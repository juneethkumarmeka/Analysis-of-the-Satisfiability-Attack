module basic_500_3000_500_30_levels_2xor_5(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
xor U0 (N_0,In_444,In_371);
nand U1 (N_1,In_421,In_28);
or U2 (N_2,In_119,In_416);
xor U3 (N_3,In_32,In_443);
nor U4 (N_4,In_472,In_65);
and U5 (N_5,In_108,In_381);
and U6 (N_6,In_365,In_336);
and U7 (N_7,In_243,In_128);
and U8 (N_8,In_245,In_202);
and U9 (N_9,In_225,In_384);
and U10 (N_10,In_209,In_271);
nor U11 (N_11,In_106,In_432);
nor U12 (N_12,In_342,In_17);
nand U13 (N_13,In_259,In_315);
nor U14 (N_14,In_356,In_36);
nor U15 (N_15,In_194,In_40);
nand U16 (N_16,In_210,In_131);
nor U17 (N_17,In_10,In_99);
xor U18 (N_18,In_41,In_0);
and U19 (N_19,In_425,In_364);
or U20 (N_20,In_164,In_470);
and U21 (N_21,In_155,In_413);
or U22 (N_22,In_308,In_35);
or U23 (N_23,In_262,In_476);
nand U24 (N_24,In_456,In_319);
xor U25 (N_25,In_335,In_58);
xnor U26 (N_26,In_217,In_494);
and U27 (N_27,In_448,In_226);
and U28 (N_28,In_45,In_96);
xnor U29 (N_29,In_81,In_244);
and U30 (N_30,In_311,In_348);
and U31 (N_31,In_485,In_94);
or U32 (N_32,In_213,In_265);
or U33 (N_33,In_475,In_269);
and U34 (N_34,In_250,In_79);
nand U35 (N_35,In_437,In_409);
xnor U36 (N_36,In_140,In_301);
nand U37 (N_37,In_25,In_346);
nor U38 (N_38,In_465,In_331);
or U39 (N_39,In_145,In_379);
nand U40 (N_40,In_439,In_26);
nor U41 (N_41,In_82,In_297);
and U42 (N_42,In_389,In_481);
and U43 (N_43,In_203,In_383);
nand U44 (N_44,In_426,In_350);
nand U45 (N_45,In_43,In_263);
nor U46 (N_46,In_102,In_248);
nand U47 (N_47,In_224,In_173);
or U48 (N_48,In_231,In_400);
xor U49 (N_49,In_423,In_33);
and U50 (N_50,In_325,In_159);
or U51 (N_51,In_281,In_30);
nor U52 (N_52,In_270,In_175);
or U53 (N_53,In_237,In_77);
and U54 (N_54,In_126,In_401);
nor U55 (N_55,In_184,In_382);
or U56 (N_56,In_487,In_132);
and U57 (N_57,In_406,In_199);
nor U58 (N_58,In_257,In_144);
nand U59 (N_59,In_85,In_332);
and U60 (N_60,In_302,In_307);
and U61 (N_61,In_14,In_362);
nor U62 (N_62,In_482,In_296);
nand U63 (N_63,In_341,In_488);
and U64 (N_64,In_172,In_97);
nand U65 (N_65,In_284,In_115);
and U66 (N_66,In_227,In_460);
and U67 (N_67,In_431,In_404);
nor U68 (N_68,In_135,In_64);
nor U69 (N_69,In_489,In_334);
or U70 (N_70,In_433,In_374);
nor U71 (N_71,In_240,In_390);
nor U72 (N_72,In_116,In_189);
nand U73 (N_73,In_181,In_451);
and U74 (N_74,In_57,In_235);
and U75 (N_75,In_300,In_124);
or U76 (N_76,In_376,In_318);
or U77 (N_77,In_282,In_415);
nand U78 (N_78,In_372,In_316);
or U79 (N_79,In_405,In_91);
or U80 (N_80,In_153,In_277);
or U81 (N_81,In_239,In_279);
or U82 (N_82,In_166,In_458);
nand U83 (N_83,In_18,In_130);
or U84 (N_84,In_123,In_320);
xor U85 (N_85,In_89,In_261);
and U86 (N_86,In_222,In_473);
nor U87 (N_87,In_42,In_138);
nor U88 (N_88,In_16,In_291);
xnor U89 (N_89,In_171,In_369);
nor U90 (N_90,In_177,In_399);
nor U91 (N_91,In_266,In_370);
and U92 (N_92,In_105,In_337);
nor U93 (N_93,In_353,In_107);
nor U94 (N_94,In_496,In_55);
and U95 (N_95,In_223,In_104);
nor U96 (N_96,In_326,In_75);
nor U97 (N_97,In_361,In_156);
nor U98 (N_98,In_367,In_21);
or U99 (N_99,In_148,In_366);
and U100 (N_100,In_76,In_27);
nand U101 (N_101,In_251,In_360);
nor U102 (N_102,In_146,N_7);
or U103 (N_103,In_446,In_230);
and U104 (N_104,In_59,In_67);
and U105 (N_105,N_71,N_94);
nor U106 (N_106,In_70,In_66);
nand U107 (N_107,In_354,In_414);
or U108 (N_108,N_88,In_93);
and U109 (N_109,In_391,N_56);
xor U110 (N_110,In_490,In_403);
or U111 (N_111,In_47,N_50);
and U112 (N_112,N_17,N_39);
nor U113 (N_113,In_388,In_359);
xor U114 (N_114,In_122,In_192);
nand U115 (N_115,In_260,In_62);
or U116 (N_116,N_36,In_411);
or U117 (N_117,In_228,In_436);
xnor U118 (N_118,In_178,In_258);
and U119 (N_119,In_478,In_154);
nand U120 (N_120,N_89,N_59);
nor U121 (N_121,N_69,In_363);
or U122 (N_122,In_295,In_63);
nand U123 (N_123,In_299,N_87);
nor U124 (N_124,N_95,N_77);
or U125 (N_125,N_2,In_141);
nand U126 (N_126,In_15,In_276);
or U127 (N_127,In_471,In_152);
or U128 (N_128,In_419,N_98);
nor U129 (N_129,In_6,In_101);
nor U130 (N_130,In_68,In_109);
nor U131 (N_131,In_170,In_100);
or U132 (N_132,In_408,In_110);
and U133 (N_133,In_92,In_118);
nand U134 (N_134,In_38,In_497);
or U135 (N_135,In_424,In_321);
and U136 (N_136,In_84,In_48);
nand U137 (N_137,In_305,In_358);
or U138 (N_138,In_339,In_254);
nand U139 (N_139,In_355,In_121);
and U140 (N_140,In_309,N_26);
or U141 (N_141,In_149,N_8);
nand U142 (N_142,In_103,In_134);
nor U143 (N_143,In_322,In_313);
nand U144 (N_144,In_351,In_442);
nand U145 (N_145,In_275,In_294);
and U146 (N_146,N_65,In_450);
nand U147 (N_147,In_137,In_338);
and U148 (N_148,In_69,N_84);
nand U149 (N_149,N_99,In_39);
nand U150 (N_150,In_9,N_63);
nand U151 (N_151,In_216,In_114);
nand U152 (N_152,In_441,In_11);
or U153 (N_153,In_272,In_255);
and U154 (N_154,In_385,N_93);
and U155 (N_155,In_264,N_29);
nor U156 (N_156,In_23,In_221);
or U157 (N_157,In_111,N_10);
nand U158 (N_158,In_2,In_232);
nand U159 (N_159,In_340,In_420);
nor U160 (N_160,In_479,In_392);
or U161 (N_161,N_64,In_143);
nand U162 (N_162,In_466,In_484);
nor U163 (N_163,In_375,N_41);
or U164 (N_164,N_14,In_24);
and U165 (N_165,N_1,In_380);
nand U166 (N_166,In_3,In_1);
nor U167 (N_167,N_51,In_19);
xor U168 (N_168,In_298,In_492);
nor U169 (N_169,In_280,In_310);
nor U170 (N_170,In_495,In_249);
xnor U171 (N_171,N_31,N_96);
or U172 (N_172,N_13,N_0);
and U173 (N_173,In_304,N_5);
and U174 (N_174,In_198,In_5);
nor U175 (N_175,In_352,N_86);
or U176 (N_176,In_438,N_54);
nand U177 (N_177,In_457,In_46);
and U178 (N_178,In_206,In_468);
and U179 (N_179,In_161,N_78);
nor U180 (N_180,In_428,N_38);
or U181 (N_181,In_20,In_205);
and U182 (N_182,N_53,In_31);
and U183 (N_183,In_56,N_19);
nand U184 (N_184,In_330,In_169);
nor U185 (N_185,In_157,In_396);
nand U186 (N_186,In_185,In_180);
and U187 (N_187,In_214,In_204);
and U188 (N_188,In_73,N_34);
nor U189 (N_189,In_477,In_312);
nand U190 (N_190,N_58,In_219);
and U191 (N_191,N_81,In_412);
nor U192 (N_192,N_20,In_434);
or U193 (N_193,In_174,In_187);
nand U194 (N_194,In_191,In_193);
nor U195 (N_195,In_133,In_86);
or U196 (N_196,In_273,In_329);
nand U197 (N_197,In_8,N_74);
or U198 (N_198,In_147,In_34);
and U199 (N_199,In_306,N_91);
or U200 (N_200,N_191,N_185);
or U201 (N_201,N_79,N_160);
nand U202 (N_202,In_333,N_72);
and U203 (N_203,In_186,In_234);
xnor U204 (N_204,In_182,N_134);
nor U205 (N_205,N_136,In_212);
or U206 (N_206,N_120,N_198);
or U207 (N_207,In_286,N_90);
nand U208 (N_208,In_327,N_190);
or U209 (N_209,N_28,In_241);
or U210 (N_210,In_54,N_57);
or U211 (N_211,N_102,N_44);
or U212 (N_212,N_199,N_109);
nand U213 (N_213,In_357,N_131);
or U214 (N_214,N_121,In_429);
nand U215 (N_215,N_155,In_256);
and U216 (N_216,In_474,In_398);
or U217 (N_217,N_60,In_207);
or U218 (N_218,N_47,N_61);
or U219 (N_219,N_145,N_23);
nand U220 (N_220,In_289,In_378);
and U221 (N_221,In_247,N_129);
and U222 (N_222,In_449,N_110);
or U223 (N_223,N_126,In_139);
and U224 (N_224,In_387,In_453);
nand U225 (N_225,In_197,N_196);
nand U226 (N_226,In_328,In_125);
and U227 (N_227,In_499,In_462);
and U228 (N_228,In_349,In_440);
or U229 (N_229,N_142,N_113);
nand U230 (N_230,N_146,In_290);
xnor U231 (N_231,N_116,In_397);
nor U232 (N_232,In_176,N_111);
nand U233 (N_233,In_422,N_37);
and U234 (N_234,In_220,In_402);
nor U235 (N_235,In_410,N_80);
nor U236 (N_236,In_188,N_169);
nor U237 (N_237,N_173,N_85);
and U238 (N_238,N_92,N_156);
nand U239 (N_239,In_150,In_129);
nor U240 (N_240,In_88,N_106);
nor U241 (N_241,N_157,N_67);
and U242 (N_242,N_119,N_76);
nor U243 (N_243,N_151,In_236);
nor U244 (N_244,N_114,In_242);
nand U245 (N_245,N_55,N_197);
and U246 (N_246,In_195,N_4);
or U247 (N_247,In_208,In_274);
nor U248 (N_248,In_83,N_179);
or U249 (N_249,N_139,N_141);
nand U250 (N_250,N_140,In_120);
nor U251 (N_251,In_491,In_87);
and U252 (N_252,In_229,N_35);
or U253 (N_253,In_394,In_452);
nor U254 (N_254,N_101,In_377);
nor U255 (N_255,In_368,N_181);
or U256 (N_256,N_118,In_293);
nand U257 (N_257,N_25,In_12);
or U258 (N_258,In_165,N_161);
and U259 (N_259,N_194,In_22);
or U260 (N_260,N_182,N_43);
and U261 (N_261,N_83,In_435);
or U262 (N_262,In_13,N_33);
and U263 (N_263,N_178,In_151);
nor U264 (N_264,In_463,N_143);
or U265 (N_265,In_7,In_288);
and U266 (N_266,In_113,In_445);
and U267 (N_267,In_343,N_104);
nand U268 (N_268,N_112,In_246);
or U269 (N_269,In_373,In_167);
nand U270 (N_270,In_317,N_15);
nand U271 (N_271,N_138,In_112);
nand U272 (N_272,N_11,In_455);
or U273 (N_273,N_167,N_123);
nor U274 (N_274,In_51,In_37);
nor U275 (N_275,In_454,N_175);
nand U276 (N_276,N_180,N_150);
nor U277 (N_277,N_177,In_53);
and U278 (N_278,N_62,N_12);
nor U279 (N_279,N_172,N_183);
xnor U280 (N_280,N_127,N_159);
nor U281 (N_281,In_427,N_147);
and U282 (N_282,In_324,In_283);
or U283 (N_283,In_469,In_183);
nand U284 (N_284,N_18,In_196);
and U285 (N_285,In_211,N_68);
nand U286 (N_286,In_314,N_70);
nor U287 (N_287,N_184,In_344);
and U288 (N_288,In_480,In_61);
or U289 (N_289,In_72,N_108);
and U290 (N_290,N_192,In_127);
and U291 (N_291,N_193,In_323);
or U292 (N_292,In_200,N_75);
nor U293 (N_293,N_45,In_467);
and U294 (N_294,In_345,In_395);
or U295 (N_295,In_201,In_303);
nand U296 (N_296,N_165,N_162);
and U297 (N_297,In_287,N_3);
nor U298 (N_298,In_417,N_154);
nand U299 (N_299,In_267,In_71);
nor U300 (N_300,N_263,N_277);
and U301 (N_301,In_78,N_253);
nand U302 (N_302,In_90,In_117);
xor U303 (N_303,N_189,N_117);
or U304 (N_304,N_166,N_187);
or U305 (N_305,N_9,In_98);
or U306 (N_306,N_278,N_30);
nand U307 (N_307,N_220,N_255);
and U308 (N_308,N_288,N_211);
nor U309 (N_309,N_296,N_271);
nand U310 (N_310,N_262,N_52);
or U311 (N_311,In_285,N_208);
or U312 (N_312,N_240,N_188);
and U313 (N_313,In_493,In_162);
and U314 (N_314,N_46,N_283);
nand U315 (N_315,N_248,N_239);
or U316 (N_316,N_276,N_207);
nand U317 (N_317,N_237,In_160);
or U318 (N_318,N_254,N_170);
and U319 (N_319,N_227,In_253);
nor U320 (N_320,N_32,N_265);
and U321 (N_321,In_461,N_176);
and U322 (N_322,In_60,N_242);
and U323 (N_323,In_407,N_256);
and U324 (N_324,N_218,N_215);
and U325 (N_325,N_292,In_464);
nand U326 (N_326,N_234,In_347);
nor U327 (N_327,N_246,N_195);
and U328 (N_328,N_209,N_201);
or U329 (N_329,N_124,N_163);
nand U330 (N_330,N_225,N_290);
and U331 (N_331,N_40,In_158);
nand U332 (N_332,N_73,In_50);
or U333 (N_333,N_249,In_393);
nand U334 (N_334,N_295,In_44);
or U335 (N_335,N_243,N_133);
nand U336 (N_336,N_200,N_149);
or U337 (N_337,N_232,N_284);
nand U338 (N_338,N_164,In_447);
or U339 (N_339,N_274,N_270);
nand U340 (N_340,N_144,In_430);
nand U341 (N_341,In_136,In_218);
and U342 (N_342,N_299,N_217);
xnor U343 (N_343,N_297,In_29);
and U344 (N_344,In_74,N_6);
nor U345 (N_345,In_179,N_272);
nand U346 (N_346,N_226,N_260);
nor U347 (N_347,N_257,In_52);
nand U348 (N_348,In_95,N_21);
and U349 (N_349,N_137,N_168);
nor U350 (N_350,N_230,In_168);
nor U351 (N_351,In_238,In_386);
or U352 (N_352,N_280,N_210);
nand U353 (N_353,N_231,N_266);
nand U354 (N_354,N_158,N_213);
or U355 (N_355,In_278,N_281);
xor U356 (N_356,N_252,N_174);
nor U357 (N_357,N_103,N_122);
or U358 (N_358,N_287,N_16);
and U359 (N_359,N_273,N_259);
nand U360 (N_360,N_238,In_268);
or U361 (N_361,N_269,N_42);
and U362 (N_362,N_152,N_275);
and U363 (N_363,N_268,N_245);
and U364 (N_364,N_148,N_219);
nand U365 (N_365,N_49,N_97);
and U366 (N_366,N_130,In_215);
or U367 (N_367,N_203,N_214);
and U368 (N_368,In_142,N_285);
xnor U369 (N_369,N_244,N_224);
nor U370 (N_370,N_298,N_229);
nand U371 (N_371,N_186,In_418);
or U372 (N_372,N_286,N_291);
nor U373 (N_373,N_212,N_202);
xnor U374 (N_374,N_258,N_132);
nor U375 (N_375,N_135,N_228);
and U376 (N_376,In_459,N_66);
and U377 (N_377,N_241,N_22);
nor U378 (N_378,N_205,N_221);
nor U379 (N_379,N_206,N_27);
or U380 (N_380,N_100,N_223);
nor U381 (N_381,N_216,N_267);
nor U382 (N_382,In_190,N_261);
and U383 (N_383,In_252,N_264);
nand U384 (N_384,In_483,N_233);
nand U385 (N_385,N_236,N_235);
nand U386 (N_386,In_163,N_105);
and U387 (N_387,N_82,N_153);
or U388 (N_388,N_222,In_498);
nor U389 (N_389,N_107,In_486);
nand U390 (N_390,N_282,N_293);
nand U391 (N_391,In_292,N_250);
nand U392 (N_392,N_204,N_294);
nand U393 (N_393,N_251,N_279);
or U394 (N_394,N_171,N_125);
or U395 (N_395,N_48,In_4);
or U396 (N_396,In_80,N_289);
nand U397 (N_397,In_49,N_128);
or U398 (N_398,N_24,N_247);
and U399 (N_399,N_115,In_233);
nor U400 (N_400,N_378,N_336);
or U401 (N_401,N_313,N_371);
or U402 (N_402,N_315,N_388);
and U403 (N_403,N_334,N_398);
nand U404 (N_404,N_357,N_306);
and U405 (N_405,N_320,N_351);
and U406 (N_406,N_300,N_356);
and U407 (N_407,N_366,N_358);
or U408 (N_408,N_399,N_374);
and U409 (N_409,N_391,N_364);
nor U410 (N_410,N_317,N_305);
and U411 (N_411,N_335,N_372);
or U412 (N_412,N_355,N_377);
nor U413 (N_413,N_344,N_393);
and U414 (N_414,N_381,N_376);
nor U415 (N_415,N_307,N_354);
nand U416 (N_416,N_311,N_360);
nor U417 (N_417,N_312,N_383);
nand U418 (N_418,N_314,N_387);
or U419 (N_419,N_353,N_369);
nor U420 (N_420,N_389,N_340);
nand U421 (N_421,N_392,N_390);
and U422 (N_422,N_347,N_341);
nand U423 (N_423,N_328,N_380);
nand U424 (N_424,N_316,N_304);
and U425 (N_425,N_321,N_396);
or U426 (N_426,N_342,N_302);
and U427 (N_427,N_384,N_329);
or U428 (N_428,N_325,N_385);
nand U429 (N_429,N_308,N_332);
nand U430 (N_430,N_368,N_324);
and U431 (N_431,N_370,N_322);
nand U432 (N_432,N_309,N_375);
nor U433 (N_433,N_337,N_339);
and U434 (N_434,N_359,N_386);
nand U435 (N_435,N_352,N_382);
nand U436 (N_436,N_379,N_365);
nand U437 (N_437,N_350,N_345);
or U438 (N_438,N_349,N_397);
or U439 (N_439,N_367,N_326);
or U440 (N_440,N_394,N_361);
nand U441 (N_441,N_318,N_303);
or U442 (N_442,N_301,N_333);
nand U443 (N_443,N_331,N_330);
and U444 (N_444,N_395,N_348);
and U445 (N_445,N_363,N_373);
and U446 (N_446,N_319,N_323);
or U447 (N_447,N_343,N_346);
or U448 (N_448,N_362,N_338);
and U449 (N_449,N_327,N_310);
nor U450 (N_450,N_342,N_365);
or U451 (N_451,N_358,N_359);
nand U452 (N_452,N_367,N_396);
nand U453 (N_453,N_395,N_343);
xnor U454 (N_454,N_340,N_375);
nor U455 (N_455,N_348,N_353);
nand U456 (N_456,N_306,N_324);
nand U457 (N_457,N_349,N_327);
nor U458 (N_458,N_336,N_374);
nor U459 (N_459,N_384,N_317);
and U460 (N_460,N_342,N_376);
or U461 (N_461,N_372,N_344);
and U462 (N_462,N_346,N_310);
nand U463 (N_463,N_367,N_378);
and U464 (N_464,N_397,N_310);
or U465 (N_465,N_316,N_326);
nor U466 (N_466,N_327,N_332);
and U467 (N_467,N_341,N_352);
nor U468 (N_468,N_315,N_375);
nor U469 (N_469,N_355,N_394);
and U470 (N_470,N_366,N_349);
nand U471 (N_471,N_336,N_300);
nor U472 (N_472,N_351,N_312);
or U473 (N_473,N_376,N_399);
nor U474 (N_474,N_394,N_353);
or U475 (N_475,N_384,N_349);
and U476 (N_476,N_365,N_362);
nand U477 (N_477,N_367,N_310);
and U478 (N_478,N_364,N_315);
nand U479 (N_479,N_375,N_310);
nor U480 (N_480,N_366,N_333);
and U481 (N_481,N_315,N_335);
or U482 (N_482,N_353,N_336);
nand U483 (N_483,N_351,N_397);
nand U484 (N_484,N_316,N_391);
xor U485 (N_485,N_368,N_392);
nor U486 (N_486,N_385,N_348);
nand U487 (N_487,N_309,N_316);
and U488 (N_488,N_316,N_300);
nor U489 (N_489,N_396,N_310);
and U490 (N_490,N_324,N_362);
or U491 (N_491,N_358,N_311);
nor U492 (N_492,N_393,N_352);
nor U493 (N_493,N_348,N_320);
nor U494 (N_494,N_383,N_359);
or U495 (N_495,N_358,N_341);
nand U496 (N_496,N_329,N_346);
nand U497 (N_497,N_359,N_353);
or U498 (N_498,N_367,N_353);
nor U499 (N_499,N_370,N_343);
nand U500 (N_500,N_473,N_422);
and U501 (N_501,N_452,N_418);
and U502 (N_502,N_429,N_407);
or U503 (N_503,N_483,N_404);
or U504 (N_504,N_431,N_403);
or U505 (N_505,N_497,N_457);
nor U506 (N_506,N_441,N_426);
and U507 (N_507,N_481,N_444);
or U508 (N_508,N_449,N_456);
nand U509 (N_509,N_458,N_450);
nand U510 (N_510,N_492,N_425);
and U511 (N_511,N_437,N_416);
or U512 (N_512,N_489,N_475);
or U513 (N_513,N_445,N_474);
nor U514 (N_514,N_484,N_411);
xnor U515 (N_515,N_463,N_482);
or U516 (N_516,N_442,N_499);
nor U517 (N_517,N_402,N_495);
or U518 (N_518,N_435,N_464);
and U519 (N_519,N_471,N_487);
nand U520 (N_520,N_432,N_455);
or U521 (N_521,N_423,N_419);
nor U522 (N_522,N_443,N_479);
nor U523 (N_523,N_400,N_434);
and U524 (N_524,N_438,N_405);
nand U525 (N_525,N_460,N_467);
or U526 (N_526,N_412,N_451);
and U527 (N_527,N_414,N_486);
nand U528 (N_528,N_417,N_478);
nand U529 (N_529,N_491,N_447);
nor U530 (N_530,N_454,N_465);
nor U531 (N_531,N_493,N_433);
and U532 (N_532,N_490,N_427);
and U533 (N_533,N_424,N_494);
nor U534 (N_534,N_470,N_496);
nand U535 (N_535,N_476,N_462);
nand U536 (N_536,N_466,N_410);
or U537 (N_537,N_477,N_408);
nor U538 (N_538,N_440,N_406);
and U539 (N_539,N_430,N_485);
and U540 (N_540,N_436,N_420);
nor U541 (N_541,N_413,N_401);
nor U542 (N_542,N_439,N_409);
nor U543 (N_543,N_480,N_446);
or U544 (N_544,N_459,N_498);
or U545 (N_545,N_488,N_461);
nand U546 (N_546,N_468,N_472);
or U547 (N_547,N_421,N_415);
xor U548 (N_548,N_428,N_469);
nor U549 (N_549,N_448,N_453);
nand U550 (N_550,N_425,N_434);
nand U551 (N_551,N_401,N_489);
or U552 (N_552,N_437,N_455);
nand U553 (N_553,N_470,N_434);
nor U554 (N_554,N_459,N_486);
nor U555 (N_555,N_495,N_470);
nor U556 (N_556,N_499,N_492);
nand U557 (N_557,N_402,N_416);
nor U558 (N_558,N_418,N_408);
nor U559 (N_559,N_474,N_473);
nand U560 (N_560,N_457,N_435);
and U561 (N_561,N_421,N_431);
or U562 (N_562,N_493,N_483);
and U563 (N_563,N_403,N_462);
nand U564 (N_564,N_440,N_479);
or U565 (N_565,N_442,N_487);
nor U566 (N_566,N_444,N_438);
or U567 (N_567,N_490,N_491);
nor U568 (N_568,N_441,N_493);
nand U569 (N_569,N_432,N_494);
or U570 (N_570,N_488,N_458);
nor U571 (N_571,N_406,N_401);
and U572 (N_572,N_499,N_410);
or U573 (N_573,N_445,N_424);
and U574 (N_574,N_468,N_441);
nor U575 (N_575,N_418,N_421);
nand U576 (N_576,N_498,N_417);
and U577 (N_577,N_453,N_401);
or U578 (N_578,N_479,N_483);
or U579 (N_579,N_474,N_487);
nand U580 (N_580,N_438,N_470);
and U581 (N_581,N_423,N_411);
xor U582 (N_582,N_444,N_418);
or U583 (N_583,N_442,N_469);
or U584 (N_584,N_460,N_478);
or U585 (N_585,N_415,N_476);
nand U586 (N_586,N_468,N_417);
nand U587 (N_587,N_498,N_490);
nand U588 (N_588,N_464,N_493);
or U589 (N_589,N_404,N_493);
and U590 (N_590,N_462,N_470);
nand U591 (N_591,N_493,N_411);
and U592 (N_592,N_414,N_427);
nor U593 (N_593,N_454,N_475);
nand U594 (N_594,N_415,N_414);
and U595 (N_595,N_445,N_459);
nor U596 (N_596,N_493,N_412);
or U597 (N_597,N_410,N_486);
and U598 (N_598,N_454,N_477);
nor U599 (N_599,N_421,N_476);
and U600 (N_600,N_531,N_526);
nor U601 (N_601,N_530,N_569);
or U602 (N_602,N_573,N_537);
nand U603 (N_603,N_556,N_585);
or U604 (N_604,N_591,N_561);
nand U605 (N_605,N_576,N_563);
and U606 (N_606,N_541,N_558);
and U607 (N_607,N_599,N_553);
nand U608 (N_608,N_583,N_567);
nand U609 (N_609,N_518,N_564);
or U610 (N_610,N_507,N_505);
and U611 (N_611,N_519,N_516);
nor U612 (N_612,N_543,N_596);
nand U613 (N_613,N_509,N_581);
nand U614 (N_614,N_506,N_560);
and U615 (N_615,N_522,N_588);
nand U616 (N_616,N_540,N_590);
and U617 (N_617,N_595,N_546);
and U618 (N_618,N_555,N_535);
and U619 (N_619,N_538,N_578);
nand U620 (N_620,N_548,N_598);
or U621 (N_621,N_554,N_597);
nor U622 (N_622,N_570,N_525);
nor U623 (N_623,N_515,N_568);
or U624 (N_624,N_508,N_529);
nor U625 (N_625,N_593,N_547);
or U626 (N_626,N_587,N_542);
nor U627 (N_627,N_503,N_521);
nor U628 (N_628,N_580,N_539);
nand U629 (N_629,N_557,N_594);
nand U630 (N_630,N_552,N_500);
and U631 (N_631,N_512,N_528);
or U632 (N_632,N_575,N_504);
nand U633 (N_633,N_545,N_524);
or U634 (N_634,N_533,N_502);
xor U635 (N_635,N_589,N_582);
nand U636 (N_636,N_513,N_571);
xor U637 (N_637,N_579,N_550);
nor U638 (N_638,N_501,N_551);
nor U639 (N_639,N_584,N_559);
and U640 (N_640,N_562,N_577);
and U641 (N_641,N_572,N_523);
and U642 (N_642,N_527,N_549);
nor U643 (N_643,N_592,N_565);
nor U644 (N_644,N_544,N_532);
nand U645 (N_645,N_510,N_534);
nor U646 (N_646,N_520,N_566);
or U647 (N_647,N_514,N_517);
or U648 (N_648,N_586,N_536);
nor U649 (N_649,N_511,N_574);
and U650 (N_650,N_572,N_569);
nor U651 (N_651,N_546,N_522);
nor U652 (N_652,N_524,N_528);
or U653 (N_653,N_528,N_544);
and U654 (N_654,N_585,N_590);
nand U655 (N_655,N_561,N_534);
nor U656 (N_656,N_548,N_572);
nor U657 (N_657,N_570,N_522);
and U658 (N_658,N_528,N_530);
and U659 (N_659,N_534,N_513);
and U660 (N_660,N_514,N_563);
or U661 (N_661,N_568,N_500);
and U662 (N_662,N_557,N_526);
and U663 (N_663,N_516,N_561);
and U664 (N_664,N_578,N_540);
nor U665 (N_665,N_583,N_520);
and U666 (N_666,N_559,N_570);
nand U667 (N_667,N_536,N_511);
or U668 (N_668,N_564,N_584);
nor U669 (N_669,N_583,N_516);
nor U670 (N_670,N_511,N_507);
and U671 (N_671,N_597,N_511);
or U672 (N_672,N_581,N_537);
nand U673 (N_673,N_577,N_594);
nand U674 (N_674,N_527,N_599);
nand U675 (N_675,N_522,N_535);
and U676 (N_676,N_590,N_577);
and U677 (N_677,N_518,N_506);
or U678 (N_678,N_504,N_582);
or U679 (N_679,N_567,N_546);
and U680 (N_680,N_585,N_543);
nor U681 (N_681,N_534,N_527);
nor U682 (N_682,N_551,N_533);
and U683 (N_683,N_505,N_510);
or U684 (N_684,N_537,N_565);
nand U685 (N_685,N_575,N_528);
nor U686 (N_686,N_578,N_586);
nand U687 (N_687,N_511,N_504);
or U688 (N_688,N_596,N_574);
or U689 (N_689,N_557,N_540);
or U690 (N_690,N_571,N_511);
nand U691 (N_691,N_593,N_560);
nor U692 (N_692,N_598,N_503);
or U693 (N_693,N_588,N_500);
or U694 (N_694,N_531,N_507);
nand U695 (N_695,N_501,N_546);
and U696 (N_696,N_544,N_561);
nand U697 (N_697,N_551,N_537);
and U698 (N_698,N_593,N_514);
and U699 (N_699,N_529,N_554);
nor U700 (N_700,N_647,N_698);
and U701 (N_701,N_626,N_650);
or U702 (N_702,N_695,N_656);
or U703 (N_703,N_651,N_690);
or U704 (N_704,N_693,N_616);
nand U705 (N_705,N_604,N_667);
nand U706 (N_706,N_654,N_648);
nor U707 (N_707,N_637,N_697);
nand U708 (N_708,N_605,N_631);
and U709 (N_709,N_611,N_630);
nand U710 (N_710,N_658,N_681);
or U711 (N_711,N_673,N_699);
and U712 (N_712,N_622,N_664);
nand U713 (N_713,N_680,N_640);
and U714 (N_714,N_612,N_666);
and U715 (N_715,N_682,N_691);
nand U716 (N_716,N_619,N_643);
nor U717 (N_717,N_607,N_657);
and U718 (N_718,N_603,N_638);
nand U719 (N_719,N_668,N_634);
nor U720 (N_720,N_674,N_602);
nor U721 (N_721,N_684,N_625);
or U722 (N_722,N_614,N_613);
nand U723 (N_723,N_610,N_679);
nor U724 (N_724,N_665,N_628);
nor U725 (N_725,N_689,N_677);
or U726 (N_726,N_688,N_669);
nor U727 (N_727,N_617,N_672);
or U728 (N_728,N_676,N_683);
nand U729 (N_729,N_636,N_608);
or U730 (N_730,N_641,N_615);
and U731 (N_731,N_633,N_671);
or U732 (N_732,N_670,N_601);
nand U733 (N_733,N_696,N_632);
nor U734 (N_734,N_675,N_663);
nor U735 (N_735,N_655,N_621);
nor U736 (N_736,N_661,N_686);
or U737 (N_737,N_646,N_649);
nor U738 (N_738,N_623,N_678);
or U739 (N_739,N_627,N_624);
and U740 (N_740,N_606,N_659);
nand U741 (N_741,N_629,N_685);
or U742 (N_742,N_662,N_652);
nor U743 (N_743,N_600,N_620);
nor U744 (N_744,N_644,N_653);
or U745 (N_745,N_642,N_694);
or U746 (N_746,N_639,N_609);
and U747 (N_747,N_660,N_618);
or U748 (N_748,N_635,N_645);
nand U749 (N_749,N_687,N_692);
or U750 (N_750,N_678,N_696);
nor U751 (N_751,N_640,N_666);
nor U752 (N_752,N_661,N_665);
nor U753 (N_753,N_695,N_672);
and U754 (N_754,N_689,N_643);
or U755 (N_755,N_665,N_681);
or U756 (N_756,N_620,N_650);
and U757 (N_757,N_630,N_682);
and U758 (N_758,N_618,N_657);
nand U759 (N_759,N_611,N_614);
nand U760 (N_760,N_672,N_658);
or U761 (N_761,N_659,N_629);
and U762 (N_762,N_691,N_609);
nand U763 (N_763,N_624,N_648);
nor U764 (N_764,N_627,N_655);
and U765 (N_765,N_620,N_601);
or U766 (N_766,N_694,N_672);
nor U767 (N_767,N_667,N_639);
and U768 (N_768,N_601,N_605);
and U769 (N_769,N_669,N_678);
nor U770 (N_770,N_630,N_681);
or U771 (N_771,N_690,N_648);
nor U772 (N_772,N_697,N_676);
nor U773 (N_773,N_627,N_679);
or U774 (N_774,N_612,N_699);
nand U775 (N_775,N_632,N_606);
and U776 (N_776,N_698,N_614);
nor U777 (N_777,N_603,N_667);
nor U778 (N_778,N_644,N_630);
and U779 (N_779,N_634,N_675);
and U780 (N_780,N_688,N_664);
and U781 (N_781,N_627,N_694);
nor U782 (N_782,N_635,N_656);
or U783 (N_783,N_629,N_636);
or U784 (N_784,N_645,N_646);
nand U785 (N_785,N_662,N_615);
nand U786 (N_786,N_684,N_616);
nand U787 (N_787,N_604,N_612);
and U788 (N_788,N_684,N_643);
nor U789 (N_789,N_655,N_693);
and U790 (N_790,N_628,N_634);
or U791 (N_791,N_630,N_668);
nand U792 (N_792,N_647,N_652);
nand U793 (N_793,N_698,N_644);
nor U794 (N_794,N_616,N_631);
or U795 (N_795,N_602,N_613);
xor U796 (N_796,N_630,N_656);
nor U797 (N_797,N_600,N_634);
and U798 (N_798,N_653,N_680);
or U799 (N_799,N_680,N_612);
nor U800 (N_800,N_734,N_713);
nor U801 (N_801,N_721,N_793);
nor U802 (N_802,N_710,N_707);
and U803 (N_803,N_760,N_757);
nand U804 (N_804,N_790,N_765);
nand U805 (N_805,N_738,N_763);
and U806 (N_806,N_798,N_762);
nor U807 (N_807,N_769,N_764);
or U808 (N_808,N_792,N_709);
nor U809 (N_809,N_786,N_720);
and U810 (N_810,N_719,N_728);
nor U811 (N_811,N_768,N_702);
nand U812 (N_812,N_741,N_736);
and U813 (N_813,N_782,N_784);
or U814 (N_814,N_799,N_725);
and U815 (N_815,N_774,N_773);
nor U816 (N_816,N_788,N_777);
nand U817 (N_817,N_732,N_703);
nor U818 (N_818,N_704,N_789);
or U819 (N_819,N_750,N_733);
or U820 (N_820,N_701,N_742);
and U821 (N_821,N_715,N_727);
or U822 (N_822,N_770,N_746);
and U823 (N_823,N_717,N_753);
nand U824 (N_824,N_795,N_708);
nor U825 (N_825,N_780,N_781);
nor U826 (N_826,N_722,N_754);
xnor U827 (N_827,N_747,N_714);
or U828 (N_828,N_723,N_752);
or U829 (N_829,N_794,N_759);
nand U830 (N_830,N_737,N_743);
nor U831 (N_831,N_772,N_756);
nand U832 (N_832,N_740,N_726);
nand U833 (N_833,N_700,N_779);
or U834 (N_834,N_745,N_724);
nor U835 (N_835,N_791,N_718);
and U836 (N_836,N_729,N_771);
nand U837 (N_837,N_730,N_749);
nor U838 (N_838,N_748,N_716);
nor U839 (N_839,N_711,N_775);
nand U840 (N_840,N_735,N_755);
or U841 (N_841,N_731,N_767);
or U842 (N_842,N_751,N_758);
xnor U843 (N_843,N_787,N_761);
nor U844 (N_844,N_744,N_796);
and U845 (N_845,N_797,N_706);
nand U846 (N_846,N_776,N_739);
and U847 (N_847,N_778,N_783);
nor U848 (N_848,N_712,N_705);
or U849 (N_849,N_785,N_766);
nor U850 (N_850,N_700,N_731);
or U851 (N_851,N_747,N_741);
or U852 (N_852,N_714,N_713);
nand U853 (N_853,N_762,N_723);
and U854 (N_854,N_763,N_724);
nand U855 (N_855,N_776,N_713);
and U856 (N_856,N_701,N_769);
nand U857 (N_857,N_787,N_769);
and U858 (N_858,N_715,N_710);
nor U859 (N_859,N_727,N_740);
nand U860 (N_860,N_701,N_775);
and U861 (N_861,N_776,N_721);
nand U862 (N_862,N_776,N_735);
nor U863 (N_863,N_749,N_707);
nor U864 (N_864,N_704,N_710);
and U865 (N_865,N_773,N_770);
or U866 (N_866,N_787,N_786);
and U867 (N_867,N_723,N_794);
nor U868 (N_868,N_797,N_703);
nand U869 (N_869,N_751,N_773);
and U870 (N_870,N_707,N_730);
or U871 (N_871,N_724,N_712);
nand U872 (N_872,N_794,N_790);
nor U873 (N_873,N_728,N_770);
nand U874 (N_874,N_781,N_797);
or U875 (N_875,N_731,N_781);
nand U876 (N_876,N_780,N_785);
nor U877 (N_877,N_721,N_777);
nand U878 (N_878,N_764,N_793);
and U879 (N_879,N_769,N_795);
nand U880 (N_880,N_767,N_751);
nand U881 (N_881,N_778,N_726);
nand U882 (N_882,N_766,N_700);
nand U883 (N_883,N_786,N_741);
and U884 (N_884,N_719,N_755);
nor U885 (N_885,N_721,N_772);
or U886 (N_886,N_768,N_761);
xor U887 (N_887,N_776,N_737);
or U888 (N_888,N_750,N_780);
nand U889 (N_889,N_795,N_725);
or U890 (N_890,N_711,N_781);
and U891 (N_891,N_718,N_729);
nor U892 (N_892,N_726,N_786);
nor U893 (N_893,N_790,N_702);
nor U894 (N_894,N_752,N_760);
nor U895 (N_895,N_769,N_731);
nor U896 (N_896,N_790,N_766);
and U897 (N_897,N_721,N_797);
nor U898 (N_898,N_733,N_714);
nor U899 (N_899,N_769,N_714);
nand U900 (N_900,N_862,N_883);
nand U901 (N_901,N_877,N_895);
or U902 (N_902,N_889,N_894);
nand U903 (N_903,N_863,N_874);
nand U904 (N_904,N_825,N_898);
and U905 (N_905,N_804,N_851);
nand U906 (N_906,N_814,N_872);
and U907 (N_907,N_846,N_890);
and U908 (N_908,N_831,N_840);
nor U909 (N_909,N_858,N_864);
nor U910 (N_910,N_822,N_870);
nor U911 (N_911,N_879,N_838);
nand U912 (N_912,N_891,N_866);
nand U913 (N_913,N_860,N_884);
or U914 (N_914,N_881,N_811);
nand U915 (N_915,N_869,N_813);
or U916 (N_916,N_844,N_893);
xnor U917 (N_917,N_803,N_865);
nand U918 (N_918,N_809,N_815);
and U919 (N_919,N_880,N_818);
nor U920 (N_920,N_807,N_854);
nand U921 (N_921,N_816,N_852);
and U922 (N_922,N_821,N_829);
nand U923 (N_923,N_849,N_859);
nand U924 (N_924,N_817,N_819);
nand U925 (N_925,N_806,N_896);
nand U926 (N_926,N_832,N_820);
or U927 (N_927,N_843,N_878);
and U928 (N_928,N_856,N_845);
nand U929 (N_929,N_830,N_828);
and U930 (N_930,N_861,N_801);
or U931 (N_931,N_823,N_808);
and U932 (N_932,N_853,N_805);
nand U933 (N_933,N_834,N_882);
and U934 (N_934,N_836,N_824);
nor U935 (N_935,N_826,N_885);
and U936 (N_936,N_802,N_871);
or U937 (N_937,N_876,N_800);
nor U938 (N_938,N_892,N_841);
or U939 (N_939,N_810,N_848);
or U940 (N_940,N_888,N_857);
and U941 (N_941,N_899,N_850);
or U942 (N_942,N_886,N_842);
or U943 (N_943,N_868,N_835);
or U944 (N_944,N_847,N_839);
nand U945 (N_945,N_887,N_812);
nor U946 (N_946,N_833,N_873);
xor U947 (N_947,N_837,N_855);
and U948 (N_948,N_875,N_827);
and U949 (N_949,N_867,N_897);
nand U950 (N_950,N_879,N_847);
xnor U951 (N_951,N_843,N_813);
and U952 (N_952,N_818,N_853);
nor U953 (N_953,N_803,N_813);
and U954 (N_954,N_891,N_884);
nand U955 (N_955,N_884,N_899);
and U956 (N_956,N_803,N_826);
nand U957 (N_957,N_875,N_888);
and U958 (N_958,N_819,N_831);
or U959 (N_959,N_886,N_831);
and U960 (N_960,N_869,N_833);
nor U961 (N_961,N_819,N_841);
and U962 (N_962,N_872,N_844);
and U963 (N_963,N_894,N_884);
xor U964 (N_964,N_859,N_832);
nor U965 (N_965,N_853,N_879);
or U966 (N_966,N_831,N_811);
or U967 (N_967,N_803,N_897);
or U968 (N_968,N_876,N_859);
or U969 (N_969,N_837,N_832);
and U970 (N_970,N_837,N_824);
nand U971 (N_971,N_878,N_810);
and U972 (N_972,N_889,N_849);
nand U973 (N_973,N_814,N_889);
and U974 (N_974,N_863,N_876);
nor U975 (N_975,N_835,N_881);
and U976 (N_976,N_866,N_875);
or U977 (N_977,N_894,N_807);
nand U978 (N_978,N_896,N_842);
and U979 (N_979,N_880,N_801);
or U980 (N_980,N_889,N_842);
nand U981 (N_981,N_826,N_881);
and U982 (N_982,N_869,N_885);
nor U983 (N_983,N_889,N_820);
nor U984 (N_984,N_839,N_809);
and U985 (N_985,N_818,N_801);
nor U986 (N_986,N_838,N_849);
or U987 (N_987,N_872,N_875);
nand U988 (N_988,N_860,N_845);
or U989 (N_989,N_825,N_835);
nand U990 (N_990,N_877,N_889);
or U991 (N_991,N_846,N_812);
and U992 (N_992,N_891,N_846);
or U993 (N_993,N_873,N_813);
and U994 (N_994,N_855,N_814);
and U995 (N_995,N_852,N_862);
nand U996 (N_996,N_801,N_885);
nand U997 (N_997,N_800,N_840);
nand U998 (N_998,N_848,N_826);
nand U999 (N_999,N_887,N_816);
nor U1000 (N_1000,N_987,N_941);
nor U1001 (N_1001,N_954,N_963);
and U1002 (N_1002,N_986,N_939);
or U1003 (N_1003,N_989,N_990);
or U1004 (N_1004,N_953,N_911);
nand U1005 (N_1005,N_956,N_983);
nor U1006 (N_1006,N_969,N_997);
or U1007 (N_1007,N_967,N_938);
or U1008 (N_1008,N_979,N_985);
and U1009 (N_1009,N_958,N_909);
and U1010 (N_1010,N_993,N_947);
nand U1011 (N_1011,N_966,N_976);
and U1012 (N_1012,N_992,N_913);
xnor U1013 (N_1013,N_931,N_935);
and U1014 (N_1014,N_934,N_906);
or U1015 (N_1015,N_927,N_903);
nand U1016 (N_1016,N_926,N_977);
nand U1017 (N_1017,N_973,N_905);
or U1018 (N_1018,N_980,N_932);
nand U1019 (N_1019,N_928,N_942);
or U1020 (N_1020,N_923,N_933);
nor U1021 (N_1021,N_916,N_944);
or U1022 (N_1022,N_924,N_920);
or U1023 (N_1023,N_975,N_970);
or U1024 (N_1024,N_918,N_945);
or U1025 (N_1025,N_991,N_937);
nor U1026 (N_1026,N_912,N_919);
nand U1027 (N_1027,N_930,N_951);
nand U1028 (N_1028,N_915,N_908);
and U1029 (N_1029,N_998,N_925);
or U1030 (N_1030,N_994,N_999);
or U1031 (N_1031,N_914,N_952);
nor U1032 (N_1032,N_972,N_971);
nand U1033 (N_1033,N_978,N_959);
or U1034 (N_1034,N_957,N_964);
or U1035 (N_1035,N_904,N_960);
or U1036 (N_1036,N_907,N_910);
or U1037 (N_1037,N_988,N_921);
or U1038 (N_1038,N_949,N_948);
nand U1039 (N_1039,N_946,N_962);
nor U1040 (N_1040,N_950,N_974);
or U1041 (N_1041,N_917,N_929);
or U1042 (N_1042,N_968,N_981);
xor U1043 (N_1043,N_922,N_900);
and U1044 (N_1044,N_902,N_936);
or U1045 (N_1045,N_995,N_965);
and U1046 (N_1046,N_901,N_955);
or U1047 (N_1047,N_943,N_982);
and U1048 (N_1048,N_940,N_996);
nor U1049 (N_1049,N_961,N_984);
nor U1050 (N_1050,N_922,N_920);
and U1051 (N_1051,N_967,N_904);
or U1052 (N_1052,N_904,N_978);
and U1053 (N_1053,N_955,N_998);
nor U1054 (N_1054,N_918,N_914);
xor U1055 (N_1055,N_905,N_948);
nand U1056 (N_1056,N_980,N_921);
and U1057 (N_1057,N_969,N_928);
and U1058 (N_1058,N_909,N_970);
and U1059 (N_1059,N_940,N_971);
nor U1060 (N_1060,N_997,N_987);
and U1061 (N_1061,N_972,N_902);
or U1062 (N_1062,N_988,N_957);
and U1063 (N_1063,N_926,N_929);
and U1064 (N_1064,N_946,N_958);
and U1065 (N_1065,N_902,N_906);
nand U1066 (N_1066,N_927,N_905);
or U1067 (N_1067,N_928,N_952);
xor U1068 (N_1068,N_909,N_955);
or U1069 (N_1069,N_906,N_965);
and U1070 (N_1070,N_993,N_992);
nand U1071 (N_1071,N_948,N_964);
and U1072 (N_1072,N_993,N_986);
nor U1073 (N_1073,N_986,N_954);
or U1074 (N_1074,N_946,N_969);
and U1075 (N_1075,N_957,N_930);
and U1076 (N_1076,N_939,N_961);
nor U1077 (N_1077,N_973,N_913);
nor U1078 (N_1078,N_912,N_955);
nor U1079 (N_1079,N_916,N_901);
and U1080 (N_1080,N_966,N_953);
nor U1081 (N_1081,N_982,N_977);
nor U1082 (N_1082,N_938,N_969);
nand U1083 (N_1083,N_931,N_972);
or U1084 (N_1084,N_934,N_998);
or U1085 (N_1085,N_929,N_910);
and U1086 (N_1086,N_945,N_935);
nor U1087 (N_1087,N_965,N_932);
nand U1088 (N_1088,N_921,N_985);
nor U1089 (N_1089,N_943,N_907);
or U1090 (N_1090,N_990,N_974);
and U1091 (N_1091,N_998,N_960);
xor U1092 (N_1092,N_972,N_941);
and U1093 (N_1093,N_948,N_908);
nor U1094 (N_1094,N_907,N_926);
nand U1095 (N_1095,N_971,N_927);
and U1096 (N_1096,N_957,N_926);
and U1097 (N_1097,N_968,N_931);
nor U1098 (N_1098,N_995,N_958);
nand U1099 (N_1099,N_982,N_933);
or U1100 (N_1100,N_1011,N_1005);
and U1101 (N_1101,N_1091,N_1079);
nor U1102 (N_1102,N_1009,N_1035);
nor U1103 (N_1103,N_1081,N_1022);
or U1104 (N_1104,N_1031,N_1095);
or U1105 (N_1105,N_1008,N_1003);
and U1106 (N_1106,N_1037,N_1020);
nand U1107 (N_1107,N_1088,N_1094);
nand U1108 (N_1108,N_1083,N_1017);
and U1109 (N_1109,N_1038,N_1047);
nand U1110 (N_1110,N_1060,N_1093);
or U1111 (N_1111,N_1065,N_1072);
or U1112 (N_1112,N_1030,N_1097);
and U1113 (N_1113,N_1080,N_1073);
nor U1114 (N_1114,N_1059,N_1069);
or U1115 (N_1115,N_1096,N_1046);
nor U1116 (N_1116,N_1034,N_1055);
or U1117 (N_1117,N_1014,N_1036);
xor U1118 (N_1118,N_1002,N_1090);
or U1119 (N_1119,N_1056,N_1012);
or U1120 (N_1120,N_1023,N_1041);
or U1121 (N_1121,N_1052,N_1067);
nand U1122 (N_1122,N_1066,N_1070);
and U1123 (N_1123,N_1010,N_1024);
nand U1124 (N_1124,N_1049,N_1075);
and U1125 (N_1125,N_1045,N_1039);
nor U1126 (N_1126,N_1015,N_1074);
nor U1127 (N_1127,N_1033,N_1044);
nand U1128 (N_1128,N_1062,N_1092);
nand U1129 (N_1129,N_1018,N_1029);
and U1130 (N_1130,N_1054,N_1042);
nor U1131 (N_1131,N_1098,N_1053);
nand U1132 (N_1132,N_1064,N_1084);
nor U1133 (N_1133,N_1087,N_1063);
and U1134 (N_1134,N_1025,N_1089);
nand U1135 (N_1135,N_1013,N_1071);
nand U1136 (N_1136,N_1027,N_1086);
nor U1137 (N_1137,N_1058,N_1019);
or U1138 (N_1138,N_1007,N_1082);
and U1139 (N_1139,N_1057,N_1068);
nand U1140 (N_1140,N_1051,N_1043);
nand U1141 (N_1141,N_1028,N_1004);
nor U1142 (N_1142,N_1050,N_1000);
and U1143 (N_1143,N_1048,N_1021);
nor U1144 (N_1144,N_1061,N_1032);
nor U1145 (N_1145,N_1077,N_1076);
or U1146 (N_1146,N_1001,N_1040);
or U1147 (N_1147,N_1026,N_1078);
nor U1148 (N_1148,N_1099,N_1016);
nor U1149 (N_1149,N_1085,N_1006);
or U1150 (N_1150,N_1079,N_1056);
nor U1151 (N_1151,N_1097,N_1073);
nor U1152 (N_1152,N_1092,N_1008);
nand U1153 (N_1153,N_1068,N_1022);
nor U1154 (N_1154,N_1021,N_1058);
nor U1155 (N_1155,N_1009,N_1071);
or U1156 (N_1156,N_1087,N_1011);
nor U1157 (N_1157,N_1029,N_1082);
and U1158 (N_1158,N_1086,N_1089);
nor U1159 (N_1159,N_1004,N_1042);
nand U1160 (N_1160,N_1080,N_1070);
nor U1161 (N_1161,N_1037,N_1083);
nor U1162 (N_1162,N_1088,N_1093);
nand U1163 (N_1163,N_1044,N_1029);
and U1164 (N_1164,N_1026,N_1017);
and U1165 (N_1165,N_1010,N_1060);
or U1166 (N_1166,N_1014,N_1040);
nand U1167 (N_1167,N_1036,N_1038);
nand U1168 (N_1168,N_1004,N_1056);
nor U1169 (N_1169,N_1043,N_1044);
and U1170 (N_1170,N_1053,N_1099);
and U1171 (N_1171,N_1076,N_1011);
or U1172 (N_1172,N_1088,N_1010);
xor U1173 (N_1173,N_1063,N_1043);
nand U1174 (N_1174,N_1048,N_1023);
nor U1175 (N_1175,N_1085,N_1007);
or U1176 (N_1176,N_1035,N_1014);
nand U1177 (N_1177,N_1002,N_1060);
nand U1178 (N_1178,N_1018,N_1031);
nand U1179 (N_1179,N_1098,N_1050);
nand U1180 (N_1180,N_1027,N_1047);
nand U1181 (N_1181,N_1065,N_1046);
and U1182 (N_1182,N_1046,N_1030);
or U1183 (N_1183,N_1062,N_1023);
and U1184 (N_1184,N_1009,N_1047);
and U1185 (N_1185,N_1014,N_1041);
nand U1186 (N_1186,N_1035,N_1038);
nor U1187 (N_1187,N_1096,N_1088);
nand U1188 (N_1188,N_1024,N_1071);
nand U1189 (N_1189,N_1049,N_1015);
and U1190 (N_1190,N_1052,N_1074);
nor U1191 (N_1191,N_1066,N_1015);
nor U1192 (N_1192,N_1071,N_1022);
nand U1193 (N_1193,N_1045,N_1014);
and U1194 (N_1194,N_1068,N_1074);
or U1195 (N_1195,N_1061,N_1029);
and U1196 (N_1196,N_1041,N_1070);
or U1197 (N_1197,N_1099,N_1003);
or U1198 (N_1198,N_1094,N_1068);
or U1199 (N_1199,N_1041,N_1080);
nor U1200 (N_1200,N_1174,N_1166);
or U1201 (N_1201,N_1147,N_1182);
nand U1202 (N_1202,N_1185,N_1191);
nand U1203 (N_1203,N_1151,N_1123);
nor U1204 (N_1204,N_1130,N_1164);
nand U1205 (N_1205,N_1179,N_1144);
nor U1206 (N_1206,N_1196,N_1171);
nor U1207 (N_1207,N_1138,N_1119);
xor U1208 (N_1208,N_1172,N_1135);
xor U1209 (N_1209,N_1107,N_1120);
or U1210 (N_1210,N_1197,N_1158);
nand U1211 (N_1211,N_1100,N_1134);
nor U1212 (N_1212,N_1188,N_1122);
or U1213 (N_1213,N_1169,N_1167);
or U1214 (N_1214,N_1110,N_1152);
or U1215 (N_1215,N_1116,N_1149);
or U1216 (N_1216,N_1163,N_1155);
and U1217 (N_1217,N_1173,N_1106);
nand U1218 (N_1218,N_1108,N_1176);
nor U1219 (N_1219,N_1192,N_1193);
or U1220 (N_1220,N_1103,N_1128);
or U1221 (N_1221,N_1181,N_1111);
xor U1222 (N_1222,N_1113,N_1170);
nand U1223 (N_1223,N_1124,N_1180);
nand U1224 (N_1224,N_1142,N_1187);
or U1225 (N_1225,N_1199,N_1194);
and U1226 (N_1226,N_1198,N_1145);
nand U1227 (N_1227,N_1125,N_1157);
nand U1228 (N_1228,N_1141,N_1162);
nor U1229 (N_1229,N_1183,N_1109);
and U1230 (N_1230,N_1190,N_1139);
or U1231 (N_1231,N_1178,N_1148);
or U1232 (N_1232,N_1156,N_1175);
nand U1233 (N_1233,N_1118,N_1126);
and U1234 (N_1234,N_1195,N_1160);
and U1235 (N_1235,N_1105,N_1153);
nor U1236 (N_1236,N_1132,N_1104);
and U1237 (N_1237,N_1186,N_1159);
and U1238 (N_1238,N_1137,N_1150);
and U1239 (N_1239,N_1154,N_1112);
or U1240 (N_1240,N_1161,N_1121);
and U1241 (N_1241,N_1165,N_1143);
nand U1242 (N_1242,N_1127,N_1136);
or U1243 (N_1243,N_1102,N_1131);
or U1244 (N_1244,N_1177,N_1133);
nand U1245 (N_1245,N_1114,N_1189);
or U1246 (N_1246,N_1184,N_1146);
or U1247 (N_1247,N_1117,N_1140);
and U1248 (N_1248,N_1129,N_1101);
nand U1249 (N_1249,N_1115,N_1168);
nand U1250 (N_1250,N_1177,N_1168);
nor U1251 (N_1251,N_1111,N_1117);
nand U1252 (N_1252,N_1126,N_1154);
nand U1253 (N_1253,N_1131,N_1111);
or U1254 (N_1254,N_1102,N_1190);
or U1255 (N_1255,N_1162,N_1154);
or U1256 (N_1256,N_1162,N_1114);
xnor U1257 (N_1257,N_1104,N_1108);
and U1258 (N_1258,N_1102,N_1149);
nand U1259 (N_1259,N_1163,N_1196);
nor U1260 (N_1260,N_1106,N_1160);
and U1261 (N_1261,N_1100,N_1187);
and U1262 (N_1262,N_1136,N_1109);
and U1263 (N_1263,N_1192,N_1143);
nand U1264 (N_1264,N_1196,N_1152);
or U1265 (N_1265,N_1119,N_1133);
nor U1266 (N_1266,N_1165,N_1185);
or U1267 (N_1267,N_1101,N_1105);
nor U1268 (N_1268,N_1163,N_1167);
and U1269 (N_1269,N_1187,N_1197);
nand U1270 (N_1270,N_1112,N_1191);
nor U1271 (N_1271,N_1117,N_1138);
nor U1272 (N_1272,N_1197,N_1156);
nand U1273 (N_1273,N_1171,N_1189);
and U1274 (N_1274,N_1167,N_1106);
and U1275 (N_1275,N_1143,N_1181);
and U1276 (N_1276,N_1146,N_1121);
nor U1277 (N_1277,N_1127,N_1171);
nand U1278 (N_1278,N_1180,N_1117);
nor U1279 (N_1279,N_1186,N_1198);
nor U1280 (N_1280,N_1146,N_1172);
or U1281 (N_1281,N_1142,N_1145);
or U1282 (N_1282,N_1167,N_1135);
nor U1283 (N_1283,N_1167,N_1125);
and U1284 (N_1284,N_1172,N_1152);
and U1285 (N_1285,N_1131,N_1141);
and U1286 (N_1286,N_1189,N_1198);
or U1287 (N_1287,N_1156,N_1109);
and U1288 (N_1288,N_1132,N_1119);
and U1289 (N_1289,N_1110,N_1191);
or U1290 (N_1290,N_1161,N_1122);
nand U1291 (N_1291,N_1101,N_1188);
and U1292 (N_1292,N_1172,N_1120);
xor U1293 (N_1293,N_1103,N_1118);
nor U1294 (N_1294,N_1169,N_1196);
or U1295 (N_1295,N_1123,N_1162);
nor U1296 (N_1296,N_1144,N_1154);
nor U1297 (N_1297,N_1181,N_1167);
nor U1298 (N_1298,N_1113,N_1145);
nor U1299 (N_1299,N_1130,N_1182);
nand U1300 (N_1300,N_1219,N_1231);
nand U1301 (N_1301,N_1216,N_1242);
or U1302 (N_1302,N_1209,N_1253);
or U1303 (N_1303,N_1266,N_1288);
and U1304 (N_1304,N_1261,N_1295);
nand U1305 (N_1305,N_1211,N_1267);
or U1306 (N_1306,N_1228,N_1260);
or U1307 (N_1307,N_1264,N_1286);
and U1308 (N_1308,N_1278,N_1238);
or U1309 (N_1309,N_1294,N_1291);
or U1310 (N_1310,N_1239,N_1262);
and U1311 (N_1311,N_1272,N_1217);
nor U1312 (N_1312,N_1281,N_1230);
nand U1313 (N_1313,N_1229,N_1221);
and U1314 (N_1314,N_1240,N_1273);
nor U1315 (N_1315,N_1279,N_1223);
and U1316 (N_1316,N_1287,N_1250);
nor U1317 (N_1317,N_1232,N_1249);
or U1318 (N_1318,N_1299,N_1212);
and U1319 (N_1319,N_1297,N_1289);
nor U1320 (N_1320,N_1298,N_1244);
xnor U1321 (N_1321,N_1213,N_1247);
nor U1322 (N_1322,N_1271,N_1265);
and U1323 (N_1323,N_1224,N_1227);
or U1324 (N_1324,N_1246,N_1233);
nand U1325 (N_1325,N_1201,N_1241);
nor U1326 (N_1326,N_1280,N_1274);
nor U1327 (N_1327,N_1277,N_1226);
and U1328 (N_1328,N_1248,N_1285);
nand U1329 (N_1329,N_1270,N_1256);
and U1330 (N_1330,N_1268,N_1283);
and U1331 (N_1331,N_1235,N_1210);
nand U1332 (N_1332,N_1258,N_1252);
nand U1333 (N_1333,N_1251,N_1208);
and U1334 (N_1334,N_1214,N_1284);
or U1335 (N_1335,N_1222,N_1259);
nor U1336 (N_1336,N_1206,N_1204);
nor U1337 (N_1337,N_1263,N_1215);
nand U1338 (N_1338,N_1269,N_1207);
and U1339 (N_1339,N_1234,N_1276);
nand U1340 (N_1340,N_1200,N_1290);
and U1341 (N_1341,N_1296,N_1257);
nor U1342 (N_1342,N_1245,N_1254);
and U1343 (N_1343,N_1275,N_1292);
nor U1344 (N_1344,N_1243,N_1205);
nor U1345 (N_1345,N_1220,N_1293);
nand U1346 (N_1346,N_1218,N_1237);
nand U1347 (N_1347,N_1236,N_1255);
or U1348 (N_1348,N_1282,N_1203);
nor U1349 (N_1349,N_1225,N_1202);
nand U1350 (N_1350,N_1261,N_1266);
and U1351 (N_1351,N_1227,N_1260);
nand U1352 (N_1352,N_1213,N_1292);
nor U1353 (N_1353,N_1282,N_1236);
or U1354 (N_1354,N_1234,N_1209);
and U1355 (N_1355,N_1265,N_1275);
or U1356 (N_1356,N_1231,N_1225);
nand U1357 (N_1357,N_1297,N_1280);
and U1358 (N_1358,N_1213,N_1215);
and U1359 (N_1359,N_1265,N_1257);
and U1360 (N_1360,N_1201,N_1243);
or U1361 (N_1361,N_1201,N_1291);
nand U1362 (N_1362,N_1264,N_1267);
nand U1363 (N_1363,N_1214,N_1291);
nand U1364 (N_1364,N_1258,N_1294);
nand U1365 (N_1365,N_1283,N_1233);
nor U1366 (N_1366,N_1269,N_1228);
or U1367 (N_1367,N_1216,N_1208);
or U1368 (N_1368,N_1261,N_1204);
and U1369 (N_1369,N_1210,N_1294);
or U1370 (N_1370,N_1205,N_1207);
and U1371 (N_1371,N_1209,N_1258);
nand U1372 (N_1372,N_1283,N_1239);
or U1373 (N_1373,N_1281,N_1293);
or U1374 (N_1374,N_1265,N_1289);
or U1375 (N_1375,N_1263,N_1285);
and U1376 (N_1376,N_1250,N_1256);
or U1377 (N_1377,N_1207,N_1250);
nand U1378 (N_1378,N_1249,N_1222);
or U1379 (N_1379,N_1248,N_1216);
and U1380 (N_1380,N_1247,N_1265);
nor U1381 (N_1381,N_1226,N_1264);
and U1382 (N_1382,N_1299,N_1253);
or U1383 (N_1383,N_1288,N_1231);
xor U1384 (N_1384,N_1249,N_1272);
xor U1385 (N_1385,N_1249,N_1276);
nor U1386 (N_1386,N_1276,N_1257);
and U1387 (N_1387,N_1219,N_1264);
or U1388 (N_1388,N_1280,N_1255);
nand U1389 (N_1389,N_1252,N_1205);
nand U1390 (N_1390,N_1212,N_1271);
nor U1391 (N_1391,N_1204,N_1299);
and U1392 (N_1392,N_1251,N_1250);
nand U1393 (N_1393,N_1219,N_1290);
nor U1394 (N_1394,N_1256,N_1269);
or U1395 (N_1395,N_1277,N_1202);
nor U1396 (N_1396,N_1223,N_1244);
nor U1397 (N_1397,N_1242,N_1251);
nor U1398 (N_1398,N_1263,N_1237);
nor U1399 (N_1399,N_1210,N_1270);
or U1400 (N_1400,N_1341,N_1351);
and U1401 (N_1401,N_1353,N_1363);
or U1402 (N_1402,N_1378,N_1388);
nor U1403 (N_1403,N_1375,N_1357);
and U1404 (N_1404,N_1344,N_1311);
or U1405 (N_1405,N_1334,N_1358);
nor U1406 (N_1406,N_1315,N_1389);
nand U1407 (N_1407,N_1310,N_1301);
nor U1408 (N_1408,N_1343,N_1323);
nor U1409 (N_1409,N_1314,N_1356);
nor U1410 (N_1410,N_1345,N_1335);
nand U1411 (N_1411,N_1379,N_1396);
and U1412 (N_1412,N_1383,N_1309);
and U1413 (N_1413,N_1370,N_1304);
and U1414 (N_1414,N_1399,N_1362);
nor U1415 (N_1415,N_1376,N_1354);
or U1416 (N_1416,N_1319,N_1333);
xor U1417 (N_1417,N_1377,N_1352);
or U1418 (N_1418,N_1337,N_1386);
and U1419 (N_1419,N_1393,N_1347);
nor U1420 (N_1420,N_1366,N_1308);
and U1421 (N_1421,N_1355,N_1329);
nand U1422 (N_1422,N_1300,N_1361);
xor U1423 (N_1423,N_1385,N_1322);
and U1424 (N_1424,N_1346,N_1348);
nand U1425 (N_1425,N_1328,N_1327);
nor U1426 (N_1426,N_1374,N_1331);
and U1427 (N_1427,N_1320,N_1340);
and U1428 (N_1428,N_1338,N_1307);
xnor U1429 (N_1429,N_1342,N_1302);
nor U1430 (N_1430,N_1398,N_1321);
xnor U1431 (N_1431,N_1395,N_1369);
and U1432 (N_1432,N_1306,N_1317);
or U1433 (N_1433,N_1324,N_1360);
xor U1434 (N_1434,N_1364,N_1391);
nor U1435 (N_1435,N_1303,N_1387);
and U1436 (N_1436,N_1330,N_1313);
nand U1437 (N_1437,N_1367,N_1382);
and U1438 (N_1438,N_1397,N_1392);
nand U1439 (N_1439,N_1384,N_1312);
and U1440 (N_1440,N_1350,N_1359);
or U1441 (N_1441,N_1326,N_1394);
nand U1442 (N_1442,N_1365,N_1349);
nand U1443 (N_1443,N_1332,N_1381);
and U1444 (N_1444,N_1339,N_1368);
and U1445 (N_1445,N_1390,N_1373);
or U1446 (N_1446,N_1371,N_1305);
nand U1447 (N_1447,N_1336,N_1380);
and U1448 (N_1448,N_1325,N_1316);
or U1449 (N_1449,N_1372,N_1318);
nor U1450 (N_1450,N_1300,N_1317);
nand U1451 (N_1451,N_1370,N_1366);
nand U1452 (N_1452,N_1312,N_1346);
or U1453 (N_1453,N_1363,N_1379);
and U1454 (N_1454,N_1330,N_1355);
or U1455 (N_1455,N_1301,N_1343);
nor U1456 (N_1456,N_1330,N_1371);
nand U1457 (N_1457,N_1318,N_1378);
and U1458 (N_1458,N_1329,N_1327);
nor U1459 (N_1459,N_1379,N_1308);
and U1460 (N_1460,N_1340,N_1390);
and U1461 (N_1461,N_1355,N_1359);
nand U1462 (N_1462,N_1311,N_1372);
and U1463 (N_1463,N_1380,N_1355);
nor U1464 (N_1464,N_1320,N_1353);
xnor U1465 (N_1465,N_1378,N_1381);
xor U1466 (N_1466,N_1372,N_1317);
or U1467 (N_1467,N_1326,N_1317);
and U1468 (N_1468,N_1392,N_1381);
or U1469 (N_1469,N_1315,N_1370);
nand U1470 (N_1470,N_1362,N_1374);
nand U1471 (N_1471,N_1388,N_1337);
nor U1472 (N_1472,N_1338,N_1358);
or U1473 (N_1473,N_1364,N_1385);
nor U1474 (N_1474,N_1339,N_1347);
or U1475 (N_1475,N_1304,N_1372);
and U1476 (N_1476,N_1315,N_1393);
nor U1477 (N_1477,N_1389,N_1366);
and U1478 (N_1478,N_1365,N_1337);
or U1479 (N_1479,N_1317,N_1358);
nand U1480 (N_1480,N_1368,N_1342);
nor U1481 (N_1481,N_1363,N_1341);
nand U1482 (N_1482,N_1336,N_1393);
and U1483 (N_1483,N_1376,N_1371);
and U1484 (N_1484,N_1304,N_1353);
nor U1485 (N_1485,N_1346,N_1320);
nand U1486 (N_1486,N_1386,N_1369);
and U1487 (N_1487,N_1334,N_1316);
and U1488 (N_1488,N_1345,N_1312);
or U1489 (N_1489,N_1331,N_1394);
and U1490 (N_1490,N_1347,N_1351);
or U1491 (N_1491,N_1312,N_1300);
and U1492 (N_1492,N_1334,N_1331);
or U1493 (N_1493,N_1349,N_1321);
nor U1494 (N_1494,N_1340,N_1338);
or U1495 (N_1495,N_1330,N_1346);
and U1496 (N_1496,N_1318,N_1369);
and U1497 (N_1497,N_1379,N_1384);
or U1498 (N_1498,N_1367,N_1388);
and U1499 (N_1499,N_1348,N_1360);
nand U1500 (N_1500,N_1459,N_1417);
and U1501 (N_1501,N_1443,N_1471);
or U1502 (N_1502,N_1400,N_1439);
nor U1503 (N_1503,N_1431,N_1495);
nand U1504 (N_1504,N_1466,N_1496);
and U1505 (N_1505,N_1447,N_1424);
nand U1506 (N_1506,N_1425,N_1448);
nor U1507 (N_1507,N_1446,N_1468);
and U1508 (N_1508,N_1430,N_1408);
nand U1509 (N_1509,N_1429,N_1467);
nand U1510 (N_1510,N_1407,N_1404);
nor U1511 (N_1511,N_1416,N_1477);
or U1512 (N_1512,N_1420,N_1465);
nand U1513 (N_1513,N_1452,N_1475);
and U1514 (N_1514,N_1445,N_1489);
or U1515 (N_1515,N_1402,N_1485);
or U1516 (N_1516,N_1487,N_1497);
or U1517 (N_1517,N_1436,N_1484);
nand U1518 (N_1518,N_1491,N_1481);
or U1519 (N_1519,N_1480,N_1435);
or U1520 (N_1520,N_1478,N_1449);
or U1521 (N_1521,N_1454,N_1426);
nor U1522 (N_1522,N_1428,N_1462);
and U1523 (N_1523,N_1434,N_1464);
and U1524 (N_1524,N_1422,N_1441);
and U1525 (N_1525,N_1499,N_1418);
or U1526 (N_1526,N_1488,N_1427);
nand U1527 (N_1527,N_1461,N_1413);
and U1528 (N_1528,N_1440,N_1483);
and U1529 (N_1529,N_1410,N_1403);
and U1530 (N_1530,N_1409,N_1493);
nand U1531 (N_1531,N_1453,N_1486);
or U1532 (N_1532,N_1470,N_1401);
and U1533 (N_1533,N_1455,N_1460);
nor U1534 (N_1534,N_1494,N_1423);
xnor U1535 (N_1535,N_1444,N_1479);
nor U1536 (N_1536,N_1456,N_1412);
and U1537 (N_1537,N_1472,N_1442);
or U1538 (N_1538,N_1437,N_1406);
nor U1539 (N_1539,N_1419,N_1405);
nand U1540 (N_1540,N_1474,N_1482);
and U1541 (N_1541,N_1498,N_1411);
or U1542 (N_1542,N_1473,N_1490);
nor U1543 (N_1543,N_1438,N_1469);
nor U1544 (N_1544,N_1492,N_1421);
and U1545 (N_1545,N_1450,N_1476);
or U1546 (N_1546,N_1433,N_1458);
nand U1547 (N_1547,N_1457,N_1414);
or U1548 (N_1548,N_1451,N_1463);
nand U1549 (N_1549,N_1432,N_1415);
and U1550 (N_1550,N_1449,N_1461);
and U1551 (N_1551,N_1425,N_1492);
and U1552 (N_1552,N_1452,N_1454);
nand U1553 (N_1553,N_1404,N_1401);
xnor U1554 (N_1554,N_1463,N_1483);
and U1555 (N_1555,N_1432,N_1426);
and U1556 (N_1556,N_1436,N_1400);
nor U1557 (N_1557,N_1401,N_1454);
and U1558 (N_1558,N_1450,N_1444);
nor U1559 (N_1559,N_1497,N_1400);
nand U1560 (N_1560,N_1468,N_1463);
nor U1561 (N_1561,N_1440,N_1417);
and U1562 (N_1562,N_1417,N_1472);
or U1563 (N_1563,N_1439,N_1481);
or U1564 (N_1564,N_1430,N_1432);
nand U1565 (N_1565,N_1451,N_1468);
nand U1566 (N_1566,N_1425,N_1414);
nor U1567 (N_1567,N_1430,N_1495);
nor U1568 (N_1568,N_1402,N_1471);
nor U1569 (N_1569,N_1437,N_1410);
nor U1570 (N_1570,N_1496,N_1453);
and U1571 (N_1571,N_1402,N_1466);
and U1572 (N_1572,N_1491,N_1477);
and U1573 (N_1573,N_1475,N_1433);
or U1574 (N_1574,N_1456,N_1459);
nand U1575 (N_1575,N_1436,N_1465);
nand U1576 (N_1576,N_1471,N_1446);
nor U1577 (N_1577,N_1493,N_1401);
nand U1578 (N_1578,N_1482,N_1476);
or U1579 (N_1579,N_1454,N_1427);
or U1580 (N_1580,N_1477,N_1412);
and U1581 (N_1581,N_1414,N_1473);
and U1582 (N_1582,N_1471,N_1435);
nor U1583 (N_1583,N_1407,N_1459);
or U1584 (N_1584,N_1422,N_1455);
nor U1585 (N_1585,N_1456,N_1465);
or U1586 (N_1586,N_1467,N_1490);
nand U1587 (N_1587,N_1475,N_1435);
nand U1588 (N_1588,N_1475,N_1482);
or U1589 (N_1589,N_1417,N_1428);
and U1590 (N_1590,N_1450,N_1487);
nand U1591 (N_1591,N_1409,N_1438);
xnor U1592 (N_1592,N_1486,N_1482);
nand U1593 (N_1593,N_1463,N_1455);
nor U1594 (N_1594,N_1437,N_1429);
or U1595 (N_1595,N_1474,N_1472);
or U1596 (N_1596,N_1488,N_1448);
and U1597 (N_1597,N_1423,N_1436);
and U1598 (N_1598,N_1494,N_1449);
nand U1599 (N_1599,N_1455,N_1492);
nand U1600 (N_1600,N_1516,N_1544);
or U1601 (N_1601,N_1510,N_1537);
nand U1602 (N_1602,N_1587,N_1527);
nor U1603 (N_1603,N_1595,N_1512);
and U1604 (N_1604,N_1579,N_1528);
or U1605 (N_1605,N_1566,N_1524);
and U1606 (N_1606,N_1523,N_1597);
xnor U1607 (N_1607,N_1565,N_1571);
or U1608 (N_1608,N_1562,N_1576);
or U1609 (N_1609,N_1503,N_1506);
and U1610 (N_1610,N_1501,N_1532);
nand U1611 (N_1611,N_1531,N_1525);
and U1612 (N_1612,N_1552,N_1545);
nor U1613 (N_1613,N_1598,N_1581);
nor U1614 (N_1614,N_1583,N_1540);
nor U1615 (N_1615,N_1547,N_1550);
nand U1616 (N_1616,N_1535,N_1559);
nor U1617 (N_1617,N_1553,N_1522);
and U1618 (N_1618,N_1574,N_1538);
or U1619 (N_1619,N_1515,N_1592);
and U1620 (N_1620,N_1578,N_1548);
and U1621 (N_1621,N_1539,N_1588);
nor U1622 (N_1622,N_1584,N_1577);
or U1623 (N_1623,N_1558,N_1533);
or U1624 (N_1624,N_1502,N_1560);
or U1625 (N_1625,N_1555,N_1546);
or U1626 (N_1626,N_1580,N_1530);
nand U1627 (N_1627,N_1543,N_1549);
nor U1628 (N_1628,N_1594,N_1591);
nand U1629 (N_1629,N_1554,N_1567);
nand U1630 (N_1630,N_1585,N_1551);
or U1631 (N_1631,N_1573,N_1582);
nand U1632 (N_1632,N_1508,N_1504);
and U1633 (N_1633,N_1536,N_1557);
and U1634 (N_1634,N_1534,N_1541);
nor U1635 (N_1635,N_1511,N_1505);
and U1636 (N_1636,N_1514,N_1529);
nand U1637 (N_1637,N_1575,N_1519);
or U1638 (N_1638,N_1572,N_1556);
or U1639 (N_1639,N_1563,N_1513);
nand U1640 (N_1640,N_1561,N_1507);
or U1641 (N_1641,N_1500,N_1570);
and U1642 (N_1642,N_1586,N_1526);
nand U1643 (N_1643,N_1517,N_1509);
nor U1644 (N_1644,N_1518,N_1599);
xor U1645 (N_1645,N_1568,N_1569);
or U1646 (N_1646,N_1521,N_1596);
nor U1647 (N_1647,N_1542,N_1520);
and U1648 (N_1648,N_1564,N_1590);
nand U1649 (N_1649,N_1589,N_1593);
and U1650 (N_1650,N_1573,N_1548);
and U1651 (N_1651,N_1572,N_1569);
or U1652 (N_1652,N_1581,N_1560);
or U1653 (N_1653,N_1537,N_1597);
nand U1654 (N_1654,N_1528,N_1537);
and U1655 (N_1655,N_1502,N_1523);
nand U1656 (N_1656,N_1543,N_1568);
and U1657 (N_1657,N_1563,N_1518);
and U1658 (N_1658,N_1588,N_1570);
nor U1659 (N_1659,N_1507,N_1596);
or U1660 (N_1660,N_1556,N_1599);
nand U1661 (N_1661,N_1512,N_1555);
or U1662 (N_1662,N_1581,N_1588);
and U1663 (N_1663,N_1585,N_1597);
nor U1664 (N_1664,N_1545,N_1541);
and U1665 (N_1665,N_1504,N_1515);
nor U1666 (N_1666,N_1507,N_1589);
and U1667 (N_1667,N_1541,N_1509);
and U1668 (N_1668,N_1529,N_1576);
nor U1669 (N_1669,N_1537,N_1580);
nand U1670 (N_1670,N_1540,N_1505);
nor U1671 (N_1671,N_1579,N_1527);
and U1672 (N_1672,N_1531,N_1546);
or U1673 (N_1673,N_1550,N_1553);
nand U1674 (N_1674,N_1561,N_1534);
or U1675 (N_1675,N_1528,N_1555);
or U1676 (N_1676,N_1575,N_1597);
nor U1677 (N_1677,N_1526,N_1519);
or U1678 (N_1678,N_1568,N_1594);
and U1679 (N_1679,N_1581,N_1566);
nor U1680 (N_1680,N_1551,N_1543);
or U1681 (N_1681,N_1577,N_1596);
nand U1682 (N_1682,N_1586,N_1560);
and U1683 (N_1683,N_1541,N_1504);
or U1684 (N_1684,N_1580,N_1512);
and U1685 (N_1685,N_1527,N_1571);
nor U1686 (N_1686,N_1540,N_1562);
or U1687 (N_1687,N_1510,N_1569);
and U1688 (N_1688,N_1565,N_1515);
and U1689 (N_1689,N_1597,N_1526);
nor U1690 (N_1690,N_1582,N_1521);
or U1691 (N_1691,N_1594,N_1523);
or U1692 (N_1692,N_1542,N_1597);
nor U1693 (N_1693,N_1595,N_1553);
or U1694 (N_1694,N_1510,N_1566);
or U1695 (N_1695,N_1502,N_1509);
or U1696 (N_1696,N_1525,N_1563);
nand U1697 (N_1697,N_1534,N_1589);
or U1698 (N_1698,N_1578,N_1571);
or U1699 (N_1699,N_1541,N_1573);
nor U1700 (N_1700,N_1638,N_1681);
nand U1701 (N_1701,N_1627,N_1618);
or U1702 (N_1702,N_1695,N_1644);
and U1703 (N_1703,N_1686,N_1658);
nor U1704 (N_1704,N_1613,N_1601);
nand U1705 (N_1705,N_1604,N_1654);
and U1706 (N_1706,N_1648,N_1661);
and U1707 (N_1707,N_1665,N_1626);
nor U1708 (N_1708,N_1679,N_1659);
and U1709 (N_1709,N_1683,N_1675);
nor U1710 (N_1710,N_1655,N_1678);
or U1711 (N_1711,N_1652,N_1673);
xnor U1712 (N_1712,N_1610,N_1685);
nand U1713 (N_1713,N_1696,N_1666);
nor U1714 (N_1714,N_1692,N_1688);
nand U1715 (N_1715,N_1625,N_1634);
nand U1716 (N_1716,N_1694,N_1642);
and U1717 (N_1717,N_1612,N_1603);
nor U1718 (N_1718,N_1630,N_1624);
nand U1719 (N_1719,N_1664,N_1615);
nand U1720 (N_1720,N_1682,N_1672);
or U1721 (N_1721,N_1670,N_1639);
or U1722 (N_1722,N_1631,N_1693);
and U1723 (N_1723,N_1640,N_1650);
xnor U1724 (N_1724,N_1632,N_1619);
nor U1725 (N_1725,N_1697,N_1636);
or U1726 (N_1726,N_1653,N_1629);
or U1727 (N_1727,N_1641,N_1622);
xor U1728 (N_1728,N_1617,N_1606);
or U1729 (N_1729,N_1623,N_1637);
nor U1730 (N_1730,N_1635,N_1607);
nor U1731 (N_1731,N_1677,N_1674);
nor U1732 (N_1732,N_1671,N_1628);
and U1733 (N_1733,N_1633,N_1600);
nor U1734 (N_1734,N_1620,N_1660);
or U1735 (N_1735,N_1646,N_1676);
nor U1736 (N_1736,N_1663,N_1602);
nand U1737 (N_1737,N_1684,N_1611);
and U1738 (N_1738,N_1662,N_1645);
nor U1739 (N_1739,N_1657,N_1621);
or U1740 (N_1740,N_1669,N_1698);
or U1741 (N_1741,N_1687,N_1605);
nand U1742 (N_1742,N_1608,N_1647);
nor U1743 (N_1743,N_1680,N_1699);
nand U1744 (N_1744,N_1690,N_1691);
and U1745 (N_1745,N_1668,N_1614);
and U1746 (N_1746,N_1616,N_1656);
or U1747 (N_1747,N_1651,N_1609);
and U1748 (N_1748,N_1667,N_1649);
and U1749 (N_1749,N_1689,N_1643);
or U1750 (N_1750,N_1681,N_1632);
and U1751 (N_1751,N_1663,N_1689);
nand U1752 (N_1752,N_1681,N_1673);
or U1753 (N_1753,N_1660,N_1624);
nand U1754 (N_1754,N_1699,N_1618);
nand U1755 (N_1755,N_1610,N_1695);
xor U1756 (N_1756,N_1608,N_1655);
nor U1757 (N_1757,N_1671,N_1619);
and U1758 (N_1758,N_1696,N_1665);
and U1759 (N_1759,N_1632,N_1646);
or U1760 (N_1760,N_1675,N_1674);
nand U1761 (N_1761,N_1667,N_1626);
and U1762 (N_1762,N_1644,N_1657);
nand U1763 (N_1763,N_1666,N_1603);
nor U1764 (N_1764,N_1678,N_1691);
and U1765 (N_1765,N_1618,N_1653);
nand U1766 (N_1766,N_1612,N_1684);
or U1767 (N_1767,N_1667,N_1636);
nand U1768 (N_1768,N_1643,N_1697);
and U1769 (N_1769,N_1642,N_1623);
nor U1770 (N_1770,N_1698,N_1659);
or U1771 (N_1771,N_1629,N_1697);
or U1772 (N_1772,N_1604,N_1689);
and U1773 (N_1773,N_1681,N_1653);
and U1774 (N_1774,N_1621,N_1680);
and U1775 (N_1775,N_1679,N_1657);
nand U1776 (N_1776,N_1618,N_1633);
and U1777 (N_1777,N_1685,N_1605);
and U1778 (N_1778,N_1674,N_1630);
nor U1779 (N_1779,N_1643,N_1601);
and U1780 (N_1780,N_1689,N_1645);
or U1781 (N_1781,N_1638,N_1616);
and U1782 (N_1782,N_1677,N_1660);
nor U1783 (N_1783,N_1673,N_1699);
nor U1784 (N_1784,N_1600,N_1611);
nor U1785 (N_1785,N_1619,N_1650);
and U1786 (N_1786,N_1682,N_1603);
nand U1787 (N_1787,N_1638,N_1605);
nor U1788 (N_1788,N_1657,N_1699);
nor U1789 (N_1789,N_1698,N_1649);
nand U1790 (N_1790,N_1648,N_1673);
and U1791 (N_1791,N_1681,N_1633);
nand U1792 (N_1792,N_1626,N_1653);
and U1793 (N_1793,N_1603,N_1642);
or U1794 (N_1794,N_1655,N_1619);
or U1795 (N_1795,N_1696,N_1654);
or U1796 (N_1796,N_1627,N_1660);
nor U1797 (N_1797,N_1609,N_1681);
nor U1798 (N_1798,N_1607,N_1630);
or U1799 (N_1799,N_1602,N_1627);
xor U1800 (N_1800,N_1764,N_1720);
or U1801 (N_1801,N_1715,N_1789);
and U1802 (N_1802,N_1723,N_1755);
and U1803 (N_1803,N_1767,N_1742);
xnor U1804 (N_1804,N_1745,N_1703);
and U1805 (N_1805,N_1726,N_1709);
or U1806 (N_1806,N_1710,N_1757);
nor U1807 (N_1807,N_1758,N_1775);
nor U1808 (N_1808,N_1766,N_1734);
nor U1809 (N_1809,N_1722,N_1704);
nor U1810 (N_1810,N_1701,N_1752);
or U1811 (N_1811,N_1744,N_1702);
and U1812 (N_1812,N_1763,N_1787);
or U1813 (N_1813,N_1753,N_1738);
or U1814 (N_1814,N_1781,N_1774);
nand U1815 (N_1815,N_1777,N_1731);
nor U1816 (N_1816,N_1732,N_1791);
and U1817 (N_1817,N_1783,N_1770);
xnor U1818 (N_1818,N_1729,N_1740);
nor U1819 (N_1819,N_1799,N_1765);
nor U1820 (N_1820,N_1776,N_1779);
nor U1821 (N_1821,N_1728,N_1793);
nand U1822 (N_1822,N_1739,N_1727);
nand U1823 (N_1823,N_1751,N_1784);
or U1824 (N_1824,N_1717,N_1713);
nor U1825 (N_1825,N_1786,N_1714);
nand U1826 (N_1826,N_1771,N_1718);
nand U1827 (N_1827,N_1756,N_1768);
nand U1828 (N_1828,N_1716,N_1721);
nor U1829 (N_1829,N_1748,N_1780);
nand U1830 (N_1830,N_1798,N_1725);
nor U1831 (N_1831,N_1733,N_1769);
nand U1832 (N_1832,N_1747,N_1792);
and U1833 (N_1833,N_1797,N_1762);
nor U1834 (N_1834,N_1754,N_1700);
nand U1835 (N_1835,N_1730,N_1778);
and U1836 (N_1836,N_1706,N_1708);
nand U1837 (N_1837,N_1750,N_1724);
or U1838 (N_1838,N_1735,N_1749);
nor U1839 (N_1839,N_1795,N_1743);
nor U1840 (N_1840,N_1707,N_1788);
and U1841 (N_1841,N_1712,N_1759);
nor U1842 (N_1842,N_1705,N_1711);
and U1843 (N_1843,N_1746,N_1737);
and U1844 (N_1844,N_1785,N_1782);
nor U1845 (N_1845,N_1794,N_1796);
nor U1846 (N_1846,N_1773,N_1736);
nand U1847 (N_1847,N_1760,N_1761);
or U1848 (N_1848,N_1741,N_1719);
or U1849 (N_1849,N_1790,N_1772);
or U1850 (N_1850,N_1726,N_1705);
nor U1851 (N_1851,N_1790,N_1789);
or U1852 (N_1852,N_1779,N_1744);
nand U1853 (N_1853,N_1781,N_1706);
or U1854 (N_1854,N_1710,N_1797);
nor U1855 (N_1855,N_1742,N_1790);
or U1856 (N_1856,N_1707,N_1737);
and U1857 (N_1857,N_1762,N_1752);
and U1858 (N_1858,N_1756,N_1791);
and U1859 (N_1859,N_1791,N_1740);
or U1860 (N_1860,N_1789,N_1762);
or U1861 (N_1861,N_1737,N_1735);
nor U1862 (N_1862,N_1732,N_1709);
and U1863 (N_1863,N_1792,N_1754);
and U1864 (N_1864,N_1777,N_1764);
nor U1865 (N_1865,N_1761,N_1790);
nor U1866 (N_1866,N_1740,N_1724);
nor U1867 (N_1867,N_1771,N_1754);
or U1868 (N_1868,N_1753,N_1727);
or U1869 (N_1869,N_1749,N_1721);
and U1870 (N_1870,N_1768,N_1714);
nor U1871 (N_1871,N_1723,N_1741);
xnor U1872 (N_1872,N_1732,N_1782);
and U1873 (N_1873,N_1753,N_1754);
and U1874 (N_1874,N_1795,N_1780);
or U1875 (N_1875,N_1772,N_1738);
or U1876 (N_1876,N_1738,N_1719);
or U1877 (N_1877,N_1706,N_1710);
xnor U1878 (N_1878,N_1790,N_1759);
nor U1879 (N_1879,N_1763,N_1735);
nor U1880 (N_1880,N_1700,N_1719);
nand U1881 (N_1881,N_1723,N_1762);
or U1882 (N_1882,N_1712,N_1710);
nand U1883 (N_1883,N_1737,N_1734);
nand U1884 (N_1884,N_1728,N_1778);
and U1885 (N_1885,N_1794,N_1789);
nor U1886 (N_1886,N_1737,N_1778);
nand U1887 (N_1887,N_1706,N_1792);
or U1888 (N_1888,N_1747,N_1766);
xnor U1889 (N_1889,N_1777,N_1712);
nor U1890 (N_1890,N_1775,N_1702);
nor U1891 (N_1891,N_1758,N_1707);
xnor U1892 (N_1892,N_1731,N_1743);
and U1893 (N_1893,N_1744,N_1733);
nand U1894 (N_1894,N_1748,N_1744);
nor U1895 (N_1895,N_1764,N_1745);
or U1896 (N_1896,N_1766,N_1726);
nand U1897 (N_1897,N_1723,N_1782);
nand U1898 (N_1898,N_1711,N_1795);
and U1899 (N_1899,N_1718,N_1760);
xnor U1900 (N_1900,N_1844,N_1819);
or U1901 (N_1901,N_1842,N_1886);
nor U1902 (N_1902,N_1885,N_1887);
and U1903 (N_1903,N_1891,N_1880);
nand U1904 (N_1904,N_1855,N_1867);
nand U1905 (N_1905,N_1898,N_1870);
nor U1906 (N_1906,N_1830,N_1850);
nor U1907 (N_1907,N_1814,N_1829);
nor U1908 (N_1908,N_1882,N_1884);
nand U1909 (N_1909,N_1853,N_1838);
and U1910 (N_1910,N_1878,N_1857);
and U1911 (N_1911,N_1862,N_1897);
and U1912 (N_1912,N_1864,N_1823);
nand U1913 (N_1913,N_1800,N_1876);
or U1914 (N_1914,N_1813,N_1883);
nand U1915 (N_1915,N_1865,N_1833);
nor U1916 (N_1916,N_1824,N_1888);
nor U1917 (N_1917,N_1854,N_1866);
and U1918 (N_1918,N_1852,N_1861);
and U1919 (N_1919,N_1805,N_1816);
nand U1920 (N_1920,N_1820,N_1863);
nand U1921 (N_1921,N_1825,N_1812);
nor U1922 (N_1922,N_1890,N_1892);
and U1923 (N_1923,N_1881,N_1843);
nor U1924 (N_1924,N_1851,N_1822);
or U1925 (N_1925,N_1874,N_1839);
or U1926 (N_1926,N_1834,N_1859);
or U1927 (N_1927,N_1858,N_1860);
and U1928 (N_1928,N_1836,N_1856);
nor U1929 (N_1929,N_1826,N_1803);
nand U1930 (N_1930,N_1889,N_1847);
and U1931 (N_1931,N_1804,N_1821);
and U1932 (N_1932,N_1815,N_1831);
nor U1933 (N_1933,N_1806,N_1873);
nand U1934 (N_1934,N_1896,N_1840);
nand U1935 (N_1935,N_1817,N_1848);
nand U1936 (N_1936,N_1810,N_1894);
nor U1937 (N_1937,N_1801,N_1849);
nand U1938 (N_1938,N_1802,N_1837);
nand U1939 (N_1939,N_1832,N_1809);
nor U1940 (N_1940,N_1879,N_1808);
and U1941 (N_1941,N_1875,N_1872);
nor U1942 (N_1942,N_1868,N_1807);
nor U1943 (N_1943,N_1895,N_1877);
nand U1944 (N_1944,N_1811,N_1869);
or U1945 (N_1945,N_1827,N_1845);
nor U1946 (N_1946,N_1841,N_1828);
nor U1947 (N_1947,N_1818,N_1899);
and U1948 (N_1948,N_1871,N_1893);
and U1949 (N_1949,N_1846,N_1835);
nand U1950 (N_1950,N_1897,N_1894);
and U1951 (N_1951,N_1869,N_1879);
or U1952 (N_1952,N_1885,N_1823);
or U1953 (N_1953,N_1898,N_1829);
nand U1954 (N_1954,N_1818,N_1808);
or U1955 (N_1955,N_1811,N_1832);
nor U1956 (N_1956,N_1822,N_1808);
and U1957 (N_1957,N_1872,N_1890);
and U1958 (N_1958,N_1850,N_1834);
nand U1959 (N_1959,N_1845,N_1813);
nand U1960 (N_1960,N_1853,N_1888);
nor U1961 (N_1961,N_1813,N_1857);
and U1962 (N_1962,N_1804,N_1819);
or U1963 (N_1963,N_1837,N_1881);
nor U1964 (N_1964,N_1810,N_1899);
and U1965 (N_1965,N_1837,N_1850);
or U1966 (N_1966,N_1837,N_1894);
nor U1967 (N_1967,N_1857,N_1864);
nor U1968 (N_1968,N_1826,N_1833);
nand U1969 (N_1969,N_1852,N_1859);
or U1970 (N_1970,N_1870,N_1860);
and U1971 (N_1971,N_1882,N_1893);
xnor U1972 (N_1972,N_1817,N_1808);
and U1973 (N_1973,N_1868,N_1865);
and U1974 (N_1974,N_1803,N_1814);
or U1975 (N_1975,N_1849,N_1818);
and U1976 (N_1976,N_1827,N_1853);
and U1977 (N_1977,N_1860,N_1869);
nor U1978 (N_1978,N_1808,N_1888);
and U1979 (N_1979,N_1869,N_1827);
nor U1980 (N_1980,N_1898,N_1872);
nor U1981 (N_1981,N_1863,N_1864);
nor U1982 (N_1982,N_1839,N_1803);
nand U1983 (N_1983,N_1873,N_1816);
nor U1984 (N_1984,N_1833,N_1897);
and U1985 (N_1985,N_1830,N_1853);
nand U1986 (N_1986,N_1869,N_1881);
nand U1987 (N_1987,N_1859,N_1880);
xnor U1988 (N_1988,N_1852,N_1830);
nor U1989 (N_1989,N_1806,N_1886);
or U1990 (N_1990,N_1840,N_1856);
and U1991 (N_1991,N_1802,N_1894);
or U1992 (N_1992,N_1833,N_1842);
and U1993 (N_1993,N_1865,N_1886);
nand U1994 (N_1994,N_1801,N_1802);
and U1995 (N_1995,N_1807,N_1873);
nor U1996 (N_1996,N_1855,N_1829);
nand U1997 (N_1997,N_1874,N_1860);
and U1998 (N_1998,N_1897,N_1808);
nand U1999 (N_1999,N_1882,N_1820);
or U2000 (N_2000,N_1926,N_1938);
or U2001 (N_2001,N_1912,N_1985);
nor U2002 (N_2002,N_1953,N_1911);
and U2003 (N_2003,N_1934,N_1909);
and U2004 (N_2004,N_1961,N_1967);
nor U2005 (N_2005,N_1930,N_1960);
and U2006 (N_2006,N_1900,N_1944);
and U2007 (N_2007,N_1988,N_1943);
nand U2008 (N_2008,N_1946,N_1939);
xnor U2009 (N_2009,N_1951,N_1927);
and U2010 (N_2010,N_1966,N_1991);
and U2011 (N_2011,N_1954,N_1940);
and U2012 (N_2012,N_1968,N_1941);
or U2013 (N_2013,N_1974,N_1996);
nor U2014 (N_2014,N_1936,N_1942);
xnor U2015 (N_2015,N_1981,N_1993);
and U2016 (N_2016,N_1972,N_1904);
nand U2017 (N_2017,N_1958,N_1965);
or U2018 (N_2018,N_1978,N_1956);
and U2019 (N_2019,N_1962,N_1905);
nand U2020 (N_2020,N_1922,N_1918);
or U2021 (N_2021,N_1950,N_1920);
nand U2022 (N_2022,N_1907,N_1915);
nor U2023 (N_2023,N_1999,N_1983);
xor U2024 (N_2024,N_1971,N_1901);
xor U2025 (N_2025,N_1921,N_1949);
nand U2026 (N_2026,N_1995,N_1903);
or U2027 (N_2027,N_1992,N_1928);
nand U2028 (N_2028,N_1979,N_1937);
nand U2029 (N_2029,N_1969,N_1917);
or U2030 (N_2030,N_1910,N_1997);
nand U2031 (N_2031,N_1919,N_1964);
nand U2032 (N_2032,N_1998,N_1929);
and U2033 (N_2033,N_1955,N_1924);
nor U2034 (N_2034,N_1990,N_1902);
and U2035 (N_2035,N_1963,N_1925);
or U2036 (N_2036,N_1952,N_1913);
or U2037 (N_2037,N_1986,N_1947);
or U2038 (N_2038,N_1970,N_1932);
nor U2039 (N_2039,N_1908,N_1957);
or U2040 (N_2040,N_1935,N_1984);
or U2041 (N_2041,N_1923,N_1987);
nand U2042 (N_2042,N_1994,N_1948);
and U2043 (N_2043,N_1916,N_1975);
or U2044 (N_2044,N_1931,N_1989);
nor U2045 (N_2045,N_1906,N_1976);
or U2046 (N_2046,N_1977,N_1959);
nand U2047 (N_2047,N_1982,N_1914);
and U2048 (N_2048,N_1933,N_1945);
nor U2049 (N_2049,N_1980,N_1973);
and U2050 (N_2050,N_1965,N_1964);
and U2051 (N_2051,N_1917,N_1902);
or U2052 (N_2052,N_1979,N_1941);
or U2053 (N_2053,N_1971,N_1979);
and U2054 (N_2054,N_1933,N_1983);
nor U2055 (N_2055,N_1926,N_1997);
and U2056 (N_2056,N_1954,N_1926);
or U2057 (N_2057,N_1956,N_1971);
and U2058 (N_2058,N_1973,N_1900);
nor U2059 (N_2059,N_1964,N_1921);
nand U2060 (N_2060,N_1960,N_1922);
or U2061 (N_2061,N_1904,N_1936);
xnor U2062 (N_2062,N_1901,N_1997);
nor U2063 (N_2063,N_1981,N_1923);
or U2064 (N_2064,N_1921,N_1952);
nand U2065 (N_2065,N_1929,N_1983);
nand U2066 (N_2066,N_1952,N_1946);
nand U2067 (N_2067,N_1961,N_1991);
nand U2068 (N_2068,N_1913,N_1924);
or U2069 (N_2069,N_1949,N_1960);
or U2070 (N_2070,N_1941,N_1932);
or U2071 (N_2071,N_1997,N_1912);
and U2072 (N_2072,N_1908,N_1920);
or U2073 (N_2073,N_1914,N_1975);
and U2074 (N_2074,N_1937,N_1993);
nor U2075 (N_2075,N_1900,N_1975);
nand U2076 (N_2076,N_1961,N_1912);
or U2077 (N_2077,N_1950,N_1942);
or U2078 (N_2078,N_1949,N_1958);
or U2079 (N_2079,N_1905,N_1986);
or U2080 (N_2080,N_1923,N_1912);
or U2081 (N_2081,N_1937,N_1926);
nor U2082 (N_2082,N_1936,N_1956);
nand U2083 (N_2083,N_1918,N_1939);
or U2084 (N_2084,N_1971,N_1931);
and U2085 (N_2085,N_1976,N_1969);
nand U2086 (N_2086,N_1990,N_1960);
nor U2087 (N_2087,N_1969,N_1913);
and U2088 (N_2088,N_1968,N_1908);
or U2089 (N_2089,N_1997,N_1962);
or U2090 (N_2090,N_1940,N_1998);
or U2091 (N_2091,N_1922,N_1981);
and U2092 (N_2092,N_1934,N_1902);
nor U2093 (N_2093,N_1932,N_1903);
or U2094 (N_2094,N_1961,N_1914);
nor U2095 (N_2095,N_1949,N_1922);
nand U2096 (N_2096,N_1953,N_1980);
nand U2097 (N_2097,N_1928,N_1951);
nor U2098 (N_2098,N_1957,N_1930);
nand U2099 (N_2099,N_1945,N_1999);
and U2100 (N_2100,N_2015,N_2044);
nand U2101 (N_2101,N_2014,N_2008);
nor U2102 (N_2102,N_2064,N_2092);
or U2103 (N_2103,N_2057,N_2009);
nand U2104 (N_2104,N_2045,N_2059);
nor U2105 (N_2105,N_2018,N_2069);
and U2106 (N_2106,N_2096,N_2035);
xor U2107 (N_2107,N_2000,N_2076);
nor U2108 (N_2108,N_2097,N_2037);
or U2109 (N_2109,N_2026,N_2062);
or U2110 (N_2110,N_2029,N_2078);
nand U2111 (N_2111,N_2066,N_2070);
and U2112 (N_2112,N_2017,N_2002);
nor U2113 (N_2113,N_2082,N_2049);
nand U2114 (N_2114,N_2001,N_2003);
or U2115 (N_2115,N_2087,N_2075);
nor U2116 (N_2116,N_2047,N_2038);
and U2117 (N_2117,N_2023,N_2021);
or U2118 (N_2118,N_2033,N_2022);
nand U2119 (N_2119,N_2031,N_2013);
or U2120 (N_2120,N_2095,N_2067);
and U2121 (N_2121,N_2077,N_2063);
or U2122 (N_2122,N_2039,N_2089);
or U2123 (N_2123,N_2004,N_2084);
nand U2124 (N_2124,N_2081,N_2036);
or U2125 (N_2125,N_2093,N_2053);
nor U2126 (N_2126,N_2074,N_2072);
nor U2127 (N_2127,N_2027,N_2088);
nand U2128 (N_2128,N_2058,N_2071);
and U2129 (N_2129,N_2065,N_2007);
nand U2130 (N_2130,N_2080,N_2073);
nand U2131 (N_2131,N_2046,N_2024);
xnor U2132 (N_2132,N_2020,N_2054);
nor U2133 (N_2133,N_2068,N_2083);
and U2134 (N_2134,N_2051,N_2060);
or U2135 (N_2135,N_2030,N_2042);
and U2136 (N_2136,N_2041,N_2061);
or U2137 (N_2137,N_2019,N_2048);
nand U2138 (N_2138,N_2034,N_2098);
or U2139 (N_2139,N_2099,N_2056);
or U2140 (N_2140,N_2090,N_2040);
and U2141 (N_2141,N_2079,N_2016);
nand U2142 (N_2142,N_2032,N_2094);
or U2143 (N_2143,N_2086,N_2010);
and U2144 (N_2144,N_2005,N_2011);
and U2145 (N_2145,N_2091,N_2055);
nor U2146 (N_2146,N_2043,N_2028);
and U2147 (N_2147,N_2006,N_2085);
nor U2148 (N_2148,N_2012,N_2050);
and U2149 (N_2149,N_2025,N_2052);
nand U2150 (N_2150,N_2067,N_2085);
nor U2151 (N_2151,N_2006,N_2095);
nor U2152 (N_2152,N_2071,N_2029);
nand U2153 (N_2153,N_2036,N_2088);
nor U2154 (N_2154,N_2043,N_2059);
or U2155 (N_2155,N_2005,N_2030);
nor U2156 (N_2156,N_2030,N_2061);
nor U2157 (N_2157,N_2005,N_2041);
and U2158 (N_2158,N_2020,N_2085);
nand U2159 (N_2159,N_2053,N_2072);
and U2160 (N_2160,N_2061,N_2073);
xnor U2161 (N_2161,N_2071,N_2055);
nand U2162 (N_2162,N_2073,N_2099);
or U2163 (N_2163,N_2034,N_2046);
or U2164 (N_2164,N_2073,N_2088);
or U2165 (N_2165,N_2048,N_2051);
or U2166 (N_2166,N_2087,N_2065);
xnor U2167 (N_2167,N_2032,N_2007);
and U2168 (N_2168,N_2000,N_2031);
nand U2169 (N_2169,N_2090,N_2039);
nand U2170 (N_2170,N_2009,N_2074);
or U2171 (N_2171,N_2014,N_2049);
nand U2172 (N_2172,N_2090,N_2044);
nor U2173 (N_2173,N_2051,N_2068);
and U2174 (N_2174,N_2061,N_2068);
and U2175 (N_2175,N_2014,N_2032);
nand U2176 (N_2176,N_2043,N_2093);
and U2177 (N_2177,N_2050,N_2084);
nor U2178 (N_2178,N_2088,N_2060);
or U2179 (N_2179,N_2006,N_2027);
nand U2180 (N_2180,N_2041,N_2054);
nor U2181 (N_2181,N_2010,N_2091);
nor U2182 (N_2182,N_2063,N_2047);
nand U2183 (N_2183,N_2058,N_2004);
nand U2184 (N_2184,N_2073,N_2042);
and U2185 (N_2185,N_2089,N_2043);
nor U2186 (N_2186,N_2011,N_2033);
or U2187 (N_2187,N_2082,N_2061);
nand U2188 (N_2188,N_2023,N_2028);
or U2189 (N_2189,N_2061,N_2069);
and U2190 (N_2190,N_2028,N_2061);
and U2191 (N_2191,N_2006,N_2044);
nor U2192 (N_2192,N_2086,N_2060);
nand U2193 (N_2193,N_2031,N_2041);
nand U2194 (N_2194,N_2063,N_2026);
xor U2195 (N_2195,N_2036,N_2050);
or U2196 (N_2196,N_2013,N_2012);
nor U2197 (N_2197,N_2052,N_2014);
and U2198 (N_2198,N_2040,N_2097);
and U2199 (N_2199,N_2024,N_2062);
nand U2200 (N_2200,N_2152,N_2112);
or U2201 (N_2201,N_2120,N_2196);
nand U2202 (N_2202,N_2125,N_2126);
and U2203 (N_2203,N_2166,N_2170);
nand U2204 (N_2204,N_2124,N_2156);
nor U2205 (N_2205,N_2182,N_2155);
or U2206 (N_2206,N_2157,N_2191);
or U2207 (N_2207,N_2146,N_2108);
and U2208 (N_2208,N_2149,N_2118);
nor U2209 (N_2209,N_2111,N_2186);
nor U2210 (N_2210,N_2178,N_2121);
nand U2211 (N_2211,N_2104,N_2110);
or U2212 (N_2212,N_2105,N_2174);
and U2213 (N_2213,N_2130,N_2188);
and U2214 (N_2214,N_2115,N_2160);
or U2215 (N_2215,N_2123,N_2107);
or U2216 (N_2216,N_2199,N_2180);
nor U2217 (N_2217,N_2154,N_2192);
and U2218 (N_2218,N_2136,N_2164);
nor U2219 (N_2219,N_2102,N_2128);
nand U2220 (N_2220,N_2193,N_2145);
nand U2221 (N_2221,N_2114,N_2172);
nor U2222 (N_2222,N_2132,N_2139);
and U2223 (N_2223,N_2138,N_2169);
xor U2224 (N_2224,N_2150,N_2147);
or U2225 (N_2225,N_2158,N_2141);
nor U2226 (N_2226,N_2106,N_2143);
nand U2227 (N_2227,N_2185,N_2163);
nand U2228 (N_2228,N_2109,N_2190);
and U2229 (N_2229,N_2116,N_2100);
nor U2230 (N_2230,N_2117,N_2161);
xor U2231 (N_2231,N_2198,N_2103);
nor U2232 (N_2232,N_2142,N_2179);
nor U2233 (N_2233,N_2151,N_2101);
or U2234 (N_2234,N_2176,N_2135);
or U2235 (N_2235,N_2144,N_2175);
and U2236 (N_2236,N_2165,N_2183);
nor U2237 (N_2237,N_2197,N_2181);
or U2238 (N_2238,N_2171,N_2187);
xnor U2239 (N_2239,N_2153,N_2133);
or U2240 (N_2240,N_2184,N_2119);
or U2241 (N_2241,N_2173,N_2194);
or U2242 (N_2242,N_2159,N_2148);
or U2243 (N_2243,N_2140,N_2137);
nand U2244 (N_2244,N_2129,N_2131);
and U2245 (N_2245,N_2168,N_2177);
nor U2246 (N_2246,N_2122,N_2134);
and U2247 (N_2247,N_2189,N_2162);
and U2248 (N_2248,N_2195,N_2113);
and U2249 (N_2249,N_2127,N_2167);
nand U2250 (N_2250,N_2149,N_2130);
and U2251 (N_2251,N_2107,N_2171);
nor U2252 (N_2252,N_2187,N_2149);
nand U2253 (N_2253,N_2187,N_2101);
or U2254 (N_2254,N_2117,N_2173);
nor U2255 (N_2255,N_2141,N_2184);
nor U2256 (N_2256,N_2198,N_2190);
or U2257 (N_2257,N_2127,N_2137);
nor U2258 (N_2258,N_2122,N_2158);
and U2259 (N_2259,N_2161,N_2137);
xnor U2260 (N_2260,N_2104,N_2164);
nor U2261 (N_2261,N_2137,N_2159);
or U2262 (N_2262,N_2134,N_2136);
and U2263 (N_2263,N_2124,N_2149);
nand U2264 (N_2264,N_2144,N_2194);
and U2265 (N_2265,N_2140,N_2132);
and U2266 (N_2266,N_2195,N_2106);
nand U2267 (N_2267,N_2146,N_2170);
and U2268 (N_2268,N_2116,N_2144);
and U2269 (N_2269,N_2106,N_2119);
and U2270 (N_2270,N_2151,N_2176);
and U2271 (N_2271,N_2120,N_2175);
nand U2272 (N_2272,N_2146,N_2115);
and U2273 (N_2273,N_2181,N_2185);
and U2274 (N_2274,N_2171,N_2152);
and U2275 (N_2275,N_2178,N_2183);
nand U2276 (N_2276,N_2177,N_2186);
nand U2277 (N_2277,N_2164,N_2193);
and U2278 (N_2278,N_2180,N_2103);
or U2279 (N_2279,N_2184,N_2155);
nor U2280 (N_2280,N_2137,N_2183);
or U2281 (N_2281,N_2100,N_2185);
nor U2282 (N_2282,N_2176,N_2179);
nand U2283 (N_2283,N_2165,N_2146);
nand U2284 (N_2284,N_2136,N_2149);
nand U2285 (N_2285,N_2151,N_2163);
and U2286 (N_2286,N_2131,N_2141);
nor U2287 (N_2287,N_2139,N_2111);
nor U2288 (N_2288,N_2129,N_2104);
and U2289 (N_2289,N_2135,N_2169);
nor U2290 (N_2290,N_2177,N_2198);
or U2291 (N_2291,N_2199,N_2132);
nor U2292 (N_2292,N_2188,N_2101);
and U2293 (N_2293,N_2145,N_2111);
nand U2294 (N_2294,N_2105,N_2179);
or U2295 (N_2295,N_2100,N_2160);
and U2296 (N_2296,N_2115,N_2142);
nand U2297 (N_2297,N_2197,N_2172);
nand U2298 (N_2298,N_2157,N_2123);
nor U2299 (N_2299,N_2122,N_2121);
nand U2300 (N_2300,N_2252,N_2242);
nor U2301 (N_2301,N_2226,N_2289);
nor U2302 (N_2302,N_2297,N_2241);
nand U2303 (N_2303,N_2223,N_2236);
nand U2304 (N_2304,N_2253,N_2215);
or U2305 (N_2305,N_2221,N_2291);
nor U2306 (N_2306,N_2284,N_2220);
and U2307 (N_2307,N_2217,N_2264);
and U2308 (N_2308,N_2248,N_2288);
or U2309 (N_2309,N_2294,N_2218);
and U2310 (N_2310,N_2200,N_2246);
nand U2311 (N_2311,N_2232,N_2270);
or U2312 (N_2312,N_2279,N_2299);
nand U2313 (N_2313,N_2251,N_2278);
nor U2314 (N_2314,N_2249,N_2213);
and U2315 (N_2315,N_2275,N_2280);
or U2316 (N_2316,N_2298,N_2245);
nor U2317 (N_2317,N_2206,N_2227);
or U2318 (N_2318,N_2269,N_2282);
or U2319 (N_2319,N_2230,N_2216);
or U2320 (N_2320,N_2208,N_2285);
nor U2321 (N_2321,N_2286,N_2202);
and U2322 (N_2322,N_2261,N_2235);
nand U2323 (N_2323,N_2281,N_2234);
nor U2324 (N_2324,N_2244,N_2201);
and U2325 (N_2325,N_2205,N_2283);
nor U2326 (N_2326,N_2287,N_2225);
nor U2327 (N_2327,N_2243,N_2290);
nor U2328 (N_2328,N_2250,N_2256);
nand U2329 (N_2329,N_2210,N_2259);
and U2330 (N_2330,N_2222,N_2247);
nand U2331 (N_2331,N_2276,N_2271);
nand U2332 (N_2332,N_2237,N_2296);
and U2333 (N_2333,N_2263,N_2209);
and U2334 (N_2334,N_2266,N_2240);
and U2335 (N_2335,N_2207,N_2273);
or U2336 (N_2336,N_2204,N_2231);
nand U2337 (N_2337,N_2211,N_2233);
xor U2338 (N_2338,N_2229,N_2238);
nor U2339 (N_2339,N_2277,N_2228);
nor U2340 (N_2340,N_2268,N_2224);
nor U2341 (N_2341,N_2267,N_2203);
nor U2342 (N_2342,N_2295,N_2265);
nand U2343 (N_2343,N_2212,N_2274);
and U2344 (N_2344,N_2219,N_2257);
or U2345 (N_2345,N_2260,N_2255);
and U2346 (N_2346,N_2239,N_2254);
or U2347 (N_2347,N_2258,N_2293);
and U2348 (N_2348,N_2292,N_2214);
nand U2349 (N_2349,N_2262,N_2272);
nand U2350 (N_2350,N_2232,N_2260);
nand U2351 (N_2351,N_2275,N_2228);
and U2352 (N_2352,N_2210,N_2296);
and U2353 (N_2353,N_2289,N_2218);
and U2354 (N_2354,N_2240,N_2263);
nor U2355 (N_2355,N_2258,N_2270);
nand U2356 (N_2356,N_2255,N_2293);
and U2357 (N_2357,N_2224,N_2201);
or U2358 (N_2358,N_2298,N_2234);
nor U2359 (N_2359,N_2212,N_2209);
and U2360 (N_2360,N_2290,N_2265);
nor U2361 (N_2361,N_2276,N_2245);
nor U2362 (N_2362,N_2234,N_2232);
nand U2363 (N_2363,N_2256,N_2293);
nand U2364 (N_2364,N_2233,N_2290);
and U2365 (N_2365,N_2279,N_2254);
nor U2366 (N_2366,N_2200,N_2284);
or U2367 (N_2367,N_2216,N_2237);
nand U2368 (N_2368,N_2280,N_2281);
nand U2369 (N_2369,N_2217,N_2230);
and U2370 (N_2370,N_2240,N_2204);
or U2371 (N_2371,N_2286,N_2245);
nor U2372 (N_2372,N_2289,N_2217);
nand U2373 (N_2373,N_2219,N_2244);
nand U2374 (N_2374,N_2203,N_2266);
and U2375 (N_2375,N_2253,N_2271);
or U2376 (N_2376,N_2251,N_2268);
xor U2377 (N_2377,N_2297,N_2242);
and U2378 (N_2378,N_2277,N_2257);
nor U2379 (N_2379,N_2217,N_2207);
nor U2380 (N_2380,N_2203,N_2259);
and U2381 (N_2381,N_2271,N_2270);
or U2382 (N_2382,N_2223,N_2255);
xnor U2383 (N_2383,N_2299,N_2238);
or U2384 (N_2384,N_2289,N_2214);
and U2385 (N_2385,N_2207,N_2210);
nand U2386 (N_2386,N_2253,N_2260);
nor U2387 (N_2387,N_2241,N_2268);
or U2388 (N_2388,N_2278,N_2201);
and U2389 (N_2389,N_2262,N_2235);
and U2390 (N_2390,N_2262,N_2269);
or U2391 (N_2391,N_2299,N_2254);
nor U2392 (N_2392,N_2228,N_2243);
nor U2393 (N_2393,N_2232,N_2202);
nor U2394 (N_2394,N_2214,N_2230);
and U2395 (N_2395,N_2278,N_2286);
nand U2396 (N_2396,N_2274,N_2297);
and U2397 (N_2397,N_2282,N_2239);
nand U2398 (N_2398,N_2261,N_2206);
and U2399 (N_2399,N_2277,N_2213);
or U2400 (N_2400,N_2362,N_2311);
and U2401 (N_2401,N_2374,N_2319);
nand U2402 (N_2402,N_2345,N_2367);
or U2403 (N_2403,N_2360,N_2387);
or U2404 (N_2404,N_2389,N_2315);
nor U2405 (N_2405,N_2347,N_2353);
and U2406 (N_2406,N_2343,N_2327);
or U2407 (N_2407,N_2392,N_2340);
nand U2408 (N_2408,N_2318,N_2329);
nor U2409 (N_2409,N_2368,N_2384);
and U2410 (N_2410,N_2373,N_2312);
nor U2411 (N_2411,N_2335,N_2304);
or U2412 (N_2412,N_2307,N_2391);
and U2413 (N_2413,N_2379,N_2321);
nand U2414 (N_2414,N_2313,N_2383);
and U2415 (N_2415,N_2394,N_2309);
nor U2416 (N_2416,N_2365,N_2322);
or U2417 (N_2417,N_2350,N_2377);
or U2418 (N_2418,N_2317,N_2328);
nand U2419 (N_2419,N_2308,N_2306);
nand U2420 (N_2420,N_2336,N_2354);
and U2421 (N_2421,N_2342,N_2395);
nor U2422 (N_2422,N_2366,N_2323);
and U2423 (N_2423,N_2301,N_2326);
xnor U2424 (N_2424,N_2316,N_2348);
nand U2425 (N_2425,N_2324,N_2355);
nand U2426 (N_2426,N_2351,N_2378);
nand U2427 (N_2427,N_2357,N_2352);
nand U2428 (N_2428,N_2396,N_2344);
or U2429 (N_2429,N_2320,N_2346);
and U2430 (N_2430,N_2314,N_2397);
and U2431 (N_2431,N_2330,N_2372);
nor U2432 (N_2432,N_2369,N_2386);
or U2433 (N_2433,N_2371,N_2302);
nor U2434 (N_2434,N_2334,N_2388);
nand U2435 (N_2435,N_2331,N_2381);
nand U2436 (N_2436,N_2337,N_2393);
or U2437 (N_2437,N_2333,N_2310);
nor U2438 (N_2438,N_2303,N_2356);
and U2439 (N_2439,N_2361,N_2305);
nand U2440 (N_2440,N_2363,N_2399);
nor U2441 (N_2441,N_2359,N_2370);
nor U2442 (N_2442,N_2385,N_2332);
or U2443 (N_2443,N_2300,N_2339);
nand U2444 (N_2444,N_2358,N_2341);
or U2445 (N_2445,N_2364,N_2338);
and U2446 (N_2446,N_2325,N_2382);
nand U2447 (N_2447,N_2349,N_2390);
or U2448 (N_2448,N_2376,N_2375);
nor U2449 (N_2449,N_2398,N_2380);
xnor U2450 (N_2450,N_2331,N_2325);
or U2451 (N_2451,N_2323,N_2328);
or U2452 (N_2452,N_2312,N_2381);
nor U2453 (N_2453,N_2333,N_2338);
and U2454 (N_2454,N_2306,N_2356);
or U2455 (N_2455,N_2326,N_2302);
nand U2456 (N_2456,N_2332,N_2381);
and U2457 (N_2457,N_2345,N_2371);
and U2458 (N_2458,N_2346,N_2336);
nor U2459 (N_2459,N_2306,N_2318);
and U2460 (N_2460,N_2319,N_2386);
nand U2461 (N_2461,N_2366,N_2354);
nor U2462 (N_2462,N_2341,N_2378);
nand U2463 (N_2463,N_2325,N_2377);
nor U2464 (N_2464,N_2396,N_2322);
and U2465 (N_2465,N_2348,N_2391);
nand U2466 (N_2466,N_2372,N_2352);
nand U2467 (N_2467,N_2326,N_2310);
nor U2468 (N_2468,N_2309,N_2326);
nor U2469 (N_2469,N_2323,N_2395);
or U2470 (N_2470,N_2349,N_2300);
or U2471 (N_2471,N_2363,N_2373);
or U2472 (N_2472,N_2379,N_2323);
or U2473 (N_2473,N_2328,N_2354);
nor U2474 (N_2474,N_2352,N_2334);
nand U2475 (N_2475,N_2373,N_2317);
or U2476 (N_2476,N_2386,N_2300);
and U2477 (N_2477,N_2390,N_2333);
and U2478 (N_2478,N_2349,N_2342);
and U2479 (N_2479,N_2325,N_2361);
or U2480 (N_2480,N_2310,N_2331);
or U2481 (N_2481,N_2330,N_2386);
nor U2482 (N_2482,N_2392,N_2379);
nor U2483 (N_2483,N_2370,N_2300);
and U2484 (N_2484,N_2362,N_2309);
and U2485 (N_2485,N_2382,N_2337);
or U2486 (N_2486,N_2340,N_2375);
nand U2487 (N_2487,N_2305,N_2310);
nor U2488 (N_2488,N_2314,N_2310);
nor U2489 (N_2489,N_2376,N_2341);
nor U2490 (N_2490,N_2397,N_2361);
nand U2491 (N_2491,N_2313,N_2334);
nor U2492 (N_2492,N_2316,N_2319);
or U2493 (N_2493,N_2374,N_2376);
or U2494 (N_2494,N_2381,N_2350);
nor U2495 (N_2495,N_2359,N_2378);
nor U2496 (N_2496,N_2377,N_2389);
and U2497 (N_2497,N_2323,N_2356);
or U2498 (N_2498,N_2318,N_2370);
nor U2499 (N_2499,N_2324,N_2387);
and U2500 (N_2500,N_2443,N_2415);
nand U2501 (N_2501,N_2488,N_2448);
or U2502 (N_2502,N_2417,N_2455);
nor U2503 (N_2503,N_2480,N_2494);
or U2504 (N_2504,N_2423,N_2467);
nand U2505 (N_2505,N_2466,N_2499);
nor U2506 (N_2506,N_2431,N_2454);
and U2507 (N_2507,N_2404,N_2496);
nand U2508 (N_2508,N_2459,N_2492);
xor U2509 (N_2509,N_2460,N_2478);
or U2510 (N_2510,N_2428,N_2487);
or U2511 (N_2511,N_2424,N_2416);
nand U2512 (N_2512,N_2408,N_2475);
and U2513 (N_2513,N_2479,N_2477);
nand U2514 (N_2514,N_2465,N_2469);
nor U2515 (N_2515,N_2485,N_2400);
or U2516 (N_2516,N_2483,N_2441);
and U2517 (N_2517,N_2420,N_2472);
nor U2518 (N_2518,N_2427,N_2445);
xnor U2519 (N_2519,N_2453,N_2457);
or U2520 (N_2520,N_2444,N_2456);
nor U2521 (N_2521,N_2405,N_2497);
or U2522 (N_2522,N_2484,N_2429);
nand U2523 (N_2523,N_2409,N_2411);
nand U2524 (N_2524,N_2437,N_2463);
and U2525 (N_2525,N_2482,N_2407);
or U2526 (N_2526,N_2462,N_2410);
and U2527 (N_2527,N_2476,N_2451);
and U2528 (N_2528,N_2433,N_2490);
nand U2529 (N_2529,N_2426,N_2471);
nor U2530 (N_2530,N_2498,N_2446);
or U2531 (N_2531,N_2413,N_2430);
or U2532 (N_2532,N_2402,N_2474);
nand U2533 (N_2533,N_2470,N_2495);
nand U2534 (N_2534,N_2425,N_2435);
and U2535 (N_2535,N_2414,N_2468);
and U2536 (N_2536,N_2418,N_2464);
nand U2537 (N_2537,N_2473,N_2489);
nand U2538 (N_2538,N_2493,N_2438);
nand U2539 (N_2539,N_2447,N_2422);
and U2540 (N_2540,N_2458,N_2449);
or U2541 (N_2541,N_2403,N_2439);
and U2542 (N_2542,N_2461,N_2406);
or U2543 (N_2543,N_2412,N_2450);
nand U2544 (N_2544,N_2419,N_2452);
nand U2545 (N_2545,N_2436,N_2486);
nand U2546 (N_2546,N_2481,N_2421);
and U2547 (N_2547,N_2491,N_2434);
nand U2548 (N_2548,N_2442,N_2440);
and U2549 (N_2549,N_2401,N_2432);
nand U2550 (N_2550,N_2417,N_2478);
or U2551 (N_2551,N_2452,N_2478);
and U2552 (N_2552,N_2446,N_2449);
or U2553 (N_2553,N_2487,N_2465);
and U2554 (N_2554,N_2493,N_2492);
nor U2555 (N_2555,N_2406,N_2475);
nor U2556 (N_2556,N_2499,N_2484);
or U2557 (N_2557,N_2422,N_2412);
or U2558 (N_2558,N_2450,N_2476);
nand U2559 (N_2559,N_2440,N_2467);
nand U2560 (N_2560,N_2461,N_2494);
or U2561 (N_2561,N_2492,N_2472);
nor U2562 (N_2562,N_2484,N_2427);
nor U2563 (N_2563,N_2495,N_2440);
nand U2564 (N_2564,N_2435,N_2431);
and U2565 (N_2565,N_2482,N_2483);
or U2566 (N_2566,N_2469,N_2490);
nor U2567 (N_2567,N_2482,N_2464);
nand U2568 (N_2568,N_2411,N_2464);
nor U2569 (N_2569,N_2469,N_2495);
nand U2570 (N_2570,N_2472,N_2462);
or U2571 (N_2571,N_2462,N_2495);
and U2572 (N_2572,N_2429,N_2455);
and U2573 (N_2573,N_2499,N_2495);
and U2574 (N_2574,N_2424,N_2443);
nand U2575 (N_2575,N_2415,N_2485);
nand U2576 (N_2576,N_2407,N_2474);
nor U2577 (N_2577,N_2457,N_2440);
and U2578 (N_2578,N_2439,N_2474);
nand U2579 (N_2579,N_2404,N_2485);
or U2580 (N_2580,N_2451,N_2423);
or U2581 (N_2581,N_2459,N_2408);
xnor U2582 (N_2582,N_2496,N_2488);
nand U2583 (N_2583,N_2479,N_2499);
nand U2584 (N_2584,N_2443,N_2489);
nand U2585 (N_2585,N_2432,N_2449);
nand U2586 (N_2586,N_2484,N_2411);
nor U2587 (N_2587,N_2445,N_2449);
and U2588 (N_2588,N_2453,N_2436);
nor U2589 (N_2589,N_2467,N_2472);
or U2590 (N_2590,N_2458,N_2416);
or U2591 (N_2591,N_2401,N_2453);
or U2592 (N_2592,N_2468,N_2495);
xnor U2593 (N_2593,N_2434,N_2418);
and U2594 (N_2594,N_2479,N_2489);
nor U2595 (N_2595,N_2462,N_2448);
nor U2596 (N_2596,N_2480,N_2457);
or U2597 (N_2597,N_2419,N_2429);
nand U2598 (N_2598,N_2404,N_2431);
nor U2599 (N_2599,N_2422,N_2475);
and U2600 (N_2600,N_2520,N_2542);
nand U2601 (N_2601,N_2518,N_2530);
nand U2602 (N_2602,N_2596,N_2588);
nor U2603 (N_2603,N_2540,N_2585);
or U2604 (N_2604,N_2567,N_2539);
and U2605 (N_2605,N_2599,N_2544);
nor U2606 (N_2606,N_2545,N_2514);
nor U2607 (N_2607,N_2536,N_2512);
nor U2608 (N_2608,N_2598,N_2572);
nor U2609 (N_2609,N_2581,N_2571);
nor U2610 (N_2610,N_2534,N_2503);
or U2611 (N_2611,N_2582,N_2575);
nand U2612 (N_2612,N_2516,N_2517);
nand U2613 (N_2613,N_2524,N_2537);
and U2614 (N_2614,N_2506,N_2553);
or U2615 (N_2615,N_2583,N_2509);
and U2616 (N_2616,N_2592,N_2521);
nor U2617 (N_2617,N_2527,N_2538);
or U2618 (N_2618,N_2558,N_2566);
and U2619 (N_2619,N_2502,N_2511);
nor U2620 (N_2620,N_2504,N_2507);
nor U2621 (N_2621,N_2528,N_2579);
and U2622 (N_2622,N_2561,N_2555);
nand U2623 (N_2623,N_2505,N_2500);
and U2624 (N_2624,N_2543,N_2529);
nor U2625 (N_2625,N_2557,N_2501);
nor U2626 (N_2626,N_2515,N_2573);
nand U2627 (N_2627,N_2584,N_2560);
nor U2628 (N_2628,N_2578,N_2577);
xnor U2629 (N_2629,N_2568,N_2548);
nand U2630 (N_2630,N_2576,N_2546);
and U2631 (N_2631,N_2513,N_2552);
and U2632 (N_2632,N_2563,N_2594);
and U2633 (N_2633,N_2565,N_2574);
nand U2634 (N_2634,N_2595,N_2549);
or U2635 (N_2635,N_2522,N_2554);
or U2636 (N_2636,N_2597,N_2589);
nor U2637 (N_2637,N_2510,N_2562);
and U2638 (N_2638,N_2590,N_2531);
or U2639 (N_2639,N_2556,N_2523);
or U2640 (N_2640,N_2535,N_2591);
and U2641 (N_2641,N_2508,N_2547);
or U2642 (N_2642,N_2570,N_2551);
nand U2643 (N_2643,N_2525,N_2559);
and U2644 (N_2644,N_2564,N_2541);
nand U2645 (N_2645,N_2569,N_2519);
nand U2646 (N_2646,N_2533,N_2586);
or U2647 (N_2647,N_2526,N_2550);
or U2648 (N_2648,N_2593,N_2532);
and U2649 (N_2649,N_2580,N_2587);
nor U2650 (N_2650,N_2580,N_2589);
and U2651 (N_2651,N_2509,N_2511);
and U2652 (N_2652,N_2598,N_2599);
and U2653 (N_2653,N_2568,N_2526);
or U2654 (N_2654,N_2544,N_2554);
nand U2655 (N_2655,N_2592,N_2517);
nand U2656 (N_2656,N_2525,N_2592);
and U2657 (N_2657,N_2526,N_2505);
and U2658 (N_2658,N_2515,N_2520);
nor U2659 (N_2659,N_2549,N_2542);
and U2660 (N_2660,N_2586,N_2566);
and U2661 (N_2661,N_2508,N_2503);
or U2662 (N_2662,N_2521,N_2502);
and U2663 (N_2663,N_2585,N_2550);
and U2664 (N_2664,N_2529,N_2573);
and U2665 (N_2665,N_2579,N_2577);
nand U2666 (N_2666,N_2521,N_2554);
nand U2667 (N_2667,N_2507,N_2515);
xor U2668 (N_2668,N_2584,N_2518);
and U2669 (N_2669,N_2512,N_2525);
xnor U2670 (N_2670,N_2540,N_2570);
xnor U2671 (N_2671,N_2533,N_2534);
or U2672 (N_2672,N_2535,N_2596);
xor U2673 (N_2673,N_2503,N_2564);
or U2674 (N_2674,N_2569,N_2534);
and U2675 (N_2675,N_2503,N_2583);
nand U2676 (N_2676,N_2531,N_2529);
and U2677 (N_2677,N_2513,N_2527);
nand U2678 (N_2678,N_2544,N_2512);
nor U2679 (N_2679,N_2597,N_2551);
or U2680 (N_2680,N_2555,N_2553);
or U2681 (N_2681,N_2587,N_2550);
nor U2682 (N_2682,N_2536,N_2517);
or U2683 (N_2683,N_2577,N_2561);
nand U2684 (N_2684,N_2550,N_2501);
nand U2685 (N_2685,N_2503,N_2592);
nand U2686 (N_2686,N_2515,N_2516);
nor U2687 (N_2687,N_2546,N_2534);
and U2688 (N_2688,N_2531,N_2539);
nor U2689 (N_2689,N_2532,N_2554);
nand U2690 (N_2690,N_2516,N_2541);
and U2691 (N_2691,N_2599,N_2514);
and U2692 (N_2692,N_2512,N_2510);
and U2693 (N_2693,N_2590,N_2546);
or U2694 (N_2694,N_2529,N_2593);
or U2695 (N_2695,N_2574,N_2591);
nand U2696 (N_2696,N_2594,N_2571);
nand U2697 (N_2697,N_2503,N_2568);
nand U2698 (N_2698,N_2533,N_2500);
nor U2699 (N_2699,N_2554,N_2545);
or U2700 (N_2700,N_2671,N_2694);
and U2701 (N_2701,N_2632,N_2636);
or U2702 (N_2702,N_2607,N_2629);
and U2703 (N_2703,N_2649,N_2628);
nand U2704 (N_2704,N_2643,N_2615);
and U2705 (N_2705,N_2630,N_2638);
and U2706 (N_2706,N_2635,N_2691);
and U2707 (N_2707,N_2623,N_2676);
nor U2708 (N_2708,N_2621,N_2692);
nand U2709 (N_2709,N_2681,N_2646);
nor U2710 (N_2710,N_2696,N_2603);
nor U2711 (N_2711,N_2631,N_2669);
and U2712 (N_2712,N_2687,N_2622);
or U2713 (N_2713,N_2642,N_2624);
and U2714 (N_2714,N_2637,N_2652);
nor U2715 (N_2715,N_2625,N_2605);
nor U2716 (N_2716,N_2677,N_2618);
nor U2717 (N_2717,N_2674,N_2699);
nand U2718 (N_2718,N_2655,N_2683);
nor U2719 (N_2719,N_2650,N_2697);
or U2720 (N_2720,N_2686,N_2657);
nor U2721 (N_2721,N_2665,N_2612);
and U2722 (N_2722,N_2658,N_2695);
and U2723 (N_2723,N_2662,N_2634);
nand U2724 (N_2724,N_2675,N_2644);
nand U2725 (N_2725,N_2664,N_2606);
nand U2726 (N_2726,N_2667,N_2660);
nand U2727 (N_2727,N_2678,N_2626);
nand U2728 (N_2728,N_2682,N_2613);
nand U2729 (N_2729,N_2684,N_2647);
nand U2730 (N_2730,N_2609,N_2641);
or U2731 (N_2731,N_2666,N_2620);
nor U2732 (N_2732,N_2698,N_2651);
or U2733 (N_2733,N_2653,N_2616);
nor U2734 (N_2734,N_2602,N_2690);
nand U2735 (N_2735,N_2619,N_2614);
nor U2736 (N_2736,N_2661,N_2659);
nor U2737 (N_2737,N_2693,N_2685);
or U2738 (N_2738,N_2617,N_2656);
or U2739 (N_2739,N_2611,N_2663);
nor U2740 (N_2740,N_2633,N_2608);
nor U2741 (N_2741,N_2680,N_2627);
nor U2742 (N_2742,N_2670,N_2645);
nor U2743 (N_2743,N_2672,N_2601);
and U2744 (N_2744,N_2679,N_2668);
or U2745 (N_2745,N_2610,N_2688);
and U2746 (N_2746,N_2654,N_2673);
or U2747 (N_2747,N_2604,N_2639);
nor U2748 (N_2748,N_2648,N_2640);
and U2749 (N_2749,N_2600,N_2689);
or U2750 (N_2750,N_2603,N_2620);
nor U2751 (N_2751,N_2658,N_2694);
nand U2752 (N_2752,N_2661,N_2674);
or U2753 (N_2753,N_2631,N_2609);
nor U2754 (N_2754,N_2692,N_2699);
or U2755 (N_2755,N_2692,N_2647);
or U2756 (N_2756,N_2658,N_2678);
nor U2757 (N_2757,N_2689,N_2688);
xnor U2758 (N_2758,N_2649,N_2654);
or U2759 (N_2759,N_2643,N_2670);
or U2760 (N_2760,N_2665,N_2653);
nand U2761 (N_2761,N_2639,N_2601);
and U2762 (N_2762,N_2668,N_2673);
or U2763 (N_2763,N_2654,N_2671);
or U2764 (N_2764,N_2678,N_2697);
xnor U2765 (N_2765,N_2618,N_2658);
or U2766 (N_2766,N_2672,N_2610);
or U2767 (N_2767,N_2676,N_2619);
and U2768 (N_2768,N_2645,N_2605);
or U2769 (N_2769,N_2629,N_2659);
nor U2770 (N_2770,N_2625,N_2689);
and U2771 (N_2771,N_2651,N_2644);
or U2772 (N_2772,N_2663,N_2632);
nand U2773 (N_2773,N_2603,N_2655);
nor U2774 (N_2774,N_2621,N_2644);
or U2775 (N_2775,N_2671,N_2617);
or U2776 (N_2776,N_2631,N_2675);
nand U2777 (N_2777,N_2679,N_2629);
or U2778 (N_2778,N_2615,N_2666);
nand U2779 (N_2779,N_2613,N_2609);
or U2780 (N_2780,N_2682,N_2609);
and U2781 (N_2781,N_2659,N_2600);
or U2782 (N_2782,N_2629,N_2685);
or U2783 (N_2783,N_2634,N_2617);
nor U2784 (N_2784,N_2645,N_2694);
nand U2785 (N_2785,N_2677,N_2649);
nor U2786 (N_2786,N_2614,N_2642);
or U2787 (N_2787,N_2697,N_2669);
and U2788 (N_2788,N_2655,N_2632);
and U2789 (N_2789,N_2627,N_2601);
nor U2790 (N_2790,N_2612,N_2621);
and U2791 (N_2791,N_2629,N_2645);
or U2792 (N_2792,N_2682,N_2670);
or U2793 (N_2793,N_2625,N_2695);
nand U2794 (N_2794,N_2622,N_2680);
nor U2795 (N_2795,N_2616,N_2637);
nor U2796 (N_2796,N_2615,N_2678);
nand U2797 (N_2797,N_2653,N_2654);
nand U2798 (N_2798,N_2671,N_2647);
or U2799 (N_2799,N_2658,N_2685);
or U2800 (N_2800,N_2746,N_2728);
and U2801 (N_2801,N_2778,N_2784);
nand U2802 (N_2802,N_2712,N_2754);
nand U2803 (N_2803,N_2735,N_2721);
or U2804 (N_2804,N_2720,N_2772);
nor U2805 (N_2805,N_2750,N_2760);
or U2806 (N_2806,N_2748,N_2763);
nand U2807 (N_2807,N_2774,N_2724);
and U2808 (N_2808,N_2734,N_2745);
and U2809 (N_2809,N_2780,N_2788);
or U2810 (N_2810,N_2704,N_2719);
or U2811 (N_2811,N_2787,N_2727);
and U2812 (N_2812,N_2789,N_2708);
nor U2813 (N_2813,N_2792,N_2781);
or U2814 (N_2814,N_2723,N_2702);
nand U2815 (N_2815,N_2798,N_2744);
nand U2816 (N_2816,N_2747,N_2762);
and U2817 (N_2817,N_2777,N_2799);
nand U2818 (N_2818,N_2740,N_2782);
or U2819 (N_2819,N_2729,N_2770);
xor U2820 (N_2820,N_2715,N_2741);
and U2821 (N_2821,N_2767,N_2786);
or U2822 (N_2822,N_2783,N_2709);
nand U2823 (N_2823,N_2707,N_2714);
and U2824 (N_2824,N_2764,N_2725);
nor U2825 (N_2825,N_2773,N_2733);
nand U2826 (N_2826,N_2706,N_2705);
or U2827 (N_2827,N_2730,N_2756);
nand U2828 (N_2828,N_2755,N_2710);
or U2829 (N_2829,N_2732,N_2713);
or U2830 (N_2830,N_2743,N_2738);
nor U2831 (N_2831,N_2739,N_2711);
nor U2832 (N_2832,N_2716,N_2717);
or U2833 (N_2833,N_2731,N_2795);
or U2834 (N_2834,N_2796,N_2752);
nor U2835 (N_2835,N_2753,N_2776);
and U2836 (N_2836,N_2790,N_2749);
nor U2837 (N_2837,N_2757,N_2779);
nor U2838 (N_2838,N_2726,N_2793);
nand U2839 (N_2839,N_2768,N_2785);
nor U2840 (N_2840,N_2797,N_2703);
and U2841 (N_2841,N_2758,N_2742);
and U2842 (N_2842,N_2761,N_2766);
nand U2843 (N_2843,N_2751,N_2737);
nand U2844 (N_2844,N_2722,N_2718);
nor U2845 (N_2845,N_2700,N_2794);
nand U2846 (N_2846,N_2736,N_2791);
or U2847 (N_2847,N_2765,N_2775);
or U2848 (N_2848,N_2701,N_2771);
nor U2849 (N_2849,N_2759,N_2769);
nor U2850 (N_2850,N_2750,N_2731);
and U2851 (N_2851,N_2781,N_2732);
or U2852 (N_2852,N_2755,N_2785);
or U2853 (N_2853,N_2765,N_2798);
and U2854 (N_2854,N_2785,N_2726);
nor U2855 (N_2855,N_2741,N_2758);
or U2856 (N_2856,N_2799,N_2703);
nor U2857 (N_2857,N_2723,N_2755);
or U2858 (N_2858,N_2705,N_2737);
nor U2859 (N_2859,N_2706,N_2709);
or U2860 (N_2860,N_2757,N_2709);
nand U2861 (N_2861,N_2745,N_2700);
nand U2862 (N_2862,N_2781,N_2704);
and U2863 (N_2863,N_2752,N_2721);
or U2864 (N_2864,N_2775,N_2733);
or U2865 (N_2865,N_2761,N_2798);
nor U2866 (N_2866,N_2711,N_2776);
and U2867 (N_2867,N_2759,N_2722);
and U2868 (N_2868,N_2771,N_2722);
and U2869 (N_2869,N_2759,N_2714);
nor U2870 (N_2870,N_2703,N_2769);
nand U2871 (N_2871,N_2736,N_2714);
and U2872 (N_2872,N_2715,N_2766);
and U2873 (N_2873,N_2710,N_2784);
or U2874 (N_2874,N_2791,N_2799);
nor U2875 (N_2875,N_2771,N_2716);
and U2876 (N_2876,N_2725,N_2788);
nand U2877 (N_2877,N_2781,N_2788);
nor U2878 (N_2878,N_2789,N_2770);
nor U2879 (N_2879,N_2790,N_2706);
nor U2880 (N_2880,N_2771,N_2768);
nand U2881 (N_2881,N_2716,N_2728);
nor U2882 (N_2882,N_2736,N_2709);
nor U2883 (N_2883,N_2717,N_2701);
nor U2884 (N_2884,N_2746,N_2731);
nor U2885 (N_2885,N_2774,N_2780);
nand U2886 (N_2886,N_2716,N_2780);
nor U2887 (N_2887,N_2750,N_2704);
nor U2888 (N_2888,N_2720,N_2775);
or U2889 (N_2889,N_2755,N_2726);
nand U2890 (N_2890,N_2742,N_2751);
or U2891 (N_2891,N_2747,N_2778);
nand U2892 (N_2892,N_2731,N_2767);
and U2893 (N_2893,N_2784,N_2799);
and U2894 (N_2894,N_2722,N_2778);
nor U2895 (N_2895,N_2774,N_2775);
nor U2896 (N_2896,N_2763,N_2759);
and U2897 (N_2897,N_2709,N_2704);
nand U2898 (N_2898,N_2704,N_2737);
or U2899 (N_2899,N_2753,N_2726);
or U2900 (N_2900,N_2817,N_2808);
nand U2901 (N_2901,N_2890,N_2805);
and U2902 (N_2902,N_2813,N_2810);
nor U2903 (N_2903,N_2872,N_2802);
and U2904 (N_2904,N_2857,N_2856);
nor U2905 (N_2905,N_2814,N_2825);
or U2906 (N_2906,N_2829,N_2807);
or U2907 (N_2907,N_2892,N_2869);
nand U2908 (N_2908,N_2812,N_2837);
nor U2909 (N_2909,N_2853,N_2809);
or U2910 (N_2910,N_2843,N_2852);
nand U2911 (N_2911,N_2891,N_2854);
nor U2912 (N_2912,N_2862,N_2887);
nand U2913 (N_2913,N_2845,N_2848);
nor U2914 (N_2914,N_2844,N_2841);
nand U2915 (N_2915,N_2840,N_2896);
or U2916 (N_2916,N_2897,N_2801);
xnor U2917 (N_2917,N_2834,N_2885);
and U2918 (N_2918,N_2831,N_2894);
or U2919 (N_2919,N_2826,N_2861);
nand U2920 (N_2920,N_2893,N_2880);
xnor U2921 (N_2921,N_2882,N_2803);
nor U2922 (N_2922,N_2835,N_2832);
nor U2923 (N_2923,N_2818,N_2827);
or U2924 (N_2924,N_2804,N_2863);
nand U2925 (N_2925,N_2849,N_2823);
and U2926 (N_2926,N_2877,N_2868);
and U2927 (N_2927,N_2884,N_2859);
or U2928 (N_2928,N_2811,N_2850);
nand U2929 (N_2929,N_2846,N_2847);
or U2930 (N_2930,N_2889,N_2816);
or U2931 (N_2931,N_2822,N_2819);
or U2932 (N_2932,N_2830,N_2867);
nor U2933 (N_2933,N_2806,N_2855);
or U2934 (N_2934,N_2899,N_2800);
nor U2935 (N_2935,N_2821,N_2888);
and U2936 (N_2936,N_2860,N_2879);
nand U2937 (N_2937,N_2870,N_2875);
nand U2938 (N_2938,N_2895,N_2864);
nor U2939 (N_2939,N_2873,N_2865);
or U2940 (N_2940,N_2883,N_2842);
and U2941 (N_2941,N_2833,N_2828);
or U2942 (N_2942,N_2815,N_2824);
and U2943 (N_2943,N_2886,N_2881);
nor U2944 (N_2944,N_2898,N_2878);
nor U2945 (N_2945,N_2851,N_2874);
nor U2946 (N_2946,N_2876,N_2866);
or U2947 (N_2947,N_2838,N_2820);
nand U2948 (N_2948,N_2836,N_2871);
xor U2949 (N_2949,N_2858,N_2839);
nand U2950 (N_2950,N_2881,N_2883);
or U2951 (N_2951,N_2828,N_2880);
nor U2952 (N_2952,N_2851,N_2858);
nor U2953 (N_2953,N_2877,N_2870);
and U2954 (N_2954,N_2813,N_2860);
and U2955 (N_2955,N_2849,N_2813);
and U2956 (N_2956,N_2866,N_2863);
and U2957 (N_2957,N_2894,N_2808);
and U2958 (N_2958,N_2875,N_2838);
xnor U2959 (N_2959,N_2816,N_2814);
or U2960 (N_2960,N_2817,N_2876);
or U2961 (N_2961,N_2884,N_2836);
nand U2962 (N_2962,N_2840,N_2842);
and U2963 (N_2963,N_2846,N_2806);
nor U2964 (N_2964,N_2848,N_2858);
and U2965 (N_2965,N_2861,N_2866);
or U2966 (N_2966,N_2834,N_2868);
nor U2967 (N_2967,N_2850,N_2898);
nand U2968 (N_2968,N_2818,N_2886);
nand U2969 (N_2969,N_2830,N_2828);
nor U2970 (N_2970,N_2811,N_2828);
nand U2971 (N_2971,N_2854,N_2813);
nand U2972 (N_2972,N_2814,N_2803);
and U2973 (N_2973,N_2851,N_2852);
or U2974 (N_2974,N_2839,N_2821);
nor U2975 (N_2975,N_2885,N_2844);
and U2976 (N_2976,N_2895,N_2852);
and U2977 (N_2977,N_2854,N_2829);
and U2978 (N_2978,N_2853,N_2897);
or U2979 (N_2979,N_2897,N_2836);
nand U2980 (N_2980,N_2821,N_2857);
nand U2981 (N_2981,N_2874,N_2883);
and U2982 (N_2982,N_2856,N_2849);
or U2983 (N_2983,N_2809,N_2874);
or U2984 (N_2984,N_2847,N_2858);
xor U2985 (N_2985,N_2835,N_2834);
and U2986 (N_2986,N_2860,N_2859);
nand U2987 (N_2987,N_2881,N_2885);
nand U2988 (N_2988,N_2891,N_2806);
nor U2989 (N_2989,N_2862,N_2854);
or U2990 (N_2990,N_2866,N_2832);
and U2991 (N_2991,N_2848,N_2870);
nand U2992 (N_2992,N_2893,N_2803);
nor U2993 (N_2993,N_2850,N_2809);
nor U2994 (N_2994,N_2851,N_2886);
and U2995 (N_2995,N_2856,N_2881);
nor U2996 (N_2996,N_2894,N_2816);
or U2997 (N_2997,N_2800,N_2834);
or U2998 (N_2998,N_2884,N_2814);
xnor U2999 (N_2999,N_2877,N_2895);
or UO_0 (O_0,N_2975,N_2979);
or UO_1 (O_1,N_2995,N_2906);
nand UO_2 (O_2,N_2940,N_2949);
or UO_3 (O_3,N_2938,N_2951);
nand UO_4 (O_4,N_2924,N_2976);
and UO_5 (O_5,N_2971,N_2939);
nor UO_6 (O_6,N_2933,N_2909);
and UO_7 (O_7,N_2968,N_2981);
or UO_8 (O_8,N_2988,N_2962);
and UO_9 (O_9,N_2918,N_2973);
nand UO_10 (O_10,N_2920,N_2930);
or UO_11 (O_11,N_2935,N_2901);
nor UO_12 (O_12,N_2946,N_2944);
nand UO_13 (O_13,N_2902,N_2982);
or UO_14 (O_14,N_2926,N_2903);
nor UO_15 (O_15,N_2934,N_2999);
nand UO_16 (O_16,N_2947,N_2991);
and UO_17 (O_17,N_2966,N_2974);
nor UO_18 (O_18,N_2956,N_2954);
nor UO_19 (O_19,N_2977,N_2916);
and UO_20 (O_20,N_2929,N_2928);
nand UO_21 (O_21,N_2927,N_2919);
and UO_22 (O_22,N_2969,N_2990);
and UO_23 (O_23,N_2952,N_2925);
nor UO_24 (O_24,N_2932,N_2972);
and UO_25 (O_25,N_2914,N_2987);
nand UO_26 (O_26,N_2986,N_2936);
nor UO_27 (O_27,N_2998,N_2942);
nor UO_28 (O_28,N_2955,N_2993);
nor UO_29 (O_29,N_2967,N_2958);
and UO_30 (O_30,N_2945,N_2941);
and UO_31 (O_31,N_2985,N_2989);
nor UO_32 (O_32,N_2915,N_2994);
and UO_33 (O_33,N_2917,N_2983);
nor UO_34 (O_34,N_2965,N_2960);
and UO_35 (O_35,N_2911,N_2912);
nor UO_36 (O_36,N_2923,N_2913);
and UO_37 (O_37,N_2970,N_2910);
nand UO_38 (O_38,N_2959,N_2908);
nand UO_39 (O_39,N_2980,N_2996);
or UO_40 (O_40,N_2904,N_2950);
nand UO_41 (O_41,N_2963,N_2953);
or UO_42 (O_42,N_2964,N_2907);
nor UO_43 (O_43,N_2943,N_2992);
nand UO_44 (O_44,N_2921,N_2961);
or UO_45 (O_45,N_2900,N_2922);
nand UO_46 (O_46,N_2957,N_2948);
nand UO_47 (O_47,N_2984,N_2931);
or UO_48 (O_48,N_2937,N_2997);
or UO_49 (O_49,N_2978,N_2905);
nand UO_50 (O_50,N_2987,N_2933);
or UO_51 (O_51,N_2905,N_2979);
or UO_52 (O_52,N_2901,N_2946);
xor UO_53 (O_53,N_2953,N_2965);
nand UO_54 (O_54,N_2998,N_2931);
nand UO_55 (O_55,N_2928,N_2901);
nor UO_56 (O_56,N_2970,N_2908);
xnor UO_57 (O_57,N_2956,N_2992);
nand UO_58 (O_58,N_2988,N_2932);
nand UO_59 (O_59,N_2997,N_2964);
nor UO_60 (O_60,N_2960,N_2909);
nand UO_61 (O_61,N_2994,N_2908);
nand UO_62 (O_62,N_2913,N_2994);
nor UO_63 (O_63,N_2985,N_2966);
or UO_64 (O_64,N_2902,N_2959);
or UO_65 (O_65,N_2993,N_2917);
or UO_66 (O_66,N_2965,N_2917);
and UO_67 (O_67,N_2929,N_2940);
and UO_68 (O_68,N_2912,N_2976);
or UO_69 (O_69,N_2966,N_2963);
nor UO_70 (O_70,N_2980,N_2975);
and UO_71 (O_71,N_2972,N_2944);
or UO_72 (O_72,N_2982,N_2948);
nor UO_73 (O_73,N_2910,N_2938);
nand UO_74 (O_74,N_2905,N_2958);
nand UO_75 (O_75,N_2982,N_2928);
and UO_76 (O_76,N_2932,N_2937);
or UO_77 (O_77,N_2914,N_2931);
and UO_78 (O_78,N_2912,N_2927);
nand UO_79 (O_79,N_2909,N_2987);
nor UO_80 (O_80,N_2992,N_2921);
nor UO_81 (O_81,N_2913,N_2973);
or UO_82 (O_82,N_2915,N_2985);
nor UO_83 (O_83,N_2901,N_2945);
nor UO_84 (O_84,N_2962,N_2946);
nor UO_85 (O_85,N_2932,N_2989);
or UO_86 (O_86,N_2989,N_2976);
nand UO_87 (O_87,N_2942,N_2908);
or UO_88 (O_88,N_2993,N_2903);
nand UO_89 (O_89,N_2990,N_2926);
or UO_90 (O_90,N_2925,N_2980);
or UO_91 (O_91,N_2945,N_2919);
and UO_92 (O_92,N_2941,N_2922);
xnor UO_93 (O_93,N_2984,N_2981);
or UO_94 (O_94,N_2994,N_2900);
nand UO_95 (O_95,N_2996,N_2909);
and UO_96 (O_96,N_2947,N_2985);
nand UO_97 (O_97,N_2998,N_2993);
or UO_98 (O_98,N_2941,N_2962);
nand UO_99 (O_99,N_2974,N_2957);
or UO_100 (O_100,N_2976,N_2903);
nor UO_101 (O_101,N_2964,N_2994);
and UO_102 (O_102,N_2942,N_2995);
nand UO_103 (O_103,N_2926,N_2928);
nor UO_104 (O_104,N_2919,N_2920);
nor UO_105 (O_105,N_2972,N_2930);
nand UO_106 (O_106,N_2900,N_2911);
nor UO_107 (O_107,N_2904,N_2985);
and UO_108 (O_108,N_2987,N_2956);
nand UO_109 (O_109,N_2968,N_2996);
and UO_110 (O_110,N_2901,N_2955);
or UO_111 (O_111,N_2920,N_2971);
nor UO_112 (O_112,N_2959,N_2931);
nand UO_113 (O_113,N_2953,N_2997);
nand UO_114 (O_114,N_2948,N_2931);
xnor UO_115 (O_115,N_2968,N_2924);
and UO_116 (O_116,N_2986,N_2948);
nor UO_117 (O_117,N_2920,N_2946);
nor UO_118 (O_118,N_2936,N_2947);
nor UO_119 (O_119,N_2983,N_2904);
or UO_120 (O_120,N_2900,N_2989);
or UO_121 (O_121,N_2983,N_2947);
xor UO_122 (O_122,N_2947,N_2923);
nor UO_123 (O_123,N_2913,N_2969);
nor UO_124 (O_124,N_2960,N_2971);
and UO_125 (O_125,N_2961,N_2979);
nand UO_126 (O_126,N_2932,N_2905);
xnor UO_127 (O_127,N_2977,N_2969);
nor UO_128 (O_128,N_2965,N_2950);
and UO_129 (O_129,N_2998,N_2976);
nor UO_130 (O_130,N_2933,N_2971);
and UO_131 (O_131,N_2916,N_2962);
nor UO_132 (O_132,N_2961,N_2954);
or UO_133 (O_133,N_2991,N_2965);
nor UO_134 (O_134,N_2903,N_2949);
nand UO_135 (O_135,N_2932,N_2987);
and UO_136 (O_136,N_2975,N_2961);
nor UO_137 (O_137,N_2950,N_2969);
or UO_138 (O_138,N_2980,N_2985);
nor UO_139 (O_139,N_2933,N_2984);
and UO_140 (O_140,N_2907,N_2979);
nor UO_141 (O_141,N_2925,N_2902);
and UO_142 (O_142,N_2995,N_2934);
xor UO_143 (O_143,N_2907,N_2981);
nand UO_144 (O_144,N_2991,N_2906);
nand UO_145 (O_145,N_2938,N_2908);
or UO_146 (O_146,N_2958,N_2969);
or UO_147 (O_147,N_2914,N_2909);
or UO_148 (O_148,N_2977,N_2918);
nand UO_149 (O_149,N_2910,N_2942);
or UO_150 (O_150,N_2918,N_2946);
or UO_151 (O_151,N_2909,N_2972);
or UO_152 (O_152,N_2988,N_2978);
or UO_153 (O_153,N_2916,N_2972);
and UO_154 (O_154,N_2993,N_2973);
or UO_155 (O_155,N_2926,N_2934);
and UO_156 (O_156,N_2976,N_2954);
or UO_157 (O_157,N_2969,N_2951);
or UO_158 (O_158,N_2935,N_2934);
and UO_159 (O_159,N_2959,N_2900);
nor UO_160 (O_160,N_2991,N_2972);
or UO_161 (O_161,N_2964,N_2987);
nand UO_162 (O_162,N_2926,N_2907);
and UO_163 (O_163,N_2959,N_2958);
nand UO_164 (O_164,N_2906,N_2964);
nand UO_165 (O_165,N_2953,N_2924);
nand UO_166 (O_166,N_2950,N_2927);
and UO_167 (O_167,N_2938,N_2954);
nor UO_168 (O_168,N_2921,N_2901);
and UO_169 (O_169,N_2945,N_2994);
and UO_170 (O_170,N_2909,N_2983);
nand UO_171 (O_171,N_2963,N_2983);
nor UO_172 (O_172,N_2993,N_2933);
and UO_173 (O_173,N_2998,N_2968);
and UO_174 (O_174,N_2927,N_2948);
nor UO_175 (O_175,N_2964,N_2967);
nor UO_176 (O_176,N_2946,N_2921);
nor UO_177 (O_177,N_2935,N_2979);
and UO_178 (O_178,N_2924,N_2994);
and UO_179 (O_179,N_2910,N_2903);
nand UO_180 (O_180,N_2958,N_2933);
and UO_181 (O_181,N_2938,N_2917);
or UO_182 (O_182,N_2992,N_2966);
nand UO_183 (O_183,N_2907,N_2984);
or UO_184 (O_184,N_2999,N_2910);
or UO_185 (O_185,N_2929,N_2997);
and UO_186 (O_186,N_2916,N_2945);
and UO_187 (O_187,N_2949,N_2966);
nand UO_188 (O_188,N_2982,N_2911);
and UO_189 (O_189,N_2959,N_2954);
nor UO_190 (O_190,N_2901,N_2911);
xnor UO_191 (O_191,N_2924,N_2993);
nor UO_192 (O_192,N_2951,N_2976);
nor UO_193 (O_193,N_2989,N_2991);
and UO_194 (O_194,N_2918,N_2965);
nand UO_195 (O_195,N_2914,N_2945);
or UO_196 (O_196,N_2963,N_2999);
and UO_197 (O_197,N_2921,N_2994);
or UO_198 (O_198,N_2916,N_2934);
nand UO_199 (O_199,N_2992,N_2970);
nor UO_200 (O_200,N_2936,N_2931);
or UO_201 (O_201,N_2918,N_2960);
or UO_202 (O_202,N_2928,N_2981);
nand UO_203 (O_203,N_2914,N_2980);
or UO_204 (O_204,N_2955,N_2935);
or UO_205 (O_205,N_2987,N_2921);
nor UO_206 (O_206,N_2981,N_2908);
xor UO_207 (O_207,N_2919,N_2903);
and UO_208 (O_208,N_2971,N_2921);
xnor UO_209 (O_209,N_2985,N_2951);
nor UO_210 (O_210,N_2973,N_2926);
or UO_211 (O_211,N_2964,N_2943);
or UO_212 (O_212,N_2939,N_2935);
nand UO_213 (O_213,N_2953,N_2970);
nand UO_214 (O_214,N_2950,N_2990);
nor UO_215 (O_215,N_2982,N_2914);
and UO_216 (O_216,N_2977,N_2975);
and UO_217 (O_217,N_2947,N_2921);
and UO_218 (O_218,N_2995,N_2968);
or UO_219 (O_219,N_2939,N_2913);
or UO_220 (O_220,N_2925,N_2946);
nor UO_221 (O_221,N_2996,N_2988);
nor UO_222 (O_222,N_2936,N_2911);
or UO_223 (O_223,N_2922,N_2909);
nand UO_224 (O_224,N_2950,N_2946);
or UO_225 (O_225,N_2952,N_2930);
nor UO_226 (O_226,N_2909,N_2910);
or UO_227 (O_227,N_2905,N_2974);
or UO_228 (O_228,N_2903,N_2954);
or UO_229 (O_229,N_2985,N_2984);
or UO_230 (O_230,N_2936,N_2914);
or UO_231 (O_231,N_2996,N_2977);
or UO_232 (O_232,N_2930,N_2993);
and UO_233 (O_233,N_2921,N_2966);
nor UO_234 (O_234,N_2943,N_2989);
nor UO_235 (O_235,N_2967,N_2974);
or UO_236 (O_236,N_2968,N_2915);
and UO_237 (O_237,N_2977,N_2982);
or UO_238 (O_238,N_2905,N_2955);
nand UO_239 (O_239,N_2958,N_2950);
nor UO_240 (O_240,N_2991,N_2918);
and UO_241 (O_241,N_2915,N_2981);
and UO_242 (O_242,N_2939,N_2986);
or UO_243 (O_243,N_2916,N_2990);
or UO_244 (O_244,N_2987,N_2954);
nor UO_245 (O_245,N_2905,N_2997);
and UO_246 (O_246,N_2991,N_2929);
and UO_247 (O_247,N_2949,N_2973);
nor UO_248 (O_248,N_2913,N_2975);
nand UO_249 (O_249,N_2930,N_2986);
nor UO_250 (O_250,N_2930,N_2917);
or UO_251 (O_251,N_2923,N_2972);
and UO_252 (O_252,N_2977,N_2960);
or UO_253 (O_253,N_2966,N_2989);
or UO_254 (O_254,N_2943,N_2909);
nor UO_255 (O_255,N_2995,N_2990);
or UO_256 (O_256,N_2988,N_2933);
nand UO_257 (O_257,N_2971,N_2905);
nor UO_258 (O_258,N_2925,N_2929);
and UO_259 (O_259,N_2943,N_2922);
nor UO_260 (O_260,N_2991,N_2930);
nor UO_261 (O_261,N_2974,N_2912);
nor UO_262 (O_262,N_2952,N_2906);
or UO_263 (O_263,N_2961,N_2908);
nor UO_264 (O_264,N_2989,N_2970);
nor UO_265 (O_265,N_2996,N_2985);
or UO_266 (O_266,N_2940,N_2980);
nand UO_267 (O_267,N_2997,N_2951);
nand UO_268 (O_268,N_2993,N_2982);
and UO_269 (O_269,N_2939,N_2944);
or UO_270 (O_270,N_2907,N_2987);
nand UO_271 (O_271,N_2984,N_2942);
nor UO_272 (O_272,N_2910,N_2986);
nand UO_273 (O_273,N_2914,N_2956);
and UO_274 (O_274,N_2977,N_2978);
and UO_275 (O_275,N_2991,N_2937);
or UO_276 (O_276,N_2916,N_2914);
and UO_277 (O_277,N_2986,N_2987);
nor UO_278 (O_278,N_2926,N_2978);
nor UO_279 (O_279,N_2913,N_2964);
nand UO_280 (O_280,N_2981,N_2983);
and UO_281 (O_281,N_2942,N_2957);
xor UO_282 (O_282,N_2917,N_2956);
or UO_283 (O_283,N_2914,N_2974);
and UO_284 (O_284,N_2977,N_2994);
and UO_285 (O_285,N_2968,N_2943);
nand UO_286 (O_286,N_2939,N_2966);
nor UO_287 (O_287,N_2928,N_2906);
or UO_288 (O_288,N_2933,N_2962);
and UO_289 (O_289,N_2974,N_2989);
xnor UO_290 (O_290,N_2964,N_2912);
and UO_291 (O_291,N_2921,N_2954);
or UO_292 (O_292,N_2951,N_2906);
nand UO_293 (O_293,N_2932,N_2943);
and UO_294 (O_294,N_2993,N_2906);
nor UO_295 (O_295,N_2941,N_2975);
and UO_296 (O_296,N_2973,N_2935);
nand UO_297 (O_297,N_2995,N_2909);
xor UO_298 (O_298,N_2981,N_2944);
and UO_299 (O_299,N_2953,N_2927);
nand UO_300 (O_300,N_2973,N_2908);
nor UO_301 (O_301,N_2939,N_2908);
or UO_302 (O_302,N_2916,N_2917);
nand UO_303 (O_303,N_2911,N_2914);
and UO_304 (O_304,N_2936,N_2925);
and UO_305 (O_305,N_2932,N_2939);
xnor UO_306 (O_306,N_2967,N_2995);
and UO_307 (O_307,N_2956,N_2919);
and UO_308 (O_308,N_2939,N_2910);
or UO_309 (O_309,N_2920,N_2994);
and UO_310 (O_310,N_2990,N_2973);
and UO_311 (O_311,N_2972,N_2996);
nor UO_312 (O_312,N_2962,N_2953);
or UO_313 (O_313,N_2975,N_2934);
xnor UO_314 (O_314,N_2952,N_2937);
nand UO_315 (O_315,N_2925,N_2913);
nand UO_316 (O_316,N_2937,N_2985);
nand UO_317 (O_317,N_2953,N_2977);
and UO_318 (O_318,N_2983,N_2960);
nand UO_319 (O_319,N_2924,N_2978);
nor UO_320 (O_320,N_2931,N_2977);
nor UO_321 (O_321,N_2951,N_2902);
or UO_322 (O_322,N_2930,N_2961);
nor UO_323 (O_323,N_2999,N_2975);
nor UO_324 (O_324,N_2951,N_2964);
nor UO_325 (O_325,N_2905,N_2943);
nor UO_326 (O_326,N_2986,N_2949);
nor UO_327 (O_327,N_2942,N_2922);
and UO_328 (O_328,N_2939,N_2958);
or UO_329 (O_329,N_2991,N_2985);
nor UO_330 (O_330,N_2945,N_2915);
nand UO_331 (O_331,N_2916,N_2975);
or UO_332 (O_332,N_2957,N_2920);
nand UO_333 (O_333,N_2945,N_2982);
nor UO_334 (O_334,N_2990,N_2945);
nor UO_335 (O_335,N_2923,N_2988);
nor UO_336 (O_336,N_2998,N_2906);
and UO_337 (O_337,N_2920,N_2955);
or UO_338 (O_338,N_2965,N_2928);
and UO_339 (O_339,N_2916,N_2996);
nor UO_340 (O_340,N_2936,N_2958);
nand UO_341 (O_341,N_2920,N_2984);
nor UO_342 (O_342,N_2964,N_2982);
and UO_343 (O_343,N_2901,N_2922);
nand UO_344 (O_344,N_2910,N_2971);
nand UO_345 (O_345,N_2951,N_2924);
and UO_346 (O_346,N_2956,N_2986);
nand UO_347 (O_347,N_2963,N_2949);
nor UO_348 (O_348,N_2990,N_2937);
or UO_349 (O_349,N_2924,N_2979);
nand UO_350 (O_350,N_2926,N_2977);
nor UO_351 (O_351,N_2953,N_2955);
nand UO_352 (O_352,N_2978,N_2982);
or UO_353 (O_353,N_2975,N_2972);
or UO_354 (O_354,N_2901,N_2963);
and UO_355 (O_355,N_2953,N_2904);
or UO_356 (O_356,N_2974,N_2993);
or UO_357 (O_357,N_2952,N_2916);
or UO_358 (O_358,N_2941,N_2998);
or UO_359 (O_359,N_2907,N_2991);
nand UO_360 (O_360,N_2980,N_2971);
nor UO_361 (O_361,N_2990,N_2961);
and UO_362 (O_362,N_2981,N_2982);
nor UO_363 (O_363,N_2976,N_2952);
nand UO_364 (O_364,N_2910,N_2992);
nand UO_365 (O_365,N_2923,N_2937);
or UO_366 (O_366,N_2943,N_2969);
and UO_367 (O_367,N_2947,N_2969);
nand UO_368 (O_368,N_2960,N_2963);
nand UO_369 (O_369,N_2923,N_2966);
or UO_370 (O_370,N_2972,N_2994);
nand UO_371 (O_371,N_2986,N_2955);
nor UO_372 (O_372,N_2997,N_2910);
nand UO_373 (O_373,N_2950,N_2978);
or UO_374 (O_374,N_2961,N_2960);
nor UO_375 (O_375,N_2928,N_2985);
xor UO_376 (O_376,N_2983,N_2968);
nor UO_377 (O_377,N_2937,N_2930);
and UO_378 (O_378,N_2964,N_2999);
xnor UO_379 (O_379,N_2927,N_2975);
nor UO_380 (O_380,N_2944,N_2943);
or UO_381 (O_381,N_2990,N_2996);
nand UO_382 (O_382,N_2905,N_2913);
or UO_383 (O_383,N_2970,N_2925);
or UO_384 (O_384,N_2993,N_2984);
nand UO_385 (O_385,N_2992,N_2974);
xor UO_386 (O_386,N_2961,N_2934);
nand UO_387 (O_387,N_2939,N_2907);
nor UO_388 (O_388,N_2934,N_2968);
nor UO_389 (O_389,N_2964,N_2920);
nor UO_390 (O_390,N_2967,N_2911);
nor UO_391 (O_391,N_2938,N_2913);
and UO_392 (O_392,N_2967,N_2902);
and UO_393 (O_393,N_2980,N_2955);
nand UO_394 (O_394,N_2975,N_2989);
and UO_395 (O_395,N_2980,N_2911);
and UO_396 (O_396,N_2988,N_2998);
nor UO_397 (O_397,N_2900,N_2906);
nor UO_398 (O_398,N_2916,N_2993);
and UO_399 (O_399,N_2961,N_2959);
or UO_400 (O_400,N_2959,N_2955);
nand UO_401 (O_401,N_2977,N_2986);
or UO_402 (O_402,N_2985,N_2987);
or UO_403 (O_403,N_2938,N_2918);
nand UO_404 (O_404,N_2987,N_2960);
nor UO_405 (O_405,N_2938,N_2967);
nor UO_406 (O_406,N_2990,N_2902);
and UO_407 (O_407,N_2952,N_2946);
nor UO_408 (O_408,N_2997,N_2977);
nand UO_409 (O_409,N_2995,N_2998);
nor UO_410 (O_410,N_2974,N_2928);
or UO_411 (O_411,N_2908,N_2983);
or UO_412 (O_412,N_2967,N_2975);
nor UO_413 (O_413,N_2985,N_2983);
or UO_414 (O_414,N_2955,N_2966);
nand UO_415 (O_415,N_2934,N_2946);
nand UO_416 (O_416,N_2945,N_2925);
nor UO_417 (O_417,N_2917,N_2928);
nor UO_418 (O_418,N_2939,N_2989);
or UO_419 (O_419,N_2982,N_2967);
or UO_420 (O_420,N_2993,N_2957);
or UO_421 (O_421,N_2967,N_2939);
or UO_422 (O_422,N_2928,N_2959);
nor UO_423 (O_423,N_2976,N_2964);
and UO_424 (O_424,N_2910,N_2916);
and UO_425 (O_425,N_2922,N_2985);
nand UO_426 (O_426,N_2999,N_2918);
and UO_427 (O_427,N_2979,N_2978);
or UO_428 (O_428,N_2916,N_2984);
nand UO_429 (O_429,N_2935,N_2952);
nand UO_430 (O_430,N_2986,N_2969);
nand UO_431 (O_431,N_2915,N_2901);
and UO_432 (O_432,N_2981,N_2954);
and UO_433 (O_433,N_2957,N_2967);
or UO_434 (O_434,N_2993,N_2915);
nand UO_435 (O_435,N_2958,N_2947);
or UO_436 (O_436,N_2968,N_2999);
nor UO_437 (O_437,N_2934,N_2933);
or UO_438 (O_438,N_2985,N_2938);
or UO_439 (O_439,N_2912,N_2910);
and UO_440 (O_440,N_2989,N_2961);
nor UO_441 (O_441,N_2918,N_2984);
or UO_442 (O_442,N_2928,N_2973);
or UO_443 (O_443,N_2907,N_2969);
or UO_444 (O_444,N_2900,N_2988);
nor UO_445 (O_445,N_2935,N_2942);
and UO_446 (O_446,N_2972,N_2940);
nor UO_447 (O_447,N_2917,N_2957);
nand UO_448 (O_448,N_2918,N_2970);
and UO_449 (O_449,N_2959,N_2921);
or UO_450 (O_450,N_2931,N_2911);
or UO_451 (O_451,N_2940,N_2941);
and UO_452 (O_452,N_2923,N_2989);
nor UO_453 (O_453,N_2992,N_2920);
and UO_454 (O_454,N_2962,N_2952);
xnor UO_455 (O_455,N_2998,N_2951);
nor UO_456 (O_456,N_2946,N_2916);
or UO_457 (O_457,N_2939,N_2911);
nor UO_458 (O_458,N_2944,N_2992);
and UO_459 (O_459,N_2926,N_2919);
nand UO_460 (O_460,N_2963,N_2944);
or UO_461 (O_461,N_2939,N_2970);
nor UO_462 (O_462,N_2983,N_2995);
and UO_463 (O_463,N_2972,N_2931);
and UO_464 (O_464,N_2916,N_2970);
nand UO_465 (O_465,N_2937,N_2904);
and UO_466 (O_466,N_2939,N_2995);
nand UO_467 (O_467,N_2934,N_2911);
and UO_468 (O_468,N_2978,N_2941);
and UO_469 (O_469,N_2969,N_2965);
nor UO_470 (O_470,N_2932,N_2963);
or UO_471 (O_471,N_2991,N_2986);
and UO_472 (O_472,N_2963,N_2903);
or UO_473 (O_473,N_2937,N_2939);
nand UO_474 (O_474,N_2952,N_2939);
nand UO_475 (O_475,N_2984,N_2923);
nor UO_476 (O_476,N_2974,N_2917);
nor UO_477 (O_477,N_2925,N_2953);
or UO_478 (O_478,N_2902,N_2950);
nor UO_479 (O_479,N_2919,N_2905);
or UO_480 (O_480,N_2905,N_2969);
nor UO_481 (O_481,N_2944,N_2987);
or UO_482 (O_482,N_2972,N_2902);
or UO_483 (O_483,N_2901,N_2944);
nor UO_484 (O_484,N_2907,N_2929);
xor UO_485 (O_485,N_2920,N_2943);
or UO_486 (O_486,N_2953,N_2947);
nor UO_487 (O_487,N_2938,N_2990);
or UO_488 (O_488,N_2932,N_2997);
and UO_489 (O_489,N_2975,N_2907);
and UO_490 (O_490,N_2929,N_2990);
or UO_491 (O_491,N_2920,N_2914);
nand UO_492 (O_492,N_2975,N_2996);
nand UO_493 (O_493,N_2999,N_2952);
or UO_494 (O_494,N_2975,N_2946);
or UO_495 (O_495,N_2903,N_2944);
xnor UO_496 (O_496,N_2937,N_2979);
nor UO_497 (O_497,N_2954,N_2917);
nand UO_498 (O_498,N_2911,N_2908);
or UO_499 (O_499,N_2930,N_2913);
endmodule