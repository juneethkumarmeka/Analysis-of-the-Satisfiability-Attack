module basic_500_3000_500_4_levels_2xor_3(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
nor U0 (N_0,In_398,In_366);
nor U1 (N_1,In_426,In_342);
and U2 (N_2,In_194,In_7);
and U3 (N_3,In_141,In_383);
nand U4 (N_4,In_328,In_369);
nor U5 (N_5,In_420,In_327);
nor U6 (N_6,In_213,In_298);
nand U7 (N_7,In_225,In_153);
nor U8 (N_8,In_46,In_283);
or U9 (N_9,In_21,In_181);
nand U10 (N_10,In_79,In_198);
or U11 (N_11,In_111,In_361);
nor U12 (N_12,In_215,In_95);
nand U13 (N_13,In_467,In_319);
nor U14 (N_14,In_97,In_156);
or U15 (N_15,In_349,In_86);
nand U16 (N_16,In_479,In_114);
nor U17 (N_17,In_131,In_78);
or U18 (N_18,In_202,In_435);
or U19 (N_19,In_295,In_494);
nor U20 (N_20,In_136,In_168);
nor U21 (N_21,In_178,In_191);
nor U22 (N_22,In_414,In_287);
nor U23 (N_23,In_105,In_499);
or U24 (N_24,In_119,In_363);
and U25 (N_25,In_2,In_410);
and U26 (N_26,In_443,In_336);
and U27 (N_27,In_109,In_474);
or U28 (N_28,In_101,In_135);
nor U29 (N_29,In_70,In_182);
or U30 (N_30,In_57,In_34);
or U31 (N_31,In_460,In_311);
nand U32 (N_32,In_160,In_1);
and U33 (N_33,In_271,In_388);
nor U34 (N_34,In_272,In_223);
nand U35 (N_35,In_227,In_496);
nand U36 (N_36,In_392,In_187);
nor U37 (N_37,In_158,In_84);
or U38 (N_38,In_347,In_453);
nor U39 (N_39,In_378,In_427);
nand U40 (N_40,In_416,In_415);
nor U41 (N_41,In_29,In_244);
nand U42 (N_42,In_399,In_455);
nand U43 (N_43,In_411,In_428);
nand U44 (N_44,In_192,In_273);
nand U45 (N_45,In_73,In_402);
nor U46 (N_46,In_441,In_102);
nor U47 (N_47,In_288,In_104);
or U48 (N_48,In_385,In_218);
xor U49 (N_49,In_165,In_395);
nor U50 (N_50,In_291,In_436);
nand U51 (N_51,In_330,In_169);
nor U52 (N_52,In_41,In_206);
nor U53 (N_53,In_275,In_180);
nand U54 (N_54,In_337,In_457);
or U55 (N_55,In_482,In_166);
nand U56 (N_56,In_140,In_210);
and U57 (N_57,In_468,In_471);
nand U58 (N_58,In_493,In_431);
nand U59 (N_59,In_144,In_299);
and U60 (N_60,In_310,In_412);
nor U61 (N_61,In_147,In_3);
nand U62 (N_62,In_315,In_145);
and U63 (N_63,In_237,In_294);
nand U64 (N_64,In_219,In_351);
and U65 (N_65,In_306,In_309);
nor U66 (N_66,In_449,In_464);
nor U67 (N_67,In_303,In_16);
or U68 (N_68,In_324,In_159);
and U69 (N_69,In_205,In_80);
and U70 (N_70,In_413,In_224);
and U71 (N_71,In_25,In_458);
nand U72 (N_72,In_157,In_430);
or U73 (N_73,In_495,In_130);
and U74 (N_74,In_233,In_172);
or U75 (N_75,In_382,In_148);
or U76 (N_76,In_329,In_211);
and U77 (N_77,In_459,In_312);
nand U78 (N_78,In_448,In_155);
xnor U79 (N_79,In_128,In_384);
and U80 (N_80,In_138,In_433);
and U81 (N_81,In_269,In_325);
and U82 (N_82,In_253,In_151);
nor U83 (N_83,In_407,In_56);
nor U84 (N_84,In_264,In_422);
nand U85 (N_85,In_132,In_401);
nor U86 (N_86,In_403,In_437);
and U87 (N_87,In_438,In_258);
or U88 (N_88,In_480,In_376);
nand U89 (N_89,In_174,In_440);
or U90 (N_90,In_9,In_353);
nand U91 (N_91,In_270,In_341);
and U92 (N_92,In_13,In_462);
xor U93 (N_93,In_381,In_344);
and U94 (N_94,In_456,In_374);
xor U95 (N_95,In_127,In_26);
or U96 (N_96,In_19,In_475);
and U97 (N_97,In_236,In_454);
nor U98 (N_98,In_358,In_217);
nand U99 (N_99,In_259,In_77);
nor U100 (N_100,In_76,In_339);
nand U101 (N_101,In_423,In_304);
nor U102 (N_102,In_20,In_164);
xnor U103 (N_103,In_72,In_481);
and U104 (N_104,In_31,In_118);
nand U105 (N_105,In_68,In_377);
and U106 (N_106,In_222,In_465);
and U107 (N_107,In_60,In_96);
nor U108 (N_108,In_445,In_55);
and U109 (N_109,In_397,In_90);
nand U110 (N_110,In_446,In_252);
nor U111 (N_111,In_150,In_92);
nand U112 (N_112,In_418,In_470);
nor U113 (N_113,In_340,In_207);
xnor U114 (N_114,In_333,In_359);
nor U115 (N_115,In_354,In_317);
nand U116 (N_116,In_11,In_254);
or U117 (N_117,In_279,In_195);
nor U118 (N_118,In_116,In_125);
and U119 (N_119,In_373,In_91);
and U120 (N_120,In_296,In_250);
and U121 (N_121,In_100,In_484);
or U122 (N_122,In_231,In_188);
and U123 (N_123,In_307,In_30);
or U124 (N_124,In_488,In_35);
or U125 (N_125,In_289,In_197);
or U126 (N_126,In_308,In_232);
and U127 (N_127,In_348,In_286);
nand U128 (N_128,In_320,In_274);
nand U129 (N_129,In_386,In_284);
nand U130 (N_130,In_99,In_408);
or U131 (N_131,In_85,In_472);
nor U132 (N_132,In_37,In_103);
or U133 (N_133,In_18,In_196);
nand U134 (N_134,In_44,In_380);
and U135 (N_135,In_214,In_24);
and U136 (N_136,In_0,In_47);
and U137 (N_137,In_62,In_179);
or U138 (N_138,In_300,In_246);
nand U139 (N_139,In_115,In_175);
or U140 (N_140,In_146,In_498);
or U141 (N_141,In_267,In_209);
and U142 (N_142,In_81,In_473);
nor U143 (N_143,In_265,In_266);
and U144 (N_144,In_372,In_282);
nor U145 (N_145,In_61,In_33);
or U146 (N_146,In_343,In_332);
nor U147 (N_147,In_38,In_45);
nand U148 (N_148,In_221,In_82);
nand U149 (N_149,In_362,In_83);
nand U150 (N_150,In_190,In_391);
nor U151 (N_151,In_208,In_15);
nand U152 (N_152,In_4,In_245);
nand U153 (N_153,In_58,In_421);
nor U154 (N_154,In_220,In_51);
and U155 (N_155,In_483,In_487);
nor U156 (N_156,In_429,In_5);
or U157 (N_157,In_120,In_485);
nor U158 (N_158,In_163,In_450);
and U159 (N_159,In_357,In_409);
nor U160 (N_160,In_491,In_256);
and U161 (N_161,In_352,In_27);
nand U162 (N_162,In_162,In_331);
or U163 (N_163,In_149,In_52);
nor U164 (N_164,In_404,In_370);
or U165 (N_165,In_368,In_261);
or U166 (N_166,In_356,In_490);
or U167 (N_167,In_154,In_117);
nand U168 (N_168,In_419,In_63);
nand U169 (N_169,In_238,In_134);
and U170 (N_170,In_387,In_177);
nand U171 (N_171,In_94,In_350);
or U172 (N_172,In_234,In_477);
or U173 (N_173,In_88,In_67);
or U174 (N_174,In_40,In_406);
nor U175 (N_175,In_365,In_439);
nor U176 (N_176,In_321,In_469);
or U177 (N_177,In_133,In_243);
or U178 (N_178,In_338,In_32);
and U179 (N_179,In_74,In_123);
nand U180 (N_180,In_476,In_121);
or U181 (N_181,In_452,In_186);
nor U182 (N_182,In_263,In_87);
or U183 (N_183,In_255,In_75);
and U184 (N_184,In_23,In_142);
or U185 (N_185,In_129,In_278);
nor U186 (N_186,In_36,In_49);
and U187 (N_187,In_48,In_65);
nand U188 (N_188,In_247,In_112);
nor U189 (N_189,In_39,In_447);
nand U190 (N_190,In_50,In_189);
or U191 (N_191,In_171,In_176);
xor U192 (N_192,In_152,In_98);
xor U193 (N_193,In_203,In_394);
nor U194 (N_194,In_110,In_239);
nor U195 (N_195,In_249,In_53);
nand U196 (N_196,In_405,In_322);
nor U197 (N_197,In_193,In_297);
and U198 (N_198,In_8,In_143);
or U199 (N_199,In_69,In_6);
nand U200 (N_200,In_451,In_290);
and U201 (N_201,In_400,In_285);
nor U202 (N_202,In_334,In_417);
nand U203 (N_203,In_242,In_241);
nor U204 (N_204,In_66,In_108);
or U205 (N_205,In_14,In_122);
and U206 (N_206,In_173,In_235);
nand U207 (N_207,In_89,In_42);
nand U208 (N_208,In_167,In_345);
and U209 (N_209,In_107,In_346);
or U210 (N_210,In_486,In_292);
nor U211 (N_211,In_126,In_22);
nor U212 (N_212,In_489,In_302);
and U213 (N_213,In_137,In_424);
and U214 (N_214,In_201,In_442);
or U215 (N_215,In_93,In_28);
nor U216 (N_216,In_161,In_314);
nand U217 (N_217,In_393,In_497);
nand U218 (N_218,In_248,In_113);
nand U219 (N_219,In_200,In_318);
nand U220 (N_220,In_228,In_281);
nor U221 (N_221,In_212,In_355);
and U222 (N_222,In_379,In_390);
nand U223 (N_223,In_371,In_17);
or U224 (N_224,In_184,In_199);
nor U225 (N_225,In_226,In_335);
nor U226 (N_226,In_396,In_316);
xor U227 (N_227,In_277,In_10);
nor U228 (N_228,In_323,In_478);
or U229 (N_229,In_257,In_59);
and U230 (N_230,In_367,In_185);
nor U231 (N_231,In_268,In_64);
or U232 (N_232,In_139,In_389);
nor U233 (N_233,In_375,In_106);
nor U234 (N_234,In_183,In_466);
xor U235 (N_235,In_276,In_251);
nand U236 (N_236,In_432,In_305);
nor U237 (N_237,In_240,In_293);
or U238 (N_238,In_313,In_364);
nand U239 (N_239,In_425,In_492);
nand U240 (N_240,In_229,In_463);
nand U241 (N_241,In_280,In_301);
nand U242 (N_242,In_54,In_262);
nand U243 (N_243,In_326,In_260);
and U244 (N_244,In_170,In_216);
nand U245 (N_245,In_12,In_43);
and U246 (N_246,In_461,In_230);
and U247 (N_247,In_360,In_434);
or U248 (N_248,In_124,In_444);
nand U249 (N_249,In_71,In_204);
or U250 (N_250,In_272,In_303);
xnor U251 (N_251,In_476,In_388);
or U252 (N_252,In_40,In_307);
and U253 (N_253,In_253,In_252);
and U254 (N_254,In_478,In_53);
nand U255 (N_255,In_428,In_265);
nand U256 (N_256,In_57,In_360);
nand U257 (N_257,In_64,In_460);
and U258 (N_258,In_56,In_211);
nor U259 (N_259,In_215,In_14);
and U260 (N_260,In_262,In_156);
nor U261 (N_261,In_210,In_228);
or U262 (N_262,In_483,In_495);
nor U263 (N_263,In_198,In_372);
and U264 (N_264,In_205,In_309);
nand U265 (N_265,In_163,In_458);
or U266 (N_266,In_185,In_265);
nand U267 (N_267,In_372,In_497);
or U268 (N_268,In_213,In_131);
or U269 (N_269,In_22,In_115);
or U270 (N_270,In_154,In_339);
nor U271 (N_271,In_104,In_499);
and U272 (N_272,In_127,In_115);
nand U273 (N_273,In_464,In_14);
nor U274 (N_274,In_259,In_406);
nor U275 (N_275,In_171,In_3);
nand U276 (N_276,In_473,In_69);
nand U277 (N_277,In_449,In_22);
and U278 (N_278,In_26,In_187);
nor U279 (N_279,In_287,In_481);
nand U280 (N_280,In_25,In_301);
or U281 (N_281,In_239,In_242);
and U282 (N_282,In_352,In_18);
nand U283 (N_283,In_291,In_77);
nor U284 (N_284,In_237,In_74);
xnor U285 (N_285,In_194,In_189);
nand U286 (N_286,In_18,In_186);
nor U287 (N_287,In_257,In_60);
and U288 (N_288,In_179,In_336);
or U289 (N_289,In_190,In_85);
nor U290 (N_290,In_493,In_24);
and U291 (N_291,In_79,In_206);
nor U292 (N_292,In_470,In_17);
nor U293 (N_293,In_69,In_293);
xnor U294 (N_294,In_333,In_250);
nand U295 (N_295,In_41,In_439);
nor U296 (N_296,In_191,In_292);
nand U297 (N_297,In_428,In_415);
or U298 (N_298,In_175,In_127);
nor U299 (N_299,In_493,In_94);
nand U300 (N_300,In_69,In_311);
or U301 (N_301,In_169,In_421);
xor U302 (N_302,In_226,In_208);
and U303 (N_303,In_498,In_92);
nand U304 (N_304,In_362,In_91);
or U305 (N_305,In_191,In_56);
nor U306 (N_306,In_358,In_364);
xor U307 (N_307,In_6,In_181);
nand U308 (N_308,In_177,In_295);
or U309 (N_309,In_393,In_265);
nand U310 (N_310,In_412,In_11);
and U311 (N_311,In_265,In_223);
nand U312 (N_312,In_216,In_267);
and U313 (N_313,In_83,In_235);
nor U314 (N_314,In_220,In_103);
nor U315 (N_315,In_476,In_432);
nor U316 (N_316,In_361,In_122);
nor U317 (N_317,In_231,In_368);
or U318 (N_318,In_134,In_77);
nor U319 (N_319,In_215,In_385);
and U320 (N_320,In_49,In_425);
or U321 (N_321,In_175,In_340);
or U322 (N_322,In_46,In_463);
xor U323 (N_323,In_452,In_209);
and U324 (N_324,In_168,In_10);
nor U325 (N_325,In_369,In_37);
or U326 (N_326,In_355,In_261);
nor U327 (N_327,In_146,In_224);
and U328 (N_328,In_114,In_377);
nor U329 (N_329,In_192,In_373);
or U330 (N_330,In_415,In_223);
nand U331 (N_331,In_171,In_409);
and U332 (N_332,In_362,In_20);
and U333 (N_333,In_183,In_182);
nand U334 (N_334,In_411,In_66);
nor U335 (N_335,In_47,In_433);
or U336 (N_336,In_225,In_403);
nand U337 (N_337,In_206,In_223);
or U338 (N_338,In_288,In_376);
and U339 (N_339,In_438,In_334);
or U340 (N_340,In_418,In_134);
nor U341 (N_341,In_95,In_257);
nand U342 (N_342,In_410,In_21);
and U343 (N_343,In_211,In_392);
nor U344 (N_344,In_65,In_324);
nor U345 (N_345,In_198,In_45);
and U346 (N_346,In_125,In_39);
nand U347 (N_347,In_185,In_397);
nand U348 (N_348,In_114,In_175);
and U349 (N_349,In_467,In_168);
or U350 (N_350,In_317,In_209);
and U351 (N_351,In_354,In_320);
nor U352 (N_352,In_348,In_342);
or U353 (N_353,In_229,In_413);
nor U354 (N_354,In_431,In_124);
and U355 (N_355,In_162,In_186);
and U356 (N_356,In_298,In_60);
or U357 (N_357,In_304,In_277);
nand U358 (N_358,In_404,In_122);
nor U359 (N_359,In_256,In_77);
nand U360 (N_360,In_135,In_434);
nand U361 (N_361,In_166,In_42);
or U362 (N_362,In_174,In_96);
nor U363 (N_363,In_443,In_437);
and U364 (N_364,In_348,In_312);
or U365 (N_365,In_23,In_480);
or U366 (N_366,In_107,In_287);
nand U367 (N_367,In_494,In_22);
or U368 (N_368,In_257,In_331);
xor U369 (N_369,In_110,In_25);
and U370 (N_370,In_174,In_496);
nand U371 (N_371,In_265,In_241);
or U372 (N_372,In_268,In_56);
nand U373 (N_373,In_66,In_30);
nand U374 (N_374,In_241,In_132);
nor U375 (N_375,In_327,In_95);
or U376 (N_376,In_26,In_471);
or U377 (N_377,In_426,In_496);
nor U378 (N_378,In_313,In_293);
or U379 (N_379,In_303,In_194);
nor U380 (N_380,In_187,In_181);
or U381 (N_381,In_304,In_406);
or U382 (N_382,In_420,In_494);
nor U383 (N_383,In_281,In_165);
or U384 (N_384,In_247,In_472);
nor U385 (N_385,In_412,In_53);
nand U386 (N_386,In_240,In_272);
nand U387 (N_387,In_334,In_139);
nor U388 (N_388,In_159,In_41);
or U389 (N_389,In_224,In_8);
or U390 (N_390,In_210,In_436);
and U391 (N_391,In_413,In_120);
nand U392 (N_392,In_254,In_461);
nand U393 (N_393,In_196,In_465);
nor U394 (N_394,In_309,In_361);
nor U395 (N_395,In_99,In_313);
nand U396 (N_396,In_114,In_58);
nand U397 (N_397,In_152,In_20);
nor U398 (N_398,In_409,In_121);
or U399 (N_399,In_369,In_32);
and U400 (N_400,In_174,In_460);
and U401 (N_401,In_170,In_63);
xor U402 (N_402,In_319,In_365);
and U403 (N_403,In_176,In_98);
nand U404 (N_404,In_331,In_322);
and U405 (N_405,In_362,In_395);
or U406 (N_406,In_142,In_397);
and U407 (N_407,In_478,In_175);
or U408 (N_408,In_372,In_208);
and U409 (N_409,In_200,In_288);
nand U410 (N_410,In_327,In_312);
nor U411 (N_411,In_464,In_496);
and U412 (N_412,In_249,In_226);
nor U413 (N_413,In_240,In_437);
and U414 (N_414,In_89,In_270);
nand U415 (N_415,In_135,In_202);
or U416 (N_416,In_54,In_309);
or U417 (N_417,In_254,In_106);
or U418 (N_418,In_280,In_217);
nor U419 (N_419,In_467,In_157);
and U420 (N_420,In_164,In_361);
nand U421 (N_421,In_76,In_219);
or U422 (N_422,In_375,In_337);
and U423 (N_423,In_486,In_156);
nand U424 (N_424,In_435,In_495);
or U425 (N_425,In_0,In_20);
or U426 (N_426,In_224,In_393);
nor U427 (N_427,In_323,In_139);
nor U428 (N_428,In_488,In_351);
nand U429 (N_429,In_91,In_23);
xor U430 (N_430,In_266,In_104);
or U431 (N_431,In_300,In_168);
nand U432 (N_432,In_445,In_311);
nor U433 (N_433,In_98,In_107);
and U434 (N_434,In_386,In_45);
and U435 (N_435,In_203,In_88);
nand U436 (N_436,In_135,In_389);
xor U437 (N_437,In_233,In_178);
or U438 (N_438,In_213,In_13);
nand U439 (N_439,In_69,In_491);
or U440 (N_440,In_212,In_346);
xor U441 (N_441,In_244,In_249);
nand U442 (N_442,In_262,In_58);
or U443 (N_443,In_258,In_88);
xor U444 (N_444,In_461,In_206);
nor U445 (N_445,In_288,In_64);
or U446 (N_446,In_110,In_206);
or U447 (N_447,In_223,In_175);
and U448 (N_448,In_216,In_255);
nand U449 (N_449,In_464,In_314);
or U450 (N_450,In_46,In_87);
and U451 (N_451,In_304,In_99);
nor U452 (N_452,In_277,In_45);
xor U453 (N_453,In_198,In_220);
or U454 (N_454,In_445,In_412);
nor U455 (N_455,In_159,In_391);
or U456 (N_456,In_119,In_472);
nand U457 (N_457,In_413,In_398);
nand U458 (N_458,In_331,In_495);
or U459 (N_459,In_347,In_380);
or U460 (N_460,In_478,In_409);
nor U461 (N_461,In_75,In_116);
nor U462 (N_462,In_84,In_295);
nor U463 (N_463,In_8,In_24);
nand U464 (N_464,In_290,In_213);
or U465 (N_465,In_130,In_207);
or U466 (N_466,In_191,In_153);
nand U467 (N_467,In_17,In_271);
nor U468 (N_468,In_486,In_490);
nand U469 (N_469,In_112,In_44);
or U470 (N_470,In_173,In_268);
or U471 (N_471,In_296,In_451);
nand U472 (N_472,In_299,In_490);
nor U473 (N_473,In_379,In_128);
nor U474 (N_474,In_498,In_477);
and U475 (N_475,In_210,In_104);
nand U476 (N_476,In_427,In_429);
xor U477 (N_477,In_72,In_202);
or U478 (N_478,In_95,In_318);
or U479 (N_479,In_177,In_416);
nand U480 (N_480,In_252,In_190);
nor U481 (N_481,In_118,In_91);
and U482 (N_482,In_423,In_48);
nand U483 (N_483,In_457,In_462);
and U484 (N_484,In_112,In_411);
or U485 (N_485,In_263,In_414);
and U486 (N_486,In_54,In_295);
nor U487 (N_487,In_281,In_289);
and U488 (N_488,In_188,In_369);
nor U489 (N_489,In_489,In_171);
nor U490 (N_490,In_18,In_329);
nor U491 (N_491,In_284,In_421);
nand U492 (N_492,In_489,In_169);
nand U493 (N_493,In_270,In_238);
nor U494 (N_494,In_262,In_371);
and U495 (N_495,In_327,In_371);
nor U496 (N_496,In_58,In_275);
nand U497 (N_497,In_364,In_187);
nand U498 (N_498,In_216,In_285);
nand U499 (N_499,In_486,In_455);
nor U500 (N_500,In_407,In_439);
or U501 (N_501,In_247,In_246);
xor U502 (N_502,In_119,In_57);
nor U503 (N_503,In_107,In_31);
and U504 (N_504,In_156,In_466);
nor U505 (N_505,In_227,In_86);
nor U506 (N_506,In_286,In_386);
and U507 (N_507,In_463,In_499);
and U508 (N_508,In_115,In_62);
nor U509 (N_509,In_321,In_490);
xnor U510 (N_510,In_139,In_466);
nand U511 (N_511,In_402,In_423);
or U512 (N_512,In_417,In_322);
nor U513 (N_513,In_431,In_54);
or U514 (N_514,In_220,In_340);
and U515 (N_515,In_253,In_30);
xor U516 (N_516,In_491,In_244);
nor U517 (N_517,In_355,In_59);
nor U518 (N_518,In_81,In_188);
nor U519 (N_519,In_71,In_296);
or U520 (N_520,In_458,In_167);
or U521 (N_521,In_85,In_141);
or U522 (N_522,In_474,In_438);
nor U523 (N_523,In_45,In_232);
nand U524 (N_524,In_288,In_197);
and U525 (N_525,In_241,In_191);
or U526 (N_526,In_269,In_116);
nand U527 (N_527,In_21,In_86);
and U528 (N_528,In_477,In_255);
nor U529 (N_529,In_26,In_202);
nand U530 (N_530,In_130,In_77);
nor U531 (N_531,In_114,In_77);
nand U532 (N_532,In_396,In_115);
nand U533 (N_533,In_44,In_496);
nor U534 (N_534,In_212,In_44);
xor U535 (N_535,In_28,In_110);
xnor U536 (N_536,In_427,In_400);
nor U537 (N_537,In_287,In_451);
or U538 (N_538,In_366,In_107);
or U539 (N_539,In_191,In_325);
and U540 (N_540,In_449,In_271);
nand U541 (N_541,In_207,In_269);
nor U542 (N_542,In_393,In_442);
nor U543 (N_543,In_78,In_372);
nand U544 (N_544,In_123,In_496);
or U545 (N_545,In_148,In_387);
or U546 (N_546,In_210,In_269);
nor U547 (N_547,In_279,In_359);
or U548 (N_548,In_244,In_0);
or U549 (N_549,In_20,In_377);
nand U550 (N_550,In_185,In_301);
nor U551 (N_551,In_486,In_218);
nand U552 (N_552,In_104,In_446);
nor U553 (N_553,In_116,In_165);
and U554 (N_554,In_239,In_328);
or U555 (N_555,In_35,In_432);
or U556 (N_556,In_54,In_112);
and U557 (N_557,In_161,In_420);
nand U558 (N_558,In_447,In_38);
and U559 (N_559,In_360,In_498);
nor U560 (N_560,In_73,In_10);
nand U561 (N_561,In_425,In_98);
and U562 (N_562,In_15,In_165);
nand U563 (N_563,In_467,In_232);
and U564 (N_564,In_64,In_201);
and U565 (N_565,In_365,In_350);
or U566 (N_566,In_121,In_282);
or U567 (N_567,In_299,In_376);
and U568 (N_568,In_333,In_152);
or U569 (N_569,In_14,In_348);
nand U570 (N_570,In_227,In_121);
or U571 (N_571,In_7,In_173);
xnor U572 (N_572,In_231,In_222);
and U573 (N_573,In_451,In_69);
nand U574 (N_574,In_231,In_451);
nor U575 (N_575,In_68,In_446);
nor U576 (N_576,In_203,In_265);
nand U577 (N_577,In_441,In_145);
nor U578 (N_578,In_147,In_269);
nor U579 (N_579,In_204,In_115);
nand U580 (N_580,In_258,In_451);
and U581 (N_581,In_446,In_177);
nor U582 (N_582,In_183,In_432);
and U583 (N_583,In_345,In_182);
nor U584 (N_584,In_29,In_20);
nand U585 (N_585,In_37,In_135);
and U586 (N_586,In_210,In_397);
nand U587 (N_587,In_484,In_335);
and U588 (N_588,In_278,In_238);
nor U589 (N_589,In_464,In_181);
nor U590 (N_590,In_256,In_46);
or U591 (N_591,In_428,In_340);
nand U592 (N_592,In_5,In_93);
and U593 (N_593,In_366,In_490);
nor U594 (N_594,In_142,In_441);
and U595 (N_595,In_2,In_495);
and U596 (N_596,In_56,In_46);
nand U597 (N_597,In_491,In_295);
or U598 (N_598,In_166,In_341);
nor U599 (N_599,In_354,In_7);
nor U600 (N_600,In_178,In_452);
or U601 (N_601,In_366,In_266);
nand U602 (N_602,In_269,In_360);
nand U603 (N_603,In_29,In_42);
and U604 (N_604,In_92,In_176);
and U605 (N_605,In_87,In_392);
or U606 (N_606,In_458,In_129);
or U607 (N_607,In_99,In_400);
nor U608 (N_608,In_3,In_5);
nor U609 (N_609,In_132,In_436);
and U610 (N_610,In_122,In_341);
nand U611 (N_611,In_494,In_292);
and U612 (N_612,In_176,In_67);
and U613 (N_613,In_438,In_0);
and U614 (N_614,In_350,In_289);
or U615 (N_615,In_487,In_460);
nand U616 (N_616,In_294,In_75);
nand U617 (N_617,In_389,In_253);
nor U618 (N_618,In_444,In_186);
nor U619 (N_619,In_136,In_213);
nand U620 (N_620,In_86,In_298);
and U621 (N_621,In_344,In_121);
nand U622 (N_622,In_478,In_200);
or U623 (N_623,In_485,In_81);
or U624 (N_624,In_339,In_402);
and U625 (N_625,In_233,In_261);
and U626 (N_626,In_177,In_202);
xor U627 (N_627,In_423,In_129);
or U628 (N_628,In_20,In_367);
and U629 (N_629,In_346,In_134);
and U630 (N_630,In_328,In_1);
nor U631 (N_631,In_267,In_129);
or U632 (N_632,In_312,In_337);
nor U633 (N_633,In_8,In_252);
and U634 (N_634,In_419,In_489);
and U635 (N_635,In_334,In_28);
and U636 (N_636,In_99,In_442);
nor U637 (N_637,In_381,In_23);
and U638 (N_638,In_6,In_378);
nor U639 (N_639,In_263,In_468);
nor U640 (N_640,In_61,In_250);
nand U641 (N_641,In_338,In_212);
nor U642 (N_642,In_403,In_325);
and U643 (N_643,In_152,In_445);
nand U644 (N_644,In_40,In_116);
or U645 (N_645,In_356,In_268);
or U646 (N_646,In_211,In_273);
xnor U647 (N_647,In_274,In_165);
nor U648 (N_648,In_267,In_384);
nand U649 (N_649,In_448,In_119);
xnor U650 (N_650,In_141,In_492);
or U651 (N_651,In_463,In_458);
and U652 (N_652,In_181,In_455);
or U653 (N_653,In_70,In_420);
nand U654 (N_654,In_28,In_337);
nand U655 (N_655,In_162,In_264);
or U656 (N_656,In_312,In_15);
and U657 (N_657,In_263,In_328);
or U658 (N_658,In_355,In_427);
nor U659 (N_659,In_481,In_271);
and U660 (N_660,In_23,In_158);
nand U661 (N_661,In_319,In_51);
nor U662 (N_662,In_164,In_85);
xnor U663 (N_663,In_318,In_19);
nor U664 (N_664,In_405,In_468);
nand U665 (N_665,In_9,In_202);
nand U666 (N_666,In_187,In_63);
nand U667 (N_667,In_58,In_307);
nor U668 (N_668,In_39,In_420);
and U669 (N_669,In_120,In_41);
and U670 (N_670,In_327,In_90);
nor U671 (N_671,In_327,In_242);
and U672 (N_672,In_344,In_6);
and U673 (N_673,In_94,In_70);
and U674 (N_674,In_171,In_45);
nor U675 (N_675,In_176,In_324);
or U676 (N_676,In_85,In_48);
nand U677 (N_677,In_343,In_215);
nor U678 (N_678,In_352,In_331);
and U679 (N_679,In_48,In_282);
or U680 (N_680,In_273,In_171);
and U681 (N_681,In_88,In_406);
nand U682 (N_682,In_43,In_65);
nor U683 (N_683,In_441,In_150);
and U684 (N_684,In_476,In_93);
nand U685 (N_685,In_155,In_221);
or U686 (N_686,In_358,In_371);
nand U687 (N_687,In_82,In_77);
xnor U688 (N_688,In_32,In_310);
nand U689 (N_689,In_284,In_263);
nand U690 (N_690,In_174,In_347);
nor U691 (N_691,In_67,In_78);
nor U692 (N_692,In_49,In_46);
nand U693 (N_693,In_27,In_376);
xnor U694 (N_694,In_81,In_292);
nor U695 (N_695,In_437,In_140);
and U696 (N_696,In_336,In_417);
and U697 (N_697,In_145,In_426);
or U698 (N_698,In_31,In_168);
nor U699 (N_699,In_179,In_438);
nor U700 (N_700,In_239,In_198);
or U701 (N_701,In_465,In_202);
or U702 (N_702,In_163,In_138);
or U703 (N_703,In_123,In_395);
and U704 (N_704,In_116,In_34);
xnor U705 (N_705,In_154,In_24);
or U706 (N_706,In_133,In_441);
and U707 (N_707,In_23,In_388);
nand U708 (N_708,In_177,In_443);
nand U709 (N_709,In_297,In_238);
or U710 (N_710,In_247,In_289);
and U711 (N_711,In_492,In_424);
or U712 (N_712,In_180,In_457);
and U713 (N_713,In_483,In_331);
nand U714 (N_714,In_47,In_428);
nor U715 (N_715,In_380,In_85);
nand U716 (N_716,In_81,In_323);
nor U717 (N_717,In_74,In_205);
nor U718 (N_718,In_373,In_33);
nand U719 (N_719,In_166,In_398);
or U720 (N_720,In_434,In_68);
nor U721 (N_721,In_88,In_229);
or U722 (N_722,In_133,In_302);
or U723 (N_723,In_199,In_116);
nor U724 (N_724,In_39,In_398);
nor U725 (N_725,In_158,In_492);
or U726 (N_726,In_34,In_88);
nand U727 (N_727,In_63,In_385);
nor U728 (N_728,In_447,In_474);
or U729 (N_729,In_351,In_328);
xor U730 (N_730,In_403,In_345);
nand U731 (N_731,In_464,In_421);
or U732 (N_732,In_175,In_142);
xnor U733 (N_733,In_430,In_466);
nand U734 (N_734,In_49,In_205);
and U735 (N_735,In_279,In_357);
nor U736 (N_736,In_476,In_421);
nor U737 (N_737,In_156,In_407);
and U738 (N_738,In_450,In_304);
or U739 (N_739,In_95,In_19);
nand U740 (N_740,In_353,In_68);
nor U741 (N_741,In_255,In_287);
or U742 (N_742,In_477,In_130);
nand U743 (N_743,In_131,In_35);
nor U744 (N_744,In_216,In_302);
or U745 (N_745,In_40,In_264);
nand U746 (N_746,In_286,In_446);
nand U747 (N_747,In_107,In_96);
nand U748 (N_748,In_463,In_6);
and U749 (N_749,In_467,In_394);
nand U750 (N_750,N_539,N_163);
or U751 (N_751,N_597,N_580);
and U752 (N_752,N_157,N_560);
or U753 (N_753,N_353,N_604);
xnor U754 (N_754,N_289,N_461);
nand U755 (N_755,N_142,N_508);
and U756 (N_756,N_374,N_527);
nand U757 (N_757,N_249,N_324);
or U758 (N_758,N_327,N_382);
or U759 (N_759,N_219,N_610);
and U760 (N_760,N_691,N_207);
and U761 (N_761,N_279,N_667);
and U762 (N_762,N_100,N_574);
and U763 (N_763,N_578,N_564);
and U764 (N_764,N_665,N_307);
nand U765 (N_765,N_136,N_350);
nand U766 (N_766,N_654,N_193);
or U767 (N_767,N_518,N_605);
and U768 (N_768,N_671,N_233);
and U769 (N_769,N_86,N_281);
nand U770 (N_770,N_134,N_402);
nor U771 (N_771,N_273,N_277);
and U772 (N_772,N_550,N_1);
nand U773 (N_773,N_436,N_173);
nand U774 (N_774,N_138,N_652);
or U775 (N_775,N_239,N_551);
or U776 (N_776,N_546,N_442);
and U777 (N_777,N_211,N_587);
or U778 (N_778,N_643,N_18);
or U779 (N_779,N_3,N_496);
or U780 (N_780,N_372,N_98);
nor U781 (N_781,N_416,N_745);
and U782 (N_782,N_127,N_76);
nand U783 (N_783,N_102,N_47);
nand U784 (N_784,N_521,N_480);
nand U785 (N_785,N_41,N_54);
and U786 (N_786,N_23,N_462);
nand U787 (N_787,N_51,N_79);
and U788 (N_788,N_427,N_81);
nor U789 (N_789,N_731,N_464);
nand U790 (N_790,N_433,N_63);
and U791 (N_791,N_391,N_642);
or U792 (N_792,N_56,N_232);
and U793 (N_793,N_257,N_178);
or U794 (N_794,N_721,N_202);
nand U795 (N_795,N_12,N_62);
and U796 (N_796,N_575,N_42);
or U797 (N_797,N_437,N_594);
or U798 (N_798,N_531,N_180);
or U799 (N_799,N_502,N_385);
and U800 (N_800,N_359,N_493);
nand U801 (N_801,N_48,N_445);
and U802 (N_802,N_245,N_241);
or U803 (N_803,N_150,N_318);
and U804 (N_804,N_291,N_513);
nor U805 (N_805,N_703,N_497);
and U806 (N_806,N_306,N_450);
and U807 (N_807,N_225,N_356);
or U808 (N_808,N_599,N_339);
and U809 (N_809,N_749,N_570);
and U810 (N_810,N_8,N_510);
nand U811 (N_811,N_485,N_203);
nor U812 (N_812,N_135,N_354);
and U813 (N_813,N_74,N_338);
nor U814 (N_814,N_617,N_545);
or U815 (N_815,N_528,N_10);
and U816 (N_816,N_495,N_524);
and U817 (N_817,N_700,N_558);
or U818 (N_818,N_105,N_491);
or U819 (N_819,N_315,N_224);
nor U820 (N_820,N_658,N_407);
nand U821 (N_821,N_607,N_474);
nand U822 (N_822,N_69,N_561);
and U823 (N_823,N_456,N_230);
and U824 (N_824,N_282,N_426);
nand U825 (N_825,N_99,N_168);
nand U826 (N_826,N_500,N_430);
nor U827 (N_827,N_261,N_598);
and U828 (N_828,N_89,N_195);
nand U829 (N_829,N_265,N_370);
nor U830 (N_830,N_419,N_670);
and U831 (N_831,N_409,N_67);
and U832 (N_832,N_97,N_35);
nand U833 (N_833,N_344,N_4);
nand U834 (N_834,N_727,N_748);
or U835 (N_835,N_144,N_68);
and U836 (N_836,N_538,N_470);
nand U837 (N_837,N_413,N_398);
nor U838 (N_838,N_634,N_153);
or U839 (N_839,N_701,N_130);
and U840 (N_840,N_141,N_638);
nand U841 (N_841,N_179,N_697);
or U842 (N_842,N_710,N_657);
and U843 (N_843,N_451,N_361);
or U844 (N_844,N_345,N_183);
nand U845 (N_845,N_684,N_739);
nor U846 (N_846,N_351,N_49);
nand U847 (N_847,N_468,N_504);
nand U848 (N_848,N_601,N_82);
and U849 (N_849,N_390,N_590);
nand U850 (N_850,N_275,N_449);
nand U851 (N_851,N_308,N_645);
or U852 (N_852,N_247,N_6);
or U853 (N_853,N_28,N_45);
and U854 (N_854,N_53,N_271);
or U855 (N_855,N_19,N_145);
nand U856 (N_856,N_268,N_228);
nor U857 (N_857,N_114,N_467);
nand U858 (N_858,N_522,N_88);
or U859 (N_859,N_91,N_322);
nor U860 (N_860,N_218,N_272);
xor U861 (N_861,N_278,N_412);
xnor U862 (N_862,N_17,N_429);
or U863 (N_863,N_410,N_443);
or U864 (N_864,N_131,N_623);
and U865 (N_865,N_613,N_536);
nor U866 (N_866,N_486,N_334);
or U867 (N_867,N_319,N_24);
and U868 (N_868,N_192,N_742);
and U869 (N_869,N_217,N_674);
or U870 (N_870,N_542,N_325);
or U871 (N_871,N_472,N_481);
or U872 (N_872,N_286,N_200);
nand U873 (N_873,N_428,N_579);
nand U874 (N_874,N_108,N_208);
nand U875 (N_875,N_596,N_563);
and U876 (N_876,N_566,N_270);
and U877 (N_877,N_376,N_688);
nor U878 (N_878,N_320,N_50);
and U879 (N_879,N_379,N_735);
or U880 (N_880,N_215,N_260);
and U881 (N_881,N_288,N_93);
or U882 (N_882,N_651,N_258);
nand U883 (N_883,N_117,N_543);
or U884 (N_884,N_120,N_169);
nor U885 (N_885,N_304,N_666);
nand U886 (N_886,N_389,N_661);
and U887 (N_887,N_300,N_75);
and U888 (N_888,N_123,N_59);
nor U889 (N_889,N_395,N_660);
nand U890 (N_890,N_582,N_712);
and U891 (N_891,N_348,N_65);
nand U892 (N_892,N_720,N_87);
or U893 (N_893,N_723,N_296);
or U894 (N_894,N_685,N_156);
and U895 (N_895,N_549,N_678);
nor U896 (N_896,N_186,N_699);
or U897 (N_897,N_534,N_212);
nor U898 (N_898,N_367,N_214);
nor U899 (N_899,N_31,N_559);
nor U900 (N_900,N_630,N_255);
or U901 (N_901,N_629,N_274);
nand U902 (N_902,N_583,N_515);
or U903 (N_903,N_83,N_611);
and U904 (N_904,N_44,N_591);
nand U905 (N_905,N_439,N_162);
and U906 (N_906,N_677,N_342);
nand U907 (N_907,N_305,N_511);
nand U908 (N_908,N_673,N_190);
nand U909 (N_909,N_741,N_175);
or U910 (N_910,N_205,N_680);
and U911 (N_911,N_718,N_418);
or U912 (N_912,N_440,N_73);
nand U913 (N_913,N_473,N_9);
nand U914 (N_914,N_593,N_541);
nand U915 (N_915,N_176,N_532);
and U916 (N_916,N_535,N_636);
or U917 (N_917,N_695,N_312);
and U918 (N_918,N_57,N_347);
nor U919 (N_919,N_111,N_196);
nor U920 (N_920,N_369,N_184);
nand U921 (N_921,N_469,N_119);
nor U922 (N_922,N_328,N_182);
and U923 (N_923,N_498,N_434);
nor U924 (N_924,N_103,N_240);
nor U925 (N_925,N_484,N_104);
or U926 (N_926,N_520,N_299);
or U927 (N_927,N_92,N_125);
nor U928 (N_928,N_415,N_447);
nand U929 (N_929,N_620,N_459);
or U930 (N_930,N_358,N_602);
and U931 (N_931,N_724,N_711);
or U932 (N_932,N_332,N_405);
nor U933 (N_933,N_95,N_106);
nand U934 (N_934,N_466,N_732);
nand U935 (N_935,N_519,N_706);
nor U936 (N_936,N_514,N_204);
nor U937 (N_937,N_113,N_687);
and U938 (N_938,N_646,N_301);
or U939 (N_939,N_734,N_383);
or U940 (N_940,N_375,N_487);
nand U941 (N_941,N_516,N_220);
nand U942 (N_942,N_309,N_198);
nand U943 (N_943,N_229,N_276);
or U944 (N_944,N_140,N_619);
and U945 (N_945,N_421,N_363);
or U946 (N_946,N_284,N_715);
nor U947 (N_947,N_562,N_606);
nor U948 (N_948,N_311,N_336);
or U949 (N_949,N_223,N_201);
nor U950 (N_950,N_115,N_483);
nand U951 (N_951,N_297,N_256);
nor U952 (N_952,N_635,N_29);
or U953 (N_953,N_171,N_343);
nand U954 (N_954,N_512,N_411);
or U955 (N_955,N_94,N_116);
nand U956 (N_956,N_717,N_235);
nand U957 (N_957,N_137,N_625);
and U958 (N_958,N_525,N_316);
nor U959 (N_959,N_733,N_244);
and U960 (N_960,N_185,N_553);
or U961 (N_961,N_631,N_747);
nor U962 (N_962,N_78,N_252);
nand U963 (N_963,N_709,N_213);
and U964 (N_964,N_431,N_80);
and U965 (N_965,N_124,N_592);
or U966 (N_966,N_38,N_565);
nand U967 (N_967,N_280,N_698);
or U968 (N_968,N_14,N_490);
nand U969 (N_969,N_554,N_321);
nand U970 (N_970,N_174,N_653);
nand U971 (N_971,N_21,N_238);
nand U972 (N_972,N_414,N_129);
nand U973 (N_973,N_346,N_32);
or U974 (N_974,N_37,N_571);
or U975 (N_975,N_567,N_373);
nand U976 (N_976,N_189,N_737);
nand U977 (N_977,N_393,N_530);
and U978 (N_978,N_614,N_479);
or U979 (N_979,N_454,N_659);
and U980 (N_980,N_509,N_11);
nand U981 (N_981,N_392,N_298);
nor U982 (N_982,N_302,N_632);
or U983 (N_983,N_128,N_387);
xor U984 (N_984,N_164,N_499);
or U985 (N_985,N_70,N_540);
or U986 (N_986,N_377,N_523);
nand U987 (N_987,N_452,N_705);
nand U988 (N_988,N_293,N_547);
or U989 (N_989,N_227,N_738);
or U990 (N_990,N_380,N_109);
nand U991 (N_991,N_259,N_595);
or U992 (N_992,N_664,N_209);
nand U993 (N_993,N_489,N_453);
nor U994 (N_994,N_696,N_133);
and U995 (N_995,N_641,N_242);
nor U996 (N_996,N_600,N_26);
nor U997 (N_997,N_647,N_526);
and U998 (N_998,N_39,N_585);
nor U999 (N_999,N_132,N_250);
nor U1000 (N_1000,N_690,N_573);
and U1001 (N_1001,N_406,N_682);
or U1002 (N_1002,N_719,N_126);
and U1003 (N_1003,N_702,N_725);
nor U1004 (N_1004,N_626,N_746);
or U1005 (N_1005,N_294,N_704);
nand U1006 (N_1006,N_388,N_736);
nor U1007 (N_1007,N_335,N_143);
nand U1008 (N_1008,N_581,N_234);
or U1009 (N_1009,N_283,N_556);
or U1010 (N_1010,N_586,N_378);
and U1011 (N_1011,N_187,N_170);
nand U1012 (N_1012,N_20,N_714);
and U1013 (N_1013,N_396,N_633);
or U1014 (N_1014,N_181,N_310);
and U1015 (N_1015,N_552,N_603);
nor U1016 (N_1016,N_381,N_161);
nand U1017 (N_1017,N_362,N_476);
nand U1018 (N_1018,N_399,N_455);
nor U1019 (N_1019,N_160,N_46);
nand U1020 (N_1020,N_77,N_609);
and U1021 (N_1021,N_615,N_649);
nand U1022 (N_1022,N_425,N_404);
nor U1023 (N_1023,N_713,N_668);
or U1024 (N_1024,N_222,N_326);
and U1025 (N_1025,N_15,N_13);
nand U1026 (N_1026,N_722,N_290);
or U1027 (N_1027,N_155,N_107);
xnor U1028 (N_1028,N_672,N_364);
and U1029 (N_1029,N_424,N_662);
and U1030 (N_1030,N_333,N_295);
nor U1031 (N_1031,N_533,N_423);
or U1032 (N_1032,N_612,N_84);
nand U1033 (N_1033,N_27,N_506);
or U1034 (N_1034,N_30,N_689);
nand U1035 (N_1035,N_122,N_269);
nor U1036 (N_1036,N_34,N_475);
xor U1037 (N_1037,N_165,N_401);
and U1038 (N_1038,N_448,N_25);
and U1039 (N_1039,N_492,N_708);
nor U1040 (N_1040,N_368,N_648);
nor U1041 (N_1041,N_314,N_251);
nand U1042 (N_1042,N_360,N_548);
or U1043 (N_1043,N_397,N_650);
and U1044 (N_1044,N_675,N_85);
nor U1045 (N_1045,N_726,N_730);
or U1046 (N_1046,N_177,N_66);
nand U1047 (N_1047,N_254,N_313);
nand U1048 (N_1048,N_569,N_655);
nor U1049 (N_1049,N_231,N_460);
and U1050 (N_1050,N_743,N_226);
nand U1051 (N_1051,N_457,N_151);
nand U1052 (N_1052,N_323,N_441);
nor U1053 (N_1053,N_216,N_477);
nand U1054 (N_1054,N_584,N_154);
or U1055 (N_1055,N_576,N_640);
nor U1056 (N_1056,N_96,N_471);
nor U1057 (N_1057,N_716,N_139);
and U1058 (N_1058,N_683,N_118);
and U1059 (N_1059,N_248,N_40);
nand U1060 (N_1060,N_331,N_110);
nor U1061 (N_1061,N_253,N_172);
nand U1062 (N_1062,N_679,N_210);
nand U1063 (N_1063,N_146,N_246);
nor U1064 (N_1064,N_588,N_420);
nor U1065 (N_1065,N_292,N_568);
nand U1066 (N_1066,N_60,N_707);
or U1067 (N_1067,N_158,N_2);
and U1068 (N_1068,N_221,N_121);
nand U1069 (N_1069,N_152,N_341);
nand U1070 (N_1070,N_400,N_693);
and U1071 (N_1071,N_494,N_0);
and U1072 (N_1072,N_644,N_616);
nand U1073 (N_1073,N_167,N_669);
and U1074 (N_1074,N_676,N_159);
or U1075 (N_1075,N_337,N_438);
nor U1076 (N_1076,N_465,N_384);
nor U1077 (N_1077,N_478,N_639);
or U1078 (N_1078,N_58,N_628);
and U1079 (N_1079,N_544,N_537);
nor U1080 (N_1080,N_728,N_744);
nor U1081 (N_1081,N_61,N_555);
nor U1082 (N_1082,N_637,N_112);
or U1083 (N_1083,N_237,N_267);
xor U1084 (N_1084,N_694,N_7);
or U1085 (N_1085,N_589,N_740);
or U1086 (N_1086,N_16,N_262);
or U1087 (N_1087,N_618,N_557);
or U1088 (N_1088,N_681,N_577);
nor U1089 (N_1089,N_529,N_501);
or U1090 (N_1090,N_355,N_352);
nor U1091 (N_1091,N_166,N_403);
nor U1092 (N_1092,N_446,N_52);
nor U1093 (N_1093,N_371,N_572);
xor U1094 (N_1094,N_357,N_394);
or U1095 (N_1095,N_36,N_317);
or U1096 (N_1096,N_488,N_287);
nor U1097 (N_1097,N_482,N_621);
nor U1098 (N_1098,N_71,N_622);
nand U1099 (N_1099,N_432,N_503);
nand U1100 (N_1100,N_148,N_101);
nand U1101 (N_1101,N_517,N_417);
nand U1102 (N_1102,N_458,N_266);
nor U1103 (N_1103,N_303,N_149);
or U1104 (N_1104,N_22,N_624);
and U1105 (N_1105,N_663,N_366);
and U1106 (N_1106,N_5,N_507);
nand U1107 (N_1107,N_197,N_72);
and U1108 (N_1108,N_692,N_627);
nand U1109 (N_1109,N_194,N_191);
nor U1110 (N_1110,N_206,N_188);
nor U1111 (N_1111,N_340,N_608);
and U1112 (N_1112,N_33,N_408);
nor U1113 (N_1113,N_505,N_422);
or U1114 (N_1114,N_729,N_463);
nand U1115 (N_1115,N_199,N_264);
xor U1116 (N_1116,N_365,N_243);
nor U1117 (N_1117,N_330,N_43);
or U1118 (N_1118,N_55,N_263);
nor U1119 (N_1119,N_686,N_656);
and U1120 (N_1120,N_64,N_147);
nand U1121 (N_1121,N_444,N_90);
or U1122 (N_1122,N_329,N_386);
or U1123 (N_1123,N_236,N_349);
nor U1124 (N_1124,N_435,N_285);
and U1125 (N_1125,N_482,N_369);
nand U1126 (N_1126,N_528,N_379);
nand U1127 (N_1127,N_654,N_125);
or U1128 (N_1128,N_35,N_640);
nor U1129 (N_1129,N_295,N_657);
or U1130 (N_1130,N_78,N_365);
or U1131 (N_1131,N_18,N_548);
nand U1132 (N_1132,N_514,N_400);
and U1133 (N_1133,N_521,N_182);
nor U1134 (N_1134,N_147,N_216);
or U1135 (N_1135,N_168,N_431);
and U1136 (N_1136,N_510,N_5);
and U1137 (N_1137,N_222,N_145);
and U1138 (N_1138,N_141,N_349);
and U1139 (N_1139,N_322,N_95);
and U1140 (N_1140,N_82,N_141);
nand U1141 (N_1141,N_64,N_249);
nand U1142 (N_1142,N_488,N_444);
nor U1143 (N_1143,N_719,N_688);
or U1144 (N_1144,N_585,N_292);
nor U1145 (N_1145,N_237,N_580);
and U1146 (N_1146,N_142,N_110);
or U1147 (N_1147,N_626,N_719);
nor U1148 (N_1148,N_738,N_114);
nor U1149 (N_1149,N_700,N_281);
nor U1150 (N_1150,N_713,N_307);
and U1151 (N_1151,N_671,N_64);
nand U1152 (N_1152,N_189,N_445);
nand U1153 (N_1153,N_536,N_249);
nor U1154 (N_1154,N_313,N_294);
nor U1155 (N_1155,N_559,N_302);
and U1156 (N_1156,N_304,N_556);
and U1157 (N_1157,N_298,N_481);
nand U1158 (N_1158,N_74,N_732);
or U1159 (N_1159,N_258,N_282);
or U1160 (N_1160,N_160,N_706);
and U1161 (N_1161,N_32,N_322);
nor U1162 (N_1162,N_105,N_258);
nand U1163 (N_1163,N_375,N_185);
or U1164 (N_1164,N_323,N_676);
and U1165 (N_1165,N_651,N_680);
and U1166 (N_1166,N_689,N_58);
nor U1167 (N_1167,N_580,N_362);
and U1168 (N_1168,N_360,N_265);
or U1169 (N_1169,N_185,N_510);
nand U1170 (N_1170,N_700,N_712);
or U1171 (N_1171,N_409,N_5);
nor U1172 (N_1172,N_303,N_452);
nand U1173 (N_1173,N_499,N_18);
nand U1174 (N_1174,N_552,N_623);
nor U1175 (N_1175,N_651,N_429);
nor U1176 (N_1176,N_322,N_452);
xor U1177 (N_1177,N_616,N_727);
or U1178 (N_1178,N_615,N_73);
or U1179 (N_1179,N_382,N_747);
nor U1180 (N_1180,N_744,N_177);
nor U1181 (N_1181,N_166,N_423);
nor U1182 (N_1182,N_703,N_577);
xor U1183 (N_1183,N_190,N_139);
xor U1184 (N_1184,N_609,N_138);
and U1185 (N_1185,N_724,N_92);
and U1186 (N_1186,N_28,N_171);
or U1187 (N_1187,N_143,N_548);
or U1188 (N_1188,N_418,N_633);
nor U1189 (N_1189,N_14,N_312);
xor U1190 (N_1190,N_289,N_442);
or U1191 (N_1191,N_605,N_614);
nor U1192 (N_1192,N_57,N_152);
or U1193 (N_1193,N_598,N_710);
and U1194 (N_1194,N_692,N_218);
or U1195 (N_1195,N_147,N_663);
nand U1196 (N_1196,N_483,N_690);
and U1197 (N_1197,N_658,N_435);
nor U1198 (N_1198,N_586,N_63);
nor U1199 (N_1199,N_17,N_597);
or U1200 (N_1200,N_425,N_553);
and U1201 (N_1201,N_488,N_560);
or U1202 (N_1202,N_376,N_132);
or U1203 (N_1203,N_559,N_734);
and U1204 (N_1204,N_558,N_664);
or U1205 (N_1205,N_169,N_107);
nand U1206 (N_1206,N_156,N_387);
and U1207 (N_1207,N_736,N_289);
or U1208 (N_1208,N_245,N_517);
nor U1209 (N_1209,N_382,N_342);
or U1210 (N_1210,N_39,N_396);
nor U1211 (N_1211,N_288,N_230);
and U1212 (N_1212,N_453,N_747);
or U1213 (N_1213,N_195,N_396);
and U1214 (N_1214,N_618,N_75);
nor U1215 (N_1215,N_151,N_306);
or U1216 (N_1216,N_24,N_177);
nor U1217 (N_1217,N_740,N_446);
nand U1218 (N_1218,N_207,N_190);
nand U1219 (N_1219,N_318,N_274);
and U1220 (N_1220,N_518,N_329);
and U1221 (N_1221,N_657,N_88);
xnor U1222 (N_1222,N_66,N_694);
and U1223 (N_1223,N_355,N_414);
or U1224 (N_1224,N_257,N_283);
or U1225 (N_1225,N_558,N_681);
nand U1226 (N_1226,N_332,N_647);
nand U1227 (N_1227,N_416,N_480);
nor U1228 (N_1228,N_56,N_678);
nand U1229 (N_1229,N_227,N_245);
and U1230 (N_1230,N_442,N_17);
nand U1231 (N_1231,N_697,N_305);
and U1232 (N_1232,N_61,N_110);
and U1233 (N_1233,N_362,N_441);
nor U1234 (N_1234,N_504,N_62);
or U1235 (N_1235,N_359,N_552);
or U1236 (N_1236,N_531,N_578);
and U1237 (N_1237,N_625,N_571);
nand U1238 (N_1238,N_295,N_527);
nand U1239 (N_1239,N_50,N_271);
nor U1240 (N_1240,N_637,N_656);
and U1241 (N_1241,N_643,N_586);
and U1242 (N_1242,N_530,N_413);
and U1243 (N_1243,N_477,N_278);
nor U1244 (N_1244,N_371,N_97);
nor U1245 (N_1245,N_316,N_624);
and U1246 (N_1246,N_60,N_368);
nand U1247 (N_1247,N_739,N_180);
nor U1248 (N_1248,N_559,N_103);
or U1249 (N_1249,N_62,N_197);
nor U1250 (N_1250,N_83,N_22);
nor U1251 (N_1251,N_224,N_144);
nand U1252 (N_1252,N_234,N_214);
nand U1253 (N_1253,N_598,N_354);
or U1254 (N_1254,N_264,N_217);
nand U1255 (N_1255,N_352,N_383);
and U1256 (N_1256,N_10,N_169);
or U1257 (N_1257,N_630,N_483);
or U1258 (N_1258,N_147,N_223);
or U1259 (N_1259,N_56,N_694);
or U1260 (N_1260,N_44,N_190);
or U1261 (N_1261,N_14,N_143);
nor U1262 (N_1262,N_681,N_425);
and U1263 (N_1263,N_519,N_695);
or U1264 (N_1264,N_548,N_242);
nand U1265 (N_1265,N_554,N_77);
or U1266 (N_1266,N_586,N_263);
and U1267 (N_1267,N_364,N_602);
or U1268 (N_1268,N_92,N_686);
or U1269 (N_1269,N_311,N_162);
nand U1270 (N_1270,N_577,N_613);
nand U1271 (N_1271,N_51,N_695);
or U1272 (N_1272,N_161,N_204);
or U1273 (N_1273,N_174,N_659);
and U1274 (N_1274,N_425,N_560);
nor U1275 (N_1275,N_736,N_339);
nor U1276 (N_1276,N_28,N_534);
or U1277 (N_1277,N_368,N_643);
or U1278 (N_1278,N_241,N_11);
or U1279 (N_1279,N_267,N_343);
nand U1280 (N_1280,N_22,N_257);
or U1281 (N_1281,N_352,N_362);
nor U1282 (N_1282,N_193,N_381);
nor U1283 (N_1283,N_232,N_634);
or U1284 (N_1284,N_389,N_221);
and U1285 (N_1285,N_686,N_105);
or U1286 (N_1286,N_59,N_666);
or U1287 (N_1287,N_243,N_610);
nand U1288 (N_1288,N_695,N_53);
nand U1289 (N_1289,N_52,N_578);
or U1290 (N_1290,N_256,N_17);
or U1291 (N_1291,N_41,N_317);
nand U1292 (N_1292,N_431,N_357);
nand U1293 (N_1293,N_33,N_655);
and U1294 (N_1294,N_319,N_274);
nand U1295 (N_1295,N_381,N_439);
xor U1296 (N_1296,N_50,N_645);
and U1297 (N_1297,N_747,N_100);
nor U1298 (N_1298,N_325,N_404);
nand U1299 (N_1299,N_586,N_402);
or U1300 (N_1300,N_491,N_498);
or U1301 (N_1301,N_201,N_700);
and U1302 (N_1302,N_176,N_397);
and U1303 (N_1303,N_488,N_416);
nor U1304 (N_1304,N_492,N_620);
xnor U1305 (N_1305,N_380,N_286);
and U1306 (N_1306,N_565,N_296);
and U1307 (N_1307,N_52,N_636);
nand U1308 (N_1308,N_372,N_197);
nand U1309 (N_1309,N_507,N_302);
or U1310 (N_1310,N_398,N_697);
or U1311 (N_1311,N_19,N_549);
nand U1312 (N_1312,N_265,N_155);
nand U1313 (N_1313,N_142,N_356);
or U1314 (N_1314,N_202,N_148);
nand U1315 (N_1315,N_442,N_135);
and U1316 (N_1316,N_296,N_411);
nand U1317 (N_1317,N_211,N_563);
nor U1318 (N_1318,N_19,N_563);
nand U1319 (N_1319,N_680,N_179);
and U1320 (N_1320,N_730,N_365);
nor U1321 (N_1321,N_527,N_288);
and U1322 (N_1322,N_438,N_43);
nand U1323 (N_1323,N_145,N_24);
xor U1324 (N_1324,N_462,N_699);
nand U1325 (N_1325,N_643,N_632);
nand U1326 (N_1326,N_222,N_161);
and U1327 (N_1327,N_491,N_523);
nand U1328 (N_1328,N_581,N_212);
or U1329 (N_1329,N_408,N_604);
nand U1330 (N_1330,N_321,N_382);
nand U1331 (N_1331,N_485,N_269);
or U1332 (N_1332,N_377,N_329);
nand U1333 (N_1333,N_9,N_322);
and U1334 (N_1334,N_679,N_314);
nand U1335 (N_1335,N_653,N_217);
and U1336 (N_1336,N_608,N_153);
nand U1337 (N_1337,N_692,N_206);
or U1338 (N_1338,N_373,N_165);
and U1339 (N_1339,N_640,N_215);
or U1340 (N_1340,N_607,N_654);
nand U1341 (N_1341,N_467,N_602);
nor U1342 (N_1342,N_515,N_685);
nand U1343 (N_1343,N_607,N_74);
or U1344 (N_1344,N_82,N_41);
or U1345 (N_1345,N_395,N_185);
nand U1346 (N_1346,N_159,N_716);
or U1347 (N_1347,N_687,N_212);
nand U1348 (N_1348,N_266,N_171);
nand U1349 (N_1349,N_278,N_289);
nor U1350 (N_1350,N_177,N_656);
and U1351 (N_1351,N_378,N_631);
or U1352 (N_1352,N_54,N_71);
nor U1353 (N_1353,N_498,N_558);
nand U1354 (N_1354,N_336,N_398);
and U1355 (N_1355,N_169,N_738);
nor U1356 (N_1356,N_100,N_333);
nand U1357 (N_1357,N_538,N_273);
or U1358 (N_1358,N_405,N_642);
and U1359 (N_1359,N_628,N_268);
or U1360 (N_1360,N_259,N_747);
and U1361 (N_1361,N_468,N_370);
or U1362 (N_1362,N_575,N_681);
nor U1363 (N_1363,N_168,N_458);
nor U1364 (N_1364,N_110,N_301);
nor U1365 (N_1365,N_136,N_202);
nor U1366 (N_1366,N_413,N_362);
nand U1367 (N_1367,N_418,N_81);
nor U1368 (N_1368,N_536,N_554);
or U1369 (N_1369,N_34,N_699);
and U1370 (N_1370,N_360,N_614);
nor U1371 (N_1371,N_54,N_674);
and U1372 (N_1372,N_219,N_27);
nor U1373 (N_1373,N_385,N_164);
and U1374 (N_1374,N_185,N_493);
nor U1375 (N_1375,N_608,N_48);
nand U1376 (N_1376,N_705,N_522);
and U1377 (N_1377,N_85,N_238);
nand U1378 (N_1378,N_499,N_663);
nand U1379 (N_1379,N_730,N_554);
or U1380 (N_1380,N_654,N_288);
nor U1381 (N_1381,N_544,N_723);
nand U1382 (N_1382,N_599,N_221);
nand U1383 (N_1383,N_339,N_232);
nand U1384 (N_1384,N_132,N_540);
nor U1385 (N_1385,N_552,N_638);
or U1386 (N_1386,N_83,N_135);
or U1387 (N_1387,N_112,N_671);
or U1388 (N_1388,N_644,N_741);
nand U1389 (N_1389,N_64,N_721);
nor U1390 (N_1390,N_446,N_90);
or U1391 (N_1391,N_748,N_371);
nand U1392 (N_1392,N_679,N_404);
or U1393 (N_1393,N_458,N_563);
nand U1394 (N_1394,N_187,N_647);
nand U1395 (N_1395,N_213,N_476);
nand U1396 (N_1396,N_375,N_479);
nand U1397 (N_1397,N_202,N_274);
nor U1398 (N_1398,N_424,N_523);
nor U1399 (N_1399,N_139,N_335);
nand U1400 (N_1400,N_699,N_377);
nand U1401 (N_1401,N_589,N_153);
or U1402 (N_1402,N_83,N_534);
or U1403 (N_1403,N_2,N_21);
or U1404 (N_1404,N_375,N_271);
nand U1405 (N_1405,N_2,N_91);
or U1406 (N_1406,N_28,N_273);
or U1407 (N_1407,N_326,N_547);
or U1408 (N_1408,N_437,N_320);
and U1409 (N_1409,N_232,N_180);
nor U1410 (N_1410,N_491,N_361);
nor U1411 (N_1411,N_85,N_331);
nand U1412 (N_1412,N_114,N_162);
and U1413 (N_1413,N_150,N_115);
nor U1414 (N_1414,N_732,N_226);
nand U1415 (N_1415,N_497,N_249);
nor U1416 (N_1416,N_81,N_632);
nand U1417 (N_1417,N_194,N_307);
nand U1418 (N_1418,N_345,N_355);
nor U1419 (N_1419,N_352,N_587);
nor U1420 (N_1420,N_550,N_567);
or U1421 (N_1421,N_377,N_105);
or U1422 (N_1422,N_244,N_425);
and U1423 (N_1423,N_280,N_369);
nand U1424 (N_1424,N_20,N_275);
or U1425 (N_1425,N_105,N_699);
and U1426 (N_1426,N_217,N_361);
or U1427 (N_1427,N_215,N_666);
nand U1428 (N_1428,N_517,N_182);
or U1429 (N_1429,N_236,N_674);
nand U1430 (N_1430,N_364,N_315);
nor U1431 (N_1431,N_566,N_526);
and U1432 (N_1432,N_671,N_345);
or U1433 (N_1433,N_445,N_203);
and U1434 (N_1434,N_283,N_468);
nand U1435 (N_1435,N_105,N_338);
xnor U1436 (N_1436,N_274,N_196);
nor U1437 (N_1437,N_450,N_195);
nand U1438 (N_1438,N_338,N_627);
nor U1439 (N_1439,N_621,N_562);
nor U1440 (N_1440,N_434,N_647);
nor U1441 (N_1441,N_2,N_479);
nand U1442 (N_1442,N_563,N_440);
nor U1443 (N_1443,N_180,N_603);
and U1444 (N_1444,N_706,N_170);
and U1445 (N_1445,N_312,N_252);
nor U1446 (N_1446,N_66,N_356);
and U1447 (N_1447,N_242,N_197);
nor U1448 (N_1448,N_156,N_579);
nor U1449 (N_1449,N_455,N_538);
or U1450 (N_1450,N_88,N_531);
or U1451 (N_1451,N_488,N_741);
nor U1452 (N_1452,N_250,N_735);
and U1453 (N_1453,N_591,N_592);
and U1454 (N_1454,N_154,N_703);
nand U1455 (N_1455,N_467,N_311);
and U1456 (N_1456,N_399,N_137);
and U1457 (N_1457,N_657,N_221);
and U1458 (N_1458,N_564,N_28);
xnor U1459 (N_1459,N_522,N_469);
nor U1460 (N_1460,N_376,N_691);
nor U1461 (N_1461,N_305,N_439);
and U1462 (N_1462,N_176,N_521);
and U1463 (N_1463,N_109,N_728);
and U1464 (N_1464,N_561,N_599);
or U1465 (N_1465,N_721,N_289);
nand U1466 (N_1466,N_116,N_674);
nor U1467 (N_1467,N_604,N_289);
nand U1468 (N_1468,N_697,N_92);
nor U1469 (N_1469,N_516,N_159);
nor U1470 (N_1470,N_363,N_689);
or U1471 (N_1471,N_633,N_117);
or U1472 (N_1472,N_513,N_403);
or U1473 (N_1473,N_139,N_396);
and U1474 (N_1474,N_386,N_45);
nand U1475 (N_1475,N_178,N_700);
nor U1476 (N_1476,N_11,N_82);
or U1477 (N_1477,N_550,N_179);
or U1478 (N_1478,N_639,N_20);
and U1479 (N_1479,N_44,N_1);
and U1480 (N_1480,N_653,N_645);
nand U1481 (N_1481,N_45,N_542);
or U1482 (N_1482,N_537,N_585);
nand U1483 (N_1483,N_547,N_168);
nand U1484 (N_1484,N_490,N_126);
or U1485 (N_1485,N_176,N_526);
and U1486 (N_1486,N_33,N_713);
nand U1487 (N_1487,N_13,N_721);
and U1488 (N_1488,N_646,N_713);
nor U1489 (N_1489,N_561,N_256);
and U1490 (N_1490,N_348,N_96);
or U1491 (N_1491,N_66,N_458);
nand U1492 (N_1492,N_136,N_443);
and U1493 (N_1493,N_568,N_7);
or U1494 (N_1494,N_41,N_390);
nand U1495 (N_1495,N_707,N_592);
or U1496 (N_1496,N_455,N_335);
and U1497 (N_1497,N_82,N_648);
nor U1498 (N_1498,N_462,N_205);
or U1499 (N_1499,N_658,N_21);
nor U1500 (N_1500,N_1424,N_1071);
nor U1501 (N_1501,N_763,N_1436);
or U1502 (N_1502,N_1272,N_1284);
nor U1503 (N_1503,N_1444,N_1435);
or U1504 (N_1504,N_1195,N_1470);
nor U1505 (N_1505,N_1129,N_1023);
nor U1506 (N_1506,N_976,N_1360);
xnor U1507 (N_1507,N_1497,N_1301);
or U1508 (N_1508,N_980,N_1221);
xnor U1509 (N_1509,N_1335,N_817);
nor U1510 (N_1510,N_885,N_814);
and U1511 (N_1511,N_1277,N_1306);
nor U1512 (N_1512,N_1329,N_1413);
nor U1513 (N_1513,N_1148,N_832);
nor U1514 (N_1514,N_872,N_1179);
nor U1515 (N_1515,N_1043,N_896);
and U1516 (N_1516,N_1483,N_1464);
nor U1517 (N_1517,N_788,N_1344);
nor U1518 (N_1518,N_1478,N_1034);
or U1519 (N_1519,N_1121,N_1332);
nor U1520 (N_1520,N_810,N_1499);
and U1521 (N_1521,N_1415,N_972);
nand U1522 (N_1522,N_908,N_997);
and U1523 (N_1523,N_1308,N_1025);
or U1524 (N_1524,N_1425,N_1219);
and U1525 (N_1525,N_1285,N_1136);
nand U1526 (N_1526,N_983,N_1217);
and U1527 (N_1527,N_784,N_1088);
nor U1528 (N_1528,N_1014,N_902);
nand U1529 (N_1529,N_1292,N_790);
nor U1530 (N_1530,N_1282,N_846);
or U1531 (N_1531,N_1107,N_1167);
and U1532 (N_1532,N_1317,N_1281);
nor U1533 (N_1533,N_804,N_840);
and U1534 (N_1534,N_1489,N_764);
nand U1535 (N_1535,N_1094,N_1190);
nand U1536 (N_1536,N_1248,N_1051);
nand U1537 (N_1537,N_1474,N_1168);
xor U1538 (N_1538,N_1283,N_871);
and U1539 (N_1539,N_1433,N_867);
nand U1540 (N_1540,N_919,N_1454);
or U1541 (N_1541,N_1357,N_865);
nor U1542 (N_1542,N_1491,N_1252);
or U1543 (N_1543,N_1054,N_1354);
nand U1544 (N_1544,N_1289,N_799);
or U1545 (N_1545,N_1368,N_1493);
nor U1546 (N_1546,N_786,N_775);
nand U1547 (N_1547,N_1141,N_883);
and U1548 (N_1548,N_1339,N_1003);
nor U1549 (N_1549,N_1211,N_1397);
xor U1550 (N_1550,N_1235,N_1274);
nor U1551 (N_1551,N_754,N_880);
nand U1552 (N_1552,N_955,N_889);
nand U1553 (N_1553,N_820,N_986);
nor U1554 (N_1554,N_922,N_1434);
and U1555 (N_1555,N_1017,N_1361);
nand U1556 (N_1556,N_778,N_1259);
nand U1557 (N_1557,N_1461,N_1314);
xor U1558 (N_1558,N_1198,N_1165);
nor U1559 (N_1559,N_1325,N_1253);
and U1560 (N_1560,N_1183,N_1075);
and U1561 (N_1561,N_989,N_1208);
and U1562 (N_1562,N_1061,N_848);
nor U1563 (N_1563,N_1185,N_916);
and U1564 (N_1564,N_1197,N_1116);
nand U1565 (N_1565,N_1093,N_1098);
or U1566 (N_1566,N_1322,N_1099);
nor U1567 (N_1567,N_774,N_1237);
nor U1568 (N_1568,N_1180,N_1084);
nand U1569 (N_1569,N_1092,N_1452);
or U1570 (N_1570,N_1374,N_1375);
or U1571 (N_1571,N_793,N_1134);
or U1572 (N_1572,N_1367,N_1053);
xnor U1573 (N_1573,N_1080,N_1076);
nand U1574 (N_1574,N_1495,N_1022);
nor U1575 (N_1575,N_1350,N_1460);
nand U1576 (N_1576,N_1112,N_1050);
nor U1577 (N_1577,N_1169,N_1422);
or U1578 (N_1578,N_1102,N_1471);
or U1579 (N_1579,N_1404,N_1070);
or U1580 (N_1580,N_1432,N_985);
nor U1581 (N_1581,N_1336,N_932);
nand U1582 (N_1582,N_994,N_981);
and U1583 (N_1583,N_1352,N_1192);
or U1584 (N_1584,N_1261,N_1320);
nand U1585 (N_1585,N_1286,N_993);
and U1586 (N_1586,N_1276,N_1095);
nand U1587 (N_1587,N_1273,N_1456);
nand U1588 (N_1588,N_868,N_789);
nand U1589 (N_1589,N_999,N_1420);
nand U1590 (N_1590,N_1480,N_767);
and U1591 (N_1591,N_966,N_1473);
nand U1592 (N_1592,N_958,N_1459);
or U1593 (N_1593,N_911,N_1482);
or U1594 (N_1594,N_940,N_937);
or U1595 (N_1595,N_1378,N_1152);
and U1596 (N_1596,N_1340,N_1194);
or U1597 (N_1597,N_806,N_783);
and U1598 (N_1598,N_855,N_801);
and U1599 (N_1599,N_1326,N_849);
nand U1600 (N_1600,N_1222,N_1319);
and U1601 (N_1601,N_1105,N_1278);
nor U1602 (N_1602,N_1427,N_1223);
nand U1603 (N_1603,N_1019,N_978);
nor U1604 (N_1604,N_828,N_1139);
nand U1605 (N_1605,N_821,N_1310);
and U1606 (N_1606,N_839,N_1036);
and U1607 (N_1607,N_1389,N_1002);
xnor U1608 (N_1608,N_960,N_1213);
nand U1609 (N_1609,N_1287,N_1077);
nor U1610 (N_1610,N_1363,N_1114);
or U1611 (N_1611,N_1202,N_1059);
nand U1612 (N_1612,N_1073,N_751);
or U1613 (N_1613,N_1067,N_1348);
or U1614 (N_1614,N_1486,N_965);
or U1615 (N_1615,N_948,N_1215);
nor U1616 (N_1616,N_1108,N_1451);
or U1617 (N_1617,N_1477,N_956);
nand U1618 (N_1618,N_1089,N_929);
and U1619 (N_1619,N_935,N_1242);
nand U1620 (N_1620,N_770,N_771);
and U1621 (N_1621,N_1041,N_1234);
and U1622 (N_1622,N_1462,N_949);
and U1623 (N_1623,N_1401,N_765);
xnor U1624 (N_1624,N_823,N_915);
xor U1625 (N_1625,N_984,N_1353);
or U1626 (N_1626,N_961,N_815);
and U1627 (N_1627,N_1411,N_1388);
or U1628 (N_1628,N_1083,N_1279);
nand U1629 (N_1629,N_1392,N_1062);
nor U1630 (N_1630,N_1164,N_1149);
nor U1631 (N_1631,N_1467,N_892);
nor U1632 (N_1632,N_1000,N_826);
nand U1633 (N_1633,N_1431,N_762);
nor U1634 (N_1634,N_1356,N_974);
and U1635 (N_1635,N_1450,N_878);
nand U1636 (N_1636,N_897,N_835);
nand U1637 (N_1637,N_1305,N_1160);
nand U1638 (N_1638,N_1366,N_1207);
nor U1639 (N_1639,N_1052,N_782);
nand U1640 (N_1640,N_1391,N_1333);
and U1641 (N_1641,N_1334,N_1072);
nand U1642 (N_1642,N_1396,N_1465);
nand U1643 (N_1643,N_1300,N_1498);
nand U1644 (N_1644,N_943,N_1091);
or U1645 (N_1645,N_863,N_1119);
or U1646 (N_1646,N_1153,N_1056);
nand U1647 (N_1647,N_1040,N_1162);
or U1648 (N_1648,N_795,N_876);
xor U1649 (N_1649,N_1176,N_777);
and U1650 (N_1650,N_1120,N_825);
or U1651 (N_1651,N_1086,N_931);
and U1652 (N_1652,N_1142,N_1426);
or U1653 (N_1653,N_1358,N_1209);
nand U1654 (N_1654,N_1214,N_964);
nand U1655 (N_1655,N_1122,N_1047);
and U1656 (N_1656,N_973,N_923);
nor U1657 (N_1657,N_1011,N_874);
and U1658 (N_1658,N_1137,N_1200);
and U1659 (N_1659,N_951,N_1245);
and U1660 (N_1660,N_977,N_870);
nor U1661 (N_1661,N_776,N_1100);
or U1662 (N_1662,N_1395,N_1417);
nor U1663 (N_1663,N_1312,N_1031);
nand U1664 (N_1664,N_1270,N_1146);
nand U1665 (N_1665,N_1403,N_845);
nand U1666 (N_1666,N_904,N_903);
nor U1667 (N_1667,N_895,N_811);
or U1668 (N_1668,N_1382,N_1265);
nand U1669 (N_1669,N_1324,N_1488);
and U1670 (N_1670,N_1455,N_1231);
and U1671 (N_1671,N_1342,N_809);
and U1672 (N_1672,N_1238,N_1163);
and U1673 (N_1673,N_1406,N_750);
nor U1674 (N_1674,N_1257,N_818);
nand U1675 (N_1675,N_785,N_780);
or U1676 (N_1676,N_1005,N_796);
nor U1677 (N_1677,N_1085,N_1386);
or U1678 (N_1678,N_1132,N_1264);
xnor U1679 (N_1679,N_873,N_1127);
and U1680 (N_1680,N_1027,N_830);
nor U1681 (N_1681,N_859,N_1079);
nand U1682 (N_1682,N_1065,N_901);
nor U1683 (N_1683,N_969,N_1158);
and U1684 (N_1684,N_864,N_1299);
or U1685 (N_1685,N_1345,N_1372);
or U1686 (N_1686,N_1428,N_1421);
and U1687 (N_1687,N_1321,N_1104);
xor U1688 (N_1688,N_1206,N_794);
nand U1689 (N_1689,N_831,N_1430);
and U1690 (N_1690,N_1410,N_1055);
or U1691 (N_1691,N_1263,N_1103);
nor U1692 (N_1692,N_1390,N_1385);
nand U1693 (N_1693,N_1013,N_1416);
and U1694 (N_1694,N_1295,N_1068);
or U1695 (N_1695,N_1302,N_875);
or U1696 (N_1696,N_1203,N_1090);
xnor U1697 (N_1697,N_879,N_1399);
nor U1698 (N_1698,N_850,N_800);
nor U1699 (N_1699,N_933,N_1443);
nor U1700 (N_1700,N_851,N_1446);
nor U1701 (N_1701,N_1131,N_1117);
and U1702 (N_1702,N_996,N_987);
nor U1703 (N_1703,N_914,N_833);
or U1704 (N_1704,N_808,N_913);
nor U1705 (N_1705,N_1193,N_1161);
or U1706 (N_1706,N_759,N_829);
nand U1707 (N_1707,N_1442,N_1479);
nor U1708 (N_1708,N_772,N_1266);
nor U1709 (N_1709,N_1196,N_1255);
or U1710 (N_1710,N_939,N_1042);
or U1711 (N_1711,N_1126,N_1384);
nor U1712 (N_1712,N_1125,N_858);
or U1713 (N_1713,N_899,N_942);
xor U1714 (N_1714,N_1124,N_1189);
nand U1715 (N_1715,N_1240,N_861);
nor U1716 (N_1716,N_930,N_1037);
nor U1717 (N_1717,N_952,N_1174);
nand U1718 (N_1718,N_1408,N_1156);
nor U1719 (N_1719,N_1081,N_834);
and U1720 (N_1720,N_1045,N_886);
nor U1721 (N_1721,N_1177,N_1186);
and U1722 (N_1722,N_1220,N_1371);
nand U1723 (N_1723,N_1307,N_970);
nand U1724 (N_1724,N_1101,N_910);
nor U1725 (N_1725,N_947,N_975);
nand U1726 (N_1726,N_852,N_1331);
nor U1727 (N_1727,N_946,N_1018);
or U1728 (N_1728,N_1337,N_926);
or U1729 (N_1729,N_1316,N_816);
nor U1730 (N_1730,N_1251,N_1106);
or U1731 (N_1731,N_1347,N_1380);
nor U1732 (N_1732,N_928,N_807);
nor U1733 (N_1733,N_798,N_779);
or U1734 (N_1734,N_805,N_971);
and U1735 (N_1735,N_802,N_1269);
nand U1736 (N_1736,N_792,N_841);
nor U1737 (N_1737,N_1074,N_1243);
nor U1738 (N_1738,N_894,N_1173);
and U1739 (N_1739,N_1323,N_1438);
nand U1740 (N_1740,N_1078,N_891);
or U1741 (N_1741,N_1063,N_1006);
nor U1742 (N_1742,N_917,N_927);
or U1743 (N_1743,N_1010,N_824);
and U1744 (N_1744,N_1191,N_945);
and U1745 (N_1745,N_1387,N_954);
nor U1746 (N_1746,N_1365,N_1212);
nor U1747 (N_1747,N_1230,N_1030);
nand U1748 (N_1748,N_1058,N_1032);
nor U1749 (N_1749,N_1138,N_1143);
nor U1750 (N_1750,N_853,N_1039);
and U1751 (N_1751,N_1327,N_1400);
nor U1752 (N_1752,N_925,N_1412);
or U1753 (N_1753,N_838,N_1241);
or U1754 (N_1754,N_1256,N_1311);
nand U1755 (N_1755,N_1267,N_1304);
nand U1756 (N_1756,N_1172,N_998);
or U1757 (N_1757,N_1181,N_1066);
nand U1758 (N_1758,N_1049,N_1439);
and U1759 (N_1759,N_950,N_843);
or U1760 (N_1760,N_1318,N_819);
and U1761 (N_1761,N_1377,N_1381);
nand U1762 (N_1762,N_1469,N_761);
nor U1763 (N_1763,N_1024,N_890);
or U1764 (N_1764,N_769,N_1171);
and U1765 (N_1765,N_968,N_860);
nor U1766 (N_1766,N_766,N_979);
or U1767 (N_1767,N_869,N_1414);
and U1768 (N_1768,N_1182,N_1496);
nand U1769 (N_1769,N_1205,N_1349);
and U1770 (N_1770,N_1250,N_1188);
nor U1771 (N_1771,N_758,N_1447);
nand U1772 (N_1772,N_1407,N_1458);
or U1773 (N_1773,N_995,N_1001);
nor U1774 (N_1774,N_1216,N_1315);
nor U1775 (N_1775,N_1096,N_1262);
nor U1776 (N_1776,N_1402,N_1369);
and U1777 (N_1777,N_755,N_1440);
nand U1778 (N_1778,N_1233,N_1110);
or U1779 (N_1779,N_1244,N_857);
nand U1780 (N_1780,N_1437,N_877);
nand U1781 (N_1781,N_847,N_1419);
and U1782 (N_1782,N_1151,N_1466);
nand U1783 (N_1783,N_1028,N_812);
nand U1784 (N_1784,N_1429,N_1135);
nand U1785 (N_1785,N_1298,N_837);
and U1786 (N_1786,N_938,N_1441);
or U1787 (N_1787,N_1330,N_1475);
nand U1788 (N_1788,N_1309,N_1409);
or U1789 (N_1789,N_753,N_1405);
nand U1790 (N_1790,N_1113,N_1170);
nand U1791 (N_1791,N_1355,N_1423);
or U1792 (N_1792,N_1115,N_881);
nor U1793 (N_1793,N_898,N_1015);
or U1794 (N_1794,N_990,N_1166);
nor U1795 (N_1795,N_1383,N_1463);
and U1796 (N_1796,N_957,N_1145);
nand U1797 (N_1797,N_1449,N_921);
nand U1798 (N_1798,N_1118,N_1044);
and U1799 (N_1799,N_1007,N_1128);
xor U1800 (N_1800,N_813,N_941);
and U1801 (N_1801,N_1236,N_1109);
nand U1802 (N_1802,N_1020,N_752);
nor U1803 (N_1803,N_1009,N_1258);
and U1804 (N_1804,N_1150,N_866);
or U1805 (N_1805,N_822,N_773);
or U1806 (N_1806,N_1069,N_1379);
and U1807 (N_1807,N_797,N_1359);
nor U1808 (N_1808,N_1485,N_1341);
or U1809 (N_1809,N_1472,N_1038);
nand U1810 (N_1810,N_988,N_1154);
nand U1811 (N_1811,N_1199,N_1016);
and U1812 (N_1812,N_1376,N_887);
nor U1813 (N_1813,N_856,N_827);
nand U1814 (N_1814,N_1296,N_1362);
and U1815 (N_1815,N_909,N_1140);
and U1816 (N_1816,N_963,N_1490);
and U1817 (N_1817,N_1260,N_1228);
or U1818 (N_1818,N_1057,N_1147);
nand U1819 (N_1819,N_1224,N_1492);
or U1820 (N_1820,N_842,N_1291);
nor U1821 (N_1821,N_1445,N_1249);
nand U1822 (N_1822,N_836,N_1394);
and U1823 (N_1823,N_1346,N_982);
xnor U1824 (N_1824,N_1364,N_991);
xor U1825 (N_1825,N_1029,N_1159);
nor U1826 (N_1826,N_1229,N_1476);
or U1827 (N_1827,N_1210,N_962);
nand U1828 (N_1828,N_1481,N_1004);
and U1829 (N_1829,N_1133,N_1453);
nand U1830 (N_1830,N_1082,N_1268);
and U1831 (N_1831,N_920,N_1111);
nand U1832 (N_1832,N_944,N_757);
and U1833 (N_1833,N_959,N_862);
or U1834 (N_1834,N_1290,N_1087);
or U1835 (N_1835,N_1157,N_1232);
or U1836 (N_1836,N_1060,N_1123);
or U1837 (N_1837,N_1184,N_1370);
nand U1838 (N_1838,N_1226,N_1175);
nand U1839 (N_1839,N_1254,N_1008);
and U1840 (N_1840,N_912,N_1201);
nand U1841 (N_1841,N_1144,N_1033);
nor U1842 (N_1842,N_900,N_1393);
nor U1843 (N_1843,N_1048,N_844);
or U1844 (N_1844,N_882,N_768);
nand U1845 (N_1845,N_893,N_905);
nor U1846 (N_1846,N_1021,N_1293);
nor U1847 (N_1847,N_1294,N_1187);
or U1848 (N_1848,N_1398,N_787);
xnor U1849 (N_1849,N_1012,N_1343);
or U1850 (N_1850,N_1484,N_1064);
and U1851 (N_1851,N_1468,N_1097);
nor U1852 (N_1852,N_1275,N_967);
nand U1853 (N_1853,N_992,N_1246);
and U1854 (N_1854,N_1313,N_907);
nor U1855 (N_1855,N_760,N_791);
nand U1856 (N_1856,N_1448,N_918);
or U1857 (N_1857,N_924,N_1225);
or U1858 (N_1858,N_934,N_1338);
nand U1859 (N_1859,N_953,N_1204);
nand U1860 (N_1860,N_1247,N_936);
nor U1861 (N_1861,N_803,N_1046);
or U1862 (N_1862,N_888,N_1487);
xor U1863 (N_1863,N_906,N_1418);
or U1864 (N_1864,N_1218,N_1288);
or U1865 (N_1865,N_1239,N_1457);
or U1866 (N_1866,N_781,N_854);
and U1867 (N_1867,N_1271,N_1026);
nor U1868 (N_1868,N_1303,N_1035);
nand U1869 (N_1869,N_1227,N_1328);
nor U1870 (N_1870,N_1494,N_884);
and U1871 (N_1871,N_1280,N_1373);
nor U1872 (N_1872,N_756,N_1297);
or U1873 (N_1873,N_1130,N_1178);
and U1874 (N_1874,N_1351,N_1155);
nor U1875 (N_1875,N_1026,N_987);
and U1876 (N_1876,N_1114,N_838);
nor U1877 (N_1877,N_1024,N_1319);
nand U1878 (N_1878,N_1206,N_1327);
nor U1879 (N_1879,N_1165,N_1235);
and U1880 (N_1880,N_1042,N_1183);
nor U1881 (N_1881,N_1408,N_916);
and U1882 (N_1882,N_1215,N_1140);
and U1883 (N_1883,N_1478,N_800);
nor U1884 (N_1884,N_985,N_1141);
and U1885 (N_1885,N_1469,N_1166);
xnor U1886 (N_1886,N_1032,N_859);
or U1887 (N_1887,N_1202,N_1418);
or U1888 (N_1888,N_1156,N_793);
or U1889 (N_1889,N_1203,N_772);
nor U1890 (N_1890,N_1460,N_1472);
and U1891 (N_1891,N_1476,N_1454);
nand U1892 (N_1892,N_1261,N_979);
and U1893 (N_1893,N_907,N_1183);
nand U1894 (N_1894,N_1254,N_1098);
nand U1895 (N_1895,N_944,N_793);
and U1896 (N_1896,N_1092,N_1210);
and U1897 (N_1897,N_1044,N_1310);
nor U1898 (N_1898,N_1016,N_1394);
or U1899 (N_1899,N_1123,N_1070);
nor U1900 (N_1900,N_1416,N_1405);
nand U1901 (N_1901,N_775,N_767);
nand U1902 (N_1902,N_924,N_1112);
nand U1903 (N_1903,N_887,N_1455);
or U1904 (N_1904,N_1189,N_1198);
or U1905 (N_1905,N_1108,N_954);
and U1906 (N_1906,N_1105,N_1082);
and U1907 (N_1907,N_932,N_1090);
nor U1908 (N_1908,N_1289,N_893);
and U1909 (N_1909,N_789,N_1496);
nor U1910 (N_1910,N_1032,N_1239);
or U1911 (N_1911,N_1126,N_1124);
or U1912 (N_1912,N_1057,N_1431);
xnor U1913 (N_1913,N_1091,N_823);
or U1914 (N_1914,N_844,N_880);
nand U1915 (N_1915,N_1432,N_1415);
nor U1916 (N_1916,N_924,N_1418);
or U1917 (N_1917,N_1323,N_1444);
and U1918 (N_1918,N_1292,N_912);
nor U1919 (N_1919,N_1445,N_1300);
nand U1920 (N_1920,N_996,N_1441);
and U1921 (N_1921,N_966,N_1392);
nor U1922 (N_1922,N_1323,N_986);
nand U1923 (N_1923,N_1000,N_1179);
or U1924 (N_1924,N_953,N_772);
and U1925 (N_1925,N_1070,N_1243);
nand U1926 (N_1926,N_1123,N_1131);
xnor U1927 (N_1927,N_1248,N_782);
or U1928 (N_1928,N_1196,N_930);
nand U1929 (N_1929,N_1397,N_984);
nand U1930 (N_1930,N_1431,N_1143);
nand U1931 (N_1931,N_1052,N_1429);
or U1932 (N_1932,N_1337,N_1316);
nor U1933 (N_1933,N_963,N_1316);
nor U1934 (N_1934,N_1009,N_1381);
nand U1935 (N_1935,N_978,N_1052);
nand U1936 (N_1936,N_1196,N_879);
nand U1937 (N_1937,N_1224,N_758);
nor U1938 (N_1938,N_1436,N_1472);
or U1939 (N_1939,N_879,N_788);
or U1940 (N_1940,N_1349,N_833);
and U1941 (N_1941,N_1497,N_910);
and U1942 (N_1942,N_1244,N_903);
nand U1943 (N_1943,N_1317,N_1482);
nand U1944 (N_1944,N_1431,N_903);
or U1945 (N_1945,N_1464,N_1330);
or U1946 (N_1946,N_1006,N_837);
nor U1947 (N_1947,N_1113,N_762);
or U1948 (N_1948,N_1269,N_1048);
nor U1949 (N_1949,N_1015,N_834);
nand U1950 (N_1950,N_1320,N_1463);
nor U1951 (N_1951,N_1084,N_1220);
and U1952 (N_1952,N_1347,N_1015);
nand U1953 (N_1953,N_887,N_1084);
or U1954 (N_1954,N_846,N_1247);
and U1955 (N_1955,N_807,N_1410);
nand U1956 (N_1956,N_1386,N_1465);
and U1957 (N_1957,N_1210,N_1114);
or U1958 (N_1958,N_1025,N_832);
nand U1959 (N_1959,N_1281,N_1102);
nand U1960 (N_1960,N_1264,N_1010);
nor U1961 (N_1961,N_791,N_1351);
nor U1962 (N_1962,N_964,N_1377);
xor U1963 (N_1963,N_896,N_1296);
nand U1964 (N_1964,N_990,N_1257);
and U1965 (N_1965,N_1045,N_1189);
or U1966 (N_1966,N_1212,N_1353);
or U1967 (N_1967,N_1361,N_1395);
and U1968 (N_1968,N_1416,N_1110);
and U1969 (N_1969,N_1384,N_941);
nor U1970 (N_1970,N_931,N_1055);
and U1971 (N_1971,N_1306,N_1029);
nand U1972 (N_1972,N_1121,N_1310);
and U1973 (N_1973,N_1111,N_1082);
and U1974 (N_1974,N_1008,N_1164);
or U1975 (N_1975,N_1483,N_1493);
nor U1976 (N_1976,N_1005,N_991);
nor U1977 (N_1977,N_1299,N_1420);
or U1978 (N_1978,N_1372,N_1152);
or U1979 (N_1979,N_993,N_982);
or U1980 (N_1980,N_1391,N_893);
nand U1981 (N_1981,N_1259,N_898);
and U1982 (N_1982,N_1253,N_1461);
or U1983 (N_1983,N_1262,N_785);
and U1984 (N_1984,N_908,N_1262);
nor U1985 (N_1985,N_849,N_1262);
and U1986 (N_1986,N_881,N_1146);
nor U1987 (N_1987,N_1286,N_1284);
and U1988 (N_1988,N_1097,N_1241);
and U1989 (N_1989,N_754,N_1177);
or U1990 (N_1990,N_816,N_1433);
and U1991 (N_1991,N_1169,N_1397);
nor U1992 (N_1992,N_1448,N_997);
or U1993 (N_1993,N_1113,N_1181);
nor U1994 (N_1994,N_904,N_993);
nor U1995 (N_1995,N_1044,N_1438);
or U1996 (N_1996,N_1450,N_1464);
and U1997 (N_1997,N_1346,N_1499);
or U1998 (N_1998,N_1143,N_1073);
nand U1999 (N_1999,N_1069,N_917);
nor U2000 (N_2000,N_931,N_972);
nand U2001 (N_2001,N_1495,N_819);
or U2002 (N_2002,N_927,N_1176);
or U2003 (N_2003,N_1420,N_959);
nand U2004 (N_2004,N_1115,N_1404);
nor U2005 (N_2005,N_1126,N_1490);
or U2006 (N_2006,N_1231,N_1473);
and U2007 (N_2007,N_844,N_1039);
nand U2008 (N_2008,N_1047,N_991);
nor U2009 (N_2009,N_1338,N_824);
and U2010 (N_2010,N_1161,N_979);
nor U2011 (N_2011,N_1015,N_986);
or U2012 (N_2012,N_969,N_765);
nor U2013 (N_2013,N_1117,N_1491);
and U2014 (N_2014,N_1495,N_1174);
nor U2015 (N_2015,N_957,N_1377);
and U2016 (N_2016,N_849,N_799);
and U2017 (N_2017,N_1451,N_1109);
nor U2018 (N_2018,N_1041,N_1313);
nand U2019 (N_2019,N_888,N_1334);
and U2020 (N_2020,N_1262,N_1076);
and U2021 (N_2021,N_967,N_1050);
and U2022 (N_2022,N_1338,N_1125);
nor U2023 (N_2023,N_863,N_1002);
nor U2024 (N_2024,N_792,N_966);
nor U2025 (N_2025,N_1028,N_1051);
nand U2026 (N_2026,N_1309,N_808);
nor U2027 (N_2027,N_1414,N_1200);
nand U2028 (N_2028,N_761,N_1043);
or U2029 (N_2029,N_1393,N_779);
nor U2030 (N_2030,N_906,N_1187);
and U2031 (N_2031,N_1092,N_1057);
nor U2032 (N_2032,N_1272,N_1065);
nand U2033 (N_2033,N_761,N_948);
nor U2034 (N_2034,N_1458,N_969);
and U2035 (N_2035,N_753,N_1186);
nand U2036 (N_2036,N_1008,N_1090);
nor U2037 (N_2037,N_1422,N_869);
or U2038 (N_2038,N_1165,N_796);
and U2039 (N_2039,N_1341,N_1370);
and U2040 (N_2040,N_1011,N_1140);
and U2041 (N_2041,N_976,N_1404);
and U2042 (N_2042,N_1011,N_1055);
and U2043 (N_2043,N_1260,N_1240);
or U2044 (N_2044,N_887,N_988);
or U2045 (N_2045,N_839,N_963);
nand U2046 (N_2046,N_777,N_780);
nand U2047 (N_2047,N_1335,N_1138);
or U2048 (N_2048,N_964,N_806);
nand U2049 (N_2049,N_923,N_816);
and U2050 (N_2050,N_1365,N_1039);
nand U2051 (N_2051,N_803,N_1000);
nand U2052 (N_2052,N_953,N_1486);
or U2053 (N_2053,N_897,N_1191);
nor U2054 (N_2054,N_1133,N_1441);
and U2055 (N_2055,N_918,N_1330);
nand U2056 (N_2056,N_1062,N_1178);
nand U2057 (N_2057,N_1098,N_1283);
or U2058 (N_2058,N_1388,N_755);
and U2059 (N_2059,N_1008,N_1392);
or U2060 (N_2060,N_1489,N_1017);
or U2061 (N_2061,N_1247,N_1185);
nor U2062 (N_2062,N_1350,N_1453);
nand U2063 (N_2063,N_1079,N_1473);
and U2064 (N_2064,N_999,N_1162);
xnor U2065 (N_2065,N_820,N_1320);
nand U2066 (N_2066,N_934,N_761);
nor U2067 (N_2067,N_863,N_1420);
nor U2068 (N_2068,N_1118,N_783);
nor U2069 (N_2069,N_1401,N_1015);
and U2070 (N_2070,N_1386,N_818);
nor U2071 (N_2071,N_1051,N_1429);
nand U2072 (N_2072,N_1230,N_1305);
or U2073 (N_2073,N_886,N_1375);
or U2074 (N_2074,N_1218,N_1463);
nor U2075 (N_2075,N_1255,N_1148);
xor U2076 (N_2076,N_1175,N_1064);
nor U2077 (N_2077,N_922,N_1254);
xor U2078 (N_2078,N_1013,N_1362);
nand U2079 (N_2079,N_1028,N_1031);
and U2080 (N_2080,N_1099,N_1141);
nor U2081 (N_2081,N_1014,N_1482);
or U2082 (N_2082,N_967,N_946);
and U2083 (N_2083,N_1338,N_847);
nor U2084 (N_2084,N_907,N_780);
or U2085 (N_2085,N_1284,N_1028);
and U2086 (N_2086,N_923,N_1160);
nand U2087 (N_2087,N_1208,N_1230);
and U2088 (N_2088,N_861,N_786);
nor U2089 (N_2089,N_1036,N_1333);
nand U2090 (N_2090,N_1401,N_1166);
nor U2091 (N_2091,N_1481,N_1270);
and U2092 (N_2092,N_836,N_1344);
nand U2093 (N_2093,N_1275,N_1484);
and U2094 (N_2094,N_1169,N_1461);
or U2095 (N_2095,N_1006,N_1286);
or U2096 (N_2096,N_985,N_839);
or U2097 (N_2097,N_1097,N_934);
and U2098 (N_2098,N_916,N_1110);
nand U2099 (N_2099,N_852,N_1220);
and U2100 (N_2100,N_1378,N_1174);
or U2101 (N_2101,N_1060,N_1498);
nand U2102 (N_2102,N_963,N_1283);
nand U2103 (N_2103,N_1196,N_1279);
and U2104 (N_2104,N_791,N_1404);
or U2105 (N_2105,N_1401,N_1053);
nand U2106 (N_2106,N_1490,N_871);
nand U2107 (N_2107,N_1139,N_779);
nor U2108 (N_2108,N_1004,N_1436);
and U2109 (N_2109,N_1138,N_836);
nand U2110 (N_2110,N_1420,N_1426);
nor U2111 (N_2111,N_1244,N_1290);
or U2112 (N_2112,N_1213,N_843);
nand U2113 (N_2113,N_1251,N_931);
and U2114 (N_2114,N_867,N_925);
and U2115 (N_2115,N_1122,N_985);
nor U2116 (N_2116,N_978,N_839);
nor U2117 (N_2117,N_1177,N_1381);
nor U2118 (N_2118,N_1285,N_1230);
nor U2119 (N_2119,N_952,N_917);
nand U2120 (N_2120,N_924,N_1065);
or U2121 (N_2121,N_1455,N_1016);
and U2122 (N_2122,N_891,N_1155);
nor U2123 (N_2123,N_1265,N_1155);
nor U2124 (N_2124,N_1148,N_1441);
or U2125 (N_2125,N_1381,N_1156);
or U2126 (N_2126,N_1251,N_879);
nor U2127 (N_2127,N_1028,N_1367);
nor U2128 (N_2128,N_1104,N_1324);
and U2129 (N_2129,N_1215,N_1411);
and U2130 (N_2130,N_911,N_1198);
nor U2131 (N_2131,N_1499,N_1008);
or U2132 (N_2132,N_1062,N_1367);
and U2133 (N_2133,N_1080,N_1138);
xnor U2134 (N_2134,N_877,N_1302);
or U2135 (N_2135,N_1135,N_1080);
or U2136 (N_2136,N_864,N_982);
xnor U2137 (N_2137,N_1193,N_1110);
and U2138 (N_2138,N_837,N_1497);
nand U2139 (N_2139,N_1379,N_1073);
nand U2140 (N_2140,N_1062,N_1263);
and U2141 (N_2141,N_1149,N_986);
and U2142 (N_2142,N_1239,N_1373);
and U2143 (N_2143,N_1370,N_1483);
nand U2144 (N_2144,N_1128,N_1416);
nand U2145 (N_2145,N_1492,N_1148);
or U2146 (N_2146,N_1153,N_1255);
and U2147 (N_2147,N_852,N_1487);
nor U2148 (N_2148,N_1095,N_1310);
xor U2149 (N_2149,N_1117,N_1450);
nor U2150 (N_2150,N_1207,N_1225);
or U2151 (N_2151,N_1113,N_862);
nor U2152 (N_2152,N_820,N_1339);
nor U2153 (N_2153,N_1305,N_992);
nor U2154 (N_2154,N_1354,N_770);
or U2155 (N_2155,N_808,N_1160);
nor U2156 (N_2156,N_1149,N_1334);
or U2157 (N_2157,N_1464,N_1443);
nor U2158 (N_2158,N_796,N_1014);
or U2159 (N_2159,N_974,N_1376);
or U2160 (N_2160,N_800,N_1299);
nor U2161 (N_2161,N_795,N_1497);
or U2162 (N_2162,N_968,N_1255);
and U2163 (N_2163,N_1457,N_920);
xnor U2164 (N_2164,N_977,N_1054);
nor U2165 (N_2165,N_1259,N_1408);
nor U2166 (N_2166,N_1207,N_1030);
nor U2167 (N_2167,N_753,N_1453);
nand U2168 (N_2168,N_1462,N_1130);
xor U2169 (N_2169,N_1039,N_1471);
and U2170 (N_2170,N_796,N_1364);
and U2171 (N_2171,N_1380,N_1104);
and U2172 (N_2172,N_1311,N_1263);
nor U2173 (N_2173,N_949,N_1094);
or U2174 (N_2174,N_772,N_1083);
nand U2175 (N_2175,N_845,N_1036);
nand U2176 (N_2176,N_1497,N_758);
nor U2177 (N_2177,N_769,N_1395);
or U2178 (N_2178,N_1273,N_928);
or U2179 (N_2179,N_876,N_1213);
nand U2180 (N_2180,N_1278,N_1139);
or U2181 (N_2181,N_1450,N_1085);
and U2182 (N_2182,N_852,N_1226);
nand U2183 (N_2183,N_1118,N_1314);
nor U2184 (N_2184,N_1179,N_797);
nand U2185 (N_2185,N_863,N_1203);
nor U2186 (N_2186,N_806,N_1266);
nand U2187 (N_2187,N_776,N_1298);
nor U2188 (N_2188,N_1223,N_1305);
xor U2189 (N_2189,N_1486,N_1040);
xor U2190 (N_2190,N_1136,N_1317);
and U2191 (N_2191,N_1368,N_1392);
and U2192 (N_2192,N_1430,N_1315);
nor U2193 (N_2193,N_1433,N_1409);
and U2194 (N_2194,N_1499,N_870);
nor U2195 (N_2195,N_1064,N_1018);
and U2196 (N_2196,N_752,N_849);
nand U2197 (N_2197,N_778,N_864);
nand U2198 (N_2198,N_1001,N_1210);
nor U2199 (N_2199,N_892,N_763);
and U2200 (N_2200,N_1321,N_1124);
nand U2201 (N_2201,N_1123,N_1419);
and U2202 (N_2202,N_1012,N_961);
and U2203 (N_2203,N_917,N_1427);
and U2204 (N_2204,N_1368,N_799);
nor U2205 (N_2205,N_1407,N_1369);
nor U2206 (N_2206,N_953,N_786);
and U2207 (N_2207,N_1037,N_935);
xor U2208 (N_2208,N_1072,N_1376);
nand U2209 (N_2209,N_852,N_903);
nand U2210 (N_2210,N_978,N_1089);
and U2211 (N_2211,N_1340,N_1011);
nor U2212 (N_2212,N_1158,N_751);
nand U2213 (N_2213,N_1103,N_838);
or U2214 (N_2214,N_1289,N_1372);
and U2215 (N_2215,N_969,N_1180);
or U2216 (N_2216,N_1362,N_1361);
or U2217 (N_2217,N_1293,N_1201);
xnor U2218 (N_2218,N_1029,N_786);
or U2219 (N_2219,N_754,N_1339);
or U2220 (N_2220,N_917,N_1204);
and U2221 (N_2221,N_1394,N_1440);
or U2222 (N_2222,N_812,N_883);
or U2223 (N_2223,N_822,N_1195);
nand U2224 (N_2224,N_1189,N_753);
and U2225 (N_2225,N_1351,N_836);
nor U2226 (N_2226,N_1030,N_1061);
or U2227 (N_2227,N_838,N_863);
and U2228 (N_2228,N_1421,N_805);
and U2229 (N_2229,N_792,N_1341);
xor U2230 (N_2230,N_928,N_844);
nor U2231 (N_2231,N_1307,N_1490);
nor U2232 (N_2232,N_1418,N_1253);
and U2233 (N_2233,N_1056,N_1011);
nor U2234 (N_2234,N_1001,N_1354);
nor U2235 (N_2235,N_1444,N_1096);
nand U2236 (N_2236,N_785,N_1077);
nor U2237 (N_2237,N_806,N_1392);
or U2238 (N_2238,N_821,N_1485);
nor U2239 (N_2239,N_1388,N_1402);
or U2240 (N_2240,N_782,N_1009);
nand U2241 (N_2241,N_1405,N_1023);
or U2242 (N_2242,N_1125,N_897);
and U2243 (N_2243,N_753,N_1377);
nand U2244 (N_2244,N_1067,N_1041);
or U2245 (N_2245,N_1125,N_1166);
and U2246 (N_2246,N_1160,N_1141);
or U2247 (N_2247,N_807,N_1154);
and U2248 (N_2248,N_1005,N_1010);
nor U2249 (N_2249,N_930,N_1042);
nand U2250 (N_2250,N_1662,N_2043);
and U2251 (N_2251,N_2037,N_2136);
or U2252 (N_2252,N_1558,N_2101);
nor U2253 (N_2253,N_1556,N_1771);
nor U2254 (N_2254,N_2002,N_2107);
and U2255 (N_2255,N_1841,N_1557);
nor U2256 (N_2256,N_1990,N_1920);
xor U2257 (N_2257,N_1524,N_1855);
and U2258 (N_2258,N_1623,N_1895);
xnor U2259 (N_2259,N_1714,N_2204);
or U2260 (N_2260,N_2062,N_1818);
nor U2261 (N_2261,N_1819,N_1859);
or U2262 (N_2262,N_1526,N_1713);
nand U2263 (N_2263,N_1608,N_1978);
nand U2264 (N_2264,N_2019,N_1531);
and U2265 (N_2265,N_1508,N_1917);
nor U2266 (N_2266,N_2081,N_1760);
nand U2267 (N_2267,N_1629,N_2125);
and U2268 (N_2268,N_2144,N_2229);
and U2269 (N_2269,N_1780,N_1597);
and U2270 (N_2270,N_2115,N_1919);
nand U2271 (N_2271,N_1875,N_2075);
nand U2272 (N_2272,N_1987,N_1973);
xor U2273 (N_2273,N_1532,N_2242);
and U2274 (N_2274,N_2235,N_1672);
and U2275 (N_2275,N_1829,N_2152);
and U2276 (N_2276,N_1507,N_1757);
nand U2277 (N_2277,N_1610,N_2195);
or U2278 (N_2278,N_1779,N_1805);
and U2279 (N_2279,N_2181,N_1918);
and U2280 (N_2280,N_1665,N_1886);
and U2281 (N_2281,N_1640,N_1799);
nand U2282 (N_2282,N_1704,N_1935);
and U2283 (N_2283,N_2032,N_1784);
nor U2284 (N_2284,N_1904,N_1809);
nand U2285 (N_2285,N_1753,N_2096);
nand U2286 (N_2286,N_1719,N_1739);
or U2287 (N_2287,N_1942,N_2063);
or U2288 (N_2288,N_1535,N_2141);
and U2289 (N_2289,N_1851,N_1647);
or U2290 (N_2290,N_2190,N_2247);
nor U2291 (N_2291,N_1677,N_1756);
or U2292 (N_2292,N_2145,N_1827);
or U2293 (N_2293,N_1939,N_1525);
nor U2294 (N_2294,N_1845,N_1907);
or U2295 (N_2295,N_2066,N_1858);
nand U2296 (N_2296,N_2087,N_1667);
nand U2297 (N_2297,N_2153,N_1601);
nand U2298 (N_2298,N_2046,N_2243);
or U2299 (N_2299,N_1506,N_1590);
and U2300 (N_2300,N_2016,N_1925);
and U2301 (N_2301,N_1947,N_1766);
nand U2302 (N_2302,N_1765,N_1706);
or U2303 (N_2303,N_1584,N_2034);
and U2304 (N_2304,N_1964,N_1847);
nor U2305 (N_2305,N_2180,N_1700);
or U2306 (N_2306,N_1835,N_1888);
nor U2307 (N_2307,N_1781,N_1878);
or U2308 (N_2308,N_2234,N_2070);
and U2309 (N_2309,N_1802,N_2124);
nor U2310 (N_2310,N_1931,N_2134);
nand U2311 (N_2311,N_2139,N_1619);
and U2312 (N_2312,N_2201,N_1566);
nor U2313 (N_2313,N_1537,N_2004);
nor U2314 (N_2314,N_1993,N_1767);
nor U2315 (N_2315,N_2020,N_1561);
and U2316 (N_2316,N_1581,N_2199);
nand U2317 (N_2317,N_2148,N_1966);
or U2318 (N_2318,N_1645,N_2011);
and U2319 (N_2319,N_1592,N_2060);
nor U2320 (N_2320,N_1881,N_1540);
and U2321 (N_2321,N_1746,N_2095);
or U2322 (N_2322,N_1902,N_1957);
xnor U2323 (N_2323,N_1913,N_1909);
nand U2324 (N_2324,N_1926,N_1960);
nor U2325 (N_2325,N_1999,N_1527);
or U2326 (N_2326,N_1981,N_1500);
and U2327 (N_2327,N_1988,N_2006);
or U2328 (N_2328,N_2179,N_1798);
nand U2329 (N_2329,N_1808,N_2098);
nor U2330 (N_2330,N_1650,N_2228);
nand U2331 (N_2331,N_1789,N_1518);
nand U2332 (N_2332,N_1785,N_1600);
or U2333 (N_2333,N_2140,N_1980);
nand U2334 (N_2334,N_1728,N_1974);
nor U2335 (N_2335,N_1937,N_1727);
or U2336 (N_2336,N_2039,N_1661);
and U2337 (N_2337,N_2240,N_2208);
nor U2338 (N_2338,N_1996,N_1961);
and U2339 (N_2339,N_1837,N_1560);
or U2340 (N_2340,N_2220,N_1534);
nor U2341 (N_2341,N_1596,N_1825);
nor U2342 (N_2342,N_2003,N_1945);
or U2343 (N_2343,N_2033,N_1657);
and U2344 (N_2344,N_1738,N_1754);
nand U2345 (N_2345,N_1834,N_2073);
nand U2346 (N_2346,N_1733,N_1620);
and U2347 (N_2347,N_1857,N_1876);
nor U2348 (N_2348,N_2216,N_1711);
and U2349 (N_2349,N_2093,N_1747);
and U2350 (N_2350,N_1529,N_2050);
nor U2351 (N_2351,N_1972,N_1811);
or U2352 (N_2352,N_1501,N_1885);
nor U2353 (N_2353,N_1502,N_2238);
nand U2354 (N_2354,N_1963,N_2080);
nor U2355 (N_2355,N_1703,N_1846);
nand U2356 (N_2356,N_1853,N_1962);
or U2357 (N_2357,N_1887,N_1669);
nor U2358 (N_2358,N_1938,N_1850);
nand U2359 (N_2359,N_2131,N_2097);
nor U2360 (N_2360,N_2083,N_2085);
nor U2361 (N_2361,N_1598,N_1530);
nor U2362 (N_2362,N_2036,N_1605);
nor U2363 (N_2363,N_1674,N_1539);
or U2364 (N_2364,N_2117,N_2106);
and U2365 (N_2365,N_1796,N_1624);
or U2366 (N_2366,N_1551,N_1787);
and U2367 (N_2367,N_2151,N_1775);
nor U2368 (N_2368,N_2028,N_1776);
and U2369 (N_2369,N_1707,N_1792);
nand U2370 (N_2370,N_1582,N_1717);
or U2371 (N_2371,N_1839,N_2076);
and U2372 (N_2372,N_1786,N_1541);
and U2373 (N_2373,N_1930,N_1737);
and U2374 (N_2374,N_1832,N_1573);
and U2375 (N_2375,N_1929,N_1759);
nor U2376 (N_2376,N_1923,N_1892);
or U2377 (N_2377,N_1628,N_2185);
nand U2378 (N_2378,N_2230,N_1870);
and U2379 (N_2379,N_2223,N_2104);
nand U2380 (N_2380,N_2114,N_1729);
and U2381 (N_2381,N_1873,N_1882);
or U2382 (N_2382,N_1511,N_1546);
or U2383 (N_2383,N_2133,N_1519);
nor U2384 (N_2384,N_1815,N_1897);
nor U2385 (N_2385,N_1977,N_1782);
and U2386 (N_2386,N_1654,N_1615);
nand U2387 (N_2387,N_2031,N_1992);
or U2388 (N_2388,N_2166,N_1614);
or U2389 (N_2389,N_2237,N_1934);
or U2390 (N_2390,N_1953,N_2162);
and U2391 (N_2391,N_2177,N_2058);
and U2392 (N_2392,N_1568,N_1922);
nand U2393 (N_2393,N_2129,N_1752);
and U2394 (N_2394,N_1595,N_2210);
or U2395 (N_2395,N_2143,N_1604);
or U2396 (N_2396,N_2024,N_1621);
nor U2397 (N_2397,N_2193,N_2150);
nand U2398 (N_2398,N_2113,N_1652);
or U2399 (N_2399,N_1646,N_2226);
nor U2400 (N_2400,N_1952,N_2218);
nor U2401 (N_2401,N_1927,N_1734);
nor U2402 (N_2402,N_1824,N_1702);
nand U2403 (N_2403,N_1843,N_2057);
nand U2404 (N_2404,N_1690,N_2198);
and U2405 (N_2405,N_2149,N_1940);
nor U2406 (N_2406,N_1635,N_1547);
or U2407 (N_2407,N_1569,N_1823);
or U2408 (N_2408,N_2209,N_2040);
nand U2409 (N_2409,N_1570,N_1762);
nor U2410 (N_2410,N_2219,N_2232);
and U2411 (N_2411,N_1583,N_1668);
or U2412 (N_2412,N_1742,N_1755);
nand U2413 (N_2413,N_1505,N_2027);
or U2414 (N_2414,N_1806,N_2064);
nor U2415 (N_2415,N_2214,N_1735);
nor U2416 (N_2416,N_1849,N_1944);
nor U2417 (N_2417,N_1585,N_1515);
nor U2418 (N_2418,N_2126,N_2164);
nand U2419 (N_2419,N_2007,N_1916);
nor U2420 (N_2420,N_1523,N_1956);
and U2421 (N_2421,N_2173,N_1777);
nand U2422 (N_2422,N_1831,N_2026);
and U2423 (N_2423,N_1687,N_2012);
nor U2424 (N_2424,N_1914,N_1783);
and U2425 (N_2425,N_1758,N_2035);
and U2426 (N_2426,N_2171,N_1833);
and U2427 (N_2427,N_1554,N_1639);
or U2428 (N_2428,N_1679,N_1716);
or U2429 (N_2429,N_1521,N_1761);
and U2430 (N_2430,N_2068,N_1543);
nor U2431 (N_2431,N_1921,N_1804);
nand U2432 (N_2432,N_1670,N_1724);
nand U2433 (N_2433,N_2183,N_2142);
nor U2434 (N_2434,N_2158,N_1503);
xnor U2435 (N_2435,N_1589,N_2059);
or U2436 (N_2436,N_1968,N_2154);
and U2437 (N_2437,N_2135,N_1671);
or U2438 (N_2438,N_2205,N_1803);
and U2439 (N_2439,N_2013,N_1691);
and U2440 (N_2440,N_2112,N_1801);
or U2441 (N_2441,N_1991,N_1958);
and U2442 (N_2442,N_1860,N_1681);
and U2443 (N_2443,N_1821,N_1522);
and U2444 (N_2444,N_2099,N_1666);
and U2445 (N_2445,N_1893,N_1591);
and U2446 (N_2446,N_1542,N_2245);
or U2447 (N_2447,N_2175,N_1842);
nand U2448 (N_2448,N_1788,N_1565);
or U2449 (N_2449,N_1730,N_1814);
or U2450 (N_2450,N_1906,N_1979);
nand U2451 (N_2451,N_1699,N_1722);
or U2452 (N_2452,N_1810,N_2090);
and U2453 (N_2453,N_1705,N_1745);
or U2454 (N_2454,N_2196,N_2191);
or U2455 (N_2455,N_1816,N_2157);
or U2456 (N_2456,N_1910,N_2174);
nand U2457 (N_2457,N_2042,N_1872);
nor U2458 (N_2458,N_1718,N_1989);
nand U2459 (N_2459,N_1509,N_1550);
nor U2460 (N_2460,N_1795,N_1869);
and U2461 (N_2461,N_1659,N_1969);
nand U2462 (N_2462,N_1763,N_1822);
and U2463 (N_2463,N_1698,N_2120);
or U2464 (N_2464,N_2137,N_1983);
and U2465 (N_2465,N_1905,N_1884);
nor U2466 (N_2466,N_2086,N_2056);
or U2467 (N_2467,N_2213,N_2212);
nor U2468 (N_2468,N_1749,N_1701);
and U2469 (N_2469,N_2221,N_1609);
nand U2470 (N_2470,N_1641,N_2023);
and U2471 (N_2471,N_1606,N_2122);
nor U2472 (N_2472,N_1588,N_2246);
nor U2473 (N_2473,N_1611,N_1517);
or U2474 (N_2474,N_1688,N_1732);
nand U2475 (N_2475,N_1813,N_1579);
nand U2476 (N_2476,N_2078,N_2203);
or U2477 (N_2477,N_1607,N_2029);
and U2478 (N_2478,N_1682,N_1778);
or U2479 (N_2479,N_1653,N_1950);
or U2480 (N_2480,N_2217,N_1683);
and U2481 (N_2481,N_1891,N_1684);
nand U2482 (N_2482,N_1625,N_2156);
nor U2483 (N_2483,N_1826,N_1695);
or U2484 (N_2484,N_1750,N_1504);
and U2485 (N_2485,N_2017,N_1678);
nand U2486 (N_2486,N_1932,N_1632);
and U2487 (N_2487,N_1998,N_1651);
or U2488 (N_2488,N_1644,N_2202);
nand U2489 (N_2489,N_1894,N_2170);
nand U2490 (N_2490,N_2110,N_1720);
nor U2491 (N_2491,N_1712,N_2021);
or U2492 (N_2492,N_1634,N_1941);
nor U2493 (N_2493,N_2244,N_2052);
and U2494 (N_2494,N_2178,N_2100);
nand U2495 (N_2495,N_1807,N_2010);
nand U2496 (N_2496,N_2000,N_1946);
nand U2497 (N_2497,N_2071,N_2051);
and U2498 (N_2498,N_1587,N_2206);
nor U2499 (N_2499,N_1726,N_2225);
or U2500 (N_2500,N_2161,N_1571);
and U2501 (N_2501,N_2118,N_2241);
or U2502 (N_2502,N_1528,N_1971);
nor U2503 (N_2503,N_2146,N_1774);
and U2504 (N_2504,N_1513,N_1797);
nand U2505 (N_2505,N_1692,N_1638);
or U2506 (N_2506,N_1854,N_1748);
or U2507 (N_2507,N_1630,N_1731);
and U2508 (N_2508,N_1627,N_2236);
nor U2509 (N_2509,N_1709,N_1626);
nor U2510 (N_2510,N_2231,N_1954);
nand U2511 (N_2511,N_2188,N_1616);
or U2512 (N_2512,N_1602,N_1984);
nor U2513 (N_2513,N_2172,N_2132);
or U2514 (N_2514,N_1648,N_2163);
nand U2515 (N_2515,N_1618,N_1577);
or U2516 (N_2516,N_2108,N_2189);
nor U2517 (N_2517,N_1764,N_1943);
nor U2518 (N_2518,N_1871,N_2008);
and U2519 (N_2519,N_2169,N_1899);
nor U2520 (N_2520,N_1613,N_1901);
nor U2521 (N_2521,N_1864,N_2111);
or U2522 (N_2522,N_1995,N_1643);
and U2523 (N_2523,N_1693,N_1715);
or U2524 (N_2524,N_1710,N_1772);
and U2525 (N_2525,N_1933,N_2168);
and U2526 (N_2526,N_1896,N_2072);
nand U2527 (N_2527,N_1911,N_2123);
or U2528 (N_2528,N_1512,N_1633);
nor U2529 (N_2529,N_2222,N_2018);
or U2530 (N_2530,N_1680,N_1673);
and U2531 (N_2531,N_1982,N_2094);
nor U2532 (N_2532,N_1578,N_2055);
and U2533 (N_2533,N_1769,N_2074);
and U2534 (N_2534,N_2130,N_1903);
nor U2535 (N_2535,N_2147,N_1617);
nor U2536 (N_2536,N_1949,N_1593);
nand U2537 (N_2537,N_1544,N_2192);
nor U2538 (N_2538,N_2103,N_1836);
and U2539 (N_2539,N_1840,N_1642);
nand U2540 (N_2540,N_1536,N_2121);
nor U2541 (N_2541,N_1708,N_1567);
nand U2542 (N_2542,N_1898,N_2084);
nor U2543 (N_2543,N_2079,N_2109);
nand U2544 (N_2544,N_2041,N_2176);
or U2545 (N_2545,N_2119,N_1852);
nor U2546 (N_2546,N_1637,N_1866);
and U2547 (N_2547,N_1865,N_1553);
and U2548 (N_2548,N_2082,N_2044);
and U2549 (N_2549,N_2005,N_1622);
or U2550 (N_2550,N_1685,N_1879);
nand U2551 (N_2551,N_2116,N_2215);
or U2552 (N_2552,N_1649,N_2182);
and U2553 (N_2553,N_1800,N_2233);
nand U2554 (N_2554,N_2054,N_2224);
nor U2555 (N_2555,N_2184,N_1516);
or U2556 (N_2556,N_2025,N_1848);
nor U2557 (N_2557,N_1889,N_1572);
nand U2558 (N_2558,N_1696,N_1868);
or U2559 (N_2559,N_1723,N_2088);
nor U2560 (N_2560,N_1686,N_2194);
and U2561 (N_2561,N_1985,N_1959);
nand U2562 (N_2562,N_1976,N_1562);
nor U2563 (N_2563,N_1861,N_2207);
or U2564 (N_2564,N_2138,N_1549);
nand U2565 (N_2565,N_1994,N_2200);
nor U2566 (N_2566,N_1689,N_2065);
and U2567 (N_2567,N_1820,N_1844);
nand U2568 (N_2568,N_1812,N_1817);
nor U2569 (N_2569,N_1768,N_1552);
or U2570 (N_2570,N_2069,N_1890);
nand U2571 (N_2571,N_2022,N_1867);
nand U2572 (N_2572,N_1948,N_1997);
nand U2573 (N_2573,N_1658,N_1883);
or U2574 (N_2574,N_1970,N_1580);
and U2575 (N_2575,N_1900,N_1603);
or U2576 (N_2576,N_1912,N_1863);
and U2577 (N_2577,N_1576,N_2160);
or U2578 (N_2578,N_1538,N_1675);
or U2579 (N_2579,N_2167,N_2045);
nor U2580 (N_2580,N_1548,N_1559);
nand U2581 (N_2581,N_2038,N_1741);
or U2582 (N_2582,N_1965,N_1676);
or U2583 (N_2583,N_2048,N_1555);
or U2584 (N_2584,N_2014,N_1928);
nand U2585 (N_2585,N_1725,N_2155);
or U2586 (N_2586,N_1563,N_2211);
nor U2587 (N_2587,N_2053,N_1533);
or U2588 (N_2588,N_2227,N_1880);
xnor U2589 (N_2589,N_1664,N_1862);
nand U2590 (N_2590,N_1564,N_1510);
and U2591 (N_2591,N_1828,N_2186);
nand U2592 (N_2592,N_1951,N_1955);
and U2593 (N_2593,N_1594,N_2102);
nand U2594 (N_2594,N_2248,N_1660);
nor U2595 (N_2595,N_1612,N_1874);
and U2596 (N_2596,N_1545,N_2197);
nor U2597 (N_2597,N_1773,N_1915);
and U2598 (N_2598,N_1986,N_2049);
and U2599 (N_2599,N_1967,N_2092);
nor U2600 (N_2600,N_1736,N_1751);
and U2601 (N_2601,N_1586,N_1740);
and U2602 (N_2602,N_2089,N_2091);
nand U2603 (N_2603,N_1877,N_1599);
or U2604 (N_2604,N_1743,N_1838);
and U2605 (N_2605,N_1514,N_1975);
nand U2606 (N_2606,N_1636,N_1656);
and U2607 (N_2607,N_1663,N_2009);
nand U2608 (N_2608,N_2165,N_2159);
xor U2609 (N_2609,N_2001,N_1655);
nand U2610 (N_2610,N_2127,N_1791);
nor U2611 (N_2611,N_1697,N_2015);
nor U2612 (N_2612,N_2187,N_2105);
and U2613 (N_2613,N_1908,N_2249);
and U2614 (N_2614,N_1721,N_1856);
and U2615 (N_2615,N_2047,N_2030);
or U2616 (N_2616,N_2128,N_2239);
or U2617 (N_2617,N_1694,N_1936);
nand U2618 (N_2618,N_1574,N_2061);
nand U2619 (N_2619,N_1790,N_1794);
nand U2620 (N_2620,N_1924,N_1744);
or U2621 (N_2621,N_1793,N_1830);
nand U2622 (N_2622,N_1520,N_2067);
or U2623 (N_2623,N_1770,N_2077);
xor U2624 (N_2624,N_1631,N_1575);
and U2625 (N_2625,N_2019,N_1576);
and U2626 (N_2626,N_2088,N_2094);
and U2627 (N_2627,N_1632,N_1622);
nor U2628 (N_2628,N_1683,N_1590);
and U2629 (N_2629,N_1838,N_2062);
and U2630 (N_2630,N_1676,N_2135);
and U2631 (N_2631,N_1912,N_1902);
and U2632 (N_2632,N_1760,N_1928);
nand U2633 (N_2633,N_1800,N_2124);
xnor U2634 (N_2634,N_1861,N_1958);
nor U2635 (N_2635,N_2147,N_1771);
or U2636 (N_2636,N_1942,N_2075);
nand U2637 (N_2637,N_2035,N_1770);
nand U2638 (N_2638,N_1742,N_1975);
nor U2639 (N_2639,N_2132,N_1735);
or U2640 (N_2640,N_1970,N_1712);
or U2641 (N_2641,N_1822,N_2039);
nand U2642 (N_2642,N_1973,N_1791);
nand U2643 (N_2643,N_1512,N_2189);
nor U2644 (N_2644,N_2177,N_2217);
and U2645 (N_2645,N_1769,N_1595);
nand U2646 (N_2646,N_1572,N_1668);
and U2647 (N_2647,N_1590,N_2182);
and U2648 (N_2648,N_2192,N_1882);
nor U2649 (N_2649,N_1541,N_1796);
and U2650 (N_2650,N_1541,N_2016);
or U2651 (N_2651,N_2167,N_1966);
nor U2652 (N_2652,N_1932,N_1508);
xor U2653 (N_2653,N_1738,N_1564);
or U2654 (N_2654,N_2241,N_1826);
nor U2655 (N_2655,N_1958,N_1736);
nand U2656 (N_2656,N_1737,N_2040);
and U2657 (N_2657,N_2122,N_2082);
nor U2658 (N_2658,N_1934,N_2099);
nor U2659 (N_2659,N_2213,N_2135);
and U2660 (N_2660,N_2041,N_2072);
nand U2661 (N_2661,N_1856,N_1886);
xnor U2662 (N_2662,N_1898,N_1702);
or U2663 (N_2663,N_2241,N_1657);
nand U2664 (N_2664,N_1930,N_1872);
and U2665 (N_2665,N_2049,N_1946);
nand U2666 (N_2666,N_1967,N_1597);
or U2667 (N_2667,N_1574,N_2009);
or U2668 (N_2668,N_1908,N_1868);
xor U2669 (N_2669,N_1659,N_2005);
and U2670 (N_2670,N_1987,N_2231);
nand U2671 (N_2671,N_1685,N_1938);
and U2672 (N_2672,N_1637,N_2060);
or U2673 (N_2673,N_1924,N_1907);
and U2674 (N_2674,N_1957,N_2067);
or U2675 (N_2675,N_1900,N_1659);
or U2676 (N_2676,N_1533,N_1560);
nor U2677 (N_2677,N_1611,N_2145);
nor U2678 (N_2678,N_1680,N_2229);
nor U2679 (N_2679,N_1527,N_1730);
nor U2680 (N_2680,N_1634,N_1648);
xnor U2681 (N_2681,N_2050,N_1644);
or U2682 (N_2682,N_1890,N_1583);
or U2683 (N_2683,N_1661,N_2243);
or U2684 (N_2684,N_1662,N_1787);
nand U2685 (N_2685,N_2212,N_1839);
nor U2686 (N_2686,N_1700,N_1948);
nor U2687 (N_2687,N_2190,N_1695);
and U2688 (N_2688,N_2063,N_1984);
or U2689 (N_2689,N_1938,N_1937);
nand U2690 (N_2690,N_1594,N_1828);
and U2691 (N_2691,N_1653,N_2067);
and U2692 (N_2692,N_1855,N_1995);
nor U2693 (N_2693,N_1905,N_1695);
nand U2694 (N_2694,N_1947,N_2247);
or U2695 (N_2695,N_1607,N_1970);
nor U2696 (N_2696,N_2176,N_2183);
nor U2697 (N_2697,N_2163,N_1927);
nand U2698 (N_2698,N_1545,N_1988);
or U2699 (N_2699,N_1871,N_1765);
and U2700 (N_2700,N_2211,N_1887);
nor U2701 (N_2701,N_2235,N_1686);
nor U2702 (N_2702,N_2117,N_1726);
and U2703 (N_2703,N_1797,N_1860);
and U2704 (N_2704,N_2194,N_2056);
or U2705 (N_2705,N_1524,N_2070);
nand U2706 (N_2706,N_1502,N_2148);
and U2707 (N_2707,N_1884,N_1767);
and U2708 (N_2708,N_1814,N_2131);
and U2709 (N_2709,N_2159,N_1799);
nand U2710 (N_2710,N_2066,N_1738);
nor U2711 (N_2711,N_2176,N_1501);
or U2712 (N_2712,N_2209,N_2226);
or U2713 (N_2713,N_1705,N_2184);
nand U2714 (N_2714,N_1782,N_1828);
or U2715 (N_2715,N_1943,N_2062);
or U2716 (N_2716,N_2061,N_1931);
or U2717 (N_2717,N_1789,N_1886);
and U2718 (N_2718,N_1567,N_1528);
nand U2719 (N_2719,N_2249,N_1564);
and U2720 (N_2720,N_1894,N_1522);
and U2721 (N_2721,N_1954,N_1814);
or U2722 (N_2722,N_2148,N_1919);
or U2723 (N_2723,N_1689,N_2176);
or U2724 (N_2724,N_1721,N_2073);
xnor U2725 (N_2725,N_2114,N_1547);
or U2726 (N_2726,N_1523,N_1741);
or U2727 (N_2727,N_1635,N_1662);
nand U2728 (N_2728,N_1542,N_2092);
and U2729 (N_2729,N_1688,N_1540);
nand U2730 (N_2730,N_2086,N_2249);
nand U2731 (N_2731,N_1602,N_2073);
or U2732 (N_2732,N_2227,N_1575);
and U2733 (N_2733,N_1619,N_2107);
and U2734 (N_2734,N_1773,N_2198);
nand U2735 (N_2735,N_1945,N_2052);
or U2736 (N_2736,N_2171,N_1800);
nor U2737 (N_2737,N_1698,N_1782);
nand U2738 (N_2738,N_1551,N_1933);
nand U2739 (N_2739,N_2161,N_2063);
nor U2740 (N_2740,N_2016,N_1916);
xnor U2741 (N_2741,N_1599,N_2205);
and U2742 (N_2742,N_1776,N_1698);
nand U2743 (N_2743,N_1935,N_1679);
nor U2744 (N_2744,N_2232,N_2025);
nor U2745 (N_2745,N_1555,N_1616);
and U2746 (N_2746,N_1758,N_1838);
nor U2747 (N_2747,N_2061,N_1971);
and U2748 (N_2748,N_1853,N_1586);
nor U2749 (N_2749,N_2122,N_1835);
or U2750 (N_2750,N_1887,N_2021);
and U2751 (N_2751,N_1975,N_1726);
or U2752 (N_2752,N_1814,N_1671);
or U2753 (N_2753,N_2060,N_1861);
and U2754 (N_2754,N_1593,N_1713);
xnor U2755 (N_2755,N_1592,N_2138);
nor U2756 (N_2756,N_1963,N_1987);
and U2757 (N_2757,N_1790,N_1797);
nor U2758 (N_2758,N_2228,N_2175);
nor U2759 (N_2759,N_1990,N_1580);
nand U2760 (N_2760,N_1988,N_1767);
nor U2761 (N_2761,N_2065,N_2169);
nor U2762 (N_2762,N_1700,N_1568);
or U2763 (N_2763,N_2113,N_1858);
nand U2764 (N_2764,N_1766,N_2057);
nor U2765 (N_2765,N_1648,N_1837);
and U2766 (N_2766,N_1742,N_1841);
nand U2767 (N_2767,N_1977,N_2132);
or U2768 (N_2768,N_2095,N_1521);
xor U2769 (N_2769,N_1682,N_2113);
xnor U2770 (N_2770,N_1683,N_2011);
nand U2771 (N_2771,N_1622,N_2227);
nor U2772 (N_2772,N_1722,N_1615);
nor U2773 (N_2773,N_1845,N_1699);
and U2774 (N_2774,N_1860,N_2064);
nor U2775 (N_2775,N_1682,N_1830);
and U2776 (N_2776,N_2145,N_1500);
nor U2777 (N_2777,N_2183,N_1969);
nor U2778 (N_2778,N_2068,N_1898);
or U2779 (N_2779,N_1965,N_1654);
and U2780 (N_2780,N_1607,N_1877);
nand U2781 (N_2781,N_1671,N_2219);
or U2782 (N_2782,N_2180,N_1951);
nor U2783 (N_2783,N_2009,N_1851);
or U2784 (N_2784,N_1534,N_1576);
and U2785 (N_2785,N_1677,N_1852);
xor U2786 (N_2786,N_1837,N_2121);
or U2787 (N_2787,N_2013,N_2058);
nor U2788 (N_2788,N_1760,N_1620);
nor U2789 (N_2789,N_1611,N_2224);
or U2790 (N_2790,N_2032,N_1858);
and U2791 (N_2791,N_2056,N_2112);
nand U2792 (N_2792,N_1716,N_2056);
and U2793 (N_2793,N_1804,N_1954);
nand U2794 (N_2794,N_1645,N_2009);
or U2795 (N_2795,N_1528,N_1917);
or U2796 (N_2796,N_2173,N_1810);
nor U2797 (N_2797,N_2050,N_1974);
or U2798 (N_2798,N_1822,N_2248);
and U2799 (N_2799,N_1963,N_1562);
nand U2800 (N_2800,N_1738,N_1654);
xnor U2801 (N_2801,N_1583,N_2074);
or U2802 (N_2802,N_1990,N_1650);
and U2803 (N_2803,N_2145,N_1855);
and U2804 (N_2804,N_2169,N_2151);
nand U2805 (N_2805,N_2093,N_1825);
or U2806 (N_2806,N_1520,N_1785);
or U2807 (N_2807,N_1897,N_2001);
or U2808 (N_2808,N_2008,N_2150);
nor U2809 (N_2809,N_2124,N_1979);
or U2810 (N_2810,N_1691,N_1938);
nand U2811 (N_2811,N_1813,N_1980);
nand U2812 (N_2812,N_1557,N_1865);
or U2813 (N_2813,N_2108,N_1893);
nand U2814 (N_2814,N_1624,N_1746);
or U2815 (N_2815,N_1657,N_1974);
or U2816 (N_2816,N_1943,N_2244);
nor U2817 (N_2817,N_2176,N_2013);
nand U2818 (N_2818,N_1975,N_1879);
or U2819 (N_2819,N_1715,N_2213);
and U2820 (N_2820,N_2141,N_2192);
nand U2821 (N_2821,N_1510,N_2013);
or U2822 (N_2822,N_1603,N_1572);
or U2823 (N_2823,N_2123,N_1953);
and U2824 (N_2824,N_1658,N_1628);
and U2825 (N_2825,N_2217,N_1861);
or U2826 (N_2826,N_1835,N_1586);
nor U2827 (N_2827,N_1784,N_2050);
nand U2828 (N_2828,N_1927,N_2004);
nand U2829 (N_2829,N_2164,N_1872);
nand U2830 (N_2830,N_2249,N_1741);
nor U2831 (N_2831,N_2104,N_1761);
or U2832 (N_2832,N_2117,N_1589);
and U2833 (N_2833,N_1961,N_2118);
or U2834 (N_2834,N_2232,N_1689);
or U2835 (N_2835,N_1639,N_1746);
or U2836 (N_2836,N_2207,N_2066);
xor U2837 (N_2837,N_2084,N_1559);
or U2838 (N_2838,N_1683,N_1639);
nand U2839 (N_2839,N_2068,N_1546);
nand U2840 (N_2840,N_1504,N_1929);
nand U2841 (N_2841,N_2181,N_1823);
nor U2842 (N_2842,N_2243,N_2226);
nand U2843 (N_2843,N_2153,N_1755);
or U2844 (N_2844,N_2183,N_2198);
nor U2845 (N_2845,N_2067,N_1900);
nor U2846 (N_2846,N_1621,N_1691);
xnor U2847 (N_2847,N_1585,N_2117);
or U2848 (N_2848,N_1874,N_2190);
or U2849 (N_2849,N_1621,N_2198);
nor U2850 (N_2850,N_1816,N_2084);
and U2851 (N_2851,N_1800,N_2098);
nor U2852 (N_2852,N_2198,N_2118);
or U2853 (N_2853,N_2042,N_1983);
nor U2854 (N_2854,N_2130,N_2181);
nand U2855 (N_2855,N_2018,N_1530);
nand U2856 (N_2856,N_2015,N_1616);
or U2857 (N_2857,N_1572,N_1569);
nor U2858 (N_2858,N_2233,N_1735);
and U2859 (N_2859,N_1806,N_2072);
or U2860 (N_2860,N_1546,N_1518);
or U2861 (N_2861,N_1909,N_1580);
nand U2862 (N_2862,N_2162,N_1699);
nor U2863 (N_2863,N_2108,N_1536);
and U2864 (N_2864,N_2066,N_1775);
or U2865 (N_2865,N_2092,N_1646);
nor U2866 (N_2866,N_2014,N_1897);
or U2867 (N_2867,N_1856,N_1549);
nand U2868 (N_2868,N_1632,N_1725);
or U2869 (N_2869,N_1729,N_1959);
nand U2870 (N_2870,N_1815,N_1559);
and U2871 (N_2871,N_1518,N_1579);
and U2872 (N_2872,N_1847,N_1942);
nand U2873 (N_2873,N_1646,N_2020);
and U2874 (N_2874,N_1848,N_2163);
or U2875 (N_2875,N_1623,N_1547);
or U2876 (N_2876,N_1574,N_1747);
and U2877 (N_2877,N_1510,N_1652);
nor U2878 (N_2878,N_1914,N_2229);
and U2879 (N_2879,N_2171,N_1929);
and U2880 (N_2880,N_1900,N_2190);
nor U2881 (N_2881,N_1761,N_1683);
nand U2882 (N_2882,N_1658,N_1923);
nor U2883 (N_2883,N_1905,N_2091);
or U2884 (N_2884,N_2096,N_2012);
xnor U2885 (N_2885,N_1790,N_1519);
or U2886 (N_2886,N_1706,N_1897);
nor U2887 (N_2887,N_1996,N_1797);
nand U2888 (N_2888,N_2063,N_1587);
or U2889 (N_2889,N_1592,N_1754);
nor U2890 (N_2890,N_1903,N_1609);
nor U2891 (N_2891,N_1735,N_2090);
nand U2892 (N_2892,N_1795,N_1984);
nand U2893 (N_2893,N_1662,N_1652);
nor U2894 (N_2894,N_2086,N_2131);
and U2895 (N_2895,N_1943,N_1542);
nand U2896 (N_2896,N_2120,N_1712);
or U2897 (N_2897,N_2024,N_2033);
nor U2898 (N_2898,N_2068,N_2218);
and U2899 (N_2899,N_1686,N_2179);
nand U2900 (N_2900,N_2168,N_1611);
nor U2901 (N_2901,N_1667,N_1976);
nor U2902 (N_2902,N_1722,N_1737);
nor U2903 (N_2903,N_1995,N_1709);
nor U2904 (N_2904,N_1951,N_2198);
or U2905 (N_2905,N_1628,N_1795);
and U2906 (N_2906,N_1611,N_1555);
nand U2907 (N_2907,N_1642,N_1792);
or U2908 (N_2908,N_2196,N_1522);
or U2909 (N_2909,N_1677,N_1552);
or U2910 (N_2910,N_1743,N_2089);
or U2911 (N_2911,N_2153,N_1979);
nor U2912 (N_2912,N_1899,N_2067);
or U2913 (N_2913,N_1857,N_1554);
nand U2914 (N_2914,N_1579,N_2140);
or U2915 (N_2915,N_1500,N_1992);
and U2916 (N_2916,N_2076,N_2246);
or U2917 (N_2917,N_1846,N_1534);
nor U2918 (N_2918,N_1506,N_1789);
and U2919 (N_2919,N_1848,N_2067);
nand U2920 (N_2920,N_1693,N_1861);
nor U2921 (N_2921,N_1753,N_1843);
nand U2922 (N_2922,N_1947,N_1789);
nand U2923 (N_2923,N_1690,N_1798);
nor U2924 (N_2924,N_2045,N_2178);
nand U2925 (N_2925,N_1676,N_1796);
nor U2926 (N_2926,N_1701,N_2075);
and U2927 (N_2927,N_2000,N_1993);
or U2928 (N_2928,N_1745,N_1727);
and U2929 (N_2929,N_1890,N_2139);
and U2930 (N_2930,N_1981,N_1990);
nand U2931 (N_2931,N_2151,N_2197);
and U2932 (N_2932,N_1636,N_2163);
nand U2933 (N_2933,N_2167,N_1601);
xnor U2934 (N_2934,N_1696,N_2214);
and U2935 (N_2935,N_1735,N_2140);
nor U2936 (N_2936,N_1645,N_2022);
nand U2937 (N_2937,N_1968,N_2010);
nor U2938 (N_2938,N_1604,N_2210);
or U2939 (N_2939,N_1922,N_1823);
and U2940 (N_2940,N_1821,N_1851);
and U2941 (N_2941,N_1978,N_1656);
nand U2942 (N_2942,N_1572,N_1592);
nand U2943 (N_2943,N_2241,N_1980);
or U2944 (N_2944,N_2134,N_1869);
or U2945 (N_2945,N_2130,N_2166);
nand U2946 (N_2946,N_2245,N_1955);
nor U2947 (N_2947,N_1599,N_1809);
nand U2948 (N_2948,N_1866,N_1640);
nand U2949 (N_2949,N_1599,N_2092);
and U2950 (N_2950,N_1645,N_1549);
nand U2951 (N_2951,N_2078,N_1636);
nand U2952 (N_2952,N_1974,N_1619);
nand U2953 (N_2953,N_1821,N_2141);
or U2954 (N_2954,N_2222,N_1698);
and U2955 (N_2955,N_2094,N_2032);
nor U2956 (N_2956,N_1911,N_1723);
and U2957 (N_2957,N_1588,N_1716);
nand U2958 (N_2958,N_1604,N_1590);
and U2959 (N_2959,N_2220,N_1626);
and U2960 (N_2960,N_2160,N_2197);
nand U2961 (N_2961,N_2055,N_1935);
nand U2962 (N_2962,N_1872,N_1938);
or U2963 (N_2963,N_1778,N_1707);
and U2964 (N_2964,N_1995,N_1810);
nor U2965 (N_2965,N_1596,N_2084);
and U2966 (N_2966,N_1762,N_1839);
nor U2967 (N_2967,N_2137,N_1987);
nor U2968 (N_2968,N_2173,N_1551);
and U2969 (N_2969,N_1575,N_2163);
nand U2970 (N_2970,N_1653,N_1946);
and U2971 (N_2971,N_1797,N_2004);
or U2972 (N_2972,N_2036,N_2035);
and U2973 (N_2973,N_1656,N_1942);
xor U2974 (N_2974,N_2054,N_2206);
and U2975 (N_2975,N_1540,N_1559);
nand U2976 (N_2976,N_1970,N_2214);
and U2977 (N_2977,N_2182,N_1794);
nand U2978 (N_2978,N_1831,N_1515);
or U2979 (N_2979,N_2010,N_1875);
or U2980 (N_2980,N_1654,N_1930);
or U2981 (N_2981,N_2088,N_1772);
and U2982 (N_2982,N_2011,N_1839);
and U2983 (N_2983,N_1917,N_1708);
and U2984 (N_2984,N_2020,N_1616);
or U2985 (N_2985,N_1782,N_1952);
and U2986 (N_2986,N_1699,N_1686);
nand U2987 (N_2987,N_1885,N_1967);
nand U2988 (N_2988,N_1870,N_1964);
xnor U2989 (N_2989,N_2200,N_1901);
nor U2990 (N_2990,N_2075,N_2184);
and U2991 (N_2991,N_1501,N_1605);
or U2992 (N_2992,N_2172,N_1555);
and U2993 (N_2993,N_2235,N_1784);
or U2994 (N_2994,N_1670,N_1514);
nand U2995 (N_2995,N_1752,N_1606);
or U2996 (N_2996,N_1959,N_1611);
nor U2997 (N_2997,N_1932,N_1859);
or U2998 (N_2998,N_1541,N_1625);
or U2999 (N_2999,N_1651,N_1686);
nand UO_0 (O_0,N_2269,N_2889);
and UO_1 (O_1,N_2766,N_2966);
or UO_2 (O_2,N_2749,N_2634);
xor UO_3 (O_3,N_2651,N_2383);
nand UO_4 (O_4,N_2747,N_2828);
nand UO_5 (O_5,N_2457,N_2489);
and UO_6 (O_6,N_2675,N_2934);
nor UO_7 (O_7,N_2759,N_2379);
and UO_8 (O_8,N_2527,N_2583);
nor UO_9 (O_9,N_2326,N_2969);
nand UO_10 (O_10,N_2328,N_2382);
or UO_11 (O_11,N_2504,N_2450);
nand UO_12 (O_12,N_2369,N_2312);
or UO_13 (O_13,N_2514,N_2748);
nand UO_14 (O_14,N_2351,N_2962);
or UO_15 (O_15,N_2851,N_2721);
or UO_16 (O_16,N_2327,N_2316);
nor UO_17 (O_17,N_2516,N_2998);
nand UO_18 (O_18,N_2591,N_2842);
and UO_19 (O_19,N_2637,N_2510);
nand UO_20 (O_20,N_2465,N_2983);
or UO_21 (O_21,N_2488,N_2371);
and UO_22 (O_22,N_2908,N_2476);
nor UO_23 (O_23,N_2907,N_2713);
nor UO_24 (O_24,N_2859,N_2306);
and UO_25 (O_25,N_2439,N_2730);
or UO_26 (O_26,N_2917,N_2463);
and UO_27 (O_27,N_2252,N_2796);
nand UO_28 (O_28,N_2590,N_2528);
nand UO_29 (O_29,N_2370,N_2911);
nor UO_30 (O_30,N_2360,N_2404);
nor UO_31 (O_31,N_2873,N_2636);
and UO_32 (O_32,N_2830,N_2879);
and UO_33 (O_33,N_2607,N_2625);
nand UO_34 (O_34,N_2319,N_2857);
and UO_35 (O_35,N_2897,N_2297);
or UO_36 (O_36,N_2931,N_2501);
nor UO_37 (O_37,N_2276,N_2596);
or UO_38 (O_38,N_2301,N_2820);
nor UO_39 (O_39,N_2535,N_2380);
or UO_40 (O_40,N_2615,N_2323);
or UO_41 (O_41,N_2937,N_2333);
nor UO_42 (O_42,N_2423,N_2671);
and UO_43 (O_43,N_2490,N_2373);
nand UO_44 (O_44,N_2774,N_2487);
nand UO_45 (O_45,N_2734,N_2445);
nor UO_46 (O_46,N_2768,N_2581);
nor UO_47 (O_47,N_2354,N_2847);
xnor UO_48 (O_48,N_2781,N_2638);
or UO_49 (O_49,N_2814,N_2999);
or UO_50 (O_50,N_2494,N_2268);
or UO_51 (O_51,N_2324,N_2309);
nor UO_52 (O_52,N_2714,N_2650);
nand UO_53 (O_53,N_2677,N_2901);
nand UO_54 (O_54,N_2341,N_2994);
nor UO_55 (O_55,N_2692,N_2419);
or UO_56 (O_56,N_2853,N_2756);
nand UO_57 (O_57,N_2807,N_2803);
xor UO_58 (O_58,N_2944,N_2927);
or UO_59 (O_59,N_2719,N_2702);
nor UO_60 (O_60,N_2732,N_2364);
or UO_61 (O_61,N_2770,N_2933);
or UO_62 (O_62,N_2881,N_2526);
nand UO_63 (O_63,N_2669,N_2554);
nor UO_64 (O_64,N_2874,N_2819);
or UO_65 (O_65,N_2695,N_2443);
and UO_66 (O_66,N_2357,N_2551);
and UO_67 (O_67,N_2885,N_2464);
xnor UO_68 (O_68,N_2542,N_2468);
and UO_69 (O_69,N_2270,N_2699);
and UO_70 (O_70,N_2684,N_2777);
or UO_71 (O_71,N_2837,N_2871);
nor UO_72 (O_72,N_2658,N_2545);
nor UO_73 (O_73,N_2454,N_2473);
nand UO_74 (O_74,N_2751,N_2785);
nor UO_75 (O_75,N_2821,N_2624);
nand UO_76 (O_76,N_2924,N_2363);
or UO_77 (O_77,N_2775,N_2530);
or UO_78 (O_78,N_2486,N_2308);
nand UO_79 (O_79,N_2891,N_2930);
nor UO_80 (O_80,N_2282,N_2986);
nor UO_81 (O_81,N_2393,N_2600);
nor UO_82 (O_82,N_2320,N_2496);
or UO_83 (O_83,N_2469,N_2818);
and UO_84 (O_84,N_2789,N_2797);
nor UO_85 (O_85,N_2694,N_2887);
nand UO_86 (O_86,N_2884,N_2670);
or UO_87 (O_87,N_2880,N_2614);
nor UO_88 (O_88,N_2532,N_2995);
or UO_89 (O_89,N_2295,N_2989);
nand UO_90 (O_90,N_2288,N_2254);
and UO_91 (O_91,N_2745,N_2421);
and UO_92 (O_92,N_2717,N_2343);
nand UO_93 (O_93,N_2648,N_2417);
nand UO_94 (O_94,N_2430,N_2949);
and UO_95 (O_95,N_2575,N_2523);
and UO_96 (O_96,N_2764,N_2864);
nor UO_97 (O_97,N_2723,N_2974);
or UO_98 (O_98,N_2654,N_2704);
nor UO_99 (O_99,N_2334,N_2460);
or UO_100 (O_100,N_2872,N_2381);
nor UO_101 (O_101,N_2398,N_2564);
or UO_102 (O_102,N_2783,N_2665);
nand UO_103 (O_103,N_2414,N_2950);
or UO_104 (O_104,N_2552,N_2757);
nand UO_105 (O_105,N_2302,N_2307);
or UO_106 (O_106,N_2791,N_2432);
or UO_107 (O_107,N_2975,N_2951);
and UO_108 (O_108,N_2505,N_2279);
and UO_109 (O_109,N_2580,N_2503);
nand UO_110 (O_110,N_2941,N_2816);
nand UO_111 (O_111,N_2291,N_2556);
and UO_112 (O_112,N_2394,N_2715);
nor UO_113 (O_113,N_2794,N_2788);
nand UO_114 (O_114,N_2280,N_2863);
nand UO_115 (O_115,N_2411,N_2305);
or UO_116 (O_116,N_2956,N_2661);
or UO_117 (O_117,N_2886,N_2706);
or UO_118 (O_118,N_2303,N_2722);
or UO_119 (O_119,N_2696,N_2627);
and UO_120 (O_120,N_2772,N_2602);
and UO_121 (O_121,N_2619,N_2700);
nor UO_122 (O_122,N_2576,N_2502);
and UO_123 (O_123,N_2338,N_2397);
nor UO_124 (O_124,N_2612,N_2459);
and UO_125 (O_125,N_2982,N_2866);
xnor UO_126 (O_126,N_2736,N_2256);
or UO_127 (O_127,N_2416,N_2954);
nor UO_128 (O_128,N_2562,N_2387);
or UO_129 (O_129,N_2507,N_2399);
xnor UO_130 (O_130,N_2988,N_2711);
nand UO_131 (O_131,N_2913,N_2958);
nor UO_132 (O_132,N_2852,N_2899);
nand UO_133 (O_133,N_2477,N_2547);
and UO_134 (O_134,N_2858,N_2606);
and UO_135 (O_135,N_2574,N_2401);
nor UO_136 (O_136,N_2760,N_2682);
or UO_137 (O_137,N_2836,N_2825);
nand UO_138 (O_138,N_2390,N_2829);
or UO_139 (O_139,N_2346,N_2391);
nor UO_140 (O_140,N_2762,N_2515);
nand UO_141 (O_141,N_2331,N_2442);
and UO_142 (O_142,N_2335,N_2867);
nor UO_143 (O_143,N_2608,N_2639);
nor UO_144 (O_144,N_2412,N_2480);
xor UO_145 (O_145,N_2935,N_2555);
nor UO_146 (O_146,N_2793,N_2928);
nand UO_147 (O_147,N_2257,N_2548);
nor UO_148 (O_148,N_2676,N_2261);
nor UO_149 (O_149,N_2446,N_2926);
or UO_150 (O_150,N_2598,N_2458);
nand UO_151 (O_151,N_2479,N_2623);
nand UO_152 (O_152,N_2895,N_2795);
nor UO_153 (O_153,N_2630,N_2253);
and UO_154 (O_154,N_2260,N_2520);
nand UO_155 (O_155,N_2595,N_2691);
nand UO_156 (O_156,N_2861,N_2498);
or UO_157 (O_157,N_2588,N_2447);
xor UO_158 (O_158,N_2893,N_2561);
nand UO_159 (O_159,N_2431,N_2940);
nor UO_160 (O_160,N_2925,N_2474);
nor UO_161 (O_161,N_2325,N_2538);
nor UO_162 (O_162,N_2452,N_2656);
and UO_163 (O_163,N_2855,N_2678);
xor UO_164 (O_164,N_2817,N_2779);
nor UO_165 (O_165,N_2663,N_2649);
xor UO_166 (O_166,N_2787,N_2844);
nand UO_167 (O_167,N_2839,N_2350);
and UO_168 (O_168,N_2299,N_2752);
nor UO_169 (O_169,N_2653,N_2921);
or UO_170 (O_170,N_2920,N_2586);
nand UO_171 (O_171,N_2876,N_2883);
or UO_172 (O_172,N_2841,N_2801);
nand UO_173 (O_173,N_2758,N_2368);
nor UO_174 (O_174,N_2693,N_2413);
or UO_175 (O_175,N_2355,N_2389);
and UO_176 (O_176,N_2262,N_2688);
nor UO_177 (O_177,N_2533,N_2977);
nor UO_178 (O_178,N_2731,N_2289);
nand UO_179 (O_179,N_2365,N_2466);
nor UO_180 (O_180,N_2961,N_2567);
nor UO_181 (O_181,N_2509,N_2963);
nor UO_182 (O_182,N_2755,N_2495);
nand UO_183 (O_183,N_2959,N_2585);
nor UO_184 (O_184,N_2686,N_2997);
nor UO_185 (O_185,N_2898,N_2618);
nand UO_186 (O_186,N_2358,N_2345);
nor UO_187 (O_187,N_2534,N_2386);
nand UO_188 (O_188,N_2806,N_2971);
nor UO_189 (O_189,N_2478,N_2415);
nor UO_190 (O_190,N_2823,N_2712);
or UO_191 (O_191,N_2666,N_2497);
or UO_192 (O_192,N_2594,N_2850);
nand UO_193 (O_193,N_2810,N_2659);
nor UO_194 (O_194,N_2640,N_2668);
nor UO_195 (O_195,N_2673,N_2293);
and UO_196 (O_196,N_2396,N_2754);
and UO_197 (O_197,N_2741,N_2838);
or UO_198 (O_198,N_2804,N_2310);
or UO_199 (O_199,N_2259,N_2792);
nor UO_200 (O_200,N_2438,N_2664);
and UO_201 (O_201,N_2738,N_2800);
or UO_202 (O_202,N_2385,N_2512);
and UO_203 (O_203,N_2970,N_2597);
or UO_204 (O_204,N_2376,N_2909);
nor UO_205 (O_205,N_2485,N_2778);
nor UO_206 (O_206,N_2361,N_2674);
nand UO_207 (O_207,N_2601,N_2264);
nand UO_208 (O_208,N_2565,N_2336);
and UO_209 (O_209,N_2923,N_2769);
nand UO_210 (O_210,N_2685,N_2629);
and UO_211 (O_211,N_2765,N_2541);
or UO_212 (O_212,N_2571,N_2318);
or UO_213 (O_213,N_2710,N_2433);
nand UO_214 (O_214,N_2577,N_2737);
nand UO_215 (O_215,N_2877,N_2395);
nor UO_216 (O_216,N_2938,N_2273);
or UO_217 (O_217,N_2916,N_2894);
xor UO_218 (O_218,N_2947,N_2508);
nand UO_219 (O_219,N_2642,N_2428);
nor UO_220 (O_220,N_2798,N_2943);
and UO_221 (O_221,N_2422,N_2643);
nand UO_222 (O_222,N_2593,N_2655);
nand UO_223 (O_223,N_2767,N_2984);
and UO_224 (O_224,N_2539,N_2388);
or UO_225 (O_225,N_2313,N_2786);
and UO_226 (O_226,N_2540,N_2753);
nand UO_227 (O_227,N_2845,N_2697);
or UO_228 (O_228,N_2645,N_2733);
or UO_229 (O_229,N_2610,N_2856);
or UO_230 (O_230,N_2315,N_2631);
xor UO_231 (O_231,N_2298,N_2739);
or UO_232 (O_232,N_2274,N_2902);
xor UO_233 (O_233,N_2266,N_2955);
nor UO_234 (O_234,N_2824,N_2742);
or UO_235 (O_235,N_2436,N_2522);
or UO_236 (O_236,N_2910,N_2996);
nand UO_237 (O_237,N_2352,N_2626);
and UO_238 (O_238,N_2740,N_2915);
nand UO_239 (O_239,N_2330,N_2846);
or UO_240 (O_240,N_2563,N_2679);
and UO_241 (O_241,N_2449,N_2890);
or UO_242 (O_242,N_2727,N_2492);
nor UO_243 (O_243,N_2356,N_2709);
and UO_244 (O_244,N_2832,N_2865);
nand UO_245 (O_245,N_2680,N_2771);
or UO_246 (O_246,N_2621,N_2833);
and UO_247 (O_247,N_2936,N_2296);
or UO_248 (O_248,N_2444,N_2725);
nand UO_249 (O_249,N_2451,N_2481);
or UO_250 (O_250,N_2744,N_2728);
or UO_251 (O_251,N_2384,N_2604);
nand UO_252 (O_252,N_2848,N_2773);
nand UO_253 (O_253,N_2491,N_2579);
and UO_254 (O_254,N_2408,N_2342);
nor UO_255 (O_255,N_2434,N_2743);
or UO_256 (O_256,N_2632,N_2347);
or UO_257 (O_257,N_2918,N_2914);
nor UO_258 (O_258,N_2426,N_2402);
or UO_259 (O_259,N_2708,N_2566);
or UO_260 (O_260,N_2475,N_2827);
nand UO_261 (O_261,N_2511,N_2633);
and UO_262 (O_262,N_2990,N_2808);
and UO_263 (O_263,N_2267,N_2493);
nand UO_264 (O_264,N_2339,N_2929);
or UO_265 (O_265,N_2647,N_2587);
xnor UO_266 (O_266,N_2687,N_2805);
nand UO_267 (O_267,N_2860,N_2763);
xnor UO_268 (O_268,N_2882,N_2531);
nor UO_269 (O_269,N_2462,N_2843);
and UO_270 (O_270,N_2482,N_2400);
or UO_271 (O_271,N_2410,N_2300);
or UO_272 (O_272,N_2972,N_2340);
and UO_273 (O_273,N_2329,N_2570);
nor UO_274 (O_274,N_2750,N_2250);
or UO_275 (O_275,N_2406,N_2952);
nand UO_276 (O_276,N_2559,N_2255);
xnor UO_277 (O_277,N_2720,N_2553);
and UO_278 (O_278,N_2967,N_2314);
xor UO_279 (O_279,N_2622,N_2584);
nand UO_280 (O_280,N_2834,N_2628);
nor UO_281 (O_281,N_2945,N_2557);
nand UO_282 (O_282,N_2278,N_2973);
xor UO_283 (O_283,N_2589,N_2448);
or UO_284 (O_284,N_2957,N_2932);
nor UO_285 (O_285,N_2662,N_2471);
nand UO_286 (O_286,N_2922,N_2407);
nand UO_287 (O_287,N_2746,N_2672);
xor UO_288 (O_288,N_2875,N_2437);
nor UO_289 (O_289,N_2440,N_2582);
or UO_290 (O_290,N_2716,N_2349);
nor UO_291 (O_291,N_2427,N_2367);
xnor UO_292 (O_292,N_2849,N_2657);
nor UO_293 (O_293,N_2689,N_2683);
nor UO_294 (O_294,N_2294,N_2521);
nor UO_295 (O_295,N_2424,N_2467);
or UO_296 (O_296,N_2646,N_2359);
nand UO_297 (O_297,N_2321,N_2617);
or UO_298 (O_298,N_2667,N_2782);
nor UO_299 (O_299,N_2946,N_2513);
nor UO_300 (O_300,N_2517,N_2549);
nor UO_301 (O_301,N_2835,N_2729);
nand UO_302 (O_302,N_2420,N_2275);
or UO_303 (O_303,N_2435,N_2644);
nand UO_304 (O_304,N_2546,N_2613);
and UO_305 (O_305,N_2472,N_2569);
and UO_306 (O_306,N_2322,N_2425);
or UO_307 (O_307,N_2811,N_2862);
nand UO_308 (O_308,N_2455,N_2284);
and UO_309 (O_309,N_2429,N_2802);
nor UO_310 (O_310,N_2537,N_2919);
nor UO_311 (O_311,N_2854,N_2550);
xor UO_312 (O_312,N_2903,N_2985);
nor UO_313 (O_313,N_2813,N_2461);
nor UO_314 (O_314,N_2506,N_2578);
nor UO_315 (O_315,N_2392,N_2263);
nor UO_316 (O_316,N_2980,N_2519);
nor UO_317 (O_317,N_2993,N_2799);
and UO_318 (O_318,N_2701,N_2718);
nor UO_319 (O_319,N_2573,N_2869);
or UO_320 (O_320,N_2942,N_2484);
nand UO_321 (O_321,N_2344,N_2609);
and UO_322 (O_322,N_2826,N_2707);
nand UO_323 (O_323,N_2529,N_2353);
nand UO_324 (O_324,N_2831,N_2780);
or UO_325 (O_325,N_2812,N_2726);
nor UO_326 (O_326,N_2251,N_2784);
and UO_327 (O_327,N_2572,N_2292);
nand UO_328 (O_328,N_2976,N_2992);
or UO_329 (O_329,N_2283,N_2815);
or UO_330 (O_330,N_2265,N_2939);
nor UO_331 (O_331,N_2978,N_2543);
or UO_332 (O_332,N_2611,N_2790);
and UO_333 (O_333,N_2603,N_2317);
and UO_334 (O_334,N_2652,N_2840);
nand UO_335 (O_335,N_2705,N_2525);
or UO_336 (O_336,N_2483,N_2500);
nor UO_337 (O_337,N_2536,N_2456);
nor UO_338 (O_338,N_2735,N_2311);
or UO_339 (O_339,N_2418,N_2912);
or UO_340 (O_340,N_2560,N_2616);
or UO_341 (O_341,N_2372,N_2968);
or UO_342 (O_342,N_2518,N_2258);
nor UO_343 (O_343,N_2660,N_2441);
or UO_344 (O_344,N_2724,N_2286);
and UO_345 (O_345,N_2375,N_2641);
or UO_346 (O_346,N_2964,N_2348);
nor UO_347 (O_347,N_2953,N_2979);
nor UO_348 (O_348,N_2960,N_2558);
and UO_349 (O_349,N_2405,N_2304);
or UO_350 (O_350,N_2332,N_2870);
and UO_351 (O_351,N_2991,N_2544);
or UO_352 (O_352,N_2965,N_2981);
nor UO_353 (O_353,N_2277,N_2272);
nand UO_354 (O_354,N_2271,N_2620);
nor UO_355 (O_355,N_2499,N_2905);
or UO_356 (O_356,N_2906,N_2888);
nor UO_357 (O_357,N_2366,N_2892);
nor UO_358 (O_358,N_2948,N_2281);
nand UO_359 (O_359,N_2681,N_2374);
nor UO_360 (O_360,N_2703,N_2592);
nor UO_361 (O_361,N_2290,N_2605);
nand UO_362 (O_362,N_2904,N_2377);
or UO_363 (O_363,N_2337,N_2868);
nor UO_364 (O_364,N_2690,N_2409);
and UO_365 (O_365,N_2809,N_2761);
and UO_366 (O_366,N_2470,N_2896);
or UO_367 (O_367,N_2900,N_2568);
and UO_368 (O_368,N_2698,N_2378);
nor UO_369 (O_369,N_2524,N_2635);
and UO_370 (O_370,N_2822,N_2362);
or UO_371 (O_371,N_2776,N_2453);
or UO_372 (O_372,N_2285,N_2987);
nor UO_373 (O_373,N_2599,N_2403);
nand UO_374 (O_374,N_2287,N_2878);
or UO_375 (O_375,N_2360,N_2282);
or UO_376 (O_376,N_2315,N_2953);
and UO_377 (O_377,N_2853,N_2803);
and UO_378 (O_378,N_2552,N_2496);
and UO_379 (O_379,N_2700,N_2358);
and UO_380 (O_380,N_2811,N_2928);
nor UO_381 (O_381,N_2621,N_2624);
nor UO_382 (O_382,N_2536,N_2459);
or UO_383 (O_383,N_2428,N_2407);
and UO_384 (O_384,N_2865,N_2333);
and UO_385 (O_385,N_2416,N_2292);
and UO_386 (O_386,N_2539,N_2688);
or UO_387 (O_387,N_2703,N_2490);
or UO_388 (O_388,N_2320,N_2842);
or UO_389 (O_389,N_2448,N_2744);
and UO_390 (O_390,N_2525,N_2612);
and UO_391 (O_391,N_2320,N_2321);
nand UO_392 (O_392,N_2674,N_2979);
nand UO_393 (O_393,N_2482,N_2734);
or UO_394 (O_394,N_2781,N_2341);
or UO_395 (O_395,N_2881,N_2838);
nor UO_396 (O_396,N_2690,N_2256);
or UO_397 (O_397,N_2966,N_2490);
nor UO_398 (O_398,N_2781,N_2775);
nor UO_399 (O_399,N_2895,N_2897);
and UO_400 (O_400,N_2253,N_2905);
nand UO_401 (O_401,N_2267,N_2950);
nand UO_402 (O_402,N_2629,N_2903);
or UO_403 (O_403,N_2552,N_2289);
and UO_404 (O_404,N_2402,N_2258);
or UO_405 (O_405,N_2346,N_2919);
nand UO_406 (O_406,N_2827,N_2492);
nand UO_407 (O_407,N_2751,N_2695);
nor UO_408 (O_408,N_2947,N_2398);
nor UO_409 (O_409,N_2771,N_2890);
or UO_410 (O_410,N_2535,N_2291);
nand UO_411 (O_411,N_2547,N_2383);
nand UO_412 (O_412,N_2582,N_2345);
nand UO_413 (O_413,N_2406,N_2495);
nand UO_414 (O_414,N_2780,N_2664);
or UO_415 (O_415,N_2617,N_2950);
nor UO_416 (O_416,N_2556,N_2262);
nand UO_417 (O_417,N_2785,N_2778);
and UO_418 (O_418,N_2753,N_2745);
nand UO_419 (O_419,N_2455,N_2722);
nor UO_420 (O_420,N_2459,N_2812);
nor UO_421 (O_421,N_2812,N_2251);
or UO_422 (O_422,N_2665,N_2327);
and UO_423 (O_423,N_2570,N_2747);
xor UO_424 (O_424,N_2458,N_2796);
or UO_425 (O_425,N_2415,N_2434);
and UO_426 (O_426,N_2394,N_2768);
and UO_427 (O_427,N_2492,N_2696);
and UO_428 (O_428,N_2990,N_2673);
nand UO_429 (O_429,N_2339,N_2789);
and UO_430 (O_430,N_2818,N_2646);
nor UO_431 (O_431,N_2874,N_2725);
nand UO_432 (O_432,N_2858,N_2423);
and UO_433 (O_433,N_2285,N_2551);
and UO_434 (O_434,N_2582,N_2846);
nor UO_435 (O_435,N_2408,N_2640);
nand UO_436 (O_436,N_2632,N_2927);
nand UO_437 (O_437,N_2261,N_2670);
or UO_438 (O_438,N_2462,N_2621);
nand UO_439 (O_439,N_2278,N_2402);
or UO_440 (O_440,N_2555,N_2311);
or UO_441 (O_441,N_2838,N_2267);
nand UO_442 (O_442,N_2835,N_2931);
nor UO_443 (O_443,N_2568,N_2646);
xnor UO_444 (O_444,N_2691,N_2367);
or UO_445 (O_445,N_2485,N_2512);
or UO_446 (O_446,N_2652,N_2417);
nand UO_447 (O_447,N_2743,N_2531);
and UO_448 (O_448,N_2653,N_2609);
and UO_449 (O_449,N_2550,N_2418);
nor UO_450 (O_450,N_2964,N_2691);
xor UO_451 (O_451,N_2690,N_2533);
nor UO_452 (O_452,N_2280,N_2557);
or UO_453 (O_453,N_2917,N_2596);
or UO_454 (O_454,N_2781,N_2360);
nor UO_455 (O_455,N_2359,N_2540);
or UO_456 (O_456,N_2468,N_2676);
nand UO_457 (O_457,N_2345,N_2442);
or UO_458 (O_458,N_2804,N_2843);
nor UO_459 (O_459,N_2548,N_2564);
nor UO_460 (O_460,N_2549,N_2952);
nand UO_461 (O_461,N_2614,N_2927);
and UO_462 (O_462,N_2895,N_2558);
nor UO_463 (O_463,N_2855,N_2277);
or UO_464 (O_464,N_2707,N_2579);
and UO_465 (O_465,N_2553,N_2816);
nand UO_466 (O_466,N_2555,N_2719);
nand UO_467 (O_467,N_2458,N_2669);
and UO_468 (O_468,N_2389,N_2957);
or UO_469 (O_469,N_2848,N_2492);
and UO_470 (O_470,N_2849,N_2786);
nor UO_471 (O_471,N_2633,N_2808);
nor UO_472 (O_472,N_2952,N_2648);
and UO_473 (O_473,N_2891,N_2518);
nor UO_474 (O_474,N_2672,N_2550);
and UO_475 (O_475,N_2590,N_2612);
nand UO_476 (O_476,N_2824,N_2738);
nor UO_477 (O_477,N_2350,N_2939);
or UO_478 (O_478,N_2889,N_2500);
nor UO_479 (O_479,N_2800,N_2870);
or UO_480 (O_480,N_2474,N_2686);
nand UO_481 (O_481,N_2683,N_2909);
and UO_482 (O_482,N_2815,N_2309);
nand UO_483 (O_483,N_2938,N_2351);
nor UO_484 (O_484,N_2504,N_2302);
nand UO_485 (O_485,N_2930,N_2825);
nor UO_486 (O_486,N_2413,N_2763);
nor UO_487 (O_487,N_2928,N_2929);
nor UO_488 (O_488,N_2394,N_2541);
or UO_489 (O_489,N_2332,N_2921);
nor UO_490 (O_490,N_2353,N_2562);
or UO_491 (O_491,N_2888,N_2743);
or UO_492 (O_492,N_2372,N_2526);
nand UO_493 (O_493,N_2812,N_2892);
nand UO_494 (O_494,N_2481,N_2869);
and UO_495 (O_495,N_2606,N_2798);
or UO_496 (O_496,N_2787,N_2678);
or UO_497 (O_497,N_2955,N_2793);
nor UO_498 (O_498,N_2315,N_2622);
nor UO_499 (O_499,N_2739,N_2865);
endmodule