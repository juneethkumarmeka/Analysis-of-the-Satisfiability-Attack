module basic_2500_25000_3000_125_levels_10xor_5(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999;
xnor U0 (N_0,In_1474,In_1727);
nor U1 (N_1,In_315,In_356);
nor U2 (N_2,In_2414,In_1725);
and U3 (N_3,In_2478,In_502);
and U4 (N_4,In_2076,In_231);
nand U5 (N_5,In_266,In_2436);
nor U6 (N_6,In_2061,In_1091);
nor U7 (N_7,In_1112,In_631);
or U8 (N_8,In_1813,In_1612);
nand U9 (N_9,In_139,In_1211);
or U10 (N_10,In_747,In_437);
or U11 (N_11,In_1618,In_1691);
or U12 (N_12,In_2130,In_2286);
nand U13 (N_13,In_1939,In_2060);
or U14 (N_14,In_2128,In_304);
and U15 (N_15,In_1759,In_1399);
or U16 (N_16,In_124,In_1374);
xor U17 (N_17,In_1600,In_1808);
nand U18 (N_18,In_1907,In_1592);
nand U19 (N_19,In_721,In_1057);
nand U20 (N_20,In_136,In_19);
xor U21 (N_21,In_900,In_1381);
nand U22 (N_22,In_1336,In_1339);
and U23 (N_23,In_1284,In_681);
or U24 (N_24,In_1240,In_451);
and U25 (N_25,In_1582,In_1253);
or U26 (N_26,In_52,In_757);
xnor U27 (N_27,In_41,In_1209);
or U28 (N_28,In_628,In_2476);
and U29 (N_29,In_250,In_2418);
xnor U30 (N_30,In_32,In_137);
xnor U31 (N_31,In_1213,In_521);
nand U32 (N_32,In_1945,In_256);
nand U33 (N_33,In_1715,In_2247);
xor U34 (N_34,In_1333,In_564);
nor U35 (N_35,In_813,In_2001);
or U36 (N_36,In_160,In_2178);
nand U37 (N_37,In_131,In_964);
xnor U38 (N_38,In_1683,In_1781);
xor U39 (N_39,In_2298,In_2135);
xor U40 (N_40,In_1466,In_7);
nor U41 (N_41,In_666,In_1826);
nand U42 (N_42,In_1358,In_1203);
or U43 (N_43,In_606,In_3);
nor U44 (N_44,In_826,In_1351);
or U45 (N_45,In_770,In_1706);
or U46 (N_46,In_180,In_656);
or U47 (N_47,In_904,In_726);
and U48 (N_48,In_950,In_1180);
nand U49 (N_49,In_591,In_611);
nor U50 (N_50,In_942,In_2116);
nor U51 (N_51,In_2392,In_486);
nand U52 (N_52,In_2275,In_1773);
and U53 (N_53,In_1941,In_252);
xnor U54 (N_54,In_1723,In_2139);
xnor U55 (N_55,In_1491,In_203);
nor U56 (N_56,In_1184,In_1287);
xnor U57 (N_57,In_556,In_2292);
nand U58 (N_58,In_712,In_1508);
nand U59 (N_59,In_1806,In_1538);
or U60 (N_60,In_76,In_313);
or U61 (N_61,In_210,In_1911);
nor U62 (N_62,In_2325,In_1972);
nor U63 (N_63,In_2170,In_1406);
nor U64 (N_64,In_2228,In_1850);
nor U65 (N_65,In_2387,In_610);
nor U66 (N_66,In_943,In_2106);
nor U67 (N_67,In_1217,In_1768);
and U68 (N_68,In_1293,In_1797);
and U69 (N_69,In_218,In_201);
nand U70 (N_70,In_2221,In_1674);
xor U71 (N_71,In_346,In_993);
xor U72 (N_72,In_906,In_1751);
and U73 (N_73,In_2199,In_1188);
and U74 (N_74,In_331,In_1126);
xnor U75 (N_75,In_838,In_1429);
and U76 (N_76,In_1397,In_1272);
nand U77 (N_77,In_293,In_154);
nand U78 (N_78,In_1274,In_1068);
nand U79 (N_79,In_2421,In_1521);
xor U80 (N_80,In_1560,In_907);
or U81 (N_81,In_848,In_796);
and U82 (N_82,In_746,In_1730);
nand U83 (N_83,In_802,In_1670);
and U84 (N_84,In_1690,In_2451);
nand U85 (N_85,In_507,In_1714);
or U86 (N_86,In_1372,In_2242);
nand U87 (N_87,In_367,In_1953);
xnor U88 (N_88,In_1915,In_596);
nor U89 (N_89,In_415,In_1377);
nor U90 (N_90,In_2013,In_1835);
xnor U91 (N_91,In_138,In_1006);
and U92 (N_92,In_2112,In_402);
nor U93 (N_93,In_2157,In_2321);
nor U94 (N_94,In_2181,In_2142);
nor U95 (N_95,In_337,In_523);
nand U96 (N_96,In_800,In_2459);
nor U97 (N_97,In_2066,In_448);
or U98 (N_98,In_2023,In_1138);
nand U99 (N_99,In_0,In_2439);
and U100 (N_100,In_417,In_347);
or U101 (N_101,In_2318,In_961);
or U102 (N_102,In_963,In_2186);
xnor U103 (N_103,In_2235,In_1022);
nor U104 (N_104,In_1663,In_209);
nand U105 (N_105,In_2332,In_1079);
or U106 (N_106,In_2261,In_249);
and U107 (N_107,In_1617,In_436);
and U108 (N_108,In_2154,In_111);
nor U109 (N_109,In_1038,In_1917);
xnor U110 (N_110,In_767,In_1831);
nand U111 (N_111,In_429,In_570);
or U112 (N_112,In_1924,In_559);
and U113 (N_113,In_1139,In_877);
xor U114 (N_114,In_853,In_50);
or U115 (N_115,In_1008,In_1601);
and U116 (N_116,In_2417,In_349);
nand U117 (N_117,In_1128,In_483);
nor U118 (N_118,In_2053,In_2007);
xnor U119 (N_119,In_953,In_60);
or U120 (N_120,In_1441,In_385);
nor U121 (N_121,In_919,In_322);
or U122 (N_122,In_2482,In_1665);
nand U123 (N_123,In_1687,In_1605);
and U124 (N_124,In_1798,In_1771);
or U125 (N_125,In_671,In_1647);
xnor U126 (N_126,In_2397,In_395);
xor U127 (N_127,In_1480,In_1559);
nand U128 (N_128,In_787,In_2264);
nand U129 (N_129,In_1923,In_194);
or U130 (N_130,In_2236,In_1111);
and U131 (N_131,In_16,In_1959);
nand U132 (N_132,In_47,In_1445);
xnor U133 (N_133,In_1968,In_1346);
xor U134 (N_134,In_2303,In_2357);
or U135 (N_135,In_695,In_1856);
or U136 (N_136,In_2343,In_994);
nand U137 (N_137,In_2259,In_912);
xor U138 (N_138,In_1942,In_790);
nor U139 (N_139,In_2164,In_985);
xor U140 (N_140,In_2168,In_949);
or U141 (N_141,In_920,In_394);
or U142 (N_142,In_884,In_75);
nand U143 (N_143,In_1570,In_1402);
or U144 (N_144,In_1844,In_2079);
or U145 (N_145,In_2209,In_2370);
or U146 (N_146,In_679,In_1711);
and U147 (N_147,In_1440,In_1081);
xor U148 (N_148,In_1634,In_286);
xor U149 (N_149,In_399,In_1210);
and U150 (N_150,In_1583,In_2102);
nor U151 (N_151,In_1815,In_1145);
xor U152 (N_152,In_982,In_1282);
or U153 (N_153,In_1565,In_1593);
xnor U154 (N_154,In_20,In_2045);
nor U155 (N_155,In_2255,In_2391);
or U156 (N_156,In_1925,In_88);
xnor U157 (N_157,In_2279,In_1719);
xor U158 (N_158,In_255,In_2485);
nor U159 (N_159,In_2337,In_2454);
nand U160 (N_160,In_680,In_2394);
nand U161 (N_161,In_1499,In_73);
xnor U162 (N_162,In_2441,In_1178);
nor U163 (N_163,In_2489,In_670);
xor U164 (N_164,In_246,In_1251);
xor U165 (N_165,In_21,In_2311);
or U166 (N_166,In_2069,In_2359);
or U167 (N_167,In_96,In_717);
or U168 (N_168,In_1303,In_2408);
xnor U169 (N_169,In_2034,In_588);
xor U170 (N_170,In_2093,In_2237);
and U171 (N_171,In_2447,In_1910);
xnor U172 (N_172,In_745,In_240);
nor U173 (N_173,In_2249,In_1395);
or U174 (N_174,In_2345,In_1443);
or U175 (N_175,In_1047,In_2257);
nor U176 (N_176,In_2351,In_1107);
nand U177 (N_177,In_234,In_1158);
or U178 (N_178,In_1183,In_2368);
or U179 (N_179,In_1795,In_511);
xnor U180 (N_180,In_922,In_959);
xnor U181 (N_181,In_1973,In_513);
and U182 (N_182,In_897,In_1660);
nand U183 (N_183,In_2118,In_157);
xnor U184 (N_184,In_1157,In_93);
and U185 (N_185,In_896,In_2223);
nor U186 (N_186,In_1985,In_1548);
and U187 (N_187,In_785,In_1710);
nand U188 (N_188,In_2248,In_1541);
or U189 (N_189,In_1896,In_881);
nor U190 (N_190,In_782,In_445);
xnor U191 (N_191,In_1919,In_1444);
xor U192 (N_192,In_2269,In_1292);
or U193 (N_193,In_1321,In_1140);
and U194 (N_194,In_176,In_363);
xnor U195 (N_195,In_918,In_1290);
or U196 (N_196,In_1702,In_334);
nand U197 (N_197,In_369,In_2348);
nand U198 (N_198,In_621,In_879);
nor U199 (N_199,In_509,In_1682);
and U200 (N_200,In_927,In_274);
xor U201 (N_201,N_10,In_1307);
nand U202 (N_202,In_663,In_1054);
or U203 (N_203,In_1023,In_1356);
nand U204 (N_204,In_1921,In_2117);
nor U205 (N_205,In_1638,In_593);
and U206 (N_206,N_125,In_771);
nand U207 (N_207,In_2159,In_1026);
and U208 (N_208,In_365,In_227);
xor U209 (N_209,In_1881,In_1712);
xor U210 (N_210,In_163,In_2466);
and U211 (N_211,In_673,In_1273);
nand U212 (N_212,N_144,In_885);
xnor U213 (N_213,In_1216,In_452);
or U214 (N_214,N_52,In_1046);
or U215 (N_215,In_1342,In_2109);
xnor U216 (N_216,In_2002,In_263);
xnor U217 (N_217,In_1802,In_338);
and U218 (N_218,In_1847,In_1500);
nand U219 (N_219,In_2008,In_2029);
nand U220 (N_220,In_192,In_2031);
xnor U221 (N_221,In_1744,In_2406);
xnor U222 (N_222,In_147,In_426);
nand U223 (N_223,In_1490,In_605);
nand U224 (N_224,N_163,In_1049);
and U225 (N_225,N_26,In_2495);
nand U226 (N_226,In_2474,In_1837);
or U227 (N_227,In_2342,In_2425);
xnor U228 (N_228,In_1830,In_1951);
nor U229 (N_229,In_1679,In_1520);
xnor U230 (N_230,In_2155,In_2470);
xnor U231 (N_231,In_2040,In_895);
nor U232 (N_232,In_2340,In_951);
nor U233 (N_233,N_166,In_2483);
nor U234 (N_234,In_1427,In_1119);
nor U235 (N_235,In_1264,In_1448);
or U236 (N_236,In_2490,In_102);
and U237 (N_237,In_668,In_744);
nor U238 (N_238,In_67,N_78);
nand U239 (N_239,In_734,In_1645);
or U240 (N_240,In_2475,In_1353);
nor U241 (N_241,In_1522,In_1453);
or U242 (N_242,In_2400,In_845);
or U243 (N_243,In_11,In_1922);
and U244 (N_244,In_1603,N_23);
and U245 (N_245,In_36,In_2143);
or U246 (N_246,In_1129,In_2028);
and U247 (N_247,In_298,In_1966);
nand U248 (N_248,In_2334,In_2022);
or U249 (N_249,N_152,In_554);
nand U250 (N_250,In_1432,In_2301);
xor U251 (N_251,In_1431,In_2115);
xor U252 (N_252,In_759,In_2014);
nand U253 (N_253,N_96,In_793);
or U254 (N_254,In_847,In_905);
nor U255 (N_255,In_1909,In_279);
and U256 (N_256,N_72,In_1132);
xor U257 (N_257,In_2051,In_760);
nor U258 (N_258,In_470,In_1355);
xnor U259 (N_259,In_1099,In_490);
xor U260 (N_260,In_1969,In_329);
nand U261 (N_261,In_756,N_60);
xnor U262 (N_262,In_1027,In_1528);
xnor U263 (N_263,N_8,In_2449);
or U264 (N_264,In_1976,In_2090);
or U265 (N_265,In_2455,In_1050);
and U266 (N_266,In_211,In_105);
or U267 (N_267,In_938,In_2444);
and U268 (N_268,In_319,N_82);
and U269 (N_269,In_23,In_1975);
xor U270 (N_270,In_2179,In_1747);
xnor U271 (N_271,In_77,In_1015);
nor U272 (N_272,In_1297,In_174);
or U273 (N_273,In_1950,In_604);
xor U274 (N_274,In_2026,In_1329);
xor U275 (N_275,In_224,In_1532);
nor U276 (N_276,In_1698,In_383);
nand U277 (N_277,In_1820,In_772);
nor U278 (N_278,In_183,In_1863);
xnor U279 (N_279,In_601,In_2212);
and U280 (N_280,In_292,In_1804);
nand U281 (N_281,In_1694,In_1062);
nor U282 (N_282,In_54,In_1940);
nor U283 (N_283,In_883,In_1437);
and U284 (N_284,In_1542,In_1035);
nor U285 (N_285,In_1625,In_856);
nand U286 (N_286,In_247,In_615);
xor U287 (N_287,In_946,In_1263);
nor U288 (N_288,In_1741,In_1231);
nand U289 (N_289,In_1078,In_2070);
and U290 (N_290,In_1799,In_35);
xnor U291 (N_291,N_22,In_328);
nor U292 (N_292,In_2147,In_187);
nand U293 (N_293,N_0,N_93);
nor U294 (N_294,In_1567,In_1754);
and U295 (N_295,In_361,In_576);
nor U296 (N_296,In_518,In_1833);
xor U297 (N_297,In_818,In_12);
nand U298 (N_298,In_1061,In_562);
nor U299 (N_299,In_1640,In_1283);
and U300 (N_300,In_241,In_1470);
nand U301 (N_301,In_2138,N_120);
or U302 (N_302,In_2125,In_318);
and U303 (N_303,In_1760,In_2);
or U304 (N_304,In_2442,In_1085);
or U305 (N_305,In_1314,In_1979);
nand U306 (N_306,In_797,In_1722);
xor U307 (N_307,In_290,In_1644);
xor U308 (N_308,In_133,In_1639);
nand U309 (N_309,In_1967,In_368);
or U310 (N_310,In_527,N_79);
xor U311 (N_311,In_2196,In_435);
nor U312 (N_312,In_1829,In_1530);
xor U313 (N_313,N_195,In_265);
nor U314 (N_314,In_1549,In_2216);
and U315 (N_315,In_1875,In_2016);
xnor U316 (N_316,In_499,In_1097);
nor U317 (N_317,In_1502,In_17);
and U318 (N_318,In_1763,N_141);
nor U319 (N_319,N_86,In_1792);
nand U320 (N_320,In_997,In_1574);
nor U321 (N_321,In_2222,In_1596);
and U322 (N_322,In_1877,In_1527);
or U323 (N_323,In_1529,In_1637);
xnor U324 (N_324,In_707,In_652);
and U325 (N_325,In_2113,In_1864);
nor U326 (N_326,In_2263,In_2011);
and U327 (N_327,In_1137,In_2119);
and U328 (N_328,In_1458,In_1425);
xnor U329 (N_329,In_852,In_1174);
and U330 (N_330,In_1566,In_398);
xor U331 (N_331,In_1254,N_185);
nand U332 (N_332,In_1124,In_2339);
and U333 (N_333,In_937,In_986);
nor U334 (N_334,In_816,In_1029);
nor U335 (N_335,In_2480,N_165);
xnor U336 (N_336,In_1746,N_131);
and U337 (N_337,In_1540,In_1030);
nand U338 (N_338,In_1226,In_1718);
or U339 (N_339,In_1367,In_832);
nor U340 (N_340,In_1676,In_291);
or U341 (N_341,In_1489,In_1051);
nor U342 (N_342,In_1033,In_25);
and U343 (N_343,In_711,In_1201);
nand U344 (N_344,In_376,In_1753);
nand U345 (N_345,N_128,In_1487);
and U346 (N_346,In_968,In_1895);
or U347 (N_347,In_104,In_1389);
nand U348 (N_348,In_2052,In_2206);
nand U349 (N_349,In_2362,In_970);
nand U350 (N_350,In_214,In_1486);
or U351 (N_351,In_645,In_236);
xnor U352 (N_352,In_870,In_980);
or U353 (N_353,In_1633,N_19);
xor U354 (N_354,In_1769,In_1621);
xor U355 (N_355,In_789,In_2322);
xor U356 (N_356,In_228,In_2457);
nand U357 (N_357,In_696,In_1767);
nand U358 (N_358,In_568,In_1931);
nand U359 (N_359,In_1277,In_321);
or U360 (N_360,In_1562,In_1385);
nor U361 (N_361,In_332,In_823);
or U362 (N_362,In_1849,In_1082);
nand U363 (N_363,In_370,In_1070);
nand U364 (N_364,In_343,In_1707);
nand U365 (N_365,In_863,In_2333);
and U366 (N_366,In_2413,In_988);
nand U367 (N_367,In_1693,In_729);
xor U368 (N_368,In_1544,In_1832);
xnor U369 (N_369,N_140,In_1879);
or U370 (N_370,In_1661,In_411);
nand U371 (N_371,In_1523,In_2190);
xnor U372 (N_372,N_127,In_2161);
xor U373 (N_373,In_1181,In_533);
nand U374 (N_374,In_1165,In_1456);
and U375 (N_375,In_1577,In_1058);
xor U376 (N_376,In_1949,In_1426);
or U377 (N_377,In_86,N_80);
and U378 (N_378,In_1249,In_2358);
and U379 (N_379,In_2405,In_525);
nand U380 (N_380,In_553,N_137);
xnor U381 (N_381,N_99,In_788);
or U382 (N_382,In_532,In_2175);
nor U383 (N_383,In_1175,In_973);
xor U384 (N_384,In_1142,In_1301);
xor U385 (N_385,In_1599,In_2122);
nand U386 (N_386,In_804,In_1214);
and U387 (N_387,In_355,In_106);
nor U388 (N_388,In_799,In_1258);
nor U389 (N_389,In_779,In_775);
xnor U390 (N_390,In_1450,In_1393);
nand U391 (N_391,In_545,In_2456);
xor U392 (N_392,In_1766,In_2384);
nand U393 (N_393,In_1415,In_1218);
or U394 (N_394,In_2153,N_3);
nand U395 (N_395,In_1853,N_122);
and U396 (N_396,In_1464,In_1224);
and U397 (N_397,In_1237,In_1227);
nor U398 (N_398,In_1598,In_421);
nand U399 (N_399,In_408,In_1092);
xor U400 (N_400,In_2166,In_1626);
nand U401 (N_401,N_118,In_1517);
nor U402 (N_402,In_1961,N_313);
xnor U403 (N_403,N_107,In_504);
or U404 (N_404,In_222,In_1629);
nor U405 (N_405,In_430,In_1247);
nor U406 (N_406,In_1186,N_150);
and U407 (N_407,In_1733,In_1518);
and U408 (N_408,In_371,N_30);
xor U409 (N_409,In_535,In_755);
nand U410 (N_410,In_95,In_1536);
nor U411 (N_411,N_130,In_2018);
nand U412 (N_412,In_217,In_646);
xnor U413 (N_413,In_330,In_1052);
nand U414 (N_414,In_1684,In_1898);
and U415 (N_415,In_1721,In_262);
and U416 (N_416,In_915,N_397);
nor U417 (N_417,In_1238,In_1403);
nand U418 (N_418,N_365,N_191);
nand U419 (N_419,In_39,N_270);
xnor U420 (N_420,In_1361,In_326);
or U421 (N_421,In_1295,In_2080);
xor U422 (N_422,In_1411,In_1048);
xnor U423 (N_423,In_1955,In_1862);
or U424 (N_424,In_864,In_763);
nand U425 (N_425,In_134,In_66);
or U426 (N_426,N_184,N_155);
nand U427 (N_427,In_205,In_2274);
and U428 (N_428,In_1954,In_508);
xor U429 (N_429,N_291,In_1981);
and U430 (N_430,N_145,In_1809);
or U431 (N_431,In_297,N_243);
xnor U432 (N_432,In_2423,N_132);
and U433 (N_433,N_360,In_1435);
and U434 (N_434,In_1348,N_4);
xor U435 (N_435,In_38,In_202);
nor U436 (N_436,In_2374,In_738);
and U437 (N_437,In_2316,In_476);
or U438 (N_438,N_157,N_362);
xnor U439 (N_439,In_2369,In_2124);
or U440 (N_440,In_1885,In_1419);
or U441 (N_441,In_819,In_2232);
or U442 (N_442,In_15,In_353);
xnor U443 (N_443,In_392,In_454);
nor U444 (N_444,In_2420,In_758);
nand U445 (N_445,In_1482,In_626);
or U446 (N_446,In_888,In_1874);
or U447 (N_447,In_1903,In_1202);
nand U448 (N_448,In_406,N_194);
nor U449 (N_449,N_357,In_2491);
xnor U450 (N_450,N_326,In_13);
nand U451 (N_451,In_2044,In_2317);
and U452 (N_452,In_1839,N_398);
or U453 (N_453,In_653,In_1784);
and U454 (N_454,In_1288,In_1865);
nand U455 (N_455,N_9,In_208);
nor U456 (N_456,N_54,In_1515);
nand U457 (N_457,In_1196,In_1788);
nand U458 (N_458,In_339,In_1986);
and U459 (N_459,In_2193,In_2471);
nand U460 (N_460,In_2030,In_2382);
and U461 (N_461,N_188,In_698);
xnor U462 (N_462,In_273,In_892);
nand U463 (N_463,In_558,In_2313);
and U464 (N_464,In_158,In_2272);
nand U465 (N_465,In_1452,In_2084);
nor U466 (N_466,In_1519,In_1589);
xnor U467 (N_467,In_1571,In_849);
or U468 (N_468,In_407,In_418);
or U469 (N_469,N_304,N_231);
and U470 (N_470,In_2050,In_2068);
nand U471 (N_471,In_1726,In_155);
nor U472 (N_472,In_635,In_914);
xor U473 (N_473,N_229,N_129);
nor U474 (N_474,In_1101,N_248);
or U475 (N_475,In_836,N_167);
xnor U476 (N_476,In_1042,In_1308);
or U477 (N_477,In_268,In_2411);
nor U478 (N_478,In_1278,In_1055);
xor U479 (N_479,N_87,In_2156);
xnor U480 (N_480,In_115,In_2494);
nor U481 (N_481,In_1117,In_846);
and U482 (N_482,In_842,In_941);
xnor U483 (N_483,In_2498,In_612);
nor U484 (N_484,In_1675,In_1155);
nand U485 (N_485,N_264,In_740);
nand U486 (N_486,In_1736,In_1999);
and U487 (N_487,In_2280,In_762);
nor U488 (N_488,In_251,In_1842);
and U489 (N_489,In_2054,In_2453);
and U490 (N_490,In_517,In_575);
nand U491 (N_491,In_1659,In_1151);
nor U492 (N_492,N_102,In_422);
or U493 (N_493,N_81,In_702);
nor U494 (N_494,In_372,N_368);
nand U495 (N_495,In_764,In_1786);
nand U496 (N_496,In_619,In_664);
and U497 (N_497,N_90,In_380);
nor U498 (N_498,In_1328,N_17);
nor U499 (N_499,In_2167,In_1539);
and U500 (N_500,In_592,In_1872);
nor U501 (N_501,In_149,In_1121);
nor U502 (N_502,In_1018,In_156);
or U503 (N_503,In_449,In_622);
and U504 (N_504,In_1906,In_1729);
nor U505 (N_505,N_88,In_1807);
or U506 (N_506,N_213,In_705);
nor U507 (N_507,N_180,N_356);
xnor U508 (N_508,N_48,In_1897);
or U509 (N_509,In_1156,In_2047);
and U510 (N_510,In_2398,In_2430);
xnor U511 (N_511,In_839,In_1056);
nand U512 (N_512,In_1244,In_627);
or U513 (N_513,In_1918,In_1028);
or U514 (N_514,In_948,In_2203);
xnor U515 (N_515,In_542,In_305);
nor U516 (N_516,In_1322,In_1988);
and U517 (N_517,In_703,In_485);
xor U518 (N_518,In_1010,In_2043);
and U519 (N_519,In_1089,In_1654);
nand U520 (N_520,N_322,In_2158);
and U521 (N_521,In_381,In_783);
or U522 (N_522,In_2165,In_1742);
xnor U523 (N_523,N_105,N_171);
or U524 (N_524,In_1267,In_373);
and U525 (N_525,In_1823,In_1428);
nand U526 (N_526,In_665,In_2208);
xor U527 (N_527,In_2049,In_204);
nor U528 (N_528,In_2277,In_1024);
nand U529 (N_529,In_2265,In_1810);
xnor U530 (N_530,In_119,In_2169);
xor U531 (N_531,N_11,In_1279);
xor U532 (N_532,In_2136,In_2213);
and U533 (N_533,In_865,N_251);
or U534 (N_534,In_2407,In_901);
xor U535 (N_535,N_266,In_78);
nor U536 (N_536,In_1845,In_971);
xor U537 (N_537,In_1868,In_784);
nand U538 (N_538,N_366,In_1388);
or U539 (N_539,In_494,N_24);
nand U540 (N_540,In_488,N_15);
nand U541 (N_541,In_390,In_63);
xor U542 (N_542,In_1934,In_1483);
and U543 (N_543,In_1590,In_2250);
nor U544 (N_544,N_115,In_2452);
xor U545 (N_545,In_1164,In_803);
nand U546 (N_546,In_1734,In_538);
nor U547 (N_547,N_240,In_301);
and U548 (N_548,N_391,N_227);
nand U549 (N_549,In_714,In_2492);
or U550 (N_550,In_1261,In_1331);
nor U551 (N_551,In_2009,N_288);
and U552 (N_552,N_233,N_234);
and U553 (N_553,N_319,In_2107);
or U554 (N_554,In_972,In_1789);
xnor U555 (N_555,N_108,In_1012);
nand U556 (N_556,In_2058,In_843);
or U557 (N_557,In_226,In_2097);
and U558 (N_558,In_1136,In_1952);
nor U559 (N_559,In_1553,In_351);
and U560 (N_560,N_176,In_1717);
or U561 (N_561,N_1,In_1298);
nor U562 (N_562,In_1606,In_1704);
or U563 (N_563,In_2104,N_35);
and U564 (N_564,In_1350,In_1154);
or U565 (N_565,N_198,In_1451);
and U566 (N_566,In_26,In_560);
or U567 (N_567,N_18,In_2177);
and U568 (N_568,In_307,In_1257);
xor U569 (N_569,In_1275,N_222);
xnor U570 (N_570,In_567,In_830);
nor U571 (N_571,N_42,In_1318);
or U572 (N_572,N_104,In_410);
nand U573 (N_573,N_385,In_530);
and U574 (N_574,In_433,In_1668);
xnor U575 (N_575,In_1587,N_289);
xor U576 (N_576,In_2020,In_2484);
or U577 (N_577,In_243,N_200);
xnor U578 (N_578,In_196,In_1713);
nor U579 (N_579,In_1572,In_1509);
nand U580 (N_580,N_29,In_235);
or U581 (N_581,N_51,In_515);
nand U582 (N_582,In_1494,In_257);
xor U583 (N_583,In_289,N_241);
and U584 (N_584,In_812,In_314);
and U585 (N_585,In_2027,N_57);
and U586 (N_586,In_1580,In_59);
or U587 (N_587,In_1400,In_1410);
and U588 (N_588,In_2245,In_733);
and U589 (N_589,N_192,In_2271);
xnor U590 (N_590,In_1748,In_489);
nand U591 (N_591,In_171,In_1800);
xor U592 (N_592,In_2246,In_1569);
or U593 (N_593,In_43,In_2253);
nand U594 (N_594,In_206,In_1360);
and U595 (N_595,In_2039,In_440);
nor U596 (N_596,In_1964,In_145);
nand U597 (N_597,In_65,In_463);
xnor U598 (N_598,In_660,In_975);
xnor U599 (N_599,In_1041,In_24);
or U600 (N_600,N_148,In_419);
xor U601 (N_601,In_1764,In_1265);
nor U602 (N_602,N_445,In_2324);
and U603 (N_603,In_724,In_2017);
nand U604 (N_604,In_1855,In_1191);
or U605 (N_605,In_1471,N_294);
xnor U606 (N_606,In_678,In_1728);
nor U607 (N_607,In_1507,N_255);
and U608 (N_608,In_1680,In_389);
nor U609 (N_609,N_562,N_259);
nor U610 (N_610,In_2312,N_375);
xor U611 (N_611,In_2380,In_1524);
or U612 (N_612,In_1783,In_1148);
nand U613 (N_613,In_1206,In_352);
nor U614 (N_614,In_1311,N_134);
xnor U615 (N_615,N_414,In_1037);
nand U616 (N_616,In_658,In_2019);
nor U617 (N_617,In_2258,In_1894);
nor U618 (N_618,In_2290,In_944);
nor U619 (N_619,N_74,In_989);
nand U620 (N_620,N_204,In_72);
nand U621 (N_621,In_2461,In_2140);
xnor U622 (N_622,N_262,In_2195);
nand U623 (N_623,In_637,In_1414);
or U624 (N_624,In_2173,In_1005);
xnor U625 (N_625,In_835,In_2440);
nand U626 (N_626,In_1072,In_1468);
xor U627 (N_627,In_2428,In_1641);
or U628 (N_628,N_216,N_377);
or U629 (N_629,N_538,In_583);
nand U630 (N_630,N_351,N_50);
and U631 (N_631,N_592,In_801);
nor U632 (N_632,In_974,In_814);
and U633 (N_633,N_524,In_1014);
xnor U634 (N_634,In_1995,In_1873);
xor U635 (N_635,In_505,N_516);
or U636 (N_636,In_1344,In_903);
nand U637 (N_637,In_1609,In_1946);
xor U638 (N_638,In_976,In_837);
nand U639 (N_639,In_2487,In_1630);
and U640 (N_640,In_1756,In_561);
or U641 (N_641,In_715,In_1838);
nor U642 (N_642,In_270,N_593);
xor U643 (N_643,In_2238,In_580);
or U644 (N_644,In_1168,N_238);
or U645 (N_645,In_2294,In_388);
nor U646 (N_646,In_1525,In_732);
and U647 (N_647,N_196,In_594);
or U648 (N_648,N_542,N_553);
nor U649 (N_649,In_1673,N_226);
nand U650 (N_650,N_566,In_1208);
or U651 (N_651,In_2373,N_491);
and U652 (N_652,In_1110,N_275);
nand U653 (N_653,N_89,N_469);
nor U654 (N_654,In_569,In_2293);
xor U655 (N_655,N_559,In_1077);
and U656 (N_656,N_170,N_455);
and U657 (N_657,N_154,N_449);
and U658 (N_658,In_1255,N_6);
nor U659 (N_659,In_1045,In_169);
nand U660 (N_660,In_550,In_1578);
or U661 (N_661,In_2033,N_350);
nand U662 (N_662,N_290,In_170);
xnor U663 (N_663,In_142,In_995);
nor U664 (N_664,N_475,In_685);
or U665 (N_665,In_977,N_512);
xor U666 (N_666,In_624,N_550);
xnor U667 (N_667,In_341,In_1642);
or U668 (N_668,In_2363,In_1433);
xnor U669 (N_669,In_484,In_2225);
and U670 (N_670,In_1602,In_2220);
or U671 (N_671,N_197,In_132);
or U672 (N_672,N_435,N_483);
xnor U673 (N_673,In_184,In_1016);
or U674 (N_674,N_558,In_172);
nor U675 (N_675,In_1758,In_644);
nor U676 (N_676,In_2335,N_109);
xor U677 (N_677,In_2415,In_1819);
nand U678 (N_678,In_2388,N_556);
and U679 (N_679,In_48,In_2032);
and U680 (N_680,In_1021,N_55);
or U681 (N_681,In_323,In_1989);
and U682 (N_682,In_1098,In_2234);
and U683 (N_683,In_1493,In_1787);
and U684 (N_684,In_2133,In_473);
and U685 (N_685,N_425,In_1310);
nor U686 (N_686,N_405,N_273);
nand U687 (N_687,In_345,In_64);
nand U688 (N_688,In_116,In_1776);
or U689 (N_689,In_74,In_774);
xor U690 (N_690,In_1666,In_269);
nand U691 (N_691,In_891,N_358);
nor U692 (N_692,N_335,N_230);
xnor U693 (N_693,In_1854,In_272);
nand U694 (N_694,In_1262,In_2469);
nand U695 (N_695,In_978,N_576);
and U696 (N_696,N_525,In_1163);
and U697 (N_697,In_1004,In_1106);
nand U698 (N_698,N_68,N_56);
xnor U699 (N_699,In_2062,In_1484);
and U700 (N_700,N_493,In_806);
nand U701 (N_701,N_409,N_12);
nor U702 (N_702,In_2329,In_428);
nor U703 (N_703,N_561,N_484);
or U704 (N_704,In_1631,In_1382);
nor U705 (N_705,In_348,In_229);
and U706 (N_706,In_765,In_992);
xnor U707 (N_707,In_278,In_177);
nor U708 (N_708,In_2055,In_917);
and U709 (N_709,In_1551,In_1416);
nor U710 (N_710,In_2121,In_1268);
xnor U711 (N_711,N_330,In_2463);
nand U712 (N_712,In_1568,In_1908);
xor U713 (N_713,In_1770,In_1000);
and U714 (N_714,In_1324,N_462);
xnor U715 (N_715,In_654,In_2085);
nand U716 (N_716,In_79,In_1313);
nor U717 (N_717,In_2488,In_129);
or U718 (N_718,In_1459,In_1620);
or U719 (N_719,N_62,In_1497);
nand U720 (N_720,In_1648,In_1891);
nor U721 (N_721,In_821,In_2493);
nand U722 (N_722,In_1364,In_1912);
and U723 (N_723,In_150,In_2273);
or U724 (N_724,In_597,In_727);
or U725 (N_725,In_1173,In_1266);
nor U726 (N_726,N_473,N_393);
nand U727 (N_727,N_201,In_2078);
or U728 (N_728,In_1011,In_1291);
xnor U729 (N_729,In_1167,N_70);
nor U730 (N_730,In_1512,In_82);
nor U731 (N_731,In_1785,In_1761);
nand U732 (N_732,In_1740,N_44);
nand U733 (N_733,In_827,N_101);
nor U734 (N_734,N_597,In_1289);
or U735 (N_735,N_271,In_1780);
or U736 (N_736,N_479,In_2176);
nand U737 (N_737,N_214,In_659);
nor U738 (N_738,N_324,N_546);
xnor U739 (N_739,In_669,In_2497);
nand U740 (N_740,In_1103,In_1134);
and U741 (N_741,In_1757,In_1828);
xnor U742 (N_742,N_419,In_1749);
xnor U743 (N_743,In_565,N_489);
or U744 (N_744,In_1883,In_965);
nand U745 (N_745,In_1672,In_1737);
or U746 (N_746,N_232,N_486);
and U747 (N_747,In_798,In_1738);
nand U748 (N_748,In_598,In_851);
nor U749 (N_749,N_329,In_551);
or U750 (N_750,In_300,N_323);
or U751 (N_751,In_2065,In_960);
nor U752 (N_752,In_873,In_1232);
nand U753 (N_753,In_2473,In_113);
or U754 (N_754,In_1204,In_2087);
or U755 (N_755,In_1446,In_42);
xor U756 (N_756,In_1146,In_809);
and U757 (N_757,N_202,N_584);
xnor U758 (N_758,In_754,In_710);
and U759 (N_759,In_1455,In_572);
nor U760 (N_760,In_1469,In_1852);
xor U761 (N_761,In_1013,N_28);
nand U762 (N_762,In_1980,In_245);
nor U763 (N_763,In_795,In_1380);
nand U764 (N_764,N_342,In_1084);
and U765 (N_765,In_478,In_1299);
nand U766 (N_766,In_2450,In_589);
xor U767 (N_767,In_1043,In_1791);
xnor U768 (N_768,In_469,In_723);
nand U769 (N_769,In_2276,N_563);
nor U770 (N_770,In_1822,In_162);
nor U771 (N_771,In_1841,In_1615);
nor U772 (N_772,In_441,In_141);
or U773 (N_773,In_90,N_139);
nor U774 (N_774,N_153,N_249);
nand U775 (N_775,In_1409,N_211);
xor U776 (N_776,N_431,In_2288);
or U777 (N_777,In_1391,In_1113);
nor U778 (N_778,In_31,In_1065);
or U779 (N_779,In_471,N_210);
nor U780 (N_780,In_825,N_492);
nor U781 (N_781,In_344,In_2194);
and U782 (N_782,N_499,N_406);
and U783 (N_783,N_476,N_502);
nor U784 (N_784,N_540,In_1235);
or U785 (N_785,N_521,N_497);
or U786 (N_786,In_1447,In_2184);
xor U787 (N_787,In_700,N_207);
nand U788 (N_788,In_786,N_236);
nor U789 (N_789,In_850,In_446);
or U790 (N_790,N_311,N_307);
nand U791 (N_791,N_169,In_1504);
or U792 (N_792,In_2056,N_199);
xnor U793 (N_793,In_1182,In_306);
nor U794 (N_794,In_175,In_1044);
nor U795 (N_795,N_535,In_2174);
and U796 (N_796,N_61,N_364);
nand U797 (N_797,N_142,In_2499);
or U798 (N_798,In_2266,In_600);
or U799 (N_799,In_585,N_494);
and U800 (N_800,N_749,In_1554);
xor U801 (N_801,N_583,N_687);
nor U802 (N_802,In_280,In_649);
or U803 (N_803,In_1479,In_197);
nor U804 (N_804,In_690,In_633);
nand U805 (N_805,In_693,N_224);
and U806 (N_806,In_258,N_443);
and U807 (N_807,N_162,N_354);
or U808 (N_808,In_362,N_717);
nand U809 (N_809,In_477,In_92);
nor U810 (N_810,In_2108,In_1439);
or U811 (N_811,In_22,In_1513);
or U812 (N_812,In_1977,In_2281);
nand U813 (N_813,In_1901,In_1153);
nor U814 (N_814,In_1177,In_4);
nor U815 (N_815,In_2012,N_551);
nor U816 (N_816,In_109,N_280);
or U817 (N_817,N_613,N_640);
or U818 (N_818,N_254,In_2077);
xor U819 (N_819,N_396,N_586);
and U820 (N_820,In_1236,N_363);
nor U821 (N_821,In_2149,In_921);
nand U822 (N_822,N_189,In_324);
and U823 (N_823,N_762,In_1884);
and U824 (N_824,In_777,N_788);
and U825 (N_825,N_208,In_2187);
or U826 (N_826,In_584,N_206);
nor U827 (N_827,In_667,N_723);
or U828 (N_828,N_708,In_5);
and U829 (N_829,In_552,In_1190);
and U830 (N_830,In_2378,In_2422);
nor U831 (N_831,In_1317,In_2123);
or U832 (N_832,In_945,In_587);
and U833 (N_833,N_685,In_336);
nor U834 (N_834,In_1557,In_534);
xor U835 (N_835,N_218,In_2296);
and U836 (N_836,In_908,In_2289);
nand U837 (N_837,In_498,In_1550);
nor U838 (N_838,In_81,In_1656);
and U839 (N_839,N_411,In_1878);
xnor U840 (N_840,In_2189,In_1162);
xor U841 (N_841,In_2073,N_440);
and U842 (N_842,N_514,In_2465);
nand U843 (N_843,N_713,In_1396);
xnor U844 (N_844,In_1696,N_545);
nor U845 (N_845,In_1457,N_178);
nor U846 (N_846,In_2285,In_603);
nand U847 (N_847,In_2446,In_730);
or U848 (N_848,N_580,In_219);
xor U849 (N_849,In_2410,In_609);
xnor U850 (N_850,In_148,In_2306);
nand U851 (N_851,N_111,In_1899);
and U852 (N_852,In_578,In_1359);
or U853 (N_853,In_62,In_573);
nor U854 (N_854,N_722,In_540);
and U855 (N_855,In_1869,In_1420);
nor U856 (N_856,In_2393,In_1228);
or U857 (N_857,In_630,In_393);
or U858 (N_858,In_85,In_1335);
and U859 (N_859,In_161,In_1271);
xor U860 (N_860,N_589,In_563);
nand U861 (N_861,In_1858,In_1430);
xor U862 (N_862,N_268,N_768);
or U863 (N_863,N_508,N_503);
xnor U864 (N_864,In_620,N_310);
xor U865 (N_865,In_861,In_472);
and U866 (N_866,In_1239,N_31);
nor U867 (N_867,N_607,In_1476);
nand U868 (N_868,In_2114,In_2260);
nand U869 (N_869,In_697,N_424);
nand U870 (N_870,In_185,In_1779);
nor U871 (N_871,In_1619,In_613);
or U872 (N_872,In_1595,N_221);
and U873 (N_873,In_1312,In_990);
or U874 (N_874,N_764,In_165);
xnor U875 (N_875,In_1160,In_223);
xor U876 (N_876,In_2320,N_217);
nand U877 (N_877,In_1765,In_238);
nor U878 (N_878,N_686,In_2419);
or U879 (N_879,In_8,N_400);
and U880 (N_880,In_984,In_120);
nor U881 (N_881,N_694,In_462);
nand U882 (N_882,N_77,In_607);
nor U883 (N_883,In_1187,N_616);
or U884 (N_884,In_2328,N_472);
xor U885 (N_885,In_2088,N_203);
nand U886 (N_886,In_629,In_780);
or U887 (N_887,N_750,In_766);
nand U888 (N_888,In_1093,N_427);
nor U889 (N_889,In_1315,N_515);
nand U890 (N_890,N_577,In_2148);
or U891 (N_891,N_113,N_729);
nand U892 (N_892,In_1563,In_80);
xor U893 (N_893,N_349,In_2129);
and U894 (N_894,In_549,In_776);
nand U895 (N_895,In_1176,N_600);
nand U896 (N_896,N_614,N_604);
nand U897 (N_897,N_735,N_117);
and U898 (N_898,In_824,In_1436);
xnor U899 (N_899,In_683,In_716);
nand U900 (N_900,In_453,In_1370);
or U901 (N_901,N_353,In_2243);
nor U902 (N_902,N_730,In_1075);
and U903 (N_903,In_1677,N_459);
and U904 (N_904,N_581,In_2426);
or U905 (N_905,In_966,In_1627);
xnor U906 (N_906,N_767,In_455);
nor U907 (N_907,In_30,N_643);
xor U908 (N_908,In_639,N_27);
nand U909 (N_909,N_632,In_493);
xnor U910 (N_910,In_110,N_645);
nand U911 (N_911,N_474,In_1962);
nand U912 (N_912,N_314,In_1205);
xor U913 (N_913,In_1564,In_2356);
xor U914 (N_914,In_1449,In_1276);
and U915 (N_915,In_768,In_514);
xnor U916 (N_916,In_1039,N_133);
xnor U917 (N_917,In_1087,N_618);
xnor U918 (N_918,N_437,In_1463);
or U919 (N_919,In_2244,In_1478);
or U920 (N_920,In_2074,N_175);
nor U921 (N_921,N_428,In_581);
and U922 (N_922,N_770,In_1782);
nand U923 (N_923,In_672,In_546);
xor U924 (N_924,N_258,In_2297);
xnor U925 (N_925,In_2205,N_596);
nor U926 (N_926,N_778,N_345);
nor U927 (N_927,N_272,In_2141);
and U928 (N_928,In_404,N_98);
or U929 (N_929,N_260,In_1379);
nand U930 (N_930,In_2204,In_2075);
nand U931 (N_931,N_705,In_1467);
nand U932 (N_932,In_2268,In_1002);
and U933 (N_933,N_564,In_1475);
xor U934 (N_934,In_898,N_573);
xnor U935 (N_935,N_151,N_530);
nor U936 (N_936,N_543,In_1750);
nand U937 (N_937,In_2137,In_1818);
nor U938 (N_938,N_712,In_46);
nor U939 (N_939,N_481,In_1131);
xnor U940 (N_940,In_577,In_2390);
xnor U941 (N_941,In_2010,In_320);
nor U942 (N_942,N_64,In_1032);
nand U943 (N_943,In_230,In_1259);
nand U944 (N_944,N_630,N_97);
and U945 (N_945,N_276,In_1122);
nor U946 (N_946,In_1658,In_2350);
nor U947 (N_947,In_2046,In_2057);
and U948 (N_948,In_225,N_334);
or U949 (N_949,In_579,In_1241);
nor U950 (N_950,N_212,N_408);
and U951 (N_951,In_357,N_156);
nor U952 (N_952,In_98,N_709);
and U953 (N_953,In_1533,N_755);
and U954 (N_954,In_178,In_2433);
and U955 (N_955,N_390,In_2146);
nand U956 (N_956,N_387,N_751);
nand U957 (N_957,In_1774,In_447);
or U958 (N_958,In_1398,In_1221);
nand U959 (N_959,In_135,In_1192);
and U960 (N_960,In_1305,In_2429);
nand U961 (N_961,N_282,In_2365);
nand U962 (N_962,In_991,N_71);
nor U963 (N_963,In_708,N_159);
and U964 (N_964,In_464,N_779);
or U965 (N_965,In_2041,In_890);
and U966 (N_966,N_183,N_124);
nand U967 (N_967,N_634,N_376);
xor U968 (N_968,N_537,In_1622);
and U969 (N_969,In_1488,In_1319);
nand U970 (N_970,N_308,In_2064);
nand U971 (N_971,In_1477,In_929);
xor U972 (N_972,In_684,N_490);
nand U973 (N_973,In_1965,N_182);
xor U974 (N_974,In_694,In_657);
xor U975 (N_975,N_511,In_2366);
and U976 (N_976,In_2101,N_570);
or U977 (N_977,N_665,In_340);
or U978 (N_978,N_690,In_2330);
and U979 (N_979,In_29,N_741);
nor U980 (N_980,N_343,N_718);
or U981 (N_981,In_1616,In_382);
nor U982 (N_982,In_200,In_2403);
and U983 (N_983,In_1584,In_1628);
or U984 (N_984,N_652,N_635);
nor U985 (N_985,In_40,In_405);
and U986 (N_986,In_1610,N_450);
nor U987 (N_987,In_1978,In_1743);
xnor U988 (N_988,N_303,In_753);
or U989 (N_989,In_181,In_244);
or U990 (N_990,N_485,In_2309);
or U991 (N_991,N_92,N_114);
nor U992 (N_992,N_347,N_526);
or U993 (N_993,N_340,In_2063);
nand U994 (N_994,N_782,In_952);
nand U995 (N_995,In_1928,In_769);
nor U996 (N_996,N_641,N_683);
xnor U997 (N_997,In_2314,In_261);
xor U998 (N_998,In_651,N_296);
and U999 (N_999,In_492,In_2424);
nor U1000 (N_1000,In_1840,N_283);
xor U1001 (N_1001,In_1586,N_766);
nand U1002 (N_1002,In_1053,N_333);
or U1003 (N_1003,In_662,In_1814);
nand U1004 (N_1004,In_1100,In_2331);
and U1005 (N_1005,N_519,N_318);
or U1006 (N_1006,In_195,N_693);
nand U1007 (N_1007,In_2395,In_1199);
nor U1008 (N_1008,In_1794,N_650);
nor U1009 (N_1009,In_2327,In_618);
nand U1010 (N_1010,In_2230,N_931);
and U1011 (N_1011,In_2364,N_316);
nor U1012 (N_1012,In_1225,N_281);
nand U1013 (N_1013,In_366,In_375);
and U1014 (N_1014,In_1581,In_1195);
nor U1015 (N_1015,N_94,In_28);
nand U1016 (N_1016,In_1120,In_1362);
nand U1017 (N_1017,In_1843,In_1836);
nand U1018 (N_1018,In_1460,N_454);
xor U1019 (N_1019,In_1069,N_807);
nand U1020 (N_1020,N_223,In_519);
or U1021 (N_1021,In_574,N_468);
nor U1022 (N_1022,In_887,In_2464);
or U1023 (N_1023,In_2458,In_2145);
nor U1024 (N_1024,N_689,In_1778);
xnor U1025 (N_1025,In_1987,N_822);
xnor U1026 (N_1026,In_642,N_315);
nor U1027 (N_1027,In_1886,In_548);
nor U1028 (N_1028,N_636,In_1492);
or U1029 (N_1029,N_681,N_267);
or U1030 (N_1030,N_803,In_61);
nand U1031 (N_1031,N_845,In_413);
or U1032 (N_1032,N_753,In_1223);
and U1033 (N_1033,N_734,In_1607);
nor U1034 (N_1034,In_1473,In_18);
or U1035 (N_1035,In_299,N_981);
or U1036 (N_1036,N_628,N_317);
nand U1037 (N_1037,In_2095,In_1933);
or U1038 (N_1038,N_528,N_531);
nor U1039 (N_1039,In_930,In_1825);
nand U1040 (N_1040,N_309,N_355);
nand U1041 (N_1041,N_886,N_5);
nor U1042 (N_1042,N_20,In_2291);
nand U1043 (N_1043,N_453,In_647);
and U1044 (N_1044,In_1330,In_528);
nor U1045 (N_1045,In_391,N_838);
or U1046 (N_1046,In_1958,In_191);
xor U1047 (N_1047,N_972,In_828);
nor U1048 (N_1048,In_1732,N_76);
and U1049 (N_1049,N_900,In_153);
or U1050 (N_1050,N_606,In_1390);
or U1051 (N_1051,In_1636,In_815);
or U1052 (N_1052,In_1269,In_2467);
xnor U1053 (N_1053,In_397,In_310);
and U1054 (N_1054,In_737,In_1159);
nor U1055 (N_1055,N_654,In_1817);
or U1056 (N_1056,In_302,N_974);
or U1057 (N_1057,N_728,In_886);
nor U1058 (N_1058,N_14,In_1892);
or U1059 (N_1059,In_2215,In_2427);
nand U1060 (N_1060,In_1304,In_1860);
and U1061 (N_1061,In_9,N_305);
or U1062 (N_1062,In_2059,In_871);
nor U1063 (N_1063,N_877,In_1543);
and U1064 (N_1064,In_1300,In_126);
nor U1065 (N_1065,In_781,N_209);
nor U1066 (N_1066,N_228,N_872);
or U1067 (N_1067,In_1546,In_1248);
or U1068 (N_1068,N_839,In_2361);
and U1069 (N_1069,N_389,In_750);
or U1070 (N_1070,In_1984,In_1588);
or U1071 (N_1071,In_741,In_1352);
nand U1072 (N_1072,In_1998,In_2383);
nor U1073 (N_1073,In_1285,In_2435);
nor U1074 (N_1074,N_648,In_198);
xor U1075 (N_1075,In_1074,N_827);
or U1076 (N_1076,N_952,N_95);
and U1077 (N_1077,In_1115,In_56);
nand U1078 (N_1078,N_664,In_571);
and U1079 (N_1079,In_1652,N_235);
or U1080 (N_1080,In_1655,In_2005);
nand U1081 (N_1081,In_1731,In_638);
and U1082 (N_1082,N_300,N_143);
nand U1083 (N_1083,N_757,In_216);
or U1084 (N_1084,In_1371,N_404);
nor U1085 (N_1085,N_667,N_13);
and U1086 (N_1086,In_634,In_510);
xor U1087 (N_1087,In_496,In_2214);
or U1088 (N_1088,N_948,In_751);
nand U1089 (N_1089,N_480,In_1608);
nor U1090 (N_1090,N_668,N_179);
xnor U1091 (N_1091,In_516,N_985);
or U1092 (N_1092,N_631,In_1664);
and U1093 (N_1093,In_2252,In_674);
and U1094 (N_1094,N_116,N_940);
xnor U1095 (N_1095,In_2081,In_1306);
and U1096 (N_1096,In_2152,N_611);
nor U1097 (N_1097,N_740,In_1219);
nor U1098 (N_1098,In_924,N_832);
and U1099 (N_1099,N_594,In_858);
nor U1100 (N_1100,In_822,In_1332);
or U1101 (N_1101,N_953,In_1944);
nor U1102 (N_1102,N_957,In_1816);
nor U1103 (N_1103,In_728,N_855);
nand U1104 (N_1104,N_529,In_438);
nor U1105 (N_1105,In_495,In_1735);
and U1106 (N_1106,In_1405,In_1495);
or U1107 (N_1107,In_2201,In_2218);
nor U1108 (N_1108,N_678,In_377);
and U1109 (N_1109,In_899,In_220);
xor U1110 (N_1110,N_656,In_2287);
nand U1111 (N_1111,N_644,N_892);
nand U1112 (N_1112,In_1555,N_568);
nor U1113 (N_1113,N_164,N_763);
nand U1114 (N_1114,N_874,In_282);
xor U1115 (N_1115,In_713,N_888);
xor U1116 (N_1116,In_1686,In_1286);
and U1117 (N_1117,In_127,N_557);
xnor U1118 (N_1118,N_798,In_179);
nor U1119 (N_1119,In_409,In_1689);
nor U1120 (N_1120,N_386,N_325);
nand U1121 (N_1121,In_2254,N_629);
or U1122 (N_1122,In_524,In_121);
xnor U1123 (N_1123,In_434,In_144);
nor U1124 (N_1124,In_2462,In_2036);
xnor U1125 (N_1125,N_801,In_1561);
nor U1126 (N_1126,In_207,In_2431);
nand U1127 (N_1127,N_620,In_936);
and U1128 (N_1128,In_735,N_914);
nor U1129 (N_1129,In_122,In_188);
and U1130 (N_1130,N_772,N_780);
and U1131 (N_1131,N_736,N_971);
nand U1132 (N_1132,In_2468,In_2126);
nor U1133 (N_1133,N_739,N_338);
nor U1134 (N_1134,In_2092,N_523);
and U1135 (N_1135,In_1623,In_2180);
and U1136 (N_1136,In_599,N_731);
or U1137 (N_1137,In_2227,In_97);
or U1138 (N_1138,N_851,In_2347);
nor U1139 (N_1139,In_1890,In_1220);
nor U1140 (N_1140,In_933,N_857);
xnor U1141 (N_1141,N_177,In_2188);
and U1142 (N_1142,In_2229,In_1392);
and U1143 (N_1143,In_1692,In_143);
and U1144 (N_1144,N_541,In_1511);
and U1145 (N_1145,N_704,N_861);
nor U1146 (N_1146,In_1697,In_1716);
nand U1147 (N_1147,N_847,In_159);
or U1148 (N_1148,In_1025,N_465);
nor U1149 (N_1149,N_599,In_271);
nand U1150 (N_1150,In_687,N_979);
or U1151 (N_1151,N_401,In_2082);
nand U1152 (N_1152,In_316,In_1537);
nor U1153 (N_1153,N_274,In_1974);
and U1154 (N_1154,N_987,In_386);
and U1155 (N_1155,N_792,In_416);
nand U1156 (N_1156,In_317,N_602);
nand U1157 (N_1157,In_2412,N_65);
and U1158 (N_1158,N_921,In_1876);
xor U1159 (N_1159,In_2172,In_1365);
nand U1160 (N_1160,N_451,In_1073);
or U1161 (N_1161,N_7,In_114);
nand U1162 (N_1162,N_929,In_70);
nor U1163 (N_1163,In_2211,In_152);
xor U1164 (N_1164,In_1059,In_1401);
nor U1165 (N_1165,In_1461,In_1579);
nand U1166 (N_1166,In_1777,In_1243);
nand U1167 (N_1167,N_899,In_536);
and U1168 (N_1168,N_902,In_1141);
nor U1169 (N_1169,In_91,N_674);
xor U1170 (N_1170,In_424,In_686);
xnor U1171 (N_1171,N_433,N_39);
xor U1172 (N_1172,In_412,In_632);
nand U1173 (N_1173,N_785,N_505);
xnor U1174 (N_1174,In_333,In_2103);
nand U1175 (N_1175,In_1423,In_253);
nand U1176 (N_1176,N_714,N_826);
and U1177 (N_1177,In_1320,In_444);
nand U1178 (N_1178,N_653,N_771);
nand U1179 (N_1179,In_909,In_1152);
nand U1180 (N_1180,In_2307,In_1604);
xor U1181 (N_1181,In_1366,In_303);
xnor U1182 (N_1182,In_1060,N_858);
nand U1183 (N_1183,In_2496,In_688);
nor U1184 (N_1184,N_312,N_488);
nor U1185 (N_1185,N_533,In_1996);
nor U1186 (N_1186,N_759,In_1172);
or U1187 (N_1187,In_807,N_370);
nand U1188 (N_1188,In_1671,In_117);
nor U1189 (N_1189,In_1558,In_1685);
nor U1190 (N_1190,N_662,N_817);
nand U1191 (N_1191,N_403,In_999);
xnor U1192 (N_1192,In_677,N_371);
and U1193 (N_1193,In_51,N_701);
and U1194 (N_1194,In_2360,In_1970);
nor U1195 (N_1195,N_744,In_233);
nor U1196 (N_1196,In_2399,In_1256);
nand U1197 (N_1197,In_1144,In_482);
or U1198 (N_1198,N_441,In_932);
nor U1199 (N_1199,In_1556,In_2282);
nand U1200 (N_1200,In_2315,N_149);
nor U1201 (N_1201,In_1669,N_715);
or U1202 (N_1202,In_1803,N_680);
nand U1203 (N_1203,N_544,N_247);
or U1204 (N_1204,N_1024,N_32);
xor U1205 (N_1205,N_256,In_625);
xnor U1206 (N_1206,In_2207,N_840);
or U1207 (N_1207,N_1012,In_1166);
or U1208 (N_1208,In_2094,N_621);
nor U1209 (N_1209,In_2402,In_423);
or U1210 (N_1210,N_1025,N_783);
and U1211 (N_1211,In_1337,In_2302);
xnor U1212 (N_1212,In_544,In_1888);
nand U1213 (N_1213,In_2341,N_1054);
or U1214 (N_1214,N_878,N_608);
and U1215 (N_1215,N_135,N_193);
nor U1216 (N_1216,In_1281,N_1089);
nand U1217 (N_1217,N_846,N_269);
nand U1218 (N_1218,In_2375,In_2000);
nor U1219 (N_1219,N_1048,In_1394);
nor U1220 (N_1220,N_889,N_672);
xor U1221 (N_1221,In_2319,N_1081);
xor U1222 (N_1222,N_898,In_1017);
nor U1223 (N_1223,N_295,N_1046);
xnor U1224 (N_1224,In_640,N_943);
nand U1225 (N_1225,In_500,In_1720);
nand U1226 (N_1226,N_1007,N_989);
or U1227 (N_1227,N_880,In_99);
and U1228 (N_1228,N_691,In_10);
nand U1229 (N_1229,N_990,N_733);
and U1230 (N_1230,N_738,N_1098);
nand U1231 (N_1231,In_1179,In_1260);
and U1232 (N_1232,N_560,In_1118);
or U1233 (N_1233,In_1993,In_1866);
nand U1234 (N_1234,N_844,N_100);
and U1235 (N_1235,In_2477,In_1861);
nand U1236 (N_1236,N_47,In_1194);
and U1237 (N_1237,N_603,N_799);
nand U1238 (N_1238,In_2048,In_2233);
nand U1239 (N_1239,In_617,In_1650);
and U1240 (N_1240,In_1932,In_2131);
nor U1241 (N_1241,N_956,In_996);
and U1242 (N_1242,In_2479,N_460);
or U1243 (N_1243,N_181,N_381);
xor U1244 (N_1244,N_639,In_283);
nor U1245 (N_1245,N_16,N_336);
xor U1246 (N_1246,N_1103,N_811);
nand U1247 (N_1247,In_288,In_1197);
nor U1248 (N_1248,In_166,N_834);
nand U1249 (N_1249,N_2,In_547);
nor U1250 (N_1250,In_1127,N_935);
xnor U1251 (N_1251,In_1347,In_1859);
or U1252 (N_1252,N_1004,In_834);
nor U1253 (N_1253,In_359,N_835);
or U1254 (N_1254,N_890,N_75);
nand U1255 (N_1255,N_1102,N_434);
nor U1256 (N_1256,N_25,N_679);
or U1257 (N_1257,N_754,In_794);
and U1258 (N_1258,In_2409,N_571);
or U1259 (N_1259,In_2270,In_89);
xor U1260 (N_1260,N_1149,N_946);
nor U1261 (N_1261,In_2006,In_168);
nor U1262 (N_1262,N_91,In_1678);
nand U1263 (N_1263,In_123,In_543);
and U1264 (N_1264,N_554,In_479);
nor U1265 (N_1265,In_1705,In_928);
nand U1266 (N_1266,N_126,In_1116);
nand U1267 (N_1267,N_784,In_1354);
nand U1268 (N_1268,N_651,N_327);
or U1269 (N_1269,N_911,N_970);
nand U1270 (N_1270,N_173,N_1055);
nor U1271 (N_1271,N_831,N_1128);
xor U1272 (N_1272,N_565,N_1188);
nand U1273 (N_1273,N_123,In_325);
nand U1274 (N_1274,N_994,In_1534);
and U1275 (N_1275,In_1947,In_342);
xor U1276 (N_1276,N_725,N_867);
and U1277 (N_1277,N_1122,N_998);
nand U1278 (N_1278,N_83,N_969);
and U1279 (N_1279,In_859,N_1067);
nor U1280 (N_1280,In_1294,In_791);
nand U1281 (N_1281,N_40,N_1143);
xor U1282 (N_1282,N_1121,In_1417);
nor U1283 (N_1283,N_1082,N_595);
or U1284 (N_1284,N_669,N_1156);
xor U1285 (N_1285,In_2202,N_1135);
nand U1286 (N_1286,In_512,N_917);
xnor U1287 (N_1287,N_816,In_164);
xor U1288 (N_1288,In_1526,N_395);
and U1289 (N_1289,In_442,N_579);
nor U1290 (N_1290,In_1323,In_1790);
and U1291 (N_1291,N_702,In_27);
nand U1292 (N_1292,In_608,In_1343);
or U1293 (N_1293,In_432,In_749);
xnor U1294 (N_1294,N_895,N_237);
and U1295 (N_1295,N_539,N_700);
nand U1296 (N_1296,N_1070,N_1120);
or U1297 (N_1297,In_876,N_1006);
and U1298 (N_1298,In_1376,N_897);
xor U1299 (N_1299,In_414,N_1178);
and U1300 (N_1300,N_1065,In_967);
or U1301 (N_1301,In_725,In_590);
nand U1302 (N_1302,N_532,In_2100);
and U1303 (N_1303,N_626,In_2105);
nor U1304 (N_1304,In_2323,N_1137);
nand U1305 (N_1305,In_520,N_697);
xor U1306 (N_1306,In_1212,N_299);
nor U1307 (N_1307,In_2355,N_410);
or U1308 (N_1308,N_1152,N_1002);
xor U1309 (N_1309,In_958,In_1130);
xor U1310 (N_1310,In_1880,In_2336);
and U1311 (N_1311,N_800,In_979);
or U1312 (N_1312,N_1040,N_1190);
or U1313 (N_1313,In_1991,In_285);
or U1314 (N_1314,In_902,N_439);
or U1315 (N_1315,In_1198,N_103);
nor U1316 (N_1316,In_364,N_302);
or U1317 (N_1317,N_789,N_293);
nor U1318 (N_1318,In_1386,In_1498);
nand U1319 (N_1319,In_190,In_602);
or U1320 (N_1320,N_756,In_1775);
xnor U1321 (N_1321,In_2445,N_1088);
nor U1322 (N_1322,N_732,N_869);
nand U1323 (N_1323,N_646,In_539);
or U1324 (N_1324,N_1184,N_242);
nor U1325 (N_1325,N_837,N_742);
nor U1326 (N_1326,In_636,N_794);
nor U1327 (N_1327,N_1196,In_2037);
nor U1328 (N_1328,In_869,N_1182);
and U1329 (N_1329,In_983,In_1325);
or U1330 (N_1330,In_910,In_242);
or U1331 (N_1331,In_691,N_982);
xor U1332 (N_1332,In_831,In_706);
nand U1333 (N_1333,N_623,In_699);
or U1334 (N_1334,N_884,N_1021);
nor U1335 (N_1335,In_1327,N_464);
nand U1336 (N_1336,N_777,In_692);
nor U1337 (N_1337,In_2300,In_1681);
or U1338 (N_1338,N_941,N_876);
nor U1339 (N_1339,In_833,In_335);
nor U1340 (N_1340,N_813,In_2200);
or U1341 (N_1341,N_417,N_1154);
xor U1342 (N_1342,N_776,In_1708);
nand U1343 (N_1343,N_879,N_699);
nand U1344 (N_1344,N_1175,N_1014);
xor U1345 (N_1345,In_720,N_1195);
and U1346 (N_1346,N_655,In_1649);
or U1347 (N_1347,N_160,In_1613);
nor U1348 (N_1348,N_510,In_475);
nand U1349 (N_1349,N_146,N_804);
nand U1350 (N_1350,In_2396,In_1904);
nand U1351 (N_1351,In_1913,In_820);
and U1352 (N_1352,N_590,In_1573);
or U1353 (N_1353,In_1349,In_1871);
and U1354 (N_1354,N_932,N_392);
nand U1355 (N_1355,N_810,N_913);
nor U1356 (N_1356,In_1215,N_1084);
and U1357 (N_1357,N_422,N_416);
xnor U1358 (N_1358,In_541,N_942);
nor U1359 (N_1359,In_2346,N_961);
or U1360 (N_1360,In_34,In_1937);
xor U1361 (N_1361,N_1126,In_1252);
nor U1362 (N_1362,N_205,In_1575);
or U1363 (N_1363,In_1334,In_57);
nand U1364 (N_1364,N_446,In_1003);
or U1365 (N_1365,In_277,N_964);
or U1366 (N_1366,N_894,In_1326);
nand U1367 (N_1367,In_1066,In_146);
nand U1368 (N_1368,In_878,N_1170);
nand U1369 (N_1369,N_225,N_1020);
nand U1370 (N_1370,N_657,N_1066);
xnor U1371 (N_1371,In_1246,N_951);
and U1372 (N_1372,In_456,N_1011);
and U1373 (N_1373,N_647,In_742);
nand U1374 (N_1374,In_2377,N_842);
nand U1375 (N_1375,N_1008,In_2448);
xor U1376 (N_1376,In_1834,N_501);
and U1377 (N_1377,In_1516,N_988);
or U1378 (N_1378,N_605,In_1552);
and U1379 (N_1379,In_648,In_1709);
and U1380 (N_1380,In_1363,In_1585);
or U1381 (N_1381,N_758,N_1181);
xnor U1382 (N_1382,N_1139,In_752);
or U1383 (N_1383,N_457,N_412);
or U1384 (N_1384,N_84,N_1198);
nand U1385 (N_1385,In_1501,In_2162);
or U1386 (N_1386,N_394,In_1418);
or U1387 (N_1387,In_1930,N_1042);
and U1388 (N_1388,In_1632,In_1905);
or U1389 (N_1389,In_1270,N_588);
nand U1390 (N_1390,In_2144,N_671);
xnor U1391 (N_1391,In_743,N_506);
and U1392 (N_1392,N_1155,N_1074);
nor U1393 (N_1393,N_337,N_860);
and U1394 (N_1394,N_1013,N_703);
nor U1395 (N_1395,In_655,In_701);
nor U1396 (N_1396,In_880,In_1368);
nand U1397 (N_1397,N_825,N_802);
nor U1398 (N_1398,In_1422,N_1174);
nand U1399 (N_1399,N_1124,N_147);
or U1400 (N_1400,N_1279,N_1211);
nand U1401 (N_1401,N_456,N_1290);
nor U1402 (N_1402,N_1230,N_676);
nor U1403 (N_1403,In_1083,N_119);
nand U1404 (N_1404,In_2024,N_1250);
xor U1405 (N_1405,In_173,N_936);
xor U1406 (N_1406,In_2354,N_666);
and U1407 (N_1407,N_761,N_1242);
nand U1408 (N_1408,N_158,N_1058);
nand U1409 (N_1409,N_1160,N_1232);
xor U1410 (N_1410,N_1083,In_1076);
nand U1411 (N_1411,N_1161,In_309);
xor U1412 (N_1412,In_2381,N_1367);
xnor U1413 (N_1413,N_983,In_287);
nor U1414 (N_1414,N_1237,In_1019);
or U1415 (N_1415,In_2486,N_1261);
or U1416 (N_1416,In_969,N_190);
nand U1417 (N_1417,N_1256,N_881);
nand U1418 (N_1418,In_33,In_1948);
nor U1419 (N_1419,N_745,In_1635);
or U1420 (N_1420,N_769,N_711);
or U1421 (N_1421,N_1354,N_1339);
nor U1422 (N_1422,N_478,N_43);
nand U1423 (N_1423,N_995,N_1043);
and U1424 (N_1424,N_1381,N_1248);
nand U1425 (N_1425,In_2183,In_829);
nor U1426 (N_1426,N_1059,In_83);
or U1427 (N_1427,N_1303,N_1390);
xnor U1428 (N_1428,N_1169,In_1762);
or U1429 (N_1429,N_1185,In_1745);
nor U1430 (N_1430,In_623,N_1313);
xnor U1431 (N_1431,In_1040,N_737);
nor U1432 (N_1432,N_341,In_327);
nand U1433 (N_1433,N_795,N_1322);
xor U1434 (N_1434,In_2226,In_889);
xor U1435 (N_1435,N_1377,N_1147);
and U1436 (N_1436,N_498,N_821);
nand U1437 (N_1437,N_1387,In_2171);
or U1438 (N_1438,In_650,N_1111);
xor U1439 (N_1439,N_172,N_569);
and U1440 (N_1440,In_497,In_221);
nand U1441 (N_1441,N_388,N_63);
xnor U1442 (N_1442,In_872,In_811);
nand U1443 (N_1443,N_849,In_2021);
or U1444 (N_1444,In_1133,In_582);
nand U1445 (N_1445,N_1252,N_1300);
xor U1446 (N_1446,N_1278,In_118);
or U1447 (N_1447,N_1353,In_112);
nand U1448 (N_1448,In_2035,N_885);
xor U1449 (N_1449,N_1085,N_806);
xor U1450 (N_1450,N_1101,N_461);
nor U1451 (N_1451,N_793,N_1123);
or U1452 (N_1452,In_151,In_2305);
nand U1453 (N_1453,N_263,N_1281);
or U1454 (N_1454,N_727,In_1207);
and U1455 (N_1455,In_1222,In_466);
nor U1456 (N_1456,N_1213,N_698);
xor U1457 (N_1457,N_1396,In_401);
and U1458 (N_1458,In_1485,In_682);
or U1459 (N_1459,N_487,In_947);
or U1460 (N_1460,In_875,N_760);
nand U1461 (N_1461,In_1369,In_2099);
or U1462 (N_1462,N_547,N_1037);
or U1463 (N_1463,N_1323,N_1249);
xnor U1464 (N_1464,In_1064,In_1701);
xnor U1465 (N_1465,N_805,N_854);
and U1466 (N_1466,In_1827,N_1286);
xnor U1467 (N_1467,In_641,In_1465);
xor U1468 (N_1468,N_1372,N_1119);
nand U1469 (N_1469,N_947,N_833);
and U1470 (N_1470,In_1535,N_1344);
or U1471 (N_1471,N_1331,In_1472);
nand U1472 (N_1472,In_1150,In_2197);
nor U1473 (N_1473,N_1157,In_2150);
or U1474 (N_1474,N_871,N_1116);
and U1475 (N_1475,N_1105,N_1192);
or U1476 (N_1476,In_212,N_1333);
or U1477 (N_1477,N_1253,N_517);
xor U1478 (N_1478,N_1221,In_1095);
and U1479 (N_1479,N_903,In_2239);
or U1480 (N_1480,In_956,N_1041);
nor U1481 (N_1481,In_867,In_2224);
and U1482 (N_1482,In_1462,N_1238);
or U1483 (N_1483,N_1057,N_1138);
nor U1484 (N_1484,N_1366,N_21);
nand U1485 (N_1485,N_278,In_384);
and U1486 (N_1486,N_1321,N_1282);
and U1487 (N_1487,In_239,In_1071);
and U1488 (N_1488,N_536,N_598);
xor U1489 (N_1489,N_1394,N_1224);
and U1490 (N_1490,In_1105,In_1643);
nand U1491 (N_1491,In_894,In_2231);
xor U1492 (N_1492,N_1327,In_862);
nor U1493 (N_1493,In_661,In_1889);
xnor U1494 (N_1494,N_458,In_1926);
nand U1495 (N_1495,In_2191,N_965);
nor U1496 (N_1496,In_940,In_2089);
xnor U1497 (N_1497,In_491,N_642);
nor U1498 (N_1498,N_1310,In_1086);
and U1499 (N_1499,In_954,In_1882);
xor U1500 (N_1500,N_843,N_1148);
nand U1501 (N_1501,In_294,In_2481);
or U1502 (N_1502,In_2185,In_103);
xor U1503 (N_1503,N_1251,In_731);
xor U1504 (N_1504,N_466,N_786);
nor U1505 (N_1505,In_350,N_1150);
nand U1506 (N_1506,In_1114,In_2389);
xor U1507 (N_1507,In_2437,In_1699);
and U1508 (N_1508,In_1250,N_920);
or U1509 (N_1509,N_612,In_199);
xor U1510 (N_1510,N_297,N_1115);
and U1511 (N_1511,In_1143,In_69);
nor U1512 (N_1512,N_1358,In_1597);
and U1513 (N_1513,N_1297,N_781);
or U1514 (N_1514,N_1193,N_958);
xor U1515 (N_1515,N_1142,N_567);
and U1516 (N_1516,N_1171,N_1254);
nand U1517 (N_1517,N_1352,In_1036);
nor U1518 (N_1518,In_962,N_908);
and U1519 (N_1519,In_817,In_718);
xor U1520 (N_1520,N_848,N_625);
nor U1521 (N_1521,N_1332,N_774);
nand U1522 (N_1522,N_1355,In_465);
and U1523 (N_1523,In_1992,N_346);
or U1524 (N_1524,In_2192,N_1291);
or U1525 (N_1525,In_2472,N_106);
or U1526 (N_1526,N_1114,In_1902);
and U1527 (N_1527,N_1334,N_724);
nor U1528 (N_1528,N_1241,N_1389);
or U1529 (N_1529,N_624,In_616);
or U1530 (N_1530,In_459,In_1034);
nor U1531 (N_1531,N_978,N_1274);
nand U1532 (N_1532,N_420,N_1240);
nor U1533 (N_1533,N_527,N_452);
nor U1534 (N_1534,N_950,In_44);
xor U1535 (N_1535,In_1094,In_1009);
xor U1536 (N_1536,N_868,N_1199);
or U1537 (N_1537,In_1434,N_572);
and U1538 (N_1538,N_1255,In_2338);
and U1539 (N_1539,In_709,N_1189);
xnor U1540 (N_1540,In_2376,N_168);
or U1541 (N_1541,In_1001,In_748);
and U1542 (N_1542,In_2299,In_2110);
and U1543 (N_1543,In_379,N_1345);
nand U1544 (N_1544,In_1772,N_1365);
and U1545 (N_1545,In_2310,N_719);
nand U1546 (N_1546,In_1357,In_1189);
nor U1547 (N_1547,In_400,In_2278);
or U1548 (N_1548,N_622,In_2353);
nor U1549 (N_1549,In_1,In_719);
or U1550 (N_1550,In_1739,N_1078);
nand U1551 (N_1551,N_841,In_586);
nand U1552 (N_1552,N_927,N_520);
or U1553 (N_1553,N_1266,N_444);
nor U1554 (N_1554,In_868,In_431);
or U1555 (N_1555,N_1306,In_1916);
or U1556 (N_1556,N_1162,In_189);
or U1557 (N_1557,N_1186,N_1273);
xnor U1558 (N_1558,N_1047,In_614);
xnor U1559 (N_1559,N_504,N_1214);
nor U1560 (N_1560,N_1270,N_332);
xnor U1561 (N_1561,N_518,In_1234);
or U1562 (N_1562,In_101,N_1293);
xnor U1563 (N_1563,In_1404,In_2003);
nand U1564 (N_1564,In_458,In_893);
nand U1565 (N_1565,In_1067,In_939);
xor U1566 (N_1566,In_1309,N_1267);
or U1567 (N_1567,N_1271,N_1319);
xnor U1568 (N_1568,N_1093,N_219);
nor U1569 (N_1569,N_1369,N_591);
nand U1570 (N_1570,In_461,N_348);
xnor U1571 (N_1571,In_125,In_2308);
or U1572 (N_1572,N_1376,N_1397);
or U1573 (N_1573,N_1109,N_907);
or U1574 (N_1574,N_285,In_1547);
and U1575 (N_1575,N_1030,N_901);
nor U1576 (N_1576,N_819,N_1315);
xnor U1577 (N_1577,In_1960,N_402);
nand U1578 (N_1578,N_747,N_534);
nand U1579 (N_1579,N_1086,In_1302);
nor U1580 (N_1580,N_1328,In_2416);
or U1581 (N_1581,N_1172,In_1938);
xor U1582 (N_1582,N_1068,N_415);
xor U1583 (N_1583,N_1316,In_1957);
xor U1584 (N_1584,N_1194,In_916);
or U1585 (N_1585,N_1312,N_407);
nor U1586 (N_1586,N_1203,In_1090);
nand U1587 (N_1587,N_1258,N_938);
nor U1588 (N_1588,N_495,N_1045);
xnor U1589 (N_1589,In_264,N_301);
and U1590 (N_1590,N_830,In_1983);
or U1591 (N_1591,In_374,N_1348);
nand U1592 (N_1592,N_548,In_1752);
or U1593 (N_1593,N_659,N_909);
and U1594 (N_1594,In_1811,N_633);
nand U1595 (N_1595,In_140,In_1412);
and U1596 (N_1596,N_1262,N_1341);
xnor U1597 (N_1597,In_1375,N_873);
nor U1598 (N_1598,N_1113,N_883);
or U1599 (N_1599,In_2240,N_1032);
nor U1600 (N_1600,N_649,In_855);
xnor U1601 (N_1601,In_276,In_1169);
nor U1602 (N_1602,N_1305,In_506);
or U1603 (N_1603,N_1320,In_761);
and U1604 (N_1604,N_1598,N_1496);
and U1605 (N_1605,In_643,N_1546);
nor U1606 (N_1606,N_1466,N_1429);
and U1607 (N_1607,In_1080,N_1260);
xor U1608 (N_1608,In_503,N_482);
or U1609 (N_1609,In_439,In_2404);
and U1610 (N_1610,N_856,In_94);
nor U1611 (N_1611,In_526,N_1410);
or U1612 (N_1612,N_773,N_399);
and U1613 (N_1613,N_1404,N_110);
nor U1614 (N_1614,N_1133,N_1452);
or U1615 (N_1615,N_1459,In_1700);
nor U1616 (N_1616,N_1536,N_1295);
and U1617 (N_1617,N_1107,In_2256);
and U1618 (N_1618,N_1212,N_1407);
or U1619 (N_1619,N_1446,In_1956);
xnor U1620 (N_1620,N_967,N_1326);
xnor U1621 (N_1621,N_1337,N_33);
xnor U1622 (N_1622,N_1499,N_1388);
nand U1623 (N_1623,N_1526,In_923);
or U1624 (N_1624,N_1229,In_934);
nand U1625 (N_1625,In_1108,N_1112);
nand U1626 (N_1626,N_1574,In_2386);
and U1627 (N_1627,In_925,N_1289);
xnor U1628 (N_1628,In_68,In_1170);
and U1629 (N_1629,In_1161,N_910);
and U1630 (N_1630,N_1060,N_1371);
nand U1631 (N_1631,N_549,N_1519);
or U1632 (N_1632,N_1514,N_1413);
or U1633 (N_1633,In_529,N_682);
xnor U1634 (N_1634,In_704,In_284);
or U1635 (N_1635,N_413,N_1209);
or U1636 (N_1636,N_609,N_1265);
and U1637 (N_1637,N_136,In_2219);
xor U1638 (N_1638,N_1379,N_928);
and U1639 (N_1639,N_1039,In_854);
nand U1640 (N_1640,In_1413,N_1027);
xor U1641 (N_1641,N_1359,In_1887);
xor U1642 (N_1642,In_955,N_1471);
nand U1643 (N_1643,N_1343,N_1483);
nor U1644 (N_1644,N_1361,N_38);
and U1645 (N_1645,N_617,N_1368);
and U1646 (N_1646,N_862,N_790);
or U1647 (N_1647,In_167,N_1475);
nand U1648 (N_1648,N_1205,In_1935);
or U1649 (N_1649,N_1210,In_1341);
nand U1650 (N_1650,N_1349,N_1426);
nor U1651 (N_1651,N_684,N_1146);
nand U1652 (N_1652,N_1385,N_352);
xnor U1653 (N_1653,In_1990,N_1228);
xnor U1654 (N_1654,In_722,In_2198);
and U1655 (N_1655,N_49,N_1547);
and U1656 (N_1656,N_1392,In_1545);
nand U1657 (N_1657,N_1357,N_58);
nand U1658 (N_1658,N_1324,In_481);
nor U1659 (N_1659,N_1523,In_248);
or U1660 (N_1660,N_829,N_968);
nand U1661 (N_1661,In_2098,In_2304);
nor U1662 (N_1662,N_1201,N_1005);
or U1663 (N_1663,N_896,N_1506);
nand U1664 (N_1664,N_986,N_252);
or U1665 (N_1665,N_1235,N_1482);
nor U1666 (N_1666,N_1460,In_87);
nand U1667 (N_1667,N_1301,N_944);
nor U1668 (N_1668,N_663,In_193);
xnor U1669 (N_1669,N_1393,N_1563);
xnor U1670 (N_1670,N_1208,In_1624);
nand U1671 (N_1671,N_1402,N_696);
nor U1672 (N_1672,In_1031,N_1503);
nand U1673 (N_1673,N_1423,N_1564);
and U1674 (N_1674,In_1496,N_1204);
nor U1675 (N_1675,N_287,N_815);
or U1676 (N_1676,In_2401,N_924);
and U1677 (N_1677,In_213,N_1573);
xor U1678 (N_1678,In_1867,In_260);
or U1679 (N_1679,In_1229,N_1136);
and U1680 (N_1680,N_992,N_865);
nor U1681 (N_1681,N_962,In_186);
or U1682 (N_1682,In_1982,N_69);
nand U1683 (N_1683,N_1480,In_2434);
nor U1684 (N_1684,In_296,N_637);
nor U1685 (N_1685,N_1543,N_1298);
or U1686 (N_1686,In_45,N_1049);
or U1687 (N_1687,N_1364,N_1072);
or U1688 (N_1688,N_1096,N_1104);
and U1689 (N_1689,N_215,In_1233);
or U1690 (N_1690,In_736,In_1280);
xor U1691 (N_1691,N_866,N_1180);
and U1692 (N_1692,In_474,In_2460);
or U1693 (N_1693,N_1223,In_2432);
and U1694 (N_1694,In_378,N_1216);
nor U1695 (N_1695,In_1801,N_1302);
or U1696 (N_1696,In_1088,N_1585);
and U1697 (N_1697,N_852,N_36);
nor U1698 (N_1698,In_130,N_1129);
nor U1699 (N_1699,N_1515,N_1582);
nand U1700 (N_1700,N_1411,N_1167);
or U1701 (N_1701,N_1414,N_1073);
xor U1702 (N_1702,In_913,In_841);
nand U1703 (N_1703,N_1003,In_1591);
xor U1704 (N_1704,N_775,N_1062);
or U1705 (N_1705,N_1053,N_477);
nand U1706 (N_1706,N_1330,N_1165);
and U1707 (N_1707,N_1568,N_1590);
nand U1708 (N_1708,N_1500,In_1020);
xor U1709 (N_1709,N_1560,N_1599);
xnor U1710 (N_1710,N_1552,In_396);
xnor U1711 (N_1711,N_1382,In_1454);
xnor U1712 (N_1712,In_312,N_1097);
xor U1713 (N_1713,N_1491,N_1050);
nand U1714 (N_1714,In_1805,N_748);
xnor U1715 (N_1715,In_2111,N_1549);
nor U1716 (N_1716,N_1340,N_1532);
nand U1717 (N_1717,N_916,In_981);
nand U1718 (N_1718,N_1000,N_585);
nor U1719 (N_1719,N_1197,N_1285);
and U1720 (N_1720,In_808,N_1473);
and U1721 (N_1721,N_1565,N_1474);
xnor U1722 (N_1722,N_710,N_1077);
nand U1723 (N_1723,N_382,N_574);
nor U1724 (N_1724,N_1487,In_537);
nand U1725 (N_1725,N_1449,In_675);
nand U1726 (N_1726,N_1541,N_418);
xnor U1727 (N_1727,In_232,In_2326);
or U1728 (N_1728,N_112,N_1106);
nor U1729 (N_1729,In_311,N_1244);
xnor U1730 (N_1730,N_1153,N_1159);
and U1731 (N_1731,N_432,N_984);
nor U1732 (N_1732,N_265,N_244);
nor U1733 (N_1733,N_1444,In_987);
xor U1734 (N_1734,N_1451,N_675);
nor U1735 (N_1735,N_1399,N_1226);
nand U1736 (N_1736,N_373,N_820);
or U1737 (N_1737,N_1158,In_1846);
nand U1738 (N_1738,In_107,N_1548);
or U1739 (N_1739,N_1569,In_53);
xor U1740 (N_1740,In_2091,In_1149);
or U1741 (N_1741,N_1380,In_1242);
nor U1742 (N_1742,N_1272,N_1516);
nand U1743 (N_1743,N_863,N_1538);
or U1744 (N_1744,N_1467,N_661);
nand U1745 (N_1745,N_507,N_619);
nor U1746 (N_1746,In_2283,N_1534);
xnor U1747 (N_1747,N_421,N_1463);
nand U1748 (N_1748,In_778,N_1477);
nor U1749 (N_1749,In_926,N_1233);
or U1750 (N_1750,N_1183,N_73);
nand U1751 (N_1751,N_555,In_295);
and U1752 (N_1752,N_1558,N_1287);
and U1753 (N_1753,N_937,N_1222);
nor U1754 (N_1754,N_1044,In_1296);
xor U1755 (N_1755,N_1257,N_339);
or U1756 (N_1756,N_186,N_1412);
nand U1757 (N_1757,In_1378,In_1316);
xnor U1758 (N_1758,N_1441,In_128);
nor U1759 (N_1759,N_1447,In_308);
or U1760 (N_1760,N_436,N_1535);
or U1761 (N_1761,N_660,N_320);
or U1762 (N_1762,In_998,N_1099);
and U1763 (N_1763,In_2132,In_1442);
and U1764 (N_1764,N_1571,In_2015);
xnor U1765 (N_1765,N_463,N_1317);
xnor U1766 (N_1766,N_1490,N_1031);
xnor U1767 (N_1767,N_1384,N_1325);
and U1768 (N_1768,N_1511,In_267);
nor U1769 (N_1769,N_1100,In_1796);
nand U1770 (N_1770,N_1508,N_1513);
xnor U1771 (N_1771,N_1061,N_582);
and U1772 (N_1772,In_254,In_1096);
nor U1773 (N_1773,N_429,In_354);
nand U1774 (N_1774,N_1507,In_957);
or U1775 (N_1775,In_1230,N_1405);
xor U1776 (N_1776,In_1614,In_1576);
nand U1777 (N_1777,N_1454,In_2438);
or U1778 (N_1778,N_321,In_1963);
xnor U1779 (N_1779,N_286,N_1567);
xnor U1780 (N_1780,N_976,N_1217);
or U1781 (N_1781,N_253,N_959);
and U1782 (N_1782,N_1069,In_420);
and U1783 (N_1783,N_1479,In_2267);
or U1784 (N_1784,N_1284,N_1362);
nand U1785 (N_1785,N_706,N_814);
nand U1786 (N_1786,N_1218,N_1443);
xnor U1787 (N_1787,In_531,N_1510);
and U1788 (N_1788,N_1438,In_1653);
or U1789 (N_1789,N_695,In_792);
and U1790 (N_1790,N_1434,N_1561);
nor U1791 (N_1791,N_1166,N_250);
nor U1792 (N_1792,N_587,In_281);
xnor U1793 (N_1793,N_1597,In_427);
nor U1794 (N_1794,In_1611,In_739);
nand U1795 (N_1795,N_997,In_2284);
or U1796 (N_1796,N_552,In_1793);
nor U1797 (N_1797,In_1900,N_374);
or U1798 (N_1798,N_1220,N_438);
and U1799 (N_1799,N_1028,N_1283);
and U1800 (N_1800,N_1743,N_905);
xnor U1801 (N_1801,N_500,In_2443);
xor U1802 (N_1802,N_1794,N_949);
and U1803 (N_1803,In_1927,N_1094);
nor U1804 (N_1804,N_1424,In_2251);
xor U1805 (N_1805,N_1386,N_1767);
and U1806 (N_1806,N_1681,N_1329);
nor U1807 (N_1807,N_367,N_1676);
nor U1808 (N_1808,N_1581,N_1610);
and U1809 (N_1809,N_1338,N_1605);
nor U1810 (N_1810,In_844,N_1742);
and U1811 (N_1811,In_773,N_161);
nor U1812 (N_1812,N_1642,N_1431);
nand U1813 (N_1813,In_1936,N_1239);
nand U1814 (N_1814,In_2217,N_578);
and U1815 (N_1815,N_442,N_1580);
or U1816 (N_1816,N_1187,N_1435);
nor U1817 (N_1817,N_298,In_1651);
xnor U1818 (N_1818,N_1033,N_1572);
or U1819 (N_1819,N_1745,In_2071);
or U1820 (N_1820,N_1545,N_1677);
xnor U1821 (N_1821,In_1193,N_1416);
xnor U1822 (N_1822,N_53,N_1036);
and U1823 (N_1823,N_677,In_55);
nand U1824 (N_1824,N_1777,N_1351);
xnor U1825 (N_1825,N_1347,In_480);
or U1826 (N_1826,In_1338,N_1621);
nand U1827 (N_1827,N_996,In_468);
nor U1828 (N_1828,N_1689,In_1102);
nor U1829 (N_1829,N_1234,N_1699);
or U1830 (N_1830,N_1502,In_360);
xor U1831 (N_1831,In_2372,N_1620);
nor U1832 (N_1832,N_1791,N_1691);
and U1833 (N_1833,N_1144,N_369);
and U1834 (N_1834,N_1601,N_1464);
or U1835 (N_1835,N_328,N_121);
and U1836 (N_1836,N_1164,N_1644);
nand U1837 (N_1837,In_1104,N_870);
nor U1838 (N_1838,N_1445,N_1645);
or U1839 (N_1839,N_1646,N_1450);
nor U1840 (N_1840,N_1417,N_1215);
nand U1841 (N_1841,N_1781,N_1163);
and U1842 (N_1842,N_918,In_1506);
nor U1843 (N_1843,N_174,In_1893);
or U1844 (N_1844,N_1420,N_1009);
and U1845 (N_1845,N_509,N_1604);
and U1846 (N_1846,N_1356,N_384);
or U1847 (N_1847,N_1462,N_1064);
or U1848 (N_1848,In_1662,In_866);
xor U1849 (N_1849,N_1653,N_1772);
nand U1850 (N_1850,N_1383,N_1501);
nand U1851 (N_1851,N_1575,In_1646);
nand U1852 (N_1852,N_1108,N_1747);
nand U1853 (N_1853,N_1750,N_812);
nor U1854 (N_1854,In_1123,In_71);
or U1855 (N_1855,N_934,N_1715);
or U1856 (N_1856,In_2134,N_1713);
nor U1857 (N_1857,N_1720,N_1314);
nor U1858 (N_1858,N_1579,N_1754);
nand U1859 (N_1859,N_45,N_1657);
nand U1860 (N_1860,N_380,N_1010);
nor U1861 (N_1861,N_1786,N_1626);
nor U1862 (N_1862,In_215,N_1727);
nand U1863 (N_1863,N_1591,In_2379);
xnor U1864 (N_1864,N_1784,N_720);
xor U1865 (N_1865,In_1994,N_1755);
xnor U1866 (N_1866,N_1264,N_960);
and U1867 (N_1867,N_1736,N_1695);
xnor U1868 (N_1868,N_1746,N_1793);
nor U1869 (N_1869,N_1292,N_726);
and U1870 (N_1870,N_716,N_41);
nor U1871 (N_1871,In_37,In_805);
or U1872 (N_1872,N_1071,N_818);
nand U1873 (N_1873,N_1583,N_1788);
or U1874 (N_1874,N_1652,N_882);
nor U1875 (N_1875,N_1711,N_809);
nand U1876 (N_1876,In_1531,N_1469);
xnor U1877 (N_1877,N_1765,In_1505);
nand U1878 (N_1878,In_2083,In_58);
or U1879 (N_1879,In_1373,N_1613);
nand U1880 (N_1880,N_1176,N_1476);
or U1881 (N_1881,N_1458,N_1650);
or U1882 (N_1882,N_1773,N_1132);
nand U1883 (N_1883,N_1517,N_1465);
xnor U1884 (N_1884,In_2038,N_1639);
nor U1885 (N_1885,N_893,N_1391);
nand U1886 (N_1886,N_1453,N_658);
nor U1887 (N_1887,N_1268,N_923);
and U1888 (N_1888,N_59,N_1732);
or U1889 (N_1889,N_1336,N_796);
and U1890 (N_1890,N_1191,N_1594);
and U1891 (N_1891,N_1553,N_1418);
or U1892 (N_1892,N_1651,In_2120);
nand U1893 (N_1893,N_1373,N_1080);
xor U1894 (N_1894,N_1633,N_1725);
or U1895 (N_1895,N_1075,In_1657);
or U1896 (N_1896,In_1384,In_450);
xnor U1897 (N_1897,In_1594,N_1311);
and U1898 (N_1898,N_1696,N_1769);
nand U1899 (N_1899,N_1015,N_1694);
nand U1900 (N_1900,N_1527,N_1735);
and U1901 (N_1901,N_1001,In_1185);
nor U1902 (N_1902,N_1798,N_1225);
xnor U1903 (N_1903,N_220,N_1436);
nor U1904 (N_1904,N_933,N_1497);
xor U1905 (N_1905,N_1529,N_993);
nor U1906 (N_1906,In_1171,N_1034);
and U1907 (N_1907,N_1687,In_2210);
and U1908 (N_1908,N_1737,N_1643);
nor U1909 (N_1909,N_1706,In_1510);
nand U1910 (N_1910,N_906,In_1703);
xor U1911 (N_1911,N_85,N_1263);
or U1912 (N_1912,N_1678,N_1087);
xnor U1913 (N_1913,N_1611,N_1422);
xnor U1914 (N_1914,N_1576,N_1578);
xor U1915 (N_1915,In_1109,N_279);
nor U1916 (N_1916,N_1638,N_1704);
and U1917 (N_1917,N_1200,In_2042);
or U1918 (N_1918,N_1664,N_1173);
or U1919 (N_1919,N_1702,In_595);
nor U1920 (N_1920,N_1723,N_1342);
nor U1921 (N_1921,N_245,In_1407);
xnor U1922 (N_1922,N_1648,In_1345);
and U1923 (N_1923,N_257,N_1247);
nor U1924 (N_1924,N_1726,N_1202);
nand U1925 (N_1925,N_1540,In_2025);
or U1926 (N_1926,In_1245,N_1022);
nor U1927 (N_1927,N_1682,In_882);
nor U1928 (N_1928,In_1135,N_1029);
nand U1929 (N_1929,N_1468,In_1147);
nand U1930 (N_1930,N_470,In_2151);
xor U1931 (N_1931,N_1596,N_1275);
or U1932 (N_1932,N_904,N_1168);
xor U1933 (N_1933,N_138,N_1647);
xnor U1934 (N_1934,N_1600,N_1577);
xor U1935 (N_1935,N_1219,N_1018);
or U1936 (N_1936,In_1340,N_37);
nor U1937 (N_1937,N_1512,N_1455);
xnor U1938 (N_1938,N_975,N_1486);
nor U1939 (N_1939,In_1857,In_1920);
xnor U1940 (N_1940,In_275,N_379);
nand U1941 (N_1941,In_501,In_1421);
xnor U1942 (N_1942,N_1607,N_1782);
nor U1943 (N_1943,N_1748,N_1672);
and U1944 (N_1944,N_1741,N_1625);
xnor U1945 (N_1945,In_1812,In_14);
and U1946 (N_1946,N_1740,N_1276);
and U1947 (N_1947,N_1588,N_1360);
and U1948 (N_1948,In_1997,In_931);
and U1949 (N_1949,N_1683,N_1494);
xnor U1950 (N_1950,In_1125,N_1131);
nand U1951 (N_1951,N_1472,N_1484);
and U1952 (N_1952,N_1026,N_1243);
or U1953 (N_1953,In_1481,N_1231);
xnor U1954 (N_1954,N_1428,N_1728);
xor U1955 (N_1955,N_1076,N_1309);
or U1956 (N_1956,N_1690,N_66);
nand U1957 (N_1957,N_1738,N_1419);
or U1958 (N_1958,N_1762,N_1721);
or U1959 (N_1959,N_1495,In_2367);
xnor U1960 (N_1960,N_331,In_237);
and U1961 (N_1961,N_1557,N_1634);
and U1962 (N_1962,N_1658,In_487);
nor U1963 (N_1963,N_922,N_1151);
nor U1964 (N_1964,N_1632,N_823);
or U1965 (N_1965,N_1685,N_1584);
xnor U1966 (N_1966,N_1437,N_601);
nor U1967 (N_1967,N_1697,In_1383);
nand U1968 (N_1968,N_1680,N_1606);
nor U1969 (N_1969,N_1245,N_1668);
and U1970 (N_1970,N_1751,N_926);
and U1971 (N_1971,N_1304,N_1731);
and U1972 (N_1972,In_676,N_1141);
or U1973 (N_1973,N_1673,In_911);
nor U1974 (N_1974,In_6,N_1640);
or U1975 (N_1975,N_791,N_1708);
xor U1976 (N_1976,N_1179,N_1378);
or U1977 (N_1977,N_1618,In_557);
nor U1978 (N_1978,N_1017,In_1387);
nand U1979 (N_1979,N_1524,N_1670);
or U1980 (N_1980,N_1662,N_1531);
or U1981 (N_1981,N_1768,N_1530);
and U1982 (N_1982,N_1641,N_610);
xnor U1983 (N_1983,N_864,N_1090);
nand U1984 (N_1984,N_1734,In_874);
and U1985 (N_1985,N_1705,In_2072);
or U1986 (N_1986,N_1749,N_1092);
nor U1987 (N_1987,N_1716,N_836);
nand U1988 (N_1988,N_1505,N_824);
nand U1989 (N_1989,N_1739,N_1616);
nand U1990 (N_1990,N_1288,N_673);
xor U1991 (N_1991,In_566,N_1439);
nand U1992 (N_1992,N_1259,N_1415);
nand U1993 (N_1993,N_1461,N_1403);
xor U1994 (N_1994,N_1448,N_467);
xnor U1995 (N_1995,N_1401,N_1679);
nor U1996 (N_1996,In_2352,N_187);
xor U1997 (N_1997,In_1695,N_423);
xnor U1998 (N_1998,In_49,N_828);
and U1999 (N_1999,N_1630,In_387);
xor U2000 (N_2000,N_1346,N_1907);
xor U2001 (N_2001,N_1970,N_1976);
and U2002 (N_2002,N_1789,N_1433);
xor U2003 (N_2003,N_1913,N_1840);
nand U2004 (N_2004,N_1982,N_1952);
nor U2005 (N_2005,N_1801,N_522);
xnor U2006 (N_2006,N_966,N_1246);
nor U2007 (N_2007,N_1615,N_1867);
nor U2008 (N_2008,N_1227,In_100);
or U2009 (N_2009,N_359,N_1766);
nand U2010 (N_2010,N_1363,N_1709);
and U2011 (N_2011,N_1872,N_1861);
nor U2012 (N_2012,N_1614,N_1879);
nand U2013 (N_2013,N_721,N_925);
xnor U2014 (N_2014,N_1566,N_1409);
nor U2015 (N_2015,N_1592,N_306);
nor U2016 (N_2016,N_1804,N_875);
xnor U2017 (N_2017,N_1299,In_810);
or U2018 (N_2018,N_1539,N_1934);
xor U2019 (N_2019,In_1929,In_457);
xor U2020 (N_2020,N_954,In_259);
nor U2021 (N_2021,N_1551,N_1985);
nand U2022 (N_2022,N_1807,N_1617);
and U2023 (N_2023,N_1847,N_1117);
nor U2024 (N_2024,N_1965,N_1528);
and U2025 (N_2025,N_1853,N_344);
nor U2026 (N_2026,N_1828,N_1799);
and U2027 (N_2027,N_471,N_1924);
or U2028 (N_2028,N_1663,N_1684);
nand U2029 (N_2029,N_1091,N_1802);
or U2030 (N_2030,N_383,N_1820);
or U2031 (N_2031,N_1555,N_372);
xor U2032 (N_2032,N_1518,N_1994);
or U2033 (N_2033,N_1134,N_670);
or U2034 (N_2034,N_1425,N_1623);
and U2035 (N_2035,N_1674,N_1821);
or U2036 (N_2036,In_860,N_1783);
nand U2037 (N_2037,N_1815,N_752);
xor U2038 (N_2038,N_1550,N_1277);
or U2039 (N_2039,N_1671,N_1335);
or U2040 (N_2040,N_1440,N_887);
or U2041 (N_2041,N_1110,N_1893);
xnor U2042 (N_2042,N_1079,N_1904);
nor U2043 (N_2043,In_108,In_1688);
and U2044 (N_2044,N_1631,In_2004);
and U2045 (N_2045,N_1882,In_689);
nand U2046 (N_2046,N_1977,N_46);
xor U2047 (N_2047,N_1854,N_1654);
and U2048 (N_2048,N_284,N_1400);
or U2049 (N_2049,N_1533,N_1812);
nor U2050 (N_2050,N_692,N_430);
and U2051 (N_2051,N_1928,N_1961);
and U2052 (N_2052,N_1967,N_1856);
or U2053 (N_2053,N_1758,N_1624);
nand U2054 (N_2054,N_1888,N_1130);
xnor U2055 (N_2055,N_1797,N_1969);
nor U2056 (N_2056,N_1978,N_930);
and U2057 (N_2057,N_1875,N_1729);
or U2058 (N_2058,N_1308,N_1757);
xnor U2059 (N_2059,N_1899,N_1921);
nand U2060 (N_2060,N_1619,N_1636);
xor U2061 (N_2061,N_1795,N_1587);
xnor U2062 (N_2062,N_1957,N_1627);
or U2063 (N_2063,N_1937,N_1819);
nor U2064 (N_2064,N_627,N_1792);
nor U2065 (N_2065,N_1843,N_1493);
and U2066 (N_2066,N_1609,N_1878);
nand U2067 (N_2067,In_1821,N_1207);
and U2068 (N_2068,N_1688,N_1125);
nor U2069 (N_2069,N_1837,In_425);
nand U2070 (N_2070,N_638,N_1895);
or U2071 (N_2071,N_1818,In_1824);
nand U2072 (N_2072,In_2241,N_496);
nor U2073 (N_2073,N_1827,In_1848);
or U2074 (N_2074,N_891,N_1876);
nor U2075 (N_2075,N_1269,N_1374);
and U2076 (N_2076,N_1889,N_1866);
xnor U2077 (N_2077,N_1778,N_1118);
or U2078 (N_2078,N_1637,In_2086);
nor U2079 (N_2079,N_1056,N_1701);
or U2080 (N_2080,In_467,N_787);
nand U2081 (N_2081,N_707,N_1955);
nor U2082 (N_2082,In_443,N_1940);
nor U2083 (N_2083,N_1554,N_1562);
nor U2084 (N_2084,N_1848,N_1883);
and U2085 (N_2085,N_447,N_1838);
nor U2086 (N_2086,N_1733,N_1813);
nor U2087 (N_2087,N_1917,N_1785);
xor U2088 (N_2088,N_1589,N_1537);
xnor U2089 (N_2089,N_1963,N_1980);
or U2090 (N_2090,N_1948,N_1722);
nor U2091 (N_2091,In_1914,N_34);
nor U2092 (N_2092,N_1752,N_1919);
xor U2093 (N_2093,N_1730,N_1911);
or U2094 (N_2094,In_1851,N_1504);
and U2095 (N_2095,N_1938,N_513);
nor U2096 (N_2096,N_1350,N_1870);
nand U2097 (N_2097,N_1912,N_1744);
and U2098 (N_2098,N_1902,N_1833);
xor U2099 (N_2099,N_1887,N_1481);
or U2100 (N_2100,N_1823,N_1831);
nor U2101 (N_2101,N_688,N_1796);
and U2102 (N_2102,N_1874,N_615);
and U2103 (N_2103,N_1628,N_1999);
or U2104 (N_2104,N_1845,N_859);
or U2105 (N_2105,N_1753,N_1909);
xor U2106 (N_2106,N_1990,N_1805);
nand U2107 (N_2107,N_955,N_1946);
xnor U2108 (N_2108,N_1520,N_1850);
xor U2109 (N_2109,N_1995,In_1943);
xor U2110 (N_2110,N_1488,N_1983);
or U2111 (N_2111,N_1478,N_1974);
nor U2112 (N_2112,N_1939,In_522);
nand U2113 (N_2113,N_1661,N_1522);
xnor U2114 (N_2114,In_358,N_1775);
nor U2115 (N_2115,N_1923,N_1457);
or U2116 (N_2116,N_1593,N_1787);
nor U2117 (N_2117,N_945,N_1926);
or U2118 (N_2118,N_1844,N_999);
nand U2119 (N_2119,N_1612,N_765);
and U2120 (N_2120,N_1915,N_1997);
xor U2121 (N_2121,N_1936,N_1900);
nand U2122 (N_2122,N_1903,In_403);
or U2123 (N_2123,N_1307,In_2371);
nor U2124 (N_2124,N_1127,N_1842);
xor U2125 (N_2125,N_1910,N_1318);
and U2126 (N_2126,N_1824,N_1774);
xnor U2127 (N_2127,N_1236,N_939);
and U2128 (N_2128,N_1972,N_1989);
xnor U2129 (N_2129,N_1993,N_1986);
and U2130 (N_2130,N_1871,N_1280);
and U2131 (N_2131,N_1906,N_1968);
nor U2132 (N_2132,N_1886,N_980);
and U2133 (N_2133,N_1951,N_1023);
xnor U2134 (N_2134,In_1438,N_1542);
xnor U2135 (N_2135,N_261,N_1712);
and U2136 (N_2136,N_1881,In_1870);
nor U2137 (N_2137,N_1489,N_1035);
or U2138 (N_2138,N_1800,N_1790);
xnor U2139 (N_2139,N_1973,N_1717);
nand U2140 (N_2140,N_1016,In_1408);
nand U2141 (N_2141,N_1862,N_1294);
or U2142 (N_2142,N_1959,N_1803);
or U2143 (N_2143,In_2385,N_1656);
or U2144 (N_2144,N_1884,N_1665);
xnor U2145 (N_2145,In_1514,In_2349);
or U2146 (N_2146,N_1897,N_1470);
xor U2147 (N_2147,N_1622,N_1177);
nand U2148 (N_2148,N_963,N_1991);
nand U2149 (N_2149,N_1485,N_1666);
or U2150 (N_2150,In_1063,In_1200);
xor U2151 (N_2151,N_246,N_1398);
nand U2152 (N_2152,N_1841,N_1395);
or U2153 (N_2153,N_797,N_1935);
xor U2154 (N_2154,N_1492,N_1981);
nor U2155 (N_2155,N_1432,N_977);
or U2156 (N_2156,N_1779,N_1817);
nor U2157 (N_2157,N_1063,N_426);
nor U2158 (N_2158,N_1498,N_1770);
xnor U2159 (N_2159,N_1570,N_1849);
nand U2160 (N_2160,N_1925,In_2262);
or U2161 (N_2161,N_1834,N_1998);
and U2162 (N_2162,N_1892,N_1038);
nor U2163 (N_2163,N_973,N_1771);
nor U2164 (N_2164,In_2295,N_1890);
or U2165 (N_2165,N_1442,N_1908);
nor U2166 (N_2166,N_1953,N_853);
nand U2167 (N_2167,N_1929,N_1806);
nor U2168 (N_2168,N_1421,N_919);
or U2169 (N_2169,N_1943,N_1865);
nand U2170 (N_2170,In_840,N_915);
xnor U2171 (N_2171,N_1296,N_1095);
nand U2172 (N_2172,N_1603,N_1916);
and U2173 (N_2173,N_1629,N_1962);
or U2174 (N_2174,N_1710,N_1808);
and U2175 (N_2175,N_1944,N_1764);
xnor U2176 (N_2176,In_857,N_1667);
nor U2177 (N_2177,N_1525,N_1675);
and U2178 (N_2178,N_1822,N_1635);
and U2179 (N_2179,N_1559,N_1932);
nand U2180 (N_2180,N_1941,N_1859);
and U2181 (N_2181,N_1992,N_1544);
nand U2182 (N_2182,In_1667,N_1933);
and U2183 (N_2183,N_1880,N_1703);
nand U2184 (N_2184,N_1988,N_1873);
nand U2185 (N_2185,N_1956,N_1898);
or U2186 (N_2186,N_1649,N_1846);
and U2187 (N_2187,N_1950,In_84);
or U2188 (N_2188,N_1914,N_1686);
xor U2189 (N_2189,N_1052,N_1140);
or U2190 (N_2190,N_1051,N_1958);
or U2191 (N_2191,N_1868,In_2182);
or U2192 (N_2192,In_2344,N_1966);
nor U2193 (N_2193,N_1145,N_1430);
or U2194 (N_2194,N_1814,N_1760);
or U2195 (N_2195,N_1869,N_1756);
nor U2196 (N_2196,In_2160,N_1971);
and U2197 (N_2197,N_1408,N_1920);
nand U2198 (N_2198,N_1816,N_1901);
and U2199 (N_2199,In_1503,N_1019);
xor U2200 (N_2200,N_1521,N_1954);
or U2201 (N_2201,N_1922,N_2147);
xor U2202 (N_2202,N_2066,N_2029);
or U2203 (N_2203,N_2043,N_2070);
or U2204 (N_2204,N_2013,N_2149);
nand U2205 (N_2205,N_1945,N_2188);
and U2206 (N_2206,N_1930,N_1960);
nor U2207 (N_2207,N_1692,N_2039);
or U2208 (N_2208,N_1809,N_2190);
nor U2209 (N_2209,In_182,N_2064);
nand U2210 (N_2210,N_1456,N_2040);
nor U2211 (N_2211,N_2067,N_1896);
xnor U2212 (N_2212,N_1855,N_1780);
nor U2213 (N_2213,N_2087,N_1700);
xnor U2214 (N_2214,N_2195,N_1586);
nor U2215 (N_2215,N_2152,N_2023);
or U2216 (N_2216,N_2176,N_2169);
nor U2217 (N_2217,N_1918,N_2093);
nor U2218 (N_2218,N_2091,N_2053);
and U2219 (N_2219,N_1942,N_808);
nand U2220 (N_2220,N_2133,N_2164);
nor U2221 (N_2221,In_935,N_1669);
nor U2222 (N_2222,N_2060,N_2128);
and U2223 (N_2223,N_2112,N_1839);
nor U2224 (N_2224,N_2055,In_555);
and U2225 (N_2225,N_2136,N_2015);
xor U2226 (N_2226,N_2009,N_2008);
nor U2227 (N_2227,N_2036,N_1836);
xnor U2228 (N_2228,N_2108,N_2031);
xor U2229 (N_2229,N_1852,N_2140);
and U2230 (N_2230,N_2062,N_2001);
xor U2231 (N_2231,N_277,N_1979);
nor U2232 (N_2232,N_1905,N_2012);
nor U2233 (N_2233,In_1971,N_1375);
or U2234 (N_2234,N_1996,N_1829);
or U2235 (N_2235,N_1987,N_1595);
and U2236 (N_2236,N_2090,N_2134);
nand U2237 (N_2237,N_2046,N_2111);
or U2238 (N_2238,N_2125,In_1424);
and U2239 (N_2239,N_2010,N_2172);
nor U2240 (N_2240,N_2170,N_2016);
or U2241 (N_2241,N_743,N_361);
or U2242 (N_2242,N_2160,N_2189);
nor U2243 (N_2243,N_2097,N_2000);
nor U2244 (N_2244,N_1964,N_2076);
or U2245 (N_2245,N_2127,N_1370);
nand U2246 (N_2246,N_2084,N_2116);
and U2247 (N_2247,N_1759,N_2022);
and U2248 (N_2248,N_2003,N_2014);
nor U2249 (N_2249,N_2044,N_1811);
nand U2250 (N_2250,N_2121,N_2194);
xnor U2251 (N_2251,N_2120,N_2032);
and U2252 (N_2252,N_2117,N_2114);
nand U2253 (N_2253,N_2148,N_1832);
nand U2254 (N_2254,N_2180,N_1698);
and U2255 (N_2255,N_2199,N_2107);
nand U2256 (N_2256,N_2085,N_1877);
or U2257 (N_2257,N_2021,In_2127);
xnor U2258 (N_2258,N_1719,N_2118);
xor U2259 (N_2259,N_2054,N_1851);
nand U2260 (N_2260,N_2030,N_2185);
and U2261 (N_2261,N_1931,In_1007);
nor U2262 (N_2262,In_2067,N_2119);
nor U2263 (N_2263,N_2028,N_2145);
nand U2264 (N_2264,N_2082,N_2146);
or U2265 (N_2265,N_1835,N_378);
nor U2266 (N_2266,N_2047,N_1860);
nand U2267 (N_2267,N_2178,N_2005);
xnor U2268 (N_2268,N_2153,N_2191);
xor U2269 (N_2269,N_2182,In_2163);
nor U2270 (N_2270,N_2196,N_2154);
xor U2271 (N_2271,N_2156,N_2072);
and U2272 (N_2272,N_2162,N_575);
nand U2273 (N_2273,N_2065,N_2109);
nor U2274 (N_2274,N_2025,N_2123);
nand U2275 (N_2275,N_1927,N_2006);
or U2276 (N_2276,N_2027,N_2035);
nor U2277 (N_2277,N_1825,N_1830);
nand U2278 (N_2278,N_2167,N_1894);
or U2279 (N_2279,N_1975,N_2129);
nor U2280 (N_2280,N_2168,N_2018);
and U2281 (N_2281,N_2088,N_2138);
and U2282 (N_2282,N_1810,N_2101);
or U2283 (N_2283,N_2096,N_2124);
nor U2284 (N_2284,N_2183,N_1693);
xor U2285 (N_2285,N_2057,N_2092);
and U2286 (N_2286,N_1406,N_2126);
and U2287 (N_2287,N_2137,N_239);
xor U2288 (N_2288,N_991,N_2115);
nand U2289 (N_2289,N_2131,N_448);
and U2290 (N_2290,N_912,N_2192);
and U2291 (N_2291,N_2144,N_2110);
or U2292 (N_2292,N_1857,N_1858);
and U2293 (N_2293,N_2049,N_1655);
and U2294 (N_2294,N_2155,N_1427);
and U2295 (N_2295,N_1659,N_2163);
nand U2296 (N_2296,N_2059,N_2068);
xnor U2297 (N_2297,N_746,N_2037);
nor U2298 (N_2298,N_1776,N_2017);
and U2299 (N_2299,In_2096,N_2019);
nor U2300 (N_2300,N_292,N_2041);
xnor U2301 (N_2301,N_2158,N_2103);
or U2302 (N_2302,N_850,In_1724);
and U2303 (N_2303,N_2151,N_2089);
or U2304 (N_2304,N_1608,N_1602);
or U2305 (N_2305,N_2034,N_2038);
or U2306 (N_2306,N_2081,N_2052);
nor U2307 (N_2307,N_2105,N_2102);
nand U2308 (N_2308,N_1947,N_2045);
nand U2309 (N_2309,N_2132,N_2026);
nor U2310 (N_2310,N_2173,N_2078);
and U2311 (N_2311,N_2157,N_2020);
or U2312 (N_2312,N_2080,N_2174);
or U2313 (N_2313,N_2056,N_2179);
and U2314 (N_2314,N_2161,N_2061);
nand U2315 (N_2315,N_2069,N_2193);
and U2316 (N_2316,N_2033,N_2142);
or U2317 (N_2317,N_2171,N_2175);
nand U2318 (N_2318,N_2048,N_2079);
xor U2319 (N_2319,N_1761,N_1509);
nor U2320 (N_2320,N_1660,N_1885);
nor U2321 (N_2321,N_2098,N_2075);
nand U2322 (N_2322,N_2074,N_2004);
nor U2323 (N_2323,In_1755,N_1707);
and U2324 (N_2324,N_2106,N_2197);
xor U2325 (N_2325,N_1826,N_1206);
nand U2326 (N_2326,N_1984,N_2077);
xnor U2327 (N_2327,N_2143,N_2095);
nand U2328 (N_2328,In_460,N_1891);
nor U2329 (N_2329,N_2104,N_2058);
nand U2330 (N_2330,N_2086,N_2094);
or U2331 (N_2331,N_2099,N_1714);
or U2332 (N_2332,N_2073,N_67);
or U2333 (N_2333,N_1724,N_2100);
or U2334 (N_2334,N_2002,N_2051);
or U2335 (N_2335,N_2050,N_1864);
and U2336 (N_2336,N_2135,N_2007);
nor U2337 (N_2337,N_2083,N_1718);
xnor U2338 (N_2338,N_2139,N_2042);
or U2339 (N_2339,N_2159,N_2186);
and U2340 (N_2340,N_2187,N_2166);
xnor U2341 (N_2341,N_2063,N_2184);
nor U2342 (N_2342,N_2150,N_2198);
xor U2343 (N_2343,N_1949,N_2165);
nand U2344 (N_2344,N_2011,N_1763);
or U2345 (N_2345,N_2141,N_1863);
nand U2346 (N_2346,N_2122,N_2024);
nand U2347 (N_2347,N_2177,N_2113);
or U2348 (N_2348,N_2181,N_2071);
and U2349 (N_2349,N_2130,N_1556);
nor U2350 (N_2350,N_1891,In_2096);
xor U2351 (N_2351,N_2018,N_2032);
and U2352 (N_2352,N_1714,N_2124);
nand U2353 (N_2353,N_2138,N_2118);
nand U2354 (N_2354,N_2047,N_1918);
nand U2355 (N_2355,N_2017,N_2085);
xor U2356 (N_2356,N_991,N_2073);
nor U2357 (N_2357,N_2052,N_2173);
xor U2358 (N_2358,N_2088,N_2065);
or U2359 (N_2359,N_575,N_2038);
or U2360 (N_2360,N_2190,N_2114);
nor U2361 (N_2361,N_1949,N_2045);
xor U2362 (N_2362,N_2147,N_2009);
xnor U2363 (N_2363,N_2183,N_2083);
and U2364 (N_2364,N_1839,N_2037);
or U2365 (N_2365,N_1698,N_1987);
and U2366 (N_2366,N_2018,N_2160);
nand U2367 (N_2367,N_1996,N_1863);
nand U2368 (N_2368,N_1714,N_1602);
and U2369 (N_2369,N_2006,N_2084);
or U2370 (N_2370,N_1718,N_1905);
nand U2371 (N_2371,N_1918,N_1945);
nor U2372 (N_2372,N_2007,N_2114);
xnor U2373 (N_2373,N_2076,N_2013);
and U2374 (N_2374,N_1829,N_1811);
xor U2375 (N_2375,N_2073,N_2043);
and U2376 (N_2376,N_2150,N_67);
and U2377 (N_2377,N_2062,N_808);
nor U2378 (N_2378,N_2173,N_1836);
nand U2379 (N_2379,N_2082,N_1693);
and U2380 (N_2380,N_1810,N_2111);
nand U2381 (N_2381,N_1945,N_277);
nor U2382 (N_2382,N_1698,N_1660);
nand U2383 (N_2383,N_2134,N_1693);
and U2384 (N_2384,N_2013,N_2178);
and U2385 (N_2385,N_2065,N_2053);
nand U2386 (N_2386,N_2138,N_1655);
or U2387 (N_2387,N_1698,N_2132);
and U2388 (N_2388,N_2111,N_2078);
and U2389 (N_2389,N_2074,N_2048);
xor U2390 (N_2390,N_2175,N_1964);
nor U2391 (N_2391,N_2100,N_2047);
and U2392 (N_2392,N_1855,N_2164);
xor U2393 (N_2393,N_2063,N_2149);
or U2394 (N_2394,N_2192,N_1669);
nor U2395 (N_2395,N_1669,N_1942);
and U2396 (N_2396,N_2005,N_2047);
and U2397 (N_2397,N_1931,N_2051);
nand U2398 (N_2398,N_2079,In_2067);
or U2399 (N_2399,N_2132,N_991);
nand U2400 (N_2400,N_2301,N_2322);
xor U2401 (N_2401,N_2367,N_2318);
nand U2402 (N_2402,N_2268,N_2285);
nor U2403 (N_2403,N_2382,N_2284);
xor U2404 (N_2404,N_2329,N_2361);
nor U2405 (N_2405,N_2257,N_2327);
or U2406 (N_2406,N_2369,N_2388);
and U2407 (N_2407,N_2358,N_2229);
and U2408 (N_2408,N_2221,N_2295);
nor U2409 (N_2409,N_2220,N_2364);
and U2410 (N_2410,N_2212,N_2302);
and U2411 (N_2411,N_2359,N_2308);
xor U2412 (N_2412,N_2218,N_2278);
xor U2413 (N_2413,N_2243,N_2303);
or U2414 (N_2414,N_2219,N_2215);
nand U2415 (N_2415,N_2351,N_2231);
nand U2416 (N_2416,N_2255,N_2336);
xor U2417 (N_2417,N_2227,N_2337);
nand U2418 (N_2418,N_2270,N_2385);
or U2419 (N_2419,N_2383,N_2201);
xor U2420 (N_2420,N_2312,N_2390);
nand U2421 (N_2421,N_2360,N_2250);
nor U2422 (N_2422,N_2328,N_2381);
or U2423 (N_2423,N_2348,N_2291);
nand U2424 (N_2424,N_2280,N_2211);
nor U2425 (N_2425,N_2392,N_2246);
or U2426 (N_2426,N_2300,N_2306);
nor U2427 (N_2427,N_2209,N_2232);
and U2428 (N_2428,N_2290,N_2325);
xnor U2429 (N_2429,N_2352,N_2240);
xor U2430 (N_2430,N_2281,N_2237);
and U2431 (N_2431,N_2338,N_2279);
xor U2432 (N_2432,N_2368,N_2216);
nand U2433 (N_2433,N_2354,N_2323);
and U2434 (N_2434,N_2294,N_2223);
nor U2435 (N_2435,N_2331,N_2272);
and U2436 (N_2436,N_2316,N_2292);
nor U2437 (N_2437,N_2313,N_2355);
nor U2438 (N_2438,N_2253,N_2203);
or U2439 (N_2439,N_2241,N_2320);
nand U2440 (N_2440,N_2311,N_2345);
or U2441 (N_2441,N_2299,N_2200);
nand U2442 (N_2442,N_2375,N_2349);
and U2443 (N_2443,N_2235,N_2386);
xor U2444 (N_2444,N_2252,N_2373);
nand U2445 (N_2445,N_2234,N_2233);
or U2446 (N_2446,N_2384,N_2387);
and U2447 (N_2447,N_2261,N_2370);
nor U2448 (N_2448,N_2330,N_2248);
nor U2449 (N_2449,N_2244,N_2260);
nor U2450 (N_2450,N_2335,N_2228);
or U2451 (N_2451,N_2210,N_2339);
nor U2452 (N_2452,N_2366,N_2242);
or U2453 (N_2453,N_2286,N_2350);
xor U2454 (N_2454,N_2399,N_2282);
nand U2455 (N_2455,N_2276,N_2363);
nand U2456 (N_2456,N_2379,N_2283);
nand U2457 (N_2457,N_2309,N_2332);
nor U2458 (N_2458,N_2256,N_2317);
nand U2459 (N_2459,N_2374,N_2347);
xor U2460 (N_2460,N_2397,N_2346);
nor U2461 (N_2461,N_2205,N_2362);
or U2462 (N_2462,N_2398,N_2289);
xor U2463 (N_2463,N_2371,N_2258);
nor U2464 (N_2464,N_2344,N_2343);
or U2465 (N_2465,N_2307,N_2263);
nand U2466 (N_2466,N_2396,N_2377);
nand U2467 (N_2467,N_2224,N_2380);
nand U2468 (N_2468,N_2230,N_2245);
nand U2469 (N_2469,N_2225,N_2378);
xor U2470 (N_2470,N_2391,N_2395);
or U2471 (N_2471,N_2259,N_2251);
nand U2472 (N_2472,N_2319,N_2334);
nor U2473 (N_2473,N_2277,N_2202);
or U2474 (N_2474,N_2266,N_2342);
and U2475 (N_2475,N_2236,N_2324);
or U2476 (N_2476,N_2265,N_2267);
xor U2477 (N_2477,N_2274,N_2271);
or U2478 (N_2478,N_2287,N_2326);
nor U2479 (N_2479,N_2222,N_2365);
nor U2480 (N_2480,N_2314,N_2247);
nand U2481 (N_2481,N_2340,N_2296);
nor U2482 (N_2482,N_2288,N_2341);
or U2483 (N_2483,N_2254,N_2305);
or U2484 (N_2484,N_2394,N_2213);
and U2485 (N_2485,N_2206,N_2269);
nor U2486 (N_2486,N_2204,N_2264);
or U2487 (N_2487,N_2217,N_2273);
nor U2488 (N_2488,N_2321,N_2353);
nand U2489 (N_2489,N_2226,N_2298);
nor U2490 (N_2490,N_2356,N_2238);
nand U2491 (N_2491,N_2357,N_2372);
nor U2492 (N_2492,N_2389,N_2333);
nor U2493 (N_2493,N_2208,N_2275);
nand U2494 (N_2494,N_2297,N_2304);
and U2495 (N_2495,N_2214,N_2376);
xor U2496 (N_2496,N_2262,N_2249);
xnor U2497 (N_2497,N_2310,N_2207);
or U2498 (N_2498,N_2293,N_2239);
and U2499 (N_2499,N_2393,N_2315);
nand U2500 (N_2500,N_2225,N_2344);
xor U2501 (N_2501,N_2270,N_2274);
xor U2502 (N_2502,N_2365,N_2344);
or U2503 (N_2503,N_2282,N_2331);
nor U2504 (N_2504,N_2342,N_2242);
or U2505 (N_2505,N_2316,N_2301);
nor U2506 (N_2506,N_2301,N_2365);
xor U2507 (N_2507,N_2324,N_2329);
nand U2508 (N_2508,N_2354,N_2340);
xnor U2509 (N_2509,N_2260,N_2308);
nor U2510 (N_2510,N_2289,N_2269);
xor U2511 (N_2511,N_2293,N_2302);
and U2512 (N_2512,N_2381,N_2215);
nor U2513 (N_2513,N_2250,N_2367);
nand U2514 (N_2514,N_2282,N_2266);
nand U2515 (N_2515,N_2222,N_2275);
nor U2516 (N_2516,N_2307,N_2361);
or U2517 (N_2517,N_2382,N_2220);
xnor U2518 (N_2518,N_2254,N_2297);
nand U2519 (N_2519,N_2292,N_2237);
xor U2520 (N_2520,N_2311,N_2226);
or U2521 (N_2521,N_2207,N_2204);
nor U2522 (N_2522,N_2316,N_2385);
xor U2523 (N_2523,N_2225,N_2246);
nor U2524 (N_2524,N_2391,N_2255);
nand U2525 (N_2525,N_2320,N_2344);
xnor U2526 (N_2526,N_2350,N_2316);
xor U2527 (N_2527,N_2279,N_2315);
xnor U2528 (N_2528,N_2327,N_2232);
xnor U2529 (N_2529,N_2325,N_2227);
nor U2530 (N_2530,N_2242,N_2353);
nor U2531 (N_2531,N_2336,N_2366);
or U2532 (N_2532,N_2315,N_2299);
xor U2533 (N_2533,N_2204,N_2326);
nand U2534 (N_2534,N_2304,N_2359);
and U2535 (N_2535,N_2329,N_2328);
or U2536 (N_2536,N_2357,N_2283);
and U2537 (N_2537,N_2222,N_2358);
or U2538 (N_2538,N_2212,N_2244);
and U2539 (N_2539,N_2364,N_2345);
nand U2540 (N_2540,N_2337,N_2375);
xor U2541 (N_2541,N_2321,N_2370);
and U2542 (N_2542,N_2389,N_2259);
xor U2543 (N_2543,N_2391,N_2376);
xor U2544 (N_2544,N_2355,N_2212);
nor U2545 (N_2545,N_2287,N_2240);
nor U2546 (N_2546,N_2219,N_2387);
or U2547 (N_2547,N_2354,N_2277);
or U2548 (N_2548,N_2284,N_2378);
nor U2549 (N_2549,N_2387,N_2270);
or U2550 (N_2550,N_2227,N_2203);
nor U2551 (N_2551,N_2294,N_2305);
or U2552 (N_2552,N_2358,N_2397);
nand U2553 (N_2553,N_2202,N_2223);
nand U2554 (N_2554,N_2235,N_2350);
or U2555 (N_2555,N_2308,N_2303);
and U2556 (N_2556,N_2201,N_2257);
nand U2557 (N_2557,N_2220,N_2294);
or U2558 (N_2558,N_2279,N_2320);
and U2559 (N_2559,N_2324,N_2372);
xor U2560 (N_2560,N_2332,N_2352);
nand U2561 (N_2561,N_2209,N_2279);
or U2562 (N_2562,N_2391,N_2261);
or U2563 (N_2563,N_2316,N_2299);
nor U2564 (N_2564,N_2351,N_2360);
nor U2565 (N_2565,N_2255,N_2352);
nand U2566 (N_2566,N_2235,N_2249);
and U2567 (N_2567,N_2261,N_2274);
and U2568 (N_2568,N_2364,N_2315);
nand U2569 (N_2569,N_2295,N_2325);
nand U2570 (N_2570,N_2379,N_2320);
nand U2571 (N_2571,N_2399,N_2369);
xnor U2572 (N_2572,N_2269,N_2299);
xor U2573 (N_2573,N_2300,N_2393);
nand U2574 (N_2574,N_2213,N_2222);
and U2575 (N_2575,N_2292,N_2322);
nand U2576 (N_2576,N_2316,N_2357);
nor U2577 (N_2577,N_2382,N_2297);
xor U2578 (N_2578,N_2333,N_2268);
nand U2579 (N_2579,N_2384,N_2314);
or U2580 (N_2580,N_2298,N_2382);
nor U2581 (N_2581,N_2204,N_2371);
nand U2582 (N_2582,N_2362,N_2213);
and U2583 (N_2583,N_2384,N_2310);
or U2584 (N_2584,N_2399,N_2308);
xnor U2585 (N_2585,N_2325,N_2367);
nand U2586 (N_2586,N_2229,N_2301);
nand U2587 (N_2587,N_2344,N_2324);
and U2588 (N_2588,N_2342,N_2391);
nor U2589 (N_2589,N_2206,N_2371);
and U2590 (N_2590,N_2291,N_2208);
nand U2591 (N_2591,N_2297,N_2316);
nor U2592 (N_2592,N_2222,N_2265);
nor U2593 (N_2593,N_2286,N_2243);
xor U2594 (N_2594,N_2387,N_2221);
xor U2595 (N_2595,N_2226,N_2334);
nand U2596 (N_2596,N_2249,N_2244);
or U2597 (N_2597,N_2260,N_2306);
nor U2598 (N_2598,N_2380,N_2282);
nand U2599 (N_2599,N_2391,N_2208);
xor U2600 (N_2600,N_2579,N_2420);
and U2601 (N_2601,N_2416,N_2500);
or U2602 (N_2602,N_2550,N_2488);
or U2603 (N_2603,N_2576,N_2408);
xor U2604 (N_2604,N_2495,N_2545);
xor U2605 (N_2605,N_2563,N_2448);
or U2606 (N_2606,N_2570,N_2566);
xnor U2607 (N_2607,N_2546,N_2454);
or U2608 (N_2608,N_2511,N_2478);
or U2609 (N_2609,N_2443,N_2598);
nor U2610 (N_2610,N_2498,N_2431);
xnor U2611 (N_2611,N_2444,N_2562);
or U2612 (N_2612,N_2527,N_2531);
or U2613 (N_2613,N_2410,N_2421);
and U2614 (N_2614,N_2536,N_2465);
nand U2615 (N_2615,N_2560,N_2440);
or U2616 (N_2616,N_2475,N_2542);
nand U2617 (N_2617,N_2569,N_2459);
and U2618 (N_2618,N_2481,N_2510);
xor U2619 (N_2619,N_2442,N_2424);
nand U2620 (N_2620,N_2505,N_2464);
xor U2621 (N_2621,N_2552,N_2514);
nor U2622 (N_2622,N_2447,N_2412);
xnor U2623 (N_2623,N_2512,N_2494);
nor U2624 (N_2624,N_2470,N_2457);
and U2625 (N_2625,N_2476,N_2596);
and U2626 (N_2626,N_2513,N_2521);
or U2627 (N_2627,N_2438,N_2485);
xnor U2628 (N_2628,N_2599,N_2544);
xor U2629 (N_2629,N_2532,N_2526);
nor U2630 (N_2630,N_2497,N_2473);
xor U2631 (N_2631,N_2418,N_2586);
and U2632 (N_2632,N_2499,N_2583);
xnor U2633 (N_2633,N_2434,N_2429);
xnor U2634 (N_2634,N_2503,N_2458);
nor U2635 (N_2635,N_2558,N_2589);
xnor U2636 (N_2636,N_2535,N_2415);
or U2637 (N_2637,N_2491,N_2405);
nand U2638 (N_2638,N_2538,N_2486);
and U2639 (N_2639,N_2400,N_2460);
nor U2640 (N_2640,N_2539,N_2413);
xor U2641 (N_2641,N_2439,N_2582);
xnor U2642 (N_2642,N_2561,N_2591);
and U2643 (N_2643,N_2441,N_2557);
and U2644 (N_2644,N_2466,N_2572);
nand U2645 (N_2645,N_2575,N_2452);
or U2646 (N_2646,N_2493,N_2568);
xnor U2647 (N_2647,N_2468,N_2422);
xor U2648 (N_2648,N_2437,N_2594);
nor U2649 (N_2649,N_2461,N_2588);
or U2650 (N_2650,N_2414,N_2403);
nand U2651 (N_2651,N_2419,N_2553);
nor U2652 (N_2652,N_2502,N_2487);
xor U2653 (N_2653,N_2573,N_2404);
xor U2654 (N_2654,N_2507,N_2492);
or U2655 (N_2655,N_2449,N_2411);
and U2656 (N_2656,N_2559,N_2428);
nand U2657 (N_2657,N_2590,N_2520);
nand U2658 (N_2658,N_2471,N_2541);
nor U2659 (N_2659,N_2417,N_2474);
or U2660 (N_2660,N_2462,N_2504);
nand U2661 (N_2661,N_2480,N_2581);
nor U2662 (N_2662,N_2402,N_2477);
and U2663 (N_2663,N_2515,N_2584);
nor U2664 (N_2664,N_2516,N_2451);
and U2665 (N_2665,N_2525,N_2574);
xor U2666 (N_2666,N_2446,N_2528);
and U2667 (N_2667,N_2472,N_2489);
xor U2668 (N_2668,N_2592,N_2463);
or U2669 (N_2669,N_2537,N_2483);
xnor U2670 (N_2670,N_2540,N_2554);
xnor U2671 (N_2671,N_2567,N_2436);
or U2672 (N_2672,N_2469,N_2533);
xor U2673 (N_2673,N_2467,N_2490);
nor U2674 (N_2674,N_2509,N_2564);
xnor U2675 (N_2675,N_2423,N_2522);
nor U2676 (N_2676,N_2530,N_2547);
or U2677 (N_2677,N_2430,N_2585);
xor U2678 (N_2678,N_2455,N_2593);
or U2679 (N_2679,N_2409,N_2549);
xnor U2680 (N_2680,N_2506,N_2496);
xnor U2681 (N_2681,N_2565,N_2450);
xor U2682 (N_2682,N_2578,N_2534);
xnor U2683 (N_2683,N_2484,N_2426);
xnor U2684 (N_2684,N_2456,N_2580);
and U2685 (N_2685,N_2548,N_2524);
nor U2686 (N_2686,N_2433,N_2501);
or U2687 (N_2687,N_2543,N_2435);
or U2688 (N_2688,N_2482,N_2529);
or U2689 (N_2689,N_2508,N_2427);
nor U2690 (N_2690,N_2406,N_2517);
nand U2691 (N_2691,N_2597,N_2479);
nand U2692 (N_2692,N_2401,N_2556);
nand U2693 (N_2693,N_2407,N_2577);
xor U2694 (N_2694,N_2555,N_2432);
nor U2695 (N_2695,N_2453,N_2518);
nor U2696 (N_2696,N_2523,N_2587);
xnor U2697 (N_2697,N_2425,N_2445);
and U2698 (N_2698,N_2551,N_2571);
nand U2699 (N_2699,N_2595,N_2519);
and U2700 (N_2700,N_2580,N_2406);
and U2701 (N_2701,N_2447,N_2451);
xor U2702 (N_2702,N_2414,N_2503);
nand U2703 (N_2703,N_2507,N_2575);
nand U2704 (N_2704,N_2458,N_2424);
or U2705 (N_2705,N_2553,N_2555);
nand U2706 (N_2706,N_2591,N_2453);
nor U2707 (N_2707,N_2452,N_2506);
and U2708 (N_2708,N_2486,N_2549);
or U2709 (N_2709,N_2447,N_2426);
or U2710 (N_2710,N_2555,N_2599);
and U2711 (N_2711,N_2514,N_2449);
nand U2712 (N_2712,N_2497,N_2490);
and U2713 (N_2713,N_2442,N_2483);
or U2714 (N_2714,N_2471,N_2509);
nand U2715 (N_2715,N_2493,N_2546);
nand U2716 (N_2716,N_2449,N_2571);
or U2717 (N_2717,N_2502,N_2469);
nand U2718 (N_2718,N_2407,N_2565);
and U2719 (N_2719,N_2580,N_2527);
nor U2720 (N_2720,N_2547,N_2582);
and U2721 (N_2721,N_2539,N_2517);
nand U2722 (N_2722,N_2463,N_2536);
or U2723 (N_2723,N_2426,N_2510);
xnor U2724 (N_2724,N_2571,N_2564);
or U2725 (N_2725,N_2537,N_2564);
nor U2726 (N_2726,N_2511,N_2451);
nand U2727 (N_2727,N_2447,N_2545);
nand U2728 (N_2728,N_2546,N_2589);
xor U2729 (N_2729,N_2501,N_2544);
nor U2730 (N_2730,N_2401,N_2525);
and U2731 (N_2731,N_2526,N_2516);
xor U2732 (N_2732,N_2522,N_2490);
nor U2733 (N_2733,N_2547,N_2448);
nand U2734 (N_2734,N_2593,N_2543);
xnor U2735 (N_2735,N_2497,N_2427);
xor U2736 (N_2736,N_2468,N_2417);
nand U2737 (N_2737,N_2554,N_2489);
xnor U2738 (N_2738,N_2526,N_2522);
xnor U2739 (N_2739,N_2528,N_2511);
nor U2740 (N_2740,N_2462,N_2589);
xor U2741 (N_2741,N_2577,N_2411);
or U2742 (N_2742,N_2538,N_2590);
and U2743 (N_2743,N_2572,N_2541);
nand U2744 (N_2744,N_2596,N_2460);
nand U2745 (N_2745,N_2411,N_2403);
nor U2746 (N_2746,N_2552,N_2448);
nor U2747 (N_2747,N_2468,N_2597);
or U2748 (N_2748,N_2428,N_2456);
nand U2749 (N_2749,N_2497,N_2478);
or U2750 (N_2750,N_2459,N_2494);
and U2751 (N_2751,N_2504,N_2463);
xnor U2752 (N_2752,N_2403,N_2447);
nand U2753 (N_2753,N_2505,N_2446);
xnor U2754 (N_2754,N_2565,N_2502);
nand U2755 (N_2755,N_2465,N_2533);
xnor U2756 (N_2756,N_2481,N_2504);
xor U2757 (N_2757,N_2550,N_2577);
nor U2758 (N_2758,N_2455,N_2432);
nor U2759 (N_2759,N_2537,N_2555);
nand U2760 (N_2760,N_2485,N_2530);
and U2761 (N_2761,N_2447,N_2433);
nand U2762 (N_2762,N_2571,N_2440);
and U2763 (N_2763,N_2464,N_2524);
nand U2764 (N_2764,N_2533,N_2579);
nand U2765 (N_2765,N_2569,N_2410);
nor U2766 (N_2766,N_2447,N_2476);
xnor U2767 (N_2767,N_2456,N_2467);
or U2768 (N_2768,N_2482,N_2560);
nand U2769 (N_2769,N_2573,N_2514);
or U2770 (N_2770,N_2562,N_2471);
and U2771 (N_2771,N_2475,N_2461);
nand U2772 (N_2772,N_2528,N_2465);
xor U2773 (N_2773,N_2583,N_2467);
or U2774 (N_2774,N_2514,N_2437);
nand U2775 (N_2775,N_2413,N_2563);
or U2776 (N_2776,N_2512,N_2450);
xor U2777 (N_2777,N_2536,N_2486);
and U2778 (N_2778,N_2502,N_2547);
or U2779 (N_2779,N_2493,N_2582);
nand U2780 (N_2780,N_2551,N_2490);
and U2781 (N_2781,N_2552,N_2451);
or U2782 (N_2782,N_2516,N_2599);
nor U2783 (N_2783,N_2405,N_2432);
and U2784 (N_2784,N_2593,N_2594);
xor U2785 (N_2785,N_2530,N_2523);
and U2786 (N_2786,N_2425,N_2435);
and U2787 (N_2787,N_2441,N_2526);
or U2788 (N_2788,N_2420,N_2505);
xnor U2789 (N_2789,N_2433,N_2559);
nor U2790 (N_2790,N_2579,N_2480);
nor U2791 (N_2791,N_2474,N_2562);
nand U2792 (N_2792,N_2482,N_2406);
and U2793 (N_2793,N_2599,N_2584);
xor U2794 (N_2794,N_2492,N_2552);
and U2795 (N_2795,N_2564,N_2451);
or U2796 (N_2796,N_2484,N_2577);
or U2797 (N_2797,N_2573,N_2554);
nand U2798 (N_2798,N_2438,N_2414);
xnor U2799 (N_2799,N_2552,N_2543);
or U2800 (N_2800,N_2709,N_2730);
or U2801 (N_2801,N_2600,N_2795);
nand U2802 (N_2802,N_2640,N_2710);
nand U2803 (N_2803,N_2720,N_2706);
xnor U2804 (N_2804,N_2743,N_2663);
or U2805 (N_2805,N_2642,N_2660);
nand U2806 (N_2806,N_2708,N_2638);
nand U2807 (N_2807,N_2656,N_2613);
and U2808 (N_2808,N_2687,N_2618);
nor U2809 (N_2809,N_2764,N_2672);
nor U2810 (N_2810,N_2679,N_2609);
or U2811 (N_2811,N_2702,N_2723);
xnor U2812 (N_2812,N_2741,N_2665);
or U2813 (N_2813,N_2655,N_2694);
nor U2814 (N_2814,N_2681,N_2667);
and U2815 (N_2815,N_2787,N_2608);
and U2816 (N_2816,N_2767,N_2654);
nor U2817 (N_2817,N_2649,N_2751);
nor U2818 (N_2818,N_2629,N_2680);
nor U2819 (N_2819,N_2716,N_2639);
nor U2820 (N_2820,N_2612,N_2688);
or U2821 (N_2821,N_2653,N_2610);
nand U2822 (N_2822,N_2760,N_2664);
and U2823 (N_2823,N_2651,N_2605);
or U2824 (N_2824,N_2633,N_2701);
and U2825 (N_2825,N_2631,N_2792);
xnor U2826 (N_2826,N_2602,N_2722);
xnor U2827 (N_2827,N_2746,N_2735);
and U2828 (N_2828,N_2673,N_2771);
nand U2829 (N_2829,N_2732,N_2617);
or U2830 (N_2830,N_2601,N_2703);
nand U2831 (N_2831,N_2791,N_2781);
nor U2832 (N_2832,N_2750,N_2621);
nand U2833 (N_2833,N_2603,N_2700);
nand U2834 (N_2834,N_2630,N_2677);
and U2835 (N_2835,N_2784,N_2676);
or U2836 (N_2836,N_2776,N_2614);
or U2837 (N_2837,N_2740,N_2756);
nor U2838 (N_2838,N_2765,N_2736);
nand U2839 (N_2839,N_2668,N_2738);
and U2840 (N_2840,N_2749,N_2674);
xor U2841 (N_2841,N_2684,N_2786);
nand U2842 (N_2842,N_2699,N_2733);
nor U2843 (N_2843,N_2695,N_2691);
nor U2844 (N_2844,N_2758,N_2755);
and U2845 (N_2845,N_2692,N_2753);
nand U2846 (N_2846,N_2624,N_2775);
nand U2847 (N_2847,N_2626,N_2693);
xor U2848 (N_2848,N_2652,N_2777);
nor U2849 (N_2849,N_2628,N_2761);
or U2850 (N_2850,N_2705,N_2728);
nand U2851 (N_2851,N_2662,N_2782);
or U2852 (N_2852,N_2607,N_2635);
nand U2853 (N_2853,N_2774,N_2697);
or U2854 (N_2854,N_2714,N_2657);
or U2855 (N_2855,N_2637,N_2698);
nor U2856 (N_2856,N_2683,N_2647);
and U2857 (N_2857,N_2779,N_2606);
or U2858 (N_2858,N_2788,N_2686);
or U2859 (N_2859,N_2796,N_2616);
nand U2860 (N_2860,N_2650,N_2744);
or U2861 (N_2861,N_2696,N_2757);
and U2862 (N_2862,N_2772,N_2636);
nor U2863 (N_2863,N_2658,N_2718);
xnor U2864 (N_2864,N_2724,N_2754);
or U2865 (N_2865,N_2646,N_2678);
xnor U2866 (N_2866,N_2762,N_2797);
or U2867 (N_2867,N_2799,N_2778);
xnor U2868 (N_2868,N_2721,N_2645);
nand U2869 (N_2869,N_2625,N_2666);
nor U2870 (N_2870,N_2766,N_2622);
or U2871 (N_2871,N_2670,N_2682);
nand U2872 (N_2872,N_2644,N_2717);
nand U2873 (N_2873,N_2742,N_2671);
xnor U2874 (N_2874,N_2737,N_2620);
nand U2875 (N_2875,N_2727,N_2739);
nand U2876 (N_2876,N_2769,N_2759);
nor U2877 (N_2877,N_2627,N_2611);
or U2878 (N_2878,N_2752,N_2748);
xor U2879 (N_2879,N_2615,N_2719);
and U2880 (N_2880,N_2734,N_2785);
or U2881 (N_2881,N_2729,N_2675);
and U2882 (N_2882,N_2713,N_2789);
or U2883 (N_2883,N_2659,N_2768);
or U2884 (N_2884,N_2623,N_2798);
or U2885 (N_2885,N_2690,N_2661);
xor U2886 (N_2886,N_2689,N_2726);
xnor U2887 (N_2887,N_2643,N_2783);
and U2888 (N_2888,N_2715,N_2634);
xnor U2889 (N_2889,N_2619,N_2794);
nand U2890 (N_2890,N_2770,N_2707);
and U2891 (N_2891,N_2648,N_2793);
and U2892 (N_2892,N_2725,N_2704);
xnor U2893 (N_2893,N_2669,N_2712);
nand U2894 (N_2894,N_2604,N_2685);
xor U2895 (N_2895,N_2747,N_2641);
nor U2896 (N_2896,N_2745,N_2773);
or U2897 (N_2897,N_2763,N_2711);
or U2898 (N_2898,N_2632,N_2790);
xnor U2899 (N_2899,N_2780,N_2731);
and U2900 (N_2900,N_2712,N_2731);
and U2901 (N_2901,N_2634,N_2694);
or U2902 (N_2902,N_2704,N_2611);
nand U2903 (N_2903,N_2780,N_2611);
and U2904 (N_2904,N_2777,N_2651);
nand U2905 (N_2905,N_2721,N_2726);
nand U2906 (N_2906,N_2627,N_2690);
nor U2907 (N_2907,N_2685,N_2696);
xnor U2908 (N_2908,N_2618,N_2614);
and U2909 (N_2909,N_2731,N_2699);
xor U2910 (N_2910,N_2719,N_2714);
and U2911 (N_2911,N_2769,N_2735);
and U2912 (N_2912,N_2617,N_2621);
nor U2913 (N_2913,N_2620,N_2732);
or U2914 (N_2914,N_2776,N_2754);
or U2915 (N_2915,N_2770,N_2680);
nand U2916 (N_2916,N_2613,N_2653);
nand U2917 (N_2917,N_2734,N_2687);
nand U2918 (N_2918,N_2741,N_2727);
nor U2919 (N_2919,N_2706,N_2766);
nor U2920 (N_2920,N_2751,N_2604);
xnor U2921 (N_2921,N_2738,N_2649);
xor U2922 (N_2922,N_2762,N_2672);
or U2923 (N_2923,N_2623,N_2794);
or U2924 (N_2924,N_2752,N_2636);
or U2925 (N_2925,N_2618,N_2774);
and U2926 (N_2926,N_2601,N_2627);
nand U2927 (N_2927,N_2740,N_2674);
or U2928 (N_2928,N_2642,N_2773);
nor U2929 (N_2929,N_2791,N_2620);
nor U2930 (N_2930,N_2797,N_2638);
xor U2931 (N_2931,N_2697,N_2733);
nand U2932 (N_2932,N_2606,N_2665);
nor U2933 (N_2933,N_2781,N_2768);
nand U2934 (N_2934,N_2755,N_2730);
nor U2935 (N_2935,N_2623,N_2631);
xor U2936 (N_2936,N_2688,N_2669);
or U2937 (N_2937,N_2734,N_2744);
xor U2938 (N_2938,N_2661,N_2618);
and U2939 (N_2939,N_2646,N_2741);
xor U2940 (N_2940,N_2665,N_2767);
nand U2941 (N_2941,N_2642,N_2760);
and U2942 (N_2942,N_2795,N_2648);
nand U2943 (N_2943,N_2612,N_2652);
or U2944 (N_2944,N_2715,N_2793);
and U2945 (N_2945,N_2719,N_2711);
xor U2946 (N_2946,N_2610,N_2646);
nor U2947 (N_2947,N_2681,N_2728);
nand U2948 (N_2948,N_2748,N_2757);
or U2949 (N_2949,N_2698,N_2752);
nand U2950 (N_2950,N_2707,N_2754);
and U2951 (N_2951,N_2623,N_2601);
nand U2952 (N_2952,N_2610,N_2741);
nand U2953 (N_2953,N_2674,N_2692);
nand U2954 (N_2954,N_2752,N_2635);
nand U2955 (N_2955,N_2608,N_2689);
nor U2956 (N_2956,N_2726,N_2729);
and U2957 (N_2957,N_2725,N_2791);
or U2958 (N_2958,N_2647,N_2717);
nor U2959 (N_2959,N_2653,N_2651);
or U2960 (N_2960,N_2628,N_2717);
or U2961 (N_2961,N_2794,N_2673);
nand U2962 (N_2962,N_2645,N_2683);
and U2963 (N_2963,N_2772,N_2631);
nor U2964 (N_2964,N_2745,N_2747);
nor U2965 (N_2965,N_2766,N_2725);
nor U2966 (N_2966,N_2696,N_2674);
nor U2967 (N_2967,N_2738,N_2774);
and U2968 (N_2968,N_2672,N_2698);
nand U2969 (N_2969,N_2797,N_2714);
xnor U2970 (N_2970,N_2786,N_2627);
nand U2971 (N_2971,N_2694,N_2798);
xor U2972 (N_2972,N_2636,N_2729);
nand U2973 (N_2973,N_2773,N_2717);
and U2974 (N_2974,N_2781,N_2636);
nand U2975 (N_2975,N_2658,N_2652);
nand U2976 (N_2976,N_2734,N_2789);
nor U2977 (N_2977,N_2792,N_2731);
nor U2978 (N_2978,N_2616,N_2687);
nor U2979 (N_2979,N_2697,N_2644);
and U2980 (N_2980,N_2646,N_2767);
or U2981 (N_2981,N_2631,N_2688);
nand U2982 (N_2982,N_2758,N_2609);
and U2983 (N_2983,N_2697,N_2735);
nand U2984 (N_2984,N_2779,N_2693);
and U2985 (N_2985,N_2716,N_2761);
xor U2986 (N_2986,N_2761,N_2711);
nor U2987 (N_2987,N_2626,N_2637);
xor U2988 (N_2988,N_2729,N_2782);
nor U2989 (N_2989,N_2687,N_2648);
nor U2990 (N_2990,N_2733,N_2624);
nor U2991 (N_2991,N_2638,N_2636);
or U2992 (N_2992,N_2674,N_2787);
or U2993 (N_2993,N_2682,N_2751);
or U2994 (N_2994,N_2771,N_2603);
nand U2995 (N_2995,N_2660,N_2603);
nor U2996 (N_2996,N_2761,N_2668);
or U2997 (N_2997,N_2760,N_2647);
and U2998 (N_2998,N_2677,N_2650);
and U2999 (N_2999,N_2640,N_2798);
or U3000 (N_3000,N_2936,N_2924);
nand U3001 (N_3001,N_2855,N_2965);
or U3002 (N_3002,N_2926,N_2847);
or U3003 (N_3003,N_2892,N_2849);
or U3004 (N_3004,N_2872,N_2851);
nor U3005 (N_3005,N_2815,N_2972);
nor U3006 (N_3006,N_2943,N_2840);
nor U3007 (N_3007,N_2876,N_2956);
and U3008 (N_3008,N_2873,N_2859);
nand U3009 (N_3009,N_2935,N_2882);
xor U3010 (N_3010,N_2838,N_2853);
nor U3011 (N_3011,N_2867,N_2973);
or U3012 (N_3012,N_2940,N_2917);
nand U3013 (N_3013,N_2870,N_2928);
xor U3014 (N_3014,N_2919,N_2885);
nand U3015 (N_3015,N_2960,N_2832);
and U3016 (N_3016,N_2805,N_2897);
or U3017 (N_3017,N_2914,N_2978);
xor U3018 (N_3018,N_2858,N_2871);
or U3019 (N_3019,N_2845,N_2984);
nand U3020 (N_3020,N_2816,N_2986);
nor U3021 (N_3021,N_2823,N_2969);
nand U3022 (N_3022,N_2971,N_2977);
or U3023 (N_3023,N_2810,N_2861);
nand U3024 (N_3024,N_2902,N_2989);
or U3025 (N_3025,N_2980,N_2942);
or U3026 (N_3026,N_2983,N_2941);
nor U3027 (N_3027,N_2958,N_2888);
nor U3028 (N_3028,N_2938,N_2891);
or U3029 (N_3029,N_2925,N_2923);
and U3030 (N_3030,N_2846,N_2804);
nand U3031 (N_3031,N_2839,N_2822);
nand U3032 (N_3032,N_2985,N_2834);
nand U3033 (N_3033,N_2961,N_2887);
and U3034 (N_3034,N_2953,N_2821);
nor U3035 (N_3035,N_2968,N_2930);
nand U3036 (N_3036,N_2869,N_2814);
nand U3037 (N_3037,N_2826,N_2974);
or U3038 (N_3038,N_2912,N_2981);
nor U3039 (N_3039,N_2905,N_2893);
and U3040 (N_3040,N_2901,N_2857);
nand U3041 (N_3041,N_2955,N_2948);
and U3042 (N_3042,N_2835,N_2864);
nor U3043 (N_3043,N_2929,N_2895);
nand U3044 (N_3044,N_2812,N_2868);
nor U3045 (N_3045,N_2806,N_2931);
or U3046 (N_3046,N_2952,N_2987);
and U3047 (N_3047,N_2970,N_2988);
or U3048 (N_3048,N_2829,N_2903);
and U3049 (N_3049,N_2862,N_2811);
and U3050 (N_3050,N_2946,N_2802);
and U3051 (N_3051,N_2852,N_2848);
xnor U3052 (N_3052,N_2863,N_2904);
and U3053 (N_3053,N_2889,N_2913);
and U3054 (N_3054,N_2896,N_2801);
xnor U3055 (N_3055,N_2898,N_2837);
nor U3056 (N_3056,N_2937,N_2825);
nand U3057 (N_3057,N_2975,N_2877);
nand U3058 (N_3058,N_2828,N_2915);
and U3059 (N_3059,N_2865,N_2909);
or U3060 (N_3060,N_2827,N_2836);
and U3061 (N_3061,N_2963,N_2800);
nor U3062 (N_3062,N_2881,N_2933);
and U3063 (N_3063,N_2886,N_2949);
or U3064 (N_3064,N_2922,N_2967);
nor U3065 (N_3065,N_2939,N_2966);
and U3066 (N_3066,N_2920,N_2842);
or U3067 (N_3067,N_2951,N_2880);
or U3068 (N_3068,N_2944,N_2950);
and U3069 (N_3069,N_2996,N_2894);
nand U3070 (N_3070,N_2844,N_2900);
or U3071 (N_3071,N_2860,N_2957);
and U3072 (N_3072,N_2982,N_2959);
and U3073 (N_3073,N_2803,N_2879);
xnor U3074 (N_3074,N_2854,N_2830);
and U3075 (N_3075,N_2874,N_2856);
nor U3076 (N_3076,N_2875,N_2850);
nand U3077 (N_3077,N_2807,N_2866);
and U3078 (N_3078,N_2918,N_2831);
and U3079 (N_3079,N_2899,N_2908);
nand U3080 (N_3080,N_2820,N_2993);
xor U3081 (N_3081,N_2910,N_2964);
and U3082 (N_3082,N_2995,N_2884);
nor U3083 (N_3083,N_2841,N_2990);
nand U3084 (N_3084,N_2819,N_2997);
and U3085 (N_3085,N_2991,N_2947);
nor U3086 (N_3086,N_2883,N_2979);
nor U3087 (N_3087,N_2999,N_2934);
and U3088 (N_3088,N_2945,N_2907);
or U3089 (N_3089,N_2906,N_2813);
or U3090 (N_3090,N_2817,N_2808);
xnor U3091 (N_3091,N_2833,N_2998);
or U3092 (N_3092,N_2976,N_2916);
nand U3093 (N_3093,N_2911,N_2878);
or U3094 (N_3094,N_2927,N_2954);
or U3095 (N_3095,N_2992,N_2921);
or U3096 (N_3096,N_2843,N_2932);
nand U3097 (N_3097,N_2994,N_2890);
nor U3098 (N_3098,N_2824,N_2818);
nor U3099 (N_3099,N_2809,N_2962);
or U3100 (N_3100,N_2864,N_2991);
nand U3101 (N_3101,N_2947,N_2975);
and U3102 (N_3102,N_2994,N_2903);
nand U3103 (N_3103,N_2889,N_2941);
or U3104 (N_3104,N_2988,N_2813);
nor U3105 (N_3105,N_2856,N_2960);
or U3106 (N_3106,N_2911,N_2940);
nand U3107 (N_3107,N_2808,N_2819);
nand U3108 (N_3108,N_2850,N_2990);
nor U3109 (N_3109,N_2956,N_2982);
nor U3110 (N_3110,N_2913,N_2912);
and U3111 (N_3111,N_2896,N_2814);
nor U3112 (N_3112,N_2851,N_2943);
and U3113 (N_3113,N_2975,N_2892);
nor U3114 (N_3114,N_2806,N_2858);
or U3115 (N_3115,N_2879,N_2954);
xor U3116 (N_3116,N_2993,N_2913);
nor U3117 (N_3117,N_2913,N_2937);
nor U3118 (N_3118,N_2874,N_2919);
nand U3119 (N_3119,N_2814,N_2998);
xnor U3120 (N_3120,N_2925,N_2999);
nor U3121 (N_3121,N_2889,N_2926);
nor U3122 (N_3122,N_2838,N_2930);
nor U3123 (N_3123,N_2895,N_2956);
or U3124 (N_3124,N_2903,N_2932);
nor U3125 (N_3125,N_2893,N_2910);
xor U3126 (N_3126,N_2883,N_2899);
nor U3127 (N_3127,N_2878,N_2876);
xnor U3128 (N_3128,N_2981,N_2923);
nor U3129 (N_3129,N_2873,N_2803);
xnor U3130 (N_3130,N_2848,N_2887);
xor U3131 (N_3131,N_2912,N_2806);
or U3132 (N_3132,N_2942,N_2945);
and U3133 (N_3133,N_2854,N_2884);
nor U3134 (N_3134,N_2801,N_2853);
nand U3135 (N_3135,N_2972,N_2800);
nand U3136 (N_3136,N_2854,N_2820);
xnor U3137 (N_3137,N_2857,N_2859);
nor U3138 (N_3138,N_2973,N_2933);
or U3139 (N_3139,N_2888,N_2996);
xnor U3140 (N_3140,N_2818,N_2910);
nor U3141 (N_3141,N_2979,N_2815);
or U3142 (N_3142,N_2907,N_2825);
nor U3143 (N_3143,N_2883,N_2849);
nor U3144 (N_3144,N_2937,N_2920);
or U3145 (N_3145,N_2977,N_2934);
xor U3146 (N_3146,N_2874,N_2801);
or U3147 (N_3147,N_2866,N_2957);
xor U3148 (N_3148,N_2962,N_2969);
nand U3149 (N_3149,N_2835,N_2856);
or U3150 (N_3150,N_2833,N_2860);
nor U3151 (N_3151,N_2865,N_2903);
nand U3152 (N_3152,N_2992,N_2968);
or U3153 (N_3153,N_2817,N_2877);
xor U3154 (N_3154,N_2851,N_2934);
xnor U3155 (N_3155,N_2981,N_2861);
nand U3156 (N_3156,N_2841,N_2904);
or U3157 (N_3157,N_2868,N_2937);
or U3158 (N_3158,N_2885,N_2815);
and U3159 (N_3159,N_2903,N_2882);
xnor U3160 (N_3160,N_2944,N_2904);
nor U3161 (N_3161,N_2938,N_2858);
nand U3162 (N_3162,N_2924,N_2919);
nand U3163 (N_3163,N_2927,N_2882);
nor U3164 (N_3164,N_2839,N_2876);
nand U3165 (N_3165,N_2970,N_2900);
nor U3166 (N_3166,N_2934,N_2969);
and U3167 (N_3167,N_2808,N_2873);
and U3168 (N_3168,N_2922,N_2911);
and U3169 (N_3169,N_2987,N_2980);
nor U3170 (N_3170,N_2980,N_2840);
nor U3171 (N_3171,N_2889,N_2835);
or U3172 (N_3172,N_2928,N_2982);
and U3173 (N_3173,N_2859,N_2853);
nand U3174 (N_3174,N_2857,N_2910);
xor U3175 (N_3175,N_2814,N_2871);
nand U3176 (N_3176,N_2808,N_2890);
or U3177 (N_3177,N_2809,N_2987);
nand U3178 (N_3178,N_2890,N_2861);
and U3179 (N_3179,N_2854,N_2806);
or U3180 (N_3180,N_2899,N_2902);
xnor U3181 (N_3181,N_2938,N_2993);
and U3182 (N_3182,N_2956,N_2991);
nand U3183 (N_3183,N_2906,N_2948);
nand U3184 (N_3184,N_2818,N_2865);
xnor U3185 (N_3185,N_2974,N_2862);
nor U3186 (N_3186,N_2817,N_2973);
or U3187 (N_3187,N_2832,N_2857);
nand U3188 (N_3188,N_2813,N_2895);
nand U3189 (N_3189,N_2925,N_2858);
or U3190 (N_3190,N_2906,N_2812);
or U3191 (N_3191,N_2863,N_2925);
xnor U3192 (N_3192,N_2831,N_2969);
xnor U3193 (N_3193,N_2862,N_2869);
and U3194 (N_3194,N_2959,N_2936);
nor U3195 (N_3195,N_2924,N_2904);
or U3196 (N_3196,N_2810,N_2884);
and U3197 (N_3197,N_2833,N_2814);
nand U3198 (N_3198,N_2942,N_2918);
and U3199 (N_3199,N_2845,N_2926);
nor U3200 (N_3200,N_3094,N_3045);
nand U3201 (N_3201,N_3020,N_3176);
and U3202 (N_3202,N_3039,N_3129);
xor U3203 (N_3203,N_3044,N_3104);
nor U3204 (N_3204,N_3037,N_3025);
nand U3205 (N_3205,N_3142,N_3080);
and U3206 (N_3206,N_3156,N_3179);
nor U3207 (N_3207,N_3090,N_3101);
xor U3208 (N_3208,N_3026,N_3173);
nor U3209 (N_3209,N_3003,N_3127);
or U3210 (N_3210,N_3190,N_3145);
nor U3211 (N_3211,N_3116,N_3018);
nand U3212 (N_3212,N_3053,N_3136);
xnor U3213 (N_3213,N_3182,N_3089);
and U3214 (N_3214,N_3012,N_3151);
nor U3215 (N_3215,N_3185,N_3017);
and U3216 (N_3216,N_3123,N_3028);
nor U3217 (N_3217,N_3174,N_3060);
and U3218 (N_3218,N_3158,N_3032);
or U3219 (N_3219,N_3167,N_3029);
xnor U3220 (N_3220,N_3027,N_3059);
and U3221 (N_3221,N_3169,N_3024);
and U3222 (N_3222,N_3146,N_3057);
nor U3223 (N_3223,N_3047,N_3164);
nor U3224 (N_3224,N_3119,N_3010);
or U3225 (N_3225,N_3105,N_3198);
nor U3226 (N_3226,N_3196,N_3021);
xnor U3227 (N_3227,N_3188,N_3177);
or U3228 (N_3228,N_3184,N_3102);
nor U3229 (N_3229,N_3132,N_3191);
or U3230 (N_3230,N_3016,N_3052);
xor U3231 (N_3231,N_3110,N_3170);
nor U3232 (N_3232,N_3139,N_3118);
nor U3233 (N_3233,N_3068,N_3138);
and U3234 (N_3234,N_3048,N_3043);
xor U3235 (N_3235,N_3165,N_3075);
nor U3236 (N_3236,N_3124,N_3058);
and U3237 (N_3237,N_3178,N_3083);
xor U3238 (N_3238,N_3041,N_3125);
xnor U3239 (N_3239,N_3064,N_3065);
nor U3240 (N_3240,N_3042,N_3189);
nor U3241 (N_3241,N_3050,N_3088);
or U3242 (N_3242,N_3008,N_3107);
and U3243 (N_3243,N_3113,N_3171);
nor U3244 (N_3244,N_3040,N_3114);
xnor U3245 (N_3245,N_3091,N_3070);
and U3246 (N_3246,N_3128,N_3194);
nand U3247 (N_3247,N_3066,N_3056);
nand U3248 (N_3248,N_3001,N_3005);
or U3249 (N_3249,N_3115,N_3004);
and U3250 (N_3250,N_3038,N_3133);
and U3251 (N_3251,N_3061,N_3015);
nor U3252 (N_3252,N_3031,N_3134);
or U3253 (N_3253,N_3095,N_3109);
nor U3254 (N_3254,N_3081,N_3195);
xor U3255 (N_3255,N_3067,N_3168);
and U3256 (N_3256,N_3126,N_3199);
or U3257 (N_3257,N_3155,N_3160);
nand U3258 (N_3258,N_3006,N_3023);
and U3259 (N_3259,N_3175,N_3181);
xor U3260 (N_3260,N_3187,N_3096);
nand U3261 (N_3261,N_3072,N_3063);
nor U3262 (N_3262,N_3073,N_3186);
nand U3263 (N_3263,N_3051,N_3033);
xnor U3264 (N_3264,N_3130,N_3148);
or U3265 (N_3265,N_3092,N_3163);
or U3266 (N_3266,N_3055,N_3085);
nand U3267 (N_3267,N_3009,N_3117);
xor U3268 (N_3268,N_3131,N_3079);
nand U3269 (N_3269,N_3049,N_3087);
and U3270 (N_3270,N_3120,N_3152);
and U3271 (N_3271,N_3108,N_3019);
xnor U3272 (N_3272,N_3197,N_3098);
and U3273 (N_3273,N_3011,N_3022);
xnor U3274 (N_3274,N_3074,N_3084);
xnor U3275 (N_3275,N_3180,N_3007);
xnor U3276 (N_3276,N_3137,N_3121);
nand U3277 (N_3277,N_3099,N_3036);
nand U3278 (N_3278,N_3154,N_3112);
nand U3279 (N_3279,N_3013,N_3157);
xor U3280 (N_3280,N_3147,N_3111);
or U3281 (N_3281,N_3030,N_3172);
nor U3282 (N_3282,N_3035,N_3166);
or U3283 (N_3283,N_3192,N_3135);
nand U3284 (N_3284,N_3183,N_3162);
nand U3285 (N_3285,N_3122,N_3144);
nand U3286 (N_3286,N_3086,N_3034);
nor U3287 (N_3287,N_3150,N_3002);
and U3288 (N_3288,N_3103,N_3062);
or U3289 (N_3289,N_3161,N_3076);
xor U3290 (N_3290,N_3097,N_3141);
nand U3291 (N_3291,N_3106,N_3078);
and U3292 (N_3292,N_3071,N_3014);
nor U3293 (N_3293,N_3046,N_3153);
xnor U3294 (N_3294,N_3054,N_3000);
nor U3295 (N_3295,N_3143,N_3082);
xnor U3296 (N_3296,N_3149,N_3140);
nor U3297 (N_3297,N_3093,N_3159);
and U3298 (N_3298,N_3100,N_3077);
xor U3299 (N_3299,N_3193,N_3069);
xnor U3300 (N_3300,N_3013,N_3082);
nand U3301 (N_3301,N_3172,N_3142);
and U3302 (N_3302,N_3154,N_3050);
nand U3303 (N_3303,N_3196,N_3183);
nand U3304 (N_3304,N_3033,N_3050);
or U3305 (N_3305,N_3116,N_3068);
nor U3306 (N_3306,N_3006,N_3105);
nand U3307 (N_3307,N_3066,N_3015);
and U3308 (N_3308,N_3029,N_3009);
nand U3309 (N_3309,N_3151,N_3039);
nand U3310 (N_3310,N_3138,N_3019);
xor U3311 (N_3311,N_3110,N_3011);
nand U3312 (N_3312,N_3025,N_3164);
xnor U3313 (N_3313,N_3003,N_3096);
and U3314 (N_3314,N_3159,N_3172);
nand U3315 (N_3315,N_3058,N_3060);
or U3316 (N_3316,N_3095,N_3072);
xnor U3317 (N_3317,N_3052,N_3013);
nor U3318 (N_3318,N_3097,N_3023);
or U3319 (N_3319,N_3191,N_3012);
and U3320 (N_3320,N_3131,N_3003);
nand U3321 (N_3321,N_3008,N_3161);
and U3322 (N_3322,N_3094,N_3132);
or U3323 (N_3323,N_3051,N_3034);
nor U3324 (N_3324,N_3051,N_3077);
xnor U3325 (N_3325,N_3115,N_3139);
nand U3326 (N_3326,N_3017,N_3014);
and U3327 (N_3327,N_3009,N_3173);
xnor U3328 (N_3328,N_3095,N_3163);
and U3329 (N_3329,N_3021,N_3121);
xnor U3330 (N_3330,N_3144,N_3102);
or U3331 (N_3331,N_3116,N_3062);
nand U3332 (N_3332,N_3039,N_3025);
or U3333 (N_3333,N_3178,N_3054);
nand U3334 (N_3334,N_3052,N_3103);
nor U3335 (N_3335,N_3131,N_3078);
nand U3336 (N_3336,N_3179,N_3074);
nand U3337 (N_3337,N_3053,N_3198);
and U3338 (N_3338,N_3191,N_3022);
and U3339 (N_3339,N_3000,N_3033);
xnor U3340 (N_3340,N_3097,N_3011);
xnor U3341 (N_3341,N_3132,N_3150);
and U3342 (N_3342,N_3024,N_3105);
nand U3343 (N_3343,N_3046,N_3158);
xor U3344 (N_3344,N_3113,N_3178);
nor U3345 (N_3345,N_3098,N_3097);
nand U3346 (N_3346,N_3167,N_3101);
and U3347 (N_3347,N_3104,N_3004);
or U3348 (N_3348,N_3199,N_3075);
xnor U3349 (N_3349,N_3164,N_3024);
or U3350 (N_3350,N_3165,N_3071);
nor U3351 (N_3351,N_3082,N_3145);
xor U3352 (N_3352,N_3137,N_3141);
nand U3353 (N_3353,N_3066,N_3198);
xnor U3354 (N_3354,N_3059,N_3084);
nand U3355 (N_3355,N_3011,N_3019);
and U3356 (N_3356,N_3152,N_3121);
and U3357 (N_3357,N_3043,N_3195);
or U3358 (N_3358,N_3103,N_3077);
xnor U3359 (N_3359,N_3122,N_3163);
xnor U3360 (N_3360,N_3104,N_3120);
and U3361 (N_3361,N_3017,N_3106);
xor U3362 (N_3362,N_3193,N_3026);
or U3363 (N_3363,N_3067,N_3135);
nand U3364 (N_3364,N_3062,N_3104);
and U3365 (N_3365,N_3129,N_3122);
xnor U3366 (N_3366,N_3115,N_3193);
nand U3367 (N_3367,N_3130,N_3004);
or U3368 (N_3368,N_3198,N_3071);
or U3369 (N_3369,N_3119,N_3118);
and U3370 (N_3370,N_3059,N_3016);
xnor U3371 (N_3371,N_3138,N_3155);
or U3372 (N_3372,N_3070,N_3175);
nand U3373 (N_3373,N_3061,N_3170);
nor U3374 (N_3374,N_3099,N_3023);
or U3375 (N_3375,N_3071,N_3024);
or U3376 (N_3376,N_3015,N_3087);
xor U3377 (N_3377,N_3127,N_3194);
xor U3378 (N_3378,N_3054,N_3110);
nor U3379 (N_3379,N_3116,N_3064);
or U3380 (N_3380,N_3066,N_3108);
or U3381 (N_3381,N_3168,N_3179);
xnor U3382 (N_3382,N_3044,N_3125);
or U3383 (N_3383,N_3073,N_3041);
or U3384 (N_3384,N_3083,N_3139);
and U3385 (N_3385,N_3119,N_3077);
nor U3386 (N_3386,N_3088,N_3024);
or U3387 (N_3387,N_3155,N_3177);
and U3388 (N_3388,N_3080,N_3039);
or U3389 (N_3389,N_3096,N_3196);
xnor U3390 (N_3390,N_3088,N_3001);
or U3391 (N_3391,N_3069,N_3140);
xnor U3392 (N_3392,N_3042,N_3070);
or U3393 (N_3393,N_3186,N_3109);
xor U3394 (N_3394,N_3187,N_3006);
and U3395 (N_3395,N_3079,N_3051);
xor U3396 (N_3396,N_3115,N_3088);
or U3397 (N_3397,N_3111,N_3033);
and U3398 (N_3398,N_3180,N_3156);
nand U3399 (N_3399,N_3093,N_3193);
nor U3400 (N_3400,N_3392,N_3301);
xnor U3401 (N_3401,N_3313,N_3354);
nand U3402 (N_3402,N_3243,N_3275);
nand U3403 (N_3403,N_3399,N_3284);
xor U3404 (N_3404,N_3246,N_3346);
xnor U3405 (N_3405,N_3223,N_3388);
or U3406 (N_3406,N_3254,N_3222);
and U3407 (N_3407,N_3324,N_3326);
or U3408 (N_3408,N_3263,N_3287);
xor U3409 (N_3409,N_3380,N_3225);
or U3410 (N_3410,N_3274,N_3312);
nor U3411 (N_3411,N_3298,N_3360);
or U3412 (N_3412,N_3364,N_3356);
and U3413 (N_3413,N_3201,N_3337);
xnor U3414 (N_3414,N_3377,N_3396);
or U3415 (N_3415,N_3256,N_3299);
or U3416 (N_3416,N_3216,N_3357);
or U3417 (N_3417,N_3343,N_3260);
nand U3418 (N_3418,N_3276,N_3368);
nor U3419 (N_3419,N_3234,N_3257);
or U3420 (N_3420,N_3255,N_3304);
and U3421 (N_3421,N_3252,N_3332);
nand U3422 (N_3422,N_3373,N_3219);
nand U3423 (N_3423,N_3325,N_3242);
or U3424 (N_3424,N_3314,N_3232);
or U3425 (N_3425,N_3310,N_3353);
xor U3426 (N_3426,N_3347,N_3221);
or U3427 (N_3427,N_3361,N_3316);
xnor U3428 (N_3428,N_3387,N_3250);
nand U3429 (N_3429,N_3210,N_3266);
or U3430 (N_3430,N_3344,N_3215);
nor U3431 (N_3431,N_3334,N_3339);
and U3432 (N_3432,N_3372,N_3345);
and U3433 (N_3433,N_3336,N_3283);
xnor U3434 (N_3434,N_3258,N_3394);
nor U3435 (N_3435,N_3262,N_3297);
and U3436 (N_3436,N_3385,N_3237);
nor U3437 (N_3437,N_3398,N_3386);
nor U3438 (N_3438,N_3350,N_3200);
nand U3439 (N_3439,N_3292,N_3281);
nand U3440 (N_3440,N_3300,N_3271);
and U3441 (N_3441,N_3329,N_3279);
xor U3442 (N_3442,N_3307,N_3319);
or U3443 (N_3443,N_3249,N_3291);
nand U3444 (N_3444,N_3247,N_3205);
and U3445 (N_3445,N_3236,N_3207);
or U3446 (N_3446,N_3395,N_3212);
nand U3447 (N_3447,N_3358,N_3251);
nor U3448 (N_3448,N_3342,N_3370);
nor U3449 (N_3449,N_3286,N_3327);
xor U3450 (N_3450,N_3366,N_3305);
xnor U3451 (N_3451,N_3230,N_3288);
or U3452 (N_3452,N_3245,N_3321);
nand U3453 (N_3453,N_3208,N_3290);
or U3454 (N_3454,N_3315,N_3265);
and U3455 (N_3455,N_3348,N_3331);
nand U3456 (N_3456,N_3390,N_3393);
and U3457 (N_3457,N_3362,N_3397);
or U3458 (N_3458,N_3235,N_3379);
and U3459 (N_3459,N_3204,N_3295);
and U3460 (N_3460,N_3311,N_3220);
nor U3461 (N_3461,N_3240,N_3277);
nand U3462 (N_3462,N_3338,N_3365);
or U3463 (N_3463,N_3268,N_3309);
and U3464 (N_3464,N_3209,N_3228);
and U3465 (N_3465,N_3293,N_3203);
and U3466 (N_3466,N_3318,N_3226);
xnor U3467 (N_3467,N_3369,N_3273);
or U3468 (N_3468,N_3375,N_3389);
nand U3469 (N_3469,N_3359,N_3306);
or U3470 (N_3470,N_3302,N_3383);
nor U3471 (N_3471,N_3206,N_3248);
nand U3472 (N_3472,N_3378,N_3280);
nor U3473 (N_3473,N_3296,N_3322);
nor U3474 (N_3474,N_3355,N_3269);
nor U3475 (N_3475,N_3239,N_3374);
and U3476 (N_3476,N_3285,N_3328);
and U3477 (N_3477,N_3253,N_3340);
nand U3478 (N_3478,N_3224,N_3282);
and U3479 (N_3479,N_3233,N_3381);
nand U3480 (N_3480,N_3211,N_3391);
nand U3481 (N_3481,N_3341,N_3363);
xor U3482 (N_3482,N_3229,N_3382);
xor U3483 (N_3483,N_3376,N_3323);
nor U3484 (N_3484,N_3227,N_3294);
and U3485 (N_3485,N_3333,N_3267);
or U3486 (N_3486,N_3330,N_3238);
nand U3487 (N_3487,N_3371,N_3351);
nor U3488 (N_3488,N_3241,N_3349);
and U3489 (N_3489,N_3218,N_3289);
nand U3490 (N_3490,N_3278,N_3384);
xnor U3491 (N_3491,N_3264,N_3261);
and U3492 (N_3492,N_3317,N_3272);
nand U3493 (N_3493,N_3367,N_3308);
nor U3494 (N_3494,N_3202,N_3213);
or U3495 (N_3495,N_3259,N_3320);
and U3496 (N_3496,N_3270,N_3231);
xor U3497 (N_3497,N_3214,N_3303);
nor U3498 (N_3498,N_3244,N_3352);
and U3499 (N_3499,N_3217,N_3335);
and U3500 (N_3500,N_3373,N_3354);
and U3501 (N_3501,N_3268,N_3380);
nor U3502 (N_3502,N_3281,N_3352);
nor U3503 (N_3503,N_3277,N_3356);
nor U3504 (N_3504,N_3244,N_3387);
nor U3505 (N_3505,N_3329,N_3350);
or U3506 (N_3506,N_3326,N_3355);
nor U3507 (N_3507,N_3310,N_3234);
nand U3508 (N_3508,N_3264,N_3356);
or U3509 (N_3509,N_3268,N_3314);
nor U3510 (N_3510,N_3263,N_3364);
xor U3511 (N_3511,N_3374,N_3327);
nor U3512 (N_3512,N_3216,N_3254);
nand U3513 (N_3513,N_3341,N_3319);
nand U3514 (N_3514,N_3272,N_3283);
nand U3515 (N_3515,N_3356,N_3271);
and U3516 (N_3516,N_3201,N_3356);
nand U3517 (N_3517,N_3230,N_3317);
xnor U3518 (N_3518,N_3273,N_3348);
nor U3519 (N_3519,N_3239,N_3392);
nand U3520 (N_3520,N_3290,N_3298);
nor U3521 (N_3521,N_3337,N_3264);
nand U3522 (N_3522,N_3339,N_3390);
xnor U3523 (N_3523,N_3214,N_3224);
or U3524 (N_3524,N_3270,N_3384);
nand U3525 (N_3525,N_3335,N_3349);
or U3526 (N_3526,N_3265,N_3386);
or U3527 (N_3527,N_3269,N_3235);
nor U3528 (N_3528,N_3327,N_3277);
xnor U3529 (N_3529,N_3362,N_3316);
nand U3530 (N_3530,N_3283,N_3251);
nor U3531 (N_3531,N_3287,N_3245);
and U3532 (N_3532,N_3390,N_3258);
nor U3533 (N_3533,N_3283,N_3235);
xnor U3534 (N_3534,N_3285,N_3232);
or U3535 (N_3535,N_3358,N_3361);
nor U3536 (N_3536,N_3271,N_3204);
nor U3537 (N_3537,N_3371,N_3246);
nor U3538 (N_3538,N_3294,N_3272);
nor U3539 (N_3539,N_3370,N_3206);
or U3540 (N_3540,N_3291,N_3342);
and U3541 (N_3541,N_3370,N_3335);
and U3542 (N_3542,N_3250,N_3364);
nand U3543 (N_3543,N_3381,N_3300);
nor U3544 (N_3544,N_3338,N_3385);
nor U3545 (N_3545,N_3220,N_3308);
and U3546 (N_3546,N_3258,N_3290);
and U3547 (N_3547,N_3286,N_3392);
xnor U3548 (N_3548,N_3346,N_3224);
and U3549 (N_3549,N_3364,N_3214);
xor U3550 (N_3550,N_3222,N_3286);
and U3551 (N_3551,N_3358,N_3310);
or U3552 (N_3552,N_3210,N_3256);
nand U3553 (N_3553,N_3229,N_3396);
and U3554 (N_3554,N_3212,N_3274);
xor U3555 (N_3555,N_3272,N_3376);
and U3556 (N_3556,N_3216,N_3388);
or U3557 (N_3557,N_3247,N_3295);
xnor U3558 (N_3558,N_3317,N_3211);
and U3559 (N_3559,N_3344,N_3246);
nor U3560 (N_3560,N_3300,N_3328);
xor U3561 (N_3561,N_3284,N_3246);
nor U3562 (N_3562,N_3395,N_3337);
or U3563 (N_3563,N_3267,N_3223);
nor U3564 (N_3564,N_3276,N_3304);
and U3565 (N_3565,N_3296,N_3286);
and U3566 (N_3566,N_3376,N_3243);
nor U3567 (N_3567,N_3213,N_3316);
nor U3568 (N_3568,N_3256,N_3261);
nand U3569 (N_3569,N_3223,N_3279);
and U3570 (N_3570,N_3354,N_3203);
xor U3571 (N_3571,N_3279,N_3272);
nor U3572 (N_3572,N_3213,N_3243);
xor U3573 (N_3573,N_3325,N_3210);
or U3574 (N_3574,N_3274,N_3269);
and U3575 (N_3575,N_3313,N_3246);
nand U3576 (N_3576,N_3348,N_3300);
and U3577 (N_3577,N_3365,N_3354);
nand U3578 (N_3578,N_3273,N_3308);
and U3579 (N_3579,N_3273,N_3219);
xor U3580 (N_3580,N_3303,N_3249);
or U3581 (N_3581,N_3201,N_3236);
and U3582 (N_3582,N_3206,N_3382);
nor U3583 (N_3583,N_3230,N_3381);
xnor U3584 (N_3584,N_3236,N_3256);
xor U3585 (N_3585,N_3288,N_3249);
and U3586 (N_3586,N_3323,N_3226);
xnor U3587 (N_3587,N_3276,N_3236);
nor U3588 (N_3588,N_3212,N_3372);
xnor U3589 (N_3589,N_3224,N_3385);
and U3590 (N_3590,N_3204,N_3291);
xnor U3591 (N_3591,N_3280,N_3302);
nor U3592 (N_3592,N_3237,N_3362);
nor U3593 (N_3593,N_3222,N_3271);
or U3594 (N_3594,N_3366,N_3279);
and U3595 (N_3595,N_3355,N_3375);
or U3596 (N_3596,N_3326,N_3367);
nor U3597 (N_3597,N_3263,N_3321);
nor U3598 (N_3598,N_3296,N_3228);
nand U3599 (N_3599,N_3211,N_3281);
or U3600 (N_3600,N_3421,N_3535);
xor U3601 (N_3601,N_3453,N_3448);
or U3602 (N_3602,N_3574,N_3445);
or U3603 (N_3603,N_3438,N_3454);
and U3604 (N_3604,N_3499,N_3546);
and U3605 (N_3605,N_3404,N_3465);
xor U3606 (N_3606,N_3464,N_3447);
nor U3607 (N_3607,N_3418,N_3451);
nor U3608 (N_3608,N_3539,N_3512);
and U3609 (N_3609,N_3565,N_3538);
nand U3610 (N_3610,N_3416,N_3548);
xnor U3611 (N_3611,N_3575,N_3544);
xnor U3612 (N_3612,N_3550,N_3414);
nand U3613 (N_3613,N_3576,N_3431);
xor U3614 (N_3614,N_3588,N_3587);
xor U3615 (N_3615,N_3592,N_3527);
xor U3616 (N_3616,N_3547,N_3551);
nor U3617 (N_3617,N_3528,N_3481);
nor U3618 (N_3618,N_3505,N_3402);
nor U3619 (N_3619,N_3482,N_3472);
nor U3620 (N_3620,N_3428,N_3480);
xnor U3621 (N_3621,N_3516,N_3566);
and U3622 (N_3622,N_3496,N_3534);
nor U3623 (N_3623,N_3561,N_3443);
xnor U3624 (N_3624,N_3570,N_3522);
or U3625 (N_3625,N_3503,N_3412);
xnor U3626 (N_3626,N_3444,N_3523);
and U3627 (N_3627,N_3457,N_3526);
nor U3628 (N_3628,N_3476,N_3468);
xor U3629 (N_3629,N_3420,N_3426);
xor U3630 (N_3630,N_3563,N_3455);
nand U3631 (N_3631,N_3517,N_3510);
and U3632 (N_3632,N_3590,N_3578);
nor U3633 (N_3633,N_3558,N_3437);
xor U3634 (N_3634,N_3530,N_3586);
nand U3635 (N_3635,N_3489,N_3542);
and U3636 (N_3636,N_3459,N_3543);
and U3637 (N_3637,N_3525,N_3596);
nor U3638 (N_3638,N_3502,N_3411);
or U3639 (N_3639,N_3440,N_3524);
xnor U3640 (N_3640,N_3433,N_3436);
or U3641 (N_3641,N_3540,N_3462);
and U3642 (N_3642,N_3556,N_3573);
nand U3643 (N_3643,N_3442,N_3562);
xor U3644 (N_3644,N_3463,N_3456);
xor U3645 (N_3645,N_3408,N_3513);
nand U3646 (N_3646,N_3429,N_3449);
nand U3647 (N_3647,N_3553,N_3477);
nor U3648 (N_3648,N_3532,N_3531);
or U3649 (N_3649,N_3529,N_3520);
nor U3650 (N_3650,N_3419,N_3460);
xnor U3651 (N_3651,N_3434,N_3492);
nand U3652 (N_3652,N_3494,N_3580);
or U3653 (N_3653,N_3432,N_3500);
nand U3654 (N_3654,N_3484,N_3403);
or U3655 (N_3655,N_3490,N_3441);
or U3656 (N_3656,N_3508,N_3582);
nor U3657 (N_3657,N_3406,N_3518);
xor U3658 (N_3658,N_3568,N_3577);
and U3659 (N_3659,N_3461,N_3506);
nor U3660 (N_3660,N_3450,N_3452);
xnor U3661 (N_3661,N_3519,N_3415);
xnor U3662 (N_3662,N_3559,N_3473);
nand U3663 (N_3663,N_3599,N_3501);
and U3664 (N_3664,N_3409,N_3424);
or U3665 (N_3665,N_3598,N_3470);
xnor U3666 (N_3666,N_3511,N_3537);
nand U3667 (N_3667,N_3549,N_3583);
or U3668 (N_3668,N_3545,N_3521);
or U3669 (N_3669,N_3514,N_3491);
xor U3670 (N_3670,N_3446,N_3597);
nand U3671 (N_3671,N_3485,N_3479);
and U3672 (N_3672,N_3585,N_3555);
nand U3673 (N_3673,N_3483,N_3487);
and U3674 (N_3674,N_3486,N_3495);
nand U3675 (N_3675,N_3422,N_3423);
and U3676 (N_3676,N_3401,N_3541);
or U3677 (N_3677,N_3504,N_3571);
and U3678 (N_3678,N_3595,N_3413);
xor U3679 (N_3679,N_3410,N_3515);
or U3680 (N_3680,N_3435,N_3498);
nand U3681 (N_3681,N_3478,N_3430);
and U3682 (N_3682,N_3581,N_3557);
or U3683 (N_3683,N_3405,N_3474);
nor U3684 (N_3684,N_3488,N_3554);
nor U3685 (N_3685,N_3417,N_3509);
and U3686 (N_3686,N_3560,N_3469);
nand U3687 (N_3687,N_3572,N_3439);
nand U3688 (N_3688,N_3407,N_3569);
xnor U3689 (N_3689,N_3567,N_3427);
nor U3690 (N_3690,N_3475,N_3507);
nand U3691 (N_3691,N_3458,N_3471);
nor U3692 (N_3692,N_3579,N_3467);
nor U3693 (N_3693,N_3584,N_3400);
and U3694 (N_3694,N_3589,N_3564);
and U3695 (N_3695,N_3466,N_3425);
xor U3696 (N_3696,N_3497,N_3533);
or U3697 (N_3697,N_3493,N_3552);
xor U3698 (N_3698,N_3591,N_3536);
nand U3699 (N_3699,N_3594,N_3593);
nor U3700 (N_3700,N_3460,N_3411);
and U3701 (N_3701,N_3571,N_3525);
and U3702 (N_3702,N_3574,N_3438);
nor U3703 (N_3703,N_3540,N_3480);
nor U3704 (N_3704,N_3565,N_3475);
nor U3705 (N_3705,N_3440,N_3589);
xor U3706 (N_3706,N_3417,N_3444);
nor U3707 (N_3707,N_3596,N_3404);
or U3708 (N_3708,N_3479,N_3402);
nor U3709 (N_3709,N_3475,N_3576);
xor U3710 (N_3710,N_3510,N_3526);
or U3711 (N_3711,N_3546,N_3572);
nand U3712 (N_3712,N_3518,N_3438);
or U3713 (N_3713,N_3539,N_3401);
or U3714 (N_3714,N_3584,N_3423);
xor U3715 (N_3715,N_3598,N_3402);
or U3716 (N_3716,N_3407,N_3531);
and U3717 (N_3717,N_3458,N_3432);
or U3718 (N_3718,N_3433,N_3530);
nand U3719 (N_3719,N_3445,N_3517);
nor U3720 (N_3720,N_3421,N_3556);
xnor U3721 (N_3721,N_3499,N_3526);
nand U3722 (N_3722,N_3558,N_3511);
and U3723 (N_3723,N_3556,N_3554);
nand U3724 (N_3724,N_3476,N_3446);
or U3725 (N_3725,N_3457,N_3507);
nand U3726 (N_3726,N_3449,N_3453);
xor U3727 (N_3727,N_3454,N_3551);
nor U3728 (N_3728,N_3488,N_3407);
nand U3729 (N_3729,N_3564,N_3568);
nand U3730 (N_3730,N_3416,N_3570);
nand U3731 (N_3731,N_3436,N_3588);
and U3732 (N_3732,N_3534,N_3463);
xor U3733 (N_3733,N_3485,N_3460);
and U3734 (N_3734,N_3509,N_3506);
nand U3735 (N_3735,N_3545,N_3482);
nor U3736 (N_3736,N_3464,N_3492);
nand U3737 (N_3737,N_3474,N_3583);
nor U3738 (N_3738,N_3577,N_3529);
and U3739 (N_3739,N_3408,N_3478);
xnor U3740 (N_3740,N_3498,N_3436);
or U3741 (N_3741,N_3436,N_3583);
xnor U3742 (N_3742,N_3445,N_3499);
or U3743 (N_3743,N_3524,N_3496);
xnor U3744 (N_3744,N_3464,N_3428);
nor U3745 (N_3745,N_3467,N_3543);
and U3746 (N_3746,N_3426,N_3500);
and U3747 (N_3747,N_3479,N_3580);
nor U3748 (N_3748,N_3450,N_3504);
and U3749 (N_3749,N_3522,N_3502);
xor U3750 (N_3750,N_3482,N_3526);
xnor U3751 (N_3751,N_3480,N_3438);
nand U3752 (N_3752,N_3567,N_3598);
nor U3753 (N_3753,N_3476,N_3547);
or U3754 (N_3754,N_3485,N_3400);
and U3755 (N_3755,N_3587,N_3433);
or U3756 (N_3756,N_3556,N_3477);
xnor U3757 (N_3757,N_3404,N_3567);
or U3758 (N_3758,N_3524,N_3577);
nand U3759 (N_3759,N_3402,N_3514);
and U3760 (N_3760,N_3562,N_3527);
and U3761 (N_3761,N_3432,N_3553);
nor U3762 (N_3762,N_3437,N_3510);
xor U3763 (N_3763,N_3450,N_3448);
or U3764 (N_3764,N_3512,N_3573);
xnor U3765 (N_3765,N_3403,N_3499);
and U3766 (N_3766,N_3560,N_3499);
or U3767 (N_3767,N_3498,N_3507);
or U3768 (N_3768,N_3562,N_3539);
or U3769 (N_3769,N_3529,N_3564);
and U3770 (N_3770,N_3504,N_3418);
and U3771 (N_3771,N_3590,N_3489);
and U3772 (N_3772,N_3550,N_3582);
and U3773 (N_3773,N_3446,N_3431);
or U3774 (N_3774,N_3459,N_3540);
xnor U3775 (N_3775,N_3541,N_3571);
or U3776 (N_3776,N_3539,N_3411);
or U3777 (N_3777,N_3462,N_3465);
or U3778 (N_3778,N_3459,N_3553);
and U3779 (N_3779,N_3450,N_3530);
and U3780 (N_3780,N_3424,N_3566);
or U3781 (N_3781,N_3463,N_3510);
nand U3782 (N_3782,N_3458,N_3518);
xor U3783 (N_3783,N_3583,N_3547);
or U3784 (N_3784,N_3565,N_3463);
and U3785 (N_3785,N_3580,N_3573);
nor U3786 (N_3786,N_3424,N_3457);
or U3787 (N_3787,N_3585,N_3420);
or U3788 (N_3788,N_3416,N_3472);
xnor U3789 (N_3789,N_3461,N_3584);
or U3790 (N_3790,N_3587,N_3458);
or U3791 (N_3791,N_3599,N_3596);
or U3792 (N_3792,N_3494,N_3411);
and U3793 (N_3793,N_3478,N_3536);
nor U3794 (N_3794,N_3576,N_3553);
nor U3795 (N_3795,N_3402,N_3470);
or U3796 (N_3796,N_3418,N_3494);
and U3797 (N_3797,N_3590,N_3548);
and U3798 (N_3798,N_3410,N_3582);
nor U3799 (N_3799,N_3429,N_3484);
or U3800 (N_3800,N_3637,N_3731);
and U3801 (N_3801,N_3794,N_3750);
nor U3802 (N_3802,N_3614,N_3751);
or U3803 (N_3803,N_3603,N_3722);
or U3804 (N_3804,N_3640,N_3627);
xor U3805 (N_3805,N_3785,N_3678);
nand U3806 (N_3806,N_3708,N_3790);
xor U3807 (N_3807,N_3647,N_3703);
nand U3808 (N_3808,N_3729,N_3670);
and U3809 (N_3809,N_3756,N_3631);
nor U3810 (N_3810,N_3629,N_3623);
xnor U3811 (N_3811,N_3721,N_3795);
nor U3812 (N_3812,N_3768,N_3797);
nand U3813 (N_3813,N_3784,N_3778);
or U3814 (N_3814,N_3608,N_3674);
nor U3815 (N_3815,N_3607,N_3688);
nor U3816 (N_3816,N_3753,N_3713);
and U3817 (N_3817,N_3626,N_3747);
and U3818 (N_3818,N_3680,N_3605);
nor U3819 (N_3819,N_3745,N_3659);
and U3820 (N_3820,N_3711,N_3666);
or U3821 (N_3821,N_3651,N_3652);
xnor U3822 (N_3822,N_3662,N_3736);
or U3823 (N_3823,N_3763,N_3767);
xor U3824 (N_3824,N_3723,N_3739);
nand U3825 (N_3825,N_3672,N_3698);
nand U3826 (N_3826,N_3696,N_3775);
xnor U3827 (N_3827,N_3783,N_3625);
xnor U3828 (N_3828,N_3692,N_3633);
and U3829 (N_3829,N_3699,N_3611);
nor U3830 (N_3830,N_3655,N_3774);
nor U3831 (N_3831,N_3691,N_3653);
and U3832 (N_3832,N_3772,N_3606);
or U3833 (N_3833,N_3601,N_3733);
xor U3834 (N_3834,N_3788,N_3757);
nand U3835 (N_3835,N_3728,N_3689);
and U3836 (N_3836,N_3730,N_3748);
or U3837 (N_3837,N_3787,N_3665);
nand U3838 (N_3838,N_3707,N_3663);
and U3839 (N_3839,N_3761,N_3643);
and U3840 (N_3840,N_3619,N_3704);
nand U3841 (N_3841,N_3616,N_3693);
or U3842 (N_3842,N_3682,N_3724);
nand U3843 (N_3843,N_3744,N_3771);
and U3844 (N_3844,N_3781,N_3634);
and U3845 (N_3845,N_3675,N_3793);
or U3846 (N_3846,N_3654,N_3765);
nand U3847 (N_3847,N_3609,N_3648);
or U3848 (N_3848,N_3734,N_3701);
nand U3849 (N_3849,N_3610,N_3741);
and U3850 (N_3850,N_3749,N_3620);
or U3851 (N_3851,N_3667,N_3770);
xnor U3852 (N_3852,N_3746,N_3602);
nor U3853 (N_3853,N_3714,N_3628);
or U3854 (N_3854,N_3684,N_3687);
or U3855 (N_3855,N_3720,N_3638);
nand U3856 (N_3856,N_3740,N_3615);
nand U3857 (N_3857,N_3719,N_3681);
xnor U3858 (N_3858,N_3773,N_3786);
nor U3859 (N_3859,N_3726,N_3668);
nor U3860 (N_3860,N_3617,N_3646);
and U3861 (N_3861,N_3649,N_3718);
and U3862 (N_3862,N_3769,N_3776);
nor U3863 (N_3863,N_3759,N_3645);
xnor U3864 (N_3864,N_3683,N_3782);
and U3865 (N_3865,N_3697,N_3676);
nand U3866 (N_3866,N_3727,N_3712);
or U3867 (N_3867,N_3762,N_3660);
and U3868 (N_3868,N_3716,N_3622);
xor U3869 (N_3869,N_3789,N_3642);
xnor U3870 (N_3870,N_3661,N_3612);
and U3871 (N_3871,N_3679,N_3658);
xnor U3872 (N_3872,N_3657,N_3656);
or U3873 (N_3873,N_3780,N_3738);
nor U3874 (N_3874,N_3752,N_3702);
xnor U3875 (N_3875,N_3630,N_3735);
xor U3876 (N_3876,N_3624,N_3725);
or U3877 (N_3877,N_3777,N_3742);
nand U3878 (N_3878,N_3700,N_3621);
or U3879 (N_3879,N_3641,N_3760);
nand U3880 (N_3880,N_3639,N_3798);
nand U3881 (N_3881,N_3796,N_3710);
or U3882 (N_3882,N_3677,N_3737);
or U3883 (N_3883,N_3715,N_3799);
and U3884 (N_3884,N_3644,N_3618);
xnor U3885 (N_3885,N_3600,N_3709);
nand U3886 (N_3886,N_3705,N_3690);
nand U3887 (N_3887,N_3717,N_3695);
xnor U3888 (N_3888,N_3604,N_3686);
nor U3889 (N_3889,N_3635,N_3650);
nor U3890 (N_3890,N_3755,N_3779);
and U3891 (N_3891,N_3743,N_3673);
and U3892 (N_3892,N_3764,N_3732);
nor U3893 (N_3893,N_3685,N_3636);
nor U3894 (N_3894,N_3792,N_3664);
xor U3895 (N_3895,N_3754,N_3613);
xnor U3896 (N_3896,N_3791,N_3632);
nand U3897 (N_3897,N_3706,N_3694);
and U3898 (N_3898,N_3766,N_3671);
xnor U3899 (N_3899,N_3758,N_3669);
nor U3900 (N_3900,N_3705,N_3656);
xnor U3901 (N_3901,N_3711,N_3785);
and U3902 (N_3902,N_3625,N_3694);
and U3903 (N_3903,N_3795,N_3707);
xnor U3904 (N_3904,N_3709,N_3707);
and U3905 (N_3905,N_3661,N_3735);
nand U3906 (N_3906,N_3624,N_3721);
and U3907 (N_3907,N_3670,N_3769);
and U3908 (N_3908,N_3671,N_3780);
or U3909 (N_3909,N_3633,N_3622);
and U3910 (N_3910,N_3658,N_3716);
or U3911 (N_3911,N_3790,N_3794);
and U3912 (N_3912,N_3774,N_3784);
nor U3913 (N_3913,N_3678,N_3671);
or U3914 (N_3914,N_3780,N_3694);
nor U3915 (N_3915,N_3766,N_3764);
nor U3916 (N_3916,N_3752,N_3622);
xor U3917 (N_3917,N_3697,N_3777);
nand U3918 (N_3918,N_3610,N_3601);
and U3919 (N_3919,N_3635,N_3714);
xor U3920 (N_3920,N_3767,N_3624);
or U3921 (N_3921,N_3738,N_3769);
nand U3922 (N_3922,N_3683,N_3655);
xnor U3923 (N_3923,N_3625,N_3715);
nand U3924 (N_3924,N_3794,N_3696);
nor U3925 (N_3925,N_3611,N_3684);
nand U3926 (N_3926,N_3626,N_3675);
and U3927 (N_3927,N_3789,N_3716);
nor U3928 (N_3928,N_3675,N_3691);
or U3929 (N_3929,N_3791,N_3681);
nor U3930 (N_3930,N_3731,N_3671);
and U3931 (N_3931,N_3641,N_3785);
or U3932 (N_3932,N_3799,N_3604);
nand U3933 (N_3933,N_3644,N_3731);
and U3934 (N_3934,N_3774,N_3669);
nand U3935 (N_3935,N_3755,N_3638);
and U3936 (N_3936,N_3654,N_3705);
nand U3937 (N_3937,N_3602,N_3625);
or U3938 (N_3938,N_3700,N_3706);
or U3939 (N_3939,N_3647,N_3772);
or U3940 (N_3940,N_3616,N_3706);
or U3941 (N_3941,N_3673,N_3731);
nor U3942 (N_3942,N_3631,N_3677);
xnor U3943 (N_3943,N_3753,N_3631);
nor U3944 (N_3944,N_3792,N_3615);
xnor U3945 (N_3945,N_3769,N_3711);
and U3946 (N_3946,N_3611,N_3655);
nand U3947 (N_3947,N_3743,N_3767);
xor U3948 (N_3948,N_3775,N_3763);
nor U3949 (N_3949,N_3604,N_3693);
xnor U3950 (N_3950,N_3670,N_3754);
xnor U3951 (N_3951,N_3703,N_3786);
and U3952 (N_3952,N_3698,N_3727);
nor U3953 (N_3953,N_3761,N_3645);
or U3954 (N_3954,N_3768,N_3750);
or U3955 (N_3955,N_3658,N_3685);
xor U3956 (N_3956,N_3608,N_3758);
and U3957 (N_3957,N_3605,N_3769);
or U3958 (N_3958,N_3675,N_3775);
or U3959 (N_3959,N_3787,N_3607);
nor U3960 (N_3960,N_3685,N_3626);
xor U3961 (N_3961,N_3741,N_3697);
and U3962 (N_3962,N_3615,N_3605);
or U3963 (N_3963,N_3724,N_3646);
nor U3964 (N_3964,N_3662,N_3759);
xor U3965 (N_3965,N_3777,N_3770);
xor U3966 (N_3966,N_3631,N_3688);
xor U3967 (N_3967,N_3628,N_3698);
and U3968 (N_3968,N_3724,N_3680);
nor U3969 (N_3969,N_3623,N_3709);
xnor U3970 (N_3970,N_3730,N_3719);
nand U3971 (N_3971,N_3625,N_3646);
or U3972 (N_3972,N_3630,N_3751);
nor U3973 (N_3973,N_3651,N_3684);
nand U3974 (N_3974,N_3721,N_3739);
xnor U3975 (N_3975,N_3714,N_3702);
nor U3976 (N_3976,N_3684,N_3602);
nand U3977 (N_3977,N_3644,N_3791);
or U3978 (N_3978,N_3708,N_3770);
nand U3979 (N_3979,N_3671,N_3779);
nand U3980 (N_3980,N_3795,N_3754);
and U3981 (N_3981,N_3749,N_3799);
or U3982 (N_3982,N_3660,N_3766);
nand U3983 (N_3983,N_3730,N_3763);
nor U3984 (N_3984,N_3634,N_3619);
nand U3985 (N_3985,N_3792,N_3655);
xor U3986 (N_3986,N_3672,N_3640);
or U3987 (N_3987,N_3662,N_3718);
nor U3988 (N_3988,N_3670,N_3607);
nand U3989 (N_3989,N_3625,N_3632);
or U3990 (N_3990,N_3781,N_3733);
and U3991 (N_3991,N_3789,N_3611);
or U3992 (N_3992,N_3773,N_3732);
nor U3993 (N_3993,N_3763,N_3667);
nand U3994 (N_3994,N_3719,N_3699);
nor U3995 (N_3995,N_3717,N_3716);
or U3996 (N_3996,N_3608,N_3736);
xor U3997 (N_3997,N_3698,N_3784);
nor U3998 (N_3998,N_3759,N_3685);
nand U3999 (N_3999,N_3626,N_3650);
nor U4000 (N_4000,N_3903,N_3925);
or U4001 (N_4001,N_3956,N_3866);
xor U4002 (N_4002,N_3951,N_3842);
and U4003 (N_4003,N_3908,N_3970);
nor U4004 (N_4004,N_3806,N_3915);
nand U4005 (N_4005,N_3934,N_3942);
and U4006 (N_4006,N_3858,N_3909);
and U4007 (N_4007,N_3962,N_3884);
xnor U4008 (N_4008,N_3876,N_3801);
xor U4009 (N_4009,N_3862,N_3971);
xnor U4010 (N_4010,N_3999,N_3813);
xor U4011 (N_4011,N_3943,N_3821);
nand U4012 (N_4012,N_3985,N_3988);
or U4013 (N_4013,N_3958,N_3946);
or U4014 (N_4014,N_3857,N_3807);
and U4015 (N_4015,N_3919,N_3816);
nor U4016 (N_4016,N_3991,N_3901);
and U4017 (N_4017,N_3945,N_3871);
xor U4018 (N_4018,N_3984,N_3822);
and U4019 (N_4019,N_3923,N_3907);
xnor U4020 (N_4020,N_3826,N_3955);
or U4021 (N_4021,N_3891,N_3900);
nand U4022 (N_4022,N_3892,N_3817);
or U4023 (N_4023,N_3912,N_3815);
and U4024 (N_4024,N_3805,N_3830);
nand U4025 (N_4025,N_3895,N_3827);
and U4026 (N_4026,N_3808,N_3990);
nor U4027 (N_4027,N_3835,N_3917);
or U4028 (N_4028,N_3926,N_3910);
nand U4029 (N_4029,N_3935,N_3864);
and U4030 (N_4030,N_3982,N_3886);
and U4031 (N_4031,N_3930,N_3928);
nor U4032 (N_4032,N_3849,N_3885);
nor U4033 (N_4033,N_3836,N_3881);
nor U4034 (N_4034,N_3947,N_3809);
and U4035 (N_4035,N_3831,N_3996);
nand U4036 (N_4036,N_3922,N_3975);
and U4037 (N_4037,N_3965,N_3921);
nor U4038 (N_4038,N_3937,N_3837);
and U4039 (N_4039,N_3848,N_3877);
nor U4040 (N_4040,N_3887,N_3904);
or U4041 (N_4041,N_3967,N_3929);
or U4042 (N_4042,N_3841,N_3932);
or U4043 (N_4043,N_3861,N_3874);
nor U4044 (N_4044,N_3977,N_3939);
and U4045 (N_4045,N_3959,N_3924);
xor U4046 (N_4046,N_3963,N_3986);
xor U4047 (N_4047,N_3875,N_3823);
xnor U4048 (N_4048,N_3960,N_3879);
xnor U4049 (N_4049,N_3838,N_3993);
nand U4050 (N_4050,N_3964,N_3902);
and U4051 (N_4051,N_3979,N_3953);
and U4052 (N_4052,N_3914,N_3906);
and U4053 (N_4053,N_3843,N_3873);
or U4054 (N_4054,N_3957,N_3825);
xnor U4055 (N_4055,N_3810,N_3828);
xor U4056 (N_4056,N_3880,N_3983);
or U4057 (N_4057,N_3941,N_3832);
nor U4058 (N_4058,N_3819,N_3860);
nand U4059 (N_4059,N_3859,N_3868);
or U4060 (N_4060,N_3918,N_3865);
nor U4061 (N_4061,N_3883,N_3969);
nor U4062 (N_4062,N_3824,N_3829);
xnor U4063 (N_4063,N_3981,N_3995);
or U4064 (N_4064,N_3853,N_3952);
nor U4065 (N_4065,N_3994,N_3944);
xor U4066 (N_4066,N_3814,N_3893);
xnor U4067 (N_4067,N_3890,N_3927);
and U4068 (N_4068,N_3992,N_3998);
and U4069 (N_4069,N_3803,N_3851);
and U4070 (N_4070,N_3933,N_3936);
nor U4071 (N_4071,N_3978,N_3974);
and U4072 (N_4072,N_3938,N_3888);
nand U4073 (N_4073,N_3882,N_3954);
nand U4074 (N_4074,N_3863,N_3839);
or U4075 (N_4075,N_3976,N_3811);
and U4076 (N_4076,N_3812,N_3897);
and U4077 (N_4077,N_3961,N_3804);
or U4078 (N_4078,N_3972,N_3973);
and U4079 (N_4079,N_3916,N_3980);
xnor U4080 (N_4080,N_3949,N_3844);
nand U4081 (N_4081,N_3854,N_3852);
and U4082 (N_4082,N_3855,N_3931);
nor U4083 (N_4083,N_3889,N_3820);
nor U4084 (N_4084,N_3894,N_3850);
nand U4085 (N_4085,N_3940,N_3950);
xor U4086 (N_4086,N_3845,N_3847);
xor U4087 (N_4087,N_3920,N_3867);
nand U4088 (N_4088,N_3878,N_3899);
and U4089 (N_4089,N_3834,N_3833);
and U4090 (N_4090,N_3846,N_3856);
xnor U4091 (N_4091,N_3905,N_3896);
nand U4092 (N_4092,N_3872,N_3968);
nand U4093 (N_4093,N_3966,N_3911);
or U4094 (N_4094,N_3818,N_3869);
or U4095 (N_4095,N_3948,N_3989);
nor U4096 (N_4096,N_3800,N_3870);
xor U4097 (N_4097,N_3987,N_3802);
and U4098 (N_4098,N_3913,N_3840);
nand U4099 (N_4099,N_3898,N_3997);
nand U4100 (N_4100,N_3826,N_3943);
nor U4101 (N_4101,N_3994,N_3899);
nor U4102 (N_4102,N_3986,N_3953);
xor U4103 (N_4103,N_3917,N_3910);
or U4104 (N_4104,N_3827,N_3972);
xnor U4105 (N_4105,N_3955,N_3844);
nor U4106 (N_4106,N_3809,N_3948);
xor U4107 (N_4107,N_3889,N_3912);
and U4108 (N_4108,N_3816,N_3896);
nor U4109 (N_4109,N_3891,N_3943);
and U4110 (N_4110,N_3976,N_3893);
nand U4111 (N_4111,N_3829,N_3939);
or U4112 (N_4112,N_3850,N_3881);
nor U4113 (N_4113,N_3954,N_3895);
and U4114 (N_4114,N_3811,N_3923);
or U4115 (N_4115,N_3853,N_3974);
or U4116 (N_4116,N_3853,N_3877);
nand U4117 (N_4117,N_3952,N_3962);
or U4118 (N_4118,N_3909,N_3931);
nor U4119 (N_4119,N_3816,N_3990);
xnor U4120 (N_4120,N_3961,N_3949);
nand U4121 (N_4121,N_3871,N_3869);
or U4122 (N_4122,N_3837,N_3816);
xnor U4123 (N_4123,N_3803,N_3861);
nor U4124 (N_4124,N_3984,N_3921);
or U4125 (N_4125,N_3851,N_3966);
or U4126 (N_4126,N_3821,N_3985);
and U4127 (N_4127,N_3933,N_3881);
and U4128 (N_4128,N_3922,N_3911);
and U4129 (N_4129,N_3820,N_3870);
xnor U4130 (N_4130,N_3808,N_3898);
or U4131 (N_4131,N_3984,N_3931);
nand U4132 (N_4132,N_3850,N_3991);
xnor U4133 (N_4133,N_3802,N_3879);
nand U4134 (N_4134,N_3926,N_3990);
nand U4135 (N_4135,N_3820,N_3888);
nand U4136 (N_4136,N_3990,N_3851);
nand U4137 (N_4137,N_3929,N_3815);
xnor U4138 (N_4138,N_3972,N_3970);
xnor U4139 (N_4139,N_3865,N_3843);
and U4140 (N_4140,N_3817,N_3835);
nand U4141 (N_4141,N_3912,N_3896);
xnor U4142 (N_4142,N_3990,N_3866);
and U4143 (N_4143,N_3848,N_3829);
or U4144 (N_4144,N_3878,N_3991);
nand U4145 (N_4145,N_3998,N_3853);
and U4146 (N_4146,N_3953,N_3881);
xnor U4147 (N_4147,N_3914,N_3894);
and U4148 (N_4148,N_3940,N_3879);
and U4149 (N_4149,N_3911,N_3909);
nor U4150 (N_4150,N_3846,N_3909);
and U4151 (N_4151,N_3911,N_3977);
and U4152 (N_4152,N_3905,N_3876);
or U4153 (N_4153,N_3960,N_3982);
nor U4154 (N_4154,N_3838,N_3862);
nor U4155 (N_4155,N_3929,N_3960);
nand U4156 (N_4156,N_3826,N_3899);
nand U4157 (N_4157,N_3924,N_3853);
and U4158 (N_4158,N_3963,N_3825);
nor U4159 (N_4159,N_3884,N_3903);
nand U4160 (N_4160,N_3937,N_3990);
and U4161 (N_4161,N_3965,N_3802);
or U4162 (N_4162,N_3838,N_3929);
nor U4163 (N_4163,N_3902,N_3944);
and U4164 (N_4164,N_3999,N_3888);
and U4165 (N_4165,N_3977,N_3867);
nand U4166 (N_4166,N_3817,N_3966);
nor U4167 (N_4167,N_3878,N_3804);
or U4168 (N_4168,N_3902,N_3978);
nand U4169 (N_4169,N_3884,N_3965);
and U4170 (N_4170,N_3835,N_3999);
xnor U4171 (N_4171,N_3927,N_3990);
or U4172 (N_4172,N_3988,N_3842);
nor U4173 (N_4173,N_3981,N_3989);
and U4174 (N_4174,N_3891,N_3918);
nor U4175 (N_4175,N_3898,N_3908);
xor U4176 (N_4176,N_3919,N_3815);
xnor U4177 (N_4177,N_3960,N_3987);
nand U4178 (N_4178,N_3934,N_3943);
xor U4179 (N_4179,N_3843,N_3962);
xor U4180 (N_4180,N_3849,N_3802);
or U4181 (N_4181,N_3882,N_3885);
nand U4182 (N_4182,N_3802,N_3808);
nor U4183 (N_4183,N_3906,N_3844);
and U4184 (N_4184,N_3831,N_3994);
xor U4185 (N_4185,N_3927,N_3982);
nand U4186 (N_4186,N_3907,N_3975);
xor U4187 (N_4187,N_3813,N_3965);
nand U4188 (N_4188,N_3991,N_3988);
xnor U4189 (N_4189,N_3956,N_3879);
and U4190 (N_4190,N_3838,N_3915);
and U4191 (N_4191,N_3902,N_3950);
or U4192 (N_4192,N_3891,N_3962);
or U4193 (N_4193,N_3944,N_3806);
and U4194 (N_4194,N_3974,N_3913);
xor U4195 (N_4195,N_3941,N_3823);
nand U4196 (N_4196,N_3803,N_3965);
and U4197 (N_4197,N_3850,N_3927);
and U4198 (N_4198,N_3876,N_3983);
and U4199 (N_4199,N_3815,N_3853);
or U4200 (N_4200,N_4007,N_4124);
and U4201 (N_4201,N_4147,N_4188);
or U4202 (N_4202,N_4129,N_4165);
xor U4203 (N_4203,N_4000,N_4051);
nand U4204 (N_4204,N_4178,N_4155);
xor U4205 (N_4205,N_4018,N_4008);
nor U4206 (N_4206,N_4162,N_4024);
nor U4207 (N_4207,N_4002,N_4092);
or U4208 (N_4208,N_4006,N_4125);
or U4209 (N_4209,N_4056,N_4140);
nand U4210 (N_4210,N_4060,N_4119);
xor U4211 (N_4211,N_4080,N_4132);
xor U4212 (N_4212,N_4020,N_4109);
xnor U4213 (N_4213,N_4148,N_4138);
nand U4214 (N_4214,N_4052,N_4016);
and U4215 (N_4215,N_4120,N_4076);
nor U4216 (N_4216,N_4185,N_4088);
or U4217 (N_4217,N_4143,N_4036);
xnor U4218 (N_4218,N_4037,N_4117);
nand U4219 (N_4219,N_4010,N_4096);
or U4220 (N_4220,N_4111,N_4174);
nand U4221 (N_4221,N_4048,N_4028);
or U4222 (N_4222,N_4061,N_4047);
nand U4223 (N_4223,N_4108,N_4160);
and U4224 (N_4224,N_4176,N_4019);
nor U4225 (N_4225,N_4089,N_4003);
and U4226 (N_4226,N_4103,N_4110);
nor U4227 (N_4227,N_4104,N_4102);
or U4228 (N_4228,N_4022,N_4070);
nor U4229 (N_4229,N_4091,N_4075);
or U4230 (N_4230,N_4121,N_4023);
and U4231 (N_4231,N_4191,N_4131);
or U4232 (N_4232,N_4163,N_4063);
nand U4233 (N_4233,N_4133,N_4149);
xor U4234 (N_4234,N_4180,N_4021);
nand U4235 (N_4235,N_4098,N_4106);
nor U4236 (N_4236,N_4194,N_4053);
xor U4237 (N_4237,N_4087,N_4164);
or U4238 (N_4238,N_4057,N_4058);
xor U4239 (N_4239,N_4077,N_4083);
nand U4240 (N_4240,N_4090,N_4025);
xnor U4241 (N_4241,N_4142,N_4179);
or U4242 (N_4242,N_4038,N_4084);
nor U4243 (N_4243,N_4095,N_4186);
nand U4244 (N_4244,N_4137,N_4099);
nand U4245 (N_4245,N_4113,N_4001);
and U4246 (N_4246,N_4141,N_4146);
nand U4247 (N_4247,N_4127,N_4190);
or U4248 (N_4248,N_4045,N_4065);
or U4249 (N_4249,N_4173,N_4115);
and U4250 (N_4250,N_4156,N_4054);
nor U4251 (N_4251,N_4112,N_4093);
xor U4252 (N_4252,N_4184,N_4050);
and U4253 (N_4253,N_4042,N_4114);
or U4254 (N_4254,N_4105,N_4150);
or U4255 (N_4255,N_4086,N_4192);
or U4256 (N_4256,N_4081,N_4066);
nand U4257 (N_4257,N_4055,N_4122);
xor U4258 (N_4258,N_4159,N_4014);
nor U4259 (N_4259,N_4015,N_4175);
nor U4260 (N_4260,N_4168,N_4074);
nor U4261 (N_4261,N_4130,N_4004);
or U4262 (N_4262,N_4177,N_4123);
and U4263 (N_4263,N_4073,N_4035);
or U4264 (N_4264,N_4139,N_4135);
xnor U4265 (N_4265,N_4079,N_4012);
nor U4266 (N_4266,N_4082,N_4161);
nor U4267 (N_4267,N_4166,N_4152);
or U4268 (N_4268,N_4072,N_4187);
nor U4269 (N_4269,N_4044,N_4198);
nor U4270 (N_4270,N_4134,N_4064);
nand U4271 (N_4271,N_4199,N_4043);
and U4272 (N_4272,N_4062,N_4011);
nor U4273 (N_4273,N_4032,N_4101);
and U4274 (N_4274,N_4026,N_4170);
xnor U4275 (N_4275,N_4033,N_4071);
nand U4276 (N_4276,N_4107,N_4069);
xnor U4277 (N_4277,N_4034,N_4040);
and U4278 (N_4278,N_4067,N_4145);
xnor U4279 (N_4279,N_4157,N_4151);
or U4280 (N_4280,N_4195,N_4017);
nor U4281 (N_4281,N_4027,N_4171);
nor U4282 (N_4282,N_4158,N_4030);
and U4283 (N_4283,N_4029,N_4059);
or U4284 (N_4284,N_4154,N_4068);
and U4285 (N_4285,N_4005,N_4169);
xor U4286 (N_4286,N_4085,N_4116);
nor U4287 (N_4287,N_4031,N_4118);
or U4288 (N_4288,N_4136,N_4167);
or U4289 (N_4289,N_4078,N_4039);
xor U4290 (N_4290,N_4046,N_4153);
nor U4291 (N_4291,N_4049,N_4144);
nor U4292 (N_4292,N_4182,N_4100);
xnor U4293 (N_4293,N_4193,N_4189);
and U4294 (N_4294,N_4197,N_4181);
or U4295 (N_4295,N_4196,N_4126);
nand U4296 (N_4296,N_4013,N_4094);
nor U4297 (N_4297,N_4009,N_4041);
or U4298 (N_4298,N_4097,N_4172);
nor U4299 (N_4299,N_4128,N_4183);
and U4300 (N_4300,N_4133,N_4062);
nand U4301 (N_4301,N_4048,N_4093);
nand U4302 (N_4302,N_4028,N_4122);
and U4303 (N_4303,N_4115,N_4007);
or U4304 (N_4304,N_4080,N_4092);
nand U4305 (N_4305,N_4116,N_4123);
or U4306 (N_4306,N_4052,N_4158);
or U4307 (N_4307,N_4075,N_4102);
and U4308 (N_4308,N_4145,N_4117);
and U4309 (N_4309,N_4136,N_4037);
nand U4310 (N_4310,N_4149,N_4024);
nor U4311 (N_4311,N_4036,N_4086);
xor U4312 (N_4312,N_4172,N_4127);
or U4313 (N_4313,N_4086,N_4091);
nand U4314 (N_4314,N_4172,N_4014);
nor U4315 (N_4315,N_4109,N_4183);
xor U4316 (N_4316,N_4181,N_4188);
nor U4317 (N_4317,N_4056,N_4166);
nor U4318 (N_4318,N_4066,N_4080);
nor U4319 (N_4319,N_4015,N_4126);
xor U4320 (N_4320,N_4173,N_4056);
and U4321 (N_4321,N_4169,N_4106);
xor U4322 (N_4322,N_4054,N_4081);
nand U4323 (N_4323,N_4165,N_4044);
nor U4324 (N_4324,N_4019,N_4075);
xnor U4325 (N_4325,N_4054,N_4020);
nor U4326 (N_4326,N_4089,N_4091);
nor U4327 (N_4327,N_4077,N_4057);
nor U4328 (N_4328,N_4094,N_4184);
and U4329 (N_4329,N_4038,N_4145);
xnor U4330 (N_4330,N_4064,N_4019);
or U4331 (N_4331,N_4035,N_4138);
and U4332 (N_4332,N_4147,N_4141);
and U4333 (N_4333,N_4176,N_4143);
xnor U4334 (N_4334,N_4112,N_4175);
xor U4335 (N_4335,N_4041,N_4062);
nor U4336 (N_4336,N_4111,N_4150);
nor U4337 (N_4337,N_4153,N_4060);
or U4338 (N_4338,N_4020,N_4167);
or U4339 (N_4339,N_4086,N_4159);
nor U4340 (N_4340,N_4173,N_4137);
xnor U4341 (N_4341,N_4087,N_4062);
and U4342 (N_4342,N_4127,N_4034);
and U4343 (N_4343,N_4105,N_4078);
nor U4344 (N_4344,N_4170,N_4066);
nand U4345 (N_4345,N_4061,N_4082);
and U4346 (N_4346,N_4148,N_4136);
nor U4347 (N_4347,N_4161,N_4045);
or U4348 (N_4348,N_4090,N_4127);
xor U4349 (N_4349,N_4119,N_4056);
nand U4350 (N_4350,N_4043,N_4001);
nor U4351 (N_4351,N_4102,N_4116);
xor U4352 (N_4352,N_4033,N_4091);
nor U4353 (N_4353,N_4106,N_4108);
and U4354 (N_4354,N_4046,N_4073);
xnor U4355 (N_4355,N_4054,N_4152);
xor U4356 (N_4356,N_4092,N_4097);
or U4357 (N_4357,N_4182,N_4027);
or U4358 (N_4358,N_4019,N_4166);
or U4359 (N_4359,N_4196,N_4045);
and U4360 (N_4360,N_4073,N_4119);
nor U4361 (N_4361,N_4036,N_4079);
or U4362 (N_4362,N_4083,N_4094);
nor U4363 (N_4363,N_4167,N_4088);
xor U4364 (N_4364,N_4027,N_4041);
or U4365 (N_4365,N_4053,N_4070);
xor U4366 (N_4366,N_4165,N_4065);
nand U4367 (N_4367,N_4041,N_4047);
nand U4368 (N_4368,N_4066,N_4162);
nor U4369 (N_4369,N_4086,N_4169);
or U4370 (N_4370,N_4101,N_4140);
nor U4371 (N_4371,N_4056,N_4109);
nor U4372 (N_4372,N_4147,N_4190);
nand U4373 (N_4373,N_4198,N_4165);
or U4374 (N_4374,N_4103,N_4087);
nor U4375 (N_4375,N_4077,N_4184);
or U4376 (N_4376,N_4150,N_4014);
nand U4377 (N_4377,N_4110,N_4167);
xor U4378 (N_4378,N_4128,N_4075);
nand U4379 (N_4379,N_4120,N_4050);
or U4380 (N_4380,N_4000,N_4146);
nor U4381 (N_4381,N_4048,N_4059);
xnor U4382 (N_4382,N_4080,N_4193);
nand U4383 (N_4383,N_4055,N_4074);
xnor U4384 (N_4384,N_4104,N_4065);
nand U4385 (N_4385,N_4127,N_4108);
and U4386 (N_4386,N_4194,N_4102);
nor U4387 (N_4387,N_4003,N_4114);
xnor U4388 (N_4388,N_4103,N_4163);
xor U4389 (N_4389,N_4161,N_4087);
or U4390 (N_4390,N_4019,N_4195);
xnor U4391 (N_4391,N_4133,N_4184);
or U4392 (N_4392,N_4157,N_4121);
or U4393 (N_4393,N_4036,N_4092);
and U4394 (N_4394,N_4010,N_4138);
and U4395 (N_4395,N_4093,N_4163);
nand U4396 (N_4396,N_4016,N_4199);
or U4397 (N_4397,N_4044,N_4006);
xnor U4398 (N_4398,N_4156,N_4080);
or U4399 (N_4399,N_4080,N_4012);
xor U4400 (N_4400,N_4254,N_4381);
or U4401 (N_4401,N_4251,N_4263);
xnor U4402 (N_4402,N_4375,N_4367);
or U4403 (N_4403,N_4359,N_4270);
xor U4404 (N_4404,N_4265,N_4313);
or U4405 (N_4405,N_4348,N_4278);
and U4406 (N_4406,N_4388,N_4389);
xor U4407 (N_4407,N_4258,N_4292);
nor U4408 (N_4408,N_4299,N_4261);
nand U4409 (N_4409,N_4245,N_4391);
nor U4410 (N_4410,N_4343,N_4316);
and U4411 (N_4411,N_4344,N_4320);
or U4412 (N_4412,N_4221,N_4330);
nor U4413 (N_4413,N_4370,N_4253);
xor U4414 (N_4414,N_4264,N_4252);
xor U4415 (N_4415,N_4218,N_4339);
and U4416 (N_4416,N_4276,N_4303);
and U4417 (N_4417,N_4345,N_4259);
nand U4418 (N_4418,N_4396,N_4200);
nor U4419 (N_4419,N_4301,N_4256);
xnor U4420 (N_4420,N_4394,N_4329);
nand U4421 (N_4421,N_4209,N_4380);
nor U4422 (N_4422,N_4277,N_4351);
nor U4423 (N_4423,N_4202,N_4268);
nor U4424 (N_4424,N_4358,N_4311);
xnor U4425 (N_4425,N_4287,N_4347);
nor U4426 (N_4426,N_4315,N_4309);
nand U4427 (N_4427,N_4314,N_4332);
xor U4428 (N_4428,N_4233,N_4338);
xnor U4429 (N_4429,N_4286,N_4235);
xor U4430 (N_4430,N_4369,N_4323);
xor U4431 (N_4431,N_4239,N_4398);
and U4432 (N_4432,N_4364,N_4217);
nand U4433 (N_4433,N_4232,N_4372);
nor U4434 (N_4434,N_4335,N_4331);
or U4435 (N_4435,N_4368,N_4360);
or U4436 (N_4436,N_4262,N_4298);
nand U4437 (N_4437,N_4291,N_4296);
nor U4438 (N_4438,N_4294,N_4207);
or U4439 (N_4439,N_4365,N_4377);
xor U4440 (N_4440,N_4322,N_4290);
and U4441 (N_4441,N_4229,N_4237);
and U4442 (N_4442,N_4336,N_4385);
xnor U4443 (N_4443,N_4272,N_4371);
or U4444 (N_4444,N_4305,N_4378);
or U4445 (N_4445,N_4242,N_4214);
nand U4446 (N_4446,N_4395,N_4234);
and U4447 (N_4447,N_4279,N_4220);
nand U4448 (N_4448,N_4241,N_4224);
xnor U4449 (N_4449,N_4350,N_4204);
nor U4450 (N_4450,N_4205,N_4379);
or U4451 (N_4451,N_4215,N_4228);
nand U4452 (N_4452,N_4310,N_4302);
nand U4453 (N_4453,N_4231,N_4297);
or U4454 (N_4454,N_4269,N_4266);
nand U4455 (N_4455,N_4333,N_4308);
xor U4456 (N_4456,N_4366,N_4295);
nor U4457 (N_4457,N_4280,N_4300);
and U4458 (N_4458,N_4293,N_4283);
and U4459 (N_4459,N_4304,N_4353);
or U4460 (N_4460,N_4206,N_4392);
nor U4461 (N_4461,N_4354,N_4376);
and U4462 (N_4462,N_4374,N_4219);
nand U4463 (N_4463,N_4230,N_4247);
nor U4464 (N_4464,N_4324,N_4307);
nand U4465 (N_4465,N_4222,N_4361);
xnor U4466 (N_4466,N_4321,N_4267);
xnor U4467 (N_4467,N_4274,N_4273);
nand U4468 (N_4468,N_4227,N_4362);
nand U4469 (N_4469,N_4225,N_4352);
nor U4470 (N_4470,N_4355,N_4238);
nor U4471 (N_4471,N_4210,N_4260);
and U4472 (N_4472,N_4211,N_4203);
xor U4473 (N_4473,N_4326,N_4208);
nor U4474 (N_4474,N_4341,N_4393);
xor U4475 (N_4475,N_4387,N_4312);
nand U4476 (N_4476,N_4281,N_4386);
nand U4477 (N_4477,N_4340,N_4243);
and U4478 (N_4478,N_4325,N_4257);
nand U4479 (N_4479,N_4216,N_4318);
nor U4480 (N_4480,N_4383,N_4342);
nor U4481 (N_4481,N_4346,N_4249);
or U4482 (N_4482,N_4373,N_4226);
nor U4483 (N_4483,N_4319,N_4271);
or U4484 (N_4484,N_4255,N_4357);
or U4485 (N_4485,N_4328,N_4288);
xnor U4486 (N_4486,N_4289,N_4334);
and U4487 (N_4487,N_4212,N_4349);
and U4488 (N_4488,N_4236,N_4284);
and U4489 (N_4489,N_4363,N_4285);
and U4490 (N_4490,N_4382,N_4201);
nand U4491 (N_4491,N_4240,N_4390);
or U4492 (N_4492,N_4246,N_4399);
nor U4493 (N_4493,N_4223,N_4306);
or U4494 (N_4494,N_4356,N_4244);
nor U4495 (N_4495,N_4248,N_4282);
nand U4496 (N_4496,N_4337,N_4213);
xnor U4497 (N_4497,N_4317,N_4327);
nor U4498 (N_4498,N_4275,N_4384);
or U4499 (N_4499,N_4397,N_4250);
and U4500 (N_4500,N_4306,N_4341);
xnor U4501 (N_4501,N_4321,N_4389);
and U4502 (N_4502,N_4274,N_4332);
or U4503 (N_4503,N_4225,N_4266);
and U4504 (N_4504,N_4278,N_4305);
and U4505 (N_4505,N_4260,N_4218);
or U4506 (N_4506,N_4294,N_4399);
nand U4507 (N_4507,N_4280,N_4398);
and U4508 (N_4508,N_4341,N_4219);
or U4509 (N_4509,N_4329,N_4335);
nor U4510 (N_4510,N_4265,N_4277);
xnor U4511 (N_4511,N_4314,N_4364);
nand U4512 (N_4512,N_4229,N_4220);
nand U4513 (N_4513,N_4391,N_4237);
xor U4514 (N_4514,N_4265,N_4352);
nor U4515 (N_4515,N_4234,N_4211);
or U4516 (N_4516,N_4335,N_4298);
nor U4517 (N_4517,N_4218,N_4315);
and U4518 (N_4518,N_4382,N_4348);
or U4519 (N_4519,N_4247,N_4313);
nand U4520 (N_4520,N_4368,N_4252);
nor U4521 (N_4521,N_4219,N_4230);
or U4522 (N_4522,N_4283,N_4303);
xnor U4523 (N_4523,N_4347,N_4207);
and U4524 (N_4524,N_4306,N_4318);
nand U4525 (N_4525,N_4238,N_4292);
nand U4526 (N_4526,N_4279,N_4253);
and U4527 (N_4527,N_4380,N_4331);
or U4528 (N_4528,N_4390,N_4224);
xnor U4529 (N_4529,N_4351,N_4394);
nand U4530 (N_4530,N_4314,N_4233);
and U4531 (N_4531,N_4392,N_4332);
nor U4532 (N_4532,N_4317,N_4323);
nor U4533 (N_4533,N_4256,N_4320);
xnor U4534 (N_4534,N_4233,N_4283);
nor U4535 (N_4535,N_4229,N_4326);
nand U4536 (N_4536,N_4224,N_4336);
or U4537 (N_4537,N_4234,N_4338);
xor U4538 (N_4538,N_4206,N_4214);
or U4539 (N_4539,N_4315,N_4213);
and U4540 (N_4540,N_4220,N_4398);
xor U4541 (N_4541,N_4238,N_4375);
nor U4542 (N_4542,N_4206,N_4270);
nor U4543 (N_4543,N_4359,N_4211);
or U4544 (N_4544,N_4358,N_4360);
or U4545 (N_4545,N_4371,N_4220);
nor U4546 (N_4546,N_4323,N_4316);
xnor U4547 (N_4547,N_4228,N_4220);
and U4548 (N_4548,N_4292,N_4306);
xnor U4549 (N_4549,N_4275,N_4250);
or U4550 (N_4550,N_4347,N_4203);
xor U4551 (N_4551,N_4232,N_4364);
xor U4552 (N_4552,N_4302,N_4204);
or U4553 (N_4553,N_4335,N_4334);
or U4554 (N_4554,N_4249,N_4366);
xor U4555 (N_4555,N_4297,N_4217);
or U4556 (N_4556,N_4383,N_4321);
and U4557 (N_4557,N_4365,N_4306);
or U4558 (N_4558,N_4277,N_4202);
or U4559 (N_4559,N_4245,N_4233);
or U4560 (N_4560,N_4370,N_4380);
and U4561 (N_4561,N_4349,N_4245);
or U4562 (N_4562,N_4210,N_4350);
and U4563 (N_4563,N_4267,N_4399);
nor U4564 (N_4564,N_4295,N_4231);
and U4565 (N_4565,N_4376,N_4331);
nor U4566 (N_4566,N_4337,N_4331);
nand U4567 (N_4567,N_4331,N_4384);
xor U4568 (N_4568,N_4272,N_4291);
nand U4569 (N_4569,N_4298,N_4247);
and U4570 (N_4570,N_4340,N_4237);
and U4571 (N_4571,N_4347,N_4379);
xnor U4572 (N_4572,N_4238,N_4366);
nand U4573 (N_4573,N_4290,N_4308);
or U4574 (N_4574,N_4267,N_4290);
and U4575 (N_4575,N_4392,N_4379);
nand U4576 (N_4576,N_4333,N_4254);
and U4577 (N_4577,N_4292,N_4280);
and U4578 (N_4578,N_4291,N_4270);
nor U4579 (N_4579,N_4231,N_4395);
or U4580 (N_4580,N_4291,N_4374);
xor U4581 (N_4581,N_4232,N_4260);
and U4582 (N_4582,N_4388,N_4218);
xnor U4583 (N_4583,N_4232,N_4345);
xnor U4584 (N_4584,N_4227,N_4271);
nand U4585 (N_4585,N_4273,N_4258);
nor U4586 (N_4586,N_4364,N_4345);
nand U4587 (N_4587,N_4306,N_4382);
and U4588 (N_4588,N_4254,N_4205);
nor U4589 (N_4589,N_4262,N_4309);
nand U4590 (N_4590,N_4279,N_4232);
nand U4591 (N_4591,N_4341,N_4394);
nand U4592 (N_4592,N_4248,N_4270);
or U4593 (N_4593,N_4375,N_4220);
and U4594 (N_4594,N_4265,N_4375);
or U4595 (N_4595,N_4257,N_4304);
nor U4596 (N_4596,N_4297,N_4293);
nor U4597 (N_4597,N_4234,N_4285);
nor U4598 (N_4598,N_4298,N_4346);
or U4599 (N_4599,N_4300,N_4342);
and U4600 (N_4600,N_4552,N_4412);
nand U4601 (N_4601,N_4463,N_4562);
nor U4602 (N_4602,N_4422,N_4477);
nor U4603 (N_4603,N_4486,N_4569);
nand U4604 (N_4604,N_4518,N_4540);
xnor U4605 (N_4605,N_4456,N_4406);
or U4606 (N_4606,N_4430,N_4564);
or U4607 (N_4607,N_4413,N_4555);
and U4608 (N_4608,N_4516,N_4590);
or U4609 (N_4609,N_4528,N_4587);
nand U4610 (N_4610,N_4597,N_4480);
or U4611 (N_4611,N_4554,N_4451);
nor U4612 (N_4612,N_4556,N_4548);
nor U4613 (N_4613,N_4592,N_4478);
or U4614 (N_4614,N_4432,N_4408);
and U4615 (N_4615,N_4561,N_4467);
xnor U4616 (N_4616,N_4433,N_4434);
nor U4617 (N_4617,N_4489,N_4424);
nand U4618 (N_4618,N_4539,N_4565);
nand U4619 (N_4619,N_4541,N_4446);
nor U4620 (N_4620,N_4466,N_4510);
and U4621 (N_4621,N_4411,N_4410);
nand U4622 (N_4622,N_4511,N_4581);
xnor U4623 (N_4623,N_4538,N_4537);
nand U4624 (N_4624,N_4496,N_4560);
nor U4625 (N_4625,N_4534,N_4574);
or U4626 (N_4626,N_4495,N_4551);
nand U4627 (N_4627,N_4567,N_4414);
nand U4628 (N_4628,N_4461,N_4519);
nand U4629 (N_4629,N_4576,N_4514);
nor U4630 (N_4630,N_4595,N_4525);
and U4631 (N_4631,N_4512,N_4490);
nor U4632 (N_4632,N_4545,N_4481);
and U4633 (N_4633,N_4521,N_4426);
or U4634 (N_4634,N_4493,N_4483);
xor U4635 (N_4635,N_4582,N_4457);
xnor U4636 (N_4636,N_4444,N_4455);
and U4637 (N_4637,N_4454,N_4515);
xor U4638 (N_4638,N_4578,N_4579);
or U4639 (N_4639,N_4400,N_4500);
or U4640 (N_4640,N_4474,N_4487);
and U4641 (N_4641,N_4476,N_4494);
nand U4642 (N_4642,N_4445,N_4558);
xnor U4643 (N_4643,N_4543,N_4584);
nor U4644 (N_4644,N_4563,N_4425);
or U4645 (N_4645,N_4462,N_4417);
and U4646 (N_4646,N_4501,N_4507);
xor U4647 (N_4647,N_4459,N_4469);
or U4648 (N_4648,N_4453,N_4404);
nor U4649 (N_4649,N_4508,N_4568);
xor U4650 (N_4650,N_4416,N_4465);
or U4651 (N_4651,N_4475,N_4547);
nor U4652 (N_4652,N_4421,N_4409);
and U4653 (N_4653,N_4530,N_4588);
or U4654 (N_4654,N_4471,N_4529);
nor U4655 (N_4655,N_4485,N_4427);
and U4656 (N_4656,N_4441,N_4403);
nor U4657 (N_4657,N_4532,N_4491);
nand U4658 (N_4658,N_4488,N_4436);
xor U4659 (N_4659,N_4492,N_4509);
nand U4660 (N_4660,N_4502,N_4513);
xor U4661 (N_4661,N_4442,N_4447);
or U4662 (N_4662,N_4520,N_4449);
or U4663 (N_4663,N_4580,N_4533);
nand U4664 (N_4664,N_4415,N_4577);
and U4665 (N_4665,N_4504,N_4591);
or U4666 (N_4666,N_4458,N_4570);
and U4667 (N_4667,N_4517,N_4499);
nand U4668 (N_4668,N_4535,N_4460);
and U4669 (N_4669,N_4448,N_4472);
and U4670 (N_4670,N_4527,N_4407);
nor U4671 (N_4671,N_4571,N_4435);
or U4672 (N_4672,N_4575,N_4573);
nand U4673 (N_4673,N_4526,N_4440);
nor U4674 (N_4674,N_4546,N_4572);
and U4675 (N_4675,N_4401,N_4549);
and U4676 (N_4676,N_4484,N_4450);
or U4677 (N_4677,N_4438,N_4420);
xor U4678 (N_4678,N_4524,N_4503);
nor U4679 (N_4679,N_4418,N_4583);
nor U4680 (N_4680,N_4522,N_4594);
nand U4681 (N_4681,N_4586,N_4531);
nor U4682 (N_4682,N_4498,N_4405);
nand U4683 (N_4683,N_4557,N_4497);
nor U4684 (N_4684,N_4599,N_4402);
xor U4685 (N_4685,N_4479,N_4593);
nand U4686 (N_4686,N_4429,N_4468);
nand U4687 (N_4687,N_4428,N_4431);
xor U4688 (N_4688,N_4423,N_4505);
xor U4689 (N_4689,N_4452,N_4523);
or U4690 (N_4690,N_4544,N_4585);
and U4691 (N_4691,N_4464,N_4550);
xnor U4692 (N_4692,N_4566,N_4506);
nand U4693 (N_4693,N_4419,N_4589);
nand U4694 (N_4694,N_4470,N_4443);
or U4695 (N_4695,N_4553,N_4559);
nand U4696 (N_4696,N_4437,N_4542);
nand U4697 (N_4697,N_4482,N_4596);
and U4698 (N_4698,N_4439,N_4598);
xnor U4699 (N_4699,N_4536,N_4473);
nand U4700 (N_4700,N_4467,N_4596);
and U4701 (N_4701,N_4462,N_4450);
and U4702 (N_4702,N_4541,N_4511);
nand U4703 (N_4703,N_4427,N_4465);
or U4704 (N_4704,N_4533,N_4598);
nor U4705 (N_4705,N_4589,N_4573);
nand U4706 (N_4706,N_4484,N_4517);
nor U4707 (N_4707,N_4506,N_4555);
or U4708 (N_4708,N_4480,N_4405);
nor U4709 (N_4709,N_4407,N_4539);
or U4710 (N_4710,N_4467,N_4563);
or U4711 (N_4711,N_4598,N_4596);
and U4712 (N_4712,N_4570,N_4416);
and U4713 (N_4713,N_4449,N_4537);
or U4714 (N_4714,N_4448,N_4587);
nor U4715 (N_4715,N_4574,N_4453);
nand U4716 (N_4716,N_4472,N_4486);
or U4717 (N_4717,N_4484,N_4594);
or U4718 (N_4718,N_4565,N_4472);
and U4719 (N_4719,N_4409,N_4506);
nand U4720 (N_4720,N_4409,N_4497);
nand U4721 (N_4721,N_4435,N_4462);
or U4722 (N_4722,N_4404,N_4539);
nand U4723 (N_4723,N_4532,N_4558);
and U4724 (N_4724,N_4499,N_4512);
xnor U4725 (N_4725,N_4485,N_4488);
and U4726 (N_4726,N_4505,N_4441);
xnor U4727 (N_4727,N_4418,N_4452);
nor U4728 (N_4728,N_4530,N_4598);
xor U4729 (N_4729,N_4484,N_4406);
xnor U4730 (N_4730,N_4456,N_4484);
or U4731 (N_4731,N_4467,N_4594);
or U4732 (N_4732,N_4499,N_4556);
nor U4733 (N_4733,N_4449,N_4455);
or U4734 (N_4734,N_4464,N_4581);
xor U4735 (N_4735,N_4482,N_4571);
xnor U4736 (N_4736,N_4478,N_4517);
nor U4737 (N_4737,N_4499,N_4432);
nor U4738 (N_4738,N_4558,N_4577);
nand U4739 (N_4739,N_4423,N_4430);
xor U4740 (N_4740,N_4405,N_4453);
xnor U4741 (N_4741,N_4412,N_4505);
nor U4742 (N_4742,N_4554,N_4536);
nor U4743 (N_4743,N_4453,N_4435);
or U4744 (N_4744,N_4490,N_4416);
nand U4745 (N_4745,N_4486,N_4423);
nor U4746 (N_4746,N_4562,N_4509);
nand U4747 (N_4747,N_4432,N_4570);
or U4748 (N_4748,N_4412,N_4492);
or U4749 (N_4749,N_4523,N_4407);
nor U4750 (N_4750,N_4501,N_4494);
nor U4751 (N_4751,N_4508,N_4533);
nor U4752 (N_4752,N_4506,N_4469);
nand U4753 (N_4753,N_4569,N_4533);
xor U4754 (N_4754,N_4501,N_4486);
or U4755 (N_4755,N_4492,N_4557);
nand U4756 (N_4756,N_4471,N_4400);
xor U4757 (N_4757,N_4598,N_4480);
xnor U4758 (N_4758,N_4509,N_4502);
nand U4759 (N_4759,N_4478,N_4461);
and U4760 (N_4760,N_4457,N_4442);
xnor U4761 (N_4761,N_4462,N_4503);
nor U4762 (N_4762,N_4518,N_4443);
nor U4763 (N_4763,N_4594,N_4570);
and U4764 (N_4764,N_4478,N_4434);
xnor U4765 (N_4765,N_4408,N_4469);
and U4766 (N_4766,N_4498,N_4502);
or U4767 (N_4767,N_4453,N_4485);
and U4768 (N_4768,N_4534,N_4502);
xor U4769 (N_4769,N_4400,N_4488);
xor U4770 (N_4770,N_4498,N_4486);
nand U4771 (N_4771,N_4493,N_4547);
nand U4772 (N_4772,N_4487,N_4484);
nand U4773 (N_4773,N_4575,N_4417);
or U4774 (N_4774,N_4419,N_4563);
xnor U4775 (N_4775,N_4581,N_4452);
nor U4776 (N_4776,N_4466,N_4517);
nor U4777 (N_4777,N_4518,N_4496);
and U4778 (N_4778,N_4498,N_4536);
or U4779 (N_4779,N_4504,N_4571);
and U4780 (N_4780,N_4528,N_4458);
nor U4781 (N_4781,N_4425,N_4434);
and U4782 (N_4782,N_4403,N_4455);
or U4783 (N_4783,N_4506,N_4479);
nor U4784 (N_4784,N_4406,N_4525);
xor U4785 (N_4785,N_4596,N_4420);
or U4786 (N_4786,N_4449,N_4575);
nor U4787 (N_4787,N_4465,N_4535);
nor U4788 (N_4788,N_4549,N_4449);
or U4789 (N_4789,N_4420,N_4552);
and U4790 (N_4790,N_4559,N_4549);
and U4791 (N_4791,N_4560,N_4408);
or U4792 (N_4792,N_4586,N_4548);
and U4793 (N_4793,N_4407,N_4541);
or U4794 (N_4794,N_4432,N_4560);
and U4795 (N_4795,N_4407,N_4492);
or U4796 (N_4796,N_4447,N_4443);
and U4797 (N_4797,N_4586,N_4583);
nand U4798 (N_4798,N_4514,N_4530);
nand U4799 (N_4799,N_4509,N_4522);
or U4800 (N_4800,N_4750,N_4612);
or U4801 (N_4801,N_4795,N_4711);
or U4802 (N_4802,N_4702,N_4746);
or U4803 (N_4803,N_4768,N_4726);
xnor U4804 (N_4804,N_4668,N_4727);
and U4805 (N_4805,N_4775,N_4794);
nand U4806 (N_4806,N_4766,N_4632);
and U4807 (N_4807,N_4622,N_4601);
or U4808 (N_4808,N_4740,N_4783);
nand U4809 (N_4809,N_4686,N_4685);
or U4810 (N_4810,N_4695,N_4673);
nor U4811 (N_4811,N_4617,N_4646);
nand U4812 (N_4812,N_4782,N_4774);
or U4813 (N_4813,N_4738,N_4614);
or U4814 (N_4814,N_4644,N_4630);
xor U4815 (N_4815,N_4762,N_4694);
or U4816 (N_4816,N_4781,N_4708);
nor U4817 (N_4817,N_4682,N_4714);
nor U4818 (N_4818,N_4643,N_4664);
nand U4819 (N_4819,N_4789,N_4628);
nand U4820 (N_4820,N_4667,N_4602);
nand U4821 (N_4821,N_4676,N_4637);
or U4822 (N_4822,N_4786,N_4733);
nand U4823 (N_4823,N_4680,N_4700);
and U4824 (N_4824,N_4732,N_4712);
nor U4825 (N_4825,N_4791,N_4716);
xor U4826 (N_4826,N_4698,N_4703);
and U4827 (N_4827,N_4736,N_4785);
xnor U4828 (N_4828,N_4689,N_4649);
and U4829 (N_4829,N_4705,N_4749);
or U4830 (N_4830,N_4769,N_4798);
or U4831 (N_4831,N_4606,N_4793);
nor U4832 (N_4832,N_4797,N_4629);
nand U4833 (N_4833,N_4745,N_4659);
and U4834 (N_4834,N_4784,N_4725);
nand U4835 (N_4835,N_4707,N_4709);
and U4836 (N_4836,N_4619,N_4600);
and U4837 (N_4837,N_4669,N_4739);
and U4838 (N_4838,N_4687,N_4743);
nand U4839 (N_4839,N_4760,N_4677);
xnor U4840 (N_4840,N_4660,N_4620);
or U4841 (N_4841,N_4672,N_4737);
nand U4842 (N_4842,N_4790,N_4603);
nor U4843 (N_4843,N_4652,N_4621);
xor U4844 (N_4844,N_4751,N_4661);
xor U4845 (N_4845,N_4616,N_4719);
xor U4846 (N_4846,N_4650,N_4615);
and U4847 (N_4847,N_4688,N_4710);
xor U4848 (N_4848,N_4610,N_4748);
nand U4849 (N_4849,N_4605,N_4720);
nand U4850 (N_4850,N_4666,N_4654);
nand U4851 (N_4851,N_4763,N_4772);
or U4852 (N_4852,N_4777,N_4640);
nor U4853 (N_4853,N_4758,N_4706);
xnor U4854 (N_4854,N_4756,N_4690);
nor U4855 (N_4855,N_4657,N_4627);
nand U4856 (N_4856,N_4773,N_4747);
nand U4857 (N_4857,N_4724,N_4771);
or U4858 (N_4858,N_4626,N_4735);
xnor U4859 (N_4859,N_4641,N_4681);
or U4860 (N_4860,N_4618,N_4665);
and U4861 (N_4861,N_4761,N_4757);
and U4862 (N_4862,N_4752,N_4679);
or U4863 (N_4863,N_4765,N_4683);
nor U4864 (N_4864,N_4638,N_4787);
nand U4865 (N_4865,N_4753,N_4729);
nand U4866 (N_4866,N_4704,N_4699);
or U4867 (N_4867,N_4730,N_4642);
nand U4868 (N_4868,N_4713,N_4647);
nand U4869 (N_4869,N_4692,N_4693);
or U4870 (N_4870,N_4697,N_4734);
or U4871 (N_4871,N_4639,N_4755);
and U4872 (N_4872,N_4754,N_4658);
and U4873 (N_4873,N_4684,N_4623);
xor U4874 (N_4874,N_4717,N_4635);
nor U4875 (N_4875,N_4744,N_4656);
nor U4876 (N_4876,N_4741,N_4633);
nor U4877 (N_4877,N_4607,N_4788);
or U4878 (N_4878,N_4721,N_4663);
or U4879 (N_4879,N_4674,N_4776);
nand U4880 (N_4880,N_4764,N_4634);
xnor U4881 (N_4881,N_4767,N_4636);
xnor U4882 (N_4882,N_4799,N_4778);
nor U4883 (N_4883,N_4651,N_4691);
nand U4884 (N_4884,N_4655,N_4731);
or U4885 (N_4885,N_4780,N_4604);
and U4886 (N_4886,N_4662,N_4624);
or U4887 (N_4887,N_4759,N_4723);
or U4888 (N_4888,N_4722,N_4609);
or U4889 (N_4889,N_4671,N_4779);
nand U4890 (N_4890,N_4670,N_4611);
and U4891 (N_4891,N_4792,N_4608);
or U4892 (N_4892,N_4701,N_4715);
nor U4893 (N_4893,N_4728,N_4696);
nand U4894 (N_4894,N_4653,N_4631);
nand U4895 (N_4895,N_4678,N_4770);
nor U4896 (N_4896,N_4645,N_4718);
or U4897 (N_4897,N_4675,N_4648);
or U4898 (N_4898,N_4625,N_4796);
and U4899 (N_4899,N_4613,N_4742);
nand U4900 (N_4900,N_4729,N_4748);
and U4901 (N_4901,N_4621,N_4634);
nand U4902 (N_4902,N_4745,N_4689);
nand U4903 (N_4903,N_4757,N_4731);
nand U4904 (N_4904,N_4714,N_4635);
and U4905 (N_4905,N_4786,N_4766);
and U4906 (N_4906,N_4688,N_4652);
and U4907 (N_4907,N_4776,N_4774);
xnor U4908 (N_4908,N_4602,N_4661);
xor U4909 (N_4909,N_4629,N_4752);
and U4910 (N_4910,N_4727,N_4784);
nor U4911 (N_4911,N_4637,N_4738);
or U4912 (N_4912,N_4794,N_4621);
nor U4913 (N_4913,N_4682,N_4698);
nor U4914 (N_4914,N_4621,N_4765);
nor U4915 (N_4915,N_4713,N_4681);
xor U4916 (N_4916,N_4697,N_4777);
nand U4917 (N_4917,N_4644,N_4759);
nand U4918 (N_4918,N_4609,N_4779);
nor U4919 (N_4919,N_4785,N_4602);
nand U4920 (N_4920,N_4623,N_4786);
xnor U4921 (N_4921,N_4798,N_4739);
or U4922 (N_4922,N_4604,N_4759);
and U4923 (N_4923,N_4639,N_4629);
xnor U4924 (N_4924,N_4648,N_4765);
and U4925 (N_4925,N_4779,N_4711);
xor U4926 (N_4926,N_4602,N_4651);
nand U4927 (N_4927,N_4695,N_4739);
nand U4928 (N_4928,N_4727,N_4685);
or U4929 (N_4929,N_4736,N_4788);
nand U4930 (N_4930,N_4634,N_4648);
or U4931 (N_4931,N_4726,N_4688);
xnor U4932 (N_4932,N_4736,N_4710);
nand U4933 (N_4933,N_4753,N_4731);
nor U4934 (N_4934,N_4786,N_4605);
xnor U4935 (N_4935,N_4773,N_4782);
or U4936 (N_4936,N_4773,N_4668);
and U4937 (N_4937,N_4642,N_4697);
nand U4938 (N_4938,N_4788,N_4716);
xnor U4939 (N_4939,N_4653,N_4629);
nor U4940 (N_4940,N_4622,N_4669);
xnor U4941 (N_4941,N_4653,N_4670);
or U4942 (N_4942,N_4776,N_4685);
or U4943 (N_4943,N_4777,N_4744);
nor U4944 (N_4944,N_4768,N_4663);
nand U4945 (N_4945,N_4614,N_4762);
xor U4946 (N_4946,N_4747,N_4739);
nand U4947 (N_4947,N_4712,N_4622);
or U4948 (N_4948,N_4768,N_4685);
and U4949 (N_4949,N_4799,N_4711);
nand U4950 (N_4950,N_4650,N_4623);
and U4951 (N_4951,N_4677,N_4708);
nor U4952 (N_4952,N_4602,N_4610);
nand U4953 (N_4953,N_4628,N_4650);
xor U4954 (N_4954,N_4679,N_4765);
or U4955 (N_4955,N_4634,N_4733);
and U4956 (N_4956,N_4628,N_4749);
nand U4957 (N_4957,N_4609,N_4683);
xnor U4958 (N_4958,N_4614,N_4681);
nand U4959 (N_4959,N_4769,N_4739);
nand U4960 (N_4960,N_4720,N_4769);
xor U4961 (N_4961,N_4631,N_4695);
nand U4962 (N_4962,N_4763,N_4730);
nand U4963 (N_4963,N_4781,N_4790);
and U4964 (N_4964,N_4668,N_4797);
nand U4965 (N_4965,N_4728,N_4713);
xor U4966 (N_4966,N_4721,N_4660);
or U4967 (N_4967,N_4702,N_4712);
nor U4968 (N_4968,N_4760,N_4739);
and U4969 (N_4969,N_4681,N_4604);
nor U4970 (N_4970,N_4672,N_4784);
or U4971 (N_4971,N_4634,N_4779);
xor U4972 (N_4972,N_4724,N_4754);
nand U4973 (N_4973,N_4747,N_4690);
nor U4974 (N_4974,N_4783,N_4676);
nor U4975 (N_4975,N_4797,N_4782);
nand U4976 (N_4976,N_4696,N_4662);
xor U4977 (N_4977,N_4768,N_4678);
and U4978 (N_4978,N_4710,N_4671);
or U4979 (N_4979,N_4663,N_4624);
xor U4980 (N_4980,N_4752,N_4725);
xnor U4981 (N_4981,N_4648,N_4728);
or U4982 (N_4982,N_4720,N_4700);
xnor U4983 (N_4983,N_4687,N_4668);
xnor U4984 (N_4984,N_4783,N_4632);
nor U4985 (N_4985,N_4631,N_4608);
nand U4986 (N_4986,N_4722,N_4788);
or U4987 (N_4987,N_4678,N_4638);
xor U4988 (N_4988,N_4772,N_4615);
or U4989 (N_4989,N_4725,N_4720);
nand U4990 (N_4990,N_4704,N_4797);
and U4991 (N_4991,N_4747,N_4734);
and U4992 (N_4992,N_4785,N_4696);
and U4993 (N_4993,N_4709,N_4649);
and U4994 (N_4994,N_4774,N_4632);
or U4995 (N_4995,N_4694,N_4689);
or U4996 (N_4996,N_4747,N_4738);
and U4997 (N_4997,N_4678,N_4692);
xnor U4998 (N_4998,N_4794,N_4690);
nand U4999 (N_4999,N_4788,N_4765);
or U5000 (N_5000,N_4824,N_4876);
or U5001 (N_5001,N_4815,N_4888);
nor U5002 (N_5002,N_4895,N_4951);
xnor U5003 (N_5003,N_4896,N_4902);
and U5004 (N_5004,N_4893,N_4991);
nand U5005 (N_5005,N_4899,N_4890);
xor U5006 (N_5006,N_4828,N_4897);
xnor U5007 (N_5007,N_4816,N_4924);
and U5008 (N_5008,N_4849,N_4865);
or U5009 (N_5009,N_4809,N_4805);
or U5010 (N_5010,N_4820,N_4814);
nand U5011 (N_5011,N_4845,N_4878);
nor U5012 (N_5012,N_4974,N_4854);
nand U5013 (N_5013,N_4968,N_4906);
or U5014 (N_5014,N_4887,N_4801);
and U5015 (N_5015,N_4918,N_4871);
or U5016 (N_5016,N_4979,N_4821);
xnor U5017 (N_5017,N_4927,N_4901);
nor U5018 (N_5018,N_4962,N_4905);
and U5019 (N_5019,N_4800,N_4920);
and U5020 (N_5020,N_4853,N_4883);
or U5021 (N_5021,N_4928,N_4898);
nand U5022 (N_5022,N_4836,N_4940);
or U5023 (N_5023,N_4839,N_4998);
and U5024 (N_5024,N_4946,N_4802);
nand U5025 (N_5025,N_4904,N_4818);
nand U5026 (N_5026,N_4808,N_4947);
nor U5027 (N_5027,N_4840,N_4967);
and U5028 (N_5028,N_4811,N_4952);
and U5029 (N_5029,N_4937,N_4838);
or U5030 (N_5030,N_4995,N_4956);
xor U5031 (N_5031,N_4882,N_4949);
nand U5032 (N_5032,N_4914,N_4859);
or U5033 (N_5033,N_4930,N_4870);
and U5034 (N_5034,N_4976,N_4855);
nor U5035 (N_5035,N_4973,N_4866);
nor U5036 (N_5036,N_4972,N_4832);
nor U5037 (N_5037,N_4803,N_4977);
nor U5038 (N_5038,N_4844,N_4997);
nor U5039 (N_5039,N_4965,N_4999);
nor U5040 (N_5040,N_4860,N_4950);
or U5041 (N_5041,N_4915,N_4987);
nand U5042 (N_5042,N_4852,N_4861);
xnor U5043 (N_5043,N_4862,N_4822);
nand U5044 (N_5044,N_4936,N_4830);
and U5045 (N_5045,N_4953,N_4960);
nor U5046 (N_5046,N_4867,N_4982);
or U5047 (N_5047,N_4963,N_4909);
or U5048 (N_5048,N_4858,N_4834);
xor U5049 (N_5049,N_4916,N_4885);
nor U5050 (N_5050,N_4863,N_4938);
nor U5051 (N_5051,N_4857,N_4945);
xor U5052 (N_5052,N_4933,N_4988);
and U5053 (N_5053,N_4819,N_4891);
and U5054 (N_5054,N_4804,N_4907);
nor U5055 (N_5055,N_4913,N_4847);
and U5056 (N_5056,N_4959,N_4978);
or U5057 (N_5057,N_4934,N_4993);
and U5058 (N_5058,N_4990,N_4848);
or U5059 (N_5059,N_4922,N_4833);
xor U5060 (N_5060,N_4986,N_4911);
nand U5061 (N_5061,N_4970,N_4975);
or U5062 (N_5062,N_4881,N_4926);
xnor U5063 (N_5063,N_4932,N_4879);
nand U5064 (N_5064,N_4908,N_4875);
xnor U5065 (N_5065,N_4971,N_4835);
and U5066 (N_5066,N_4964,N_4869);
nand U5067 (N_5067,N_4825,N_4837);
or U5068 (N_5068,N_4826,N_4985);
nor U5069 (N_5069,N_4877,N_4910);
and U5070 (N_5070,N_4892,N_4996);
nand U5071 (N_5071,N_4942,N_4864);
or U5072 (N_5072,N_4884,N_4983);
xnor U5073 (N_5073,N_4827,N_4812);
xnor U5074 (N_5074,N_4900,N_4846);
xor U5075 (N_5075,N_4874,N_4894);
and U5076 (N_5076,N_4813,N_4903);
or U5077 (N_5077,N_4851,N_4980);
xnor U5078 (N_5078,N_4954,N_4931);
nor U5079 (N_5079,N_4806,N_4957);
nand U5080 (N_5080,N_4984,N_4925);
and U5081 (N_5081,N_4955,N_4966);
nand U5082 (N_5082,N_4941,N_4944);
nand U5083 (N_5083,N_4843,N_4886);
xor U5084 (N_5084,N_4856,N_4823);
nor U5085 (N_5085,N_4917,N_4948);
or U5086 (N_5086,N_4989,N_4842);
nand U5087 (N_5087,N_4912,N_4872);
or U5088 (N_5088,N_4810,N_4939);
and U5089 (N_5089,N_4850,N_4981);
and U5090 (N_5090,N_4817,N_4829);
or U5091 (N_5091,N_4994,N_4919);
nand U5092 (N_5092,N_4969,N_4807);
xor U5093 (N_5093,N_4923,N_4873);
nand U5094 (N_5094,N_4868,N_4992);
nor U5095 (N_5095,N_4935,N_4929);
or U5096 (N_5096,N_4961,N_4958);
xnor U5097 (N_5097,N_4921,N_4880);
nor U5098 (N_5098,N_4841,N_4889);
and U5099 (N_5099,N_4943,N_4831);
or U5100 (N_5100,N_4812,N_4990);
nand U5101 (N_5101,N_4834,N_4848);
and U5102 (N_5102,N_4879,N_4892);
nand U5103 (N_5103,N_4804,N_4886);
nand U5104 (N_5104,N_4883,N_4879);
nor U5105 (N_5105,N_4808,N_4994);
xor U5106 (N_5106,N_4992,N_4861);
and U5107 (N_5107,N_4885,N_4861);
or U5108 (N_5108,N_4943,N_4986);
xor U5109 (N_5109,N_4987,N_4875);
nand U5110 (N_5110,N_4886,N_4968);
and U5111 (N_5111,N_4882,N_4995);
nor U5112 (N_5112,N_4991,N_4844);
nor U5113 (N_5113,N_4833,N_4970);
nand U5114 (N_5114,N_4838,N_4856);
and U5115 (N_5115,N_4918,N_4937);
or U5116 (N_5116,N_4809,N_4973);
nand U5117 (N_5117,N_4878,N_4992);
nor U5118 (N_5118,N_4972,N_4960);
nand U5119 (N_5119,N_4876,N_4875);
nand U5120 (N_5120,N_4820,N_4823);
xnor U5121 (N_5121,N_4972,N_4996);
nand U5122 (N_5122,N_4877,N_4980);
nor U5123 (N_5123,N_4905,N_4844);
and U5124 (N_5124,N_4858,N_4978);
nand U5125 (N_5125,N_4859,N_4878);
nand U5126 (N_5126,N_4944,N_4979);
nand U5127 (N_5127,N_4898,N_4831);
nand U5128 (N_5128,N_4805,N_4956);
or U5129 (N_5129,N_4938,N_4987);
and U5130 (N_5130,N_4930,N_4941);
or U5131 (N_5131,N_4881,N_4864);
nand U5132 (N_5132,N_4833,N_4821);
xor U5133 (N_5133,N_4997,N_4968);
xnor U5134 (N_5134,N_4892,N_4979);
nor U5135 (N_5135,N_4943,N_4879);
and U5136 (N_5136,N_4877,N_4833);
xnor U5137 (N_5137,N_4928,N_4945);
nand U5138 (N_5138,N_4902,N_4942);
nand U5139 (N_5139,N_4816,N_4989);
nand U5140 (N_5140,N_4918,N_4882);
nand U5141 (N_5141,N_4933,N_4828);
xnor U5142 (N_5142,N_4814,N_4845);
or U5143 (N_5143,N_4803,N_4926);
and U5144 (N_5144,N_4912,N_4947);
and U5145 (N_5145,N_4965,N_4948);
or U5146 (N_5146,N_4970,N_4838);
nand U5147 (N_5147,N_4977,N_4926);
or U5148 (N_5148,N_4948,N_4995);
xnor U5149 (N_5149,N_4926,N_4801);
nand U5150 (N_5150,N_4938,N_4828);
nand U5151 (N_5151,N_4840,N_4906);
or U5152 (N_5152,N_4856,N_4976);
xor U5153 (N_5153,N_4859,N_4983);
nand U5154 (N_5154,N_4910,N_4826);
nand U5155 (N_5155,N_4815,N_4802);
xnor U5156 (N_5156,N_4949,N_4912);
or U5157 (N_5157,N_4971,N_4927);
nor U5158 (N_5158,N_4821,N_4859);
nand U5159 (N_5159,N_4928,N_4818);
or U5160 (N_5160,N_4930,N_4981);
and U5161 (N_5161,N_4903,N_4802);
nor U5162 (N_5162,N_4809,N_4934);
nand U5163 (N_5163,N_4965,N_4987);
and U5164 (N_5164,N_4940,N_4895);
nand U5165 (N_5165,N_4970,N_4969);
xor U5166 (N_5166,N_4824,N_4804);
nand U5167 (N_5167,N_4819,N_4928);
nor U5168 (N_5168,N_4965,N_4956);
nor U5169 (N_5169,N_4825,N_4935);
nor U5170 (N_5170,N_4889,N_4984);
or U5171 (N_5171,N_4947,N_4924);
xnor U5172 (N_5172,N_4901,N_4824);
nor U5173 (N_5173,N_4994,N_4861);
nand U5174 (N_5174,N_4857,N_4978);
and U5175 (N_5175,N_4864,N_4919);
xor U5176 (N_5176,N_4806,N_4852);
nand U5177 (N_5177,N_4819,N_4925);
or U5178 (N_5178,N_4871,N_4955);
and U5179 (N_5179,N_4894,N_4973);
and U5180 (N_5180,N_4925,N_4935);
nand U5181 (N_5181,N_4995,N_4908);
or U5182 (N_5182,N_4870,N_4943);
or U5183 (N_5183,N_4988,N_4941);
and U5184 (N_5184,N_4925,N_4855);
and U5185 (N_5185,N_4962,N_4990);
nor U5186 (N_5186,N_4843,N_4912);
or U5187 (N_5187,N_4852,N_4825);
or U5188 (N_5188,N_4833,N_4897);
xnor U5189 (N_5189,N_4898,N_4911);
xor U5190 (N_5190,N_4964,N_4998);
nor U5191 (N_5191,N_4936,N_4801);
or U5192 (N_5192,N_4825,N_4905);
xnor U5193 (N_5193,N_4852,N_4888);
nor U5194 (N_5194,N_4974,N_4992);
nand U5195 (N_5195,N_4842,N_4866);
nand U5196 (N_5196,N_4901,N_4964);
xnor U5197 (N_5197,N_4926,N_4847);
xor U5198 (N_5198,N_4802,N_4929);
xnor U5199 (N_5199,N_4955,N_4801);
nand U5200 (N_5200,N_5108,N_5016);
nor U5201 (N_5201,N_5196,N_5177);
nor U5202 (N_5202,N_5048,N_5129);
and U5203 (N_5203,N_5059,N_5098);
nor U5204 (N_5204,N_5037,N_5142);
and U5205 (N_5205,N_5044,N_5136);
xor U5206 (N_5206,N_5124,N_5138);
nand U5207 (N_5207,N_5058,N_5022);
and U5208 (N_5208,N_5085,N_5112);
or U5209 (N_5209,N_5121,N_5091);
or U5210 (N_5210,N_5027,N_5053);
or U5211 (N_5211,N_5092,N_5135);
nand U5212 (N_5212,N_5070,N_5102);
nand U5213 (N_5213,N_5054,N_5150);
xnor U5214 (N_5214,N_5090,N_5103);
or U5215 (N_5215,N_5012,N_5191);
nor U5216 (N_5216,N_5179,N_5021);
xor U5217 (N_5217,N_5107,N_5080);
nor U5218 (N_5218,N_5197,N_5097);
or U5219 (N_5219,N_5031,N_5141);
nor U5220 (N_5220,N_5050,N_5189);
nor U5221 (N_5221,N_5167,N_5006);
xor U5222 (N_5222,N_5030,N_5187);
nor U5223 (N_5223,N_5019,N_5083);
nand U5224 (N_5224,N_5106,N_5130);
xor U5225 (N_5225,N_5005,N_5077);
and U5226 (N_5226,N_5143,N_5152);
nor U5227 (N_5227,N_5011,N_5133);
and U5228 (N_5228,N_5056,N_5109);
xor U5229 (N_5229,N_5008,N_5188);
nand U5230 (N_5230,N_5115,N_5029);
nor U5231 (N_5231,N_5186,N_5182);
and U5232 (N_5232,N_5120,N_5162);
and U5233 (N_5233,N_5176,N_5153);
and U5234 (N_5234,N_5057,N_5064);
and U5235 (N_5235,N_5013,N_5066);
nor U5236 (N_5236,N_5194,N_5084);
nor U5237 (N_5237,N_5158,N_5146);
xor U5238 (N_5238,N_5018,N_5192);
or U5239 (N_5239,N_5072,N_5000);
nor U5240 (N_5240,N_5122,N_5126);
xnor U5241 (N_5241,N_5104,N_5052);
xor U5242 (N_5242,N_5161,N_5026);
and U5243 (N_5243,N_5079,N_5172);
and U5244 (N_5244,N_5131,N_5045);
xor U5245 (N_5245,N_5028,N_5035);
nor U5246 (N_5246,N_5055,N_5125);
xnor U5247 (N_5247,N_5137,N_5139);
nand U5248 (N_5248,N_5081,N_5199);
nor U5249 (N_5249,N_5051,N_5170);
nor U5250 (N_5250,N_5003,N_5039);
xor U5251 (N_5251,N_5165,N_5068);
nor U5252 (N_5252,N_5195,N_5060);
or U5253 (N_5253,N_5157,N_5183);
nand U5254 (N_5254,N_5010,N_5149);
or U5255 (N_5255,N_5134,N_5069);
xor U5256 (N_5256,N_5113,N_5078);
or U5257 (N_5257,N_5042,N_5144);
nor U5258 (N_5258,N_5096,N_5111);
or U5259 (N_5259,N_5047,N_5178);
xnor U5260 (N_5260,N_5190,N_5118);
nand U5261 (N_5261,N_5036,N_5156);
or U5262 (N_5262,N_5004,N_5105);
xnor U5263 (N_5263,N_5065,N_5095);
xor U5264 (N_5264,N_5099,N_5128);
nand U5265 (N_5265,N_5063,N_5087);
or U5266 (N_5266,N_5094,N_5015);
and U5267 (N_5267,N_5074,N_5034);
and U5268 (N_5268,N_5132,N_5155);
nand U5269 (N_5269,N_5151,N_5020);
xnor U5270 (N_5270,N_5171,N_5088);
nor U5271 (N_5271,N_5007,N_5127);
nor U5272 (N_5272,N_5154,N_5169);
or U5273 (N_5273,N_5180,N_5086);
nand U5274 (N_5274,N_5145,N_5025);
nor U5275 (N_5275,N_5017,N_5076);
or U5276 (N_5276,N_5093,N_5173);
nand U5277 (N_5277,N_5009,N_5116);
xnor U5278 (N_5278,N_5123,N_5001);
nor U5279 (N_5279,N_5175,N_5163);
or U5280 (N_5280,N_5023,N_5160);
and U5281 (N_5281,N_5061,N_5164);
nand U5282 (N_5282,N_5114,N_5089);
nor U5283 (N_5283,N_5071,N_5148);
nand U5284 (N_5284,N_5166,N_5075);
or U5285 (N_5285,N_5100,N_5140);
nor U5286 (N_5286,N_5073,N_5185);
or U5287 (N_5287,N_5117,N_5043);
or U5288 (N_5288,N_5049,N_5184);
nand U5289 (N_5289,N_5024,N_5159);
nand U5290 (N_5290,N_5002,N_5082);
and U5291 (N_5291,N_5101,N_5014);
and U5292 (N_5292,N_5067,N_5181);
and U5293 (N_5293,N_5168,N_5174);
xor U5294 (N_5294,N_5193,N_5147);
xnor U5295 (N_5295,N_5110,N_5046);
nand U5296 (N_5296,N_5032,N_5040);
and U5297 (N_5297,N_5119,N_5198);
or U5298 (N_5298,N_5038,N_5062);
xor U5299 (N_5299,N_5041,N_5033);
or U5300 (N_5300,N_5167,N_5192);
or U5301 (N_5301,N_5191,N_5167);
nand U5302 (N_5302,N_5103,N_5189);
nor U5303 (N_5303,N_5025,N_5157);
xor U5304 (N_5304,N_5139,N_5007);
and U5305 (N_5305,N_5033,N_5053);
nor U5306 (N_5306,N_5105,N_5035);
nor U5307 (N_5307,N_5137,N_5111);
nand U5308 (N_5308,N_5189,N_5166);
or U5309 (N_5309,N_5148,N_5040);
nor U5310 (N_5310,N_5069,N_5050);
or U5311 (N_5311,N_5077,N_5134);
nand U5312 (N_5312,N_5084,N_5092);
nand U5313 (N_5313,N_5012,N_5043);
or U5314 (N_5314,N_5059,N_5166);
and U5315 (N_5315,N_5037,N_5119);
xnor U5316 (N_5316,N_5067,N_5162);
nand U5317 (N_5317,N_5022,N_5124);
and U5318 (N_5318,N_5152,N_5122);
or U5319 (N_5319,N_5135,N_5074);
nor U5320 (N_5320,N_5122,N_5129);
nor U5321 (N_5321,N_5136,N_5021);
xnor U5322 (N_5322,N_5048,N_5051);
xor U5323 (N_5323,N_5182,N_5050);
xnor U5324 (N_5324,N_5101,N_5172);
or U5325 (N_5325,N_5069,N_5122);
and U5326 (N_5326,N_5140,N_5026);
nand U5327 (N_5327,N_5055,N_5038);
xnor U5328 (N_5328,N_5048,N_5054);
nor U5329 (N_5329,N_5088,N_5188);
and U5330 (N_5330,N_5081,N_5046);
and U5331 (N_5331,N_5195,N_5049);
nor U5332 (N_5332,N_5073,N_5135);
or U5333 (N_5333,N_5097,N_5092);
nand U5334 (N_5334,N_5164,N_5118);
nor U5335 (N_5335,N_5183,N_5015);
or U5336 (N_5336,N_5042,N_5139);
and U5337 (N_5337,N_5113,N_5082);
or U5338 (N_5338,N_5039,N_5164);
or U5339 (N_5339,N_5156,N_5087);
and U5340 (N_5340,N_5057,N_5087);
or U5341 (N_5341,N_5191,N_5063);
nand U5342 (N_5342,N_5141,N_5073);
nand U5343 (N_5343,N_5070,N_5176);
xnor U5344 (N_5344,N_5035,N_5175);
xor U5345 (N_5345,N_5052,N_5038);
and U5346 (N_5346,N_5190,N_5074);
or U5347 (N_5347,N_5122,N_5154);
and U5348 (N_5348,N_5098,N_5091);
or U5349 (N_5349,N_5009,N_5137);
or U5350 (N_5350,N_5059,N_5013);
or U5351 (N_5351,N_5071,N_5129);
or U5352 (N_5352,N_5130,N_5070);
xnor U5353 (N_5353,N_5149,N_5186);
xor U5354 (N_5354,N_5127,N_5155);
or U5355 (N_5355,N_5179,N_5005);
or U5356 (N_5356,N_5156,N_5042);
and U5357 (N_5357,N_5142,N_5081);
or U5358 (N_5358,N_5083,N_5030);
xnor U5359 (N_5359,N_5076,N_5176);
or U5360 (N_5360,N_5187,N_5137);
nor U5361 (N_5361,N_5185,N_5095);
nand U5362 (N_5362,N_5137,N_5164);
nor U5363 (N_5363,N_5147,N_5022);
and U5364 (N_5364,N_5087,N_5163);
or U5365 (N_5365,N_5150,N_5099);
xnor U5366 (N_5366,N_5164,N_5147);
or U5367 (N_5367,N_5086,N_5037);
or U5368 (N_5368,N_5101,N_5092);
or U5369 (N_5369,N_5017,N_5068);
and U5370 (N_5370,N_5140,N_5023);
nand U5371 (N_5371,N_5144,N_5143);
or U5372 (N_5372,N_5176,N_5164);
xnor U5373 (N_5373,N_5137,N_5199);
xor U5374 (N_5374,N_5082,N_5128);
or U5375 (N_5375,N_5114,N_5060);
and U5376 (N_5376,N_5167,N_5021);
or U5377 (N_5377,N_5089,N_5145);
nand U5378 (N_5378,N_5104,N_5107);
and U5379 (N_5379,N_5129,N_5013);
xnor U5380 (N_5380,N_5069,N_5142);
xnor U5381 (N_5381,N_5138,N_5028);
nand U5382 (N_5382,N_5037,N_5004);
and U5383 (N_5383,N_5053,N_5076);
nor U5384 (N_5384,N_5046,N_5104);
nor U5385 (N_5385,N_5140,N_5135);
nand U5386 (N_5386,N_5188,N_5079);
nand U5387 (N_5387,N_5165,N_5071);
and U5388 (N_5388,N_5124,N_5158);
or U5389 (N_5389,N_5042,N_5198);
and U5390 (N_5390,N_5105,N_5166);
nand U5391 (N_5391,N_5156,N_5192);
or U5392 (N_5392,N_5062,N_5026);
nor U5393 (N_5393,N_5096,N_5163);
or U5394 (N_5394,N_5054,N_5076);
and U5395 (N_5395,N_5055,N_5058);
nand U5396 (N_5396,N_5111,N_5142);
xor U5397 (N_5397,N_5147,N_5183);
nor U5398 (N_5398,N_5156,N_5124);
nand U5399 (N_5399,N_5039,N_5092);
xnor U5400 (N_5400,N_5370,N_5254);
and U5401 (N_5401,N_5276,N_5389);
or U5402 (N_5402,N_5343,N_5341);
and U5403 (N_5403,N_5204,N_5352);
xnor U5404 (N_5404,N_5248,N_5252);
or U5405 (N_5405,N_5292,N_5260);
nor U5406 (N_5406,N_5388,N_5360);
nor U5407 (N_5407,N_5259,N_5322);
and U5408 (N_5408,N_5369,N_5330);
nor U5409 (N_5409,N_5217,N_5349);
nor U5410 (N_5410,N_5226,N_5235);
nand U5411 (N_5411,N_5263,N_5396);
nand U5412 (N_5412,N_5220,N_5347);
or U5413 (N_5413,N_5209,N_5211);
nand U5414 (N_5414,N_5356,N_5309);
and U5415 (N_5415,N_5261,N_5355);
xor U5416 (N_5416,N_5326,N_5201);
and U5417 (N_5417,N_5375,N_5223);
and U5418 (N_5418,N_5218,N_5277);
or U5419 (N_5419,N_5214,N_5271);
or U5420 (N_5420,N_5284,N_5222);
and U5421 (N_5421,N_5288,N_5257);
and U5422 (N_5422,N_5390,N_5212);
nand U5423 (N_5423,N_5240,N_5242);
and U5424 (N_5424,N_5304,N_5364);
xor U5425 (N_5425,N_5300,N_5287);
or U5426 (N_5426,N_5342,N_5251);
or U5427 (N_5427,N_5381,N_5250);
xor U5428 (N_5428,N_5238,N_5306);
or U5429 (N_5429,N_5397,N_5382);
and U5430 (N_5430,N_5282,N_5331);
and U5431 (N_5431,N_5358,N_5395);
nor U5432 (N_5432,N_5233,N_5392);
xor U5433 (N_5433,N_5279,N_5350);
nand U5434 (N_5434,N_5387,N_5371);
and U5435 (N_5435,N_5264,N_5362);
nor U5436 (N_5436,N_5312,N_5307);
and U5437 (N_5437,N_5268,N_5359);
and U5438 (N_5438,N_5372,N_5286);
nand U5439 (N_5439,N_5200,N_5267);
nor U5440 (N_5440,N_5269,N_5230);
xnor U5441 (N_5441,N_5353,N_5344);
nand U5442 (N_5442,N_5376,N_5225);
or U5443 (N_5443,N_5354,N_5329);
nor U5444 (N_5444,N_5310,N_5208);
and U5445 (N_5445,N_5272,N_5265);
or U5446 (N_5446,N_5219,N_5386);
or U5447 (N_5447,N_5302,N_5246);
nand U5448 (N_5448,N_5320,N_5294);
and U5449 (N_5449,N_5202,N_5351);
or U5450 (N_5450,N_5262,N_5256);
or U5451 (N_5451,N_5270,N_5399);
nor U5452 (N_5452,N_5346,N_5335);
or U5453 (N_5453,N_5290,N_5237);
nor U5454 (N_5454,N_5241,N_5232);
and U5455 (N_5455,N_5236,N_5316);
or U5456 (N_5456,N_5303,N_5377);
nor U5457 (N_5457,N_5273,N_5361);
and U5458 (N_5458,N_5244,N_5365);
nand U5459 (N_5459,N_5301,N_5357);
xnor U5460 (N_5460,N_5274,N_5367);
nor U5461 (N_5461,N_5337,N_5207);
xor U5462 (N_5462,N_5228,N_5332);
xnor U5463 (N_5463,N_5229,N_5366);
or U5464 (N_5464,N_5317,N_5391);
and U5465 (N_5465,N_5368,N_5280);
or U5466 (N_5466,N_5323,N_5224);
or U5467 (N_5467,N_5385,N_5333);
or U5468 (N_5468,N_5278,N_5339);
nor U5469 (N_5469,N_5311,N_5319);
or U5470 (N_5470,N_5345,N_5383);
nand U5471 (N_5471,N_5253,N_5336);
or U5472 (N_5472,N_5215,N_5231);
xnor U5473 (N_5473,N_5308,N_5293);
nor U5474 (N_5474,N_5379,N_5318);
nor U5475 (N_5475,N_5394,N_5213);
xnor U5476 (N_5476,N_5239,N_5393);
nor U5477 (N_5477,N_5289,N_5299);
or U5478 (N_5478,N_5321,N_5243);
and U5479 (N_5479,N_5285,N_5314);
nor U5480 (N_5480,N_5297,N_5340);
nand U5481 (N_5481,N_5283,N_5373);
nand U5482 (N_5482,N_5315,N_5334);
and U5483 (N_5483,N_5206,N_5281);
or U5484 (N_5484,N_5398,N_5324);
xnor U5485 (N_5485,N_5363,N_5221);
nor U5486 (N_5486,N_5227,N_5210);
nor U5487 (N_5487,N_5313,N_5205);
or U5488 (N_5488,N_5328,N_5374);
and U5489 (N_5489,N_5291,N_5384);
or U5490 (N_5490,N_5216,N_5295);
or U5491 (N_5491,N_5203,N_5380);
nand U5492 (N_5492,N_5348,N_5247);
or U5493 (N_5493,N_5338,N_5296);
nor U5494 (N_5494,N_5245,N_5266);
or U5495 (N_5495,N_5378,N_5298);
xor U5496 (N_5496,N_5255,N_5249);
xor U5497 (N_5497,N_5327,N_5275);
xnor U5498 (N_5498,N_5325,N_5258);
and U5499 (N_5499,N_5234,N_5305);
or U5500 (N_5500,N_5290,N_5370);
or U5501 (N_5501,N_5381,N_5355);
or U5502 (N_5502,N_5247,N_5397);
xnor U5503 (N_5503,N_5230,N_5379);
nand U5504 (N_5504,N_5306,N_5286);
xnor U5505 (N_5505,N_5246,N_5299);
and U5506 (N_5506,N_5379,N_5330);
and U5507 (N_5507,N_5360,N_5357);
or U5508 (N_5508,N_5293,N_5212);
xnor U5509 (N_5509,N_5372,N_5231);
nor U5510 (N_5510,N_5354,N_5303);
nand U5511 (N_5511,N_5351,N_5205);
xnor U5512 (N_5512,N_5275,N_5205);
nand U5513 (N_5513,N_5251,N_5378);
or U5514 (N_5514,N_5322,N_5378);
xor U5515 (N_5515,N_5221,N_5365);
or U5516 (N_5516,N_5314,N_5351);
xnor U5517 (N_5517,N_5293,N_5222);
and U5518 (N_5518,N_5386,N_5277);
or U5519 (N_5519,N_5295,N_5236);
nand U5520 (N_5520,N_5215,N_5279);
nor U5521 (N_5521,N_5330,N_5288);
nand U5522 (N_5522,N_5300,N_5285);
or U5523 (N_5523,N_5272,N_5380);
nor U5524 (N_5524,N_5385,N_5398);
nand U5525 (N_5525,N_5384,N_5217);
nor U5526 (N_5526,N_5319,N_5363);
nor U5527 (N_5527,N_5209,N_5363);
nand U5528 (N_5528,N_5232,N_5252);
xor U5529 (N_5529,N_5398,N_5254);
nand U5530 (N_5530,N_5281,N_5224);
nand U5531 (N_5531,N_5251,N_5236);
and U5532 (N_5532,N_5247,N_5227);
nor U5533 (N_5533,N_5225,N_5310);
or U5534 (N_5534,N_5286,N_5327);
or U5535 (N_5535,N_5263,N_5231);
xor U5536 (N_5536,N_5325,N_5242);
nor U5537 (N_5537,N_5340,N_5365);
nor U5538 (N_5538,N_5394,N_5352);
and U5539 (N_5539,N_5363,N_5200);
nor U5540 (N_5540,N_5277,N_5321);
nand U5541 (N_5541,N_5286,N_5281);
or U5542 (N_5542,N_5288,N_5328);
or U5543 (N_5543,N_5360,N_5200);
nor U5544 (N_5544,N_5273,N_5263);
and U5545 (N_5545,N_5217,N_5345);
or U5546 (N_5546,N_5300,N_5341);
or U5547 (N_5547,N_5363,N_5394);
and U5548 (N_5548,N_5260,N_5270);
xor U5549 (N_5549,N_5328,N_5245);
nand U5550 (N_5550,N_5287,N_5339);
xnor U5551 (N_5551,N_5228,N_5273);
nor U5552 (N_5552,N_5228,N_5296);
nand U5553 (N_5553,N_5203,N_5361);
or U5554 (N_5554,N_5316,N_5201);
and U5555 (N_5555,N_5208,N_5281);
nor U5556 (N_5556,N_5312,N_5213);
and U5557 (N_5557,N_5390,N_5264);
or U5558 (N_5558,N_5344,N_5327);
and U5559 (N_5559,N_5342,N_5285);
or U5560 (N_5560,N_5361,N_5256);
and U5561 (N_5561,N_5296,N_5394);
xnor U5562 (N_5562,N_5359,N_5319);
nor U5563 (N_5563,N_5236,N_5384);
nor U5564 (N_5564,N_5308,N_5256);
nand U5565 (N_5565,N_5356,N_5394);
or U5566 (N_5566,N_5301,N_5314);
xnor U5567 (N_5567,N_5298,N_5386);
nor U5568 (N_5568,N_5344,N_5263);
and U5569 (N_5569,N_5241,N_5312);
nand U5570 (N_5570,N_5212,N_5317);
xor U5571 (N_5571,N_5316,N_5265);
nor U5572 (N_5572,N_5345,N_5307);
or U5573 (N_5573,N_5306,N_5347);
nor U5574 (N_5574,N_5311,N_5378);
xor U5575 (N_5575,N_5343,N_5393);
and U5576 (N_5576,N_5243,N_5376);
nand U5577 (N_5577,N_5370,N_5390);
xnor U5578 (N_5578,N_5291,N_5216);
xor U5579 (N_5579,N_5209,N_5226);
and U5580 (N_5580,N_5386,N_5295);
xor U5581 (N_5581,N_5359,N_5349);
nor U5582 (N_5582,N_5334,N_5292);
nand U5583 (N_5583,N_5293,N_5270);
or U5584 (N_5584,N_5354,N_5290);
or U5585 (N_5585,N_5374,N_5217);
xor U5586 (N_5586,N_5232,N_5399);
xor U5587 (N_5587,N_5328,N_5280);
nor U5588 (N_5588,N_5327,N_5265);
nor U5589 (N_5589,N_5261,N_5393);
nand U5590 (N_5590,N_5311,N_5323);
nand U5591 (N_5591,N_5297,N_5312);
nor U5592 (N_5592,N_5390,N_5379);
or U5593 (N_5593,N_5217,N_5318);
or U5594 (N_5594,N_5294,N_5220);
or U5595 (N_5595,N_5208,N_5269);
nor U5596 (N_5596,N_5248,N_5398);
xnor U5597 (N_5597,N_5325,N_5393);
or U5598 (N_5598,N_5333,N_5310);
and U5599 (N_5599,N_5310,N_5294);
nand U5600 (N_5600,N_5586,N_5415);
or U5601 (N_5601,N_5482,N_5401);
nor U5602 (N_5602,N_5511,N_5486);
nand U5603 (N_5603,N_5558,N_5460);
xor U5604 (N_5604,N_5456,N_5520);
xor U5605 (N_5605,N_5425,N_5561);
and U5606 (N_5606,N_5458,N_5419);
xnor U5607 (N_5607,N_5515,N_5470);
nor U5608 (N_5608,N_5573,N_5473);
and U5609 (N_5609,N_5525,N_5542);
nand U5610 (N_5610,N_5541,N_5469);
nor U5611 (N_5611,N_5567,N_5403);
or U5612 (N_5612,N_5509,N_5557);
or U5613 (N_5613,N_5537,N_5487);
and U5614 (N_5614,N_5568,N_5516);
or U5615 (N_5615,N_5485,N_5582);
nand U5616 (N_5616,N_5451,N_5570);
xnor U5617 (N_5617,N_5575,N_5472);
xor U5618 (N_5618,N_5497,N_5481);
nand U5619 (N_5619,N_5414,N_5423);
nand U5620 (N_5620,N_5556,N_5409);
or U5621 (N_5621,N_5534,N_5440);
nand U5622 (N_5622,N_5416,N_5547);
nand U5623 (N_5623,N_5549,N_5554);
or U5624 (N_5624,N_5421,N_5464);
or U5625 (N_5625,N_5408,N_5592);
and U5626 (N_5626,N_5426,N_5475);
nand U5627 (N_5627,N_5533,N_5591);
or U5628 (N_5628,N_5430,N_5531);
nor U5629 (N_5629,N_5590,N_5406);
xor U5630 (N_5630,N_5495,N_5468);
xnor U5631 (N_5631,N_5407,N_5536);
xnor U5632 (N_5632,N_5597,N_5502);
xor U5633 (N_5633,N_5506,N_5523);
xnor U5634 (N_5634,N_5429,N_5553);
xor U5635 (N_5635,N_5545,N_5513);
or U5636 (N_5636,N_5550,N_5500);
nand U5637 (N_5637,N_5462,N_5574);
or U5638 (N_5638,N_5484,N_5461);
or U5639 (N_5639,N_5422,N_5587);
nand U5640 (N_5640,N_5552,N_5455);
nor U5641 (N_5641,N_5512,N_5427);
nand U5642 (N_5642,N_5585,N_5593);
nor U5643 (N_5643,N_5527,N_5524);
xor U5644 (N_5644,N_5420,N_5435);
nor U5645 (N_5645,N_5504,N_5476);
xor U5646 (N_5646,N_5563,N_5599);
nor U5647 (N_5647,N_5596,N_5565);
nand U5648 (N_5648,N_5471,N_5442);
or U5649 (N_5649,N_5494,N_5595);
or U5650 (N_5650,N_5438,N_5457);
xor U5651 (N_5651,N_5480,N_5463);
nand U5652 (N_5652,N_5560,N_5410);
nor U5653 (N_5653,N_5579,N_5514);
nor U5654 (N_5654,N_5483,N_5432);
nor U5655 (N_5655,N_5535,N_5503);
or U5656 (N_5656,N_5402,N_5443);
and U5657 (N_5657,N_5418,N_5564);
nand U5658 (N_5658,N_5433,N_5530);
xor U5659 (N_5659,N_5400,N_5517);
nor U5660 (N_5660,N_5526,N_5439);
or U5661 (N_5661,N_5584,N_5546);
xor U5662 (N_5662,N_5583,N_5447);
xor U5663 (N_5663,N_5405,N_5507);
nand U5664 (N_5664,N_5572,N_5488);
nor U5665 (N_5665,N_5580,N_5539);
nand U5666 (N_5666,N_5522,N_5478);
and U5667 (N_5667,N_5413,N_5519);
and U5668 (N_5668,N_5551,N_5446);
and U5669 (N_5669,N_5412,N_5559);
or U5670 (N_5670,N_5538,N_5465);
nand U5671 (N_5671,N_5467,N_5577);
or U5672 (N_5672,N_5459,N_5581);
and U5673 (N_5673,N_5417,N_5449);
xnor U5674 (N_5674,N_5445,N_5466);
or U5675 (N_5675,N_5431,N_5444);
xnor U5676 (N_5676,N_5428,N_5543);
and U5677 (N_5677,N_5404,N_5411);
or U5678 (N_5678,N_5540,N_5498);
nand U5679 (N_5679,N_5424,N_5529);
and U5680 (N_5680,N_5491,N_5493);
xnor U5681 (N_5681,N_5548,N_5578);
nor U5682 (N_5682,N_5588,N_5594);
or U5683 (N_5683,N_5452,N_5555);
or U5684 (N_5684,N_5598,N_5450);
or U5685 (N_5685,N_5436,N_5448);
or U5686 (N_5686,N_5571,N_5518);
or U5687 (N_5687,N_5544,N_5441);
or U5688 (N_5688,N_5490,N_5453);
nor U5689 (N_5689,N_5510,N_5477);
nand U5690 (N_5690,N_5505,N_5521);
or U5691 (N_5691,N_5528,N_5499);
and U5692 (N_5692,N_5562,N_5492);
or U5693 (N_5693,N_5479,N_5454);
nor U5694 (N_5694,N_5508,N_5566);
xnor U5695 (N_5695,N_5489,N_5569);
and U5696 (N_5696,N_5496,N_5532);
and U5697 (N_5697,N_5474,N_5437);
and U5698 (N_5698,N_5576,N_5501);
nor U5699 (N_5699,N_5434,N_5589);
or U5700 (N_5700,N_5469,N_5484);
or U5701 (N_5701,N_5455,N_5457);
and U5702 (N_5702,N_5462,N_5529);
or U5703 (N_5703,N_5504,N_5427);
nor U5704 (N_5704,N_5492,N_5495);
xnor U5705 (N_5705,N_5443,N_5540);
nand U5706 (N_5706,N_5463,N_5457);
xnor U5707 (N_5707,N_5465,N_5460);
nand U5708 (N_5708,N_5530,N_5561);
xor U5709 (N_5709,N_5448,N_5527);
or U5710 (N_5710,N_5597,N_5511);
or U5711 (N_5711,N_5444,N_5533);
and U5712 (N_5712,N_5541,N_5508);
nand U5713 (N_5713,N_5430,N_5447);
nor U5714 (N_5714,N_5586,N_5539);
or U5715 (N_5715,N_5588,N_5472);
xnor U5716 (N_5716,N_5467,N_5491);
xnor U5717 (N_5717,N_5484,N_5525);
or U5718 (N_5718,N_5565,N_5534);
nor U5719 (N_5719,N_5425,N_5597);
nor U5720 (N_5720,N_5453,N_5541);
and U5721 (N_5721,N_5520,N_5469);
xnor U5722 (N_5722,N_5463,N_5559);
and U5723 (N_5723,N_5446,N_5424);
xor U5724 (N_5724,N_5511,N_5438);
nor U5725 (N_5725,N_5476,N_5553);
nor U5726 (N_5726,N_5403,N_5466);
nand U5727 (N_5727,N_5531,N_5466);
nand U5728 (N_5728,N_5596,N_5444);
nand U5729 (N_5729,N_5446,N_5420);
and U5730 (N_5730,N_5497,N_5454);
xnor U5731 (N_5731,N_5408,N_5577);
and U5732 (N_5732,N_5560,N_5513);
or U5733 (N_5733,N_5462,N_5581);
or U5734 (N_5734,N_5467,N_5514);
nor U5735 (N_5735,N_5510,N_5550);
nor U5736 (N_5736,N_5414,N_5437);
nor U5737 (N_5737,N_5512,N_5433);
nor U5738 (N_5738,N_5402,N_5571);
xnor U5739 (N_5739,N_5434,N_5497);
nor U5740 (N_5740,N_5405,N_5414);
nand U5741 (N_5741,N_5515,N_5546);
or U5742 (N_5742,N_5577,N_5426);
and U5743 (N_5743,N_5579,N_5559);
nor U5744 (N_5744,N_5569,N_5401);
nand U5745 (N_5745,N_5529,N_5496);
xor U5746 (N_5746,N_5501,N_5516);
and U5747 (N_5747,N_5421,N_5422);
xor U5748 (N_5748,N_5520,N_5412);
xnor U5749 (N_5749,N_5534,N_5424);
or U5750 (N_5750,N_5496,N_5412);
nor U5751 (N_5751,N_5465,N_5530);
nor U5752 (N_5752,N_5594,N_5491);
nor U5753 (N_5753,N_5504,N_5410);
or U5754 (N_5754,N_5476,N_5550);
nor U5755 (N_5755,N_5522,N_5463);
and U5756 (N_5756,N_5419,N_5407);
and U5757 (N_5757,N_5400,N_5454);
xor U5758 (N_5758,N_5599,N_5451);
or U5759 (N_5759,N_5438,N_5503);
and U5760 (N_5760,N_5425,N_5592);
or U5761 (N_5761,N_5546,N_5474);
nor U5762 (N_5762,N_5599,N_5473);
or U5763 (N_5763,N_5568,N_5515);
nor U5764 (N_5764,N_5473,N_5471);
or U5765 (N_5765,N_5592,N_5470);
nor U5766 (N_5766,N_5450,N_5585);
and U5767 (N_5767,N_5570,N_5546);
xnor U5768 (N_5768,N_5589,N_5591);
or U5769 (N_5769,N_5506,N_5470);
or U5770 (N_5770,N_5465,N_5534);
nand U5771 (N_5771,N_5545,N_5428);
xnor U5772 (N_5772,N_5447,N_5461);
nand U5773 (N_5773,N_5490,N_5464);
nand U5774 (N_5774,N_5584,N_5583);
or U5775 (N_5775,N_5499,N_5457);
nor U5776 (N_5776,N_5419,N_5520);
and U5777 (N_5777,N_5406,N_5428);
or U5778 (N_5778,N_5443,N_5556);
and U5779 (N_5779,N_5457,N_5459);
nand U5780 (N_5780,N_5599,N_5404);
or U5781 (N_5781,N_5505,N_5402);
nor U5782 (N_5782,N_5496,N_5485);
or U5783 (N_5783,N_5467,N_5419);
xnor U5784 (N_5784,N_5472,N_5493);
xnor U5785 (N_5785,N_5417,N_5568);
or U5786 (N_5786,N_5472,N_5596);
nor U5787 (N_5787,N_5477,N_5481);
nor U5788 (N_5788,N_5575,N_5457);
xnor U5789 (N_5789,N_5485,N_5547);
nor U5790 (N_5790,N_5407,N_5598);
or U5791 (N_5791,N_5452,N_5549);
and U5792 (N_5792,N_5501,N_5570);
xnor U5793 (N_5793,N_5512,N_5406);
or U5794 (N_5794,N_5465,N_5514);
nand U5795 (N_5795,N_5405,N_5553);
or U5796 (N_5796,N_5500,N_5470);
nor U5797 (N_5797,N_5432,N_5544);
nand U5798 (N_5798,N_5416,N_5441);
xor U5799 (N_5799,N_5404,N_5589);
and U5800 (N_5800,N_5611,N_5651);
or U5801 (N_5801,N_5739,N_5682);
nand U5802 (N_5802,N_5796,N_5631);
nand U5803 (N_5803,N_5795,N_5637);
and U5804 (N_5804,N_5767,N_5718);
and U5805 (N_5805,N_5766,N_5799);
nand U5806 (N_5806,N_5632,N_5711);
xnor U5807 (N_5807,N_5636,N_5649);
and U5808 (N_5808,N_5645,N_5797);
xor U5809 (N_5809,N_5701,N_5624);
nand U5810 (N_5810,N_5757,N_5613);
nand U5811 (N_5811,N_5657,N_5748);
xnor U5812 (N_5812,N_5740,N_5686);
or U5813 (N_5813,N_5627,N_5689);
xnor U5814 (N_5814,N_5623,N_5702);
and U5815 (N_5815,N_5704,N_5736);
and U5816 (N_5816,N_5693,N_5674);
nand U5817 (N_5817,N_5776,N_5699);
nand U5818 (N_5818,N_5724,N_5610);
or U5819 (N_5819,N_5644,N_5625);
or U5820 (N_5820,N_5738,N_5786);
nand U5821 (N_5821,N_5727,N_5607);
and U5822 (N_5822,N_5703,N_5617);
xor U5823 (N_5823,N_5681,N_5665);
or U5824 (N_5824,N_5714,N_5603);
or U5825 (N_5825,N_5609,N_5654);
nand U5826 (N_5826,N_5634,N_5774);
nor U5827 (N_5827,N_5778,N_5755);
and U5828 (N_5828,N_5679,N_5735);
nand U5829 (N_5829,N_5694,N_5761);
and U5830 (N_5830,N_5673,N_5769);
nor U5831 (N_5831,N_5785,N_5692);
or U5832 (N_5832,N_5648,N_5770);
or U5833 (N_5833,N_5783,N_5667);
or U5834 (N_5834,N_5655,N_5771);
nand U5835 (N_5835,N_5798,N_5784);
and U5836 (N_5836,N_5661,N_5787);
nand U5837 (N_5837,N_5688,N_5615);
and U5838 (N_5838,N_5647,N_5700);
and U5839 (N_5839,N_5746,N_5780);
or U5840 (N_5840,N_5602,N_5656);
or U5841 (N_5841,N_5731,N_5690);
nand U5842 (N_5842,N_5762,N_5768);
nor U5843 (N_5843,N_5640,N_5628);
and U5844 (N_5844,N_5750,N_5683);
or U5845 (N_5845,N_5601,N_5663);
nor U5846 (N_5846,N_5729,N_5781);
or U5847 (N_5847,N_5659,N_5764);
and U5848 (N_5848,N_5638,N_5664);
nor U5849 (N_5849,N_5777,N_5772);
nand U5850 (N_5850,N_5790,N_5705);
and U5851 (N_5851,N_5723,N_5743);
nor U5852 (N_5852,N_5629,N_5765);
nor U5853 (N_5853,N_5733,N_5745);
nor U5854 (N_5854,N_5660,N_5635);
nand U5855 (N_5855,N_5653,N_5706);
nor U5856 (N_5856,N_5759,N_5794);
and U5857 (N_5857,N_5698,N_5707);
and U5858 (N_5858,N_5675,N_5708);
or U5859 (N_5859,N_5639,N_5604);
or U5860 (N_5860,N_5684,N_5753);
xor U5861 (N_5861,N_5788,N_5747);
or U5862 (N_5862,N_5622,N_5721);
xnor U5863 (N_5863,N_5773,N_5671);
nor U5864 (N_5864,N_5717,N_5658);
and U5865 (N_5865,N_5630,N_5676);
nand U5866 (N_5866,N_5722,N_5728);
xor U5867 (N_5867,N_5605,N_5691);
xor U5868 (N_5868,N_5716,N_5709);
and U5869 (N_5869,N_5715,N_5677);
nor U5870 (N_5870,N_5782,N_5760);
nand U5871 (N_5871,N_5652,N_5744);
nand U5872 (N_5872,N_5793,N_5670);
nor U5873 (N_5873,N_5775,N_5720);
nand U5874 (N_5874,N_5719,N_5616);
and U5875 (N_5875,N_5646,N_5792);
nand U5876 (N_5876,N_5618,N_5685);
and U5877 (N_5877,N_5696,N_5741);
xnor U5878 (N_5878,N_5791,N_5666);
and U5879 (N_5879,N_5643,N_5668);
xor U5880 (N_5880,N_5606,N_5712);
and U5881 (N_5881,N_5756,N_5710);
xor U5882 (N_5882,N_5620,N_5742);
nand U5883 (N_5883,N_5725,N_5678);
nor U5884 (N_5884,N_5752,N_5672);
nand U5885 (N_5885,N_5726,N_5695);
nor U5886 (N_5886,N_5600,N_5732);
or U5887 (N_5887,N_5734,N_5626);
or U5888 (N_5888,N_5730,N_5789);
nor U5889 (N_5889,N_5614,N_5641);
and U5890 (N_5890,N_5680,N_5763);
xnor U5891 (N_5891,N_5633,N_5621);
and U5892 (N_5892,N_5758,N_5713);
or U5893 (N_5893,N_5612,N_5751);
nor U5894 (N_5894,N_5697,N_5749);
and U5895 (N_5895,N_5608,N_5642);
xor U5896 (N_5896,N_5669,N_5650);
xnor U5897 (N_5897,N_5779,N_5619);
and U5898 (N_5898,N_5737,N_5662);
xnor U5899 (N_5899,N_5754,N_5687);
and U5900 (N_5900,N_5762,N_5744);
xor U5901 (N_5901,N_5645,N_5616);
or U5902 (N_5902,N_5714,N_5666);
or U5903 (N_5903,N_5734,N_5612);
and U5904 (N_5904,N_5701,N_5646);
xnor U5905 (N_5905,N_5706,N_5714);
and U5906 (N_5906,N_5779,N_5640);
xnor U5907 (N_5907,N_5727,N_5675);
nor U5908 (N_5908,N_5760,N_5736);
or U5909 (N_5909,N_5677,N_5746);
or U5910 (N_5910,N_5612,N_5630);
xnor U5911 (N_5911,N_5635,N_5663);
nand U5912 (N_5912,N_5679,N_5604);
nor U5913 (N_5913,N_5719,N_5702);
or U5914 (N_5914,N_5701,N_5703);
nand U5915 (N_5915,N_5713,N_5679);
xnor U5916 (N_5916,N_5746,N_5796);
nor U5917 (N_5917,N_5647,N_5606);
or U5918 (N_5918,N_5718,N_5652);
nor U5919 (N_5919,N_5750,N_5698);
nor U5920 (N_5920,N_5768,N_5664);
xnor U5921 (N_5921,N_5707,N_5638);
or U5922 (N_5922,N_5658,N_5780);
or U5923 (N_5923,N_5639,N_5614);
and U5924 (N_5924,N_5618,N_5632);
nand U5925 (N_5925,N_5661,N_5673);
xor U5926 (N_5926,N_5701,N_5630);
or U5927 (N_5927,N_5794,N_5748);
or U5928 (N_5928,N_5782,N_5748);
and U5929 (N_5929,N_5681,N_5739);
xor U5930 (N_5930,N_5756,N_5730);
nand U5931 (N_5931,N_5687,N_5705);
nor U5932 (N_5932,N_5719,N_5687);
and U5933 (N_5933,N_5632,N_5653);
nand U5934 (N_5934,N_5659,N_5797);
nor U5935 (N_5935,N_5640,N_5726);
nand U5936 (N_5936,N_5600,N_5746);
and U5937 (N_5937,N_5675,N_5615);
and U5938 (N_5938,N_5752,N_5666);
and U5939 (N_5939,N_5613,N_5723);
and U5940 (N_5940,N_5771,N_5645);
and U5941 (N_5941,N_5751,N_5642);
nand U5942 (N_5942,N_5706,N_5749);
and U5943 (N_5943,N_5602,N_5660);
nand U5944 (N_5944,N_5762,N_5702);
nand U5945 (N_5945,N_5634,N_5666);
nor U5946 (N_5946,N_5687,N_5600);
and U5947 (N_5947,N_5788,N_5655);
nand U5948 (N_5948,N_5607,N_5605);
nand U5949 (N_5949,N_5727,N_5653);
xnor U5950 (N_5950,N_5680,N_5749);
nand U5951 (N_5951,N_5648,N_5662);
and U5952 (N_5952,N_5756,N_5620);
nand U5953 (N_5953,N_5681,N_5772);
nor U5954 (N_5954,N_5684,N_5795);
nor U5955 (N_5955,N_5768,N_5632);
nand U5956 (N_5956,N_5660,N_5624);
xnor U5957 (N_5957,N_5612,N_5617);
xnor U5958 (N_5958,N_5671,N_5640);
or U5959 (N_5959,N_5675,N_5652);
nand U5960 (N_5960,N_5717,N_5631);
xor U5961 (N_5961,N_5735,N_5694);
nand U5962 (N_5962,N_5751,N_5602);
or U5963 (N_5963,N_5763,N_5667);
and U5964 (N_5964,N_5609,N_5639);
nand U5965 (N_5965,N_5721,N_5701);
xor U5966 (N_5966,N_5649,N_5619);
nand U5967 (N_5967,N_5624,N_5780);
nor U5968 (N_5968,N_5690,N_5728);
nor U5969 (N_5969,N_5731,N_5783);
and U5970 (N_5970,N_5699,N_5695);
nand U5971 (N_5971,N_5755,N_5754);
or U5972 (N_5972,N_5749,N_5730);
xor U5973 (N_5973,N_5647,N_5743);
or U5974 (N_5974,N_5677,N_5724);
nand U5975 (N_5975,N_5600,N_5724);
and U5976 (N_5976,N_5737,N_5733);
and U5977 (N_5977,N_5604,N_5709);
and U5978 (N_5978,N_5750,N_5688);
nand U5979 (N_5979,N_5746,N_5674);
and U5980 (N_5980,N_5626,N_5704);
nand U5981 (N_5981,N_5764,N_5781);
nor U5982 (N_5982,N_5655,N_5710);
nand U5983 (N_5983,N_5636,N_5789);
nand U5984 (N_5984,N_5614,N_5779);
and U5985 (N_5985,N_5662,N_5774);
or U5986 (N_5986,N_5654,N_5699);
nand U5987 (N_5987,N_5714,N_5721);
xor U5988 (N_5988,N_5799,N_5665);
nor U5989 (N_5989,N_5601,N_5643);
or U5990 (N_5990,N_5653,N_5607);
or U5991 (N_5991,N_5630,N_5686);
nor U5992 (N_5992,N_5739,N_5765);
xnor U5993 (N_5993,N_5780,N_5642);
and U5994 (N_5994,N_5679,N_5768);
nor U5995 (N_5995,N_5797,N_5746);
xnor U5996 (N_5996,N_5735,N_5709);
or U5997 (N_5997,N_5661,N_5641);
xor U5998 (N_5998,N_5636,N_5717);
xor U5999 (N_5999,N_5652,N_5607);
nor U6000 (N_6000,N_5882,N_5893);
or U6001 (N_6001,N_5889,N_5996);
or U6002 (N_6002,N_5952,N_5898);
xnor U6003 (N_6003,N_5878,N_5899);
nand U6004 (N_6004,N_5844,N_5880);
nor U6005 (N_6005,N_5817,N_5873);
and U6006 (N_6006,N_5860,N_5959);
xnor U6007 (N_6007,N_5886,N_5857);
xor U6008 (N_6008,N_5928,N_5947);
nand U6009 (N_6009,N_5840,N_5842);
and U6010 (N_6010,N_5975,N_5865);
or U6011 (N_6011,N_5832,N_5940);
nand U6012 (N_6012,N_5993,N_5820);
or U6013 (N_6013,N_5989,N_5931);
and U6014 (N_6014,N_5963,N_5872);
nand U6015 (N_6015,N_5866,N_5845);
nor U6016 (N_6016,N_5977,N_5911);
nor U6017 (N_6017,N_5968,N_5864);
nand U6018 (N_6018,N_5969,N_5901);
nor U6019 (N_6019,N_5988,N_5896);
and U6020 (N_6020,N_5935,N_5834);
or U6021 (N_6021,N_5822,N_5847);
nor U6022 (N_6022,N_5828,N_5978);
nor U6023 (N_6023,N_5868,N_5909);
nor U6024 (N_6024,N_5831,N_5819);
xnor U6025 (N_6025,N_5894,N_5926);
nand U6026 (N_6026,N_5803,N_5971);
nand U6027 (N_6027,N_5836,N_5964);
nor U6028 (N_6028,N_5994,N_5821);
and U6029 (N_6029,N_5841,N_5802);
and U6030 (N_6030,N_5995,N_5907);
xnor U6031 (N_6031,N_5801,N_5922);
or U6032 (N_6032,N_5936,N_5867);
or U6033 (N_6033,N_5932,N_5812);
nand U6034 (N_6034,N_5891,N_5892);
and U6035 (N_6035,N_5957,N_5917);
nor U6036 (N_6036,N_5815,N_5955);
nor U6037 (N_6037,N_5863,N_5854);
xor U6038 (N_6038,N_5944,N_5980);
nor U6039 (N_6039,N_5972,N_5982);
nor U6040 (N_6040,N_5902,N_5870);
xor U6041 (N_6041,N_5998,N_5883);
and U6042 (N_6042,N_5851,N_5999);
nand U6043 (N_6043,N_5943,N_5816);
nand U6044 (N_6044,N_5976,N_5987);
and U6045 (N_6045,N_5924,N_5912);
nand U6046 (N_6046,N_5833,N_5927);
nor U6047 (N_6047,N_5981,N_5914);
or U6048 (N_6048,N_5890,N_5948);
and U6049 (N_6049,N_5861,N_5965);
nor U6050 (N_6050,N_5973,N_5904);
nor U6051 (N_6051,N_5910,N_5921);
or U6052 (N_6052,N_5869,N_5837);
xnor U6053 (N_6053,N_5849,N_5915);
and U6054 (N_6054,N_5923,N_5941);
and U6055 (N_6055,N_5920,N_5954);
xnor U6056 (N_6056,N_5852,N_5877);
and U6057 (N_6057,N_5983,N_5949);
nor U6058 (N_6058,N_5974,N_5908);
and U6059 (N_6059,N_5830,N_5925);
nor U6060 (N_6060,N_5990,N_5827);
or U6061 (N_6061,N_5826,N_5905);
xor U6062 (N_6062,N_5811,N_5951);
and U6063 (N_6063,N_5960,N_5934);
and U6064 (N_6064,N_5810,N_5906);
xnor U6065 (N_6065,N_5884,N_5875);
and U6066 (N_6066,N_5945,N_5824);
xor U6067 (N_6067,N_5850,N_5853);
xor U6068 (N_6068,N_5813,N_5895);
or U6069 (N_6069,N_5806,N_5839);
nand U6070 (N_6070,N_5823,N_5956);
nor U6071 (N_6071,N_5871,N_5997);
or U6072 (N_6072,N_5809,N_5862);
xor U6073 (N_6073,N_5942,N_5825);
and U6074 (N_6074,N_5808,N_5966);
nand U6075 (N_6075,N_5967,N_5919);
and U6076 (N_6076,N_5953,N_5938);
nand U6077 (N_6077,N_5958,N_5804);
and U6078 (N_6078,N_5846,N_5986);
or U6079 (N_6079,N_5930,N_5876);
nor U6080 (N_6080,N_5929,N_5885);
nand U6081 (N_6081,N_5881,N_5835);
or U6082 (N_6082,N_5937,N_5887);
or U6083 (N_6083,N_5879,N_5918);
xor U6084 (N_6084,N_5979,N_5985);
and U6085 (N_6085,N_5962,N_5903);
and U6086 (N_6086,N_5939,N_5991);
and U6087 (N_6087,N_5848,N_5900);
nand U6088 (N_6088,N_5814,N_5800);
xnor U6089 (N_6089,N_5961,N_5888);
and U6090 (N_6090,N_5829,N_5897);
or U6091 (N_6091,N_5913,N_5843);
xor U6092 (N_6092,N_5807,N_5859);
and U6093 (N_6093,N_5805,N_5916);
nor U6094 (N_6094,N_5818,N_5874);
or U6095 (N_6095,N_5933,N_5858);
and U6096 (N_6096,N_5984,N_5970);
xor U6097 (N_6097,N_5946,N_5856);
nor U6098 (N_6098,N_5950,N_5992);
xnor U6099 (N_6099,N_5838,N_5855);
or U6100 (N_6100,N_5895,N_5846);
or U6101 (N_6101,N_5814,N_5914);
xnor U6102 (N_6102,N_5880,N_5888);
xnor U6103 (N_6103,N_5956,N_5827);
or U6104 (N_6104,N_5911,N_5945);
and U6105 (N_6105,N_5858,N_5943);
nor U6106 (N_6106,N_5833,N_5847);
and U6107 (N_6107,N_5934,N_5976);
xnor U6108 (N_6108,N_5871,N_5989);
or U6109 (N_6109,N_5847,N_5925);
nor U6110 (N_6110,N_5948,N_5876);
nand U6111 (N_6111,N_5981,N_5835);
and U6112 (N_6112,N_5927,N_5822);
nor U6113 (N_6113,N_5931,N_5854);
nor U6114 (N_6114,N_5849,N_5978);
xor U6115 (N_6115,N_5940,N_5908);
or U6116 (N_6116,N_5935,N_5928);
nand U6117 (N_6117,N_5945,N_5951);
and U6118 (N_6118,N_5868,N_5964);
nor U6119 (N_6119,N_5815,N_5962);
nor U6120 (N_6120,N_5888,N_5954);
nand U6121 (N_6121,N_5931,N_5884);
or U6122 (N_6122,N_5960,N_5867);
or U6123 (N_6123,N_5996,N_5918);
nand U6124 (N_6124,N_5861,N_5872);
nor U6125 (N_6125,N_5920,N_5951);
nand U6126 (N_6126,N_5802,N_5975);
nor U6127 (N_6127,N_5919,N_5996);
nand U6128 (N_6128,N_5886,N_5921);
or U6129 (N_6129,N_5828,N_5858);
or U6130 (N_6130,N_5820,N_5880);
xor U6131 (N_6131,N_5991,N_5903);
or U6132 (N_6132,N_5876,N_5891);
xnor U6133 (N_6133,N_5873,N_5942);
xnor U6134 (N_6134,N_5943,N_5879);
or U6135 (N_6135,N_5843,N_5882);
xor U6136 (N_6136,N_5840,N_5907);
and U6137 (N_6137,N_5864,N_5979);
or U6138 (N_6138,N_5821,N_5941);
or U6139 (N_6139,N_5866,N_5823);
xnor U6140 (N_6140,N_5929,N_5928);
or U6141 (N_6141,N_5835,N_5848);
xnor U6142 (N_6142,N_5844,N_5881);
nor U6143 (N_6143,N_5838,N_5944);
nand U6144 (N_6144,N_5891,N_5939);
nand U6145 (N_6145,N_5847,N_5877);
or U6146 (N_6146,N_5950,N_5834);
nand U6147 (N_6147,N_5825,N_5895);
and U6148 (N_6148,N_5836,N_5985);
nor U6149 (N_6149,N_5931,N_5852);
xor U6150 (N_6150,N_5800,N_5991);
or U6151 (N_6151,N_5892,N_5915);
xor U6152 (N_6152,N_5973,N_5821);
nand U6153 (N_6153,N_5900,N_5827);
xnor U6154 (N_6154,N_5890,N_5836);
and U6155 (N_6155,N_5976,N_5824);
nand U6156 (N_6156,N_5930,N_5933);
or U6157 (N_6157,N_5851,N_5823);
and U6158 (N_6158,N_5926,N_5944);
or U6159 (N_6159,N_5864,N_5803);
and U6160 (N_6160,N_5994,N_5967);
xnor U6161 (N_6161,N_5892,N_5908);
and U6162 (N_6162,N_5969,N_5866);
xnor U6163 (N_6163,N_5968,N_5887);
nand U6164 (N_6164,N_5826,N_5875);
and U6165 (N_6165,N_5955,N_5868);
xnor U6166 (N_6166,N_5965,N_5866);
xor U6167 (N_6167,N_5951,N_5977);
nand U6168 (N_6168,N_5876,N_5908);
and U6169 (N_6169,N_5997,N_5994);
nand U6170 (N_6170,N_5928,N_5836);
xnor U6171 (N_6171,N_5995,N_5874);
or U6172 (N_6172,N_5829,N_5985);
or U6173 (N_6173,N_5884,N_5990);
xor U6174 (N_6174,N_5904,N_5843);
or U6175 (N_6175,N_5817,N_5846);
and U6176 (N_6176,N_5930,N_5808);
nor U6177 (N_6177,N_5910,N_5828);
nor U6178 (N_6178,N_5943,N_5912);
nor U6179 (N_6179,N_5824,N_5998);
nand U6180 (N_6180,N_5862,N_5887);
nand U6181 (N_6181,N_5966,N_5811);
nand U6182 (N_6182,N_5814,N_5995);
and U6183 (N_6183,N_5825,N_5923);
nor U6184 (N_6184,N_5916,N_5827);
and U6185 (N_6185,N_5919,N_5891);
nand U6186 (N_6186,N_5937,N_5892);
nand U6187 (N_6187,N_5880,N_5861);
xnor U6188 (N_6188,N_5807,N_5919);
or U6189 (N_6189,N_5808,N_5944);
nand U6190 (N_6190,N_5946,N_5986);
nor U6191 (N_6191,N_5887,N_5809);
xor U6192 (N_6192,N_5905,N_5893);
or U6193 (N_6193,N_5802,N_5998);
xor U6194 (N_6194,N_5865,N_5921);
and U6195 (N_6195,N_5814,N_5969);
nand U6196 (N_6196,N_5821,N_5859);
nand U6197 (N_6197,N_5913,N_5873);
and U6198 (N_6198,N_5930,N_5804);
or U6199 (N_6199,N_5883,N_5864);
and U6200 (N_6200,N_6107,N_6061);
xnor U6201 (N_6201,N_6159,N_6000);
and U6202 (N_6202,N_6125,N_6162);
or U6203 (N_6203,N_6084,N_6197);
nand U6204 (N_6204,N_6196,N_6103);
nor U6205 (N_6205,N_6041,N_6127);
or U6206 (N_6206,N_6053,N_6095);
or U6207 (N_6207,N_6078,N_6019);
xor U6208 (N_6208,N_6088,N_6072);
nor U6209 (N_6209,N_6155,N_6080);
and U6210 (N_6210,N_6097,N_6066);
nand U6211 (N_6211,N_6176,N_6089);
nand U6212 (N_6212,N_6025,N_6005);
xnor U6213 (N_6213,N_6062,N_6108);
xnor U6214 (N_6214,N_6178,N_6016);
nor U6215 (N_6215,N_6166,N_6052);
and U6216 (N_6216,N_6049,N_6115);
nor U6217 (N_6217,N_6094,N_6035);
and U6218 (N_6218,N_6112,N_6135);
xor U6219 (N_6219,N_6104,N_6050);
nor U6220 (N_6220,N_6132,N_6079);
nor U6221 (N_6221,N_6101,N_6153);
or U6222 (N_6222,N_6075,N_6065);
and U6223 (N_6223,N_6007,N_6188);
and U6224 (N_6224,N_6038,N_6147);
nor U6225 (N_6225,N_6128,N_6064);
xnor U6226 (N_6226,N_6169,N_6146);
xnor U6227 (N_6227,N_6008,N_6027);
nand U6228 (N_6228,N_6122,N_6001);
nor U6229 (N_6229,N_6023,N_6119);
xnor U6230 (N_6230,N_6124,N_6189);
nor U6231 (N_6231,N_6192,N_6165);
or U6232 (N_6232,N_6054,N_6154);
or U6233 (N_6233,N_6024,N_6018);
xnor U6234 (N_6234,N_6140,N_6026);
nand U6235 (N_6235,N_6193,N_6130);
or U6236 (N_6236,N_6134,N_6173);
or U6237 (N_6237,N_6068,N_6172);
nor U6238 (N_6238,N_6092,N_6056);
xnor U6239 (N_6239,N_6170,N_6199);
and U6240 (N_6240,N_6070,N_6006);
nor U6241 (N_6241,N_6136,N_6100);
xnor U6242 (N_6242,N_6090,N_6151);
or U6243 (N_6243,N_6149,N_6185);
xor U6244 (N_6244,N_6057,N_6150);
and U6245 (N_6245,N_6022,N_6037);
and U6246 (N_6246,N_6017,N_6116);
xnor U6247 (N_6247,N_6020,N_6120);
nor U6248 (N_6248,N_6141,N_6129);
or U6249 (N_6249,N_6142,N_6010);
or U6250 (N_6250,N_6114,N_6043);
nand U6251 (N_6251,N_6152,N_6156);
xnor U6252 (N_6252,N_6144,N_6060);
nand U6253 (N_6253,N_6164,N_6081);
nand U6254 (N_6254,N_6163,N_6003);
nor U6255 (N_6255,N_6031,N_6184);
nand U6256 (N_6256,N_6091,N_6028);
nand U6257 (N_6257,N_6113,N_6085);
xnor U6258 (N_6258,N_6167,N_6182);
nor U6259 (N_6259,N_6076,N_6045);
or U6260 (N_6260,N_6137,N_6123);
xor U6261 (N_6261,N_6157,N_6133);
nand U6262 (N_6262,N_6039,N_6121);
nor U6263 (N_6263,N_6083,N_6187);
xor U6264 (N_6264,N_6033,N_6058);
nand U6265 (N_6265,N_6004,N_6109);
xnor U6266 (N_6266,N_6086,N_6082);
and U6267 (N_6267,N_6161,N_6047);
nor U6268 (N_6268,N_6105,N_6021);
xor U6269 (N_6269,N_6190,N_6071);
nand U6270 (N_6270,N_6012,N_6106);
xor U6271 (N_6271,N_6069,N_6015);
nand U6272 (N_6272,N_6096,N_6171);
nor U6273 (N_6273,N_6143,N_6148);
xor U6274 (N_6274,N_6181,N_6186);
xnor U6275 (N_6275,N_6139,N_6046);
nor U6276 (N_6276,N_6048,N_6118);
or U6277 (N_6277,N_6168,N_6032);
nand U6278 (N_6278,N_6051,N_6111);
and U6279 (N_6279,N_6117,N_6175);
xnor U6280 (N_6280,N_6110,N_6158);
nor U6281 (N_6281,N_6067,N_6055);
and U6282 (N_6282,N_6063,N_6177);
nand U6283 (N_6283,N_6042,N_6138);
xnor U6284 (N_6284,N_6093,N_6180);
nor U6285 (N_6285,N_6073,N_6098);
nand U6286 (N_6286,N_6099,N_6040);
and U6287 (N_6287,N_6145,N_6102);
or U6288 (N_6288,N_6077,N_6191);
xor U6289 (N_6289,N_6002,N_6074);
xor U6290 (N_6290,N_6087,N_6160);
or U6291 (N_6291,N_6183,N_6011);
or U6292 (N_6292,N_6126,N_6034);
xor U6293 (N_6293,N_6198,N_6044);
xor U6294 (N_6294,N_6030,N_6194);
nand U6295 (N_6295,N_6059,N_6131);
nor U6296 (N_6296,N_6195,N_6174);
nand U6297 (N_6297,N_6029,N_6014);
or U6298 (N_6298,N_6036,N_6013);
nand U6299 (N_6299,N_6179,N_6009);
nor U6300 (N_6300,N_6188,N_6193);
and U6301 (N_6301,N_6060,N_6102);
xor U6302 (N_6302,N_6085,N_6179);
nor U6303 (N_6303,N_6078,N_6108);
nand U6304 (N_6304,N_6029,N_6153);
xnor U6305 (N_6305,N_6040,N_6198);
or U6306 (N_6306,N_6039,N_6093);
or U6307 (N_6307,N_6183,N_6199);
nand U6308 (N_6308,N_6050,N_6030);
and U6309 (N_6309,N_6197,N_6004);
and U6310 (N_6310,N_6058,N_6045);
xnor U6311 (N_6311,N_6116,N_6040);
or U6312 (N_6312,N_6050,N_6160);
or U6313 (N_6313,N_6061,N_6133);
and U6314 (N_6314,N_6153,N_6074);
nor U6315 (N_6315,N_6101,N_6080);
nand U6316 (N_6316,N_6044,N_6103);
and U6317 (N_6317,N_6174,N_6163);
and U6318 (N_6318,N_6028,N_6004);
and U6319 (N_6319,N_6081,N_6137);
nand U6320 (N_6320,N_6033,N_6150);
or U6321 (N_6321,N_6137,N_6028);
xor U6322 (N_6322,N_6043,N_6111);
xnor U6323 (N_6323,N_6173,N_6050);
or U6324 (N_6324,N_6136,N_6193);
and U6325 (N_6325,N_6020,N_6046);
nand U6326 (N_6326,N_6095,N_6008);
xor U6327 (N_6327,N_6026,N_6195);
nand U6328 (N_6328,N_6098,N_6085);
or U6329 (N_6329,N_6068,N_6040);
nor U6330 (N_6330,N_6024,N_6016);
nor U6331 (N_6331,N_6153,N_6061);
nand U6332 (N_6332,N_6093,N_6011);
or U6333 (N_6333,N_6174,N_6008);
xor U6334 (N_6334,N_6051,N_6113);
nand U6335 (N_6335,N_6065,N_6086);
xnor U6336 (N_6336,N_6199,N_6014);
and U6337 (N_6337,N_6079,N_6187);
or U6338 (N_6338,N_6091,N_6153);
xor U6339 (N_6339,N_6099,N_6049);
and U6340 (N_6340,N_6029,N_6056);
nor U6341 (N_6341,N_6043,N_6044);
and U6342 (N_6342,N_6104,N_6112);
or U6343 (N_6343,N_6115,N_6113);
nand U6344 (N_6344,N_6095,N_6017);
xor U6345 (N_6345,N_6035,N_6104);
and U6346 (N_6346,N_6135,N_6194);
or U6347 (N_6347,N_6034,N_6147);
nand U6348 (N_6348,N_6045,N_6031);
nand U6349 (N_6349,N_6107,N_6045);
and U6350 (N_6350,N_6069,N_6019);
nor U6351 (N_6351,N_6129,N_6198);
or U6352 (N_6352,N_6119,N_6172);
xnor U6353 (N_6353,N_6049,N_6119);
or U6354 (N_6354,N_6051,N_6075);
nor U6355 (N_6355,N_6078,N_6011);
and U6356 (N_6356,N_6083,N_6019);
nand U6357 (N_6357,N_6148,N_6183);
nand U6358 (N_6358,N_6035,N_6149);
xor U6359 (N_6359,N_6131,N_6176);
and U6360 (N_6360,N_6057,N_6084);
xnor U6361 (N_6361,N_6100,N_6006);
or U6362 (N_6362,N_6195,N_6070);
nor U6363 (N_6363,N_6058,N_6070);
and U6364 (N_6364,N_6093,N_6136);
nor U6365 (N_6365,N_6134,N_6129);
nand U6366 (N_6366,N_6115,N_6037);
and U6367 (N_6367,N_6027,N_6119);
or U6368 (N_6368,N_6117,N_6002);
nand U6369 (N_6369,N_6127,N_6023);
nand U6370 (N_6370,N_6032,N_6138);
and U6371 (N_6371,N_6151,N_6190);
or U6372 (N_6372,N_6071,N_6134);
xor U6373 (N_6373,N_6081,N_6015);
nor U6374 (N_6374,N_6096,N_6052);
and U6375 (N_6375,N_6194,N_6175);
nor U6376 (N_6376,N_6172,N_6178);
and U6377 (N_6377,N_6003,N_6116);
nand U6378 (N_6378,N_6166,N_6102);
nor U6379 (N_6379,N_6063,N_6193);
and U6380 (N_6380,N_6043,N_6171);
or U6381 (N_6381,N_6004,N_6177);
nor U6382 (N_6382,N_6035,N_6076);
nor U6383 (N_6383,N_6136,N_6151);
xnor U6384 (N_6384,N_6024,N_6165);
nand U6385 (N_6385,N_6066,N_6077);
nor U6386 (N_6386,N_6075,N_6187);
nor U6387 (N_6387,N_6113,N_6136);
or U6388 (N_6388,N_6183,N_6076);
or U6389 (N_6389,N_6105,N_6189);
nor U6390 (N_6390,N_6065,N_6048);
xor U6391 (N_6391,N_6066,N_6120);
nor U6392 (N_6392,N_6083,N_6156);
and U6393 (N_6393,N_6095,N_6060);
nand U6394 (N_6394,N_6034,N_6187);
xor U6395 (N_6395,N_6149,N_6051);
and U6396 (N_6396,N_6101,N_6065);
or U6397 (N_6397,N_6190,N_6116);
nand U6398 (N_6398,N_6028,N_6055);
or U6399 (N_6399,N_6144,N_6079);
nand U6400 (N_6400,N_6302,N_6240);
xor U6401 (N_6401,N_6299,N_6369);
or U6402 (N_6402,N_6384,N_6362);
xor U6403 (N_6403,N_6378,N_6395);
nor U6404 (N_6404,N_6211,N_6271);
nor U6405 (N_6405,N_6263,N_6320);
or U6406 (N_6406,N_6340,N_6322);
nor U6407 (N_6407,N_6326,N_6393);
xor U6408 (N_6408,N_6351,N_6266);
xnor U6409 (N_6409,N_6390,N_6377);
xor U6410 (N_6410,N_6366,N_6279);
and U6411 (N_6411,N_6282,N_6231);
nor U6412 (N_6412,N_6288,N_6388);
nand U6413 (N_6413,N_6298,N_6215);
or U6414 (N_6414,N_6248,N_6249);
nor U6415 (N_6415,N_6373,N_6316);
nand U6416 (N_6416,N_6386,N_6353);
and U6417 (N_6417,N_6260,N_6338);
or U6418 (N_6418,N_6250,N_6284);
or U6419 (N_6419,N_6281,N_6274);
or U6420 (N_6420,N_6308,N_6254);
nor U6421 (N_6421,N_6247,N_6348);
or U6422 (N_6422,N_6257,N_6355);
xor U6423 (N_6423,N_6214,N_6262);
xnor U6424 (N_6424,N_6224,N_6333);
or U6425 (N_6425,N_6295,N_6331);
nor U6426 (N_6426,N_6312,N_6341);
and U6427 (N_6427,N_6327,N_6309);
nor U6428 (N_6428,N_6286,N_6365);
nand U6429 (N_6429,N_6229,N_6216);
xor U6430 (N_6430,N_6367,N_6237);
and U6431 (N_6431,N_6354,N_6346);
or U6432 (N_6432,N_6336,N_6324);
nor U6433 (N_6433,N_6251,N_6310);
nor U6434 (N_6434,N_6283,N_6379);
nor U6435 (N_6435,N_6387,N_6398);
xor U6436 (N_6436,N_6317,N_6360);
or U6437 (N_6437,N_6217,N_6313);
nand U6438 (N_6438,N_6218,N_6246);
nor U6439 (N_6439,N_6370,N_6287);
nand U6440 (N_6440,N_6226,N_6212);
and U6441 (N_6441,N_6293,N_6272);
and U6442 (N_6442,N_6396,N_6306);
xor U6443 (N_6443,N_6368,N_6305);
xnor U6444 (N_6444,N_6359,N_6397);
and U6445 (N_6445,N_6399,N_6383);
and U6446 (N_6446,N_6256,N_6374);
or U6447 (N_6447,N_6297,N_6380);
or U6448 (N_6448,N_6291,N_6385);
or U6449 (N_6449,N_6208,N_6227);
nor U6450 (N_6450,N_6325,N_6392);
nor U6451 (N_6451,N_6372,N_6290);
nor U6452 (N_6452,N_6278,N_6352);
and U6453 (N_6453,N_6311,N_6394);
and U6454 (N_6454,N_6233,N_6364);
or U6455 (N_6455,N_6277,N_6264);
and U6456 (N_6456,N_6234,N_6381);
or U6457 (N_6457,N_6332,N_6307);
xor U6458 (N_6458,N_6343,N_6301);
xor U6459 (N_6459,N_6220,N_6253);
or U6460 (N_6460,N_6222,N_6201);
and U6461 (N_6461,N_6202,N_6389);
nand U6462 (N_6462,N_6314,N_6319);
and U6463 (N_6463,N_6328,N_6382);
and U6464 (N_6464,N_6252,N_6329);
or U6465 (N_6465,N_6344,N_6221);
nand U6466 (N_6466,N_6391,N_6267);
nand U6467 (N_6467,N_6375,N_6228);
nor U6468 (N_6468,N_6371,N_6330);
xor U6469 (N_6469,N_6357,N_6206);
or U6470 (N_6470,N_6323,N_6356);
nor U6471 (N_6471,N_6361,N_6350);
or U6472 (N_6472,N_6294,N_6261);
nor U6473 (N_6473,N_6347,N_6349);
xnor U6474 (N_6474,N_6243,N_6245);
nor U6475 (N_6475,N_6230,N_6270);
and U6476 (N_6476,N_6363,N_6321);
nor U6477 (N_6477,N_6225,N_6303);
xor U6478 (N_6478,N_6276,N_6376);
or U6479 (N_6479,N_6315,N_6219);
xnor U6480 (N_6480,N_6345,N_6213);
or U6481 (N_6481,N_6318,N_6242);
nor U6482 (N_6482,N_6280,N_6304);
or U6483 (N_6483,N_6241,N_6238);
xnor U6484 (N_6484,N_6210,N_6235);
xnor U6485 (N_6485,N_6232,N_6209);
xor U6486 (N_6486,N_6275,N_6204);
nand U6487 (N_6487,N_6258,N_6265);
nand U6488 (N_6488,N_6335,N_6200);
xor U6489 (N_6489,N_6236,N_6239);
nor U6490 (N_6490,N_6339,N_6269);
and U6491 (N_6491,N_6337,N_6300);
or U6492 (N_6492,N_6223,N_6296);
and U6493 (N_6493,N_6203,N_6205);
and U6494 (N_6494,N_6358,N_6285);
nor U6495 (N_6495,N_6292,N_6259);
or U6496 (N_6496,N_6268,N_6255);
and U6497 (N_6497,N_6334,N_6342);
xor U6498 (N_6498,N_6289,N_6207);
nor U6499 (N_6499,N_6273,N_6244);
nand U6500 (N_6500,N_6227,N_6379);
xor U6501 (N_6501,N_6233,N_6294);
or U6502 (N_6502,N_6351,N_6282);
nand U6503 (N_6503,N_6388,N_6212);
nor U6504 (N_6504,N_6361,N_6378);
nor U6505 (N_6505,N_6283,N_6265);
and U6506 (N_6506,N_6313,N_6238);
or U6507 (N_6507,N_6302,N_6249);
nor U6508 (N_6508,N_6329,N_6333);
nor U6509 (N_6509,N_6323,N_6294);
nand U6510 (N_6510,N_6217,N_6218);
or U6511 (N_6511,N_6230,N_6330);
nand U6512 (N_6512,N_6382,N_6258);
and U6513 (N_6513,N_6227,N_6315);
or U6514 (N_6514,N_6309,N_6325);
or U6515 (N_6515,N_6287,N_6340);
xor U6516 (N_6516,N_6391,N_6340);
nand U6517 (N_6517,N_6374,N_6262);
xnor U6518 (N_6518,N_6261,N_6311);
xor U6519 (N_6519,N_6311,N_6335);
and U6520 (N_6520,N_6234,N_6361);
or U6521 (N_6521,N_6235,N_6360);
and U6522 (N_6522,N_6318,N_6203);
nor U6523 (N_6523,N_6353,N_6241);
nand U6524 (N_6524,N_6370,N_6277);
or U6525 (N_6525,N_6341,N_6226);
or U6526 (N_6526,N_6319,N_6343);
or U6527 (N_6527,N_6232,N_6336);
and U6528 (N_6528,N_6313,N_6389);
and U6529 (N_6529,N_6320,N_6288);
and U6530 (N_6530,N_6374,N_6235);
nor U6531 (N_6531,N_6338,N_6227);
or U6532 (N_6532,N_6346,N_6264);
nand U6533 (N_6533,N_6319,N_6396);
nand U6534 (N_6534,N_6234,N_6311);
and U6535 (N_6535,N_6246,N_6330);
or U6536 (N_6536,N_6396,N_6323);
or U6537 (N_6537,N_6283,N_6304);
xor U6538 (N_6538,N_6235,N_6303);
or U6539 (N_6539,N_6391,N_6345);
and U6540 (N_6540,N_6380,N_6299);
xnor U6541 (N_6541,N_6297,N_6398);
nor U6542 (N_6542,N_6221,N_6312);
and U6543 (N_6543,N_6349,N_6336);
xnor U6544 (N_6544,N_6293,N_6309);
or U6545 (N_6545,N_6342,N_6263);
and U6546 (N_6546,N_6382,N_6314);
nor U6547 (N_6547,N_6376,N_6298);
nor U6548 (N_6548,N_6240,N_6259);
or U6549 (N_6549,N_6391,N_6295);
or U6550 (N_6550,N_6274,N_6389);
and U6551 (N_6551,N_6265,N_6292);
or U6552 (N_6552,N_6285,N_6397);
or U6553 (N_6553,N_6265,N_6384);
or U6554 (N_6554,N_6297,N_6296);
and U6555 (N_6555,N_6388,N_6335);
xnor U6556 (N_6556,N_6398,N_6301);
or U6557 (N_6557,N_6359,N_6347);
nand U6558 (N_6558,N_6281,N_6354);
xnor U6559 (N_6559,N_6395,N_6351);
or U6560 (N_6560,N_6211,N_6347);
xor U6561 (N_6561,N_6253,N_6204);
nand U6562 (N_6562,N_6266,N_6215);
nand U6563 (N_6563,N_6300,N_6352);
nor U6564 (N_6564,N_6294,N_6309);
or U6565 (N_6565,N_6359,N_6374);
xnor U6566 (N_6566,N_6268,N_6295);
nand U6567 (N_6567,N_6317,N_6316);
xor U6568 (N_6568,N_6246,N_6252);
nor U6569 (N_6569,N_6378,N_6348);
or U6570 (N_6570,N_6327,N_6374);
nand U6571 (N_6571,N_6268,N_6378);
and U6572 (N_6572,N_6226,N_6374);
and U6573 (N_6573,N_6250,N_6306);
nor U6574 (N_6574,N_6265,N_6204);
and U6575 (N_6575,N_6209,N_6245);
nor U6576 (N_6576,N_6334,N_6250);
nor U6577 (N_6577,N_6285,N_6327);
nand U6578 (N_6578,N_6374,N_6309);
xnor U6579 (N_6579,N_6327,N_6335);
or U6580 (N_6580,N_6334,N_6341);
or U6581 (N_6581,N_6224,N_6374);
xnor U6582 (N_6582,N_6222,N_6312);
nor U6583 (N_6583,N_6333,N_6264);
and U6584 (N_6584,N_6370,N_6271);
nand U6585 (N_6585,N_6349,N_6361);
nor U6586 (N_6586,N_6339,N_6233);
nand U6587 (N_6587,N_6350,N_6365);
and U6588 (N_6588,N_6353,N_6272);
or U6589 (N_6589,N_6352,N_6320);
and U6590 (N_6590,N_6336,N_6383);
or U6591 (N_6591,N_6355,N_6293);
and U6592 (N_6592,N_6338,N_6273);
nor U6593 (N_6593,N_6264,N_6295);
nand U6594 (N_6594,N_6389,N_6248);
xnor U6595 (N_6595,N_6321,N_6294);
nor U6596 (N_6596,N_6232,N_6219);
or U6597 (N_6597,N_6331,N_6325);
nand U6598 (N_6598,N_6358,N_6316);
and U6599 (N_6599,N_6380,N_6307);
or U6600 (N_6600,N_6510,N_6563);
nand U6601 (N_6601,N_6432,N_6555);
xor U6602 (N_6602,N_6568,N_6448);
nor U6603 (N_6603,N_6523,N_6478);
or U6604 (N_6604,N_6522,N_6530);
nand U6605 (N_6605,N_6470,N_6415);
nand U6606 (N_6606,N_6508,N_6519);
nand U6607 (N_6607,N_6583,N_6550);
and U6608 (N_6608,N_6484,N_6474);
nand U6609 (N_6609,N_6412,N_6562);
and U6610 (N_6610,N_6435,N_6401);
and U6611 (N_6611,N_6536,N_6431);
xnor U6612 (N_6612,N_6503,N_6535);
xnor U6613 (N_6613,N_6586,N_6572);
or U6614 (N_6614,N_6445,N_6512);
nand U6615 (N_6615,N_6529,N_6417);
nor U6616 (N_6616,N_6579,N_6488);
nor U6617 (N_6617,N_6442,N_6569);
xor U6618 (N_6618,N_6476,N_6539);
or U6619 (N_6619,N_6520,N_6564);
or U6620 (N_6620,N_6594,N_6558);
xnor U6621 (N_6621,N_6490,N_6407);
nand U6622 (N_6622,N_6596,N_6425);
nor U6623 (N_6623,N_6597,N_6500);
and U6624 (N_6624,N_6440,N_6495);
nor U6625 (N_6625,N_6492,N_6505);
and U6626 (N_6626,N_6411,N_6454);
and U6627 (N_6627,N_6494,N_6537);
and U6628 (N_6628,N_6464,N_6557);
or U6629 (N_6629,N_6541,N_6590);
and U6630 (N_6630,N_6414,N_6592);
xor U6631 (N_6631,N_6554,N_6466);
xnor U6632 (N_6632,N_6540,N_6424);
nor U6633 (N_6633,N_6433,N_6497);
nor U6634 (N_6634,N_6422,N_6444);
or U6635 (N_6635,N_6589,N_6434);
nand U6636 (N_6636,N_6524,N_6504);
or U6637 (N_6637,N_6566,N_6410);
and U6638 (N_6638,N_6588,N_6599);
nand U6639 (N_6639,N_6450,N_6573);
xnor U6640 (N_6640,N_6518,N_6409);
xor U6641 (N_6641,N_6570,N_6514);
nor U6642 (N_6642,N_6565,N_6577);
xor U6643 (N_6643,N_6534,N_6493);
nor U6644 (N_6644,N_6501,N_6453);
nand U6645 (N_6645,N_6451,N_6449);
or U6646 (N_6646,N_6413,N_6416);
xnor U6647 (N_6647,N_6427,N_6489);
or U6648 (N_6648,N_6538,N_6582);
or U6649 (N_6649,N_6404,N_6581);
nor U6650 (N_6650,N_6515,N_6471);
or U6651 (N_6651,N_6468,N_6461);
or U6652 (N_6652,N_6467,N_6498);
nand U6653 (N_6653,N_6487,N_6446);
or U6654 (N_6654,N_6456,N_6548);
or U6655 (N_6655,N_6525,N_6420);
nor U6656 (N_6656,N_6400,N_6481);
or U6657 (N_6657,N_6511,N_6598);
nand U6658 (N_6658,N_6463,N_6560);
and U6659 (N_6659,N_6595,N_6408);
and U6660 (N_6660,N_6496,N_6426);
or U6661 (N_6661,N_6419,N_6475);
nand U6662 (N_6662,N_6593,N_6437);
and U6663 (N_6663,N_6587,N_6521);
or U6664 (N_6664,N_6513,N_6459);
or U6665 (N_6665,N_6472,N_6559);
nand U6666 (N_6666,N_6546,N_6452);
or U6667 (N_6667,N_6567,N_6439);
nor U6668 (N_6668,N_6547,N_6552);
or U6669 (N_6669,N_6473,N_6516);
nor U6670 (N_6670,N_6491,N_6580);
or U6671 (N_6671,N_6502,N_6509);
nor U6672 (N_6672,N_6418,N_6527);
xnor U6673 (N_6673,N_6578,N_6405);
and U6674 (N_6674,N_6479,N_6460);
nand U6675 (N_6675,N_6455,N_6545);
xor U6676 (N_6676,N_6441,N_6421);
nor U6677 (N_6677,N_6480,N_6483);
nand U6678 (N_6678,N_6486,N_6543);
nand U6679 (N_6679,N_6465,N_6533);
or U6680 (N_6680,N_6403,N_6576);
xor U6681 (N_6681,N_6436,N_6402);
nand U6682 (N_6682,N_6585,N_6561);
and U6683 (N_6683,N_6458,N_6499);
nor U6684 (N_6684,N_6584,N_6429);
nor U6685 (N_6685,N_6430,N_6556);
or U6686 (N_6686,N_6469,N_6542);
nor U6687 (N_6687,N_6443,N_6591);
or U6688 (N_6688,N_6571,N_6438);
or U6689 (N_6689,N_6447,N_6406);
xor U6690 (N_6690,N_6532,N_6477);
xnor U6691 (N_6691,N_6506,N_6482);
nor U6692 (N_6692,N_6457,N_6544);
nor U6693 (N_6693,N_6549,N_6485);
and U6694 (N_6694,N_6462,N_6428);
xnor U6695 (N_6695,N_6528,N_6531);
nor U6696 (N_6696,N_6507,N_6551);
xor U6697 (N_6697,N_6526,N_6517);
nand U6698 (N_6698,N_6575,N_6574);
nand U6699 (N_6699,N_6423,N_6553);
or U6700 (N_6700,N_6552,N_6585);
or U6701 (N_6701,N_6516,N_6414);
xnor U6702 (N_6702,N_6592,N_6566);
nand U6703 (N_6703,N_6579,N_6576);
nand U6704 (N_6704,N_6436,N_6443);
and U6705 (N_6705,N_6487,N_6402);
nor U6706 (N_6706,N_6514,N_6455);
and U6707 (N_6707,N_6415,N_6469);
and U6708 (N_6708,N_6412,N_6427);
nand U6709 (N_6709,N_6536,N_6580);
or U6710 (N_6710,N_6583,N_6516);
nand U6711 (N_6711,N_6463,N_6490);
and U6712 (N_6712,N_6566,N_6428);
nor U6713 (N_6713,N_6583,N_6452);
nand U6714 (N_6714,N_6548,N_6477);
or U6715 (N_6715,N_6461,N_6490);
nor U6716 (N_6716,N_6561,N_6440);
nand U6717 (N_6717,N_6427,N_6501);
or U6718 (N_6718,N_6593,N_6568);
nand U6719 (N_6719,N_6543,N_6565);
nor U6720 (N_6720,N_6516,N_6513);
and U6721 (N_6721,N_6474,N_6406);
nand U6722 (N_6722,N_6403,N_6571);
nand U6723 (N_6723,N_6521,N_6428);
xor U6724 (N_6724,N_6406,N_6554);
and U6725 (N_6725,N_6446,N_6567);
nor U6726 (N_6726,N_6554,N_6562);
nor U6727 (N_6727,N_6521,N_6545);
or U6728 (N_6728,N_6430,N_6422);
nor U6729 (N_6729,N_6483,N_6470);
or U6730 (N_6730,N_6587,N_6575);
nand U6731 (N_6731,N_6462,N_6437);
xnor U6732 (N_6732,N_6414,N_6529);
nor U6733 (N_6733,N_6542,N_6539);
xor U6734 (N_6734,N_6424,N_6447);
nor U6735 (N_6735,N_6475,N_6513);
nor U6736 (N_6736,N_6412,N_6417);
nor U6737 (N_6737,N_6467,N_6563);
nand U6738 (N_6738,N_6509,N_6429);
and U6739 (N_6739,N_6553,N_6506);
nor U6740 (N_6740,N_6589,N_6459);
or U6741 (N_6741,N_6549,N_6480);
nand U6742 (N_6742,N_6441,N_6565);
nand U6743 (N_6743,N_6435,N_6424);
and U6744 (N_6744,N_6544,N_6576);
nor U6745 (N_6745,N_6579,N_6559);
nor U6746 (N_6746,N_6447,N_6506);
xor U6747 (N_6747,N_6479,N_6544);
and U6748 (N_6748,N_6599,N_6561);
nor U6749 (N_6749,N_6581,N_6442);
nor U6750 (N_6750,N_6425,N_6570);
or U6751 (N_6751,N_6555,N_6595);
nand U6752 (N_6752,N_6451,N_6417);
and U6753 (N_6753,N_6497,N_6412);
xnor U6754 (N_6754,N_6590,N_6538);
nand U6755 (N_6755,N_6588,N_6533);
or U6756 (N_6756,N_6548,N_6553);
xor U6757 (N_6757,N_6417,N_6423);
and U6758 (N_6758,N_6555,N_6404);
nand U6759 (N_6759,N_6495,N_6526);
nor U6760 (N_6760,N_6446,N_6414);
or U6761 (N_6761,N_6579,N_6511);
and U6762 (N_6762,N_6599,N_6495);
nor U6763 (N_6763,N_6406,N_6582);
nand U6764 (N_6764,N_6442,N_6449);
and U6765 (N_6765,N_6564,N_6422);
and U6766 (N_6766,N_6546,N_6436);
nor U6767 (N_6767,N_6529,N_6587);
or U6768 (N_6768,N_6571,N_6447);
nand U6769 (N_6769,N_6575,N_6507);
xor U6770 (N_6770,N_6587,N_6431);
or U6771 (N_6771,N_6555,N_6552);
or U6772 (N_6772,N_6447,N_6587);
xor U6773 (N_6773,N_6559,N_6538);
xnor U6774 (N_6774,N_6461,N_6564);
and U6775 (N_6775,N_6485,N_6471);
nand U6776 (N_6776,N_6444,N_6497);
xor U6777 (N_6777,N_6440,N_6489);
and U6778 (N_6778,N_6544,N_6488);
nor U6779 (N_6779,N_6561,N_6453);
xor U6780 (N_6780,N_6516,N_6486);
and U6781 (N_6781,N_6525,N_6441);
xor U6782 (N_6782,N_6436,N_6540);
nor U6783 (N_6783,N_6449,N_6528);
nand U6784 (N_6784,N_6527,N_6476);
nand U6785 (N_6785,N_6575,N_6543);
xor U6786 (N_6786,N_6560,N_6480);
nand U6787 (N_6787,N_6537,N_6457);
or U6788 (N_6788,N_6507,N_6577);
nor U6789 (N_6789,N_6553,N_6488);
xor U6790 (N_6790,N_6597,N_6452);
nor U6791 (N_6791,N_6519,N_6514);
and U6792 (N_6792,N_6516,N_6542);
xnor U6793 (N_6793,N_6580,N_6515);
xnor U6794 (N_6794,N_6450,N_6560);
or U6795 (N_6795,N_6544,N_6542);
or U6796 (N_6796,N_6474,N_6599);
or U6797 (N_6797,N_6512,N_6424);
and U6798 (N_6798,N_6533,N_6598);
or U6799 (N_6799,N_6412,N_6479);
xor U6800 (N_6800,N_6648,N_6761);
xnor U6801 (N_6801,N_6713,N_6773);
nand U6802 (N_6802,N_6751,N_6609);
xor U6803 (N_6803,N_6606,N_6607);
xor U6804 (N_6804,N_6744,N_6700);
or U6805 (N_6805,N_6786,N_6624);
nand U6806 (N_6806,N_6680,N_6762);
and U6807 (N_6807,N_6633,N_6640);
nand U6808 (N_6808,N_6637,N_6676);
nand U6809 (N_6809,N_6741,N_6667);
and U6810 (N_6810,N_6675,N_6707);
nor U6811 (N_6811,N_6757,N_6652);
or U6812 (N_6812,N_6706,N_6692);
xnor U6813 (N_6813,N_6691,N_6725);
xnor U6814 (N_6814,N_6695,N_6778);
nand U6815 (N_6815,N_6669,N_6622);
xor U6816 (N_6816,N_6765,N_6797);
nand U6817 (N_6817,N_6779,N_6715);
or U6818 (N_6818,N_6618,N_6641);
or U6819 (N_6819,N_6623,N_6681);
xor U6820 (N_6820,N_6730,N_6662);
nand U6821 (N_6821,N_6718,N_6722);
xor U6822 (N_6822,N_6697,N_6738);
nand U6823 (N_6823,N_6732,N_6764);
and U6824 (N_6824,N_6754,N_6705);
nor U6825 (N_6825,N_6702,N_6616);
and U6826 (N_6826,N_6763,N_6717);
nor U6827 (N_6827,N_6704,N_6690);
nand U6828 (N_6828,N_6739,N_6785);
nor U6829 (N_6829,N_6649,N_6740);
and U6830 (N_6830,N_6798,N_6708);
or U6831 (N_6831,N_6632,N_6639);
or U6832 (N_6832,N_6612,N_6716);
and U6833 (N_6833,N_6677,N_6694);
nor U6834 (N_6834,N_6682,N_6627);
or U6835 (N_6835,N_6656,N_6769);
nand U6836 (N_6836,N_6613,N_6636);
and U6837 (N_6837,N_6768,N_6683);
nand U6838 (N_6838,N_6767,N_6789);
nand U6839 (N_6839,N_6614,N_6696);
xor U6840 (N_6840,N_6657,N_6688);
and U6841 (N_6841,N_6653,N_6780);
or U6842 (N_6842,N_6787,N_6745);
xnor U6843 (N_6843,N_6790,N_6794);
and U6844 (N_6844,N_6734,N_6693);
xor U6845 (N_6845,N_6660,N_6748);
or U6846 (N_6846,N_6753,N_6645);
nor U6847 (N_6847,N_6710,N_6635);
xnor U6848 (N_6848,N_6735,N_6668);
or U6849 (N_6849,N_6631,N_6755);
or U6850 (N_6850,N_6665,N_6759);
xor U6851 (N_6851,N_6726,N_6719);
and U6852 (N_6852,N_6630,N_6781);
and U6853 (N_6853,N_6663,N_6777);
nand U6854 (N_6854,N_6658,N_6721);
nand U6855 (N_6855,N_6600,N_6699);
nor U6856 (N_6856,N_6720,N_6603);
nand U6857 (N_6857,N_6617,N_6711);
nor U6858 (N_6858,N_6771,N_6724);
or U6859 (N_6859,N_6604,N_6770);
xor U6860 (N_6860,N_6701,N_6642);
nand U6861 (N_6861,N_6601,N_6664);
and U6862 (N_6862,N_6698,N_6742);
and U6863 (N_6863,N_6685,N_6774);
nand U6864 (N_6864,N_6793,N_6673);
nand U6865 (N_6865,N_6611,N_6625);
nand U6866 (N_6866,N_6647,N_6799);
xnor U6867 (N_6867,N_6709,N_6703);
nand U6868 (N_6868,N_6621,N_6791);
or U6869 (N_6869,N_6752,N_6687);
or U6870 (N_6870,N_6784,N_6608);
xor U6871 (N_6871,N_6758,N_6650);
xnor U6872 (N_6872,N_6733,N_6629);
and U6873 (N_6873,N_6646,N_6638);
nor U6874 (N_6874,N_6729,N_6736);
and U6875 (N_6875,N_6788,N_6746);
or U6876 (N_6876,N_6689,N_6750);
xnor U6877 (N_6877,N_6731,N_6659);
or U6878 (N_6878,N_6626,N_6766);
and U6879 (N_6879,N_6655,N_6644);
nand U6880 (N_6880,N_6783,N_6686);
and U6881 (N_6881,N_6670,N_6723);
nand U6882 (N_6882,N_6678,N_6605);
or U6883 (N_6883,N_6634,N_6672);
nand U6884 (N_6884,N_6772,N_6792);
and U6885 (N_6885,N_6619,N_6756);
xnor U6886 (N_6886,N_6679,N_6747);
or U6887 (N_6887,N_6796,N_6674);
xor U6888 (N_6888,N_6712,N_6749);
or U6889 (N_6889,N_6743,N_6727);
xnor U6890 (N_6890,N_6671,N_6661);
nor U6891 (N_6891,N_6654,N_6620);
nand U6892 (N_6892,N_6760,N_6737);
nor U6893 (N_6893,N_6728,N_6643);
nor U6894 (N_6894,N_6651,N_6615);
or U6895 (N_6895,N_6776,N_6628);
nor U6896 (N_6896,N_6782,N_6775);
nand U6897 (N_6897,N_6666,N_6795);
nand U6898 (N_6898,N_6610,N_6684);
nor U6899 (N_6899,N_6714,N_6602);
nand U6900 (N_6900,N_6640,N_6791);
nor U6901 (N_6901,N_6776,N_6793);
xnor U6902 (N_6902,N_6603,N_6635);
nand U6903 (N_6903,N_6661,N_6732);
or U6904 (N_6904,N_6659,N_6746);
or U6905 (N_6905,N_6752,N_6728);
nand U6906 (N_6906,N_6666,N_6744);
and U6907 (N_6907,N_6747,N_6761);
and U6908 (N_6908,N_6636,N_6626);
xor U6909 (N_6909,N_6752,N_6769);
nor U6910 (N_6910,N_6755,N_6685);
nand U6911 (N_6911,N_6700,N_6774);
xnor U6912 (N_6912,N_6622,N_6664);
nand U6913 (N_6913,N_6699,N_6602);
xor U6914 (N_6914,N_6774,N_6617);
nor U6915 (N_6915,N_6625,N_6692);
or U6916 (N_6916,N_6799,N_6678);
or U6917 (N_6917,N_6653,N_6748);
nand U6918 (N_6918,N_6697,N_6764);
nor U6919 (N_6919,N_6741,N_6754);
and U6920 (N_6920,N_6621,N_6673);
nand U6921 (N_6921,N_6700,N_6786);
nor U6922 (N_6922,N_6692,N_6651);
or U6923 (N_6923,N_6687,N_6692);
or U6924 (N_6924,N_6721,N_6737);
and U6925 (N_6925,N_6620,N_6607);
nor U6926 (N_6926,N_6784,N_6641);
and U6927 (N_6927,N_6723,N_6614);
or U6928 (N_6928,N_6685,N_6788);
xnor U6929 (N_6929,N_6619,N_6655);
nor U6930 (N_6930,N_6628,N_6642);
nand U6931 (N_6931,N_6718,N_6723);
and U6932 (N_6932,N_6633,N_6641);
nand U6933 (N_6933,N_6782,N_6712);
or U6934 (N_6934,N_6680,N_6683);
xor U6935 (N_6935,N_6793,N_6612);
or U6936 (N_6936,N_6629,N_6796);
nand U6937 (N_6937,N_6748,N_6605);
nor U6938 (N_6938,N_6640,N_6761);
nand U6939 (N_6939,N_6703,N_6777);
nand U6940 (N_6940,N_6760,N_6619);
xor U6941 (N_6941,N_6633,N_6757);
nor U6942 (N_6942,N_6693,N_6692);
nor U6943 (N_6943,N_6791,N_6675);
nand U6944 (N_6944,N_6752,N_6713);
or U6945 (N_6945,N_6788,N_6698);
nor U6946 (N_6946,N_6710,N_6676);
and U6947 (N_6947,N_6757,N_6778);
nand U6948 (N_6948,N_6743,N_6700);
nand U6949 (N_6949,N_6750,N_6795);
and U6950 (N_6950,N_6621,N_6661);
xor U6951 (N_6951,N_6708,N_6607);
or U6952 (N_6952,N_6657,N_6665);
nand U6953 (N_6953,N_6664,N_6780);
and U6954 (N_6954,N_6790,N_6730);
and U6955 (N_6955,N_6740,N_6623);
and U6956 (N_6956,N_6759,N_6662);
and U6957 (N_6957,N_6777,N_6702);
nand U6958 (N_6958,N_6748,N_6611);
and U6959 (N_6959,N_6670,N_6660);
nand U6960 (N_6960,N_6625,N_6640);
xnor U6961 (N_6961,N_6723,N_6631);
or U6962 (N_6962,N_6707,N_6602);
nand U6963 (N_6963,N_6748,N_6682);
or U6964 (N_6964,N_6743,N_6726);
and U6965 (N_6965,N_6609,N_6779);
xnor U6966 (N_6966,N_6773,N_6712);
and U6967 (N_6967,N_6607,N_6794);
or U6968 (N_6968,N_6776,N_6725);
or U6969 (N_6969,N_6771,N_6607);
xnor U6970 (N_6970,N_6647,N_6759);
nor U6971 (N_6971,N_6716,N_6699);
nor U6972 (N_6972,N_6781,N_6785);
xor U6973 (N_6973,N_6706,N_6665);
nor U6974 (N_6974,N_6713,N_6617);
nor U6975 (N_6975,N_6674,N_6709);
xnor U6976 (N_6976,N_6761,N_6763);
nor U6977 (N_6977,N_6795,N_6689);
and U6978 (N_6978,N_6642,N_6671);
nor U6979 (N_6979,N_6758,N_6735);
and U6980 (N_6980,N_6737,N_6612);
or U6981 (N_6981,N_6773,N_6753);
or U6982 (N_6982,N_6650,N_6666);
and U6983 (N_6983,N_6778,N_6728);
or U6984 (N_6984,N_6767,N_6758);
nor U6985 (N_6985,N_6695,N_6648);
or U6986 (N_6986,N_6799,N_6753);
nand U6987 (N_6987,N_6619,N_6673);
and U6988 (N_6988,N_6629,N_6621);
nand U6989 (N_6989,N_6652,N_6755);
xor U6990 (N_6990,N_6740,N_6726);
nand U6991 (N_6991,N_6645,N_6679);
xnor U6992 (N_6992,N_6706,N_6672);
nand U6993 (N_6993,N_6767,N_6765);
or U6994 (N_6994,N_6755,N_6731);
xor U6995 (N_6995,N_6641,N_6631);
and U6996 (N_6996,N_6742,N_6643);
nand U6997 (N_6997,N_6711,N_6633);
nand U6998 (N_6998,N_6712,N_6682);
xnor U6999 (N_6999,N_6749,N_6670);
or U7000 (N_7000,N_6819,N_6927);
nand U7001 (N_7001,N_6835,N_6985);
xor U7002 (N_7002,N_6931,N_6847);
nor U7003 (N_7003,N_6823,N_6955);
nor U7004 (N_7004,N_6850,N_6887);
or U7005 (N_7005,N_6936,N_6858);
and U7006 (N_7006,N_6893,N_6923);
and U7007 (N_7007,N_6979,N_6908);
nor U7008 (N_7008,N_6922,N_6997);
nand U7009 (N_7009,N_6902,N_6929);
nor U7010 (N_7010,N_6899,N_6951);
or U7011 (N_7011,N_6990,N_6945);
nand U7012 (N_7012,N_6943,N_6926);
and U7013 (N_7013,N_6888,N_6980);
xor U7014 (N_7014,N_6941,N_6813);
and U7015 (N_7015,N_6866,N_6839);
nand U7016 (N_7016,N_6881,N_6965);
xnor U7017 (N_7017,N_6915,N_6801);
nor U7018 (N_7018,N_6934,N_6986);
or U7019 (N_7019,N_6999,N_6960);
nor U7020 (N_7020,N_6844,N_6972);
nand U7021 (N_7021,N_6889,N_6911);
xor U7022 (N_7022,N_6946,N_6851);
xnor U7023 (N_7023,N_6861,N_6831);
nor U7024 (N_7024,N_6803,N_6937);
xnor U7025 (N_7025,N_6935,N_6838);
nor U7026 (N_7026,N_6870,N_6868);
xor U7027 (N_7027,N_6996,N_6959);
nand U7028 (N_7028,N_6932,N_6846);
and U7029 (N_7029,N_6900,N_6871);
or U7030 (N_7030,N_6865,N_6805);
xnor U7031 (N_7031,N_6974,N_6857);
xnor U7032 (N_7032,N_6834,N_6907);
xnor U7033 (N_7033,N_6978,N_6919);
xor U7034 (N_7034,N_6942,N_6944);
or U7035 (N_7035,N_6872,N_6869);
xor U7036 (N_7036,N_6967,N_6895);
nor U7037 (N_7037,N_6879,N_6976);
and U7038 (N_7038,N_6827,N_6949);
nand U7039 (N_7039,N_6892,N_6836);
or U7040 (N_7040,N_6921,N_6817);
or U7041 (N_7041,N_6856,N_6859);
xnor U7042 (N_7042,N_6826,N_6948);
or U7043 (N_7043,N_6940,N_6958);
or U7044 (N_7044,N_6939,N_6977);
xor U7045 (N_7045,N_6989,N_6809);
xnor U7046 (N_7046,N_6909,N_6849);
and U7047 (N_7047,N_6837,N_6961);
or U7048 (N_7048,N_6854,N_6906);
nand U7049 (N_7049,N_6905,N_6933);
or U7050 (N_7050,N_6903,N_6918);
nor U7051 (N_7051,N_6885,N_6842);
xor U7052 (N_7052,N_6828,N_6896);
nor U7053 (N_7053,N_6833,N_6963);
nand U7054 (N_7054,N_6877,N_6822);
nor U7055 (N_7055,N_6832,N_6882);
and U7056 (N_7056,N_6820,N_6966);
nor U7057 (N_7057,N_6925,N_6800);
nand U7058 (N_7058,N_6912,N_6864);
and U7059 (N_7059,N_6901,N_6930);
xor U7060 (N_7060,N_6971,N_6969);
xor U7061 (N_7061,N_6987,N_6910);
and U7062 (N_7062,N_6884,N_6954);
xnor U7063 (N_7063,N_6878,N_6818);
nand U7064 (N_7064,N_6886,N_6862);
or U7065 (N_7065,N_6814,N_6920);
nand U7066 (N_7066,N_6983,N_6897);
nor U7067 (N_7067,N_6880,N_6968);
xnor U7068 (N_7068,N_6916,N_6970);
nor U7069 (N_7069,N_6975,N_6873);
xor U7070 (N_7070,N_6904,N_6840);
nor U7071 (N_7071,N_6876,N_6852);
nor U7072 (N_7072,N_6810,N_6848);
and U7073 (N_7073,N_6988,N_6962);
nor U7074 (N_7074,N_6947,N_6917);
nor U7075 (N_7075,N_6894,N_6995);
and U7076 (N_7076,N_6811,N_6825);
and U7077 (N_7077,N_6824,N_6956);
or U7078 (N_7078,N_6982,N_6841);
and U7079 (N_7079,N_6874,N_6853);
and U7080 (N_7080,N_6928,N_6993);
xnor U7081 (N_7081,N_6860,N_6924);
and U7082 (N_7082,N_6830,N_6891);
or U7083 (N_7083,N_6821,N_6863);
or U7084 (N_7084,N_6802,N_6957);
nor U7085 (N_7085,N_6964,N_6950);
xnor U7086 (N_7086,N_6914,N_6984);
nor U7087 (N_7087,N_6812,N_6807);
nor U7088 (N_7088,N_6898,N_6998);
nor U7089 (N_7089,N_6991,N_6845);
nor U7090 (N_7090,N_6815,N_6981);
xnor U7091 (N_7091,N_6804,N_6883);
and U7092 (N_7092,N_6994,N_6992);
or U7093 (N_7093,N_6829,N_6867);
or U7094 (N_7094,N_6973,N_6855);
nand U7095 (N_7095,N_6913,N_6875);
nor U7096 (N_7096,N_6806,N_6843);
nor U7097 (N_7097,N_6953,N_6816);
xnor U7098 (N_7098,N_6952,N_6890);
nand U7099 (N_7099,N_6938,N_6808);
nand U7100 (N_7100,N_6995,N_6909);
xor U7101 (N_7101,N_6810,N_6861);
xnor U7102 (N_7102,N_6867,N_6814);
or U7103 (N_7103,N_6813,N_6884);
and U7104 (N_7104,N_6970,N_6897);
nor U7105 (N_7105,N_6995,N_6835);
nor U7106 (N_7106,N_6843,N_6829);
nand U7107 (N_7107,N_6825,N_6974);
and U7108 (N_7108,N_6854,N_6862);
or U7109 (N_7109,N_6921,N_6884);
xor U7110 (N_7110,N_6811,N_6994);
nand U7111 (N_7111,N_6997,N_6852);
nand U7112 (N_7112,N_6825,N_6954);
and U7113 (N_7113,N_6998,N_6958);
or U7114 (N_7114,N_6802,N_6974);
or U7115 (N_7115,N_6851,N_6913);
and U7116 (N_7116,N_6913,N_6931);
xnor U7117 (N_7117,N_6992,N_6847);
nand U7118 (N_7118,N_6905,N_6830);
and U7119 (N_7119,N_6961,N_6877);
nand U7120 (N_7120,N_6894,N_6838);
or U7121 (N_7121,N_6812,N_6849);
nor U7122 (N_7122,N_6863,N_6932);
and U7123 (N_7123,N_6900,N_6874);
or U7124 (N_7124,N_6856,N_6917);
and U7125 (N_7125,N_6847,N_6899);
xnor U7126 (N_7126,N_6963,N_6920);
and U7127 (N_7127,N_6813,N_6892);
xor U7128 (N_7128,N_6831,N_6902);
xor U7129 (N_7129,N_6915,N_6996);
nand U7130 (N_7130,N_6963,N_6836);
xnor U7131 (N_7131,N_6831,N_6939);
or U7132 (N_7132,N_6934,N_6971);
nor U7133 (N_7133,N_6823,N_6927);
and U7134 (N_7134,N_6830,N_6946);
nor U7135 (N_7135,N_6800,N_6802);
nor U7136 (N_7136,N_6902,N_6880);
nand U7137 (N_7137,N_6889,N_6906);
or U7138 (N_7138,N_6968,N_6819);
nor U7139 (N_7139,N_6936,N_6927);
xor U7140 (N_7140,N_6980,N_6924);
xnor U7141 (N_7141,N_6961,N_6866);
or U7142 (N_7142,N_6860,N_6917);
and U7143 (N_7143,N_6952,N_6821);
xnor U7144 (N_7144,N_6923,N_6852);
nor U7145 (N_7145,N_6908,N_6826);
nand U7146 (N_7146,N_6815,N_6885);
or U7147 (N_7147,N_6897,N_6826);
and U7148 (N_7148,N_6830,N_6828);
or U7149 (N_7149,N_6973,N_6988);
nor U7150 (N_7150,N_6971,N_6837);
xnor U7151 (N_7151,N_6872,N_6994);
nand U7152 (N_7152,N_6817,N_6927);
nand U7153 (N_7153,N_6879,N_6950);
or U7154 (N_7154,N_6926,N_6952);
nor U7155 (N_7155,N_6859,N_6933);
xor U7156 (N_7156,N_6968,N_6871);
and U7157 (N_7157,N_6821,N_6838);
nor U7158 (N_7158,N_6909,N_6893);
xor U7159 (N_7159,N_6946,N_6877);
nand U7160 (N_7160,N_6827,N_6840);
and U7161 (N_7161,N_6856,N_6891);
nand U7162 (N_7162,N_6900,N_6915);
or U7163 (N_7163,N_6905,N_6904);
nor U7164 (N_7164,N_6983,N_6952);
and U7165 (N_7165,N_6838,N_6933);
xor U7166 (N_7166,N_6926,N_6832);
xnor U7167 (N_7167,N_6998,N_6973);
nor U7168 (N_7168,N_6930,N_6938);
nand U7169 (N_7169,N_6932,N_6878);
or U7170 (N_7170,N_6980,N_6970);
or U7171 (N_7171,N_6814,N_6990);
nor U7172 (N_7172,N_6808,N_6948);
or U7173 (N_7173,N_6820,N_6902);
nand U7174 (N_7174,N_6961,N_6993);
or U7175 (N_7175,N_6832,N_6808);
nand U7176 (N_7176,N_6876,N_6980);
or U7177 (N_7177,N_6989,N_6954);
or U7178 (N_7178,N_6942,N_6930);
and U7179 (N_7179,N_6801,N_6905);
xor U7180 (N_7180,N_6991,N_6807);
or U7181 (N_7181,N_6873,N_6915);
nand U7182 (N_7182,N_6910,N_6966);
or U7183 (N_7183,N_6807,N_6897);
and U7184 (N_7184,N_6921,N_6829);
xnor U7185 (N_7185,N_6854,N_6948);
nor U7186 (N_7186,N_6959,N_6871);
nor U7187 (N_7187,N_6917,N_6916);
nand U7188 (N_7188,N_6898,N_6921);
and U7189 (N_7189,N_6998,N_6893);
and U7190 (N_7190,N_6812,N_6974);
or U7191 (N_7191,N_6892,N_6840);
and U7192 (N_7192,N_6804,N_6869);
nand U7193 (N_7193,N_6932,N_6895);
nand U7194 (N_7194,N_6947,N_6869);
or U7195 (N_7195,N_6862,N_6887);
xor U7196 (N_7196,N_6953,N_6844);
nor U7197 (N_7197,N_6949,N_6917);
nand U7198 (N_7198,N_6950,N_6893);
nand U7199 (N_7199,N_6812,N_6808);
or U7200 (N_7200,N_7109,N_7125);
xnor U7201 (N_7201,N_7132,N_7083);
nor U7202 (N_7202,N_7182,N_7012);
xor U7203 (N_7203,N_7094,N_7003);
xnor U7204 (N_7204,N_7199,N_7146);
or U7205 (N_7205,N_7150,N_7031);
nand U7206 (N_7206,N_7034,N_7063);
nor U7207 (N_7207,N_7194,N_7035);
or U7208 (N_7208,N_7000,N_7127);
xor U7209 (N_7209,N_7015,N_7197);
and U7210 (N_7210,N_7143,N_7129);
or U7211 (N_7211,N_7048,N_7032);
and U7212 (N_7212,N_7160,N_7080);
nand U7213 (N_7213,N_7156,N_7191);
nand U7214 (N_7214,N_7095,N_7178);
or U7215 (N_7215,N_7070,N_7076);
nor U7216 (N_7216,N_7114,N_7198);
or U7217 (N_7217,N_7128,N_7118);
nand U7218 (N_7218,N_7057,N_7061);
nor U7219 (N_7219,N_7002,N_7107);
nand U7220 (N_7220,N_7131,N_7085);
xnor U7221 (N_7221,N_7013,N_7120);
nor U7222 (N_7222,N_7009,N_7110);
or U7223 (N_7223,N_7195,N_7175);
and U7224 (N_7224,N_7078,N_7140);
xor U7225 (N_7225,N_7130,N_7168);
or U7226 (N_7226,N_7186,N_7187);
nor U7227 (N_7227,N_7097,N_7139);
xor U7228 (N_7228,N_7176,N_7027);
nand U7229 (N_7229,N_7006,N_7189);
nand U7230 (N_7230,N_7081,N_7111);
nor U7231 (N_7231,N_7026,N_7045);
and U7232 (N_7232,N_7053,N_7193);
and U7233 (N_7233,N_7166,N_7014);
nand U7234 (N_7234,N_7038,N_7071);
and U7235 (N_7235,N_7105,N_7054);
nand U7236 (N_7236,N_7134,N_7077);
or U7237 (N_7237,N_7161,N_7181);
xor U7238 (N_7238,N_7052,N_7196);
xnor U7239 (N_7239,N_7060,N_7001);
or U7240 (N_7240,N_7135,N_7163);
xnor U7241 (N_7241,N_7041,N_7152);
or U7242 (N_7242,N_7119,N_7157);
or U7243 (N_7243,N_7158,N_7092);
nand U7244 (N_7244,N_7155,N_7117);
xnor U7245 (N_7245,N_7016,N_7018);
xor U7246 (N_7246,N_7147,N_7104);
xnor U7247 (N_7247,N_7180,N_7039);
nor U7248 (N_7248,N_7082,N_7164);
nand U7249 (N_7249,N_7170,N_7144);
nand U7250 (N_7250,N_7086,N_7100);
and U7251 (N_7251,N_7165,N_7112);
and U7252 (N_7252,N_7089,N_7021);
and U7253 (N_7253,N_7159,N_7123);
nor U7254 (N_7254,N_7004,N_7074);
or U7255 (N_7255,N_7066,N_7096);
and U7256 (N_7256,N_7108,N_7087);
nor U7257 (N_7257,N_7093,N_7102);
and U7258 (N_7258,N_7064,N_7029);
nand U7259 (N_7259,N_7044,N_7185);
nand U7260 (N_7260,N_7103,N_7149);
or U7261 (N_7261,N_7024,N_7124);
and U7262 (N_7262,N_7073,N_7042);
nand U7263 (N_7263,N_7058,N_7040);
nor U7264 (N_7264,N_7137,N_7173);
nor U7265 (N_7265,N_7148,N_7153);
or U7266 (N_7266,N_7005,N_7017);
nand U7267 (N_7267,N_7142,N_7033);
nor U7268 (N_7268,N_7169,N_7046);
nand U7269 (N_7269,N_7008,N_7030);
nand U7270 (N_7270,N_7084,N_7101);
nor U7271 (N_7271,N_7098,N_7145);
or U7272 (N_7272,N_7162,N_7067);
xnor U7273 (N_7273,N_7065,N_7036);
xnor U7274 (N_7274,N_7190,N_7072);
and U7275 (N_7275,N_7113,N_7043);
nand U7276 (N_7276,N_7099,N_7037);
nand U7277 (N_7277,N_7126,N_7011);
nand U7278 (N_7278,N_7019,N_7188);
xnor U7279 (N_7279,N_7133,N_7055);
nand U7280 (N_7280,N_7116,N_7088);
nand U7281 (N_7281,N_7141,N_7179);
nor U7282 (N_7282,N_7121,N_7154);
nand U7283 (N_7283,N_7106,N_7183);
or U7284 (N_7284,N_7050,N_7007);
nand U7285 (N_7285,N_7151,N_7172);
and U7286 (N_7286,N_7047,N_7192);
or U7287 (N_7287,N_7023,N_7059);
and U7288 (N_7288,N_7136,N_7184);
or U7289 (N_7289,N_7091,N_7022);
nand U7290 (N_7290,N_7069,N_7056);
or U7291 (N_7291,N_7079,N_7025);
nor U7292 (N_7292,N_7167,N_7028);
xnor U7293 (N_7293,N_7051,N_7090);
nand U7294 (N_7294,N_7171,N_7122);
nor U7295 (N_7295,N_7138,N_7068);
or U7296 (N_7296,N_7020,N_7075);
and U7297 (N_7297,N_7049,N_7062);
nor U7298 (N_7298,N_7115,N_7010);
xor U7299 (N_7299,N_7174,N_7177);
and U7300 (N_7300,N_7144,N_7187);
or U7301 (N_7301,N_7135,N_7191);
xnor U7302 (N_7302,N_7179,N_7171);
nor U7303 (N_7303,N_7043,N_7072);
nor U7304 (N_7304,N_7065,N_7100);
or U7305 (N_7305,N_7093,N_7030);
nor U7306 (N_7306,N_7104,N_7185);
nand U7307 (N_7307,N_7110,N_7012);
or U7308 (N_7308,N_7051,N_7077);
nand U7309 (N_7309,N_7085,N_7169);
xor U7310 (N_7310,N_7184,N_7155);
and U7311 (N_7311,N_7087,N_7130);
or U7312 (N_7312,N_7047,N_7154);
or U7313 (N_7313,N_7167,N_7088);
and U7314 (N_7314,N_7032,N_7135);
and U7315 (N_7315,N_7128,N_7159);
or U7316 (N_7316,N_7047,N_7135);
nand U7317 (N_7317,N_7112,N_7008);
xor U7318 (N_7318,N_7031,N_7070);
or U7319 (N_7319,N_7151,N_7193);
nor U7320 (N_7320,N_7155,N_7157);
and U7321 (N_7321,N_7166,N_7027);
nand U7322 (N_7322,N_7162,N_7074);
and U7323 (N_7323,N_7090,N_7087);
nor U7324 (N_7324,N_7074,N_7154);
nor U7325 (N_7325,N_7029,N_7117);
xor U7326 (N_7326,N_7045,N_7189);
nor U7327 (N_7327,N_7123,N_7065);
nand U7328 (N_7328,N_7094,N_7113);
and U7329 (N_7329,N_7030,N_7102);
and U7330 (N_7330,N_7090,N_7105);
or U7331 (N_7331,N_7002,N_7042);
nand U7332 (N_7332,N_7147,N_7178);
or U7333 (N_7333,N_7029,N_7081);
xor U7334 (N_7334,N_7020,N_7051);
xor U7335 (N_7335,N_7196,N_7035);
xnor U7336 (N_7336,N_7146,N_7050);
or U7337 (N_7337,N_7105,N_7099);
or U7338 (N_7338,N_7010,N_7018);
and U7339 (N_7339,N_7173,N_7114);
or U7340 (N_7340,N_7130,N_7135);
nor U7341 (N_7341,N_7127,N_7089);
xor U7342 (N_7342,N_7135,N_7181);
and U7343 (N_7343,N_7116,N_7000);
or U7344 (N_7344,N_7147,N_7105);
nand U7345 (N_7345,N_7137,N_7073);
nor U7346 (N_7346,N_7046,N_7091);
nor U7347 (N_7347,N_7084,N_7020);
xnor U7348 (N_7348,N_7159,N_7068);
nand U7349 (N_7349,N_7106,N_7006);
nor U7350 (N_7350,N_7047,N_7168);
or U7351 (N_7351,N_7177,N_7182);
nand U7352 (N_7352,N_7075,N_7184);
xnor U7353 (N_7353,N_7113,N_7128);
nor U7354 (N_7354,N_7090,N_7073);
xnor U7355 (N_7355,N_7178,N_7196);
or U7356 (N_7356,N_7193,N_7125);
nor U7357 (N_7357,N_7096,N_7188);
nand U7358 (N_7358,N_7106,N_7009);
nand U7359 (N_7359,N_7104,N_7179);
xor U7360 (N_7360,N_7057,N_7166);
and U7361 (N_7361,N_7100,N_7077);
nor U7362 (N_7362,N_7146,N_7034);
nand U7363 (N_7363,N_7058,N_7060);
nor U7364 (N_7364,N_7030,N_7129);
and U7365 (N_7365,N_7082,N_7105);
and U7366 (N_7366,N_7190,N_7146);
nor U7367 (N_7367,N_7005,N_7111);
xor U7368 (N_7368,N_7007,N_7087);
xor U7369 (N_7369,N_7012,N_7149);
or U7370 (N_7370,N_7048,N_7190);
and U7371 (N_7371,N_7011,N_7185);
nor U7372 (N_7372,N_7147,N_7013);
nor U7373 (N_7373,N_7190,N_7161);
and U7374 (N_7374,N_7052,N_7080);
nor U7375 (N_7375,N_7103,N_7131);
xnor U7376 (N_7376,N_7194,N_7114);
or U7377 (N_7377,N_7013,N_7095);
nand U7378 (N_7378,N_7139,N_7131);
nor U7379 (N_7379,N_7119,N_7049);
nor U7380 (N_7380,N_7077,N_7086);
or U7381 (N_7381,N_7120,N_7192);
xor U7382 (N_7382,N_7013,N_7066);
nand U7383 (N_7383,N_7155,N_7000);
nor U7384 (N_7384,N_7118,N_7080);
nor U7385 (N_7385,N_7007,N_7091);
or U7386 (N_7386,N_7168,N_7029);
nor U7387 (N_7387,N_7117,N_7069);
and U7388 (N_7388,N_7050,N_7128);
and U7389 (N_7389,N_7122,N_7088);
nand U7390 (N_7390,N_7176,N_7186);
or U7391 (N_7391,N_7136,N_7104);
and U7392 (N_7392,N_7025,N_7041);
or U7393 (N_7393,N_7158,N_7058);
or U7394 (N_7394,N_7167,N_7166);
or U7395 (N_7395,N_7111,N_7136);
nand U7396 (N_7396,N_7027,N_7159);
and U7397 (N_7397,N_7170,N_7176);
nand U7398 (N_7398,N_7086,N_7058);
nor U7399 (N_7399,N_7161,N_7196);
or U7400 (N_7400,N_7246,N_7348);
nand U7401 (N_7401,N_7288,N_7290);
or U7402 (N_7402,N_7365,N_7363);
nor U7403 (N_7403,N_7207,N_7219);
or U7404 (N_7404,N_7324,N_7238);
or U7405 (N_7405,N_7320,N_7368);
and U7406 (N_7406,N_7223,N_7367);
xor U7407 (N_7407,N_7251,N_7374);
nor U7408 (N_7408,N_7375,N_7228);
nor U7409 (N_7409,N_7226,N_7258);
or U7410 (N_7410,N_7333,N_7215);
and U7411 (N_7411,N_7329,N_7347);
or U7412 (N_7412,N_7350,N_7237);
nand U7413 (N_7413,N_7201,N_7321);
xnor U7414 (N_7414,N_7345,N_7235);
nor U7415 (N_7415,N_7269,N_7222);
nor U7416 (N_7416,N_7245,N_7311);
or U7417 (N_7417,N_7332,N_7315);
and U7418 (N_7418,N_7309,N_7287);
nor U7419 (N_7419,N_7384,N_7319);
xnor U7420 (N_7420,N_7276,N_7252);
and U7421 (N_7421,N_7386,N_7244);
nand U7422 (N_7422,N_7227,N_7230);
nand U7423 (N_7423,N_7255,N_7385);
nor U7424 (N_7424,N_7229,N_7307);
nor U7425 (N_7425,N_7356,N_7282);
xnor U7426 (N_7426,N_7205,N_7303);
or U7427 (N_7427,N_7317,N_7360);
and U7428 (N_7428,N_7273,N_7259);
xnor U7429 (N_7429,N_7369,N_7373);
nor U7430 (N_7430,N_7262,N_7202);
and U7431 (N_7431,N_7381,N_7275);
nor U7432 (N_7432,N_7279,N_7383);
or U7433 (N_7433,N_7218,N_7323);
nor U7434 (N_7434,N_7220,N_7265);
and U7435 (N_7435,N_7336,N_7289);
nor U7436 (N_7436,N_7300,N_7212);
and U7437 (N_7437,N_7297,N_7340);
nor U7438 (N_7438,N_7210,N_7271);
xnor U7439 (N_7439,N_7310,N_7326);
or U7440 (N_7440,N_7281,N_7388);
nand U7441 (N_7441,N_7301,N_7254);
nand U7442 (N_7442,N_7351,N_7377);
nand U7443 (N_7443,N_7291,N_7380);
xor U7444 (N_7444,N_7308,N_7295);
nand U7445 (N_7445,N_7208,N_7217);
and U7446 (N_7446,N_7357,N_7398);
nor U7447 (N_7447,N_7216,N_7240);
and U7448 (N_7448,N_7200,N_7312);
nand U7449 (N_7449,N_7391,N_7266);
nor U7450 (N_7450,N_7243,N_7305);
nand U7451 (N_7451,N_7392,N_7247);
and U7452 (N_7452,N_7278,N_7270);
nor U7453 (N_7453,N_7304,N_7213);
and U7454 (N_7454,N_7344,N_7327);
xnor U7455 (N_7455,N_7382,N_7358);
xor U7456 (N_7456,N_7296,N_7221);
xor U7457 (N_7457,N_7299,N_7280);
nand U7458 (N_7458,N_7387,N_7359);
nor U7459 (N_7459,N_7274,N_7285);
and U7460 (N_7460,N_7233,N_7314);
xor U7461 (N_7461,N_7372,N_7371);
nor U7462 (N_7462,N_7379,N_7337);
nor U7463 (N_7463,N_7306,N_7263);
xnor U7464 (N_7464,N_7264,N_7354);
nor U7465 (N_7465,N_7267,N_7394);
and U7466 (N_7466,N_7376,N_7396);
or U7467 (N_7467,N_7362,N_7231);
and U7468 (N_7468,N_7204,N_7214);
nand U7469 (N_7469,N_7328,N_7316);
xnor U7470 (N_7470,N_7261,N_7389);
xnor U7471 (N_7471,N_7283,N_7206);
nor U7472 (N_7472,N_7260,N_7342);
xnor U7473 (N_7473,N_7352,N_7395);
xnor U7474 (N_7474,N_7397,N_7313);
nor U7475 (N_7475,N_7343,N_7366);
or U7476 (N_7476,N_7256,N_7225);
xnor U7477 (N_7477,N_7268,N_7298);
or U7478 (N_7478,N_7293,N_7239);
or U7479 (N_7479,N_7234,N_7322);
nor U7480 (N_7480,N_7203,N_7232);
and U7481 (N_7481,N_7339,N_7284);
nand U7482 (N_7482,N_7353,N_7399);
or U7483 (N_7483,N_7209,N_7241);
or U7484 (N_7484,N_7248,N_7378);
or U7485 (N_7485,N_7341,N_7361);
nand U7486 (N_7486,N_7224,N_7302);
or U7487 (N_7487,N_7277,N_7364);
and U7488 (N_7488,N_7292,N_7257);
or U7489 (N_7489,N_7236,N_7330);
nor U7490 (N_7490,N_7390,N_7211);
or U7491 (N_7491,N_7249,N_7334);
xor U7492 (N_7492,N_7286,N_7318);
and U7493 (N_7493,N_7335,N_7370);
xnor U7494 (N_7494,N_7338,N_7253);
nor U7495 (N_7495,N_7325,N_7331);
nand U7496 (N_7496,N_7294,N_7242);
xor U7497 (N_7497,N_7349,N_7346);
or U7498 (N_7498,N_7272,N_7250);
nand U7499 (N_7499,N_7355,N_7393);
or U7500 (N_7500,N_7278,N_7227);
or U7501 (N_7501,N_7389,N_7371);
and U7502 (N_7502,N_7380,N_7336);
nor U7503 (N_7503,N_7329,N_7223);
nand U7504 (N_7504,N_7256,N_7382);
nor U7505 (N_7505,N_7360,N_7334);
nor U7506 (N_7506,N_7363,N_7369);
nor U7507 (N_7507,N_7247,N_7373);
and U7508 (N_7508,N_7324,N_7303);
nor U7509 (N_7509,N_7241,N_7386);
or U7510 (N_7510,N_7318,N_7337);
nand U7511 (N_7511,N_7256,N_7315);
xor U7512 (N_7512,N_7228,N_7387);
nor U7513 (N_7513,N_7284,N_7355);
xor U7514 (N_7514,N_7218,N_7333);
xnor U7515 (N_7515,N_7280,N_7275);
or U7516 (N_7516,N_7388,N_7354);
or U7517 (N_7517,N_7221,N_7247);
nor U7518 (N_7518,N_7358,N_7220);
or U7519 (N_7519,N_7288,N_7235);
or U7520 (N_7520,N_7379,N_7203);
and U7521 (N_7521,N_7318,N_7218);
or U7522 (N_7522,N_7218,N_7293);
or U7523 (N_7523,N_7201,N_7223);
nand U7524 (N_7524,N_7281,N_7253);
nor U7525 (N_7525,N_7237,N_7385);
nand U7526 (N_7526,N_7303,N_7345);
or U7527 (N_7527,N_7239,N_7222);
xor U7528 (N_7528,N_7257,N_7284);
nand U7529 (N_7529,N_7319,N_7388);
and U7530 (N_7530,N_7202,N_7235);
or U7531 (N_7531,N_7321,N_7366);
and U7532 (N_7532,N_7347,N_7378);
nor U7533 (N_7533,N_7281,N_7212);
nand U7534 (N_7534,N_7339,N_7253);
and U7535 (N_7535,N_7200,N_7262);
xor U7536 (N_7536,N_7379,N_7312);
or U7537 (N_7537,N_7224,N_7212);
or U7538 (N_7538,N_7331,N_7330);
xnor U7539 (N_7539,N_7335,N_7350);
xnor U7540 (N_7540,N_7364,N_7308);
nand U7541 (N_7541,N_7342,N_7257);
or U7542 (N_7542,N_7240,N_7241);
or U7543 (N_7543,N_7234,N_7373);
or U7544 (N_7544,N_7206,N_7236);
and U7545 (N_7545,N_7253,N_7372);
nor U7546 (N_7546,N_7364,N_7233);
or U7547 (N_7547,N_7331,N_7200);
nor U7548 (N_7548,N_7332,N_7351);
and U7549 (N_7549,N_7374,N_7358);
nand U7550 (N_7550,N_7351,N_7376);
nand U7551 (N_7551,N_7383,N_7288);
nor U7552 (N_7552,N_7224,N_7326);
and U7553 (N_7553,N_7295,N_7218);
xnor U7554 (N_7554,N_7222,N_7309);
xor U7555 (N_7555,N_7236,N_7359);
xnor U7556 (N_7556,N_7399,N_7300);
nand U7557 (N_7557,N_7248,N_7336);
or U7558 (N_7558,N_7315,N_7271);
nor U7559 (N_7559,N_7205,N_7337);
nor U7560 (N_7560,N_7289,N_7364);
and U7561 (N_7561,N_7373,N_7308);
xor U7562 (N_7562,N_7389,N_7315);
xnor U7563 (N_7563,N_7388,N_7269);
or U7564 (N_7564,N_7231,N_7399);
and U7565 (N_7565,N_7362,N_7268);
nand U7566 (N_7566,N_7360,N_7379);
nand U7567 (N_7567,N_7268,N_7334);
xor U7568 (N_7568,N_7362,N_7247);
nand U7569 (N_7569,N_7206,N_7391);
nand U7570 (N_7570,N_7219,N_7350);
nand U7571 (N_7571,N_7341,N_7377);
or U7572 (N_7572,N_7344,N_7337);
xnor U7573 (N_7573,N_7330,N_7286);
or U7574 (N_7574,N_7314,N_7245);
nor U7575 (N_7575,N_7334,N_7269);
nand U7576 (N_7576,N_7284,N_7383);
and U7577 (N_7577,N_7365,N_7210);
nand U7578 (N_7578,N_7319,N_7230);
xor U7579 (N_7579,N_7333,N_7316);
and U7580 (N_7580,N_7231,N_7294);
or U7581 (N_7581,N_7307,N_7398);
and U7582 (N_7582,N_7239,N_7298);
xnor U7583 (N_7583,N_7232,N_7324);
nand U7584 (N_7584,N_7257,N_7258);
xnor U7585 (N_7585,N_7322,N_7276);
nor U7586 (N_7586,N_7378,N_7264);
nor U7587 (N_7587,N_7211,N_7336);
or U7588 (N_7588,N_7260,N_7353);
nand U7589 (N_7589,N_7285,N_7220);
nor U7590 (N_7590,N_7214,N_7241);
and U7591 (N_7591,N_7213,N_7263);
nand U7592 (N_7592,N_7360,N_7358);
nor U7593 (N_7593,N_7292,N_7326);
xor U7594 (N_7594,N_7298,N_7330);
nor U7595 (N_7595,N_7218,N_7382);
xor U7596 (N_7596,N_7338,N_7207);
and U7597 (N_7597,N_7272,N_7210);
and U7598 (N_7598,N_7340,N_7291);
or U7599 (N_7599,N_7232,N_7339);
nor U7600 (N_7600,N_7571,N_7434);
and U7601 (N_7601,N_7495,N_7568);
and U7602 (N_7602,N_7575,N_7456);
nor U7603 (N_7603,N_7570,N_7523);
xor U7604 (N_7604,N_7479,N_7553);
xnor U7605 (N_7605,N_7594,N_7518);
and U7606 (N_7606,N_7593,N_7535);
xor U7607 (N_7607,N_7406,N_7443);
nor U7608 (N_7608,N_7449,N_7522);
nand U7609 (N_7609,N_7559,N_7428);
and U7610 (N_7610,N_7563,N_7551);
xnor U7611 (N_7611,N_7521,N_7595);
xnor U7612 (N_7612,N_7576,N_7539);
xor U7613 (N_7613,N_7425,N_7515);
nand U7614 (N_7614,N_7466,N_7492);
xor U7615 (N_7615,N_7436,N_7582);
nand U7616 (N_7616,N_7459,N_7565);
nand U7617 (N_7617,N_7526,N_7411);
nand U7618 (N_7618,N_7502,N_7550);
and U7619 (N_7619,N_7421,N_7536);
xor U7620 (N_7620,N_7572,N_7438);
xor U7621 (N_7621,N_7498,N_7566);
or U7622 (N_7622,N_7497,N_7440);
or U7623 (N_7623,N_7400,N_7417);
xor U7624 (N_7624,N_7410,N_7501);
nand U7625 (N_7625,N_7591,N_7562);
or U7626 (N_7626,N_7533,N_7488);
nand U7627 (N_7627,N_7464,N_7445);
nor U7628 (N_7628,N_7493,N_7460);
nor U7629 (N_7629,N_7403,N_7473);
or U7630 (N_7630,N_7580,N_7467);
and U7631 (N_7631,N_7447,N_7404);
and U7632 (N_7632,N_7454,N_7474);
and U7633 (N_7633,N_7499,N_7458);
nand U7634 (N_7634,N_7418,N_7435);
or U7635 (N_7635,N_7446,N_7416);
nand U7636 (N_7636,N_7525,N_7412);
or U7637 (N_7637,N_7481,N_7577);
and U7638 (N_7638,N_7484,N_7511);
nor U7639 (N_7639,N_7527,N_7503);
nor U7640 (N_7640,N_7509,N_7487);
or U7641 (N_7641,N_7544,N_7452);
and U7642 (N_7642,N_7524,N_7538);
nand U7643 (N_7643,N_7437,N_7426);
or U7644 (N_7644,N_7472,N_7468);
nor U7645 (N_7645,N_7429,N_7541);
nand U7646 (N_7646,N_7424,N_7549);
xnor U7647 (N_7647,N_7587,N_7537);
nand U7648 (N_7648,N_7442,N_7494);
nand U7649 (N_7649,N_7598,N_7457);
nor U7650 (N_7650,N_7554,N_7433);
or U7651 (N_7651,N_7486,N_7530);
or U7652 (N_7652,N_7470,N_7430);
and U7653 (N_7653,N_7439,N_7561);
nor U7654 (N_7654,N_7422,N_7547);
nand U7655 (N_7655,N_7556,N_7508);
nand U7656 (N_7656,N_7490,N_7528);
or U7657 (N_7657,N_7504,N_7405);
nor U7658 (N_7658,N_7564,N_7461);
or U7659 (N_7659,N_7529,N_7574);
and U7660 (N_7660,N_7427,N_7597);
nand U7661 (N_7661,N_7542,N_7478);
and U7662 (N_7662,N_7599,N_7489);
nor U7663 (N_7663,N_7402,N_7476);
xor U7664 (N_7664,N_7413,N_7555);
or U7665 (N_7665,N_7540,N_7414);
and U7666 (N_7666,N_7420,N_7465);
xor U7667 (N_7667,N_7480,N_7408);
or U7668 (N_7668,N_7471,N_7507);
xnor U7669 (N_7669,N_7512,N_7482);
or U7670 (N_7670,N_7506,N_7589);
nand U7671 (N_7671,N_7432,N_7453);
or U7672 (N_7672,N_7573,N_7516);
nand U7673 (N_7673,N_7548,N_7531);
or U7674 (N_7674,N_7514,N_7462);
and U7675 (N_7675,N_7552,N_7532);
xnor U7676 (N_7676,N_7444,N_7448);
or U7677 (N_7677,N_7578,N_7546);
nand U7678 (N_7678,N_7579,N_7505);
xnor U7679 (N_7679,N_7517,N_7431);
nand U7680 (N_7680,N_7519,N_7401);
xnor U7681 (N_7681,N_7500,N_7451);
or U7682 (N_7682,N_7584,N_7485);
or U7683 (N_7683,N_7567,N_7409);
or U7684 (N_7684,N_7534,N_7423);
or U7685 (N_7685,N_7585,N_7491);
xnor U7686 (N_7686,N_7590,N_7583);
or U7687 (N_7687,N_7513,N_7586);
xnor U7688 (N_7688,N_7455,N_7415);
nor U7689 (N_7689,N_7545,N_7510);
xor U7690 (N_7690,N_7569,N_7592);
xnor U7691 (N_7691,N_7450,N_7469);
nor U7692 (N_7692,N_7557,N_7441);
xor U7693 (N_7693,N_7558,N_7483);
nor U7694 (N_7694,N_7419,N_7477);
or U7695 (N_7695,N_7475,N_7596);
xor U7696 (N_7696,N_7581,N_7520);
and U7697 (N_7697,N_7407,N_7496);
nor U7698 (N_7698,N_7463,N_7588);
nor U7699 (N_7699,N_7560,N_7543);
or U7700 (N_7700,N_7470,N_7433);
nand U7701 (N_7701,N_7530,N_7406);
and U7702 (N_7702,N_7523,N_7464);
nand U7703 (N_7703,N_7425,N_7479);
nor U7704 (N_7704,N_7448,N_7452);
nand U7705 (N_7705,N_7430,N_7406);
nor U7706 (N_7706,N_7560,N_7420);
and U7707 (N_7707,N_7555,N_7412);
xnor U7708 (N_7708,N_7596,N_7458);
nand U7709 (N_7709,N_7473,N_7523);
xnor U7710 (N_7710,N_7585,N_7542);
xor U7711 (N_7711,N_7484,N_7516);
xnor U7712 (N_7712,N_7590,N_7423);
and U7713 (N_7713,N_7580,N_7530);
and U7714 (N_7714,N_7557,N_7456);
nand U7715 (N_7715,N_7400,N_7501);
nor U7716 (N_7716,N_7491,N_7409);
and U7717 (N_7717,N_7446,N_7597);
nor U7718 (N_7718,N_7547,N_7569);
xnor U7719 (N_7719,N_7572,N_7587);
xnor U7720 (N_7720,N_7435,N_7547);
or U7721 (N_7721,N_7572,N_7440);
and U7722 (N_7722,N_7564,N_7479);
nor U7723 (N_7723,N_7448,N_7506);
and U7724 (N_7724,N_7432,N_7478);
and U7725 (N_7725,N_7500,N_7447);
xnor U7726 (N_7726,N_7420,N_7562);
nand U7727 (N_7727,N_7550,N_7547);
nand U7728 (N_7728,N_7449,N_7581);
nand U7729 (N_7729,N_7568,N_7539);
or U7730 (N_7730,N_7577,N_7480);
xnor U7731 (N_7731,N_7448,N_7413);
nor U7732 (N_7732,N_7450,N_7583);
or U7733 (N_7733,N_7459,N_7591);
xor U7734 (N_7734,N_7522,N_7480);
or U7735 (N_7735,N_7547,N_7400);
and U7736 (N_7736,N_7557,N_7483);
nor U7737 (N_7737,N_7446,N_7454);
nor U7738 (N_7738,N_7446,N_7453);
or U7739 (N_7739,N_7491,N_7541);
nand U7740 (N_7740,N_7551,N_7436);
nand U7741 (N_7741,N_7581,N_7477);
and U7742 (N_7742,N_7532,N_7586);
nand U7743 (N_7743,N_7538,N_7407);
nand U7744 (N_7744,N_7457,N_7510);
nor U7745 (N_7745,N_7520,N_7458);
nand U7746 (N_7746,N_7517,N_7528);
nor U7747 (N_7747,N_7574,N_7493);
nand U7748 (N_7748,N_7449,N_7535);
xnor U7749 (N_7749,N_7414,N_7476);
nor U7750 (N_7750,N_7555,N_7501);
nand U7751 (N_7751,N_7434,N_7477);
xor U7752 (N_7752,N_7429,N_7551);
nor U7753 (N_7753,N_7505,N_7464);
xor U7754 (N_7754,N_7593,N_7594);
nand U7755 (N_7755,N_7502,N_7544);
xor U7756 (N_7756,N_7421,N_7443);
or U7757 (N_7757,N_7450,N_7477);
nand U7758 (N_7758,N_7497,N_7519);
and U7759 (N_7759,N_7471,N_7544);
and U7760 (N_7760,N_7552,N_7470);
xnor U7761 (N_7761,N_7486,N_7418);
and U7762 (N_7762,N_7450,N_7570);
and U7763 (N_7763,N_7561,N_7498);
and U7764 (N_7764,N_7525,N_7485);
nor U7765 (N_7765,N_7591,N_7582);
and U7766 (N_7766,N_7507,N_7453);
and U7767 (N_7767,N_7444,N_7530);
nand U7768 (N_7768,N_7596,N_7442);
xnor U7769 (N_7769,N_7561,N_7517);
xnor U7770 (N_7770,N_7510,N_7466);
xor U7771 (N_7771,N_7566,N_7553);
or U7772 (N_7772,N_7411,N_7404);
nor U7773 (N_7773,N_7544,N_7442);
nand U7774 (N_7774,N_7461,N_7488);
nand U7775 (N_7775,N_7504,N_7414);
xnor U7776 (N_7776,N_7550,N_7492);
or U7777 (N_7777,N_7511,N_7469);
xor U7778 (N_7778,N_7450,N_7448);
xor U7779 (N_7779,N_7481,N_7594);
nor U7780 (N_7780,N_7447,N_7499);
nor U7781 (N_7781,N_7444,N_7472);
xnor U7782 (N_7782,N_7514,N_7494);
or U7783 (N_7783,N_7452,N_7541);
nor U7784 (N_7784,N_7597,N_7418);
nand U7785 (N_7785,N_7589,N_7550);
nand U7786 (N_7786,N_7532,N_7512);
and U7787 (N_7787,N_7447,N_7562);
or U7788 (N_7788,N_7401,N_7516);
and U7789 (N_7789,N_7498,N_7425);
and U7790 (N_7790,N_7514,N_7568);
and U7791 (N_7791,N_7567,N_7416);
and U7792 (N_7792,N_7583,N_7491);
xnor U7793 (N_7793,N_7486,N_7522);
xnor U7794 (N_7794,N_7487,N_7485);
and U7795 (N_7795,N_7485,N_7583);
nand U7796 (N_7796,N_7406,N_7487);
or U7797 (N_7797,N_7572,N_7531);
xnor U7798 (N_7798,N_7585,N_7430);
and U7799 (N_7799,N_7596,N_7542);
xor U7800 (N_7800,N_7773,N_7727);
or U7801 (N_7801,N_7652,N_7707);
nor U7802 (N_7802,N_7708,N_7699);
nand U7803 (N_7803,N_7644,N_7697);
or U7804 (N_7804,N_7758,N_7687);
and U7805 (N_7805,N_7779,N_7756);
and U7806 (N_7806,N_7767,N_7615);
nand U7807 (N_7807,N_7729,N_7704);
xor U7808 (N_7808,N_7663,N_7744);
xnor U7809 (N_7809,N_7765,N_7701);
or U7810 (N_7810,N_7761,N_7664);
and U7811 (N_7811,N_7705,N_7629);
xnor U7812 (N_7812,N_7753,N_7624);
nand U7813 (N_7813,N_7643,N_7711);
or U7814 (N_7814,N_7741,N_7619);
and U7815 (N_7815,N_7608,N_7791);
or U7816 (N_7816,N_7734,N_7649);
and U7817 (N_7817,N_7690,N_7626);
or U7818 (N_7818,N_7755,N_7654);
nand U7819 (N_7819,N_7787,N_7634);
or U7820 (N_7820,N_7674,N_7722);
nand U7821 (N_7821,N_7723,N_7766);
or U7822 (N_7822,N_7647,N_7694);
nor U7823 (N_7823,N_7743,N_7648);
and U7824 (N_7824,N_7782,N_7739);
nor U7825 (N_7825,N_7622,N_7712);
nand U7826 (N_7826,N_7631,N_7784);
xnor U7827 (N_7827,N_7688,N_7798);
or U7828 (N_7828,N_7680,N_7627);
and U7829 (N_7829,N_7632,N_7630);
nor U7830 (N_7830,N_7611,N_7736);
nand U7831 (N_7831,N_7796,N_7786);
and U7832 (N_7832,N_7726,N_7793);
nor U7833 (N_7833,N_7660,N_7760);
or U7834 (N_7834,N_7702,N_7716);
nor U7835 (N_7835,N_7692,N_7733);
or U7836 (N_7836,N_7745,N_7613);
or U7837 (N_7837,N_7651,N_7730);
nand U7838 (N_7838,N_7724,N_7768);
nand U7839 (N_7839,N_7686,N_7637);
and U7840 (N_7840,N_7763,N_7728);
nor U7841 (N_7841,N_7754,N_7602);
nand U7842 (N_7842,N_7625,N_7703);
or U7843 (N_7843,N_7683,N_7670);
nand U7844 (N_7844,N_7689,N_7742);
nand U7845 (N_7845,N_7770,N_7789);
nand U7846 (N_7846,N_7673,N_7678);
xor U7847 (N_7847,N_7646,N_7696);
nand U7848 (N_7848,N_7671,N_7628);
nand U7849 (N_7849,N_7623,N_7693);
and U7850 (N_7850,N_7620,N_7797);
xnor U7851 (N_7851,N_7601,N_7607);
xor U7852 (N_7852,N_7679,N_7667);
and U7853 (N_7853,N_7783,N_7788);
nor U7854 (N_7854,N_7609,N_7762);
or U7855 (N_7855,N_7617,N_7621);
xor U7856 (N_7856,N_7672,N_7605);
or U7857 (N_7857,N_7792,N_7706);
nor U7858 (N_7858,N_7700,N_7769);
and U7859 (N_7859,N_7731,N_7669);
nor U7860 (N_7860,N_7655,N_7650);
xnor U7861 (N_7861,N_7799,N_7633);
or U7862 (N_7862,N_7748,N_7618);
xnor U7863 (N_7863,N_7616,N_7676);
or U7864 (N_7864,N_7720,N_7719);
xor U7865 (N_7865,N_7685,N_7738);
xnor U7866 (N_7866,N_7638,N_7750);
nand U7867 (N_7867,N_7603,N_7732);
or U7868 (N_7868,N_7635,N_7777);
nand U7869 (N_7869,N_7653,N_7721);
and U7870 (N_7870,N_7642,N_7610);
nor U7871 (N_7871,N_7764,N_7640);
and U7872 (N_7872,N_7639,N_7606);
nor U7873 (N_7873,N_7675,N_7775);
nand U7874 (N_7874,N_7668,N_7600);
and U7875 (N_7875,N_7781,N_7661);
xor U7876 (N_7876,N_7659,N_7656);
nor U7877 (N_7877,N_7771,N_7698);
nor U7878 (N_7878,N_7785,N_7662);
and U7879 (N_7879,N_7776,N_7735);
or U7880 (N_7880,N_7752,N_7658);
xnor U7881 (N_7881,N_7737,N_7695);
and U7882 (N_7882,N_7612,N_7657);
nor U7883 (N_7883,N_7725,N_7717);
xnor U7884 (N_7884,N_7718,N_7759);
nand U7885 (N_7885,N_7681,N_7780);
nand U7886 (N_7886,N_7746,N_7772);
and U7887 (N_7887,N_7709,N_7636);
nor U7888 (N_7888,N_7740,N_7795);
or U7889 (N_7889,N_7790,N_7778);
or U7890 (N_7890,N_7604,N_7682);
or U7891 (N_7891,N_7774,N_7641);
xor U7892 (N_7892,N_7614,N_7747);
or U7893 (N_7893,N_7710,N_7713);
or U7894 (N_7894,N_7666,N_7715);
nand U7895 (N_7895,N_7677,N_7749);
nor U7896 (N_7896,N_7714,N_7665);
nand U7897 (N_7897,N_7757,N_7794);
xor U7898 (N_7898,N_7691,N_7645);
or U7899 (N_7899,N_7684,N_7751);
xnor U7900 (N_7900,N_7798,N_7780);
and U7901 (N_7901,N_7735,N_7602);
xnor U7902 (N_7902,N_7615,N_7756);
nand U7903 (N_7903,N_7787,N_7786);
nand U7904 (N_7904,N_7644,N_7658);
nand U7905 (N_7905,N_7758,N_7757);
xnor U7906 (N_7906,N_7768,N_7786);
nand U7907 (N_7907,N_7794,N_7746);
xor U7908 (N_7908,N_7652,N_7788);
and U7909 (N_7909,N_7784,N_7673);
or U7910 (N_7910,N_7725,N_7683);
nand U7911 (N_7911,N_7729,N_7714);
xnor U7912 (N_7912,N_7764,N_7627);
xor U7913 (N_7913,N_7673,N_7785);
xnor U7914 (N_7914,N_7785,N_7754);
and U7915 (N_7915,N_7613,N_7641);
or U7916 (N_7916,N_7612,N_7682);
or U7917 (N_7917,N_7696,N_7615);
nand U7918 (N_7918,N_7686,N_7623);
or U7919 (N_7919,N_7646,N_7637);
nor U7920 (N_7920,N_7780,N_7781);
nor U7921 (N_7921,N_7699,N_7621);
and U7922 (N_7922,N_7668,N_7690);
nand U7923 (N_7923,N_7609,N_7698);
nor U7924 (N_7924,N_7609,N_7660);
or U7925 (N_7925,N_7761,N_7658);
or U7926 (N_7926,N_7743,N_7777);
and U7927 (N_7927,N_7795,N_7746);
nand U7928 (N_7928,N_7706,N_7784);
xor U7929 (N_7929,N_7785,N_7784);
or U7930 (N_7930,N_7673,N_7796);
nand U7931 (N_7931,N_7641,N_7603);
and U7932 (N_7932,N_7727,N_7673);
nand U7933 (N_7933,N_7631,N_7720);
xnor U7934 (N_7934,N_7738,N_7699);
nor U7935 (N_7935,N_7602,N_7601);
nand U7936 (N_7936,N_7793,N_7666);
xnor U7937 (N_7937,N_7792,N_7649);
and U7938 (N_7938,N_7662,N_7795);
or U7939 (N_7939,N_7686,N_7785);
xor U7940 (N_7940,N_7684,N_7710);
xor U7941 (N_7941,N_7774,N_7692);
nor U7942 (N_7942,N_7686,N_7607);
or U7943 (N_7943,N_7739,N_7795);
xnor U7944 (N_7944,N_7700,N_7786);
nand U7945 (N_7945,N_7680,N_7719);
nor U7946 (N_7946,N_7718,N_7791);
and U7947 (N_7947,N_7699,N_7615);
xor U7948 (N_7948,N_7781,N_7649);
xor U7949 (N_7949,N_7695,N_7652);
or U7950 (N_7950,N_7609,N_7791);
or U7951 (N_7951,N_7680,N_7603);
nand U7952 (N_7952,N_7735,N_7665);
nand U7953 (N_7953,N_7716,N_7733);
and U7954 (N_7954,N_7689,N_7725);
and U7955 (N_7955,N_7782,N_7784);
and U7956 (N_7956,N_7765,N_7792);
nand U7957 (N_7957,N_7763,N_7784);
xor U7958 (N_7958,N_7685,N_7674);
nor U7959 (N_7959,N_7603,N_7672);
nand U7960 (N_7960,N_7768,N_7796);
nor U7961 (N_7961,N_7645,N_7646);
and U7962 (N_7962,N_7674,N_7667);
xnor U7963 (N_7963,N_7700,N_7624);
and U7964 (N_7964,N_7687,N_7734);
nor U7965 (N_7965,N_7714,N_7628);
nand U7966 (N_7966,N_7784,N_7676);
and U7967 (N_7967,N_7729,N_7673);
or U7968 (N_7968,N_7741,N_7646);
or U7969 (N_7969,N_7775,N_7710);
nor U7970 (N_7970,N_7609,N_7757);
or U7971 (N_7971,N_7744,N_7785);
or U7972 (N_7972,N_7768,N_7755);
nor U7973 (N_7973,N_7610,N_7723);
or U7974 (N_7974,N_7750,N_7633);
and U7975 (N_7975,N_7708,N_7652);
xnor U7976 (N_7976,N_7692,N_7797);
nor U7977 (N_7977,N_7640,N_7636);
xor U7978 (N_7978,N_7642,N_7735);
nand U7979 (N_7979,N_7660,N_7615);
and U7980 (N_7980,N_7663,N_7714);
nor U7981 (N_7981,N_7633,N_7790);
or U7982 (N_7982,N_7712,N_7653);
and U7983 (N_7983,N_7704,N_7775);
xnor U7984 (N_7984,N_7761,N_7789);
nor U7985 (N_7985,N_7718,N_7617);
nor U7986 (N_7986,N_7780,N_7733);
and U7987 (N_7987,N_7650,N_7773);
nor U7988 (N_7988,N_7697,N_7778);
and U7989 (N_7989,N_7682,N_7611);
and U7990 (N_7990,N_7793,N_7619);
or U7991 (N_7991,N_7797,N_7796);
nand U7992 (N_7992,N_7691,N_7678);
or U7993 (N_7993,N_7798,N_7603);
nor U7994 (N_7994,N_7603,N_7697);
nand U7995 (N_7995,N_7723,N_7617);
nor U7996 (N_7996,N_7762,N_7777);
and U7997 (N_7997,N_7608,N_7762);
nand U7998 (N_7998,N_7748,N_7753);
or U7999 (N_7999,N_7690,N_7636);
xor U8000 (N_8000,N_7996,N_7814);
nor U8001 (N_8001,N_7987,N_7958);
nor U8002 (N_8002,N_7990,N_7992);
and U8003 (N_8003,N_7913,N_7827);
and U8004 (N_8004,N_7875,N_7868);
nand U8005 (N_8005,N_7872,N_7835);
xnor U8006 (N_8006,N_7993,N_7801);
nor U8007 (N_8007,N_7809,N_7943);
nor U8008 (N_8008,N_7976,N_7933);
xnor U8009 (N_8009,N_7966,N_7876);
nor U8010 (N_8010,N_7956,N_7911);
nand U8011 (N_8011,N_7923,N_7982);
or U8012 (N_8012,N_7878,N_7959);
nor U8013 (N_8013,N_7965,N_7852);
xor U8014 (N_8014,N_7877,N_7915);
or U8015 (N_8015,N_7845,N_7887);
xnor U8016 (N_8016,N_7816,N_7847);
nor U8017 (N_8017,N_7984,N_7920);
nand U8018 (N_8018,N_7999,N_7804);
and U8019 (N_8019,N_7865,N_7897);
nor U8020 (N_8020,N_7994,N_7997);
xnor U8021 (N_8021,N_7922,N_7889);
xnor U8022 (N_8022,N_7867,N_7926);
nand U8023 (N_8023,N_7942,N_7960);
nand U8024 (N_8024,N_7813,N_7885);
or U8025 (N_8025,N_7921,N_7907);
nor U8026 (N_8026,N_7856,N_7928);
nand U8027 (N_8027,N_7914,N_7981);
nor U8028 (N_8028,N_7910,N_7961);
or U8029 (N_8029,N_7912,N_7930);
nand U8030 (N_8030,N_7833,N_7846);
and U8031 (N_8031,N_7870,N_7843);
nand U8032 (N_8032,N_7848,N_7851);
or U8033 (N_8033,N_7844,N_7849);
and U8034 (N_8034,N_7803,N_7939);
xor U8035 (N_8035,N_7919,N_7881);
nor U8036 (N_8036,N_7973,N_7941);
xnor U8037 (N_8037,N_7900,N_7892);
xnor U8038 (N_8038,N_7904,N_7972);
or U8039 (N_8039,N_7879,N_7883);
nand U8040 (N_8040,N_7838,N_7829);
nand U8041 (N_8041,N_7975,N_7974);
and U8042 (N_8042,N_7986,N_7950);
or U8043 (N_8043,N_7998,N_7896);
nor U8044 (N_8044,N_7839,N_7812);
nor U8045 (N_8045,N_7822,N_7924);
and U8046 (N_8046,N_7902,N_7891);
nand U8047 (N_8047,N_7931,N_7862);
or U8048 (N_8048,N_7895,N_7890);
and U8049 (N_8049,N_7906,N_7898);
nor U8050 (N_8050,N_7825,N_7935);
nor U8051 (N_8051,N_7936,N_7841);
and U8052 (N_8052,N_7916,N_7944);
nand U8053 (N_8053,N_7854,N_7991);
nor U8054 (N_8054,N_7925,N_7828);
xor U8055 (N_8055,N_7945,N_7858);
and U8056 (N_8056,N_7929,N_7908);
nor U8057 (N_8057,N_7983,N_7882);
or U8058 (N_8058,N_7899,N_7818);
or U8059 (N_8059,N_7863,N_7927);
or U8060 (N_8060,N_7819,N_7861);
or U8061 (N_8061,N_7810,N_7864);
nor U8062 (N_8062,N_7824,N_7970);
or U8063 (N_8063,N_7903,N_7817);
nor U8064 (N_8064,N_7980,N_7869);
and U8065 (N_8065,N_7962,N_7918);
xnor U8066 (N_8066,N_7946,N_7808);
or U8067 (N_8067,N_7859,N_7953);
nor U8068 (N_8068,N_7871,N_7947);
or U8069 (N_8069,N_7886,N_7917);
or U8070 (N_8070,N_7971,N_7909);
nor U8071 (N_8071,N_7855,N_7954);
nand U8072 (N_8072,N_7938,N_7949);
and U8073 (N_8073,N_7951,N_7989);
or U8074 (N_8074,N_7830,N_7940);
nand U8075 (N_8075,N_7880,N_7837);
xor U8076 (N_8076,N_7932,N_7952);
xor U8077 (N_8077,N_7826,N_7957);
and U8078 (N_8078,N_7857,N_7995);
nand U8079 (N_8079,N_7836,N_7831);
and U8080 (N_8080,N_7964,N_7866);
nand U8081 (N_8081,N_7834,N_7821);
nand U8082 (N_8082,N_7805,N_7888);
nand U8083 (N_8083,N_7967,N_7905);
xor U8084 (N_8084,N_7800,N_7894);
and U8085 (N_8085,N_7901,N_7874);
nand U8086 (N_8086,N_7937,N_7955);
nor U8087 (N_8087,N_7806,N_7820);
xor U8088 (N_8088,N_7884,N_7815);
nand U8089 (N_8089,N_7842,N_7979);
and U8090 (N_8090,N_7823,N_7968);
and U8091 (N_8091,N_7850,N_7802);
or U8092 (N_8092,N_7977,N_7873);
nand U8093 (N_8093,N_7893,N_7860);
and U8094 (N_8094,N_7948,N_7934);
and U8095 (N_8095,N_7963,N_7988);
and U8096 (N_8096,N_7969,N_7807);
nand U8097 (N_8097,N_7978,N_7840);
and U8098 (N_8098,N_7832,N_7985);
xnor U8099 (N_8099,N_7811,N_7853);
and U8100 (N_8100,N_7889,N_7872);
or U8101 (N_8101,N_7880,N_7956);
and U8102 (N_8102,N_7963,N_7816);
nor U8103 (N_8103,N_7808,N_7840);
and U8104 (N_8104,N_7943,N_7959);
nor U8105 (N_8105,N_7818,N_7801);
nand U8106 (N_8106,N_7830,N_7973);
or U8107 (N_8107,N_7893,N_7949);
nand U8108 (N_8108,N_7827,N_7929);
or U8109 (N_8109,N_7998,N_7856);
nor U8110 (N_8110,N_7968,N_7936);
xnor U8111 (N_8111,N_7920,N_7998);
nand U8112 (N_8112,N_7949,N_7806);
and U8113 (N_8113,N_7975,N_7968);
nor U8114 (N_8114,N_7817,N_7829);
nor U8115 (N_8115,N_7961,N_7860);
and U8116 (N_8116,N_7818,N_7891);
or U8117 (N_8117,N_7939,N_7908);
nand U8118 (N_8118,N_7838,N_7840);
xor U8119 (N_8119,N_7936,N_7960);
and U8120 (N_8120,N_7991,N_7806);
or U8121 (N_8121,N_7868,N_7985);
or U8122 (N_8122,N_7924,N_7949);
and U8123 (N_8123,N_7875,N_7913);
xnor U8124 (N_8124,N_7831,N_7902);
nor U8125 (N_8125,N_7997,N_7938);
nor U8126 (N_8126,N_7831,N_7811);
and U8127 (N_8127,N_7836,N_7859);
xor U8128 (N_8128,N_7955,N_7915);
nor U8129 (N_8129,N_7878,N_7989);
or U8130 (N_8130,N_7829,N_7971);
nor U8131 (N_8131,N_7939,N_7951);
nor U8132 (N_8132,N_7816,N_7886);
xor U8133 (N_8133,N_7933,N_7814);
xnor U8134 (N_8134,N_7813,N_7900);
or U8135 (N_8135,N_7926,N_7998);
nor U8136 (N_8136,N_7917,N_7810);
nor U8137 (N_8137,N_7997,N_7849);
nor U8138 (N_8138,N_7805,N_7901);
xnor U8139 (N_8139,N_7825,N_7910);
and U8140 (N_8140,N_7932,N_7867);
nor U8141 (N_8141,N_7910,N_7841);
nand U8142 (N_8142,N_7903,N_7913);
and U8143 (N_8143,N_7917,N_7895);
and U8144 (N_8144,N_7854,N_7813);
nor U8145 (N_8145,N_7850,N_7917);
nor U8146 (N_8146,N_7890,N_7918);
and U8147 (N_8147,N_7989,N_7835);
nand U8148 (N_8148,N_7990,N_7939);
nor U8149 (N_8149,N_7981,N_7989);
nand U8150 (N_8150,N_7884,N_7941);
xor U8151 (N_8151,N_7882,N_7863);
xor U8152 (N_8152,N_7864,N_7882);
or U8153 (N_8153,N_7876,N_7954);
nand U8154 (N_8154,N_7900,N_7878);
nor U8155 (N_8155,N_7923,N_7910);
xnor U8156 (N_8156,N_7968,N_7885);
and U8157 (N_8157,N_7945,N_7990);
nor U8158 (N_8158,N_7993,N_7804);
or U8159 (N_8159,N_7974,N_7837);
xnor U8160 (N_8160,N_7913,N_7918);
xor U8161 (N_8161,N_7801,N_7969);
and U8162 (N_8162,N_7812,N_7919);
nor U8163 (N_8163,N_7829,N_7865);
nor U8164 (N_8164,N_7991,N_7850);
xnor U8165 (N_8165,N_7912,N_7956);
nand U8166 (N_8166,N_7815,N_7809);
or U8167 (N_8167,N_7810,N_7952);
nor U8168 (N_8168,N_7934,N_7829);
nor U8169 (N_8169,N_7849,N_7839);
nor U8170 (N_8170,N_7830,N_7823);
and U8171 (N_8171,N_7977,N_7893);
nand U8172 (N_8172,N_7980,N_7897);
and U8173 (N_8173,N_7877,N_7895);
and U8174 (N_8174,N_7875,N_7975);
nor U8175 (N_8175,N_7867,N_7929);
or U8176 (N_8176,N_7942,N_7974);
nor U8177 (N_8177,N_7819,N_7878);
xor U8178 (N_8178,N_7868,N_7986);
and U8179 (N_8179,N_7890,N_7900);
nor U8180 (N_8180,N_7944,N_7863);
xnor U8181 (N_8181,N_7830,N_7851);
or U8182 (N_8182,N_7834,N_7988);
xor U8183 (N_8183,N_7984,N_7859);
nand U8184 (N_8184,N_7954,N_7923);
and U8185 (N_8185,N_7879,N_7914);
and U8186 (N_8186,N_7893,N_7824);
nor U8187 (N_8187,N_7978,N_7943);
xor U8188 (N_8188,N_7997,N_7925);
or U8189 (N_8189,N_7828,N_7947);
xor U8190 (N_8190,N_7822,N_7913);
nand U8191 (N_8191,N_7994,N_7963);
nor U8192 (N_8192,N_7963,N_7991);
nand U8193 (N_8193,N_7900,N_7948);
xor U8194 (N_8194,N_7902,N_7825);
or U8195 (N_8195,N_7811,N_7908);
nor U8196 (N_8196,N_7955,N_7841);
or U8197 (N_8197,N_7816,N_7931);
xor U8198 (N_8198,N_7816,N_7823);
and U8199 (N_8199,N_7949,N_7820);
or U8200 (N_8200,N_8197,N_8112);
nand U8201 (N_8201,N_8135,N_8131);
or U8202 (N_8202,N_8132,N_8175);
xnor U8203 (N_8203,N_8183,N_8091);
nand U8204 (N_8204,N_8076,N_8096);
or U8205 (N_8205,N_8128,N_8032);
xnor U8206 (N_8206,N_8066,N_8017);
nor U8207 (N_8207,N_8038,N_8015);
or U8208 (N_8208,N_8051,N_8063);
nor U8209 (N_8209,N_8044,N_8125);
and U8210 (N_8210,N_8192,N_8115);
xor U8211 (N_8211,N_8190,N_8193);
nor U8212 (N_8212,N_8155,N_8013);
or U8213 (N_8213,N_8179,N_8176);
nor U8214 (N_8214,N_8011,N_8100);
and U8215 (N_8215,N_8198,N_8158);
nand U8216 (N_8216,N_8094,N_8110);
or U8217 (N_8217,N_8064,N_8180);
nand U8218 (N_8218,N_8120,N_8058);
nand U8219 (N_8219,N_8178,N_8170);
nor U8220 (N_8220,N_8107,N_8068);
or U8221 (N_8221,N_8195,N_8097);
and U8222 (N_8222,N_8102,N_8114);
or U8223 (N_8223,N_8134,N_8137);
or U8224 (N_8224,N_8073,N_8159);
xnor U8225 (N_8225,N_8016,N_8008);
nor U8226 (N_8226,N_8023,N_8113);
xnor U8227 (N_8227,N_8109,N_8092);
nor U8228 (N_8228,N_8024,N_8182);
xnor U8229 (N_8229,N_8117,N_8030);
nor U8230 (N_8230,N_8150,N_8065);
nor U8231 (N_8231,N_8174,N_8034);
or U8232 (N_8232,N_8162,N_8140);
and U8233 (N_8233,N_8136,N_8143);
and U8234 (N_8234,N_8083,N_8001);
xnor U8235 (N_8235,N_8042,N_8028);
and U8236 (N_8236,N_8098,N_8168);
or U8237 (N_8237,N_8111,N_8090);
xnor U8238 (N_8238,N_8037,N_8084);
and U8239 (N_8239,N_8133,N_8152);
or U8240 (N_8240,N_8149,N_8104);
or U8241 (N_8241,N_8087,N_8022);
xnor U8242 (N_8242,N_8021,N_8148);
and U8243 (N_8243,N_8039,N_8194);
or U8244 (N_8244,N_8025,N_8081);
xnor U8245 (N_8245,N_8167,N_8086);
nand U8246 (N_8246,N_8046,N_8103);
nand U8247 (N_8247,N_8181,N_8018);
or U8248 (N_8248,N_8072,N_8164);
nand U8249 (N_8249,N_8138,N_8186);
nor U8250 (N_8250,N_8123,N_8003);
nor U8251 (N_8251,N_8053,N_8043);
or U8252 (N_8252,N_8082,N_8040);
nor U8253 (N_8253,N_8020,N_8071);
nor U8254 (N_8254,N_8169,N_8002);
nor U8255 (N_8255,N_8163,N_8057);
nand U8256 (N_8256,N_8031,N_8077);
nand U8257 (N_8257,N_8118,N_8041);
and U8258 (N_8258,N_8060,N_8045);
nand U8259 (N_8259,N_8156,N_8172);
nand U8260 (N_8260,N_8165,N_8056);
or U8261 (N_8261,N_8079,N_8101);
and U8262 (N_8262,N_8035,N_8067);
nor U8263 (N_8263,N_8062,N_8173);
nand U8264 (N_8264,N_8145,N_8089);
or U8265 (N_8265,N_8129,N_8055);
or U8266 (N_8266,N_8151,N_8099);
and U8267 (N_8267,N_8093,N_8187);
nand U8268 (N_8268,N_8106,N_8061);
nor U8269 (N_8269,N_8124,N_8177);
and U8270 (N_8270,N_8116,N_8007);
nand U8271 (N_8271,N_8027,N_8160);
nand U8272 (N_8272,N_8070,N_8154);
nor U8273 (N_8273,N_8119,N_8142);
and U8274 (N_8274,N_8019,N_8012);
xnor U8275 (N_8275,N_8157,N_8185);
nand U8276 (N_8276,N_8188,N_8147);
and U8277 (N_8277,N_8080,N_8054);
nor U8278 (N_8278,N_8052,N_8000);
nand U8279 (N_8279,N_8139,N_8075);
nand U8280 (N_8280,N_8004,N_8122);
or U8281 (N_8281,N_8171,N_8085);
or U8282 (N_8282,N_8078,N_8161);
xnor U8283 (N_8283,N_8026,N_8184);
or U8284 (N_8284,N_8009,N_8130);
and U8285 (N_8285,N_8049,N_8189);
and U8286 (N_8286,N_8059,N_8141);
and U8287 (N_8287,N_8014,N_8095);
nor U8288 (N_8288,N_8048,N_8006);
xnor U8289 (N_8289,N_8010,N_8144);
xor U8290 (N_8290,N_8069,N_8036);
xor U8291 (N_8291,N_8121,N_8047);
nor U8292 (N_8292,N_8196,N_8005);
nand U8293 (N_8293,N_8126,N_8146);
xor U8294 (N_8294,N_8029,N_8033);
nor U8295 (N_8295,N_8199,N_8108);
or U8296 (N_8296,N_8191,N_8127);
nand U8297 (N_8297,N_8050,N_8105);
or U8298 (N_8298,N_8088,N_8166);
or U8299 (N_8299,N_8153,N_8074);
xnor U8300 (N_8300,N_8060,N_8135);
xnor U8301 (N_8301,N_8184,N_8115);
nand U8302 (N_8302,N_8174,N_8056);
or U8303 (N_8303,N_8175,N_8052);
xnor U8304 (N_8304,N_8047,N_8022);
nand U8305 (N_8305,N_8141,N_8043);
xor U8306 (N_8306,N_8197,N_8099);
or U8307 (N_8307,N_8044,N_8056);
or U8308 (N_8308,N_8068,N_8039);
and U8309 (N_8309,N_8130,N_8146);
nand U8310 (N_8310,N_8066,N_8129);
nand U8311 (N_8311,N_8109,N_8026);
nor U8312 (N_8312,N_8061,N_8099);
nand U8313 (N_8313,N_8098,N_8036);
or U8314 (N_8314,N_8081,N_8179);
nand U8315 (N_8315,N_8196,N_8020);
nor U8316 (N_8316,N_8125,N_8048);
nor U8317 (N_8317,N_8132,N_8074);
nor U8318 (N_8318,N_8138,N_8017);
xor U8319 (N_8319,N_8188,N_8198);
nor U8320 (N_8320,N_8037,N_8000);
or U8321 (N_8321,N_8029,N_8196);
nor U8322 (N_8322,N_8182,N_8065);
xor U8323 (N_8323,N_8191,N_8120);
xor U8324 (N_8324,N_8133,N_8078);
xnor U8325 (N_8325,N_8199,N_8000);
nor U8326 (N_8326,N_8078,N_8131);
and U8327 (N_8327,N_8135,N_8191);
nor U8328 (N_8328,N_8129,N_8054);
nand U8329 (N_8329,N_8180,N_8110);
xnor U8330 (N_8330,N_8103,N_8064);
nor U8331 (N_8331,N_8160,N_8057);
xnor U8332 (N_8332,N_8187,N_8141);
or U8333 (N_8333,N_8077,N_8041);
and U8334 (N_8334,N_8165,N_8101);
nor U8335 (N_8335,N_8069,N_8173);
nand U8336 (N_8336,N_8087,N_8008);
and U8337 (N_8337,N_8129,N_8125);
or U8338 (N_8338,N_8183,N_8064);
nor U8339 (N_8339,N_8128,N_8113);
or U8340 (N_8340,N_8016,N_8023);
nand U8341 (N_8341,N_8192,N_8152);
nand U8342 (N_8342,N_8074,N_8046);
or U8343 (N_8343,N_8007,N_8096);
or U8344 (N_8344,N_8157,N_8189);
nand U8345 (N_8345,N_8046,N_8163);
nand U8346 (N_8346,N_8112,N_8110);
xor U8347 (N_8347,N_8195,N_8052);
and U8348 (N_8348,N_8099,N_8062);
xor U8349 (N_8349,N_8048,N_8152);
or U8350 (N_8350,N_8084,N_8111);
xnor U8351 (N_8351,N_8021,N_8059);
or U8352 (N_8352,N_8016,N_8180);
nand U8353 (N_8353,N_8117,N_8020);
and U8354 (N_8354,N_8030,N_8033);
nor U8355 (N_8355,N_8053,N_8067);
xnor U8356 (N_8356,N_8139,N_8154);
nand U8357 (N_8357,N_8156,N_8013);
or U8358 (N_8358,N_8119,N_8192);
and U8359 (N_8359,N_8086,N_8079);
and U8360 (N_8360,N_8101,N_8013);
xnor U8361 (N_8361,N_8078,N_8166);
nand U8362 (N_8362,N_8021,N_8117);
nand U8363 (N_8363,N_8044,N_8062);
and U8364 (N_8364,N_8084,N_8152);
nand U8365 (N_8365,N_8101,N_8034);
nor U8366 (N_8366,N_8071,N_8104);
xnor U8367 (N_8367,N_8188,N_8031);
and U8368 (N_8368,N_8177,N_8180);
xnor U8369 (N_8369,N_8051,N_8028);
nand U8370 (N_8370,N_8007,N_8155);
nor U8371 (N_8371,N_8111,N_8182);
or U8372 (N_8372,N_8160,N_8118);
nand U8373 (N_8373,N_8132,N_8006);
nor U8374 (N_8374,N_8035,N_8045);
nor U8375 (N_8375,N_8179,N_8048);
and U8376 (N_8376,N_8115,N_8187);
nor U8377 (N_8377,N_8101,N_8046);
nor U8378 (N_8378,N_8093,N_8047);
or U8379 (N_8379,N_8156,N_8139);
nor U8380 (N_8380,N_8187,N_8053);
and U8381 (N_8381,N_8197,N_8080);
nor U8382 (N_8382,N_8024,N_8003);
or U8383 (N_8383,N_8146,N_8184);
and U8384 (N_8384,N_8133,N_8020);
nor U8385 (N_8385,N_8160,N_8162);
nor U8386 (N_8386,N_8133,N_8155);
nor U8387 (N_8387,N_8097,N_8019);
nand U8388 (N_8388,N_8120,N_8060);
and U8389 (N_8389,N_8067,N_8080);
or U8390 (N_8390,N_8133,N_8007);
xnor U8391 (N_8391,N_8034,N_8112);
and U8392 (N_8392,N_8136,N_8184);
and U8393 (N_8393,N_8125,N_8045);
nand U8394 (N_8394,N_8027,N_8050);
xnor U8395 (N_8395,N_8181,N_8005);
nor U8396 (N_8396,N_8006,N_8053);
nand U8397 (N_8397,N_8087,N_8029);
xnor U8398 (N_8398,N_8111,N_8055);
nor U8399 (N_8399,N_8148,N_8083);
nor U8400 (N_8400,N_8331,N_8391);
and U8401 (N_8401,N_8269,N_8325);
nor U8402 (N_8402,N_8213,N_8254);
xor U8403 (N_8403,N_8312,N_8366);
and U8404 (N_8404,N_8282,N_8291);
and U8405 (N_8405,N_8201,N_8262);
nor U8406 (N_8406,N_8316,N_8354);
and U8407 (N_8407,N_8294,N_8383);
and U8408 (N_8408,N_8328,N_8252);
or U8409 (N_8409,N_8271,N_8364);
nand U8410 (N_8410,N_8244,N_8327);
or U8411 (N_8411,N_8289,N_8314);
and U8412 (N_8412,N_8394,N_8200);
nand U8413 (N_8413,N_8335,N_8317);
nand U8414 (N_8414,N_8227,N_8236);
and U8415 (N_8415,N_8398,N_8225);
nor U8416 (N_8416,N_8384,N_8353);
xor U8417 (N_8417,N_8358,N_8237);
nand U8418 (N_8418,N_8250,N_8303);
nand U8419 (N_8419,N_8382,N_8318);
and U8420 (N_8420,N_8336,N_8320);
xnor U8421 (N_8421,N_8390,N_8330);
nor U8422 (N_8422,N_8315,N_8329);
and U8423 (N_8423,N_8243,N_8239);
nand U8424 (N_8424,N_8210,N_8334);
or U8425 (N_8425,N_8286,N_8298);
nand U8426 (N_8426,N_8324,N_8321);
and U8427 (N_8427,N_8229,N_8277);
nand U8428 (N_8428,N_8204,N_8295);
xor U8429 (N_8429,N_8265,N_8309);
or U8430 (N_8430,N_8385,N_8326);
or U8431 (N_8431,N_8238,N_8249);
or U8432 (N_8432,N_8297,N_8278);
and U8433 (N_8433,N_8258,N_8226);
and U8434 (N_8434,N_8395,N_8344);
nand U8435 (N_8435,N_8389,N_8284);
xor U8436 (N_8436,N_8206,N_8251);
nor U8437 (N_8437,N_8220,N_8281);
or U8438 (N_8438,N_8323,N_8274);
nor U8439 (N_8439,N_8349,N_8346);
nor U8440 (N_8440,N_8362,N_8370);
xor U8441 (N_8441,N_8203,N_8386);
nand U8442 (N_8442,N_8228,N_8372);
nand U8443 (N_8443,N_8290,N_8368);
nand U8444 (N_8444,N_8319,N_8221);
xor U8445 (N_8445,N_8342,N_8369);
nand U8446 (N_8446,N_8339,N_8270);
nor U8447 (N_8447,N_8300,N_8245);
nor U8448 (N_8448,N_8343,N_8365);
and U8449 (N_8449,N_8264,N_8256);
or U8450 (N_8450,N_8241,N_8235);
nor U8451 (N_8451,N_8363,N_8311);
and U8452 (N_8452,N_8257,N_8380);
or U8453 (N_8453,N_8373,N_8287);
nor U8454 (N_8454,N_8340,N_8224);
or U8455 (N_8455,N_8367,N_8378);
nor U8456 (N_8456,N_8234,N_8253);
nor U8457 (N_8457,N_8355,N_8360);
nand U8458 (N_8458,N_8299,N_8379);
nor U8459 (N_8459,N_8218,N_8397);
and U8460 (N_8460,N_8233,N_8399);
nand U8461 (N_8461,N_8306,N_8375);
xor U8462 (N_8462,N_8308,N_8293);
or U8463 (N_8463,N_8248,N_8280);
nor U8464 (N_8464,N_8279,N_8333);
or U8465 (N_8465,N_8381,N_8301);
xor U8466 (N_8466,N_8232,N_8352);
and U8467 (N_8467,N_8223,N_8214);
nand U8468 (N_8468,N_8307,N_8338);
or U8469 (N_8469,N_8255,N_8351);
xor U8470 (N_8470,N_8357,N_8212);
and U8471 (N_8471,N_8275,N_8350);
nand U8472 (N_8472,N_8261,N_8377);
or U8473 (N_8473,N_8292,N_8374);
xor U8474 (N_8474,N_8208,N_8231);
nor U8475 (N_8475,N_8209,N_8216);
and U8476 (N_8476,N_8361,N_8273);
nand U8477 (N_8477,N_8205,N_8242);
or U8478 (N_8478,N_8387,N_8345);
and U8479 (N_8479,N_8288,N_8359);
or U8480 (N_8480,N_8240,N_8313);
nand U8481 (N_8481,N_8371,N_8393);
nor U8482 (N_8482,N_8230,N_8259);
and U8483 (N_8483,N_8348,N_8272);
and U8484 (N_8484,N_8332,N_8388);
or U8485 (N_8485,N_8347,N_8267);
or U8486 (N_8486,N_8296,N_8211);
and U8487 (N_8487,N_8246,N_8302);
and U8488 (N_8488,N_8376,N_8322);
xnor U8489 (N_8489,N_8276,N_8207);
xnor U8490 (N_8490,N_8283,N_8341);
nand U8491 (N_8491,N_8217,N_8285);
xnor U8492 (N_8492,N_8337,N_8305);
and U8493 (N_8493,N_8268,N_8310);
xnor U8494 (N_8494,N_8202,N_8247);
and U8495 (N_8495,N_8219,N_8215);
nor U8496 (N_8496,N_8260,N_8356);
or U8497 (N_8497,N_8396,N_8266);
and U8498 (N_8498,N_8304,N_8392);
or U8499 (N_8499,N_8222,N_8263);
nor U8500 (N_8500,N_8274,N_8228);
nor U8501 (N_8501,N_8347,N_8262);
and U8502 (N_8502,N_8230,N_8361);
nand U8503 (N_8503,N_8243,N_8348);
xor U8504 (N_8504,N_8397,N_8314);
or U8505 (N_8505,N_8317,N_8242);
and U8506 (N_8506,N_8260,N_8337);
nor U8507 (N_8507,N_8295,N_8395);
and U8508 (N_8508,N_8276,N_8264);
nor U8509 (N_8509,N_8398,N_8312);
or U8510 (N_8510,N_8247,N_8372);
xnor U8511 (N_8511,N_8368,N_8332);
nor U8512 (N_8512,N_8207,N_8353);
nor U8513 (N_8513,N_8282,N_8326);
or U8514 (N_8514,N_8255,N_8222);
and U8515 (N_8515,N_8323,N_8266);
nor U8516 (N_8516,N_8219,N_8293);
xnor U8517 (N_8517,N_8211,N_8311);
nor U8518 (N_8518,N_8371,N_8399);
nor U8519 (N_8519,N_8256,N_8351);
xor U8520 (N_8520,N_8221,N_8365);
nand U8521 (N_8521,N_8335,N_8322);
nand U8522 (N_8522,N_8337,N_8277);
or U8523 (N_8523,N_8205,N_8351);
nand U8524 (N_8524,N_8219,N_8247);
xor U8525 (N_8525,N_8325,N_8225);
nor U8526 (N_8526,N_8206,N_8361);
and U8527 (N_8527,N_8353,N_8222);
xor U8528 (N_8528,N_8340,N_8217);
or U8529 (N_8529,N_8219,N_8303);
and U8530 (N_8530,N_8302,N_8341);
xnor U8531 (N_8531,N_8222,N_8366);
and U8532 (N_8532,N_8310,N_8351);
nor U8533 (N_8533,N_8278,N_8202);
nor U8534 (N_8534,N_8304,N_8346);
nand U8535 (N_8535,N_8247,N_8255);
nor U8536 (N_8536,N_8354,N_8287);
or U8537 (N_8537,N_8242,N_8392);
nor U8538 (N_8538,N_8286,N_8235);
or U8539 (N_8539,N_8349,N_8335);
xor U8540 (N_8540,N_8344,N_8323);
nor U8541 (N_8541,N_8342,N_8219);
and U8542 (N_8542,N_8255,N_8362);
nor U8543 (N_8543,N_8274,N_8343);
xnor U8544 (N_8544,N_8353,N_8395);
xor U8545 (N_8545,N_8367,N_8216);
and U8546 (N_8546,N_8386,N_8263);
and U8547 (N_8547,N_8255,N_8288);
xnor U8548 (N_8548,N_8263,N_8373);
and U8549 (N_8549,N_8354,N_8368);
xor U8550 (N_8550,N_8302,N_8276);
and U8551 (N_8551,N_8264,N_8331);
or U8552 (N_8552,N_8294,N_8321);
or U8553 (N_8553,N_8240,N_8281);
nand U8554 (N_8554,N_8345,N_8248);
nand U8555 (N_8555,N_8294,N_8274);
nor U8556 (N_8556,N_8328,N_8361);
nor U8557 (N_8557,N_8386,N_8255);
or U8558 (N_8558,N_8210,N_8363);
or U8559 (N_8559,N_8326,N_8210);
or U8560 (N_8560,N_8340,N_8216);
or U8561 (N_8561,N_8334,N_8312);
xor U8562 (N_8562,N_8211,N_8275);
and U8563 (N_8563,N_8361,N_8324);
nor U8564 (N_8564,N_8381,N_8310);
and U8565 (N_8565,N_8275,N_8376);
nor U8566 (N_8566,N_8301,N_8306);
and U8567 (N_8567,N_8318,N_8364);
and U8568 (N_8568,N_8268,N_8389);
and U8569 (N_8569,N_8202,N_8312);
nand U8570 (N_8570,N_8313,N_8383);
xnor U8571 (N_8571,N_8388,N_8289);
or U8572 (N_8572,N_8212,N_8368);
nand U8573 (N_8573,N_8304,N_8237);
nand U8574 (N_8574,N_8309,N_8389);
and U8575 (N_8575,N_8331,N_8355);
nor U8576 (N_8576,N_8285,N_8355);
xor U8577 (N_8577,N_8331,N_8203);
nor U8578 (N_8578,N_8348,N_8264);
xnor U8579 (N_8579,N_8201,N_8360);
xor U8580 (N_8580,N_8307,N_8213);
and U8581 (N_8581,N_8255,N_8398);
and U8582 (N_8582,N_8321,N_8277);
or U8583 (N_8583,N_8236,N_8336);
or U8584 (N_8584,N_8337,N_8358);
and U8585 (N_8585,N_8324,N_8314);
and U8586 (N_8586,N_8225,N_8222);
and U8587 (N_8587,N_8240,N_8389);
xnor U8588 (N_8588,N_8274,N_8223);
or U8589 (N_8589,N_8261,N_8200);
and U8590 (N_8590,N_8263,N_8220);
nor U8591 (N_8591,N_8396,N_8285);
nand U8592 (N_8592,N_8260,N_8201);
nor U8593 (N_8593,N_8362,N_8394);
and U8594 (N_8594,N_8209,N_8239);
or U8595 (N_8595,N_8207,N_8360);
and U8596 (N_8596,N_8342,N_8399);
and U8597 (N_8597,N_8338,N_8332);
nand U8598 (N_8598,N_8380,N_8322);
nor U8599 (N_8599,N_8238,N_8301);
nand U8600 (N_8600,N_8470,N_8430);
or U8601 (N_8601,N_8561,N_8433);
nor U8602 (N_8602,N_8511,N_8528);
or U8603 (N_8603,N_8480,N_8440);
or U8604 (N_8604,N_8596,N_8504);
or U8605 (N_8605,N_8478,N_8424);
and U8606 (N_8606,N_8557,N_8565);
and U8607 (N_8607,N_8505,N_8562);
or U8608 (N_8608,N_8442,N_8556);
nor U8609 (N_8609,N_8537,N_8581);
nand U8610 (N_8610,N_8541,N_8506);
or U8611 (N_8611,N_8590,N_8498);
or U8612 (N_8612,N_8490,N_8444);
and U8613 (N_8613,N_8499,N_8534);
nand U8614 (N_8614,N_8507,N_8571);
or U8615 (N_8615,N_8420,N_8486);
or U8616 (N_8616,N_8594,N_8418);
and U8617 (N_8617,N_8475,N_8543);
nand U8618 (N_8618,N_8595,N_8449);
and U8619 (N_8619,N_8404,N_8587);
and U8620 (N_8620,N_8495,N_8539);
nor U8621 (N_8621,N_8593,N_8538);
and U8622 (N_8622,N_8567,N_8456);
nand U8623 (N_8623,N_8542,N_8533);
and U8624 (N_8624,N_8431,N_8483);
xor U8625 (N_8625,N_8484,N_8407);
and U8626 (N_8626,N_8471,N_8578);
nor U8627 (N_8627,N_8513,N_8580);
nand U8628 (N_8628,N_8474,N_8441);
and U8629 (N_8629,N_8568,N_8510);
and U8630 (N_8630,N_8428,N_8454);
nand U8631 (N_8631,N_8517,N_8588);
or U8632 (N_8632,N_8438,N_8447);
and U8633 (N_8633,N_8419,N_8555);
xnor U8634 (N_8634,N_8560,N_8577);
or U8635 (N_8635,N_8405,N_8477);
nor U8636 (N_8636,N_8481,N_8563);
nand U8637 (N_8637,N_8417,N_8497);
nor U8638 (N_8638,N_8421,N_8451);
nand U8639 (N_8639,N_8525,N_8466);
or U8640 (N_8640,N_8552,N_8502);
nand U8641 (N_8641,N_8529,N_8408);
nor U8642 (N_8642,N_8452,N_8515);
or U8643 (N_8643,N_8463,N_8423);
nand U8644 (N_8644,N_8462,N_8592);
nor U8645 (N_8645,N_8485,N_8548);
or U8646 (N_8646,N_8482,N_8461);
nand U8647 (N_8647,N_8446,N_8468);
nor U8648 (N_8648,N_8429,N_8514);
nor U8649 (N_8649,N_8576,N_8455);
and U8650 (N_8650,N_8526,N_8439);
nor U8651 (N_8651,N_8489,N_8573);
and U8652 (N_8652,N_8472,N_8450);
xnor U8653 (N_8653,N_8564,N_8467);
and U8654 (N_8654,N_8530,N_8547);
or U8655 (N_8655,N_8518,N_8558);
nor U8656 (N_8656,N_8569,N_8512);
and U8657 (N_8657,N_8412,N_8524);
and U8658 (N_8658,N_8527,N_8414);
or U8659 (N_8659,N_8535,N_8584);
xor U8660 (N_8660,N_8453,N_8591);
or U8661 (N_8661,N_8436,N_8536);
or U8662 (N_8662,N_8491,N_8473);
nor U8663 (N_8663,N_8501,N_8425);
nand U8664 (N_8664,N_8476,N_8409);
and U8665 (N_8665,N_8597,N_8574);
and U8666 (N_8666,N_8410,N_8411);
nand U8667 (N_8667,N_8540,N_8523);
nor U8668 (N_8668,N_8458,N_8583);
xnor U8669 (N_8669,N_8457,N_8549);
or U8670 (N_8670,N_8402,N_8599);
xnor U8671 (N_8671,N_8532,N_8500);
and U8672 (N_8672,N_8516,N_8544);
or U8673 (N_8673,N_8546,N_8437);
or U8674 (N_8674,N_8508,N_8415);
xor U8675 (N_8675,N_8403,N_8521);
and U8676 (N_8676,N_8492,N_8509);
xor U8677 (N_8677,N_8531,N_8487);
or U8678 (N_8678,N_8503,N_8579);
and U8679 (N_8679,N_8493,N_8427);
xnor U8680 (N_8680,N_8426,N_8422);
nor U8681 (N_8681,N_8464,N_8416);
and U8682 (N_8682,N_8589,N_8519);
nand U8683 (N_8683,N_8460,N_8432);
nand U8684 (N_8684,N_8570,N_8494);
or U8685 (N_8685,N_8553,N_8496);
nand U8686 (N_8686,N_8448,N_8443);
and U8687 (N_8687,N_8401,N_8445);
nor U8688 (N_8688,N_8520,N_8434);
or U8689 (N_8689,N_8465,N_8559);
xor U8690 (N_8690,N_8598,N_8585);
or U8691 (N_8691,N_8406,N_8413);
xor U8692 (N_8692,N_8575,N_8545);
or U8693 (N_8693,N_8551,N_8566);
and U8694 (N_8694,N_8400,N_8586);
nor U8695 (N_8695,N_8550,N_8469);
and U8696 (N_8696,N_8459,N_8554);
xnor U8697 (N_8697,N_8435,N_8572);
or U8698 (N_8698,N_8522,N_8582);
and U8699 (N_8699,N_8479,N_8488);
nor U8700 (N_8700,N_8573,N_8484);
or U8701 (N_8701,N_8576,N_8535);
xnor U8702 (N_8702,N_8443,N_8465);
and U8703 (N_8703,N_8589,N_8403);
or U8704 (N_8704,N_8580,N_8543);
and U8705 (N_8705,N_8503,N_8594);
nand U8706 (N_8706,N_8561,N_8484);
and U8707 (N_8707,N_8550,N_8562);
nor U8708 (N_8708,N_8599,N_8557);
and U8709 (N_8709,N_8483,N_8561);
or U8710 (N_8710,N_8439,N_8400);
and U8711 (N_8711,N_8496,N_8415);
or U8712 (N_8712,N_8597,N_8404);
nor U8713 (N_8713,N_8469,N_8586);
nor U8714 (N_8714,N_8591,N_8444);
nand U8715 (N_8715,N_8419,N_8537);
or U8716 (N_8716,N_8410,N_8487);
nor U8717 (N_8717,N_8566,N_8511);
or U8718 (N_8718,N_8478,N_8555);
nor U8719 (N_8719,N_8538,N_8434);
xnor U8720 (N_8720,N_8403,N_8576);
nor U8721 (N_8721,N_8433,N_8485);
xor U8722 (N_8722,N_8578,N_8476);
xor U8723 (N_8723,N_8448,N_8455);
xor U8724 (N_8724,N_8405,N_8509);
nor U8725 (N_8725,N_8478,N_8519);
nand U8726 (N_8726,N_8430,N_8547);
or U8727 (N_8727,N_8411,N_8466);
xor U8728 (N_8728,N_8497,N_8588);
or U8729 (N_8729,N_8560,N_8452);
nor U8730 (N_8730,N_8456,N_8480);
and U8731 (N_8731,N_8413,N_8553);
or U8732 (N_8732,N_8416,N_8420);
nand U8733 (N_8733,N_8491,N_8520);
and U8734 (N_8734,N_8460,N_8478);
or U8735 (N_8735,N_8537,N_8480);
nand U8736 (N_8736,N_8568,N_8592);
xnor U8737 (N_8737,N_8475,N_8420);
nand U8738 (N_8738,N_8404,N_8457);
nand U8739 (N_8739,N_8407,N_8427);
and U8740 (N_8740,N_8566,N_8403);
and U8741 (N_8741,N_8555,N_8584);
and U8742 (N_8742,N_8550,N_8592);
and U8743 (N_8743,N_8594,N_8448);
nor U8744 (N_8744,N_8434,N_8506);
nor U8745 (N_8745,N_8491,N_8421);
nor U8746 (N_8746,N_8486,N_8591);
nand U8747 (N_8747,N_8594,N_8515);
nand U8748 (N_8748,N_8494,N_8475);
nor U8749 (N_8749,N_8492,N_8409);
nand U8750 (N_8750,N_8438,N_8546);
and U8751 (N_8751,N_8584,N_8541);
or U8752 (N_8752,N_8594,N_8552);
and U8753 (N_8753,N_8407,N_8447);
xnor U8754 (N_8754,N_8550,N_8489);
nor U8755 (N_8755,N_8533,N_8517);
nor U8756 (N_8756,N_8595,N_8567);
or U8757 (N_8757,N_8466,N_8533);
nor U8758 (N_8758,N_8555,N_8510);
nor U8759 (N_8759,N_8441,N_8581);
and U8760 (N_8760,N_8424,N_8499);
and U8761 (N_8761,N_8454,N_8481);
nand U8762 (N_8762,N_8589,N_8442);
or U8763 (N_8763,N_8597,N_8417);
xor U8764 (N_8764,N_8565,N_8455);
and U8765 (N_8765,N_8429,N_8495);
xnor U8766 (N_8766,N_8457,N_8471);
or U8767 (N_8767,N_8598,N_8593);
and U8768 (N_8768,N_8561,N_8479);
xnor U8769 (N_8769,N_8453,N_8409);
or U8770 (N_8770,N_8572,N_8404);
xor U8771 (N_8771,N_8417,N_8409);
and U8772 (N_8772,N_8491,N_8547);
xor U8773 (N_8773,N_8518,N_8519);
or U8774 (N_8774,N_8532,N_8587);
nor U8775 (N_8775,N_8497,N_8473);
nand U8776 (N_8776,N_8522,N_8413);
xor U8777 (N_8777,N_8555,N_8420);
xor U8778 (N_8778,N_8556,N_8541);
or U8779 (N_8779,N_8555,N_8561);
nor U8780 (N_8780,N_8477,N_8559);
or U8781 (N_8781,N_8422,N_8455);
nor U8782 (N_8782,N_8446,N_8439);
and U8783 (N_8783,N_8559,N_8515);
nand U8784 (N_8784,N_8586,N_8440);
nor U8785 (N_8785,N_8488,N_8481);
nor U8786 (N_8786,N_8464,N_8518);
or U8787 (N_8787,N_8486,N_8595);
nand U8788 (N_8788,N_8572,N_8538);
and U8789 (N_8789,N_8439,N_8459);
or U8790 (N_8790,N_8532,N_8525);
xor U8791 (N_8791,N_8526,N_8515);
or U8792 (N_8792,N_8408,N_8468);
or U8793 (N_8793,N_8466,N_8517);
and U8794 (N_8794,N_8597,N_8431);
nand U8795 (N_8795,N_8401,N_8575);
xnor U8796 (N_8796,N_8517,N_8438);
nor U8797 (N_8797,N_8451,N_8450);
and U8798 (N_8798,N_8425,N_8468);
nor U8799 (N_8799,N_8556,N_8450);
xnor U8800 (N_8800,N_8714,N_8618);
or U8801 (N_8801,N_8743,N_8752);
nand U8802 (N_8802,N_8732,N_8796);
xor U8803 (N_8803,N_8734,N_8682);
nor U8804 (N_8804,N_8718,N_8730);
nor U8805 (N_8805,N_8620,N_8698);
nor U8806 (N_8806,N_8601,N_8612);
or U8807 (N_8807,N_8735,N_8717);
or U8808 (N_8808,N_8750,N_8627);
or U8809 (N_8809,N_8753,N_8629);
xor U8810 (N_8810,N_8652,N_8688);
or U8811 (N_8811,N_8793,N_8617);
xor U8812 (N_8812,N_8733,N_8690);
and U8813 (N_8813,N_8628,N_8630);
or U8814 (N_8814,N_8740,N_8788);
nand U8815 (N_8815,N_8692,N_8670);
or U8816 (N_8816,N_8705,N_8797);
nand U8817 (N_8817,N_8710,N_8660);
nand U8818 (N_8818,N_8722,N_8765);
xnor U8819 (N_8819,N_8696,N_8699);
or U8820 (N_8820,N_8642,N_8745);
nor U8821 (N_8821,N_8623,N_8742);
nor U8822 (N_8822,N_8639,N_8654);
nor U8823 (N_8823,N_8604,N_8686);
or U8824 (N_8824,N_8697,N_8731);
and U8825 (N_8825,N_8641,N_8727);
nor U8826 (N_8826,N_8616,N_8606);
and U8827 (N_8827,N_8744,N_8781);
nor U8828 (N_8828,N_8792,N_8636);
and U8829 (N_8829,N_8761,N_8737);
xnor U8830 (N_8830,N_8725,N_8706);
nand U8831 (N_8831,N_8785,N_8665);
and U8832 (N_8832,N_8762,N_8709);
nand U8833 (N_8833,N_8695,N_8694);
xnor U8834 (N_8834,N_8779,N_8608);
nor U8835 (N_8835,N_8666,N_8702);
and U8836 (N_8836,N_8640,N_8783);
and U8837 (N_8837,N_8789,N_8647);
nor U8838 (N_8838,N_8767,N_8751);
nor U8839 (N_8839,N_8650,N_8776);
nand U8840 (N_8840,N_8600,N_8659);
nor U8841 (N_8841,N_8687,N_8609);
or U8842 (N_8842,N_8724,N_8790);
or U8843 (N_8843,N_8635,N_8798);
nand U8844 (N_8844,N_8782,N_8712);
and U8845 (N_8845,N_8678,N_8703);
or U8846 (N_8846,N_8748,N_8738);
and U8847 (N_8847,N_8631,N_8757);
xnor U8848 (N_8848,N_8602,N_8637);
or U8849 (N_8849,N_8615,N_8624);
xor U8850 (N_8850,N_8683,N_8746);
xnor U8851 (N_8851,N_8786,N_8739);
or U8852 (N_8852,N_8663,N_8685);
and U8853 (N_8853,N_8708,N_8649);
xor U8854 (N_8854,N_8784,N_8726);
xnor U8855 (N_8855,N_8653,N_8671);
nor U8856 (N_8856,N_8773,N_8775);
nor U8857 (N_8857,N_8626,N_8681);
or U8858 (N_8858,N_8759,N_8684);
nand U8859 (N_8859,N_8655,N_8672);
or U8860 (N_8860,N_8611,N_8704);
nor U8861 (N_8861,N_8673,N_8643);
or U8862 (N_8862,N_8674,N_8677);
and U8863 (N_8863,N_8768,N_8758);
or U8864 (N_8864,N_8664,N_8719);
nand U8865 (N_8865,N_8648,N_8772);
nor U8866 (N_8866,N_8614,N_8770);
xnor U8867 (N_8867,N_8621,N_8676);
and U8868 (N_8868,N_8749,N_8736);
nor U8869 (N_8869,N_8774,N_8713);
or U8870 (N_8870,N_8787,N_8691);
and U8871 (N_8871,N_8632,N_8657);
nor U8872 (N_8872,N_8610,N_8667);
nor U8873 (N_8873,N_8689,N_8754);
nor U8874 (N_8874,N_8680,N_8651);
nor U8875 (N_8875,N_8755,N_8646);
and U8876 (N_8876,N_8668,N_8716);
and U8877 (N_8877,N_8658,N_8720);
and U8878 (N_8878,N_8605,N_8723);
nand U8879 (N_8879,N_8700,N_8645);
or U8880 (N_8880,N_8721,N_8766);
xor U8881 (N_8881,N_8729,N_8633);
nand U8882 (N_8882,N_8661,N_8791);
and U8883 (N_8883,N_8728,N_8662);
or U8884 (N_8884,N_8613,N_8763);
and U8885 (N_8885,N_8669,N_8771);
or U8886 (N_8886,N_8634,N_8675);
xor U8887 (N_8887,N_8656,N_8638);
xor U8888 (N_8888,N_8780,N_8794);
and U8889 (N_8889,N_8619,N_8707);
nor U8890 (N_8890,N_8701,N_8607);
or U8891 (N_8891,N_8644,N_8711);
and U8892 (N_8892,N_8777,N_8693);
and U8893 (N_8893,N_8715,N_8625);
or U8894 (N_8894,N_8679,N_8622);
nor U8895 (N_8895,N_8747,N_8756);
xnor U8896 (N_8896,N_8769,N_8764);
and U8897 (N_8897,N_8795,N_8760);
and U8898 (N_8898,N_8799,N_8741);
or U8899 (N_8899,N_8603,N_8778);
and U8900 (N_8900,N_8629,N_8726);
nor U8901 (N_8901,N_8767,N_8748);
nor U8902 (N_8902,N_8621,N_8764);
xor U8903 (N_8903,N_8727,N_8635);
nor U8904 (N_8904,N_8777,N_8673);
xor U8905 (N_8905,N_8787,N_8660);
xor U8906 (N_8906,N_8744,N_8652);
or U8907 (N_8907,N_8654,N_8647);
nand U8908 (N_8908,N_8714,N_8712);
nor U8909 (N_8909,N_8787,N_8770);
xnor U8910 (N_8910,N_8624,N_8638);
and U8911 (N_8911,N_8736,N_8747);
nor U8912 (N_8912,N_8753,N_8685);
xnor U8913 (N_8913,N_8699,N_8702);
nand U8914 (N_8914,N_8782,N_8676);
xnor U8915 (N_8915,N_8785,N_8716);
nand U8916 (N_8916,N_8761,N_8779);
xor U8917 (N_8917,N_8686,N_8601);
nor U8918 (N_8918,N_8702,N_8747);
xnor U8919 (N_8919,N_8796,N_8795);
xor U8920 (N_8920,N_8777,N_8677);
xor U8921 (N_8921,N_8712,N_8723);
or U8922 (N_8922,N_8620,N_8714);
nand U8923 (N_8923,N_8731,N_8673);
nor U8924 (N_8924,N_8652,N_8766);
nor U8925 (N_8925,N_8694,N_8626);
and U8926 (N_8926,N_8797,N_8703);
nand U8927 (N_8927,N_8786,N_8747);
and U8928 (N_8928,N_8789,N_8788);
nor U8929 (N_8929,N_8732,N_8689);
or U8930 (N_8930,N_8685,N_8679);
nand U8931 (N_8931,N_8799,N_8625);
and U8932 (N_8932,N_8661,N_8756);
nor U8933 (N_8933,N_8659,N_8708);
nand U8934 (N_8934,N_8612,N_8649);
nor U8935 (N_8935,N_8641,N_8773);
and U8936 (N_8936,N_8633,N_8695);
and U8937 (N_8937,N_8758,N_8653);
xor U8938 (N_8938,N_8643,N_8727);
xor U8939 (N_8939,N_8632,N_8763);
nor U8940 (N_8940,N_8728,N_8722);
xor U8941 (N_8941,N_8712,N_8611);
xnor U8942 (N_8942,N_8687,N_8619);
or U8943 (N_8943,N_8676,N_8641);
nor U8944 (N_8944,N_8683,N_8689);
or U8945 (N_8945,N_8759,N_8778);
xnor U8946 (N_8946,N_8613,N_8737);
nor U8947 (N_8947,N_8603,N_8647);
nand U8948 (N_8948,N_8643,N_8732);
or U8949 (N_8949,N_8698,N_8796);
and U8950 (N_8950,N_8685,N_8713);
xor U8951 (N_8951,N_8690,N_8765);
nand U8952 (N_8952,N_8742,N_8727);
or U8953 (N_8953,N_8683,N_8740);
nor U8954 (N_8954,N_8625,N_8731);
nand U8955 (N_8955,N_8777,N_8782);
xor U8956 (N_8956,N_8601,N_8635);
nor U8957 (N_8957,N_8687,N_8757);
nand U8958 (N_8958,N_8613,N_8614);
xnor U8959 (N_8959,N_8602,N_8793);
nor U8960 (N_8960,N_8662,N_8743);
or U8961 (N_8961,N_8750,N_8734);
xnor U8962 (N_8962,N_8617,N_8603);
xor U8963 (N_8963,N_8768,N_8775);
or U8964 (N_8964,N_8615,N_8600);
or U8965 (N_8965,N_8788,N_8647);
or U8966 (N_8966,N_8798,N_8618);
and U8967 (N_8967,N_8692,N_8723);
or U8968 (N_8968,N_8775,N_8654);
nand U8969 (N_8969,N_8776,N_8714);
xnor U8970 (N_8970,N_8705,N_8618);
or U8971 (N_8971,N_8799,N_8716);
nand U8972 (N_8972,N_8788,N_8739);
nor U8973 (N_8973,N_8621,N_8719);
nor U8974 (N_8974,N_8699,N_8771);
nor U8975 (N_8975,N_8741,N_8618);
and U8976 (N_8976,N_8775,N_8727);
or U8977 (N_8977,N_8768,N_8766);
xor U8978 (N_8978,N_8613,N_8709);
nand U8979 (N_8979,N_8651,N_8799);
and U8980 (N_8980,N_8705,N_8694);
and U8981 (N_8981,N_8609,N_8683);
nand U8982 (N_8982,N_8702,N_8642);
xnor U8983 (N_8983,N_8734,N_8641);
nand U8984 (N_8984,N_8703,N_8782);
nand U8985 (N_8985,N_8662,N_8708);
and U8986 (N_8986,N_8626,N_8757);
xor U8987 (N_8987,N_8635,N_8756);
and U8988 (N_8988,N_8700,N_8660);
nand U8989 (N_8989,N_8756,N_8714);
xor U8990 (N_8990,N_8721,N_8786);
xnor U8991 (N_8991,N_8730,N_8650);
nand U8992 (N_8992,N_8754,N_8706);
nand U8993 (N_8993,N_8621,N_8732);
nand U8994 (N_8994,N_8793,N_8761);
nand U8995 (N_8995,N_8638,N_8798);
or U8996 (N_8996,N_8674,N_8681);
and U8997 (N_8997,N_8713,N_8782);
or U8998 (N_8998,N_8727,N_8648);
or U8999 (N_8999,N_8736,N_8710);
nor U9000 (N_9000,N_8946,N_8967);
or U9001 (N_9001,N_8915,N_8923);
nand U9002 (N_9002,N_8969,N_8890);
or U9003 (N_9003,N_8876,N_8879);
nor U9004 (N_9004,N_8857,N_8958);
xor U9005 (N_9005,N_8892,N_8907);
and U9006 (N_9006,N_8964,N_8850);
xor U9007 (N_9007,N_8985,N_8819);
xnor U9008 (N_9008,N_8831,N_8941);
and U9009 (N_9009,N_8904,N_8851);
nor U9010 (N_9010,N_8837,N_8947);
nand U9011 (N_9011,N_8852,N_8838);
nand U9012 (N_9012,N_8827,N_8900);
nor U9013 (N_9013,N_8822,N_8954);
nand U9014 (N_9014,N_8963,N_8942);
nand U9015 (N_9015,N_8883,N_8880);
or U9016 (N_9016,N_8898,N_8856);
nor U9017 (N_9017,N_8965,N_8800);
nor U9018 (N_9018,N_8834,N_8878);
and U9019 (N_9019,N_8829,N_8918);
nor U9020 (N_9020,N_8801,N_8846);
or U9021 (N_9021,N_8867,N_8914);
nand U9022 (N_9022,N_8853,N_8917);
and U9023 (N_9023,N_8974,N_8833);
or U9024 (N_9024,N_8908,N_8866);
and U9025 (N_9025,N_8806,N_8889);
nand U9026 (N_9026,N_8938,N_8960);
or U9027 (N_9027,N_8805,N_8988);
nand U9028 (N_9028,N_8979,N_8976);
xnor U9029 (N_9029,N_8865,N_8920);
xnor U9030 (N_9030,N_8845,N_8933);
or U9031 (N_9031,N_8888,N_8913);
nand U9032 (N_9032,N_8841,N_8821);
nand U9033 (N_9033,N_8980,N_8818);
nor U9034 (N_9034,N_8926,N_8869);
xnor U9035 (N_9035,N_8839,N_8951);
nand U9036 (N_9036,N_8996,N_8897);
nand U9037 (N_9037,N_8968,N_8925);
xnor U9038 (N_9038,N_8940,N_8986);
nor U9039 (N_9039,N_8971,N_8952);
xnor U9040 (N_9040,N_8957,N_8993);
nand U9041 (N_9041,N_8981,N_8950);
nand U9042 (N_9042,N_8901,N_8916);
nand U9043 (N_9043,N_8902,N_8828);
and U9044 (N_9044,N_8847,N_8959);
and U9045 (N_9045,N_8843,N_8953);
nand U9046 (N_9046,N_8861,N_8945);
nor U9047 (N_9047,N_8803,N_8875);
nand U9048 (N_9048,N_8810,N_8882);
nand U9049 (N_9049,N_8874,N_8944);
or U9050 (N_9050,N_8840,N_8909);
or U9051 (N_9051,N_8977,N_8895);
and U9052 (N_9052,N_8804,N_8932);
and U9053 (N_9053,N_8886,N_8929);
and U9054 (N_9054,N_8807,N_8802);
nor U9055 (N_9055,N_8826,N_8830);
xnor U9056 (N_9056,N_8911,N_8864);
nor U9057 (N_9057,N_8935,N_8991);
nor U9058 (N_9058,N_8884,N_8924);
and U9059 (N_9059,N_8842,N_8893);
nor U9060 (N_9060,N_8870,N_8984);
nor U9061 (N_9061,N_8956,N_8948);
nor U9062 (N_9062,N_8975,N_8860);
xor U9063 (N_9063,N_8949,N_8814);
nand U9064 (N_9064,N_8813,N_8823);
xnor U9065 (N_9065,N_8885,N_8905);
nor U9066 (N_9066,N_8930,N_8997);
and U9067 (N_9067,N_8812,N_8855);
nor U9068 (N_9068,N_8836,N_8961);
nand U9069 (N_9069,N_8899,N_8863);
nand U9070 (N_9070,N_8848,N_8972);
or U9071 (N_9071,N_8809,N_8921);
nor U9072 (N_9072,N_8927,N_8983);
nand U9073 (N_9073,N_8858,N_8825);
xnor U9074 (N_9074,N_8928,N_8824);
and U9075 (N_9075,N_8811,N_8835);
nand U9076 (N_9076,N_8910,N_8817);
and U9077 (N_9077,N_8919,N_8990);
xnor U9078 (N_9078,N_8808,N_8989);
or U9079 (N_9079,N_8982,N_8887);
xnor U9080 (N_9080,N_8859,N_8896);
or U9081 (N_9081,N_8820,N_8936);
nand U9082 (N_9082,N_8881,N_8937);
nand U9083 (N_9083,N_8922,N_8970);
xnor U9084 (N_9084,N_8931,N_8854);
nor U9085 (N_9085,N_8832,N_8877);
xor U9086 (N_9086,N_8816,N_8872);
xor U9087 (N_9087,N_8962,N_8939);
xnor U9088 (N_9088,N_8891,N_8998);
xnor U9089 (N_9089,N_8871,N_8994);
nor U9090 (N_9090,N_8868,N_8992);
nand U9091 (N_9091,N_8966,N_8862);
nand U9092 (N_9092,N_8844,N_8912);
xnor U9093 (N_9093,N_8955,N_8894);
nand U9094 (N_9094,N_8849,N_8903);
nand U9095 (N_9095,N_8978,N_8934);
nand U9096 (N_9096,N_8906,N_8815);
nor U9097 (N_9097,N_8987,N_8943);
nor U9098 (N_9098,N_8995,N_8999);
and U9099 (N_9099,N_8973,N_8873);
or U9100 (N_9100,N_8889,N_8844);
nor U9101 (N_9101,N_8957,N_8841);
xnor U9102 (N_9102,N_8897,N_8951);
and U9103 (N_9103,N_8984,N_8891);
nand U9104 (N_9104,N_8823,N_8922);
nor U9105 (N_9105,N_8991,N_8800);
nand U9106 (N_9106,N_8865,N_8939);
and U9107 (N_9107,N_8806,N_8937);
and U9108 (N_9108,N_8853,N_8825);
or U9109 (N_9109,N_8894,N_8901);
nand U9110 (N_9110,N_8915,N_8977);
and U9111 (N_9111,N_8879,N_8913);
and U9112 (N_9112,N_8810,N_8884);
xor U9113 (N_9113,N_8806,N_8939);
nor U9114 (N_9114,N_8813,N_8850);
and U9115 (N_9115,N_8989,N_8818);
nor U9116 (N_9116,N_8932,N_8837);
xnor U9117 (N_9117,N_8995,N_8864);
nand U9118 (N_9118,N_8948,N_8965);
and U9119 (N_9119,N_8893,N_8936);
nor U9120 (N_9120,N_8892,N_8912);
nor U9121 (N_9121,N_8839,N_8872);
nor U9122 (N_9122,N_8905,N_8933);
and U9123 (N_9123,N_8943,N_8985);
or U9124 (N_9124,N_8811,N_8922);
and U9125 (N_9125,N_8832,N_8857);
or U9126 (N_9126,N_8994,N_8980);
or U9127 (N_9127,N_8928,N_8814);
and U9128 (N_9128,N_8851,N_8903);
and U9129 (N_9129,N_8850,N_8867);
xnor U9130 (N_9130,N_8826,N_8889);
or U9131 (N_9131,N_8977,N_8835);
or U9132 (N_9132,N_8974,N_8964);
nor U9133 (N_9133,N_8894,N_8938);
xor U9134 (N_9134,N_8910,N_8994);
nand U9135 (N_9135,N_8954,N_8818);
xnor U9136 (N_9136,N_8839,N_8857);
or U9137 (N_9137,N_8845,N_8968);
and U9138 (N_9138,N_8843,N_8940);
and U9139 (N_9139,N_8875,N_8865);
nor U9140 (N_9140,N_8952,N_8805);
nor U9141 (N_9141,N_8899,N_8865);
or U9142 (N_9142,N_8919,N_8892);
and U9143 (N_9143,N_8835,N_8965);
nand U9144 (N_9144,N_8960,N_8977);
nand U9145 (N_9145,N_8995,N_8841);
and U9146 (N_9146,N_8879,N_8816);
or U9147 (N_9147,N_8906,N_8810);
nor U9148 (N_9148,N_8836,N_8994);
or U9149 (N_9149,N_8940,N_8887);
and U9150 (N_9150,N_8901,N_8918);
nor U9151 (N_9151,N_8874,N_8912);
nand U9152 (N_9152,N_8881,N_8847);
nand U9153 (N_9153,N_8922,N_8865);
or U9154 (N_9154,N_8828,N_8834);
nor U9155 (N_9155,N_8874,N_8910);
nand U9156 (N_9156,N_8848,N_8968);
nor U9157 (N_9157,N_8920,N_8810);
nand U9158 (N_9158,N_8838,N_8846);
nor U9159 (N_9159,N_8975,N_8926);
or U9160 (N_9160,N_8821,N_8935);
and U9161 (N_9161,N_8950,N_8922);
xnor U9162 (N_9162,N_8842,N_8809);
nand U9163 (N_9163,N_8956,N_8984);
xnor U9164 (N_9164,N_8827,N_8843);
nand U9165 (N_9165,N_8829,N_8901);
nand U9166 (N_9166,N_8883,N_8957);
or U9167 (N_9167,N_8842,N_8865);
nor U9168 (N_9168,N_8857,N_8831);
and U9169 (N_9169,N_8992,N_8827);
xor U9170 (N_9170,N_8997,N_8982);
xor U9171 (N_9171,N_8828,N_8865);
xor U9172 (N_9172,N_8938,N_8885);
nand U9173 (N_9173,N_8955,N_8983);
xor U9174 (N_9174,N_8927,N_8890);
nand U9175 (N_9175,N_8982,N_8828);
or U9176 (N_9176,N_8867,N_8825);
nand U9177 (N_9177,N_8923,N_8943);
and U9178 (N_9178,N_8945,N_8820);
nor U9179 (N_9179,N_8902,N_8895);
xor U9180 (N_9180,N_8890,N_8821);
nand U9181 (N_9181,N_8924,N_8806);
nand U9182 (N_9182,N_8976,N_8984);
nand U9183 (N_9183,N_8882,N_8971);
nor U9184 (N_9184,N_8961,N_8967);
or U9185 (N_9185,N_8999,N_8803);
nor U9186 (N_9186,N_8816,N_8887);
xnor U9187 (N_9187,N_8943,N_8986);
nor U9188 (N_9188,N_8905,N_8977);
or U9189 (N_9189,N_8967,N_8968);
or U9190 (N_9190,N_8861,N_8870);
xor U9191 (N_9191,N_8936,N_8917);
xor U9192 (N_9192,N_8969,N_8989);
xnor U9193 (N_9193,N_8866,N_8890);
xnor U9194 (N_9194,N_8828,N_8924);
nor U9195 (N_9195,N_8932,N_8830);
nor U9196 (N_9196,N_8961,N_8812);
nor U9197 (N_9197,N_8829,N_8810);
or U9198 (N_9198,N_8825,N_8988);
nor U9199 (N_9199,N_8876,N_8992);
and U9200 (N_9200,N_9079,N_9096);
nor U9201 (N_9201,N_9155,N_9082);
xor U9202 (N_9202,N_9195,N_9023);
or U9203 (N_9203,N_9090,N_9036);
nor U9204 (N_9204,N_9051,N_9194);
nor U9205 (N_9205,N_9144,N_9028);
nor U9206 (N_9206,N_9131,N_9069);
nor U9207 (N_9207,N_9008,N_9054);
nor U9208 (N_9208,N_9192,N_9127);
and U9209 (N_9209,N_9122,N_9197);
xnor U9210 (N_9210,N_9035,N_9093);
nand U9211 (N_9211,N_9040,N_9166);
nor U9212 (N_9212,N_9141,N_9123);
nand U9213 (N_9213,N_9180,N_9150);
and U9214 (N_9214,N_9129,N_9032);
nand U9215 (N_9215,N_9189,N_9016);
xnor U9216 (N_9216,N_9080,N_9047);
nor U9217 (N_9217,N_9067,N_9117);
nor U9218 (N_9218,N_9085,N_9038);
or U9219 (N_9219,N_9030,N_9113);
nand U9220 (N_9220,N_9136,N_9169);
or U9221 (N_9221,N_9039,N_9184);
and U9222 (N_9222,N_9041,N_9092);
and U9223 (N_9223,N_9125,N_9049);
xor U9224 (N_9224,N_9073,N_9172);
nor U9225 (N_9225,N_9132,N_9002);
and U9226 (N_9226,N_9171,N_9089);
and U9227 (N_9227,N_9074,N_9108);
nand U9228 (N_9228,N_9161,N_9095);
and U9229 (N_9229,N_9020,N_9027);
nor U9230 (N_9230,N_9182,N_9115);
or U9231 (N_9231,N_9181,N_9013);
xnor U9232 (N_9232,N_9101,N_9012);
xor U9233 (N_9233,N_9176,N_9071);
nand U9234 (N_9234,N_9138,N_9170);
nand U9235 (N_9235,N_9139,N_9137);
xor U9236 (N_9236,N_9151,N_9188);
and U9237 (N_9237,N_9061,N_9102);
xnor U9238 (N_9238,N_9072,N_9015);
or U9239 (N_9239,N_9050,N_9057);
and U9240 (N_9240,N_9199,N_9066);
nor U9241 (N_9241,N_9034,N_9059);
or U9242 (N_9242,N_9070,N_9168);
or U9243 (N_9243,N_9097,N_9118);
nand U9244 (N_9244,N_9135,N_9116);
nor U9245 (N_9245,N_9156,N_9065);
nand U9246 (N_9246,N_9109,N_9000);
nor U9247 (N_9247,N_9026,N_9148);
nand U9248 (N_9248,N_9100,N_9142);
and U9249 (N_9249,N_9005,N_9063);
and U9250 (N_9250,N_9190,N_9133);
nor U9251 (N_9251,N_9037,N_9178);
and U9252 (N_9252,N_9045,N_9044);
or U9253 (N_9253,N_9078,N_9186);
nand U9254 (N_9254,N_9198,N_9031);
nand U9255 (N_9255,N_9140,N_9152);
xor U9256 (N_9256,N_9087,N_9098);
nor U9257 (N_9257,N_9009,N_9105);
nand U9258 (N_9258,N_9185,N_9162);
nand U9259 (N_9259,N_9058,N_9042);
or U9260 (N_9260,N_9025,N_9126);
or U9261 (N_9261,N_9173,N_9165);
or U9262 (N_9262,N_9158,N_9111);
nor U9263 (N_9263,N_9106,N_9154);
nand U9264 (N_9264,N_9104,N_9048);
or U9265 (N_9265,N_9088,N_9147);
and U9266 (N_9266,N_9145,N_9064);
xor U9267 (N_9267,N_9004,N_9068);
and U9268 (N_9268,N_9052,N_9014);
xnor U9269 (N_9269,N_9177,N_9120);
nand U9270 (N_9270,N_9112,N_9083);
xnor U9271 (N_9271,N_9157,N_9022);
and U9272 (N_9272,N_9110,N_9010);
nand U9273 (N_9273,N_9159,N_9060);
and U9274 (N_9274,N_9077,N_9076);
and U9275 (N_9275,N_9174,N_9033);
xnor U9276 (N_9276,N_9196,N_9011);
or U9277 (N_9277,N_9018,N_9075);
nor U9278 (N_9278,N_9124,N_9006);
or U9279 (N_9279,N_9107,N_9175);
xor U9280 (N_9280,N_9084,N_9001);
and U9281 (N_9281,N_9029,N_9146);
or U9282 (N_9282,N_9119,N_9163);
nand U9283 (N_9283,N_9149,N_9021);
nand U9284 (N_9284,N_9007,N_9164);
nor U9285 (N_9285,N_9183,N_9056);
xor U9286 (N_9286,N_9179,N_9046);
xnor U9287 (N_9287,N_9160,N_9167);
and U9288 (N_9288,N_9134,N_9128);
and U9289 (N_9289,N_9114,N_9103);
and U9290 (N_9290,N_9143,N_9017);
nor U9291 (N_9291,N_9024,N_9099);
and U9292 (N_9292,N_9121,N_9081);
or U9293 (N_9293,N_9094,N_9153);
nor U9294 (N_9294,N_9053,N_9086);
and U9295 (N_9295,N_9187,N_9193);
and U9296 (N_9296,N_9019,N_9043);
nand U9297 (N_9297,N_9062,N_9130);
or U9298 (N_9298,N_9191,N_9055);
or U9299 (N_9299,N_9003,N_9091);
xor U9300 (N_9300,N_9089,N_9115);
xnor U9301 (N_9301,N_9039,N_9165);
nand U9302 (N_9302,N_9048,N_9138);
or U9303 (N_9303,N_9040,N_9137);
nand U9304 (N_9304,N_9162,N_9066);
or U9305 (N_9305,N_9013,N_9049);
nor U9306 (N_9306,N_9193,N_9136);
nor U9307 (N_9307,N_9026,N_9082);
xnor U9308 (N_9308,N_9092,N_9159);
nand U9309 (N_9309,N_9169,N_9004);
and U9310 (N_9310,N_9104,N_9022);
and U9311 (N_9311,N_9088,N_9154);
nor U9312 (N_9312,N_9053,N_9148);
or U9313 (N_9313,N_9074,N_9096);
nand U9314 (N_9314,N_9024,N_9191);
nand U9315 (N_9315,N_9063,N_9032);
or U9316 (N_9316,N_9094,N_9198);
or U9317 (N_9317,N_9198,N_9037);
nor U9318 (N_9318,N_9081,N_9102);
and U9319 (N_9319,N_9185,N_9104);
nand U9320 (N_9320,N_9026,N_9037);
or U9321 (N_9321,N_9048,N_9074);
nand U9322 (N_9322,N_9181,N_9175);
nand U9323 (N_9323,N_9080,N_9139);
and U9324 (N_9324,N_9014,N_9085);
and U9325 (N_9325,N_9046,N_9103);
xnor U9326 (N_9326,N_9170,N_9177);
nand U9327 (N_9327,N_9140,N_9053);
nand U9328 (N_9328,N_9151,N_9096);
xor U9329 (N_9329,N_9173,N_9026);
or U9330 (N_9330,N_9148,N_9107);
nor U9331 (N_9331,N_9126,N_9019);
nor U9332 (N_9332,N_9078,N_9053);
or U9333 (N_9333,N_9021,N_9170);
nor U9334 (N_9334,N_9078,N_9190);
nand U9335 (N_9335,N_9197,N_9089);
nor U9336 (N_9336,N_9157,N_9174);
and U9337 (N_9337,N_9063,N_9194);
nand U9338 (N_9338,N_9096,N_9189);
xor U9339 (N_9339,N_9072,N_9170);
or U9340 (N_9340,N_9090,N_9092);
nand U9341 (N_9341,N_9100,N_9063);
nand U9342 (N_9342,N_9057,N_9012);
and U9343 (N_9343,N_9064,N_9148);
or U9344 (N_9344,N_9182,N_9128);
nand U9345 (N_9345,N_9127,N_9161);
nand U9346 (N_9346,N_9000,N_9147);
nor U9347 (N_9347,N_9046,N_9148);
and U9348 (N_9348,N_9024,N_9169);
or U9349 (N_9349,N_9193,N_9129);
or U9350 (N_9350,N_9157,N_9035);
and U9351 (N_9351,N_9182,N_9188);
xor U9352 (N_9352,N_9195,N_9199);
xor U9353 (N_9353,N_9072,N_9043);
and U9354 (N_9354,N_9008,N_9129);
nor U9355 (N_9355,N_9140,N_9190);
and U9356 (N_9356,N_9002,N_9063);
nand U9357 (N_9357,N_9108,N_9011);
nor U9358 (N_9358,N_9143,N_9015);
nand U9359 (N_9359,N_9107,N_9164);
and U9360 (N_9360,N_9196,N_9111);
xnor U9361 (N_9361,N_9170,N_9095);
or U9362 (N_9362,N_9102,N_9071);
xor U9363 (N_9363,N_9034,N_9071);
nor U9364 (N_9364,N_9141,N_9179);
and U9365 (N_9365,N_9144,N_9006);
and U9366 (N_9366,N_9152,N_9150);
and U9367 (N_9367,N_9115,N_9049);
nand U9368 (N_9368,N_9061,N_9069);
or U9369 (N_9369,N_9017,N_9165);
and U9370 (N_9370,N_9161,N_9056);
and U9371 (N_9371,N_9164,N_9009);
nand U9372 (N_9372,N_9152,N_9188);
and U9373 (N_9373,N_9044,N_9027);
nand U9374 (N_9374,N_9136,N_9065);
xor U9375 (N_9375,N_9147,N_9025);
and U9376 (N_9376,N_9029,N_9008);
nor U9377 (N_9377,N_9185,N_9166);
or U9378 (N_9378,N_9153,N_9145);
xnor U9379 (N_9379,N_9160,N_9115);
nor U9380 (N_9380,N_9073,N_9039);
nor U9381 (N_9381,N_9066,N_9107);
and U9382 (N_9382,N_9142,N_9159);
nor U9383 (N_9383,N_9187,N_9134);
nor U9384 (N_9384,N_9182,N_9102);
or U9385 (N_9385,N_9061,N_9143);
and U9386 (N_9386,N_9178,N_9082);
or U9387 (N_9387,N_9189,N_9186);
nand U9388 (N_9388,N_9101,N_9130);
or U9389 (N_9389,N_9177,N_9116);
xor U9390 (N_9390,N_9180,N_9026);
nor U9391 (N_9391,N_9182,N_9181);
or U9392 (N_9392,N_9101,N_9141);
and U9393 (N_9393,N_9086,N_9084);
and U9394 (N_9394,N_9017,N_9122);
nor U9395 (N_9395,N_9095,N_9032);
and U9396 (N_9396,N_9155,N_9190);
xnor U9397 (N_9397,N_9087,N_9013);
nand U9398 (N_9398,N_9177,N_9142);
xnor U9399 (N_9399,N_9071,N_9086);
xnor U9400 (N_9400,N_9216,N_9232);
or U9401 (N_9401,N_9291,N_9264);
or U9402 (N_9402,N_9347,N_9219);
nor U9403 (N_9403,N_9339,N_9290);
nand U9404 (N_9404,N_9314,N_9317);
or U9405 (N_9405,N_9340,N_9354);
and U9406 (N_9406,N_9235,N_9334);
nand U9407 (N_9407,N_9330,N_9297);
nand U9408 (N_9408,N_9213,N_9221);
xor U9409 (N_9409,N_9214,N_9274);
xnor U9410 (N_9410,N_9272,N_9395);
or U9411 (N_9411,N_9326,N_9351);
nand U9412 (N_9412,N_9391,N_9217);
nor U9413 (N_9413,N_9335,N_9275);
or U9414 (N_9414,N_9323,N_9236);
nor U9415 (N_9415,N_9390,N_9293);
or U9416 (N_9416,N_9252,N_9386);
xor U9417 (N_9417,N_9228,N_9307);
nor U9418 (N_9418,N_9229,N_9282);
or U9419 (N_9419,N_9284,N_9300);
nand U9420 (N_9420,N_9355,N_9318);
nand U9421 (N_9421,N_9273,N_9346);
or U9422 (N_9422,N_9369,N_9200);
nor U9423 (N_9423,N_9234,N_9279);
and U9424 (N_9424,N_9315,N_9220);
xnor U9425 (N_9425,N_9376,N_9289);
xor U9426 (N_9426,N_9356,N_9254);
xor U9427 (N_9427,N_9247,N_9375);
nor U9428 (N_9428,N_9338,N_9305);
and U9429 (N_9429,N_9287,N_9206);
xor U9430 (N_9430,N_9222,N_9238);
and U9431 (N_9431,N_9371,N_9246);
and U9432 (N_9432,N_9364,N_9295);
and U9433 (N_9433,N_9202,N_9309);
nand U9434 (N_9434,N_9208,N_9283);
nand U9435 (N_9435,N_9316,N_9336);
and U9436 (N_9436,N_9262,N_9261);
xnor U9437 (N_9437,N_9393,N_9327);
and U9438 (N_9438,N_9313,N_9243);
and U9439 (N_9439,N_9268,N_9223);
and U9440 (N_9440,N_9399,N_9227);
or U9441 (N_9441,N_9368,N_9259);
xnor U9442 (N_9442,N_9245,N_9203);
and U9443 (N_9443,N_9266,N_9251);
and U9444 (N_9444,N_9281,N_9392);
or U9445 (N_9445,N_9280,N_9269);
nor U9446 (N_9446,N_9302,N_9348);
nor U9447 (N_9447,N_9296,N_9384);
or U9448 (N_9448,N_9398,N_9212);
and U9449 (N_9449,N_9341,N_9304);
or U9450 (N_9450,N_9357,N_9366);
xor U9451 (N_9451,N_9237,N_9270);
nor U9452 (N_9452,N_9210,N_9358);
or U9453 (N_9453,N_9311,N_9207);
nand U9454 (N_9454,N_9324,N_9362);
xnor U9455 (N_9455,N_9382,N_9342);
xnor U9456 (N_9456,N_9383,N_9285);
and U9457 (N_9457,N_9301,N_9380);
xor U9458 (N_9458,N_9263,N_9396);
or U9459 (N_9459,N_9292,N_9226);
nor U9460 (N_9460,N_9265,N_9388);
xor U9461 (N_9461,N_9288,N_9225);
or U9462 (N_9462,N_9378,N_9387);
nor U9463 (N_9463,N_9278,N_9240);
or U9464 (N_9464,N_9257,N_9394);
nand U9465 (N_9465,N_9361,N_9353);
and U9466 (N_9466,N_9255,N_9244);
and U9467 (N_9467,N_9271,N_9201);
xnor U9468 (N_9468,N_9322,N_9385);
or U9469 (N_9469,N_9320,N_9211);
nand U9470 (N_9470,N_9333,N_9360);
nor U9471 (N_9471,N_9294,N_9205);
and U9472 (N_9472,N_9381,N_9329);
xor U9473 (N_9473,N_9312,N_9250);
nor U9474 (N_9474,N_9258,N_9242);
nand U9475 (N_9475,N_9204,N_9350);
and U9476 (N_9476,N_9260,N_9332);
xnor U9477 (N_9477,N_9215,N_9343);
or U9478 (N_9478,N_9373,N_9321);
or U9479 (N_9479,N_9352,N_9359);
and U9480 (N_9480,N_9276,N_9256);
or U9481 (N_9481,N_9224,N_9370);
nand U9482 (N_9482,N_9377,N_9241);
and U9483 (N_9483,N_9349,N_9298);
or U9484 (N_9484,N_9389,N_9218);
xnor U9485 (N_9485,N_9367,N_9286);
nor U9486 (N_9486,N_9209,N_9253);
xor U9487 (N_9487,N_9397,N_9233);
or U9488 (N_9488,N_9345,N_9308);
nor U9489 (N_9489,N_9249,N_9303);
and U9490 (N_9490,N_9379,N_9363);
xnor U9491 (N_9491,N_9319,N_9344);
nand U9492 (N_9492,N_9306,N_9248);
nand U9493 (N_9493,N_9328,N_9372);
nand U9494 (N_9494,N_9337,N_9277);
and U9495 (N_9495,N_9365,N_9267);
nor U9496 (N_9496,N_9230,N_9310);
nand U9497 (N_9497,N_9239,N_9325);
or U9498 (N_9498,N_9231,N_9299);
and U9499 (N_9499,N_9331,N_9374);
nand U9500 (N_9500,N_9233,N_9268);
and U9501 (N_9501,N_9336,N_9216);
and U9502 (N_9502,N_9308,N_9334);
and U9503 (N_9503,N_9393,N_9218);
xnor U9504 (N_9504,N_9230,N_9278);
nand U9505 (N_9505,N_9241,N_9353);
or U9506 (N_9506,N_9307,N_9264);
nand U9507 (N_9507,N_9200,N_9327);
and U9508 (N_9508,N_9263,N_9214);
or U9509 (N_9509,N_9369,N_9259);
and U9510 (N_9510,N_9307,N_9252);
xnor U9511 (N_9511,N_9215,N_9275);
xnor U9512 (N_9512,N_9304,N_9331);
or U9513 (N_9513,N_9371,N_9292);
nand U9514 (N_9514,N_9242,N_9206);
or U9515 (N_9515,N_9343,N_9286);
or U9516 (N_9516,N_9388,N_9253);
nand U9517 (N_9517,N_9232,N_9282);
xor U9518 (N_9518,N_9299,N_9338);
nor U9519 (N_9519,N_9213,N_9382);
and U9520 (N_9520,N_9383,N_9229);
or U9521 (N_9521,N_9201,N_9376);
and U9522 (N_9522,N_9304,N_9384);
or U9523 (N_9523,N_9272,N_9313);
nor U9524 (N_9524,N_9209,N_9248);
or U9525 (N_9525,N_9273,N_9307);
and U9526 (N_9526,N_9353,N_9214);
or U9527 (N_9527,N_9203,N_9210);
nor U9528 (N_9528,N_9352,N_9307);
nand U9529 (N_9529,N_9366,N_9219);
or U9530 (N_9530,N_9291,N_9364);
nand U9531 (N_9531,N_9292,N_9257);
and U9532 (N_9532,N_9365,N_9303);
nand U9533 (N_9533,N_9292,N_9385);
nor U9534 (N_9534,N_9348,N_9384);
or U9535 (N_9535,N_9399,N_9398);
nand U9536 (N_9536,N_9364,N_9356);
and U9537 (N_9537,N_9381,N_9393);
and U9538 (N_9538,N_9366,N_9359);
nand U9539 (N_9539,N_9265,N_9254);
and U9540 (N_9540,N_9334,N_9348);
xor U9541 (N_9541,N_9374,N_9369);
xnor U9542 (N_9542,N_9311,N_9281);
nor U9543 (N_9543,N_9379,N_9259);
or U9544 (N_9544,N_9272,N_9355);
xor U9545 (N_9545,N_9250,N_9232);
and U9546 (N_9546,N_9221,N_9318);
xnor U9547 (N_9547,N_9310,N_9330);
nand U9548 (N_9548,N_9398,N_9358);
nand U9549 (N_9549,N_9274,N_9332);
and U9550 (N_9550,N_9229,N_9276);
or U9551 (N_9551,N_9314,N_9334);
xnor U9552 (N_9552,N_9346,N_9215);
and U9553 (N_9553,N_9315,N_9319);
nand U9554 (N_9554,N_9336,N_9369);
and U9555 (N_9555,N_9316,N_9245);
nor U9556 (N_9556,N_9307,N_9208);
or U9557 (N_9557,N_9217,N_9247);
or U9558 (N_9558,N_9377,N_9355);
xnor U9559 (N_9559,N_9282,N_9201);
or U9560 (N_9560,N_9321,N_9280);
or U9561 (N_9561,N_9315,N_9296);
nand U9562 (N_9562,N_9365,N_9208);
nor U9563 (N_9563,N_9335,N_9222);
and U9564 (N_9564,N_9351,N_9362);
xnor U9565 (N_9565,N_9364,N_9377);
xor U9566 (N_9566,N_9242,N_9302);
or U9567 (N_9567,N_9215,N_9296);
nor U9568 (N_9568,N_9311,N_9350);
or U9569 (N_9569,N_9364,N_9248);
or U9570 (N_9570,N_9368,N_9340);
nor U9571 (N_9571,N_9239,N_9315);
and U9572 (N_9572,N_9375,N_9248);
nand U9573 (N_9573,N_9282,N_9386);
xor U9574 (N_9574,N_9356,N_9375);
and U9575 (N_9575,N_9256,N_9242);
nand U9576 (N_9576,N_9247,N_9219);
xor U9577 (N_9577,N_9285,N_9200);
and U9578 (N_9578,N_9245,N_9343);
xnor U9579 (N_9579,N_9383,N_9272);
nor U9580 (N_9580,N_9370,N_9249);
and U9581 (N_9581,N_9296,N_9279);
nand U9582 (N_9582,N_9383,N_9231);
or U9583 (N_9583,N_9391,N_9340);
and U9584 (N_9584,N_9343,N_9291);
and U9585 (N_9585,N_9216,N_9252);
nor U9586 (N_9586,N_9394,N_9300);
xnor U9587 (N_9587,N_9248,N_9293);
nand U9588 (N_9588,N_9218,N_9376);
and U9589 (N_9589,N_9375,N_9262);
xnor U9590 (N_9590,N_9335,N_9283);
xor U9591 (N_9591,N_9206,N_9224);
xor U9592 (N_9592,N_9274,N_9324);
nand U9593 (N_9593,N_9274,N_9397);
nand U9594 (N_9594,N_9307,N_9318);
and U9595 (N_9595,N_9338,N_9366);
nand U9596 (N_9596,N_9386,N_9288);
nand U9597 (N_9597,N_9275,N_9207);
nand U9598 (N_9598,N_9350,N_9242);
xnor U9599 (N_9599,N_9358,N_9246);
nor U9600 (N_9600,N_9526,N_9454);
xnor U9601 (N_9601,N_9580,N_9474);
xnor U9602 (N_9602,N_9553,N_9442);
and U9603 (N_9603,N_9486,N_9570);
nand U9604 (N_9604,N_9517,N_9531);
xor U9605 (N_9605,N_9552,N_9471);
nor U9606 (N_9606,N_9484,N_9549);
nor U9607 (N_9607,N_9511,N_9573);
and U9608 (N_9608,N_9406,N_9502);
nor U9609 (N_9609,N_9566,N_9451);
nand U9610 (N_9610,N_9492,N_9404);
nor U9611 (N_9611,N_9488,N_9555);
xor U9612 (N_9612,N_9528,N_9495);
xnor U9613 (N_9613,N_9537,N_9550);
nand U9614 (N_9614,N_9463,N_9575);
nand U9615 (N_9615,N_9587,N_9571);
xor U9616 (N_9616,N_9548,N_9532);
nor U9617 (N_9617,N_9411,N_9529);
or U9618 (N_9618,N_9408,N_9512);
xor U9619 (N_9619,N_9522,N_9459);
or U9620 (N_9620,N_9591,N_9400);
nor U9621 (N_9621,N_9498,N_9579);
nor U9622 (N_9622,N_9556,N_9534);
nor U9623 (N_9623,N_9443,N_9530);
nand U9624 (N_9624,N_9428,N_9562);
xor U9625 (N_9625,N_9516,N_9569);
nor U9626 (N_9626,N_9405,N_9494);
or U9627 (N_9627,N_9563,N_9430);
nand U9628 (N_9628,N_9567,N_9527);
nor U9629 (N_9629,N_9559,N_9444);
nand U9630 (N_9630,N_9506,N_9477);
xnor U9631 (N_9631,N_9478,N_9423);
nand U9632 (N_9632,N_9499,N_9476);
and U9633 (N_9633,N_9427,N_9447);
nand U9634 (N_9634,N_9504,N_9541);
or U9635 (N_9635,N_9565,N_9435);
and U9636 (N_9636,N_9433,N_9581);
and U9637 (N_9637,N_9588,N_9401);
and U9638 (N_9638,N_9544,N_9479);
xnor U9639 (N_9639,N_9420,N_9410);
xor U9640 (N_9640,N_9460,N_9578);
and U9641 (N_9641,N_9542,N_9576);
or U9642 (N_9642,N_9409,N_9590);
nor U9643 (N_9643,N_9585,N_9449);
xor U9644 (N_9644,N_9545,N_9521);
xor U9645 (N_9645,N_9437,N_9536);
nand U9646 (N_9646,N_9508,N_9535);
nor U9647 (N_9647,N_9465,N_9461);
nor U9648 (N_9648,N_9558,N_9543);
and U9649 (N_9649,N_9472,N_9574);
nor U9650 (N_9650,N_9414,N_9593);
xor U9651 (N_9651,N_9418,N_9524);
nand U9652 (N_9652,N_9490,N_9462);
and U9653 (N_9653,N_9547,N_9491);
or U9654 (N_9654,N_9525,N_9440);
or U9655 (N_9655,N_9425,N_9557);
xnor U9656 (N_9656,N_9583,N_9452);
nand U9657 (N_9657,N_9515,N_9470);
xnor U9658 (N_9658,N_9469,N_9586);
nand U9659 (N_9659,N_9480,N_9501);
and U9660 (N_9660,N_9450,N_9482);
nor U9661 (N_9661,N_9468,N_9592);
or U9662 (N_9662,N_9466,N_9483);
xnor U9663 (N_9663,N_9438,N_9513);
and U9664 (N_9664,N_9467,N_9445);
or U9665 (N_9665,N_9432,N_9439);
or U9666 (N_9666,N_9599,N_9485);
xor U9667 (N_9667,N_9458,N_9510);
and U9668 (N_9668,N_9596,N_9407);
and U9669 (N_9669,N_9598,N_9554);
and U9670 (N_9670,N_9572,N_9497);
xor U9671 (N_9671,N_9518,N_9520);
and U9672 (N_9672,N_9503,N_9533);
xnor U9673 (N_9673,N_9514,N_9403);
or U9674 (N_9674,N_9446,N_9582);
nor U9675 (N_9675,N_9546,N_9561);
or U9676 (N_9676,N_9594,N_9424);
and U9677 (N_9677,N_9584,N_9496);
and U9678 (N_9678,N_9489,N_9473);
and U9679 (N_9679,N_9422,N_9412);
nor U9680 (N_9680,N_9507,N_9419);
nand U9681 (N_9681,N_9595,N_9568);
nand U9682 (N_9682,N_9481,N_9500);
xor U9683 (N_9683,N_9413,N_9417);
nor U9684 (N_9684,N_9589,N_9402);
xor U9685 (N_9685,N_9577,N_9509);
or U9686 (N_9686,N_9453,N_9539);
or U9687 (N_9687,N_9421,N_9416);
and U9688 (N_9688,N_9597,N_9505);
nand U9689 (N_9689,N_9540,N_9434);
nand U9690 (N_9690,N_9415,N_9441);
xor U9691 (N_9691,N_9551,N_9564);
and U9692 (N_9692,N_9431,N_9523);
nor U9693 (N_9693,N_9464,N_9426);
nand U9694 (N_9694,N_9448,N_9538);
or U9695 (N_9695,N_9457,N_9436);
xnor U9696 (N_9696,N_9456,N_9429);
nand U9697 (N_9697,N_9519,N_9475);
nor U9698 (N_9698,N_9487,N_9455);
xnor U9699 (N_9699,N_9493,N_9560);
or U9700 (N_9700,N_9403,N_9439);
and U9701 (N_9701,N_9433,N_9563);
nor U9702 (N_9702,N_9490,N_9467);
xnor U9703 (N_9703,N_9595,N_9485);
nand U9704 (N_9704,N_9584,N_9502);
nor U9705 (N_9705,N_9445,N_9503);
and U9706 (N_9706,N_9483,N_9590);
or U9707 (N_9707,N_9501,N_9447);
nand U9708 (N_9708,N_9481,N_9483);
nor U9709 (N_9709,N_9464,N_9568);
nand U9710 (N_9710,N_9476,N_9514);
xor U9711 (N_9711,N_9498,N_9593);
or U9712 (N_9712,N_9452,N_9489);
nand U9713 (N_9713,N_9515,N_9487);
xor U9714 (N_9714,N_9403,N_9550);
nand U9715 (N_9715,N_9565,N_9503);
or U9716 (N_9716,N_9561,N_9524);
nand U9717 (N_9717,N_9532,N_9493);
and U9718 (N_9718,N_9533,N_9577);
nand U9719 (N_9719,N_9463,N_9514);
nand U9720 (N_9720,N_9510,N_9473);
or U9721 (N_9721,N_9521,N_9514);
and U9722 (N_9722,N_9590,N_9551);
and U9723 (N_9723,N_9539,N_9457);
or U9724 (N_9724,N_9498,N_9562);
nand U9725 (N_9725,N_9498,N_9496);
nand U9726 (N_9726,N_9440,N_9435);
nor U9727 (N_9727,N_9420,N_9400);
nor U9728 (N_9728,N_9521,N_9458);
nor U9729 (N_9729,N_9465,N_9544);
xnor U9730 (N_9730,N_9465,N_9558);
or U9731 (N_9731,N_9464,N_9441);
xnor U9732 (N_9732,N_9430,N_9468);
nor U9733 (N_9733,N_9440,N_9595);
nand U9734 (N_9734,N_9540,N_9478);
nor U9735 (N_9735,N_9446,N_9400);
or U9736 (N_9736,N_9493,N_9438);
and U9737 (N_9737,N_9454,N_9562);
and U9738 (N_9738,N_9584,N_9551);
and U9739 (N_9739,N_9545,N_9467);
and U9740 (N_9740,N_9564,N_9585);
or U9741 (N_9741,N_9448,N_9572);
nand U9742 (N_9742,N_9507,N_9452);
and U9743 (N_9743,N_9481,N_9475);
xnor U9744 (N_9744,N_9514,N_9536);
nand U9745 (N_9745,N_9582,N_9467);
or U9746 (N_9746,N_9526,N_9570);
or U9747 (N_9747,N_9518,N_9494);
nor U9748 (N_9748,N_9545,N_9446);
nand U9749 (N_9749,N_9429,N_9586);
nor U9750 (N_9750,N_9415,N_9463);
xor U9751 (N_9751,N_9438,N_9445);
xor U9752 (N_9752,N_9437,N_9559);
or U9753 (N_9753,N_9466,N_9462);
or U9754 (N_9754,N_9420,N_9497);
nor U9755 (N_9755,N_9542,N_9451);
nand U9756 (N_9756,N_9486,N_9489);
nor U9757 (N_9757,N_9549,N_9459);
or U9758 (N_9758,N_9499,N_9540);
or U9759 (N_9759,N_9561,N_9462);
and U9760 (N_9760,N_9429,N_9599);
xor U9761 (N_9761,N_9538,N_9572);
xnor U9762 (N_9762,N_9576,N_9512);
or U9763 (N_9763,N_9401,N_9410);
nand U9764 (N_9764,N_9551,N_9431);
nor U9765 (N_9765,N_9446,N_9530);
xor U9766 (N_9766,N_9474,N_9539);
or U9767 (N_9767,N_9457,N_9475);
or U9768 (N_9768,N_9503,N_9464);
and U9769 (N_9769,N_9494,N_9520);
xor U9770 (N_9770,N_9584,N_9463);
xor U9771 (N_9771,N_9568,N_9482);
nand U9772 (N_9772,N_9524,N_9488);
nor U9773 (N_9773,N_9451,N_9523);
nand U9774 (N_9774,N_9450,N_9547);
and U9775 (N_9775,N_9585,N_9424);
nor U9776 (N_9776,N_9436,N_9495);
or U9777 (N_9777,N_9410,N_9460);
nand U9778 (N_9778,N_9494,N_9577);
nor U9779 (N_9779,N_9421,N_9502);
or U9780 (N_9780,N_9437,N_9586);
and U9781 (N_9781,N_9471,N_9425);
nand U9782 (N_9782,N_9567,N_9554);
xor U9783 (N_9783,N_9462,N_9481);
or U9784 (N_9784,N_9497,N_9536);
and U9785 (N_9785,N_9487,N_9517);
nor U9786 (N_9786,N_9521,N_9443);
or U9787 (N_9787,N_9429,N_9425);
nor U9788 (N_9788,N_9475,N_9442);
xnor U9789 (N_9789,N_9574,N_9515);
and U9790 (N_9790,N_9586,N_9438);
nand U9791 (N_9791,N_9464,N_9518);
nand U9792 (N_9792,N_9444,N_9463);
nand U9793 (N_9793,N_9428,N_9559);
xnor U9794 (N_9794,N_9435,N_9473);
and U9795 (N_9795,N_9440,N_9540);
nand U9796 (N_9796,N_9517,N_9490);
and U9797 (N_9797,N_9457,N_9462);
xnor U9798 (N_9798,N_9556,N_9480);
nor U9799 (N_9799,N_9479,N_9428);
xor U9800 (N_9800,N_9755,N_9642);
or U9801 (N_9801,N_9756,N_9781);
nor U9802 (N_9802,N_9796,N_9789);
xnor U9803 (N_9803,N_9744,N_9695);
nor U9804 (N_9804,N_9670,N_9646);
nor U9805 (N_9805,N_9636,N_9624);
and U9806 (N_9806,N_9658,N_9737);
or U9807 (N_9807,N_9612,N_9640);
nand U9808 (N_9808,N_9703,N_9627);
nand U9809 (N_9809,N_9792,N_9600);
or U9810 (N_9810,N_9671,N_9641);
nor U9811 (N_9811,N_9794,N_9793);
nand U9812 (N_9812,N_9639,N_9678);
xor U9813 (N_9813,N_9607,N_9662);
xor U9814 (N_9814,N_9654,N_9777);
or U9815 (N_9815,N_9606,N_9660);
and U9816 (N_9816,N_9644,N_9619);
and U9817 (N_9817,N_9667,N_9690);
and U9818 (N_9818,N_9725,N_9766);
nand U9819 (N_9819,N_9790,N_9706);
or U9820 (N_9820,N_9668,N_9778);
nand U9821 (N_9821,N_9645,N_9738);
and U9822 (N_9822,N_9773,N_9722);
or U9823 (N_9823,N_9760,N_9724);
nor U9824 (N_9824,N_9783,N_9776);
nor U9825 (N_9825,N_9748,N_9715);
nor U9826 (N_9826,N_9700,N_9797);
or U9827 (N_9827,N_9677,N_9732);
or U9828 (N_9828,N_9689,N_9665);
or U9829 (N_9829,N_9650,N_9702);
nand U9830 (N_9830,N_9649,N_9674);
nand U9831 (N_9831,N_9617,N_9782);
or U9832 (N_9832,N_9740,N_9770);
and U9833 (N_9833,N_9692,N_9618);
or U9834 (N_9834,N_9684,N_9635);
or U9835 (N_9835,N_9746,N_9727);
nand U9836 (N_9836,N_9716,N_9758);
nor U9837 (N_9837,N_9704,N_9799);
nor U9838 (N_9838,N_9752,N_9780);
xnor U9839 (N_9839,N_9775,N_9718);
xor U9840 (N_9840,N_9651,N_9736);
nand U9841 (N_9841,N_9643,N_9714);
or U9842 (N_9842,N_9628,N_9767);
nand U9843 (N_9843,N_9669,N_9763);
nor U9844 (N_9844,N_9726,N_9620);
nand U9845 (N_9845,N_9647,N_9601);
or U9846 (N_9846,N_9788,N_9705);
and U9847 (N_9847,N_9629,N_9675);
xnor U9848 (N_9848,N_9786,N_9753);
xor U9849 (N_9849,N_9663,N_9656);
xor U9850 (N_9850,N_9698,N_9623);
or U9851 (N_9851,N_9791,N_9614);
xnor U9852 (N_9852,N_9679,N_9608);
or U9853 (N_9853,N_9648,N_9734);
and U9854 (N_9854,N_9661,N_9685);
and U9855 (N_9855,N_9739,N_9731);
nand U9856 (N_9856,N_9632,N_9615);
or U9857 (N_9857,N_9723,N_9613);
nor U9858 (N_9858,N_9733,N_9762);
nor U9859 (N_9859,N_9750,N_9621);
and U9860 (N_9860,N_9699,N_9764);
and U9861 (N_9861,N_9701,N_9697);
and U9862 (N_9862,N_9728,N_9754);
and U9863 (N_9863,N_9603,N_9779);
nor U9864 (N_9864,N_9798,N_9693);
nand U9865 (N_9865,N_9711,N_9719);
nand U9866 (N_9866,N_9768,N_9771);
nor U9867 (N_9867,N_9659,N_9729);
nand U9868 (N_9868,N_9712,N_9741);
xor U9869 (N_9869,N_9696,N_9717);
xor U9870 (N_9870,N_9604,N_9682);
nand U9871 (N_9871,N_9652,N_9747);
nand U9872 (N_9872,N_9631,N_9630);
or U9873 (N_9873,N_9676,N_9673);
nor U9874 (N_9874,N_9681,N_9683);
xnor U9875 (N_9875,N_9655,N_9795);
and U9876 (N_9876,N_9657,N_9672);
nand U9877 (N_9877,N_9721,N_9765);
nand U9878 (N_9878,N_9785,N_9745);
or U9879 (N_9879,N_9759,N_9616);
xor U9880 (N_9880,N_9713,N_9694);
or U9881 (N_9881,N_9602,N_9708);
xnor U9882 (N_9882,N_9749,N_9634);
or U9883 (N_9883,N_9688,N_9720);
xnor U9884 (N_9884,N_9743,N_9687);
and U9885 (N_9885,N_9735,N_9730);
nor U9886 (N_9886,N_9761,N_9680);
or U9887 (N_9887,N_9769,N_9751);
or U9888 (N_9888,N_9691,N_9638);
xnor U9889 (N_9889,N_9653,N_9742);
and U9890 (N_9890,N_9710,N_9707);
nand U9891 (N_9891,N_9633,N_9686);
nand U9892 (N_9892,N_9622,N_9637);
and U9893 (N_9893,N_9787,N_9757);
or U9894 (N_9894,N_9609,N_9610);
and U9895 (N_9895,N_9772,N_9625);
nand U9896 (N_9896,N_9666,N_9774);
and U9897 (N_9897,N_9611,N_9605);
nor U9898 (N_9898,N_9709,N_9664);
and U9899 (N_9899,N_9626,N_9784);
or U9900 (N_9900,N_9726,N_9652);
or U9901 (N_9901,N_9655,N_9736);
and U9902 (N_9902,N_9673,N_9681);
nor U9903 (N_9903,N_9607,N_9675);
nand U9904 (N_9904,N_9669,N_9689);
xor U9905 (N_9905,N_9712,N_9685);
xnor U9906 (N_9906,N_9682,N_9727);
xnor U9907 (N_9907,N_9716,N_9655);
or U9908 (N_9908,N_9724,N_9711);
and U9909 (N_9909,N_9747,N_9609);
or U9910 (N_9910,N_9689,N_9605);
xor U9911 (N_9911,N_9633,N_9750);
or U9912 (N_9912,N_9696,N_9610);
nand U9913 (N_9913,N_9748,N_9673);
and U9914 (N_9914,N_9783,N_9668);
or U9915 (N_9915,N_9701,N_9765);
nor U9916 (N_9916,N_9634,N_9779);
nor U9917 (N_9917,N_9788,N_9734);
and U9918 (N_9918,N_9738,N_9719);
or U9919 (N_9919,N_9782,N_9765);
xor U9920 (N_9920,N_9657,N_9752);
or U9921 (N_9921,N_9612,N_9723);
nor U9922 (N_9922,N_9664,N_9726);
xnor U9923 (N_9923,N_9638,N_9761);
nor U9924 (N_9924,N_9755,N_9784);
xnor U9925 (N_9925,N_9695,N_9715);
nor U9926 (N_9926,N_9799,N_9616);
and U9927 (N_9927,N_9703,N_9676);
or U9928 (N_9928,N_9797,N_9705);
nand U9929 (N_9929,N_9714,N_9783);
nand U9930 (N_9930,N_9670,N_9796);
and U9931 (N_9931,N_9655,N_9772);
and U9932 (N_9932,N_9673,N_9749);
xor U9933 (N_9933,N_9692,N_9735);
xnor U9934 (N_9934,N_9685,N_9782);
xor U9935 (N_9935,N_9601,N_9761);
and U9936 (N_9936,N_9741,N_9784);
nor U9937 (N_9937,N_9735,N_9637);
and U9938 (N_9938,N_9721,N_9629);
xor U9939 (N_9939,N_9714,N_9650);
nor U9940 (N_9940,N_9692,N_9600);
xor U9941 (N_9941,N_9623,N_9619);
and U9942 (N_9942,N_9753,N_9715);
xnor U9943 (N_9943,N_9612,N_9675);
xor U9944 (N_9944,N_9705,N_9752);
or U9945 (N_9945,N_9669,N_9775);
or U9946 (N_9946,N_9697,N_9728);
nor U9947 (N_9947,N_9677,N_9769);
nor U9948 (N_9948,N_9643,N_9632);
and U9949 (N_9949,N_9642,N_9617);
and U9950 (N_9950,N_9742,N_9738);
or U9951 (N_9951,N_9725,N_9732);
xor U9952 (N_9952,N_9772,N_9759);
and U9953 (N_9953,N_9663,N_9688);
nor U9954 (N_9954,N_9616,N_9627);
nand U9955 (N_9955,N_9770,N_9722);
nand U9956 (N_9956,N_9754,N_9722);
nand U9957 (N_9957,N_9744,N_9760);
and U9958 (N_9958,N_9780,N_9694);
nor U9959 (N_9959,N_9635,N_9716);
nand U9960 (N_9960,N_9749,N_9645);
nand U9961 (N_9961,N_9765,N_9746);
nand U9962 (N_9962,N_9614,N_9751);
nand U9963 (N_9963,N_9609,N_9670);
nor U9964 (N_9964,N_9636,N_9726);
xnor U9965 (N_9965,N_9724,N_9766);
and U9966 (N_9966,N_9608,N_9683);
and U9967 (N_9967,N_9727,N_9626);
xor U9968 (N_9968,N_9729,N_9760);
or U9969 (N_9969,N_9765,N_9757);
xor U9970 (N_9970,N_9659,N_9658);
nand U9971 (N_9971,N_9671,N_9610);
xor U9972 (N_9972,N_9623,N_9728);
nand U9973 (N_9973,N_9707,N_9699);
or U9974 (N_9974,N_9644,N_9774);
or U9975 (N_9975,N_9643,N_9624);
xnor U9976 (N_9976,N_9749,N_9649);
or U9977 (N_9977,N_9751,N_9686);
xnor U9978 (N_9978,N_9612,N_9737);
nand U9979 (N_9979,N_9619,N_9667);
or U9980 (N_9980,N_9725,N_9737);
nor U9981 (N_9981,N_9709,N_9712);
and U9982 (N_9982,N_9653,N_9610);
or U9983 (N_9983,N_9675,N_9710);
nand U9984 (N_9984,N_9659,N_9776);
and U9985 (N_9985,N_9684,N_9788);
and U9986 (N_9986,N_9602,N_9749);
and U9987 (N_9987,N_9638,N_9620);
nand U9988 (N_9988,N_9638,N_9696);
nand U9989 (N_9989,N_9757,N_9706);
and U9990 (N_9990,N_9668,N_9638);
xnor U9991 (N_9991,N_9757,N_9728);
nor U9992 (N_9992,N_9669,N_9734);
xor U9993 (N_9993,N_9773,N_9726);
or U9994 (N_9994,N_9704,N_9758);
nor U9995 (N_9995,N_9642,N_9637);
nor U9996 (N_9996,N_9682,N_9601);
or U9997 (N_9997,N_9722,N_9641);
or U9998 (N_9998,N_9705,N_9612);
or U9999 (N_9999,N_9643,N_9705);
xnor U10000 (N_10000,N_9971,N_9962);
nor U10001 (N_10001,N_9934,N_9931);
nand U10002 (N_10002,N_9841,N_9875);
or U10003 (N_10003,N_9929,N_9982);
nand U10004 (N_10004,N_9944,N_9958);
nor U10005 (N_10005,N_9967,N_9925);
and U10006 (N_10006,N_9866,N_9919);
or U10007 (N_10007,N_9988,N_9899);
nor U10008 (N_10008,N_9935,N_9990);
xor U10009 (N_10009,N_9815,N_9942);
xnor U10010 (N_10010,N_9861,N_9822);
or U10011 (N_10011,N_9854,N_9953);
nand U10012 (N_10012,N_9821,N_9945);
and U10013 (N_10013,N_9874,N_9985);
or U10014 (N_10014,N_9845,N_9909);
and U10015 (N_10015,N_9825,N_9957);
nor U10016 (N_10016,N_9829,N_9817);
nand U10017 (N_10017,N_9946,N_9968);
nor U10018 (N_10018,N_9921,N_9824);
xnor U10019 (N_10019,N_9893,N_9905);
or U10020 (N_10020,N_9923,N_9897);
or U10021 (N_10021,N_9871,N_9812);
nor U10022 (N_10022,N_9873,N_9926);
nor U10023 (N_10023,N_9865,N_9890);
nand U10024 (N_10024,N_9853,N_9917);
nand U10025 (N_10025,N_9974,N_9859);
or U10026 (N_10026,N_9963,N_9870);
or U10027 (N_10027,N_9930,N_9912);
nand U10028 (N_10028,N_9947,N_9885);
and U10029 (N_10029,N_9862,N_9832);
nor U10030 (N_10030,N_9833,N_9936);
nor U10031 (N_10031,N_9847,N_9973);
xnor U10032 (N_10032,N_9869,N_9916);
xnor U10033 (N_10033,N_9999,N_9902);
and U10034 (N_10034,N_9959,N_9867);
xor U10035 (N_10035,N_9801,N_9882);
nand U10036 (N_10036,N_9927,N_9907);
xnor U10037 (N_10037,N_9978,N_9852);
nor U10038 (N_10038,N_9810,N_9880);
and U10039 (N_10039,N_9881,N_9955);
or U10040 (N_10040,N_9964,N_9920);
and U10041 (N_10041,N_9995,N_9858);
nand U10042 (N_10042,N_9922,N_9911);
or U10043 (N_10043,N_9928,N_9887);
and U10044 (N_10044,N_9932,N_9992);
and U10045 (N_10045,N_9969,N_9949);
or U10046 (N_10046,N_9918,N_9804);
nand U10047 (N_10047,N_9828,N_9908);
and U10048 (N_10048,N_9996,N_9965);
xnor U10049 (N_10049,N_9901,N_9888);
or U10050 (N_10050,N_9831,N_9826);
nand U10051 (N_10051,N_9997,N_9864);
or U10052 (N_10052,N_9950,N_9876);
xor U10053 (N_10053,N_9814,N_9809);
xnor U10054 (N_10054,N_9842,N_9802);
nand U10055 (N_10055,N_9898,N_9910);
nor U10056 (N_10056,N_9807,N_9894);
xor U10057 (N_10057,N_9966,N_9933);
and U10058 (N_10058,N_9857,N_9954);
nor U10059 (N_10059,N_9986,N_9889);
or U10060 (N_10060,N_9983,N_9850);
and U10061 (N_10061,N_9848,N_9872);
nor U10062 (N_10062,N_9837,N_9913);
xor U10063 (N_10063,N_9903,N_9904);
nor U10064 (N_10064,N_9972,N_9827);
and U10065 (N_10065,N_9951,N_9886);
and U10066 (N_10066,N_9879,N_9977);
nor U10067 (N_10067,N_9851,N_9868);
nand U10068 (N_10068,N_9993,N_9840);
nor U10069 (N_10069,N_9943,N_9820);
and U10070 (N_10070,N_9856,N_9844);
nand U10071 (N_10071,N_9952,N_9948);
and U10072 (N_10072,N_9924,N_9830);
nor U10073 (N_10073,N_9994,N_9883);
xor U10074 (N_10074,N_9823,N_9998);
or U10075 (N_10075,N_9991,N_9940);
and U10076 (N_10076,N_9849,N_9813);
nand U10077 (N_10077,N_9860,N_9895);
or U10078 (N_10078,N_9980,N_9855);
or U10079 (N_10079,N_9884,N_9878);
or U10080 (N_10080,N_9839,N_9987);
and U10081 (N_10081,N_9984,N_9818);
xnor U10082 (N_10082,N_9976,N_9960);
and U10083 (N_10083,N_9938,N_9835);
nor U10084 (N_10084,N_9819,N_9805);
nand U10085 (N_10085,N_9808,N_9979);
and U10086 (N_10086,N_9811,N_9836);
and U10087 (N_10087,N_9896,N_9906);
xor U10088 (N_10088,N_9975,N_9834);
xor U10089 (N_10089,N_9800,N_9863);
nand U10090 (N_10090,N_9941,N_9900);
or U10091 (N_10091,N_9877,N_9989);
nor U10092 (N_10092,N_9803,N_9937);
nand U10093 (N_10093,N_9846,N_9981);
nand U10094 (N_10094,N_9806,N_9970);
nor U10095 (N_10095,N_9961,N_9892);
nor U10096 (N_10096,N_9914,N_9915);
xnor U10097 (N_10097,N_9939,N_9838);
nor U10098 (N_10098,N_9816,N_9843);
and U10099 (N_10099,N_9891,N_9956);
and U10100 (N_10100,N_9806,N_9908);
or U10101 (N_10101,N_9977,N_9856);
or U10102 (N_10102,N_9843,N_9849);
and U10103 (N_10103,N_9940,N_9892);
xor U10104 (N_10104,N_9913,N_9876);
nor U10105 (N_10105,N_9843,N_9886);
nand U10106 (N_10106,N_9889,N_9905);
nor U10107 (N_10107,N_9967,N_9964);
xor U10108 (N_10108,N_9900,N_9911);
nor U10109 (N_10109,N_9938,N_9992);
nand U10110 (N_10110,N_9820,N_9893);
and U10111 (N_10111,N_9837,N_9889);
xor U10112 (N_10112,N_9940,N_9931);
and U10113 (N_10113,N_9895,N_9976);
xor U10114 (N_10114,N_9881,N_9832);
or U10115 (N_10115,N_9877,N_9966);
and U10116 (N_10116,N_9922,N_9875);
nand U10117 (N_10117,N_9866,N_9898);
or U10118 (N_10118,N_9822,N_9895);
and U10119 (N_10119,N_9884,N_9928);
and U10120 (N_10120,N_9828,N_9932);
and U10121 (N_10121,N_9851,N_9845);
and U10122 (N_10122,N_9853,N_9873);
nand U10123 (N_10123,N_9950,N_9940);
nor U10124 (N_10124,N_9903,N_9936);
xor U10125 (N_10125,N_9998,N_9903);
xor U10126 (N_10126,N_9937,N_9925);
or U10127 (N_10127,N_9835,N_9968);
nor U10128 (N_10128,N_9933,N_9965);
nand U10129 (N_10129,N_9894,N_9947);
and U10130 (N_10130,N_9885,N_9879);
xnor U10131 (N_10131,N_9888,N_9991);
nand U10132 (N_10132,N_9965,N_9872);
and U10133 (N_10133,N_9851,N_9908);
xor U10134 (N_10134,N_9828,N_9991);
and U10135 (N_10135,N_9817,N_9871);
nor U10136 (N_10136,N_9960,N_9912);
nand U10137 (N_10137,N_9938,N_9920);
xor U10138 (N_10138,N_9956,N_9933);
or U10139 (N_10139,N_9834,N_9813);
nand U10140 (N_10140,N_9916,N_9970);
or U10141 (N_10141,N_9975,N_9880);
xor U10142 (N_10142,N_9824,N_9965);
xnor U10143 (N_10143,N_9806,N_9977);
or U10144 (N_10144,N_9886,N_9945);
xor U10145 (N_10145,N_9931,N_9936);
xnor U10146 (N_10146,N_9929,N_9875);
xnor U10147 (N_10147,N_9957,N_9916);
nand U10148 (N_10148,N_9935,N_9923);
or U10149 (N_10149,N_9910,N_9949);
xnor U10150 (N_10150,N_9901,N_9985);
nor U10151 (N_10151,N_9833,N_9932);
and U10152 (N_10152,N_9857,N_9925);
xor U10153 (N_10153,N_9820,N_9901);
nand U10154 (N_10154,N_9923,N_9904);
or U10155 (N_10155,N_9861,N_9838);
or U10156 (N_10156,N_9969,N_9970);
nand U10157 (N_10157,N_9819,N_9842);
nor U10158 (N_10158,N_9822,N_9814);
and U10159 (N_10159,N_9964,N_9902);
nor U10160 (N_10160,N_9853,N_9988);
and U10161 (N_10161,N_9949,N_9894);
and U10162 (N_10162,N_9980,N_9954);
and U10163 (N_10163,N_9837,N_9848);
nor U10164 (N_10164,N_9869,N_9989);
xnor U10165 (N_10165,N_9936,N_9847);
or U10166 (N_10166,N_9870,N_9948);
or U10167 (N_10167,N_9972,N_9950);
nor U10168 (N_10168,N_9818,N_9865);
nor U10169 (N_10169,N_9827,N_9873);
nand U10170 (N_10170,N_9813,N_9995);
nand U10171 (N_10171,N_9983,N_9936);
or U10172 (N_10172,N_9950,N_9860);
xnor U10173 (N_10173,N_9837,N_9959);
xnor U10174 (N_10174,N_9914,N_9873);
nand U10175 (N_10175,N_9929,N_9817);
nand U10176 (N_10176,N_9927,N_9987);
and U10177 (N_10177,N_9888,N_9935);
nand U10178 (N_10178,N_9937,N_9946);
and U10179 (N_10179,N_9827,N_9942);
and U10180 (N_10180,N_9820,N_9926);
or U10181 (N_10181,N_9922,N_9823);
or U10182 (N_10182,N_9890,N_9953);
xor U10183 (N_10183,N_9949,N_9919);
xnor U10184 (N_10184,N_9984,N_9856);
nor U10185 (N_10185,N_9913,N_9882);
or U10186 (N_10186,N_9811,N_9990);
nor U10187 (N_10187,N_9838,N_9948);
or U10188 (N_10188,N_9993,N_9958);
xor U10189 (N_10189,N_9800,N_9936);
or U10190 (N_10190,N_9838,N_9932);
and U10191 (N_10191,N_9994,N_9898);
and U10192 (N_10192,N_9938,N_9907);
or U10193 (N_10193,N_9919,N_9819);
xor U10194 (N_10194,N_9863,N_9830);
xnor U10195 (N_10195,N_9905,N_9930);
xnor U10196 (N_10196,N_9957,N_9936);
and U10197 (N_10197,N_9800,N_9914);
nand U10198 (N_10198,N_9971,N_9879);
xnor U10199 (N_10199,N_9941,N_9901);
nand U10200 (N_10200,N_10145,N_10004);
or U10201 (N_10201,N_10131,N_10022);
nand U10202 (N_10202,N_10067,N_10073);
xnor U10203 (N_10203,N_10006,N_10020);
or U10204 (N_10204,N_10116,N_10138);
nand U10205 (N_10205,N_10181,N_10052);
nor U10206 (N_10206,N_10146,N_10109);
and U10207 (N_10207,N_10009,N_10064);
xnor U10208 (N_10208,N_10185,N_10007);
or U10209 (N_10209,N_10005,N_10158);
nand U10210 (N_10210,N_10169,N_10096);
or U10211 (N_10211,N_10032,N_10072);
nor U10212 (N_10212,N_10081,N_10175);
and U10213 (N_10213,N_10115,N_10031);
nand U10214 (N_10214,N_10055,N_10193);
xnor U10215 (N_10215,N_10154,N_10156);
nand U10216 (N_10216,N_10026,N_10039);
and U10217 (N_10217,N_10155,N_10104);
nor U10218 (N_10218,N_10177,N_10092);
or U10219 (N_10219,N_10088,N_10082);
nor U10220 (N_10220,N_10123,N_10120);
or U10221 (N_10221,N_10140,N_10013);
and U10222 (N_10222,N_10148,N_10179);
nor U10223 (N_10223,N_10170,N_10149);
nand U10224 (N_10224,N_10030,N_10141);
or U10225 (N_10225,N_10098,N_10172);
or U10226 (N_10226,N_10083,N_10037);
nor U10227 (N_10227,N_10184,N_10126);
nand U10228 (N_10228,N_10113,N_10074);
or U10229 (N_10229,N_10017,N_10183);
and U10230 (N_10230,N_10065,N_10134);
nand U10231 (N_10231,N_10060,N_10047);
xor U10232 (N_10232,N_10122,N_10010);
xor U10233 (N_10233,N_10014,N_10199);
xor U10234 (N_10234,N_10024,N_10135);
and U10235 (N_10235,N_10105,N_10080);
nand U10236 (N_10236,N_10130,N_10164);
and U10237 (N_10237,N_10062,N_10027);
nand U10238 (N_10238,N_10044,N_10068);
nand U10239 (N_10239,N_10132,N_10159);
nand U10240 (N_10240,N_10054,N_10069);
xor U10241 (N_10241,N_10050,N_10076);
nand U10242 (N_10242,N_10127,N_10021);
nor U10243 (N_10243,N_10114,N_10150);
or U10244 (N_10244,N_10139,N_10023);
xor U10245 (N_10245,N_10090,N_10157);
nor U10246 (N_10246,N_10153,N_10182);
and U10247 (N_10247,N_10119,N_10110);
or U10248 (N_10248,N_10129,N_10108);
or U10249 (N_10249,N_10051,N_10056);
and U10250 (N_10250,N_10042,N_10118);
nand U10251 (N_10251,N_10136,N_10049);
and U10252 (N_10252,N_10143,N_10176);
nand U10253 (N_10253,N_10086,N_10034);
or U10254 (N_10254,N_10035,N_10171);
or U10255 (N_10255,N_10059,N_10137);
and U10256 (N_10256,N_10058,N_10198);
nor U10257 (N_10257,N_10187,N_10189);
xnor U10258 (N_10258,N_10011,N_10190);
or U10259 (N_10259,N_10028,N_10097);
and U10260 (N_10260,N_10008,N_10087);
nor U10261 (N_10261,N_10029,N_10012);
or U10262 (N_10262,N_10071,N_10016);
and U10263 (N_10263,N_10048,N_10040);
nor U10264 (N_10264,N_10038,N_10142);
or U10265 (N_10265,N_10151,N_10002);
nand U10266 (N_10266,N_10188,N_10018);
nand U10267 (N_10267,N_10043,N_10085);
nor U10268 (N_10268,N_10195,N_10101);
xor U10269 (N_10269,N_10173,N_10124);
and U10270 (N_10270,N_10194,N_10168);
xor U10271 (N_10271,N_10089,N_10019);
nor U10272 (N_10272,N_10041,N_10077);
or U10273 (N_10273,N_10102,N_10152);
xnor U10274 (N_10274,N_10166,N_10015);
xnor U10275 (N_10275,N_10186,N_10165);
nor U10276 (N_10276,N_10066,N_10001);
and U10277 (N_10277,N_10084,N_10111);
or U10278 (N_10278,N_10161,N_10107);
xor U10279 (N_10279,N_10178,N_10112);
xor U10280 (N_10280,N_10128,N_10162);
nor U10281 (N_10281,N_10079,N_10003);
and U10282 (N_10282,N_10075,N_10197);
nand U10283 (N_10283,N_10025,N_10045);
xor U10284 (N_10284,N_10000,N_10046);
nand U10285 (N_10285,N_10036,N_10133);
and U10286 (N_10286,N_10103,N_10091);
and U10287 (N_10287,N_10094,N_10078);
nand U10288 (N_10288,N_10061,N_10093);
nand U10289 (N_10289,N_10192,N_10163);
nor U10290 (N_10290,N_10106,N_10144);
xnor U10291 (N_10291,N_10167,N_10147);
nand U10292 (N_10292,N_10100,N_10174);
or U10293 (N_10293,N_10063,N_10053);
and U10294 (N_10294,N_10125,N_10099);
xnor U10295 (N_10295,N_10121,N_10033);
nand U10296 (N_10296,N_10070,N_10160);
nand U10297 (N_10297,N_10117,N_10180);
xnor U10298 (N_10298,N_10196,N_10095);
or U10299 (N_10299,N_10057,N_10191);
or U10300 (N_10300,N_10036,N_10002);
and U10301 (N_10301,N_10044,N_10031);
and U10302 (N_10302,N_10010,N_10150);
or U10303 (N_10303,N_10064,N_10110);
xnor U10304 (N_10304,N_10047,N_10142);
and U10305 (N_10305,N_10028,N_10136);
or U10306 (N_10306,N_10011,N_10166);
nor U10307 (N_10307,N_10003,N_10034);
nor U10308 (N_10308,N_10019,N_10003);
xnor U10309 (N_10309,N_10149,N_10038);
nand U10310 (N_10310,N_10048,N_10150);
nor U10311 (N_10311,N_10092,N_10014);
nand U10312 (N_10312,N_10085,N_10198);
nand U10313 (N_10313,N_10040,N_10036);
or U10314 (N_10314,N_10142,N_10126);
and U10315 (N_10315,N_10149,N_10191);
and U10316 (N_10316,N_10119,N_10050);
and U10317 (N_10317,N_10177,N_10157);
and U10318 (N_10318,N_10010,N_10025);
nand U10319 (N_10319,N_10042,N_10125);
and U10320 (N_10320,N_10163,N_10195);
nand U10321 (N_10321,N_10083,N_10124);
nor U10322 (N_10322,N_10129,N_10174);
nand U10323 (N_10323,N_10122,N_10194);
and U10324 (N_10324,N_10131,N_10108);
nand U10325 (N_10325,N_10150,N_10127);
or U10326 (N_10326,N_10066,N_10043);
or U10327 (N_10327,N_10033,N_10050);
xor U10328 (N_10328,N_10004,N_10047);
or U10329 (N_10329,N_10047,N_10090);
and U10330 (N_10330,N_10166,N_10190);
nor U10331 (N_10331,N_10085,N_10014);
and U10332 (N_10332,N_10160,N_10059);
and U10333 (N_10333,N_10199,N_10192);
nand U10334 (N_10334,N_10124,N_10194);
or U10335 (N_10335,N_10034,N_10072);
nand U10336 (N_10336,N_10151,N_10078);
xnor U10337 (N_10337,N_10082,N_10178);
nand U10338 (N_10338,N_10069,N_10049);
xor U10339 (N_10339,N_10003,N_10188);
nand U10340 (N_10340,N_10135,N_10154);
nand U10341 (N_10341,N_10128,N_10072);
xnor U10342 (N_10342,N_10052,N_10024);
and U10343 (N_10343,N_10032,N_10082);
nand U10344 (N_10344,N_10196,N_10182);
xor U10345 (N_10345,N_10090,N_10031);
xor U10346 (N_10346,N_10127,N_10044);
nor U10347 (N_10347,N_10025,N_10154);
nand U10348 (N_10348,N_10166,N_10098);
or U10349 (N_10349,N_10019,N_10027);
or U10350 (N_10350,N_10182,N_10174);
nor U10351 (N_10351,N_10107,N_10005);
nor U10352 (N_10352,N_10176,N_10066);
and U10353 (N_10353,N_10032,N_10141);
nand U10354 (N_10354,N_10199,N_10044);
nor U10355 (N_10355,N_10001,N_10178);
or U10356 (N_10356,N_10183,N_10180);
xnor U10357 (N_10357,N_10034,N_10020);
nand U10358 (N_10358,N_10198,N_10164);
or U10359 (N_10359,N_10008,N_10078);
xor U10360 (N_10360,N_10074,N_10015);
and U10361 (N_10361,N_10171,N_10198);
nand U10362 (N_10362,N_10052,N_10065);
and U10363 (N_10363,N_10025,N_10112);
nor U10364 (N_10364,N_10059,N_10023);
xor U10365 (N_10365,N_10194,N_10095);
nand U10366 (N_10366,N_10143,N_10171);
nor U10367 (N_10367,N_10058,N_10031);
nand U10368 (N_10368,N_10010,N_10090);
and U10369 (N_10369,N_10015,N_10168);
and U10370 (N_10370,N_10020,N_10100);
xor U10371 (N_10371,N_10043,N_10186);
and U10372 (N_10372,N_10197,N_10146);
nor U10373 (N_10373,N_10153,N_10107);
nor U10374 (N_10374,N_10187,N_10118);
or U10375 (N_10375,N_10196,N_10104);
nor U10376 (N_10376,N_10181,N_10145);
and U10377 (N_10377,N_10092,N_10015);
xor U10378 (N_10378,N_10189,N_10149);
xnor U10379 (N_10379,N_10053,N_10148);
or U10380 (N_10380,N_10145,N_10057);
xnor U10381 (N_10381,N_10136,N_10011);
nor U10382 (N_10382,N_10033,N_10088);
xor U10383 (N_10383,N_10073,N_10093);
xnor U10384 (N_10384,N_10063,N_10177);
and U10385 (N_10385,N_10071,N_10026);
nor U10386 (N_10386,N_10068,N_10142);
nand U10387 (N_10387,N_10077,N_10155);
nand U10388 (N_10388,N_10197,N_10024);
nand U10389 (N_10389,N_10120,N_10039);
xnor U10390 (N_10390,N_10032,N_10010);
nand U10391 (N_10391,N_10160,N_10164);
xor U10392 (N_10392,N_10145,N_10165);
and U10393 (N_10393,N_10134,N_10076);
xor U10394 (N_10394,N_10036,N_10154);
xnor U10395 (N_10395,N_10156,N_10043);
xnor U10396 (N_10396,N_10188,N_10011);
and U10397 (N_10397,N_10036,N_10018);
or U10398 (N_10398,N_10077,N_10094);
and U10399 (N_10399,N_10134,N_10097);
or U10400 (N_10400,N_10322,N_10394);
or U10401 (N_10401,N_10396,N_10341);
and U10402 (N_10402,N_10287,N_10200);
and U10403 (N_10403,N_10211,N_10225);
or U10404 (N_10404,N_10397,N_10326);
and U10405 (N_10405,N_10398,N_10345);
or U10406 (N_10406,N_10390,N_10228);
xnor U10407 (N_10407,N_10284,N_10314);
nor U10408 (N_10408,N_10353,N_10253);
xor U10409 (N_10409,N_10378,N_10386);
or U10410 (N_10410,N_10221,N_10309);
xor U10411 (N_10411,N_10291,N_10273);
and U10412 (N_10412,N_10364,N_10327);
xnor U10413 (N_10413,N_10348,N_10382);
nor U10414 (N_10414,N_10389,N_10263);
nand U10415 (N_10415,N_10380,N_10393);
nor U10416 (N_10416,N_10363,N_10204);
or U10417 (N_10417,N_10395,N_10366);
nor U10418 (N_10418,N_10301,N_10346);
nor U10419 (N_10419,N_10313,N_10274);
nor U10420 (N_10420,N_10238,N_10245);
or U10421 (N_10421,N_10249,N_10283);
nor U10422 (N_10422,N_10234,N_10320);
xor U10423 (N_10423,N_10205,N_10239);
or U10424 (N_10424,N_10206,N_10236);
and U10425 (N_10425,N_10377,N_10336);
nor U10426 (N_10426,N_10329,N_10367);
and U10427 (N_10427,N_10271,N_10357);
xnor U10428 (N_10428,N_10210,N_10347);
and U10429 (N_10429,N_10246,N_10230);
nor U10430 (N_10430,N_10351,N_10276);
xnor U10431 (N_10431,N_10269,N_10317);
and U10432 (N_10432,N_10244,N_10312);
and U10433 (N_10433,N_10222,N_10227);
or U10434 (N_10434,N_10358,N_10290);
or U10435 (N_10435,N_10342,N_10265);
nand U10436 (N_10436,N_10279,N_10354);
xor U10437 (N_10437,N_10315,N_10224);
xnor U10438 (N_10438,N_10201,N_10330);
xnor U10439 (N_10439,N_10350,N_10392);
nor U10440 (N_10440,N_10250,N_10267);
xor U10441 (N_10441,N_10212,N_10337);
nor U10442 (N_10442,N_10262,N_10310);
and U10443 (N_10443,N_10302,N_10308);
or U10444 (N_10444,N_10241,N_10359);
and U10445 (N_10445,N_10334,N_10275);
nand U10446 (N_10446,N_10305,N_10349);
nor U10447 (N_10447,N_10281,N_10272);
nand U10448 (N_10448,N_10338,N_10376);
nor U10449 (N_10449,N_10307,N_10261);
and U10450 (N_10450,N_10370,N_10369);
nand U10451 (N_10451,N_10237,N_10384);
nand U10452 (N_10452,N_10203,N_10332);
nand U10453 (N_10453,N_10375,N_10372);
xnor U10454 (N_10454,N_10352,N_10216);
or U10455 (N_10455,N_10311,N_10259);
nor U10456 (N_10456,N_10202,N_10277);
nor U10457 (N_10457,N_10297,N_10217);
and U10458 (N_10458,N_10218,N_10242);
xor U10459 (N_10459,N_10318,N_10356);
nand U10460 (N_10460,N_10252,N_10233);
nor U10461 (N_10461,N_10232,N_10381);
xor U10462 (N_10462,N_10316,N_10243);
nor U10463 (N_10463,N_10325,N_10256);
or U10464 (N_10464,N_10240,N_10319);
xnor U10465 (N_10465,N_10391,N_10264);
xnor U10466 (N_10466,N_10304,N_10368);
nor U10467 (N_10467,N_10247,N_10298);
xnor U10468 (N_10468,N_10255,N_10254);
and U10469 (N_10469,N_10362,N_10388);
or U10470 (N_10470,N_10344,N_10379);
and U10471 (N_10471,N_10223,N_10248);
nor U10472 (N_10472,N_10299,N_10340);
xor U10473 (N_10473,N_10324,N_10303);
nand U10474 (N_10474,N_10278,N_10360);
or U10475 (N_10475,N_10226,N_10383);
xor U10476 (N_10476,N_10333,N_10335);
nor U10477 (N_10477,N_10339,N_10328);
nor U10478 (N_10478,N_10258,N_10220);
and U10479 (N_10479,N_10219,N_10300);
xor U10480 (N_10480,N_10293,N_10289);
nand U10481 (N_10481,N_10343,N_10282);
xor U10482 (N_10482,N_10355,N_10209);
nor U10483 (N_10483,N_10323,N_10280);
and U10484 (N_10484,N_10295,N_10286);
nor U10485 (N_10485,N_10387,N_10215);
or U10486 (N_10486,N_10294,N_10207);
or U10487 (N_10487,N_10361,N_10231);
nor U10488 (N_10488,N_10213,N_10399);
nand U10489 (N_10489,N_10365,N_10292);
xnor U10490 (N_10490,N_10285,N_10385);
or U10491 (N_10491,N_10296,N_10288);
or U10492 (N_10492,N_10208,N_10260);
xnor U10493 (N_10493,N_10229,N_10214);
and U10494 (N_10494,N_10251,N_10374);
or U10495 (N_10495,N_10266,N_10373);
xnor U10496 (N_10496,N_10321,N_10306);
and U10497 (N_10497,N_10235,N_10331);
or U10498 (N_10498,N_10257,N_10270);
xor U10499 (N_10499,N_10268,N_10371);
nor U10500 (N_10500,N_10355,N_10263);
and U10501 (N_10501,N_10253,N_10242);
nor U10502 (N_10502,N_10256,N_10263);
nor U10503 (N_10503,N_10274,N_10322);
nand U10504 (N_10504,N_10253,N_10222);
or U10505 (N_10505,N_10378,N_10290);
nand U10506 (N_10506,N_10343,N_10341);
nor U10507 (N_10507,N_10241,N_10360);
nor U10508 (N_10508,N_10210,N_10254);
nor U10509 (N_10509,N_10311,N_10301);
nor U10510 (N_10510,N_10384,N_10239);
nor U10511 (N_10511,N_10270,N_10231);
and U10512 (N_10512,N_10265,N_10219);
nor U10513 (N_10513,N_10317,N_10242);
and U10514 (N_10514,N_10366,N_10301);
nor U10515 (N_10515,N_10212,N_10211);
nor U10516 (N_10516,N_10254,N_10360);
and U10517 (N_10517,N_10388,N_10282);
nor U10518 (N_10518,N_10217,N_10357);
nor U10519 (N_10519,N_10257,N_10291);
nor U10520 (N_10520,N_10291,N_10254);
nand U10521 (N_10521,N_10325,N_10210);
and U10522 (N_10522,N_10347,N_10308);
xor U10523 (N_10523,N_10202,N_10313);
nor U10524 (N_10524,N_10371,N_10298);
and U10525 (N_10525,N_10333,N_10314);
xnor U10526 (N_10526,N_10262,N_10220);
nand U10527 (N_10527,N_10300,N_10353);
or U10528 (N_10528,N_10227,N_10287);
or U10529 (N_10529,N_10272,N_10260);
nor U10530 (N_10530,N_10375,N_10351);
and U10531 (N_10531,N_10342,N_10279);
xnor U10532 (N_10532,N_10274,N_10351);
and U10533 (N_10533,N_10362,N_10221);
nand U10534 (N_10534,N_10362,N_10208);
and U10535 (N_10535,N_10360,N_10376);
xnor U10536 (N_10536,N_10307,N_10315);
xnor U10537 (N_10537,N_10228,N_10216);
and U10538 (N_10538,N_10326,N_10209);
nor U10539 (N_10539,N_10324,N_10265);
xor U10540 (N_10540,N_10208,N_10221);
and U10541 (N_10541,N_10258,N_10302);
xor U10542 (N_10542,N_10397,N_10287);
or U10543 (N_10543,N_10273,N_10355);
and U10544 (N_10544,N_10371,N_10315);
nor U10545 (N_10545,N_10290,N_10314);
xor U10546 (N_10546,N_10302,N_10293);
nor U10547 (N_10547,N_10354,N_10332);
nand U10548 (N_10548,N_10279,N_10312);
and U10549 (N_10549,N_10203,N_10230);
xnor U10550 (N_10550,N_10279,N_10200);
nand U10551 (N_10551,N_10396,N_10397);
xor U10552 (N_10552,N_10235,N_10217);
and U10553 (N_10553,N_10398,N_10364);
or U10554 (N_10554,N_10333,N_10301);
nor U10555 (N_10555,N_10252,N_10341);
nand U10556 (N_10556,N_10303,N_10369);
nand U10557 (N_10557,N_10343,N_10248);
nand U10558 (N_10558,N_10370,N_10317);
and U10559 (N_10559,N_10390,N_10216);
nor U10560 (N_10560,N_10315,N_10250);
nand U10561 (N_10561,N_10358,N_10268);
nor U10562 (N_10562,N_10319,N_10368);
and U10563 (N_10563,N_10200,N_10213);
or U10564 (N_10564,N_10313,N_10311);
nand U10565 (N_10565,N_10314,N_10390);
or U10566 (N_10566,N_10328,N_10271);
xor U10567 (N_10567,N_10343,N_10328);
or U10568 (N_10568,N_10320,N_10344);
and U10569 (N_10569,N_10239,N_10307);
or U10570 (N_10570,N_10318,N_10250);
nand U10571 (N_10571,N_10220,N_10229);
and U10572 (N_10572,N_10290,N_10271);
or U10573 (N_10573,N_10375,N_10305);
or U10574 (N_10574,N_10300,N_10247);
and U10575 (N_10575,N_10327,N_10381);
nor U10576 (N_10576,N_10230,N_10365);
and U10577 (N_10577,N_10243,N_10330);
or U10578 (N_10578,N_10303,N_10351);
nand U10579 (N_10579,N_10237,N_10337);
or U10580 (N_10580,N_10373,N_10265);
and U10581 (N_10581,N_10235,N_10369);
and U10582 (N_10582,N_10308,N_10273);
nand U10583 (N_10583,N_10351,N_10314);
or U10584 (N_10584,N_10339,N_10308);
and U10585 (N_10585,N_10353,N_10352);
or U10586 (N_10586,N_10316,N_10248);
nor U10587 (N_10587,N_10229,N_10353);
nand U10588 (N_10588,N_10307,N_10255);
nor U10589 (N_10589,N_10310,N_10268);
xnor U10590 (N_10590,N_10398,N_10265);
xor U10591 (N_10591,N_10252,N_10293);
xor U10592 (N_10592,N_10311,N_10338);
nand U10593 (N_10593,N_10253,N_10236);
nor U10594 (N_10594,N_10278,N_10226);
xor U10595 (N_10595,N_10246,N_10285);
nor U10596 (N_10596,N_10293,N_10393);
and U10597 (N_10597,N_10221,N_10391);
xor U10598 (N_10598,N_10329,N_10219);
nor U10599 (N_10599,N_10287,N_10347);
or U10600 (N_10600,N_10419,N_10437);
nor U10601 (N_10601,N_10495,N_10445);
xor U10602 (N_10602,N_10539,N_10403);
or U10603 (N_10603,N_10448,N_10594);
nand U10604 (N_10604,N_10597,N_10505);
xnor U10605 (N_10605,N_10479,N_10477);
xnor U10606 (N_10606,N_10489,N_10475);
or U10607 (N_10607,N_10493,N_10410);
nor U10608 (N_10608,N_10460,N_10596);
or U10609 (N_10609,N_10428,N_10543);
xor U10610 (N_10610,N_10532,N_10402);
and U10611 (N_10611,N_10484,N_10440);
nor U10612 (N_10612,N_10449,N_10537);
or U10613 (N_10613,N_10506,N_10457);
and U10614 (N_10614,N_10455,N_10551);
and U10615 (N_10615,N_10525,N_10508);
and U10616 (N_10616,N_10500,N_10544);
or U10617 (N_10617,N_10527,N_10464);
nor U10618 (N_10618,N_10542,N_10408);
nand U10619 (N_10619,N_10462,N_10516);
nor U10620 (N_10620,N_10503,N_10514);
or U10621 (N_10621,N_10468,N_10404);
nor U10622 (N_10622,N_10487,N_10469);
or U10623 (N_10623,N_10576,N_10534);
nor U10624 (N_10624,N_10434,N_10549);
and U10625 (N_10625,N_10540,N_10577);
nand U10626 (N_10626,N_10444,N_10583);
xor U10627 (N_10627,N_10560,N_10423);
and U10628 (N_10628,N_10548,N_10558);
xnor U10629 (N_10629,N_10414,N_10461);
or U10630 (N_10630,N_10535,N_10530);
xnor U10631 (N_10631,N_10592,N_10492);
nor U10632 (N_10632,N_10523,N_10565);
xnor U10633 (N_10633,N_10411,N_10572);
nand U10634 (N_10634,N_10520,N_10555);
nand U10635 (N_10635,N_10578,N_10407);
xnor U10636 (N_10636,N_10453,N_10429);
nand U10637 (N_10637,N_10439,N_10424);
and U10638 (N_10638,N_10531,N_10526);
or U10639 (N_10639,N_10422,N_10485);
and U10640 (N_10640,N_10433,N_10454);
xor U10641 (N_10641,N_10405,N_10478);
xnor U10642 (N_10642,N_10401,N_10447);
nor U10643 (N_10643,N_10563,N_10470);
nor U10644 (N_10644,N_10467,N_10575);
nand U10645 (N_10645,N_10581,N_10427);
nand U10646 (N_10646,N_10426,N_10472);
nand U10647 (N_10647,N_10588,N_10546);
xnor U10648 (N_10648,N_10412,N_10502);
or U10649 (N_10649,N_10490,N_10463);
and U10650 (N_10650,N_10491,N_10498);
or U10651 (N_10651,N_10459,N_10599);
nor U10652 (N_10652,N_10512,N_10590);
and U10653 (N_10653,N_10519,N_10473);
or U10654 (N_10654,N_10415,N_10579);
xor U10655 (N_10655,N_10566,N_10584);
and U10656 (N_10656,N_10413,N_10483);
and U10657 (N_10657,N_10511,N_10561);
and U10658 (N_10658,N_10541,N_10436);
nand U10659 (N_10659,N_10458,N_10451);
and U10660 (N_10660,N_10421,N_10559);
xor U10661 (N_10661,N_10533,N_10450);
xor U10662 (N_10662,N_10417,N_10418);
nor U10663 (N_10663,N_10488,N_10513);
or U10664 (N_10664,N_10420,N_10510);
nand U10665 (N_10665,N_10480,N_10482);
nand U10666 (N_10666,N_10430,N_10443);
and U10667 (N_10667,N_10476,N_10589);
xnor U10668 (N_10668,N_10524,N_10598);
nor U10669 (N_10669,N_10538,N_10466);
and U10670 (N_10670,N_10554,N_10580);
and U10671 (N_10671,N_10501,N_10562);
nor U10672 (N_10672,N_10446,N_10518);
and U10673 (N_10673,N_10529,N_10552);
nor U10674 (N_10674,N_10441,N_10509);
xor U10675 (N_10675,N_10571,N_10573);
nand U10676 (N_10676,N_10587,N_10557);
or U10677 (N_10677,N_10582,N_10567);
or U10678 (N_10678,N_10496,N_10591);
or U10679 (N_10679,N_10586,N_10406);
and U10680 (N_10680,N_10585,N_10465);
xor U10681 (N_10681,N_10517,N_10547);
or U10682 (N_10682,N_10435,N_10452);
nand U10683 (N_10683,N_10550,N_10536);
or U10684 (N_10684,N_10494,N_10593);
nor U10685 (N_10685,N_10471,N_10416);
or U10686 (N_10686,N_10556,N_10522);
and U10687 (N_10687,N_10595,N_10570);
xor U10688 (N_10688,N_10521,N_10425);
xnor U10689 (N_10689,N_10474,N_10574);
nor U10690 (N_10690,N_10432,N_10409);
nand U10691 (N_10691,N_10456,N_10569);
nand U10692 (N_10692,N_10553,N_10481);
nand U10693 (N_10693,N_10438,N_10486);
nor U10694 (N_10694,N_10507,N_10431);
xnor U10695 (N_10695,N_10528,N_10499);
and U10696 (N_10696,N_10564,N_10504);
xor U10697 (N_10697,N_10400,N_10442);
and U10698 (N_10698,N_10545,N_10568);
nor U10699 (N_10699,N_10497,N_10515);
and U10700 (N_10700,N_10428,N_10425);
and U10701 (N_10701,N_10561,N_10431);
nand U10702 (N_10702,N_10532,N_10412);
xnor U10703 (N_10703,N_10489,N_10482);
and U10704 (N_10704,N_10499,N_10444);
nand U10705 (N_10705,N_10535,N_10571);
or U10706 (N_10706,N_10512,N_10594);
or U10707 (N_10707,N_10471,N_10572);
or U10708 (N_10708,N_10476,N_10433);
nor U10709 (N_10709,N_10416,N_10504);
and U10710 (N_10710,N_10412,N_10547);
nand U10711 (N_10711,N_10546,N_10564);
nand U10712 (N_10712,N_10489,N_10531);
and U10713 (N_10713,N_10553,N_10565);
nor U10714 (N_10714,N_10575,N_10557);
nor U10715 (N_10715,N_10573,N_10544);
or U10716 (N_10716,N_10461,N_10538);
nand U10717 (N_10717,N_10507,N_10576);
xor U10718 (N_10718,N_10419,N_10493);
nor U10719 (N_10719,N_10462,N_10518);
nor U10720 (N_10720,N_10576,N_10448);
xnor U10721 (N_10721,N_10588,N_10574);
nor U10722 (N_10722,N_10589,N_10415);
or U10723 (N_10723,N_10501,N_10486);
and U10724 (N_10724,N_10550,N_10449);
and U10725 (N_10725,N_10550,N_10599);
nor U10726 (N_10726,N_10423,N_10500);
and U10727 (N_10727,N_10557,N_10508);
nand U10728 (N_10728,N_10468,N_10521);
or U10729 (N_10729,N_10410,N_10439);
xnor U10730 (N_10730,N_10405,N_10569);
nor U10731 (N_10731,N_10544,N_10418);
xnor U10732 (N_10732,N_10581,N_10521);
xor U10733 (N_10733,N_10483,N_10479);
xor U10734 (N_10734,N_10492,N_10568);
or U10735 (N_10735,N_10549,N_10471);
nand U10736 (N_10736,N_10524,N_10427);
or U10737 (N_10737,N_10563,N_10459);
nor U10738 (N_10738,N_10572,N_10413);
nor U10739 (N_10739,N_10465,N_10410);
or U10740 (N_10740,N_10538,N_10567);
nand U10741 (N_10741,N_10473,N_10429);
nand U10742 (N_10742,N_10526,N_10478);
and U10743 (N_10743,N_10513,N_10440);
nor U10744 (N_10744,N_10593,N_10458);
nand U10745 (N_10745,N_10584,N_10494);
xor U10746 (N_10746,N_10591,N_10470);
xnor U10747 (N_10747,N_10553,N_10418);
xor U10748 (N_10748,N_10466,N_10421);
nor U10749 (N_10749,N_10481,N_10544);
xnor U10750 (N_10750,N_10535,N_10424);
nor U10751 (N_10751,N_10412,N_10446);
nor U10752 (N_10752,N_10489,N_10402);
and U10753 (N_10753,N_10441,N_10571);
nor U10754 (N_10754,N_10590,N_10406);
nand U10755 (N_10755,N_10537,N_10423);
or U10756 (N_10756,N_10561,N_10425);
and U10757 (N_10757,N_10514,N_10586);
xnor U10758 (N_10758,N_10570,N_10511);
nor U10759 (N_10759,N_10491,N_10594);
or U10760 (N_10760,N_10406,N_10417);
xnor U10761 (N_10761,N_10430,N_10489);
xnor U10762 (N_10762,N_10437,N_10482);
nor U10763 (N_10763,N_10547,N_10485);
nand U10764 (N_10764,N_10598,N_10549);
nor U10765 (N_10765,N_10507,N_10458);
or U10766 (N_10766,N_10414,N_10583);
xor U10767 (N_10767,N_10566,N_10434);
nor U10768 (N_10768,N_10526,N_10424);
or U10769 (N_10769,N_10424,N_10405);
or U10770 (N_10770,N_10590,N_10479);
xor U10771 (N_10771,N_10537,N_10531);
xor U10772 (N_10772,N_10576,N_10542);
nor U10773 (N_10773,N_10461,N_10453);
and U10774 (N_10774,N_10572,N_10567);
xnor U10775 (N_10775,N_10419,N_10455);
nor U10776 (N_10776,N_10519,N_10415);
nor U10777 (N_10777,N_10569,N_10517);
xor U10778 (N_10778,N_10443,N_10543);
or U10779 (N_10779,N_10501,N_10548);
or U10780 (N_10780,N_10497,N_10596);
xor U10781 (N_10781,N_10520,N_10519);
xor U10782 (N_10782,N_10419,N_10594);
nor U10783 (N_10783,N_10500,N_10415);
xnor U10784 (N_10784,N_10598,N_10466);
xor U10785 (N_10785,N_10449,N_10406);
nor U10786 (N_10786,N_10438,N_10460);
or U10787 (N_10787,N_10493,N_10425);
and U10788 (N_10788,N_10513,N_10567);
nand U10789 (N_10789,N_10477,N_10551);
and U10790 (N_10790,N_10518,N_10428);
nor U10791 (N_10791,N_10499,N_10517);
and U10792 (N_10792,N_10586,N_10530);
xnor U10793 (N_10793,N_10485,N_10421);
and U10794 (N_10794,N_10549,N_10520);
xor U10795 (N_10795,N_10440,N_10481);
nand U10796 (N_10796,N_10596,N_10416);
nor U10797 (N_10797,N_10487,N_10497);
and U10798 (N_10798,N_10525,N_10565);
and U10799 (N_10799,N_10404,N_10562);
and U10800 (N_10800,N_10759,N_10762);
nor U10801 (N_10801,N_10776,N_10714);
nand U10802 (N_10802,N_10634,N_10653);
and U10803 (N_10803,N_10683,N_10725);
nand U10804 (N_10804,N_10682,N_10620);
or U10805 (N_10805,N_10644,N_10732);
and U10806 (N_10806,N_10752,N_10718);
xor U10807 (N_10807,N_10754,N_10645);
nand U10808 (N_10808,N_10789,N_10758);
nand U10809 (N_10809,N_10618,N_10643);
or U10810 (N_10810,N_10747,N_10727);
and U10811 (N_10811,N_10771,N_10749);
and U10812 (N_10812,N_10631,N_10703);
and U10813 (N_10813,N_10724,N_10687);
nand U10814 (N_10814,N_10666,N_10605);
nor U10815 (N_10815,N_10709,N_10711);
or U10816 (N_10816,N_10716,N_10782);
and U10817 (N_10817,N_10673,N_10788);
xnor U10818 (N_10818,N_10681,N_10627);
and U10819 (N_10819,N_10744,N_10722);
or U10820 (N_10820,N_10674,N_10751);
nor U10821 (N_10821,N_10662,N_10773);
or U10822 (N_10822,N_10787,N_10700);
nor U10823 (N_10823,N_10690,N_10667);
nor U10824 (N_10824,N_10770,N_10632);
xnor U10825 (N_10825,N_10661,N_10704);
and U10826 (N_10826,N_10622,N_10604);
or U10827 (N_10827,N_10616,N_10783);
nand U10828 (N_10828,N_10742,N_10723);
nand U10829 (N_10829,N_10637,N_10708);
or U10830 (N_10830,N_10772,N_10701);
xnor U10831 (N_10831,N_10707,N_10774);
nand U10832 (N_10832,N_10623,N_10713);
or U10833 (N_10833,N_10646,N_10781);
nand U10834 (N_10834,N_10730,N_10729);
or U10835 (N_10835,N_10735,N_10615);
nand U10836 (N_10836,N_10763,N_10686);
and U10837 (N_10837,N_10785,N_10746);
or U10838 (N_10838,N_10670,N_10769);
and U10839 (N_10839,N_10733,N_10657);
or U10840 (N_10840,N_10710,N_10639);
nand U10841 (N_10841,N_10606,N_10678);
and U10842 (N_10842,N_10736,N_10706);
and U10843 (N_10843,N_10750,N_10790);
nand U10844 (N_10844,N_10755,N_10702);
nor U10845 (N_10845,N_10654,N_10617);
and U10846 (N_10846,N_10726,N_10717);
nand U10847 (N_10847,N_10797,N_10640);
nand U10848 (N_10848,N_10663,N_10794);
and U10849 (N_10849,N_10664,N_10760);
nor U10850 (N_10850,N_10695,N_10614);
xor U10851 (N_10851,N_10731,N_10669);
nor U10852 (N_10852,N_10638,N_10636);
and U10853 (N_10853,N_10607,N_10768);
nand U10854 (N_10854,N_10780,N_10625);
nand U10855 (N_10855,N_10680,N_10697);
or U10856 (N_10856,N_10734,N_10608);
and U10857 (N_10857,N_10737,N_10764);
nand U10858 (N_10858,N_10748,N_10688);
nor U10859 (N_10859,N_10675,N_10753);
and U10860 (N_10860,N_10660,N_10671);
nor U10861 (N_10861,N_10611,N_10791);
nand U10862 (N_10862,N_10610,N_10626);
nor U10863 (N_10863,N_10738,N_10635);
nor U10864 (N_10864,N_10628,N_10619);
and U10865 (N_10865,N_10629,N_10777);
xor U10866 (N_10866,N_10656,N_10792);
or U10867 (N_10867,N_10677,N_10658);
and U10868 (N_10868,N_10765,N_10798);
xnor U10869 (N_10869,N_10601,N_10728);
or U10870 (N_10870,N_10679,N_10712);
nand U10871 (N_10871,N_10757,N_10756);
xnor U10872 (N_10872,N_10786,N_10676);
and U10873 (N_10873,N_10766,N_10715);
xnor U10874 (N_10874,N_10633,N_10668);
and U10875 (N_10875,N_10796,N_10652);
nor U10876 (N_10876,N_10743,N_10696);
nor U10877 (N_10877,N_10659,N_10689);
nor U10878 (N_10878,N_10799,N_10705);
nor U10879 (N_10879,N_10795,N_10693);
nand U10880 (N_10880,N_10665,N_10613);
nor U10881 (N_10881,N_10603,N_10612);
or U10882 (N_10882,N_10624,N_10784);
or U10883 (N_10883,N_10698,N_10651);
and U10884 (N_10884,N_10694,N_10775);
nor U10885 (N_10885,N_10721,N_10699);
nand U10886 (N_10886,N_10685,N_10650);
nor U10887 (N_10887,N_10647,N_10655);
nand U10888 (N_10888,N_10630,N_10691);
and U10889 (N_10889,N_10741,N_10621);
or U10890 (N_10890,N_10609,N_10779);
nor U10891 (N_10891,N_10719,N_10642);
xor U10892 (N_10892,N_10648,N_10649);
and U10893 (N_10893,N_10761,N_10740);
nor U10894 (N_10894,N_10672,N_10745);
or U10895 (N_10895,N_10602,N_10641);
nor U10896 (N_10896,N_10684,N_10692);
and U10897 (N_10897,N_10720,N_10600);
xnor U10898 (N_10898,N_10778,N_10767);
xnor U10899 (N_10899,N_10793,N_10739);
nand U10900 (N_10900,N_10721,N_10683);
or U10901 (N_10901,N_10682,N_10692);
or U10902 (N_10902,N_10705,N_10695);
nor U10903 (N_10903,N_10694,N_10701);
and U10904 (N_10904,N_10661,N_10756);
nor U10905 (N_10905,N_10729,N_10696);
and U10906 (N_10906,N_10650,N_10623);
nor U10907 (N_10907,N_10704,N_10659);
or U10908 (N_10908,N_10734,N_10745);
nand U10909 (N_10909,N_10715,N_10695);
and U10910 (N_10910,N_10696,N_10651);
nor U10911 (N_10911,N_10706,N_10746);
or U10912 (N_10912,N_10703,N_10683);
nor U10913 (N_10913,N_10600,N_10645);
nor U10914 (N_10914,N_10721,N_10746);
xnor U10915 (N_10915,N_10684,N_10781);
or U10916 (N_10916,N_10635,N_10632);
and U10917 (N_10917,N_10753,N_10709);
xor U10918 (N_10918,N_10723,N_10666);
and U10919 (N_10919,N_10651,N_10747);
nor U10920 (N_10920,N_10755,N_10796);
or U10921 (N_10921,N_10603,N_10647);
and U10922 (N_10922,N_10789,N_10734);
nand U10923 (N_10923,N_10722,N_10632);
xnor U10924 (N_10924,N_10784,N_10728);
nand U10925 (N_10925,N_10746,N_10655);
or U10926 (N_10926,N_10687,N_10613);
and U10927 (N_10927,N_10619,N_10659);
or U10928 (N_10928,N_10618,N_10798);
nor U10929 (N_10929,N_10628,N_10693);
or U10930 (N_10930,N_10713,N_10665);
and U10931 (N_10931,N_10628,N_10685);
and U10932 (N_10932,N_10732,N_10716);
xor U10933 (N_10933,N_10782,N_10692);
or U10934 (N_10934,N_10759,N_10778);
and U10935 (N_10935,N_10786,N_10617);
or U10936 (N_10936,N_10685,N_10787);
xor U10937 (N_10937,N_10702,N_10741);
or U10938 (N_10938,N_10702,N_10678);
or U10939 (N_10939,N_10619,N_10714);
nor U10940 (N_10940,N_10772,N_10627);
nor U10941 (N_10941,N_10685,N_10765);
xor U10942 (N_10942,N_10774,N_10639);
nor U10943 (N_10943,N_10781,N_10668);
and U10944 (N_10944,N_10714,N_10783);
xor U10945 (N_10945,N_10654,N_10704);
and U10946 (N_10946,N_10666,N_10714);
nor U10947 (N_10947,N_10691,N_10713);
and U10948 (N_10948,N_10691,N_10711);
or U10949 (N_10949,N_10772,N_10787);
nor U10950 (N_10950,N_10745,N_10639);
xnor U10951 (N_10951,N_10771,N_10734);
xnor U10952 (N_10952,N_10645,N_10709);
nor U10953 (N_10953,N_10697,N_10690);
nor U10954 (N_10954,N_10623,N_10756);
nand U10955 (N_10955,N_10697,N_10674);
xor U10956 (N_10956,N_10617,N_10702);
nor U10957 (N_10957,N_10658,N_10637);
xnor U10958 (N_10958,N_10744,N_10697);
nand U10959 (N_10959,N_10667,N_10740);
nor U10960 (N_10960,N_10756,N_10753);
nor U10961 (N_10961,N_10602,N_10777);
and U10962 (N_10962,N_10769,N_10709);
and U10963 (N_10963,N_10685,N_10659);
nand U10964 (N_10964,N_10672,N_10702);
xor U10965 (N_10965,N_10665,N_10716);
or U10966 (N_10966,N_10768,N_10616);
nand U10967 (N_10967,N_10605,N_10786);
and U10968 (N_10968,N_10745,N_10612);
nor U10969 (N_10969,N_10620,N_10747);
nand U10970 (N_10970,N_10646,N_10757);
nand U10971 (N_10971,N_10666,N_10751);
or U10972 (N_10972,N_10757,N_10658);
and U10973 (N_10973,N_10630,N_10702);
nor U10974 (N_10974,N_10785,N_10618);
xnor U10975 (N_10975,N_10634,N_10666);
or U10976 (N_10976,N_10621,N_10701);
and U10977 (N_10977,N_10675,N_10775);
nor U10978 (N_10978,N_10686,N_10734);
or U10979 (N_10979,N_10606,N_10715);
and U10980 (N_10980,N_10797,N_10623);
xnor U10981 (N_10981,N_10650,N_10645);
and U10982 (N_10982,N_10670,N_10728);
nor U10983 (N_10983,N_10636,N_10734);
and U10984 (N_10984,N_10716,N_10713);
or U10985 (N_10985,N_10717,N_10654);
and U10986 (N_10986,N_10785,N_10651);
or U10987 (N_10987,N_10671,N_10631);
nand U10988 (N_10988,N_10632,N_10757);
and U10989 (N_10989,N_10636,N_10646);
xor U10990 (N_10990,N_10670,N_10727);
xnor U10991 (N_10991,N_10729,N_10673);
or U10992 (N_10992,N_10642,N_10671);
xnor U10993 (N_10993,N_10738,N_10615);
or U10994 (N_10994,N_10703,N_10685);
nor U10995 (N_10995,N_10698,N_10702);
or U10996 (N_10996,N_10603,N_10655);
nor U10997 (N_10997,N_10799,N_10630);
and U10998 (N_10998,N_10789,N_10663);
nand U10999 (N_10999,N_10692,N_10781);
or U11000 (N_11000,N_10869,N_10925);
and U11001 (N_11001,N_10996,N_10861);
nor U11002 (N_11002,N_10857,N_10949);
or U11003 (N_11003,N_10938,N_10962);
and U11004 (N_11004,N_10830,N_10875);
and U11005 (N_11005,N_10905,N_10918);
xor U11006 (N_11006,N_10853,N_10849);
and U11007 (N_11007,N_10812,N_10851);
nor U11008 (N_11008,N_10976,N_10865);
nand U11009 (N_11009,N_10921,N_10864);
and U11010 (N_11010,N_10872,N_10874);
nand U11011 (N_11011,N_10970,N_10951);
and U11012 (N_11012,N_10955,N_10889);
nand U11013 (N_11013,N_10840,N_10928);
or U11014 (N_11014,N_10901,N_10934);
and U11015 (N_11015,N_10994,N_10960);
nor U11016 (N_11016,N_10837,N_10937);
nor U11017 (N_11017,N_10866,N_10992);
or U11018 (N_11018,N_10913,N_10917);
nand U11019 (N_11019,N_10805,N_10900);
nor U11020 (N_11020,N_10977,N_10884);
nor U11021 (N_11021,N_10856,N_10859);
nor U11022 (N_11022,N_10825,N_10882);
nand U11023 (N_11023,N_10932,N_10969);
or U11024 (N_11024,N_10867,N_10898);
and U11025 (N_11025,N_10950,N_10893);
nand U11026 (N_11026,N_10959,N_10923);
nor U11027 (N_11027,N_10968,N_10904);
nand U11028 (N_11028,N_10891,N_10933);
xnor U11029 (N_11029,N_10852,N_10868);
xor U11030 (N_11030,N_10924,N_10886);
nand U11031 (N_11031,N_10873,N_10836);
xnor U11032 (N_11032,N_10802,N_10888);
or U11033 (N_11033,N_10834,N_10972);
xnor U11034 (N_11034,N_10974,N_10943);
and U11035 (N_11035,N_10847,N_10870);
and U11036 (N_11036,N_10820,N_10916);
nand U11037 (N_11037,N_10803,N_10824);
and U11038 (N_11038,N_10899,N_10926);
nand U11039 (N_11039,N_10848,N_10823);
nor U11040 (N_11040,N_10881,N_10871);
nor U11041 (N_11041,N_10858,N_10897);
nand U11042 (N_11042,N_10930,N_10843);
nand U11043 (N_11043,N_10966,N_10818);
nor U11044 (N_11044,N_10999,N_10844);
nand U11045 (N_11045,N_10984,N_10832);
nand U11046 (N_11046,N_10936,N_10841);
or U11047 (N_11047,N_10961,N_10952);
and U11048 (N_11048,N_10817,N_10997);
and U11049 (N_11049,N_10995,N_10815);
and U11050 (N_11050,N_10998,N_10915);
and U11051 (N_11051,N_10821,N_10816);
nor U11052 (N_11052,N_10947,N_10806);
nor U11053 (N_11053,N_10954,N_10981);
nor U11054 (N_11054,N_10819,N_10850);
nand U11055 (N_11055,N_10831,N_10914);
xor U11056 (N_11056,N_10929,N_10906);
nor U11057 (N_11057,N_10903,N_10983);
or U11058 (N_11058,N_10879,N_10944);
or U11059 (N_11059,N_10896,N_10880);
nor U11060 (N_11060,N_10854,N_10946);
and U11061 (N_11061,N_10978,N_10833);
nand U11062 (N_11062,N_10971,N_10911);
and U11063 (N_11063,N_10876,N_10839);
or U11064 (N_11064,N_10892,N_10967);
nor U11065 (N_11065,N_10842,N_10993);
xor U11066 (N_11066,N_10940,N_10982);
xor U11067 (N_11067,N_10883,N_10988);
nand U11068 (N_11068,N_10907,N_10885);
or U11069 (N_11069,N_10939,N_10878);
xnor U11070 (N_11070,N_10927,N_10807);
or U11071 (N_11071,N_10964,N_10801);
xor U11072 (N_11072,N_10942,N_10813);
nand U11073 (N_11073,N_10908,N_10826);
nor U11074 (N_11074,N_10987,N_10920);
nor U11075 (N_11075,N_10910,N_10835);
xnor U11076 (N_11076,N_10945,N_10931);
nor U11077 (N_11077,N_10845,N_10975);
nand U11078 (N_11078,N_10980,N_10846);
and U11079 (N_11079,N_10958,N_10935);
or U11080 (N_11080,N_10828,N_10811);
and U11081 (N_11081,N_10822,N_10827);
and U11082 (N_11082,N_10810,N_10894);
or U11083 (N_11083,N_10963,N_10838);
nand U11084 (N_11084,N_10922,N_10979);
nor U11085 (N_11085,N_10887,N_10829);
and U11086 (N_11086,N_10941,N_10953);
xnor U11087 (N_11087,N_10948,N_10877);
xor U11088 (N_11088,N_10814,N_10890);
xor U11089 (N_11089,N_10912,N_10990);
xor U11090 (N_11090,N_10991,N_10989);
or U11091 (N_11091,N_10800,N_10985);
nor U11092 (N_11092,N_10860,N_10862);
nand U11093 (N_11093,N_10863,N_10956);
xnor U11094 (N_11094,N_10855,N_10902);
or U11095 (N_11095,N_10986,N_10973);
and U11096 (N_11096,N_10957,N_10919);
and U11097 (N_11097,N_10895,N_10909);
nor U11098 (N_11098,N_10808,N_10804);
and U11099 (N_11099,N_10809,N_10965);
xnor U11100 (N_11100,N_10848,N_10961);
nor U11101 (N_11101,N_10885,N_10879);
xor U11102 (N_11102,N_10818,N_10804);
nand U11103 (N_11103,N_10814,N_10803);
xor U11104 (N_11104,N_10868,N_10826);
nand U11105 (N_11105,N_10848,N_10858);
xnor U11106 (N_11106,N_10911,N_10909);
or U11107 (N_11107,N_10961,N_10932);
and U11108 (N_11108,N_10879,N_10849);
nor U11109 (N_11109,N_10850,N_10824);
xor U11110 (N_11110,N_10967,N_10946);
xor U11111 (N_11111,N_10886,N_10887);
nand U11112 (N_11112,N_10891,N_10888);
or U11113 (N_11113,N_10947,N_10990);
nor U11114 (N_11114,N_10987,N_10873);
nand U11115 (N_11115,N_10992,N_10917);
nor U11116 (N_11116,N_10971,N_10939);
nor U11117 (N_11117,N_10831,N_10817);
nand U11118 (N_11118,N_10945,N_10940);
xor U11119 (N_11119,N_10933,N_10819);
and U11120 (N_11120,N_10840,N_10871);
and U11121 (N_11121,N_10857,N_10959);
xor U11122 (N_11122,N_10950,N_10963);
and U11123 (N_11123,N_10818,N_10891);
or U11124 (N_11124,N_10916,N_10808);
nand U11125 (N_11125,N_10958,N_10831);
nor U11126 (N_11126,N_10927,N_10965);
xnor U11127 (N_11127,N_10939,N_10934);
xor U11128 (N_11128,N_10919,N_10818);
or U11129 (N_11129,N_10948,N_10882);
nor U11130 (N_11130,N_10868,N_10978);
and U11131 (N_11131,N_10987,N_10967);
or U11132 (N_11132,N_10986,N_10828);
xor U11133 (N_11133,N_10940,N_10929);
nand U11134 (N_11134,N_10905,N_10916);
nor U11135 (N_11135,N_10833,N_10890);
nand U11136 (N_11136,N_10882,N_10935);
and U11137 (N_11137,N_10819,N_10821);
and U11138 (N_11138,N_10900,N_10862);
or U11139 (N_11139,N_10829,N_10872);
or U11140 (N_11140,N_10839,N_10919);
or U11141 (N_11141,N_10923,N_10958);
xor U11142 (N_11142,N_10849,N_10808);
nand U11143 (N_11143,N_10976,N_10943);
and U11144 (N_11144,N_10974,N_10843);
or U11145 (N_11145,N_10992,N_10865);
xor U11146 (N_11146,N_10843,N_10943);
and U11147 (N_11147,N_10839,N_10970);
xor U11148 (N_11148,N_10879,N_10953);
and U11149 (N_11149,N_10998,N_10986);
or U11150 (N_11150,N_10979,N_10842);
nor U11151 (N_11151,N_10902,N_10875);
nor U11152 (N_11152,N_10855,N_10920);
and U11153 (N_11153,N_10802,N_10930);
and U11154 (N_11154,N_10901,N_10930);
and U11155 (N_11155,N_10915,N_10804);
nor U11156 (N_11156,N_10893,N_10981);
nor U11157 (N_11157,N_10873,N_10977);
or U11158 (N_11158,N_10889,N_10929);
or U11159 (N_11159,N_10903,N_10976);
or U11160 (N_11160,N_10901,N_10913);
and U11161 (N_11161,N_10899,N_10937);
nor U11162 (N_11162,N_10873,N_10868);
or U11163 (N_11163,N_10988,N_10935);
nand U11164 (N_11164,N_10804,N_10914);
xnor U11165 (N_11165,N_10972,N_10992);
nor U11166 (N_11166,N_10950,N_10895);
or U11167 (N_11167,N_10937,N_10828);
and U11168 (N_11168,N_10827,N_10817);
nand U11169 (N_11169,N_10861,N_10807);
nand U11170 (N_11170,N_10979,N_10892);
nand U11171 (N_11171,N_10825,N_10868);
nor U11172 (N_11172,N_10826,N_10964);
nor U11173 (N_11173,N_10920,N_10883);
or U11174 (N_11174,N_10949,N_10877);
or U11175 (N_11175,N_10878,N_10926);
nor U11176 (N_11176,N_10963,N_10997);
xor U11177 (N_11177,N_10913,N_10937);
xor U11178 (N_11178,N_10944,N_10907);
or U11179 (N_11179,N_10986,N_10886);
xor U11180 (N_11180,N_10975,N_10860);
xnor U11181 (N_11181,N_10885,N_10966);
and U11182 (N_11182,N_10970,N_10858);
nand U11183 (N_11183,N_10973,N_10818);
xor U11184 (N_11184,N_10882,N_10872);
or U11185 (N_11185,N_10917,N_10994);
nor U11186 (N_11186,N_10936,N_10823);
nor U11187 (N_11187,N_10952,N_10908);
or U11188 (N_11188,N_10804,N_10962);
nand U11189 (N_11189,N_10800,N_10867);
nor U11190 (N_11190,N_10920,N_10884);
and U11191 (N_11191,N_10949,N_10972);
and U11192 (N_11192,N_10993,N_10853);
nand U11193 (N_11193,N_10976,N_10994);
nor U11194 (N_11194,N_10966,N_10809);
and U11195 (N_11195,N_10883,N_10801);
nor U11196 (N_11196,N_10919,N_10960);
xnor U11197 (N_11197,N_10887,N_10984);
nor U11198 (N_11198,N_10996,N_10926);
xnor U11199 (N_11199,N_10991,N_10935);
xor U11200 (N_11200,N_11052,N_11134);
xnor U11201 (N_11201,N_11161,N_11009);
nor U11202 (N_11202,N_11101,N_11124);
and U11203 (N_11203,N_11165,N_11006);
nand U11204 (N_11204,N_11064,N_11176);
and U11205 (N_11205,N_11028,N_11164);
and U11206 (N_11206,N_11104,N_11139);
nand U11207 (N_11207,N_11157,N_11199);
xnor U11208 (N_11208,N_11019,N_11093);
nor U11209 (N_11209,N_11098,N_11057);
xnor U11210 (N_11210,N_11041,N_11198);
and U11211 (N_11211,N_11092,N_11170);
or U11212 (N_11212,N_11062,N_11177);
nor U11213 (N_11213,N_11027,N_11070);
or U11214 (N_11214,N_11127,N_11130);
nand U11215 (N_11215,N_11071,N_11103);
xnor U11216 (N_11216,N_11003,N_11094);
or U11217 (N_11217,N_11194,N_11049);
and U11218 (N_11218,N_11081,N_11033);
or U11219 (N_11219,N_11079,N_11126);
nor U11220 (N_11220,N_11097,N_11043);
nor U11221 (N_11221,N_11158,N_11122);
xnor U11222 (N_11222,N_11020,N_11059);
nand U11223 (N_11223,N_11102,N_11036);
nor U11224 (N_11224,N_11100,N_11148);
nor U11225 (N_11225,N_11105,N_11016);
or U11226 (N_11226,N_11015,N_11132);
xnor U11227 (N_11227,N_11114,N_11083);
and U11228 (N_11228,N_11002,N_11011);
and U11229 (N_11229,N_11150,N_11060);
nor U11230 (N_11230,N_11187,N_11076);
or U11231 (N_11231,N_11146,N_11024);
and U11232 (N_11232,N_11125,N_11069);
and U11233 (N_11233,N_11107,N_11029);
nor U11234 (N_11234,N_11193,N_11090);
nor U11235 (N_11235,N_11075,N_11053);
nand U11236 (N_11236,N_11007,N_11018);
or U11237 (N_11237,N_11044,N_11188);
or U11238 (N_11238,N_11035,N_11182);
nand U11239 (N_11239,N_11032,N_11109);
nor U11240 (N_11240,N_11144,N_11121);
xnor U11241 (N_11241,N_11168,N_11038);
xnor U11242 (N_11242,N_11115,N_11112);
nor U11243 (N_11243,N_11023,N_11078);
or U11244 (N_11244,N_11026,N_11137);
xnor U11245 (N_11245,N_11159,N_11108);
nand U11246 (N_11246,N_11034,N_11117);
and U11247 (N_11247,N_11166,N_11012);
nand U11248 (N_11248,N_11197,N_11140);
or U11249 (N_11249,N_11185,N_11192);
nand U11250 (N_11250,N_11180,N_11095);
and U11251 (N_11251,N_11087,N_11088);
or U11252 (N_11252,N_11047,N_11152);
xnor U11253 (N_11253,N_11025,N_11084);
xnor U11254 (N_11254,N_11173,N_11174);
and U11255 (N_11255,N_11119,N_11138);
nand U11256 (N_11256,N_11040,N_11172);
nand U11257 (N_11257,N_11133,N_11195);
xor U11258 (N_11258,N_11054,N_11042);
and U11259 (N_11259,N_11067,N_11058);
nor U11260 (N_11260,N_11068,N_11111);
nor U11261 (N_11261,N_11149,N_11000);
nor U11262 (N_11262,N_11051,N_11056);
or U11263 (N_11263,N_11145,N_11129);
or U11264 (N_11264,N_11156,N_11116);
nand U11265 (N_11265,N_11143,N_11151);
xor U11266 (N_11266,N_11022,N_11106);
or U11267 (N_11267,N_11160,N_11037);
nand U11268 (N_11268,N_11089,N_11186);
nor U11269 (N_11269,N_11014,N_11030);
nor U11270 (N_11270,N_11162,N_11163);
and U11271 (N_11271,N_11021,N_11113);
and U11272 (N_11272,N_11013,N_11167);
nor U11273 (N_11273,N_11061,N_11120);
nand U11274 (N_11274,N_11055,N_11169);
nor U11275 (N_11275,N_11179,N_11017);
or U11276 (N_11276,N_11072,N_11189);
or U11277 (N_11277,N_11110,N_11183);
xnor U11278 (N_11278,N_11099,N_11171);
and U11279 (N_11279,N_11141,N_11031);
nor U11280 (N_11280,N_11001,N_11050);
and U11281 (N_11281,N_11153,N_11123);
and U11282 (N_11282,N_11048,N_11147);
nand U11283 (N_11283,N_11005,N_11080);
xnor U11284 (N_11284,N_11046,N_11155);
nor U11285 (N_11285,N_11190,N_11136);
nand U11286 (N_11286,N_11010,N_11039);
xor U11287 (N_11287,N_11096,N_11175);
or U11288 (N_11288,N_11074,N_11184);
nand U11289 (N_11289,N_11045,N_11086);
nand U11290 (N_11290,N_11154,N_11066);
nand U11291 (N_11291,N_11091,N_11142);
xor U11292 (N_11292,N_11131,N_11073);
xor U11293 (N_11293,N_11063,N_11135);
nand U11294 (N_11294,N_11181,N_11196);
nor U11295 (N_11295,N_11085,N_11118);
and U11296 (N_11296,N_11178,N_11191);
or U11297 (N_11297,N_11082,N_11004);
or U11298 (N_11298,N_11065,N_11077);
or U11299 (N_11299,N_11128,N_11008);
and U11300 (N_11300,N_11199,N_11098);
and U11301 (N_11301,N_11035,N_11015);
or U11302 (N_11302,N_11073,N_11082);
nand U11303 (N_11303,N_11127,N_11132);
and U11304 (N_11304,N_11109,N_11079);
nor U11305 (N_11305,N_11034,N_11042);
or U11306 (N_11306,N_11051,N_11134);
nand U11307 (N_11307,N_11021,N_11189);
xnor U11308 (N_11308,N_11047,N_11164);
nor U11309 (N_11309,N_11009,N_11084);
nand U11310 (N_11310,N_11144,N_11140);
nand U11311 (N_11311,N_11064,N_11011);
and U11312 (N_11312,N_11043,N_11191);
and U11313 (N_11313,N_11138,N_11084);
nor U11314 (N_11314,N_11139,N_11007);
or U11315 (N_11315,N_11161,N_11063);
nor U11316 (N_11316,N_11027,N_11017);
nor U11317 (N_11317,N_11086,N_11052);
and U11318 (N_11318,N_11186,N_11002);
and U11319 (N_11319,N_11181,N_11018);
and U11320 (N_11320,N_11186,N_11166);
or U11321 (N_11321,N_11080,N_11099);
and U11322 (N_11322,N_11157,N_11068);
nor U11323 (N_11323,N_11147,N_11146);
xor U11324 (N_11324,N_11191,N_11007);
xnor U11325 (N_11325,N_11164,N_11042);
or U11326 (N_11326,N_11091,N_11036);
xnor U11327 (N_11327,N_11187,N_11064);
and U11328 (N_11328,N_11053,N_11084);
nor U11329 (N_11329,N_11022,N_11072);
or U11330 (N_11330,N_11099,N_11084);
and U11331 (N_11331,N_11063,N_11110);
nor U11332 (N_11332,N_11033,N_11025);
nor U11333 (N_11333,N_11128,N_11023);
and U11334 (N_11334,N_11135,N_11114);
nand U11335 (N_11335,N_11112,N_11146);
nand U11336 (N_11336,N_11113,N_11157);
nor U11337 (N_11337,N_11149,N_11181);
nor U11338 (N_11338,N_11179,N_11008);
nor U11339 (N_11339,N_11182,N_11189);
or U11340 (N_11340,N_11106,N_11090);
nand U11341 (N_11341,N_11186,N_11138);
nand U11342 (N_11342,N_11188,N_11162);
xor U11343 (N_11343,N_11047,N_11030);
nand U11344 (N_11344,N_11171,N_11169);
and U11345 (N_11345,N_11176,N_11093);
nand U11346 (N_11346,N_11027,N_11195);
nor U11347 (N_11347,N_11122,N_11184);
xor U11348 (N_11348,N_11118,N_11180);
xnor U11349 (N_11349,N_11169,N_11162);
and U11350 (N_11350,N_11065,N_11089);
nand U11351 (N_11351,N_11102,N_11067);
or U11352 (N_11352,N_11187,N_11057);
nand U11353 (N_11353,N_11059,N_11105);
and U11354 (N_11354,N_11190,N_11154);
nor U11355 (N_11355,N_11120,N_11032);
and U11356 (N_11356,N_11106,N_11069);
or U11357 (N_11357,N_11122,N_11166);
nand U11358 (N_11358,N_11189,N_11047);
nand U11359 (N_11359,N_11114,N_11016);
and U11360 (N_11360,N_11086,N_11105);
or U11361 (N_11361,N_11143,N_11186);
and U11362 (N_11362,N_11199,N_11039);
xor U11363 (N_11363,N_11043,N_11166);
nor U11364 (N_11364,N_11131,N_11113);
xnor U11365 (N_11365,N_11012,N_11097);
xnor U11366 (N_11366,N_11053,N_11177);
xor U11367 (N_11367,N_11028,N_11178);
xnor U11368 (N_11368,N_11167,N_11162);
nor U11369 (N_11369,N_11109,N_11014);
and U11370 (N_11370,N_11004,N_11053);
or U11371 (N_11371,N_11104,N_11133);
xor U11372 (N_11372,N_11084,N_11061);
xor U11373 (N_11373,N_11007,N_11151);
and U11374 (N_11374,N_11070,N_11107);
or U11375 (N_11375,N_11164,N_11155);
nor U11376 (N_11376,N_11168,N_11031);
nand U11377 (N_11377,N_11131,N_11156);
nand U11378 (N_11378,N_11004,N_11007);
nor U11379 (N_11379,N_11068,N_11057);
nor U11380 (N_11380,N_11186,N_11006);
nor U11381 (N_11381,N_11101,N_11075);
and U11382 (N_11382,N_11062,N_11083);
xor U11383 (N_11383,N_11093,N_11082);
nand U11384 (N_11384,N_11006,N_11162);
and U11385 (N_11385,N_11001,N_11003);
or U11386 (N_11386,N_11089,N_11192);
nor U11387 (N_11387,N_11054,N_11073);
nand U11388 (N_11388,N_11088,N_11130);
or U11389 (N_11389,N_11128,N_11187);
or U11390 (N_11390,N_11078,N_11199);
or U11391 (N_11391,N_11084,N_11085);
or U11392 (N_11392,N_11115,N_11015);
and U11393 (N_11393,N_11146,N_11000);
and U11394 (N_11394,N_11062,N_11022);
and U11395 (N_11395,N_11051,N_11067);
xnor U11396 (N_11396,N_11105,N_11017);
nand U11397 (N_11397,N_11006,N_11121);
or U11398 (N_11398,N_11046,N_11086);
or U11399 (N_11399,N_11077,N_11005);
and U11400 (N_11400,N_11264,N_11387);
or U11401 (N_11401,N_11205,N_11254);
and U11402 (N_11402,N_11275,N_11230);
and U11403 (N_11403,N_11386,N_11296);
or U11404 (N_11404,N_11299,N_11348);
nor U11405 (N_11405,N_11220,N_11247);
nand U11406 (N_11406,N_11289,N_11242);
and U11407 (N_11407,N_11306,N_11326);
nor U11408 (N_11408,N_11375,N_11227);
nand U11409 (N_11409,N_11384,N_11245);
or U11410 (N_11410,N_11368,N_11244);
nand U11411 (N_11411,N_11365,N_11304);
nand U11412 (N_11412,N_11251,N_11257);
xnor U11413 (N_11413,N_11288,N_11223);
nand U11414 (N_11414,N_11248,N_11323);
nor U11415 (N_11415,N_11284,N_11294);
or U11416 (N_11416,N_11238,N_11313);
nand U11417 (N_11417,N_11253,N_11331);
nand U11418 (N_11418,N_11338,N_11249);
and U11419 (N_11419,N_11312,N_11369);
xnor U11420 (N_11420,N_11340,N_11382);
nand U11421 (N_11421,N_11266,N_11291);
xnor U11422 (N_11422,N_11315,N_11351);
nand U11423 (N_11423,N_11224,N_11317);
or U11424 (N_11424,N_11343,N_11236);
and U11425 (N_11425,N_11268,N_11350);
and U11426 (N_11426,N_11240,N_11255);
nand U11427 (N_11427,N_11283,N_11363);
or U11428 (N_11428,N_11278,N_11208);
nand U11429 (N_11429,N_11209,N_11393);
xnor U11430 (N_11430,N_11341,N_11307);
or U11431 (N_11431,N_11310,N_11217);
nand U11432 (N_11432,N_11328,N_11346);
nor U11433 (N_11433,N_11392,N_11279);
nand U11434 (N_11434,N_11308,N_11243);
nand U11435 (N_11435,N_11270,N_11259);
nand U11436 (N_11436,N_11290,N_11221);
nand U11437 (N_11437,N_11399,N_11324);
nand U11438 (N_11438,N_11287,N_11394);
or U11439 (N_11439,N_11318,N_11335);
or U11440 (N_11440,N_11303,N_11272);
xnor U11441 (N_11441,N_11252,N_11214);
nor U11442 (N_11442,N_11302,N_11206);
xnor U11443 (N_11443,N_11321,N_11200);
xor U11444 (N_11444,N_11362,N_11219);
xnor U11445 (N_11445,N_11202,N_11261);
and U11446 (N_11446,N_11285,N_11235);
and U11447 (N_11447,N_11391,N_11273);
and U11448 (N_11448,N_11396,N_11234);
xor U11449 (N_11449,N_11329,N_11352);
or U11450 (N_11450,N_11359,N_11280);
nor U11451 (N_11451,N_11383,N_11311);
nor U11452 (N_11452,N_11390,N_11305);
nand U11453 (N_11453,N_11357,N_11298);
xnor U11454 (N_11454,N_11366,N_11228);
and U11455 (N_11455,N_11314,N_11262);
xor U11456 (N_11456,N_11211,N_11295);
nor U11457 (N_11457,N_11374,N_11241);
or U11458 (N_11458,N_11376,N_11388);
nand U11459 (N_11459,N_11334,N_11322);
and U11460 (N_11460,N_11282,N_11381);
nand U11461 (N_11461,N_11395,N_11274);
nor U11462 (N_11462,N_11319,N_11316);
nor U11463 (N_11463,N_11336,N_11256);
nor U11464 (N_11464,N_11300,N_11226);
and U11465 (N_11465,N_11276,N_11372);
xnor U11466 (N_11466,N_11309,N_11229);
xor U11467 (N_11467,N_11373,N_11207);
xnor U11468 (N_11468,N_11397,N_11201);
nor U11469 (N_11469,N_11204,N_11320);
nand U11470 (N_11470,N_11237,N_11339);
or U11471 (N_11471,N_11398,N_11250);
nor U11472 (N_11472,N_11233,N_11286);
and U11473 (N_11473,N_11337,N_11216);
nor U11474 (N_11474,N_11330,N_11239);
and U11475 (N_11475,N_11263,N_11360);
and U11476 (N_11476,N_11378,N_11342);
nand U11477 (N_11477,N_11379,N_11364);
xor U11478 (N_11478,N_11349,N_11277);
nor U11479 (N_11479,N_11327,N_11325);
nor U11480 (N_11480,N_11213,N_11267);
xnor U11481 (N_11481,N_11222,N_11377);
nor U11482 (N_11482,N_11370,N_11269);
xnor U11483 (N_11483,N_11260,N_11218);
nand U11484 (N_11484,N_11225,N_11347);
xor U11485 (N_11485,N_11345,N_11265);
and U11486 (N_11486,N_11212,N_11271);
and U11487 (N_11487,N_11215,N_11354);
nand U11488 (N_11488,N_11353,N_11297);
and U11489 (N_11489,N_11344,N_11385);
nor U11490 (N_11490,N_11301,N_11281);
or U11491 (N_11491,N_11293,N_11231);
or U11492 (N_11492,N_11389,N_11380);
nor U11493 (N_11493,N_11358,N_11333);
or U11494 (N_11494,N_11203,N_11355);
or U11495 (N_11495,N_11361,N_11332);
and U11496 (N_11496,N_11292,N_11367);
or U11497 (N_11497,N_11210,N_11232);
nand U11498 (N_11498,N_11246,N_11371);
nor U11499 (N_11499,N_11356,N_11258);
nor U11500 (N_11500,N_11285,N_11322);
nor U11501 (N_11501,N_11277,N_11262);
nand U11502 (N_11502,N_11360,N_11342);
or U11503 (N_11503,N_11261,N_11209);
xor U11504 (N_11504,N_11348,N_11200);
or U11505 (N_11505,N_11266,N_11392);
xor U11506 (N_11506,N_11388,N_11239);
nand U11507 (N_11507,N_11304,N_11378);
or U11508 (N_11508,N_11361,N_11318);
nor U11509 (N_11509,N_11310,N_11360);
or U11510 (N_11510,N_11347,N_11387);
or U11511 (N_11511,N_11364,N_11279);
xnor U11512 (N_11512,N_11223,N_11250);
and U11513 (N_11513,N_11311,N_11378);
nand U11514 (N_11514,N_11347,N_11290);
nand U11515 (N_11515,N_11206,N_11301);
nor U11516 (N_11516,N_11264,N_11323);
xor U11517 (N_11517,N_11363,N_11217);
xnor U11518 (N_11518,N_11350,N_11314);
and U11519 (N_11519,N_11233,N_11295);
or U11520 (N_11520,N_11258,N_11245);
and U11521 (N_11521,N_11335,N_11239);
or U11522 (N_11522,N_11291,N_11276);
xor U11523 (N_11523,N_11369,N_11339);
xor U11524 (N_11524,N_11211,N_11390);
or U11525 (N_11525,N_11327,N_11224);
nor U11526 (N_11526,N_11348,N_11283);
nor U11527 (N_11527,N_11302,N_11225);
and U11528 (N_11528,N_11216,N_11320);
nor U11529 (N_11529,N_11255,N_11253);
nor U11530 (N_11530,N_11393,N_11227);
and U11531 (N_11531,N_11275,N_11239);
or U11532 (N_11532,N_11373,N_11394);
xnor U11533 (N_11533,N_11346,N_11361);
nand U11534 (N_11534,N_11307,N_11355);
xnor U11535 (N_11535,N_11362,N_11363);
nand U11536 (N_11536,N_11380,N_11219);
or U11537 (N_11537,N_11274,N_11391);
and U11538 (N_11538,N_11370,N_11307);
nand U11539 (N_11539,N_11345,N_11256);
and U11540 (N_11540,N_11382,N_11375);
nand U11541 (N_11541,N_11390,N_11357);
nor U11542 (N_11542,N_11320,N_11287);
and U11543 (N_11543,N_11399,N_11292);
or U11544 (N_11544,N_11270,N_11362);
nor U11545 (N_11545,N_11213,N_11251);
xnor U11546 (N_11546,N_11378,N_11352);
nor U11547 (N_11547,N_11275,N_11359);
and U11548 (N_11548,N_11201,N_11365);
or U11549 (N_11549,N_11391,N_11362);
xnor U11550 (N_11550,N_11386,N_11269);
nand U11551 (N_11551,N_11209,N_11258);
nand U11552 (N_11552,N_11226,N_11391);
and U11553 (N_11553,N_11295,N_11334);
xor U11554 (N_11554,N_11373,N_11335);
nor U11555 (N_11555,N_11259,N_11320);
nor U11556 (N_11556,N_11264,N_11334);
nor U11557 (N_11557,N_11317,N_11244);
and U11558 (N_11558,N_11219,N_11329);
nor U11559 (N_11559,N_11387,N_11213);
nand U11560 (N_11560,N_11361,N_11249);
nor U11561 (N_11561,N_11383,N_11361);
and U11562 (N_11562,N_11395,N_11371);
nor U11563 (N_11563,N_11380,N_11383);
xor U11564 (N_11564,N_11339,N_11305);
or U11565 (N_11565,N_11209,N_11255);
nor U11566 (N_11566,N_11398,N_11286);
nor U11567 (N_11567,N_11365,N_11227);
nand U11568 (N_11568,N_11398,N_11356);
and U11569 (N_11569,N_11257,N_11260);
nand U11570 (N_11570,N_11224,N_11245);
nor U11571 (N_11571,N_11335,N_11249);
nor U11572 (N_11572,N_11249,N_11214);
xnor U11573 (N_11573,N_11378,N_11234);
nor U11574 (N_11574,N_11285,N_11341);
or U11575 (N_11575,N_11248,N_11285);
nand U11576 (N_11576,N_11256,N_11238);
nand U11577 (N_11577,N_11383,N_11350);
xor U11578 (N_11578,N_11272,N_11389);
and U11579 (N_11579,N_11203,N_11397);
or U11580 (N_11580,N_11243,N_11379);
xnor U11581 (N_11581,N_11298,N_11394);
or U11582 (N_11582,N_11351,N_11221);
nor U11583 (N_11583,N_11322,N_11262);
xnor U11584 (N_11584,N_11267,N_11245);
or U11585 (N_11585,N_11237,N_11352);
and U11586 (N_11586,N_11313,N_11249);
or U11587 (N_11587,N_11231,N_11291);
nor U11588 (N_11588,N_11214,N_11229);
and U11589 (N_11589,N_11279,N_11354);
and U11590 (N_11590,N_11247,N_11377);
nand U11591 (N_11591,N_11318,N_11259);
xor U11592 (N_11592,N_11230,N_11308);
and U11593 (N_11593,N_11215,N_11336);
nor U11594 (N_11594,N_11359,N_11216);
and U11595 (N_11595,N_11206,N_11316);
or U11596 (N_11596,N_11282,N_11348);
xnor U11597 (N_11597,N_11360,N_11201);
nand U11598 (N_11598,N_11249,N_11207);
and U11599 (N_11599,N_11255,N_11237);
xnor U11600 (N_11600,N_11406,N_11469);
xnor U11601 (N_11601,N_11586,N_11513);
and U11602 (N_11602,N_11403,N_11501);
xnor U11603 (N_11603,N_11477,N_11490);
xnor U11604 (N_11604,N_11457,N_11499);
or U11605 (N_11605,N_11575,N_11409);
or U11606 (N_11606,N_11464,N_11565);
or U11607 (N_11607,N_11421,N_11502);
or U11608 (N_11608,N_11574,N_11595);
xor U11609 (N_11609,N_11436,N_11516);
xor U11610 (N_11610,N_11488,N_11413);
or U11611 (N_11611,N_11466,N_11536);
or U11612 (N_11612,N_11440,N_11431);
xor U11613 (N_11613,N_11582,N_11590);
or U11614 (N_11614,N_11437,N_11427);
and U11615 (N_11615,N_11529,N_11493);
xnor U11616 (N_11616,N_11562,N_11423);
or U11617 (N_11617,N_11564,N_11571);
nand U11618 (N_11618,N_11456,N_11503);
and U11619 (N_11619,N_11504,N_11510);
nand U11620 (N_11620,N_11455,N_11468);
and U11621 (N_11621,N_11434,N_11446);
nand U11622 (N_11622,N_11400,N_11439);
xnor U11623 (N_11623,N_11546,N_11535);
xnor U11624 (N_11624,N_11572,N_11581);
nand U11625 (N_11625,N_11524,N_11452);
or U11626 (N_11626,N_11419,N_11540);
nand U11627 (N_11627,N_11578,N_11459);
xnor U11628 (N_11628,N_11460,N_11521);
nand U11629 (N_11629,N_11476,N_11541);
nor U11630 (N_11630,N_11430,N_11465);
or U11631 (N_11631,N_11569,N_11560);
and U11632 (N_11632,N_11515,N_11534);
xor U11633 (N_11633,N_11444,N_11483);
and U11634 (N_11634,N_11544,N_11429);
or U11635 (N_11635,N_11495,N_11438);
or U11636 (N_11636,N_11550,N_11485);
nand U11637 (N_11637,N_11432,N_11507);
and U11638 (N_11638,N_11486,N_11598);
or U11639 (N_11639,N_11551,N_11523);
or U11640 (N_11640,N_11599,N_11472);
xnor U11641 (N_11641,N_11553,N_11498);
xnor U11642 (N_11642,N_11487,N_11597);
nor U11643 (N_11643,N_11505,N_11508);
or U11644 (N_11644,N_11518,N_11528);
or U11645 (N_11645,N_11412,N_11527);
or U11646 (N_11646,N_11484,N_11537);
xor U11647 (N_11647,N_11454,N_11407);
or U11648 (N_11648,N_11414,N_11522);
nor U11649 (N_11649,N_11426,N_11471);
xnor U11650 (N_11650,N_11568,N_11566);
xnor U11651 (N_11651,N_11418,N_11467);
xnor U11652 (N_11652,N_11428,N_11447);
nor U11653 (N_11653,N_11593,N_11482);
and U11654 (N_11654,N_11470,N_11496);
xnor U11655 (N_11655,N_11538,N_11517);
nor U11656 (N_11656,N_11443,N_11579);
and U11657 (N_11657,N_11549,N_11494);
and U11658 (N_11658,N_11405,N_11547);
xor U11659 (N_11659,N_11401,N_11449);
and U11660 (N_11660,N_11417,N_11463);
or U11661 (N_11661,N_11570,N_11489);
and U11662 (N_11662,N_11475,N_11596);
nand U11663 (N_11663,N_11461,N_11552);
nand U11664 (N_11664,N_11448,N_11500);
or U11665 (N_11665,N_11577,N_11583);
and U11666 (N_11666,N_11585,N_11411);
xor U11667 (N_11667,N_11458,N_11531);
and U11668 (N_11668,N_11408,N_11556);
xnor U11669 (N_11669,N_11480,N_11402);
nor U11670 (N_11670,N_11543,N_11462);
nor U11671 (N_11671,N_11587,N_11433);
nor U11672 (N_11672,N_11545,N_11514);
nand U11673 (N_11673,N_11591,N_11559);
or U11674 (N_11674,N_11453,N_11473);
and U11675 (N_11675,N_11592,N_11584);
or U11676 (N_11676,N_11520,N_11506);
xor U11677 (N_11677,N_11404,N_11410);
or U11678 (N_11678,N_11451,N_11424);
nor U11679 (N_11679,N_11563,N_11573);
or U11680 (N_11680,N_11415,N_11512);
nand U11681 (N_11681,N_11532,N_11533);
nand U11682 (N_11682,N_11478,N_11557);
or U11683 (N_11683,N_11479,N_11555);
nand U11684 (N_11684,N_11554,N_11526);
nand U11685 (N_11685,N_11511,N_11588);
xor U11686 (N_11686,N_11558,N_11491);
xor U11687 (N_11687,N_11576,N_11441);
nand U11688 (N_11688,N_11580,N_11567);
nor U11689 (N_11689,N_11519,N_11497);
nor U11690 (N_11690,N_11525,N_11450);
and U11691 (N_11691,N_11589,N_11492);
or U11692 (N_11692,N_11561,N_11420);
nor U11693 (N_11693,N_11481,N_11425);
nor U11694 (N_11694,N_11509,N_11416);
xor U11695 (N_11695,N_11539,N_11435);
or U11696 (N_11696,N_11542,N_11594);
nand U11697 (N_11697,N_11474,N_11548);
or U11698 (N_11698,N_11530,N_11422);
nand U11699 (N_11699,N_11445,N_11442);
or U11700 (N_11700,N_11403,N_11547);
or U11701 (N_11701,N_11411,N_11509);
xor U11702 (N_11702,N_11595,N_11472);
nand U11703 (N_11703,N_11576,N_11515);
nor U11704 (N_11704,N_11504,N_11419);
nor U11705 (N_11705,N_11595,N_11540);
and U11706 (N_11706,N_11405,N_11531);
xnor U11707 (N_11707,N_11571,N_11552);
nand U11708 (N_11708,N_11496,N_11508);
nor U11709 (N_11709,N_11432,N_11537);
nor U11710 (N_11710,N_11447,N_11455);
or U11711 (N_11711,N_11540,N_11477);
nor U11712 (N_11712,N_11595,N_11514);
nand U11713 (N_11713,N_11505,N_11477);
xnor U11714 (N_11714,N_11589,N_11493);
and U11715 (N_11715,N_11459,N_11531);
and U11716 (N_11716,N_11446,N_11420);
nand U11717 (N_11717,N_11551,N_11492);
or U11718 (N_11718,N_11521,N_11406);
xnor U11719 (N_11719,N_11429,N_11403);
or U11720 (N_11720,N_11551,N_11516);
nand U11721 (N_11721,N_11413,N_11469);
xnor U11722 (N_11722,N_11539,N_11529);
nor U11723 (N_11723,N_11535,N_11515);
xnor U11724 (N_11724,N_11456,N_11577);
nand U11725 (N_11725,N_11416,N_11557);
or U11726 (N_11726,N_11591,N_11435);
nor U11727 (N_11727,N_11402,N_11561);
xor U11728 (N_11728,N_11526,N_11486);
and U11729 (N_11729,N_11526,N_11445);
nand U11730 (N_11730,N_11521,N_11556);
nand U11731 (N_11731,N_11583,N_11514);
nand U11732 (N_11732,N_11569,N_11457);
nor U11733 (N_11733,N_11485,N_11470);
xor U11734 (N_11734,N_11531,N_11543);
or U11735 (N_11735,N_11598,N_11434);
xnor U11736 (N_11736,N_11452,N_11443);
xor U11737 (N_11737,N_11489,N_11579);
xnor U11738 (N_11738,N_11450,N_11487);
nand U11739 (N_11739,N_11538,N_11503);
xnor U11740 (N_11740,N_11461,N_11596);
nor U11741 (N_11741,N_11479,N_11498);
xor U11742 (N_11742,N_11590,N_11439);
and U11743 (N_11743,N_11549,N_11525);
and U11744 (N_11744,N_11553,N_11423);
xor U11745 (N_11745,N_11527,N_11469);
or U11746 (N_11746,N_11458,N_11420);
and U11747 (N_11747,N_11525,N_11594);
and U11748 (N_11748,N_11540,N_11444);
nand U11749 (N_11749,N_11450,N_11401);
and U11750 (N_11750,N_11427,N_11483);
and U11751 (N_11751,N_11471,N_11419);
and U11752 (N_11752,N_11481,N_11599);
nor U11753 (N_11753,N_11584,N_11583);
and U11754 (N_11754,N_11537,N_11493);
or U11755 (N_11755,N_11499,N_11525);
nor U11756 (N_11756,N_11508,N_11461);
xor U11757 (N_11757,N_11554,N_11569);
or U11758 (N_11758,N_11475,N_11400);
nand U11759 (N_11759,N_11513,N_11408);
nor U11760 (N_11760,N_11526,N_11563);
nand U11761 (N_11761,N_11450,N_11559);
nand U11762 (N_11762,N_11533,N_11407);
nand U11763 (N_11763,N_11447,N_11505);
or U11764 (N_11764,N_11492,N_11482);
or U11765 (N_11765,N_11409,N_11437);
and U11766 (N_11766,N_11553,N_11566);
nor U11767 (N_11767,N_11525,N_11555);
xnor U11768 (N_11768,N_11431,N_11497);
and U11769 (N_11769,N_11468,N_11595);
xnor U11770 (N_11770,N_11491,N_11537);
nand U11771 (N_11771,N_11555,N_11419);
xor U11772 (N_11772,N_11439,N_11586);
nand U11773 (N_11773,N_11566,N_11520);
nand U11774 (N_11774,N_11511,N_11583);
or U11775 (N_11775,N_11485,N_11510);
or U11776 (N_11776,N_11572,N_11554);
or U11777 (N_11777,N_11449,N_11472);
or U11778 (N_11778,N_11506,N_11437);
and U11779 (N_11779,N_11474,N_11587);
nor U11780 (N_11780,N_11466,N_11470);
and U11781 (N_11781,N_11425,N_11525);
or U11782 (N_11782,N_11408,N_11450);
and U11783 (N_11783,N_11594,N_11469);
nor U11784 (N_11784,N_11485,N_11489);
nor U11785 (N_11785,N_11421,N_11413);
or U11786 (N_11786,N_11529,N_11528);
nor U11787 (N_11787,N_11509,N_11408);
or U11788 (N_11788,N_11578,N_11591);
or U11789 (N_11789,N_11561,N_11560);
nor U11790 (N_11790,N_11567,N_11471);
and U11791 (N_11791,N_11492,N_11572);
xnor U11792 (N_11792,N_11578,N_11570);
xnor U11793 (N_11793,N_11474,N_11460);
xnor U11794 (N_11794,N_11419,N_11432);
nand U11795 (N_11795,N_11436,N_11465);
nor U11796 (N_11796,N_11573,N_11593);
and U11797 (N_11797,N_11528,N_11448);
nand U11798 (N_11798,N_11539,N_11442);
xnor U11799 (N_11799,N_11562,N_11558);
or U11800 (N_11800,N_11688,N_11708);
xor U11801 (N_11801,N_11697,N_11640);
and U11802 (N_11802,N_11775,N_11644);
nor U11803 (N_11803,N_11729,N_11645);
nand U11804 (N_11804,N_11751,N_11766);
nor U11805 (N_11805,N_11611,N_11612);
or U11806 (N_11806,N_11764,N_11681);
and U11807 (N_11807,N_11632,N_11713);
or U11808 (N_11808,N_11723,N_11687);
xnor U11809 (N_11809,N_11718,N_11701);
and U11810 (N_11810,N_11670,N_11780);
xnor U11811 (N_11811,N_11761,N_11743);
nor U11812 (N_11812,N_11606,N_11756);
and U11813 (N_11813,N_11628,N_11745);
and U11814 (N_11814,N_11702,N_11750);
or U11815 (N_11815,N_11652,N_11758);
nor U11816 (N_11816,N_11667,N_11793);
or U11817 (N_11817,N_11621,N_11658);
nand U11818 (N_11818,N_11655,N_11608);
and U11819 (N_11819,N_11796,N_11774);
and U11820 (N_11820,N_11685,N_11748);
xor U11821 (N_11821,N_11777,N_11619);
or U11822 (N_11822,N_11650,N_11671);
xnor U11823 (N_11823,N_11740,N_11782);
nand U11824 (N_11824,N_11613,N_11733);
or U11825 (N_11825,N_11771,N_11705);
or U11826 (N_11826,N_11712,N_11639);
nor U11827 (N_11827,N_11629,N_11770);
xnor U11828 (N_11828,N_11785,N_11732);
nor U11829 (N_11829,N_11675,N_11624);
or U11830 (N_11830,N_11676,N_11604);
nor U11831 (N_11831,N_11794,N_11679);
or U11832 (N_11832,N_11616,N_11772);
nand U11833 (N_11833,N_11752,N_11762);
nand U11834 (N_11834,N_11672,N_11668);
or U11835 (N_11835,N_11631,N_11678);
xor U11836 (N_11836,N_11686,N_11765);
nor U11837 (N_11837,N_11635,N_11703);
xor U11838 (N_11838,N_11790,N_11614);
nor U11839 (N_11839,N_11789,N_11783);
nand U11840 (N_11840,N_11634,N_11649);
and U11841 (N_11841,N_11730,N_11754);
nand U11842 (N_11842,N_11601,N_11735);
nand U11843 (N_11843,N_11673,N_11623);
or U11844 (N_11844,N_11647,N_11636);
xnor U11845 (N_11845,N_11725,N_11674);
and U11846 (N_11846,N_11746,N_11788);
xnor U11847 (N_11847,N_11741,N_11615);
xor U11848 (N_11848,N_11798,N_11714);
or U11849 (N_11849,N_11602,N_11659);
xnor U11850 (N_11850,N_11707,N_11792);
nand U11851 (N_11851,N_11749,N_11727);
xnor U11852 (N_11852,N_11695,N_11620);
or U11853 (N_11853,N_11776,N_11609);
nand U11854 (N_11854,N_11737,N_11665);
and U11855 (N_11855,N_11654,N_11779);
and U11856 (N_11856,N_11747,N_11716);
xor U11857 (N_11857,N_11691,N_11637);
or U11858 (N_11858,N_11662,N_11651);
nor U11859 (N_11859,N_11700,N_11719);
nor U11860 (N_11860,N_11696,N_11753);
nand U11861 (N_11861,N_11627,N_11784);
nor U11862 (N_11862,N_11622,N_11757);
xnor U11863 (N_11863,N_11607,N_11680);
and U11864 (N_11864,N_11664,N_11663);
or U11865 (N_11865,N_11646,N_11641);
xor U11866 (N_11866,N_11699,N_11692);
nor U11867 (N_11867,N_11630,N_11661);
xnor U11868 (N_11868,N_11638,N_11739);
nor U11869 (N_11869,N_11689,N_11722);
nand U11870 (N_11870,N_11666,N_11715);
and U11871 (N_11871,N_11724,N_11642);
nor U11872 (N_11872,N_11797,N_11768);
xor U11873 (N_11873,N_11605,N_11726);
nand U11874 (N_11874,N_11781,N_11704);
xnor U11875 (N_11875,N_11738,N_11684);
nand U11876 (N_11876,N_11709,N_11791);
xnor U11877 (N_11877,N_11690,N_11734);
nand U11878 (N_11878,N_11698,N_11767);
and U11879 (N_11879,N_11603,N_11710);
and U11880 (N_11880,N_11760,N_11677);
nand U11881 (N_11881,N_11643,N_11693);
and U11882 (N_11882,N_11653,N_11633);
and U11883 (N_11883,N_11769,N_11625);
or U11884 (N_11884,N_11755,N_11763);
and U11885 (N_11885,N_11600,N_11682);
xnor U11886 (N_11886,N_11799,N_11660);
nand U11887 (N_11887,N_11717,N_11711);
nand U11888 (N_11888,N_11618,N_11683);
and U11889 (N_11889,N_11742,N_11610);
nand U11890 (N_11890,N_11731,N_11795);
or U11891 (N_11891,N_11720,N_11626);
nand U11892 (N_11892,N_11694,N_11617);
and U11893 (N_11893,N_11773,N_11706);
xor U11894 (N_11894,N_11786,N_11669);
nand U11895 (N_11895,N_11759,N_11656);
nand U11896 (N_11896,N_11736,N_11744);
and U11897 (N_11897,N_11657,N_11721);
nand U11898 (N_11898,N_11648,N_11728);
or U11899 (N_11899,N_11787,N_11778);
nand U11900 (N_11900,N_11735,N_11708);
and U11901 (N_11901,N_11691,N_11798);
or U11902 (N_11902,N_11621,N_11724);
and U11903 (N_11903,N_11628,N_11729);
and U11904 (N_11904,N_11661,N_11732);
nand U11905 (N_11905,N_11723,N_11656);
xor U11906 (N_11906,N_11769,N_11708);
or U11907 (N_11907,N_11721,N_11755);
nand U11908 (N_11908,N_11708,N_11611);
or U11909 (N_11909,N_11684,N_11669);
nor U11910 (N_11910,N_11798,N_11771);
or U11911 (N_11911,N_11791,N_11755);
nand U11912 (N_11912,N_11600,N_11641);
xnor U11913 (N_11913,N_11790,N_11742);
or U11914 (N_11914,N_11708,N_11782);
nand U11915 (N_11915,N_11777,N_11607);
and U11916 (N_11916,N_11742,N_11786);
xor U11917 (N_11917,N_11794,N_11625);
nor U11918 (N_11918,N_11763,N_11659);
and U11919 (N_11919,N_11624,N_11653);
nand U11920 (N_11920,N_11618,N_11645);
nor U11921 (N_11921,N_11784,N_11619);
and U11922 (N_11922,N_11660,N_11762);
nand U11923 (N_11923,N_11688,N_11723);
and U11924 (N_11924,N_11611,N_11671);
and U11925 (N_11925,N_11608,N_11611);
xnor U11926 (N_11926,N_11670,N_11685);
or U11927 (N_11927,N_11741,N_11772);
xnor U11928 (N_11928,N_11717,N_11684);
and U11929 (N_11929,N_11619,N_11656);
xor U11930 (N_11930,N_11620,N_11636);
or U11931 (N_11931,N_11799,N_11650);
nor U11932 (N_11932,N_11755,N_11752);
or U11933 (N_11933,N_11648,N_11631);
nand U11934 (N_11934,N_11690,N_11697);
xnor U11935 (N_11935,N_11602,N_11677);
and U11936 (N_11936,N_11621,N_11628);
xor U11937 (N_11937,N_11680,N_11714);
nand U11938 (N_11938,N_11671,N_11734);
xnor U11939 (N_11939,N_11642,N_11665);
nor U11940 (N_11940,N_11604,N_11697);
nand U11941 (N_11941,N_11651,N_11762);
xnor U11942 (N_11942,N_11667,N_11773);
or U11943 (N_11943,N_11725,N_11697);
nand U11944 (N_11944,N_11652,N_11600);
nor U11945 (N_11945,N_11764,N_11617);
nor U11946 (N_11946,N_11739,N_11759);
nor U11947 (N_11947,N_11725,N_11614);
and U11948 (N_11948,N_11788,N_11648);
nand U11949 (N_11949,N_11611,N_11659);
nand U11950 (N_11950,N_11671,N_11779);
xnor U11951 (N_11951,N_11751,N_11605);
or U11952 (N_11952,N_11687,N_11699);
nor U11953 (N_11953,N_11781,N_11706);
or U11954 (N_11954,N_11721,N_11775);
nand U11955 (N_11955,N_11661,N_11750);
or U11956 (N_11956,N_11712,N_11749);
xor U11957 (N_11957,N_11623,N_11691);
nand U11958 (N_11958,N_11702,N_11785);
nor U11959 (N_11959,N_11674,N_11618);
or U11960 (N_11960,N_11619,N_11737);
or U11961 (N_11961,N_11714,N_11653);
nand U11962 (N_11962,N_11795,N_11685);
and U11963 (N_11963,N_11617,N_11681);
and U11964 (N_11964,N_11794,N_11702);
and U11965 (N_11965,N_11648,N_11611);
nor U11966 (N_11966,N_11747,N_11619);
and U11967 (N_11967,N_11727,N_11647);
nor U11968 (N_11968,N_11610,N_11691);
and U11969 (N_11969,N_11725,N_11798);
xor U11970 (N_11970,N_11741,N_11678);
xnor U11971 (N_11971,N_11706,N_11736);
nand U11972 (N_11972,N_11708,N_11731);
and U11973 (N_11973,N_11703,N_11637);
xor U11974 (N_11974,N_11775,N_11656);
and U11975 (N_11975,N_11653,N_11781);
xor U11976 (N_11976,N_11712,N_11693);
xnor U11977 (N_11977,N_11790,N_11744);
nor U11978 (N_11978,N_11650,N_11771);
or U11979 (N_11979,N_11616,N_11683);
nor U11980 (N_11980,N_11615,N_11630);
and U11981 (N_11981,N_11764,N_11780);
nand U11982 (N_11982,N_11650,N_11730);
and U11983 (N_11983,N_11702,N_11796);
nor U11984 (N_11984,N_11695,N_11765);
and U11985 (N_11985,N_11624,N_11781);
and U11986 (N_11986,N_11695,N_11797);
or U11987 (N_11987,N_11773,N_11795);
or U11988 (N_11988,N_11788,N_11651);
nor U11989 (N_11989,N_11714,N_11604);
nor U11990 (N_11990,N_11633,N_11671);
nor U11991 (N_11991,N_11720,N_11773);
nand U11992 (N_11992,N_11679,N_11788);
nand U11993 (N_11993,N_11670,N_11671);
or U11994 (N_11994,N_11742,N_11777);
nand U11995 (N_11995,N_11711,N_11747);
or U11996 (N_11996,N_11714,N_11740);
xor U11997 (N_11997,N_11634,N_11728);
or U11998 (N_11998,N_11704,N_11608);
and U11999 (N_11999,N_11755,N_11646);
nand U12000 (N_12000,N_11840,N_11952);
or U12001 (N_12001,N_11881,N_11839);
xor U12002 (N_12002,N_11927,N_11871);
nand U12003 (N_12003,N_11940,N_11959);
nor U12004 (N_12004,N_11936,N_11833);
and U12005 (N_12005,N_11815,N_11864);
or U12006 (N_12006,N_11931,N_11924);
xnor U12007 (N_12007,N_11846,N_11895);
or U12008 (N_12008,N_11963,N_11961);
and U12009 (N_12009,N_11879,N_11908);
or U12010 (N_12010,N_11844,N_11910);
xor U12011 (N_12011,N_11855,N_11824);
xor U12012 (N_12012,N_11980,N_11923);
or U12013 (N_12013,N_11872,N_11907);
nand U12014 (N_12014,N_11922,N_11889);
or U12015 (N_12015,N_11865,N_11848);
nor U12016 (N_12016,N_11987,N_11949);
xor U12017 (N_12017,N_11983,N_11991);
nand U12018 (N_12018,N_11878,N_11828);
nand U12019 (N_12019,N_11918,N_11974);
and U12020 (N_12020,N_11926,N_11929);
and U12021 (N_12021,N_11985,N_11984);
nor U12022 (N_12022,N_11847,N_11986);
or U12023 (N_12023,N_11867,N_11838);
and U12024 (N_12024,N_11802,N_11831);
nor U12025 (N_12025,N_11965,N_11860);
nand U12026 (N_12026,N_11972,N_11995);
and U12027 (N_12027,N_11957,N_11836);
nor U12028 (N_12028,N_11964,N_11928);
nand U12029 (N_12029,N_11829,N_11905);
or U12030 (N_12030,N_11874,N_11958);
xnor U12031 (N_12031,N_11885,N_11883);
or U12032 (N_12032,N_11887,N_11911);
nor U12033 (N_12033,N_11835,N_11812);
xor U12034 (N_12034,N_11989,N_11863);
nor U12035 (N_12035,N_11932,N_11937);
xor U12036 (N_12036,N_11998,N_11997);
or U12037 (N_12037,N_11808,N_11853);
and U12038 (N_12038,N_11953,N_11942);
or U12039 (N_12039,N_11822,N_11904);
nand U12040 (N_12040,N_11884,N_11934);
or U12041 (N_12041,N_11823,N_11852);
xnor U12042 (N_12042,N_11819,N_11925);
or U12043 (N_12043,N_11996,N_11939);
or U12044 (N_12044,N_11968,N_11956);
and U12045 (N_12045,N_11827,N_11891);
nand U12046 (N_12046,N_11975,N_11903);
and U12047 (N_12047,N_11811,N_11805);
nand U12048 (N_12048,N_11806,N_11966);
and U12049 (N_12049,N_11861,N_11919);
or U12050 (N_12050,N_11892,N_11821);
nand U12051 (N_12051,N_11859,N_11917);
and U12052 (N_12052,N_11899,N_11938);
nand U12053 (N_12053,N_11837,N_11877);
and U12054 (N_12054,N_11994,N_11981);
xnor U12055 (N_12055,N_11870,N_11955);
and U12056 (N_12056,N_11843,N_11820);
nor U12057 (N_12057,N_11976,N_11888);
and U12058 (N_12058,N_11933,N_11803);
xnor U12059 (N_12059,N_11954,N_11982);
nor U12060 (N_12060,N_11943,N_11830);
nand U12061 (N_12061,N_11886,N_11945);
nand U12062 (N_12062,N_11944,N_11947);
or U12063 (N_12063,N_11915,N_11979);
nand U12064 (N_12064,N_11857,N_11897);
nor U12065 (N_12065,N_11901,N_11898);
or U12066 (N_12066,N_11893,N_11988);
or U12067 (N_12067,N_11967,N_11970);
nand U12068 (N_12068,N_11800,N_11842);
nor U12069 (N_12069,N_11999,N_11946);
and U12070 (N_12070,N_11825,N_11813);
and U12071 (N_12071,N_11935,N_11973);
xnor U12072 (N_12072,N_11950,N_11900);
and U12073 (N_12073,N_11890,N_11801);
nor U12074 (N_12074,N_11809,N_11832);
and U12075 (N_12075,N_11882,N_11948);
and U12076 (N_12076,N_11914,N_11941);
xor U12077 (N_12077,N_11849,N_11909);
xnor U12078 (N_12078,N_11845,N_11894);
nor U12079 (N_12079,N_11807,N_11810);
nand U12080 (N_12080,N_11866,N_11873);
or U12081 (N_12081,N_11921,N_11913);
xnor U12082 (N_12082,N_11978,N_11977);
or U12083 (N_12083,N_11969,N_11993);
nand U12084 (N_12084,N_11868,N_11960);
nand U12085 (N_12085,N_11876,N_11916);
nand U12086 (N_12086,N_11862,N_11851);
nor U12087 (N_12087,N_11826,N_11856);
nor U12088 (N_12088,N_11816,N_11869);
xnor U12089 (N_12089,N_11858,N_11841);
nor U12090 (N_12090,N_11804,N_11875);
xor U12091 (N_12091,N_11930,N_11912);
or U12092 (N_12092,N_11880,N_11854);
nand U12093 (N_12093,N_11906,N_11850);
xnor U12094 (N_12094,N_11896,N_11902);
nand U12095 (N_12095,N_11951,N_11817);
and U12096 (N_12096,N_11814,N_11992);
nor U12097 (N_12097,N_11971,N_11920);
nand U12098 (N_12098,N_11962,N_11834);
and U12099 (N_12099,N_11990,N_11818);
or U12100 (N_12100,N_11992,N_11925);
and U12101 (N_12101,N_11841,N_11943);
nand U12102 (N_12102,N_11937,N_11983);
nand U12103 (N_12103,N_11927,N_11935);
nor U12104 (N_12104,N_11809,N_11976);
nor U12105 (N_12105,N_11953,N_11869);
and U12106 (N_12106,N_11994,N_11872);
nor U12107 (N_12107,N_11922,N_11988);
and U12108 (N_12108,N_11867,N_11849);
nand U12109 (N_12109,N_11831,N_11998);
or U12110 (N_12110,N_11983,N_11965);
or U12111 (N_12111,N_11947,N_11980);
or U12112 (N_12112,N_11915,N_11884);
nand U12113 (N_12113,N_11893,N_11856);
and U12114 (N_12114,N_11985,N_11972);
and U12115 (N_12115,N_11945,N_11831);
xnor U12116 (N_12116,N_11805,N_11981);
nand U12117 (N_12117,N_11813,N_11847);
nor U12118 (N_12118,N_11963,N_11807);
and U12119 (N_12119,N_11973,N_11852);
and U12120 (N_12120,N_11986,N_11857);
nand U12121 (N_12121,N_11850,N_11914);
and U12122 (N_12122,N_11869,N_11994);
nor U12123 (N_12123,N_11990,N_11858);
or U12124 (N_12124,N_11855,N_11984);
or U12125 (N_12125,N_11838,N_11907);
nand U12126 (N_12126,N_11884,N_11802);
xnor U12127 (N_12127,N_11832,N_11858);
or U12128 (N_12128,N_11874,N_11936);
and U12129 (N_12129,N_11913,N_11839);
or U12130 (N_12130,N_11932,N_11802);
nor U12131 (N_12131,N_11863,N_11892);
and U12132 (N_12132,N_11974,N_11948);
nand U12133 (N_12133,N_11898,N_11916);
xnor U12134 (N_12134,N_11841,N_11907);
xor U12135 (N_12135,N_11960,N_11863);
nor U12136 (N_12136,N_11895,N_11827);
nor U12137 (N_12137,N_11975,N_11995);
xnor U12138 (N_12138,N_11869,N_11821);
or U12139 (N_12139,N_11883,N_11917);
xnor U12140 (N_12140,N_11911,N_11890);
nor U12141 (N_12141,N_11906,N_11810);
and U12142 (N_12142,N_11939,N_11877);
and U12143 (N_12143,N_11867,N_11958);
and U12144 (N_12144,N_11859,N_11897);
nand U12145 (N_12145,N_11996,N_11872);
or U12146 (N_12146,N_11833,N_11991);
and U12147 (N_12147,N_11941,N_11833);
xor U12148 (N_12148,N_11886,N_11955);
or U12149 (N_12149,N_11826,N_11912);
nand U12150 (N_12150,N_11975,N_11897);
or U12151 (N_12151,N_11804,N_11866);
and U12152 (N_12152,N_11978,N_11848);
or U12153 (N_12153,N_11904,N_11846);
and U12154 (N_12154,N_11928,N_11936);
xor U12155 (N_12155,N_11853,N_11930);
nor U12156 (N_12156,N_11926,N_11821);
or U12157 (N_12157,N_11847,N_11816);
and U12158 (N_12158,N_11843,N_11937);
or U12159 (N_12159,N_11820,N_11866);
nand U12160 (N_12160,N_11928,N_11963);
xnor U12161 (N_12161,N_11987,N_11842);
or U12162 (N_12162,N_11915,N_11987);
or U12163 (N_12163,N_11911,N_11812);
and U12164 (N_12164,N_11868,N_11919);
and U12165 (N_12165,N_11932,N_11813);
and U12166 (N_12166,N_11977,N_11960);
nand U12167 (N_12167,N_11816,N_11814);
nor U12168 (N_12168,N_11882,N_11880);
nand U12169 (N_12169,N_11904,N_11848);
nor U12170 (N_12170,N_11891,N_11885);
and U12171 (N_12171,N_11878,N_11939);
nand U12172 (N_12172,N_11845,N_11885);
nand U12173 (N_12173,N_11976,N_11814);
nor U12174 (N_12174,N_11814,N_11911);
xnor U12175 (N_12175,N_11977,N_11935);
nor U12176 (N_12176,N_11854,N_11935);
nor U12177 (N_12177,N_11800,N_11813);
or U12178 (N_12178,N_11833,N_11827);
xnor U12179 (N_12179,N_11995,N_11832);
nand U12180 (N_12180,N_11815,N_11932);
and U12181 (N_12181,N_11860,N_11986);
xnor U12182 (N_12182,N_11934,N_11984);
nor U12183 (N_12183,N_11879,N_11990);
or U12184 (N_12184,N_11899,N_11971);
or U12185 (N_12185,N_11887,N_11897);
and U12186 (N_12186,N_11941,N_11932);
xor U12187 (N_12187,N_11982,N_11910);
nand U12188 (N_12188,N_11884,N_11855);
or U12189 (N_12189,N_11906,N_11899);
and U12190 (N_12190,N_11924,N_11893);
xor U12191 (N_12191,N_11818,N_11904);
xor U12192 (N_12192,N_11966,N_11882);
or U12193 (N_12193,N_11800,N_11836);
xnor U12194 (N_12194,N_11973,N_11824);
and U12195 (N_12195,N_11953,N_11894);
xnor U12196 (N_12196,N_11802,N_11946);
nand U12197 (N_12197,N_11933,N_11832);
nor U12198 (N_12198,N_11861,N_11903);
and U12199 (N_12199,N_11962,N_11960);
and U12200 (N_12200,N_12168,N_12117);
and U12201 (N_12201,N_12003,N_12016);
or U12202 (N_12202,N_12010,N_12000);
and U12203 (N_12203,N_12136,N_12163);
nor U12204 (N_12204,N_12082,N_12035);
or U12205 (N_12205,N_12189,N_12126);
or U12206 (N_12206,N_12066,N_12042);
nor U12207 (N_12207,N_12161,N_12172);
nand U12208 (N_12208,N_12080,N_12186);
and U12209 (N_12209,N_12167,N_12093);
nor U12210 (N_12210,N_12132,N_12142);
xor U12211 (N_12211,N_12028,N_12194);
or U12212 (N_12212,N_12155,N_12064);
and U12213 (N_12213,N_12113,N_12158);
nand U12214 (N_12214,N_12012,N_12007);
nand U12215 (N_12215,N_12190,N_12027);
nand U12216 (N_12216,N_12157,N_12149);
nand U12217 (N_12217,N_12191,N_12184);
or U12218 (N_12218,N_12097,N_12051);
xor U12219 (N_12219,N_12101,N_12046);
or U12220 (N_12220,N_12015,N_12160);
or U12221 (N_12221,N_12134,N_12043);
nor U12222 (N_12222,N_12129,N_12078);
or U12223 (N_12223,N_12183,N_12112);
xor U12224 (N_12224,N_12197,N_12063);
nand U12225 (N_12225,N_12122,N_12150);
and U12226 (N_12226,N_12032,N_12029);
nand U12227 (N_12227,N_12009,N_12055);
nor U12228 (N_12228,N_12198,N_12061);
nand U12229 (N_12229,N_12020,N_12094);
and U12230 (N_12230,N_12037,N_12038);
or U12231 (N_12231,N_12090,N_12079);
nand U12232 (N_12232,N_12076,N_12065);
nand U12233 (N_12233,N_12067,N_12119);
and U12234 (N_12234,N_12192,N_12127);
or U12235 (N_12235,N_12060,N_12047);
or U12236 (N_12236,N_12185,N_12144);
xnor U12237 (N_12237,N_12104,N_12008);
xnor U12238 (N_12238,N_12138,N_12092);
nand U12239 (N_12239,N_12024,N_12018);
and U12240 (N_12240,N_12131,N_12011);
nor U12241 (N_12241,N_12114,N_12188);
xnor U12242 (N_12242,N_12033,N_12173);
and U12243 (N_12243,N_12077,N_12199);
xnor U12244 (N_12244,N_12128,N_12026);
nor U12245 (N_12245,N_12048,N_12145);
nor U12246 (N_12246,N_12193,N_12187);
and U12247 (N_12247,N_12105,N_12116);
xor U12248 (N_12248,N_12133,N_12143);
and U12249 (N_12249,N_12195,N_12098);
and U12250 (N_12250,N_12087,N_12130);
xor U12251 (N_12251,N_12156,N_12170);
nand U12252 (N_12252,N_12177,N_12086);
or U12253 (N_12253,N_12071,N_12180);
nand U12254 (N_12254,N_12091,N_12013);
nand U12255 (N_12255,N_12152,N_12106);
or U12256 (N_12256,N_12154,N_12153);
nand U12257 (N_12257,N_12075,N_12006);
and U12258 (N_12258,N_12109,N_12084);
and U12259 (N_12259,N_12021,N_12054);
or U12260 (N_12260,N_12014,N_12118);
and U12261 (N_12261,N_12089,N_12030);
xnor U12262 (N_12262,N_12059,N_12169);
nand U12263 (N_12263,N_12107,N_12081);
nand U12264 (N_12264,N_12120,N_12056);
and U12265 (N_12265,N_12062,N_12110);
nand U12266 (N_12266,N_12031,N_12096);
or U12267 (N_12267,N_12017,N_12135);
nor U12268 (N_12268,N_12068,N_12057);
xor U12269 (N_12269,N_12001,N_12005);
nor U12270 (N_12270,N_12103,N_12179);
nand U12271 (N_12271,N_12019,N_12099);
xnor U12272 (N_12272,N_12023,N_12069);
or U12273 (N_12273,N_12141,N_12052);
or U12274 (N_12274,N_12004,N_12095);
xor U12275 (N_12275,N_12178,N_12159);
xor U12276 (N_12276,N_12088,N_12121);
and U12277 (N_12277,N_12123,N_12111);
nand U12278 (N_12278,N_12050,N_12040);
xor U12279 (N_12279,N_12045,N_12147);
xor U12280 (N_12280,N_12022,N_12025);
and U12281 (N_12281,N_12176,N_12058);
or U12282 (N_12282,N_12181,N_12182);
nor U12283 (N_12283,N_12036,N_12137);
nor U12284 (N_12284,N_12146,N_12151);
nand U12285 (N_12285,N_12102,N_12085);
and U12286 (N_12286,N_12072,N_12074);
xnor U12287 (N_12287,N_12165,N_12164);
or U12288 (N_12288,N_12034,N_12196);
nor U12289 (N_12289,N_12041,N_12139);
nor U12290 (N_12290,N_12166,N_12049);
and U12291 (N_12291,N_12124,N_12175);
nand U12292 (N_12292,N_12174,N_12125);
and U12293 (N_12293,N_12140,N_12108);
xor U12294 (N_12294,N_12070,N_12073);
and U12295 (N_12295,N_12115,N_12039);
nand U12296 (N_12296,N_12171,N_12162);
or U12297 (N_12297,N_12044,N_12148);
nand U12298 (N_12298,N_12053,N_12100);
nand U12299 (N_12299,N_12002,N_12083);
nand U12300 (N_12300,N_12118,N_12096);
nor U12301 (N_12301,N_12067,N_12180);
nor U12302 (N_12302,N_12110,N_12071);
xor U12303 (N_12303,N_12184,N_12088);
or U12304 (N_12304,N_12044,N_12112);
nor U12305 (N_12305,N_12143,N_12086);
or U12306 (N_12306,N_12048,N_12014);
and U12307 (N_12307,N_12141,N_12070);
nand U12308 (N_12308,N_12068,N_12009);
nor U12309 (N_12309,N_12132,N_12072);
or U12310 (N_12310,N_12155,N_12158);
nor U12311 (N_12311,N_12074,N_12174);
nor U12312 (N_12312,N_12106,N_12150);
nand U12313 (N_12313,N_12122,N_12014);
nand U12314 (N_12314,N_12130,N_12142);
and U12315 (N_12315,N_12159,N_12042);
or U12316 (N_12316,N_12011,N_12177);
and U12317 (N_12317,N_12088,N_12104);
xnor U12318 (N_12318,N_12047,N_12089);
nand U12319 (N_12319,N_12167,N_12082);
nand U12320 (N_12320,N_12118,N_12139);
xor U12321 (N_12321,N_12155,N_12122);
and U12322 (N_12322,N_12051,N_12167);
nor U12323 (N_12323,N_12043,N_12180);
and U12324 (N_12324,N_12090,N_12143);
or U12325 (N_12325,N_12122,N_12059);
nor U12326 (N_12326,N_12142,N_12053);
or U12327 (N_12327,N_12101,N_12085);
xnor U12328 (N_12328,N_12163,N_12183);
xnor U12329 (N_12329,N_12052,N_12095);
nor U12330 (N_12330,N_12090,N_12164);
and U12331 (N_12331,N_12064,N_12145);
and U12332 (N_12332,N_12122,N_12113);
nor U12333 (N_12333,N_12197,N_12154);
nand U12334 (N_12334,N_12005,N_12144);
nand U12335 (N_12335,N_12002,N_12006);
xnor U12336 (N_12336,N_12100,N_12047);
and U12337 (N_12337,N_12170,N_12105);
and U12338 (N_12338,N_12197,N_12059);
xnor U12339 (N_12339,N_12123,N_12054);
nor U12340 (N_12340,N_12141,N_12067);
xnor U12341 (N_12341,N_12163,N_12175);
xnor U12342 (N_12342,N_12101,N_12076);
or U12343 (N_12343,N_12069,N_12129);
nand U12344 (N_12344,N_12132,N_12140);
xor U12345 (N_12345,N_12103,N_12101);
or U12346 (N_12346,N_12009,N_12088);
xor U12347 (N_12347,N_12186,N_12032);
nor U12348 (N_12348,N_12193,N_12054);
and U12349 (N_12349,N_12129,N_12038);
xnor U12350 (N_12350,N_12021,N_12128);
xnor U12351 (N_12351,N_12180,N_12162);
and U12352 (N_12352,N_12130,N_12085);
nor U12353 (N_12353,N_12160,N_12132);
nand U12354 (N_12354,N_12015,N_12076);
xor U12355 (N_12355,N_12036,N_12142);
and U12356 (N_12356,N_12152,N_12053);
nor U12357 (N_12357,N_12191,N_12192);
nor U12358 (N_12358,N_12109,N_12044);
xor U12359 (N_12359,N_12066,N_12181);
nand U12360 (N_12360,N_12085,N_12120);
xor U12361 (N_12361,N_12107,N_12161);
xnor U12362 (N_12362,N_12120,N_12139);
nand U12363 (N_12363,N_12140,N_12021);
nand U12364 (N_12364,N_12193,N_12045);
xnor U12365 (N_12365,N_12072,N_12169);
nor U12366 (N_12366,N_12022,N_12008);
and U12367 (N_12367,N_12057,N_12120);
or U12368 (N_12368,N_12053,N_12198);
nand U12369 (N_12369,N_12177,N_12136);
or U12370 (N_12370,N_12035,N_12028);
and U12371 (N_12371,N_12028,N_12178);
nand U12372 (N_12372,N_12030,N_12011);
nand U12373 (N_12373,N_12095,N_12120);
and U12374 (N_12374,N_12041,N_12044);
and U12375 (N_12375,N_12043,N_12155);
nor U12376 (N_12376,N_12070,N_12015);
and U12377 (N_12377,N_12170,N_12196);
or U12378 (N_12378,N_12122,N_12111);
or U12379 (N_12379,N_12120,N_12081);
nor U12380 (N_12380,N_12114,N_12054);
nand U12381 (N_12381,N_12080,N_12044);
nand U12382 (N_12382,N_12006,N_12128);
or U12383 (N_12383,N_12124,N_12061);
or U12384 (N_12384,N_12058,N_12098);
or U12385 (N_12385,N_12124,N_12121);
xor U12386 (N_12386,N_12156,N_12088);
nor U12387 (N_12387,N_12055,N_12023);
xnor U12388 (N_12388,N_12139,N_12062);
xor U12389 (N_12389,N_12096,N_12134);
nand U12390 (N_12390,N_12088,N_12185);
and U12391 (N_12391,N_12074,N_12102);
nor U12392 (N_12392,N_12102,N_12070);
nor U12393 (N_12393,N_12126,N_12042);
nor U12394 (N_12394,N_12152,N_12128);
or U12395 (N_12395,N_12182,N_12024);
nand U12396 (N_12396,N_12191,N_12180);
nor U12397 (N_12397,N_12068,N_12167);
xnor U12398 (N_12398,N_12178,N_12044);
nor U12399 (N_12399,N_12035,N_12093);
nand U12400 (N_12400,N_12342,N_12252);
xor U12401 (N_12401,N_12309,N_12306);
and U12402 (N_12402,N_12301,N_12293);
nand U12403 (N_12403,N_12250,N_12258);
nor U12404 (N_12404,N_12224,N_12275);
xnor U12405 (N_12405,N_12269,N_12251);
nand U12406 (N_12406,N_12282,N_12346);
and U12407 (N_12407,N_12241,N_12383);
and U12408 (N_12408,N_12382,N_12375);
nor U12409 (N_12409,N_12229,N_12392);
xnor U12410 (N_12410,N_12295,N_12374);
xnor U12411 (N_12411,N_12261,N_12298);
xnor U12412 (N_12412,N_12323,N_12368);
nand U12413 (N_12413,N_12276,N_12287);
nor U12414 (N_12414,N_12203,N_12313);
and U12415 (N_12415,N_12249,N_12201);
nor U12416 (N_12416,N_12314,N_12321);
xnor U12417 (N_12417,N_12360,N_12316);
or U12418 (N_12418,N_12359,N_12354);
nand U12419 (N_12419,N_12333,N_12396);
nor U12420 (N_12420,N_12286,N_12345);
and U12421 (N_12421,N_12256,N_12222);
and U12422 (N_12422,N_12334,N_12384);
and U12423 (N_12423,N_12200,N_12253);
xor U12424 (N_12424,N_12364,N_12358);
xor U12425 (N_12425,N_12202,N_12255);
nand U12426 (N_12426,N_12300,N_12219);
xnor U12427 (N_12427,N_12367,N_12355);
xnor U12428 (N_12428,N_12373,N_12296);
or U12429 (N_12429,N_12325,N_12277);
nand U12430 (N_12430,N_12220,N_12370);
or U12431 (N_12431,N_12225,N_12362);
and U12432 (N_12432,N_12240,N_12338);
and U12433 (N_12433,N_12238,N_12239);
and U12434 (N_12434,N_12242,N_12208);
nor U12435 (N_12435,N_12307,N_12218);
nand U12436 (N_12436,N_12206,N_12365);
and U12437 (N_12437,N_12317,N_12343);
xor U12438 (N_12438,N_12221,N_12381);
and U12439 (N_12439,N_12291,N_12347);
xor U12440 (N_12440,N_12337,N_12332);
and U12441 (N_12441,N_12356,N_12284);
nor U12442 (N_12442,N_12312,N_12271);
and U12443 (N_12443,N_12265,N_12273);
nor U12444 (N_12444,N_12243,N_12272);
nor U12445 (N_12445,N_12386,N_12237);
nor U12446 (N_12446,N_12214,N_12246);
and U12447 (N_12447,N_12315,N_12235);
nand U12448 (N_12448,N_12311,N_12213);
nor U12449 (N_12449,N_12394,N_12299);
xnor U12450 (N_12450,N_12232,N_12283);
xor U12451 (N_12451,N_12371,N_12260);
or U12452 (N_12452,N_12245,N_12353);
or U12453 (N_12453,N_12344,N_12230);
or U12454 (N_12454,N_12327,N_12270);
and U12455 (N_12455,N_12376,N_12335);
xor U12456 (N_12456,N_12308,N_12310);
and U12457 (N_12457,N_12331,N_12352);
nor U12458 (N_12458,N_12215,N_12350);
xor U12459 (N_12459,N_12278,N_12209);
nand U12460 (N_12460,N_12378,N_12290);
or U12461 (N_12461,N_12318,N_12330);
xor U12462 (N_12462,N_12336,N_12267);
or U12463 (N_12463,N_12211,N_12379);
nor U12464 (N_12464,N_12259,N_12393);
nand U12465 (N_12465,N_12366,N_12289);
or U12466 (N_12466,N_12385,N_12216);
xnor U12467 (N_12467,N_12341,N_12328);
or U12468 (N_12468,N_12248,N_12390);
nand U12469 (N_12469,N_12326,N_12339);
or U12470 (N_12470,N_12349,N_12263);
nor U12471 (N_12471,N_12304,N_12236);
or U12472 (N_12472,N_12357,N_12377);
xnor U12473 (N_12473,N_12234,N_12207);
nor U12474 (N_12474,N_12247,N_12320);
nand U12475 (N_12475,N_12285,N_12329);
or U12476 (N_12476,N_12305,N_12340);
nor U12477 (N_12477,N_12205,N_12228);
nor U12478 (N_12478,N_12324,N_12369);
xnor U12479 (N_12479,N_12244,N_12303);
or U12480 (N_12480,N_12227,N_12380);
and U12481 (N_12481,N_12372,N_12288);
xor U12482 (N_12482,N_12351,N_12361);
or U12483 (N_12483,N_12231,N_12217);
xnor U12484 (N_12484,N_12348,N_12280);
or U12485 (N_12485,N_12399,N_12257);
nand U12486 (N_12486,N_12281,N_12292);
nand U12487 (N_12487,N_12398,N_12387);
and U12488 (N_12488,N_12388,N_12210);
nand U12489 (N_12489,N_12389,N_12274);
xnor U12490 (N_12490,N_12268,N_12294);
or U12491 (N_12491,N_12204,N_12397);
or U12492 (N_12492,N_12212,N_12223);
xnor U12493 (N_12493,N_12391,N_12264);
xnor U12494 (N_12494,N_12279,N_12262);
nand U12495 (N_12495,N_12266,N_12226);
nor U12496 (N_12496,N_12302,N_12395);
nor U12497 (N_12497,N_12254,N_12363);
nand U12498 (N_12498,N_12297,N_12319);
and U12499 (N_12499,N_12233,N_12322);
and U12500 (N_12500,N_12334,N_12288);
or U12501 (N_12501,N_12291,N_12214);
xnor U12502 (N_12502,N_12342,N_12399);
or U12503 (N_12503,N_12215,N_12341);
nand U12504 (N_12504,N_12292,N_12222);
nor U12505 (N_12505,N_12351,N_12224);
nand U12506 (N_12506,N_12342,N_12236);
or U12507 (N_12507,N_12240,N_12394);
and U12508 (N_12508,N_12240,N_12257);
nor U12509 (N_12509,N_12313,N_12284);
nor U12510 (N_12510,N_12385,N_12224);
or U12511 (N_12511,N_12350,N_12270);
or U12512 (N_12512,N_12280,N_12342);
or U12513 (N_12513,N_12340,N_12291);
xnor U12514 (N_12514,N_12210,N_12339);
nor U12515 (N_12515,N_12204,N_12362);
xor U12516 (N_12516,N_12322,N_12215);
nor U12517 (N_12517,N_12338,N_12344);
xnor U12518 (N_12518,N_12323,N_12356);
nor U12519 (N_12519,N_12304,N_12256);
xor U12520 (N_12520,N_12387,N_12317);
nand U12521 (N_12521,N_12256,N_12303);
and U12522 (N_12522,N_12330,N_12370);
or U12523 (N_12523,N_12314,N_12220);
or U12524 (N_12524,N_12372,N_12305);
xnor U12525 (N_12525,N_12311,N_12350);
and U12526 (N_12526,N_12391,N_12341);
xnor U12527 (N_12527,N_12347,N_12261);
or U12528 (N_12528,N_12313,N_12338);
xnor U12529 (N_12529,N_12259,N_12357);
nand U12530 (N_12530,N_12359,N_12335);
and U12531 (N_12531,N_12261,N_12306);
and U12532 (N_12532,N_12321,N_12210);
or U12533 (N_12533,N_12399,N_12357);
nand U12534 (N_12534,N_12376,N_12301);
nor U12535 (N_12535,N_12348,N_12356);
or U12536 (N_12536,N_12268,N_12288);
or U12537 (N_12537,N_12239,N_12354);
or U12538 (N_12538,N_12382,N_12319);
or U12539 (N_12539,N_12227,N_12213);
nor U12540 (N_12540,N_12385,N_12259);
or U12541 (N_12541,N_12315,N_12294);
nand U12542 (N_12542,N_12235,N_12203);
nand U12543 (N_12543,N_12299,N_12371);
and U12544 (N_12544,N_12330,N_12338);
or U12545 (N_12545,N_12245,N_12396);
nor U12546 (N_12546,N_12233,N_12271);
nor U12547 (N_12547,N_12375,N_12330);
nor U12548 (N_12548,N_12397,N_12317);
nor U12549 (N_12549,N_12355,N_12235);
and U12550 (N_12550,N_12200,N_12288);
and U12551 (N_12551,N_12357,N_12281);
and U12552 (N_12552,N_12245,N_12286);
nand U12553 (N_12553,N_12356,N_12212);
and U12554 (N_12554,N_12310,N_12239);
xor U12555 (N_12555,N_12272,N_12295);
or U12556 (N_12556,N_12375,N_12301);
or U12557 (N_12557,N_12239,N_12300);
and U12558 (N_12558,N_12283,N_12258);
nand U12559 (N_12559,N_12217,N_12304);
and U12560 (N_12560,N_12240,N_12340);
and U12561 (N_12561,N_12285,N_12343);
nand U12562 (N_12562,N_12263,N_12302);
nor U12563 (N_12563,N_12266,N_12373);
and U12564 (N_12564,N_12309,N_12295);
nand U12565 (N_12565,N_12319,N_12367);
nand U12566 (N_12566,N_12329,N_12276);
and U12567 (N_12567,N_12378,N_12357);
xor U12568 (N_12568,N_12214,N_12278);
or U12569 (N_12569,N_12301,N_12230);
nor U12570 (N_12570,N_12390,N_12332);
nor U12571 (N_12571,N_12368,N_12232);
or U12572 (N_12572,N_12354,N_12209);
and U12573 (N_12573,N_12340,N_12277);
nand U12574 (N_12574,N_12258,N_12387);
and U12575 (N_12575,N_12318,N_12362);
xor U12576 (N_12576,N_12350,N_12321);
or U12577 (N_12577,N_12268,N_12202);
nor U12578 (N_12578,N_12309,N_12399);
and U12579 (N_12579,N_12367,N_12364);
or U12580 (N_12580,N_12311,N_12293);
nand U12581 (N_12581,N_12340,N_12268);
nand U12582 (N_12582,N_12358,N_12215);
xnor U12583 (N_12583,N_12368,N_12259);
nand U12584 (N_12584,N_12344,N_12220);
nand U12585 (N_12585,N_12336,N_12298);
nor U12586 (N_12586,N_12368,N_12216);
nand U12587 (N_12587,N_12373,N_12387);
xnor U12588 (N_12588,N_12253,N_12229);
nor U12589 (N_12589,N_12243,N_12325);
nand U12590 (N_12590,N_12338,N_12304);
nand U12591 (N_12591,N_12345,N_12240);
nor U12592 (N_12592,N_12358,N_12283);
xor U12593 (N_12593,N_12204,N_12375);
and U12594 (N_12594,N_12389,N_12343);
nor U12595 (N_12595,N_12224,N_12226);
or U12596 (N_12596,N_12381,N_12306);
or U12597 (N_12597,N_12210,N_12289);
or U12598 (N_12598,N_12308,N_12265);
or U12599 (N_12599,N_12200,N_12314);
or U12600 (N_12600,N_12493,N_12439);
or U12601 (N_12601,N_12558,N_12413);
nor U12602 (N_12602,N_12543,N_12504);
or U12603 (N_12603,N_12408,N_12488);
xnor U12604 (N_12604,N_12464,N_12564);
or U12605 (N_12605,N_12553,N_12497);
nand U12606 (N_12606,N_12457,N_12409);
nand U12607 (N_12607,N_12563,N_12523);
or U12608 (N_12608,N_12438,N_12516);
nand U12609 (N_12609,N_12566,N_12572);
nand U12610 (N_12610,N_12425,N_12557);
nand U12611 (N_12611,N_12471,N_12552);
nand U12612 (N_12612,N_12437,N_12595);
nor U12613 (N_12613,N_12580,N_12594);
nand U12614 (N_12614,N_12578,N_12562);
or U12615 (N_12615,N_12401,N_12421);
nand U12616 (N_12616,N_12524,N_12577);
xnor U12617 (N_12617,N_12522,N_12585);
or U12618 (N_12618,N_12546,N_12508);
nand U12619 (N_12619,N_12427,N_12515);
nor U12620 (N_12620,N_12452,N_12486);
xnor U12621 (N_12621,N_12410,N_12416);
xnor U12622 (N_12622,N_12473,N_12591);
nand U12623 (N_12623,N_12514,N_12529);
xor U12624 (N_12624,N_12411,N_12592);
or U12625 (N_12625,N_12412,N_12554);
nor U12626 (N_12626,N_12598,N_12590);
nand U12627 (N_12627,N_12478,N_12474);
nand U12628 (N_12628,N_12458,N_12510);
or U12629 (N_12629,N_12431,N_12426);
or U12630 (N_12630,N_12480,N_12432);
or U12631 (N_12631,N_12537,N_12544);
or U12632 (N_12632,N_12453,N_12476);
nor U12633 (N_12633,N_12555,N_12404);
xnor U12634 (N_12634,N_12593,N_12501);
nand U12635 (N_12635,N_12527,N_12455);
or U12636 (N_12636,N_12534,N_12467);
or U12637 (N_12637,N_12550,N_12433);
nand U12638 (N_12638,N_12539,N_12491);
nand U12639 (N_12639,N_12519,N_12528);
nand U12640 (N_12640,N_12587,N_12445);
nor U12641 (N_12641,N_12570,N_12436);
nor U12642 (N_12642,N_12469,N_12470);
and U12643 (N_12643,N_12406,N_12463);
and U12644 (N_12644,N_12481,N_12441);
or U12645 (N_12645,N_12400,N_12582);
nor U12646 (N_12646,N_12583,N_12547);
xnor U12647 (N_12647,N_12414,N_12540);
and U12648 (N_12648,N_12442,N_12509);
nor U12649 (N_12649,N_12517,N_12456);
xor U12650 (N_12650,N_12494,N_12448);
and U12651 (N_12651,N_12446,N_12521);
and U12652 (N_12652,N_12533,N_12477);
xor U12653 (N_12653,N_12506,N_12512);
xnor U12654 (N_12654,N_12405,N_12454);
xor U12655 (N_12655,N_12444,N_12526);
and U12656 (N_12656,N_12475,N_12556);
xnor U12657 (N_12657,N_12451,N_12472);
and U12658 (N_12658,N_12545,N_12489);
xor U12659 (N_12659,N_12490,N_12576);
and U12660 (N_12660,N_12492,N_12468);
nor U12661 (N_12661,N_12485,N_12466);
or U12662 (N_12662,N_12597,N_12505);
nand U12663 (N_12663,N_12599,N_12483);
xnor U12664 (N_12664,N_12541,N_12429);
and U12665 (N_12665,N_12465,N_12417);
and U12666 (N_12666,N_12542,N_12575);
xnor U12667 (N_12667,N_12443,N_12571);
or U12668 (N_12668,N_12484,N_12422);
xnor U12669 (N_12669,N_12459,N_12503);
xnor U12670 (N_12670,N_12535,N_12507);
nor U12671 (N_12671,N_12407,N_12532);
and U12672 (N_12672,N_12435,N_12415);
or U12673 (N_12673,N_12551,N_12513);
nand U12674 (N_12674,N_12420,N_12560);
xor U12675 (N_12675,N_12447,N_12581);
nand U12676 (N_12676,N_12561,N_12482);
nor U12677 (N_12677,N_12428,N_12536);
and U12678 (N_12678,N_12525,N_12487);
nor U12679 (N_12679,N_12434,N_12530);
nor U12680 (N_12680,N_12419,N_12567);
or U12681 (N_12681,N_12462,N_12449);
and U12682 (N_12682,N_12548,N_12520);
nor U12683 (N_12683,N_12402,N_12579);
nor U12684 (N_12684,N_12568,N_12403);
and U12685 (N_12685,N_12518,N_12461);
or U12686 (N_12686,N_12496,N_12589);
xnor U12687 (N_12687,N_12596,N_12498);
nor U12688 (N_12688,N_12418,N_12573);
or U12689 (N_12689,N_12588,N_12499);
nand U12690 (N_12690,N_12565,N_12559);
nor U12691 (N_12691,N_12538,N_12430);
nor U12692 (N_12692,N_12423,N_12460);
or U12693 (N_12693,N_12586,N_12502);
or U12694 (N_12694,N_12479,N_12574);
or U12695 (N_12695,N_12584,N_12495);
nor U12696 (N_12696,N_12424,N_12531);
and U12697 (N_12697,N_12569,N_12500);
xnor U12698 (N_12698,N_12511,N_12440);
nand U12699 (N_12699,N_12450,N_12549);
nand U12700 (N_12700,N_12572,N_12537);
nor U12701 (N_12701,N_12531,N_12436);
or U12702 (N_12702,N_12467,N_12414);
nand U12703 (N_12703,N_12552,N_12492);
xnor U12704 (N_12704,N_12524,N_12579);
xor U12705 (N_12705,N_12496,N_12401);
and U12706 (N_12706,N_12486,N_12550);
or U12707 (N_12707,N_12447,N_12549);
nand U12708 (N_12708,N_12459,N_12507);
xor U12709 (N_12709,N_12462,N_12456);
and U12710 (N_12710,N_12482,N_12589);
or U12711 (N_12711,N_12490,N_12434);
and U12712 (N_12712,N_12536,N_12438);
or U12713 (N_12713,N_12536,N_12576);
and U12714 (N_12714,N_12485,N_12486);
xnor U12715 (N_12715,N_12544,N_12431);
and U12716 (N_12716,N_12566,N_12487);
or U12717 (N_12717,N_12588,N_12440);
nor U12718 (N_12718,N_12547,N_12593);
or U12719 (N_12719,N_12522,N_12567);
or U12720 (N_12720,N_12532,N_12421);
xnor U12721 (N_12721,N_12453,N_12528);
nand U12722 (N_12722,N_12426,N_12416);
xor U12723 (N_12723,N_12497,N_12545);
and U12724 (N_12724,N_12521,N_12414);
nor U12725 (N_12725,N_12420,N_12417);
or U12726 (N_12726,N_12477,N_12404);
xor U12727 (N_12727,N_12586,N_12531);
and U12728 (N_12728,N_12598,N_12550);
and U12729 (N_12729,N_12568,N_12417);
or U12730 (N_12730,N_12437,N_12579);
or U12731 (N_12731,N_12579,N_12442);
nor U12732 (N_12732,N_12533,N_12514);
or U12733 (N_12733,N_12527,N_12481);
and U12734 (N_12734,N_12584,N_12494);
or U12735 (N_12735,N_12466,N_12576);
nand U12736 (N_12736,N_12599,N_12487);
or U12737 (N_12737,N_12425,N_12457);
or U12738 (N_12738,N_12439,N_12556);
nand U12739 (N_12739,N_12551,N_12524);
and U12740 (N_12740,N_12595,N_12583);
and U12741 (N_12741,N_12578,N_12549);
or U12742 (N_12742,N_12560,N_12575);
and U12743 (N_12743,N_12426,N_12494);
nand U12744 (N_12744,N_12570,N_12401);
or U12745 (N_12745,N_12541,N_12454);
and U12746 (N_12746,N_12537,N_12564);
or U12747 (N_12747,N_12541,N_12508);
and U12748 (N_12748,N_12437,N_12499);
or U12749 (N_12749,N_12558,N_12496);
or U12750 (N_12750,N_12498,N_12494);
or U12751 (N_12751,N_12596,N_12546);
or U12752 (N_12752,N_12570,N_12542);
or U12753 (N_12753,N_12407,N_12537);
nor U12754 (N_12754,N_12490,N_12458);
nand U12755 (N_12755,N_12598,N_12440);
nor U12756 (N_12756,N_12489,N_12498);
or U12757 (N_12757,N_12572,N_12420);
nand U12758 (N_12758,N_12435,N_12479);
and U12759 (N_12759,N_12413,N_12564);
nor U12760 (N_12760,N_12433,N_12517);
nand U12761 (N_12761,N_12595,N_12556);
xnor U12762 (N_12762,N_12431,N_12400);
xor U12763 (N_12763,N_12487,N_12513);
or U12764 (N_12764,N_12556,N_12441);
nand U12765 (N_12765,N_12521,N_12403);
nor U12766 (N_12766,N_12508,N_12536);
nor U12767 (N_12767,N_12436,N_12580);
nor U12768 (N_12768,N_12532,N_12448);
nand U12769 (N_12769,N_12467,N_12579);
and U12770 (N_12770,N_12498,N_12591);
or U12771 (N_12771,N_12450,N_12418);
and U12772 (N_12772,N_12440,N_12537);
nand U12773 (N_12773,N_12527,N_12511);
and U12774 (N_12774,N_12558,N_12545);
nand U12775 (N_12775,N_12416,N_12477);
xor U12776 (N_12776,N_12588,N_12472);
or U12777 (N_12777,N_12590,N_12523);
and U12778 (N_12778,N_12464,N_12475);
nand U12779 (N_12779,N_12522,N_12410);
nor U12780 (N_12780,N_12475,N_12522);
xnor U12781 (N_12781,N_12487,N_12508);
nand U12782 (N_12782,N_12563,N_12525);
or U12783 (N_12783,N_12440,N_12412);
and U12784 (N_12784,N_12560,N_12569);
nor U12785 (N_12785,N_12438,N_12532);
and U12786 (N_12786,N_12467,N_12410);
nor U12787 (N_12787,N_12441,N_12462);
or U12788 (N_12788,N_12421,N_12490);
xnor U12789 (N_12789,N_12419,N_12539);
or U12790 (N_12790,N_12539,N_12478);
and U12791 (N_12791,N_12526,N_12403);
xor U12792 (N_12792,N_12421,N_12437);
nor U12793 (N_12793,N_12593,N_12583);
nand U12794 (N_12794,N_12456,N_12563);
xor U12795 (N_12795,N_12475,N_12413);
and U12796 (N_12796,N_12573,N_12508);
nand U12797 (N_12797,N_12466,N_12436);
nor U12798 (N_12798,N_12462,N_12508);
nand U12799 (N_12799,N_12490,N_12562);
nand U12800 (N_12800,N_12633,N_12611);
xor U12801 (N_12801,N_12773,N_12610);
nor U12802 (N_12802,N_12718,N_12690);
nor U12803 (N_12803,N_12758,N_12609);
or U12804 (N_12804,N_12641,N_12664);
nor U12805 (N_12805,N_12646,N_12766);
xnor U12806 (N_12806,N_12696,N_12793);
xor U12807 (N_12807,N_12782,N_12765);
nand U12808 (N_12808,N_12635,N_12704);
or U12809 (N_12809,N_12666,N_12791);
or U12810 (N_12810,N_12686,N_12768);
nand U12811 (N_12811,N_12654,N_12778);
nor U12812 (N_12812,N_12628,N_12668);
nand U12813 (N_12813,N_12781,N_12753);
xnor U12814 (N_12814,N_12794,N_12630);
or U12815 (N_12815,N_12740,N_12614);
xor U12816 (N_12816,N_12680,N_12745);
nand U12817 (N_12817,N_12669,N_12706);
xnor U12818 (N_12818,N_12601,N_12695);
nor U12819 (N_12819,N_12678,N_12729);
xor U12820 (N_12820,N_12709,N_12776);
nand U12821 (N_12821,N_12600,N_12651);
or U12822 (N_12822,N_12632,N_12667);
and U12823 (N_12823,N_12629,N_12619);
nor U12824 (N_12824,N_12756,N_12659);
and U12825 (N_12825,N_12688,N_12725);
and U12826 (N_12826,N_12606,N_12790);
nor U12827 (N_12827,N_12604,N_12760);
and U12828 (N_12828,N_12750,N_12770);
xnor U12829 (N_12829,N_12780,N_12661);
and U12830 (N_12830,N_12761,N_12707);
nand U12831 (N_12831,N_12692,N_12764);
and U12832 (N_12832,N_12620,N_12603);
nor U12833 (N_12833,N_12639,N_12700);
nand U12834 (N_12834,N_12728,N_12674);
nand U12835 (N_12835,N_12703,N_12712);
nor U12836 (N_12836,N_12784,N_12657);
or U12837 (N_12837,N_12687,N_12705);
nor U12838 (N_12838,N_12751,N_12731);
and U12839 (N_12839,N_12749,N_12658);
nor U12840 (N_12840,N_12681,N_12638);
and U12841 (N_12841,N_12757,N_12612);
or U12842 (N_12842,N_12671,N_12733);
or U12843 (N_12843,N_12792,N_12735);
xnor U12844 (N_12844,N_12679,N_12631);
xnor U12845 (N_12845,N_12755,N_12789);
xor U12846 (N_12846,N_12787,N_12713);
xor U12847 (N_12847,N_12724,N_12741);
or U12848 (N_12848,N_12621,N_12702);
and U12849 (N_12849,N_12672,N_12662);
nor U12850 (N_12850,N_12650,N_12767);
and U12851 (N_12851,N_12626,N_12783);
nor U12852 (N_12852,N_12618,N_12625);
and U12853 (N_12853,N_12649,N_12798);
or U12854 (N_12854,N_12608,N_12648);
or U12855 (N_12855,N_12653,N_12786);
nor U12856 (N_12856,N_12747,N_12655);
or U12857 (N_12857,N_12665,N_12605);
and U12858 (N_12858,N_12615,N_12613);
xor U12859 (N_12859,N_12683,N_12742);
xor U12860 (N_12860,N_12624,N_12645);
nand U12861 (N_12861,N_12797,N_12698);
or U12862 (N_12862,N_12723,N_12737);
nand U12863 (N_12863,N_12714,N_12616);
xnor U12864 (N_12864,N_12701,N_12720);
or U12865 (N_12865,N_12732,N_12799);
nor U12866 (N_12866,N_12697,N_12677);
or U12867 (N_12867,N_12711,N_12746);
or U12868 (N_12868,N_12779,N_12642);
nand U12869 (N_12869,N_12673,N_12736);
or U12870 (N_12870,N_12663,N_12644);
or U12871 (N_12871,N_12694,N_12689);
xor U12872 (N_12872,N_12777,N_12656);
and U12873 (N_12873,N_12623,N_12684);
nor U12874 (N_12874,N_12717,N_12785);
and U12875 (N_12875,N_12774,N_12676);
nor U12876 (N_12876,N_12795,N_12738);
nand U12877 (N_12877,N_12772,N_12739);
nand U12878 (N_12878,N_12759,N_12754);
nor U12879 (N_12879,N_12652,N_12775);
nor U12880 (N_12880,N_12607,N_12762);
or U12881 (N_12881,N_12637,N_12643);
nor U12882 (N_12882,N_12685,N_12716);
nor U12883 (N_12883,N_12675,N_12743);
and U12884 (N_12884,N_12682,N_12660);
and U12885 (N_12885,N_12730,N_12691);
nand U12886 (N_12886,N_12771,N_12788);
xnor U12887 (N_12887,N_12710,N_12721);
nand U12888 (N_12888,N_12670,N_12715);
nand U12889 (N_12889,N_12752,N_12726);
or U12890 (N_12890,N_12693,N_12734);
or U12891 (N_12891,N_12708,N_12722);
and U12892 (N_12892,N_12622,N_12719);
and U12893 (N_12893,N_12796,N_12727);
and U12894 (N_12894,N_12617,N_12647);
nor U12895 (N_12895,N_12627,N_12634);
and U12896 (N_12896,N_12699,N_12636);
nor U12897 (N_12897,N_12769,N_12602);
nand U12898 (N_12898,N_12763,N_12640);
and U12899 (N_12899,N_12748,N_12744);
and U12900 (N_12900,N_12711,N_12663);
nor U12901 (N_12901,N_12756,N_12623);
nand U12902 (N_12902,N_12689,N_12676);
or U12903 (N_12903,N_12771,N_12631);
xor U12904 (N_12904,N_12608,N_12668);
nor U12905 (N_12905,N_12759,N_12693);
or U12906 (N_12906,N_12637,N_12651);
or U12907 (N_12907,N_12799,N_12648);
and U12908 (N_12908,N_12635,N_12634);
nand U12909 (N_12909,N_12613,N_12711);
nor U12910 (N_12910,N_12678,N_12602);
or U12911 (N_12911,N_12645,N_12639);
xor U12912 (N_12912,N_12716,N_12726);
xor U12913 (N_12913,N_12736,N_12757);
or U12914 (N_12914,N_12765,N_12797);
nor U12915 (N_12915,N_12607,N_12796);
nand U12916 (N_12916,N_12723,N_12646);
or U12917 (N_12917,N_12763,N_12785);
nand U12918 (N_12918,N_12647,N_12650);
nor U12919 (N_12919,N_12659,N_12673);
and U12920 (N_12920,N_12653,N_12678);
nand U12921 (N_12921,N_12636,N_12739);
or U12922 (N_12922,N_12652,N_12740);
nand U12923 (N_12923,N_12706,N_12683);
and U12924 (N_12924,N_12795,N_12791);
or U12925 (N_12925,N_12793,N_12689);
and U12926 (N_12926,N_12762,N_12638);
xor U12927 (N_12927,N_12625,N_12609);
and U12928 (N_12928,N_12600,N_12761);
xor U12929 (N_12929,N_12620,N_12637);
and U12930 (N_12930,N_12772,N_12798);
nor U12931 (N_12931,N_12765,N_12710);
and U12932 (N_12932,N_12739,N_12684);
nor U12933 (N_12933,N_12796,N_12783);
and U12934 (N_12934,N_12668,N_12679);
nor U12935 (N_12935,N_12738,N_12719);
nand U12936 (N_12936,N_12745,N_12640);
or U12937 (N_12937,N_12737,N_12682);
nor U12938 (N_12938,N_12790,N_12672);
xnor U12939 (N_12939,N_12657,N_12727);
and U12940 (N_12940,N_12661,N_12769);
or U12941 (N_12941,N_12723,N_12627);
and U12942 (N_12942,N_12724,N_12745);
nand U12943 (N_12943,N_12738,N_12665);
xnor U12944 (N_12944,N_12781,N_12793);
nor U12945 (N_12945,N_12730,N_12646);
nand U12946 (N_12946,N_12612,N_12712);
nor U12947 (N_12947,N_12602,N_12661);
and U12948 (N_12948,N_12632,N_12612);
and U12949 (N_12949,N_12773,N_12672);
xnor U12950 (N_12950,N_12695,N_12720);
nand U12951 (N_12951,N_12777,N_12601);
or U12952 (N_12952,N_12728,N_12696);
xnor U12953 (N_12953,N_12775,N_12751);
nand U12954 (N_12954,N_12733,N_12635);
nor U12955 (N_12955,N_12785,N_12602);
and U12956 (N_12956,N_12678,N_12739);
xnor U12957 (N_12957,N_12735,N_12758);
nand U12958 (N_12958,N_12603,N_12674);
nand U12959 (N_12959,N_12682,N_12715);
nor U12960 (N_12960,N_12696,N_12638);
and U12961 (N_12961,N_12776,N_12674);
xnor U12962 (N_12962,N_12629,N_12758);
and U12963 (N_12963,N_12735,N_12695);
nand U12964 (N_12964,N_12628,N_12680);
nand U12965 (N_12965,N_12746,N_12785);
or U12966 (N_12966,N_12777,N_12708);
nor U12967 (N_12967,N_12657,N_12643);
or U12968 (N_12968,N_12795,N_12743);
and U12969 (N_12969,N_12625,N_12795);
xor U12970 (N_12970,N_12696,N_12764);
or U12971 (N_12971,N_12645,N_12700);
or U12972 (N_12972,N_12606,N_12781);
nand U12973 (N_12973,N_12604,N_12717);
nor U12974 (N_12974,N_12710,N_12770);
and U12975 (N_12975,N_12623,N_12649);
xnor U12976 (N_12976,N_12650,N_12758);
xnor U12977 (N_12977,N_12607,N_12653);
nand U12978 (N_12978,N_12735,N_12713);
nor U12979 (N_12979,N_12741,N_12627);
nand U12980 (N_12980,N_12612,N_12798);
or U12981 (N_12981,N_12775,N_12778);
xnor U12982 (N_12982,N_12630,N_12707);
and U12983 (N_12983,N_12634,N_12784);
xor U12984 (N_12984,N_12655,N_12767);
or U12985 (N_12985,N_12691,N_12782);
nand U12986 (N_12986,N_12725,N_12785);
nand U12987 (N_12987,N_12732,N_12722);
or U12988 (N_12988,N_12673,N_12671);
nor U12989 (N_12989,N_12710,N_12796);
or U12990 (N_12990,N_12770,N_12790);
and U12991 (N_12991,N_12762,N_12703);
nor U12992 (N_12992,N_12629,N_12774);
xor U12993 (N_12993,N_12717,N_12732);
and U12994 (N_12994,N_12641,N_12673);
or U12995 (N_12995,N_12792,N_12720);
xor U12996 (N_12996,N_12773,N_12731);
nand U12997 (N_12997,N_12739,N_12641);
nand U12998 (N_12998,N_12657,N_12630);
nand U12999 (N_12999,N_12672,N_12715);
or U13000 (N_13000,N_12939,N_12996);
or U13001 (N_13001,N_12918,N_12800);
or U13002 (N_13002,N_12861,N_12898);
and U13003 (N_13003,N_12862,N_12826);
nor U13004 (N_13004,N_12936,N_12959);
and U13005 (N_13005,N_12889,N_12969);
nand U13006 (N_13006,N_12967,N_12841);
nor U13007 (N_13007,N_12986,N_12827);
or U13008 (N_13008,N_12966,N_12821);
and U13009 (N_13009,N_12857,N_12883);
and U13010 (N_13010,N_12946,N_12956);
nand U13011 (N_13011,N_12984,N_12963);
nor U13012 (N_13012,N_12972,N_12863);
nand U13013 (N_13013,N_12887,N_12845);
and U13014 (N_13014,N_12839,N_12854);
xor U13015 (N_13015,N_12948,N_12825);
nor U13016 (N_13016,N_12869,N_12823);
and U13017 (N_13017,N_12953,N_12893);
nand U13018 (N_13018,N_12904,N_12961);
or U13019 (N_13019,N_12916,N_12924);
or U13020 (N_13020,N_12885,N_12962);
xor U13021 (N_13021,N_12960,N_12949);
or U13022 (N_13022,N_12835,N_12899);
xnor U13023 (N_13023,N_12818,N_12850);
nor U13024 (N_13024,N_12968,N_12942);
or U13025 (N_13025,N_12927,N_12994);
or U13026 (N_13026,N_12832,N_12859);
nor U13027 (N_13027,N_12941,N_12804);
xor U13028 (N_13028,N_12932,N_12888);
and U13029 (N_13029,N_12999,N_12910);
xor U13030 (N_13030,N_12976,N_12983);
xor U13031 (N_13031,N_12938,N_12882);
nor U13032 (N_13032,N_12914,N_12877);
or U13033 (N_13033,N_12834,N_12803);
and U13034 (N_13034,N_12971,N_12801);
or U13035 (N_13035,N_12843,N_12846);
or U13036 (N_13036,N_12987,N_12828);
and U13037 (N_13037,N_12940,N_12920);
nand U13038 (N_13038,N_12922,N_12952);
nand U13039 (N_13039,N_12802,N_12809);
or U13040 (N_13040,N_12830,N_12909);
nor U13041 (N_13041,N_12937,N_12955);
or U13042 (N_13042,N_12903,N_12997);
or U13043 (N_13043,N_12964,N_12917);
xor U13044 (N_13044,N_12831,N_12868);
and U13045 (N_13045,N_12853,N_12896);
xor U13046 (N_13046,N_12891,N_12978);
or U13047 (N_13047,N_12934,N_12926);
nor U13048 (N_13048,N_12897,N_12833);
nand U13049 (N_13049,N_12816,N_12973);
nor U13050 (N_13050,N_12923,N_12880);
nor U13051 (N_13051,N_12944,N_12858);
and U13052 (N_13052,N_12847,N_12866);
nand U13053 (N_13053,N_12931,N_12849);
or U13054 (N_13054,N_12989,N_12954);
and U13055 (N_13055,N_12945,N_12811);
nand U13056 (N_13056,N_12873,N_12837);
nand U13057 (N_13057,N_12865,N_12958);
xnor U13058 (N_13058,N_12982,N_12894);
or U13059 (N_13059,N_12881,N_12814);
or U13060 (N_13060,N_12965,N_12806);
nand U13061 (N_13061,N_12810,N_12950);
xor U13062 (N_13062,N_12840,N_12870);
nor U13063 (N_13063,N_12879,N_12844);
xor U13064 (N_13064,N_12943,N_12975);
nor U13065 (N_13065,N_12933,N_12848);
and U13066 (N_13066,N_12842,N_12928);
or U13067 (N_13067,N_12895,N_12991);
xor U13068 (N_13068,N_12892,N_12957);
xnor U13069 (N_13069,N_12988,N_12929);
and U13070 (N_13070,N_12981,N_12979);
nand U13071 (N_13071,N_12815,N_12808);
xnor U13072 (N_13072,N_12992,N_12915);
or U13073 (N_13073,N_12817,N_12913);
nand U13074 (N_13074,N_12900,N_12947);
nand U13075 (N_13075,N_12890,N_12860);
xnor U13076 (N_13076,N_12902,N_12875);
or U13077 (N_13077,N_12820,N_12985);
xnor U13078 (N_13078,N_12867,N_12930);
and U13079 (N_13079,N_12886,N_12919);
and U13080 (N_13080,N_12977,N_12876);
xnor U13081 (N_13081,N_12874,N_12824);
and U13082 (N_13082,N_12912,N_12878);
nand U13083 (N_13083,N_12907,N_12884);
nand U13084 (N_13084,N_12905,N_12813);
or U13085 (N_13085,N_12871,N_12911);
nand U13086 (N_13086,N_12864,N_12995);
nor U13087 (N_13087,N_12993,N_12851);
nand U13088 (N_13088,N_12855,N_12807);
nand U13089 (N_13089,N_12990,N_12901);
nor U13090 (N_13090,N_12856,N_12838);
xor U13091 (N_13091,N_12980,N_12935);
and U13092 (N_13092,N_12970,N_12998);
and U13093 (N_13093,N_12829,N_12908);
nor U13094 (N_13094,N_12872,N_12852);
nand U13095 (N_13095,N_12822,N_12925);
xor U13096 (N_13096,N_12812,N_12836);
nor U13097 (N_13097,N_12906,N_12819);
or U13098 (N_13098,N_12921,N_12951);
nor U13099 (N_13099,N_12974,N_12805);
nor U13100 (N_13100,N_12983,N_12910);
nor U13101 (N_13101,N_12838,N_12960);
or U13102 (N_13102,N_12892,N_12955);
xnor U13103 (N_13103,N_12808,N_12975);
and U13104 (N_13104,N_12896,N_12878);
or U13105 (N_13105,N_12832,N_12875);
nand U13106 (N_13106,N_12830,N_12943);
xnor U13107 (N_13107,N_12962,N_12851);
nand U13108 (N_13108,N_12806,N_12856);
nor U13109 (N_13109,N_12949,N_12983);
and U13110 (N_13110,N_12824,N_12891);
or U13111 (N_13111,N_12936,N_12985);
or U13112 (N_13112,N_12948,N_12942);
nand U13113 (N_13113,N_12897,N_12857);
or U13114 (N_13114,N_12901,N_12866);
and U13115 (N_13115,N_12997,N_12902);
or U13116 (N_13116,N_12929,N_12832);
and U13117 (N_13117,N_12950,N_12983);
nor U13118 (N_13118,N_12945,N_12952);
nor U13119 (N_13119,N_12966,N_12867);
nor U13120 (N_13120,N_12860,N_12939);
xor U13121 (N_13121,N_12838,N_12878);
and U13122 (N_13122,N_12950,N_12825);
nor U13123 (N_13123,N_12876,N_12923);
and U13124 (N_13124,N_12821,N_12998);
or U13125 (N_13125,N_12861,N_12987);
xor U13126 (N_13126,N_12921,N_12820);
nor U13127 (N_13127,N_12892,N_12876);
nand U13128 (N_13128,N_12984,N_12891);
nand U13129 (N_13129,N_12857,N_12971);
nor U13130 (N_13130,N_12803,N_12899);
or U13131 (N_13131,N_12902,N_12927);
and U13132 (N_13132,N_12989,N_12857);
xnor U13133 (N_13133,N_12943,N_12974);
nand U13134 (N_13134,N_12872,N_12858);
and U13135 (N_13135,N_12912,N_12815);
or U13136 (N_13136,N_12924,N_12849);
nor U13137 (N_13137,N_12977,N_12887);
nand U13138 (N_13138,N_12926,N_12807);
and U13139 (N_13139,N_12800,N_12915);
xnor U13140 (N_13140,N_12816,N_12883);
and U13141 (N_13141,N_12869,N_12856);
nor U13142 (N_13142,N_12806,N_12932);
nor U13143 (N_13143,N_12888,N_12835);
nor U13144 (N_13144,N_12876,N_12859);
nor U13145 (N_13145,N_12897,N_12893);
xor U13146 (N_13146,N_12986,N_12907);
and U13147 (N_13147,N_12982,N_12960);
xnor U13148 (N_13148,N_12904,N_12840);
and U13149 (N_13149,N_12942,N_12901);
and U13150 (N_13150,N_12852,N_12815);
nand U13151 (N_13151,N_12871,N_12805);
nand U13152 (N_13152,N_12947,N_12971);
and U13153 (N_13153,N_12910,N_12878);
or U13154 (N_13154,N_12914,N_12818);
and U13155 (N_13155,N_12840,N_12964);
nor U13156 (N_13156,N_12967,N_12932);
or U13157 (N_13157,N_12871,N_12989);
or U13158 (N_13158,N_12830,N_12896);
or U13159 (N_13159,N_12937,N_12817);
nand U13160 (N_13160,N_12943,N_12961);
and U13161 (N_13161,N_12983,N_12815);
or U13162 (N_13162,N_12992,N_12822);
xor U13163 (N_13163,N_12812,N_12994);
xor U13164 (N_13164,N_12957,N_12970);
or U13165 (N_13165,N_12878,N_12925);
xor U13166 (N_13166,N_12881,N_12940);
or U13167 (N_13167,N_12841,N_12905);
and U13168 (N_13168,N_12901,N_12921);
and U13169 (N_13169,N_12979,N_12846);
xnor U13170 (N_13170,N_12901,N_12884);
nand U13171 (N_13171,N_12809,N_12855);
and U13172 (N_13172,N_12919,N_12943);
or U13173 (N_13173,N_12846,N_12919);
nor U13174 (N_13174,N_12837,N_12834);
nand U13175 (N_13175,N_12952,N_12909);
nor U13176 (N_13176,N_12839,N_12862);
nand U13177 (N_13177,N_12808,N_12962);
and U13178 (N_13178,N_12885,N_12920);
or U13179 (N_13179,N_12875,N_12992);
and U13180 (N_13180,N_12909,N_12919);
or U13181 (N_13181,N_12872,N_12916);
nor U13182 (N_13182,N_12870,N_12811);
and U13183 (N_13183,N_12905,N_12864);
nor U13184 (N_13184,N_12967,N_12933);
and U13185 (N_13185,N_12995,N_12990);
nand U13186 (N_13186,N_12930,N_12917);
and U13187 (N_13187,N_12990,N_12973);
nand U13188 (N_13188,N_12902,N_12973);
and U13189 (N_13189,N_12875,N_12912);
xor U13190 (N_13190,N_12934,N_12992);
nor U13191 (N_13191,N_12864,N_12993);
or U13192 (N_13192,N_12962,N_12837);
xor U13193 (N_13193,N_12901,N_12952);
nor U13194 (N_13194,N_12865,N_12815);
nor U13195 (N_13195,N_12800,N_12927);
or U13196 (N_13196,N_12943,N_12840);
and U13197 (N_13197,N_12988,N_12903);
xor U13198 (N_13198,N_12823,N_12877);
nor U13199 (N_13199,N_12946,N_12820);
nand U13200 (N_13200,N_13109,N_13196);
nand U13201 (N_13201,N_13115,N_13172);
nand U13202 (N_13202,N_13170,N_13079);
and U13203 (N_13203,N_13005,N_13125);
or U13204 (N_13204,N_13039,N_13015);
and U13205 (N_13205,N_13001,N_13089);
or U13206 (N_13206,N_13037,N_13138);
nor U13207 (N_13207,N_13038,N_13028);
nor U13208 (N_13208,N_13073,N_13169);
and U13209 (N_13209,N_13076,N_13108);
xor U13210 (N_13210,N_13052,N_13097);
xnor U13211 (N_13211,N_13116,N_13021);
nor U13212 (N_13212,N_13103,N_13132);
or U13213 (N_13213,N_13189,N_13093);
nor U13214 (N_13214,N_13051,N_13153);
or U13215 (N_13215,N_13091,N_13130);
nor U13216 (N_13216,N_13148,N_13023);
and U13217 (N_13217,N_13110,N_13107);
xnor U13218 (N_13218,N_13111,N_13141);
nor U13219 (N_13219,N_13187,N_13128);
or U13220 (N_13220,N_13029,N_13086);
nor U13221 (N_13221,N_13166,N_13071);
nand U13222 (N_13222,N_13040,N_13085);
nor U13223 (N_13223,N_13198,N_13106);
nor U13224 (N_13224,N_13178,N_13131);
nor U13225 (N_13225,N_13161,N_13041);
xnor U13226 (N_13226,N_13179,N_13155);
xor U13227 (N_13227,N_13143,N_13112);
nand U13228 (N_13228,N_13065,N_13018);
and U13229 (N_13229,N_13199,N_13014);
and U13230 (N_13230,N_13067,N_13195);
and U13231 (N_13231,N_13006,N_13083);
xor U13232 (N_13232,N_13000,N_13171);
or U13233 (N_13233,N_13154,N_13026);
or U13234 (N_13234,N_13173,N_13059);
nand U13235 (N_13235,N_13082,N_13008);
or U13236 (N_13236,N_13139,N_13042);
and U13237 (N_13237,N_13032,N_13055);
xnor U13238 (N_13238,N_13197,N_13184);
nor U13239 (N_13239,N_13105,N_13190);
nor U13240 (N_13240,N_13165,N_13194);
and U13241 (N_13241,N_13122,N_13124);
nand U13242 (N_13242,N_13099,N_13078);
or U13243 (N_13243,N_13164,N_13060);
xor U13244 (N_13244,N_13080,N_13019);
nor U13245 (N_13245,N_13145,N_13017);
nand U13246 (N_13246,N_13003,N_13188);
and U13247 (N_13247,N_13177,N_13104);
and U13248 (N_13248,N_13077,N_13035);
and U13249 (N_13249,N_13157,N_13118);
nor U13250 (N_13250,N_13183,N_13149);
xor U13251 (N_13251,N_13140,N_13119);
or U13252 (N_13252,N_13013,N_13114);
or U13253 (N_13253,N_13063,N_13117);
or U13254 (N_13254,N_13069,N_13016);
xnor U13255 (N_13255,N_13088,N_13053);
or U13256 (N_13256,N_13162,N_13121);
and U13257 (N_13257,N_13185,N_13075);
nor U13258 (N_13258,N_13048,N_13176);
and U13259 (N_13259,N_13027,N_13084);
nor U13260 (N_13260,N_13113,N_13129);
nor U13261 (N_13261,N_13127,N_13096);
nor U13262 (N_13262,N_13066,N_13168);
and U13263 (N_13263,N_13180,N_13031);
or U13264 (N_13264,N_13150,N_13090);
or U13265 (N_13265,N_13046,N_13036);
xnor U13266 (N_13266,N_13020,N_13047);
xnor U13267 (N_13267,N_13133,N_13009);
or U13268 (N_13268,N_13012,N_13142);
and U13269 (N_13269,N_13182,N_13152);
nor U13270 (N_13270,N_13004,N_13101);
nor U13271 (N_13271,N_13081,N_13191);
and U13272 (N_13272,N_13057,N_13193);
and U13273 (N_13273,N_13072,N_13025);
and U13274 (N_13274,N_13174,N_13123);
xnor U13275 (N_13275,N_13022,N_13054);
xnor U13276 (N_13276,N_13163,N_13098);
or U13277 (N_13277,N_13137,N_13030);
and U13278 (N_13278,N_13062,N_13160);
xnor U13279 (N_13279,N_13011,N_13050);
nand U13280 (N_13280,N_13146,N_13058);
and U13281 (N_13281,N_13049,N_13181);
xor U13282 (N_13282,N_13044,N_13100);
xnor U13283 (N_13283,N_13002,N_13094);
xnor U13284 (N_13284,N_13144,N_13192);
xor U13285 (N_13285,N_13156,N_13061);
nor U13286 (N_13286,N_13167,N_13064);
and U13287 (N_13287,N_13034,N_13033);
nand U13288 (N_13288,N_13087,N_13135);
and U13289 (N_13289,N_13147,N_13056);
nor U13290 (N_13290,N_13134,N_13007);
xor U13291 (N_13291,N_13092,N_13024);
xor U13292 (N_13292,N_13095,N_13070);
or U13293 (N_13293,N_13010,N_13043);
nand U13294 (N_13294,N_13102,N_13045);
nand U13295 (N_13295,N_13068,N_13120);
and U13296 (N_13296,N_13151,N_13175);
or U13297 (N_13297,N_13074,N_13186);
nand U13298 (N_13298,N_13159,N_13126);
and U13299 (N_13299,N_13136,N_13158);
xnor U13300 (N_13300,N_13143,N_13043);
nor U13301 (N_13301,N_13052,N_13127);
or U13302 (N_13302,N_13062,N_13029);
xor U13303 (N_13303,N_13019,N_13172);
xnor U13304 (N_13304,N_13096,N_13114);
or U13305 (N_13305,N_13176,N_13120);
nand U13306 (N_13306,N_13112,N_13028);
nor U13307 (N_13307,N_13064,N_13005);
xnor U13308 (N_13308,N_13063,N_13135);
nand U13309 (N_13309,N_13031,N_13052);
xnor U13310 (N_13310,N_13135,N_13111);
xor U13311 (N_13311,N_13167,N_13090);
or U13312 (N_13312,N_13164,N_13175);
nor U13313 (N_13313,N_13118,N_13189);
nor U13314 (N_13314,N_13090,N_13046);
and U13315 (N_13315,N_13194,N_13140);
nor U13316 (N_13316,N_13044,N_13180);
nor U13317 (N_13317,N_13109,N_13081);
or U13318 (N_13318,N_13132,N_13033);
and U13319 (N_13319,N_13069,N_13189);
nor U13320 (N_13320,N_13129,N_13116);
or U13321 (N_13321,N_13123,N_13049);
xnor U13322 (N_13322,N_13091,N_13150);
or U13323 (N_13323,N_13068,N_13011);
nor U13324 (N_13324,N_13111,N_13189);
and U13325 (N_13325,N_13086,N_13069);
xor U13326 (N_13326,N_13094,N_13122);
nor U13327 (N_13327,N_13050,N_13167);
nor U13328 (N_13328,N_13133,N_13170);
or U13329 (N_13329,N_13118,N_13169);
xor U13330 (N_13330,N_13070,N_13140);
nor U13331 (N_13331,N_13064,N_13062);
nor U13332 (N_13332,N_13008,N_13123);
and U13333 (N_13333,N_13118,N_13063);
or U13334 (N_13334,N_13118,N_13192);
or U13335 (N_13335,N_13087,N_13131);
or U13336 (N_13336,N_13172,N_13015);
xor U13337 (N_13337,N_13093,N_13072);
xnor U13338 (N_13338,N_13133,N_13136);
or U13339 (N_13339,N_13073,N_13043);
nand U13340 (N_13340,N_13101,N_13162);
nand U13341 (N_13341,N_13176,N_13174);
or U13342 (N_13342,N_13193,N_13082);
xor U13343 (N_13343,N_13046,N_13173);
nand U13344 (N_13344,N_13043,N_13078);
or U13345 (N_13345,N_13035,N_13012);
nand U13346 (N_13346,N_13015,N_13001);
nor U13347 (N_13347,N_13126,N_13132);
xnor U13348 (N_13348,N_13080,N_13137);
nor U13349 (N_13349,N_13158,N_13071);
nand U13350 (N_13350,N_13067,N_13116);
and U13351 (N_13351,N_13193,N_13187);
xor U13352 (N_13352,N_13052,N_13143);
or U13353 (N_13353,N_13055,N_13139);
nor U13354 (N_13354,N_13123,N_13036);
and U13355 (N_13355,N_13048,N_13115);
and U13356 (N_13356,N_13165,N_13074);
xnor U13357 (N_13357,N_13045,N_13087);
or U13358 (N_13358,N_13042,N_13183);
nor U13359 (N_13359,N_13072,N_13089);
or U13360 (N_13360,N_13012,N_13134);
and U13361 (N_13361,N_13091,N_13149);
nand U13362 (N_13362,N_13181,N_13157);
nand U13363 (N_13363,N_13016,N_13058);
and U13364 (N_13364,N_13190,N_13059);
xnor U13365 (N_13365,N_13148,N_13188);
nand U13366 (N_13366,N_13137,N_13189);
xnor U13367 (N_13367,N_13106,N_13124);
and U13368 (N_13368,N_13001,N_13088);
xnor U13369 (N_13369,N_13071,N_13061);
xor U13370 (N_13370,N_13141,N_13158);
nor U13371 (N_13371,N_13096,N_13046);
xnor U13372 (N_13372,N_13103,N_13081);
nor U13373 (N_13373,N_13098,N_13077);
xnor U13374 (N_13374,N_13133,N_13068);
or U13375 (N_13375,N_13134,N_13154);
and U13376 (N_13376,N_13169,N_13187);
nand U13377 (N_13377,N_13088,N_13115);
xnor U13378 (N_13378,N_13019,N_13126);
or U13379 (N_13379,N_13111,N_13151);
xor U13380 (N_13380,N_13189,N_13168);
nand U13381 (N_13381,N_13062,N_13169);
nor U13382 (N_13382,N_13185,N_13035);
xnor U13383 (N_13383,N_13147,N_13163);
or U13384 (N_13384,N_13090,N_13008);
and U13385 (N_13385,N_13197,N_13140);
nand U13386 (N_13386,N_13064,N_13031);
nor U13387 (N_13387,N_13096,N_13188);
nand U13388 (N_13388,N_13091,N_13005);
and U13389 (N_13389,N_13112,N_13119);
and U13390 (N_13390,N_13128,N_13165);
and U13391 (N_13391,N_13088,N_13010);
nor U13392 (N_13392,N_13193,N_13066);
xnor U13393 (N_13393,N_13006,N_13169);
and U13394 (N_13394,N_13101,N_13092);
or U13395 (N_13395,N_13170,N_13167);
or U13396 (N_13396,N_13163,N_13086);
nor U13397 (N_13397,N_13152,N_13130);
nand U13398 (N_13398,N_13025,N_13099);
nand U13399 (N_13399,N_13158,N_13163);
or U13400 (N_13400,N_13216,N_13311);
nand U13401 (N_13401,N_13234,N_13301);
or U13402 (N_13402,N_13351,N_13207);
or U13403 (N_13403,N_13223,N_13215);
and U13404 (N_13404,N_13332,N_13343);
nor U13405 (N_13405,N_13239,N_13208);
nand U13406 (N_13406,N_13380,N_13305);
nor U13407 (N_13407,N_13302,N_13206);
or U13408 (N_13408,N_13290,N_13367);
xor U13409 (N_13409,N_13204,N_13396);
nand U13410 (N_13410,N_13210,N_13378);
nand U13411 (N_13411,N_13266,N_13219);
and U13412 (N_13412,N_13300,N_13362);
nand U13413 (N_13413,N_13379,N_13303);
nand U13414 (N_13414,N_13359,N_13316);
and U13415 (N_13415,N_13338,N_13254);
and U13416 (N_13416,N_13317,N_13320);
nor U13417 (N_13417,N_13275,N_13237);
or U13418 (N_13418,N_13389,N_13296);
nor U13419 (N_13419,N_13306,N_13361);
nor U13420 (N_13420,N_13383,N_13323);
nand U13421 (N_13421,N_13333,N_13256);
nand U13422 (N_13422,N_13279,N_13214);
nand U13423 (N_13423,N_13213,N_13288);
and U13424 (N_13424,N_13315,N_13203);
and U13425 (N_13425,N_13201,N_13335);
or U13426 (N_13426,N_13329,N_13269);
and U13427 (N_13427,N_13337,N_13393);
nand U13428 (N_13428,N_13372,N_13248);
nor U13429 (N_13429,N_13265,N_13340);
nand U13430 (N_13430,N_13261,N_13344);
or U13431 (N_13431,N_13264,N_13373);
xnor U13432 (N_13432,N_13330,N_13233);
or U13433 (N_13433,N_13224,N_13345);
and U13434 (N_13434,N_13384,N_13246);
nand U13435 (N_13435,N_13394,N_13352);
or U13436 (N_13436,N_13310,N_13211);
xnor U13437 (N_13437,N_13291,N_13358);
or U13438 (N_13438,N_13342,N_13238);
nand U13439 (N_13439,N_13293,N_13326);
xor U13440 (N_13440,N_13247,N_13241);
xor U13441 (N_13441,N_13220,N_13309);
and U13442 (N_13442,N_13390,N_13334);
nand U13443 (N_13443,N_13307,N_13205);
xnor U13444 (N_13444,N_13331,N_13245);
or U13445 (N_13445,N_13325,N_13282);
nand U13446 (N_13446,N_13386,N_13212);
xnor U13447 (N_13447,N_13382,N_13381);
or U13448 (N_13448,N_13298,N_13267);
nor U13449 (N_13449,N_13395,N_13263);
and U13450 (N_13450,N_13328,N_13365);
nor U13451 (N_13451,N_13257,N_13366);
xor U13452 (N_13452,N_13369,N_13304);
nand U13453 (N_13453,N_13376,N_13284);
xnor U13454 (N_13454,N_13251,N_13385);
or U13455 (N_13455,N_13285,N_13295);
xnor U13456 (N_13456,N_13363,N_13324);
nor U13457 (N_13457,N_13218,N_13322);
or U13458 (N_13458,N_13312,N_13370);
nand U13459 (N_13459,N_13286,N_13348);
xnor U13460 (N_13460,N_13364,N_13314);
xnor U13461 (N_13461,N_13287,N_13276);
nand U13462 (N_13462,N_13240,N_13388);
nand U13463 (N_13463,N_13355,N_13268);
or U13464 (N_13464,N_13375,N_13244);
xnor U13465 (N_13465,N_13374,N_13230);
or U13466 (N_13466,N_13226,N_13258);
and U13467 (N_13467,N_13371,N_13368);
nand U13468 (N_13468,N_13354,N_13341);
nor U13469 (N_13469,N_13231,N_13283);
xnor U13470 (N_13470,N_13274,N_13217);
or U13471 (N_13471,N_13399,N_13387);
nor U13472 (N_13472,N_13277,N_13350);
nor U13473 (N_13473,N_13232,N_13236);
nand U13474 (N_13474,N_13225,N_13260);
or U13475 (N_13475,N_13278,N_13255);
nand U13476 (N_13476,N_13259,N_13271);
xnor U13477 (N_13477,N_13228,N_13377);
xor U13478 (N_13478,N_13202,N_13292);
and U13479 (N_13479,N_13281,N_13346);
and U13480 (N_13480,N_13313,N_13347);
or U13481 (N_13481,N_13321,N_13280);
or U13482 (N_13482,N_13392,N_13270);
xor U13483 (N_13483,N_13398,N_13327);
or U13484 (N_13484,N_13222,N_13391);
or U13485 (N_13485,N_13397,N_13357);
or U13486 (N_13486,N_13242,N_13297);
nand U13487 (N_13487,N_13308,N_13360);
xor U13488 (N_13488,N_13252,N_13349);
nand U13489 (N_13489,N_13262,N_13319);
and U13490 (N_13490,N_13221,N_13273);
nand U13491 (N_13491,N_13227,N_13249);
xor U13492 (N_13492,N_13235,N_13356);
nand U13493 (N_13493,N_13353,N_13253);
and U13494 (N_13494,N_13272,N_13229);
xor U13495 (N_13495,N_13200,N_13339);
and U13496 (N_13496,N_13336,N_13318);
and U13497 (N_13497,N_13243,N_13294);
nor U13498 (N_13498,N_13299,N_13289);
nand U13499 (N_13499,N_13250,N_13209);
nor U13500 (N_13500,N_13349,N_13360);
xor U13501 (N_13501,N_13343,N_13338);
xnor U13502 (N_13502,N_13397,N_13242);
nand U13503 (N_13503,N_13362,N_13200);
nor U13504 (N_13504,N_13301,N_13368);
and U13505 (N_13505,N_13393,N_13308);
xor U13506 (N_13506,N_13360,N_13336);
or U13507 (N_13507,N_13203,N_13350);
xor U13508 (N_13508,N_13210,N_13289);
nor U13509 (N_13509,N_13374,N_13300);
or U13510 (N_13510,N_13348,N_13208);
and U13511 (N_13511,N_13290,N_13271);
or U13512 (N_13512,N_13346,N_13340);
and U13513 (N_13513,N_13296,N_13223);
nand U13514 (N_13514,N_13373,N_13275);
nor U13515 (N_13515,N_13247,N_13248);
xor U13516 (N_13516,N_13339,N_13290);
xor U13517 (N_13517,N_13321,N_13317);
nand U13518 (N_13518,N_13353,N_13277);
nand U13519 (N_13519,N_13368,N_13264);
nor U13520 (N_13520,N_13295,N_13363);
or U13521 (N_13521,N_13202,N_13286);
and U13522 (N_13522,N_13335,N_13363);
and U13523 (N_13523,N_13394,N_13323);
nor U13524 (N_13524,N_13317,N_13297);
or U13525 (N_13525,N_13388,N_13268);
and U13526 (N_13526,N_13231,N_13280);
xor U13527 (N_13527,N_13317,N_13398);
nor U13528 (N_13528,N_13347,N_13352);
and U13529 (N_13529,N_13205,N_13319);
xor U13530 (N_13530,N_13301,N_13278);
and U13531 (N_13531,N_13289,N_13282);
or U13532 (N_13532,N_13368,N_13321);
nor U13533 (N_13533,N_13319,N_13307);
xnor U13534 (N_13534,N_13364,N_13250);
or U13535 (N_13535,N_13342,N_13345);
or U13536 (N_13536,N_13390,N_13294);
and U13537 (N_13537,N_13278,N_13215);
nor U13538 (N_13538,N_13211,N_13390);
or U13539 (N_13539,N_13352,N_13270);
or U13540 (N_13540,N_13313,N_13320);
or U13541 (N_13541,N_13395,N_13363);
nand U13542 (N_13542,N_13392,N_13296);
and U13543 (N_13543,N_13202,N_13265);
or U13544 (N_13544,N_13200,N_13226);
xor U13545 (N_13545,N_13340,N_13399);
and U13546 (N_13546,N_13288,N_13218);
and U13547 (N_13547,N_13291,N_13301);
or U13548 (N_13548,N_13202,N_13285);
nand U13549 (N_13549,N_13249,N_13246);
nor U13550 (N_13550,N_13272,N_13342);
nor U13551 (N_13551,N_13221,N_13272);
nor U13552 (N_13552,N_13213,N_13381);
and U13553 (N_13553,N_13351,N_13374);
or U13554 (N_13554,N_13216,N_13246);
and U13555 (N_13555,N_13341,N_13256);
or U13556 (N_13556,N_13237,N_13305);
xnor U13557 (N_13557,N_13314,N_13233);
or U13558 (N_13558,N_13277,N_13300);
and U13559 (N_13559,N_13214,N_13350);
nor U13560 (N_13560,N_13276,N_13214);
nand U13561 (N_13561,N_13289,N_13304);
nor U13562 (N_13562,N_13248,N_13349);
and U13563 (N_13563,N_13263,N_13281);
nor U13564 (N_13564,N_13393,N_13286);
and U13565 (N_13565,N_13278,N_13307);
xnor U13566 (N_13566,N_13271,N_13307);
or U13567 (N_13567,N_13216,N_13232);
and U13568 (N_13568,N_13321,N_13255);
and U13569 (N_13569,N_13295,N_13273);
xnor U13570 (N_13570,N_13318,N_13213);
xnor U13571 (N_13571,N_13241,N_13307);
nand U13572 (N_13572,N_13247,N_13272);
nand U13573 (N_13573,N_13240,N_13276);
or U13574 (N_13574,N_13359,N_13377);
or U13575 (N_13575,N_13335,N_13372);
nand U13576 (N_13576,N_13267,N_13302);
nand U13577 (N_13577,N_13231,N_13309);
xnor U13578 (N_13578,N_13239,N_13288);
nor U13579 (N_13579,N_13349,N_13251);
and U13580 (N_13580,N_13263,N_13372);
and U13581 (N_13581,N_13316,N_13375);
nand U13582 (N_13582,N_13358,N_13286);
nand U13583 (N_13583,N_13305,N_13257);
nand U13584 (N_13584,N_13269,N_13233);
nor U13585 (N_13585,N_13276,N_13345);
and U13586 (N_13586,N_13211,N_13345);
or U13587 (N_13587,N_13386,N_13246);
xnor U13588 (N_13588,N_13393,N_13277);
and U13589 (N_13589,N_13258,N_13212);
and U13590 (N_13590,N_13396,N_13319);
nand U13591 (N_13591,N_13226,N_13399);
xor U13592 (N_13592,N_13352,N_13237);
xor U13593 (N_13593,N_13253,N_13315);
nand U13594 (N_13594,N_13329,N_13201);
nor U13595 (N_13595,N_13323,N_13274);
nand U13596 (N_13596,N_13224,N_13236);
nand U13597 (N_13597,N_13315,N_13351);
nor U13598 (N_13598,N_13237,N_13262);
xor U13599 (N_13599,N_13206,N_13332);
nor U13600 (N_13600,N_13531,N_13542);
and U13601 (N_13601,N_13515,N_13514);
nor U13602 (N_13602,N_13401,N_13464);
nor U13603 (N_13603,N_13403,N_13416);
and U13604 (N_13604,N_13442,N_13410);
xor U13605 (N_13605,N_13582,N_13441);
nand U13606 (N_13606,N_13587,N_13507);
or U13607 (N_13607,N_13517,N_13585);
nand U13608 (N_13608,N_13497,N_13419);
nor U13609 (N_13609,N_13492,N_13570);
and U13610 (N_13610,N_13539,N_13415);
nand U13611 (N_13611,N_13460,N_13448);
nand U13612 (N_13612,N_13576,N_13523);
nor U13613 (N_13613,N_13411,N_13427);
nand U13614 (N_13614,N_13499,N_13599);
xnor U13615 (N_13615,N_13463,N_13553);
nand U13616 (N_13616,N_13589,N_13597);
nand U13617 (N_13617,N_13583,N_13491);
or U13618 (N_13618,N_13483,N_13516);
nand U13619 (N_13619,N_13575,N_13557);
or U13620 (N_13620,N_13472,N_13417);
and U13621 (N_13621,N_13511,N_13462);
nand U13622 (N_13622,N_13406,N_13530);
nor U13623 (N_13623,N_13565,N_13588);
nor U13624 (N_13624,N_13494,N_13535);
xnor U13625 (N_13625,N_13524,N_13509);
or U13626 (N_13626,N_13452,N_13493);
nor U13627 (N_13627,N_13573,N_13598);
xnor U13628 (N_13628,N_13446,N_13421);
nand U13629 (N_13629,N_13490,N_13581);
nor U13630 (N_13630,N_13420,N_13590);
xnor U13631 (N_13631,N_13536,N_13593);
or U13632 (N_13632,N_13434,N_13487);
or U13633 (N_13633,N_13432,N_13486);
nor U13634 (N_13634,N_13512,N_13540);
nand U13635 (N_13635,N_13484,N_13546);
nor U13636 (N_13636,N_13586,N_13549);
nor U13637 (N_13637,N_13554,N_13456);
xnor U13638 (N_13638,N_13471,N_13505);
nand U13639 (N_13639,N_13558,N_13412);
xnor U13640 (N_13640,N_13532,N_13481);
and U13641 (N_13641,N_13564,N_13454);
or U13642 (N_13642,N_13596,N_13444);
nor U13643 (N_13643,N_13469,N_13467);
nor U13644 (N_13644,N_13485,N_13508);
xor U13645 (N_13645,N_13578,N_13574);
or U13646 (N_13646,N_13474,N_13522);
xnor U13647 (N_13647,N_13468,N_13520);
or U13648 (N_13648,N_13513,N_13488);
nand U13649 (N_13649,N_13451,N_13525);
nand U13650 (N_13650,N_13592,N_13449);
or U13651 (N_13651,N_13569,N_13436);
xnor U13652 (N_13652,N_13433,N_13521);
and U13653 (N_13653,N_13430,N_13437);
and U13654 (N_13654,N_13550,N_13591);
or U13655 (N_13655,N_13547,N_13537);
xnor U13656 (N_13656,N_13404,N_13453);
or U13657 (N_13657,N_13527,N_13482);
or U13658 (N_13658,N_13450,N_13435);
xor U13659 (N_13659,N_13478,N_13510);
nor U13660 (N_13660,N_13526,N_13429);
nand U13661 (N_13661,N_13476,N_13504);
nor U13662 (N_13662,N_13461,N_13551);
and U13663 (N_13663,N_13584,N_13562);
or U13664 (N_13664,N_13480,N_13423);
nand U13665 (N_13665,N_13457,N_13545);
nand U13666 (N_13666,N_13555,N_13519);
nand U13667 (N_13667,N_13479,N_13402);
or U13668 (N_13668,N_13466,N_13568);
xnor U13669 (N_13669,N_13455,N_13572);
nor U13670 (N_13670,N_13529,N_13566);
nor U13671 (N_13671,N_13475,N_13563);
and U13672 (N_13672,N_13459,N_13595);
nor U13673 (N_13673,N_13424,N_13445);
or U13674 (N_13674,N_13458,N_13556);
nand U13675 (N_13675,N_13561,N_13405);
and U13676 (N_13676,N_13470,N_13489);
nor U13677 (N_13677,N_13571,N_13534);
and U13678 (N_13678,N_13500,N_13501);
nor U13679 (N_13679,N_13477,N_13408);
nand U13680 (N_13680,N_13594,N_13506);
nand U13681 (N_13681,N_13422,N_13496);
or U13682 (N_13682,N_13438,N_13447);
xnor U13683 (N_13683,N_13538,N_13425);
nand U13684 (N_13684,N_13407,N_13552);
nand U13685 (N_13685,N_13413,N_13465);
or U13686 (N_13686,N_13414,N_13560);
nor U13687 (N_13687,N_13503,N_13528);
and U13688 (N_13688,N_13567,N_13577);
xor U13689 (N_13689,N_13559,N_13518);
nand U13690 (N_13690,N_13443,N_13426);
nand U13691 (N_13691,N_13431,N_13400);
and U13692 (N_13692,N_13439,N_13418);
nand U13693 (N_13693,N_13580,N_13428);
nand U13694 (N_13694,N_13543,N_13498);
nand U13695 (N_13695,N_13544,N_13548);
nor U13696 (N_13696,N_13502,N_13579);
xor U13697 (N_13697,N_13473,N_13409);
nand U13698 (N_13698,N_13440,N_13541);
and U13699 (N_13699,N_13533,N_13495);
or U13700 (N_13700,N_13418,N_13597);
nand U13701 (N_13701,N_13513,N_13570);
or U13702 (N_13702,N_13500,N_13595);
or U13703 (N_13703,N_13533,N_13497);
nand U13704 (N_13704,N_13560,N_13525);
xor U13705 (N_13705,N_13568,N_13528);
nand U13706 (N_13706,N_13472,N_13532);
nor U13707 (N_13707,N_13429,N_13430);
nand U13708 (N_13708,N_13444,N_13445);
nor U13709 (N_13709,N_13549,N_13437);
xnor U13710 (N_13710,N_13555,N_13593);
nand U13711 (N_13711,N_13513,N_13492);
xnor U13712 (N_13712,N_13555,N_13508);
nand U13713 (N_13713,N_13431,N_13537);
nor U13714 (N_13714,N_13446,N_13479);
nand U13715 (N_13715,N_13446,N_13524);
nand U13716 (N_13716,N_13451,N_13401);
and U13717 (N_13717,N_13535,N_13558);
and U13718 (N_13718,N_13518,N_13486);
or U13719 (N_13719,N_13518,N_13426);
and U13720 (N_13720,N_13551,N_13450);
xor U13721 (N_13721,N_13420,N_13511);
and U13722 (N_13722,N_13512,N_13553);
and U13723 (N_13723,N_13500,N_13476);
nor U13724 (N_13724,N_13494,N_13466);
nand U13725 (N_13725,N_13507,N_13521);
xor U13726 (N_13726,N_13409,N_13480);
and U13727 (N_13727,N_13578,N_13589);
nand U13728 (N_13728,N_13444,N_13524);
xnor U13729 (N_13729,N_13425,N_13524);
and U13730 (N_13730,N_13568,N_13414);
xor U13731 (N_13731,N_13512,N_13500);
or U13732 (N_13732,N_13430,N_13439);
and U13733 (N_13733,N_13470,N_13498);
and U13734 (N_13734,N_13460,N_13583);
and U13735 (N_13735,N_13562,N_13400);
and U13736 (N_13736,N_13586,N_13591);
and U13737 (N_13737,N_13427,N_13581);
or U13738 (N_13738,N_13429,N_13473);
nand U13739 (N_13739,N_13453,N_13507);
and U13740 (N_13740,N_13464,N_13518);
and U13741 (N_13741,N_13476,N_13409);
nand U13742 (N_13742,N_13518,N_13568);
and U13743 (N_13743,N_13540,N_13554);
nor U13744 (N_13744,N_13541,N_13445);
and U13745 (N_13745,N_13551,N_13516);
and U13746 (N_13746,N_13443,N_13438);
or U13747 (N_13747,N_13445,N_13590);
xor U13748 (N_13748,N_13556,N_13535);
or U13749 (N_13749,N_13585,N_13456);
nand U13750 (N_13750,N_13511,N_13521);
nand U13751 (N_13751,N_13557,N_13479);
or U13752 (N_13752,N_13484,N_13457);
or U13753 (N_13753,N_13410,N_13412);
xnor U13754 (N_13754,N_13589,N_13421);
and U13755 (N_13755,N_13481,N_13514);
and U13756 (N_13756,N_13494,N_13455);
xor U13757 (N_13757,N_13475,N_13549);
nand U13758 (N_13758,N_13431,N_13518);
and U13759 (N_13759,N_13480,N_13473);
nand U13760 (N_13760,N_13565,N_13417);
nand U13761 (N_13761,N_13452,N_13489);
xnor U13762 (N_13762,N_13462,N_13574);
nor U13763 (N_13763,N_13466,N_13598);
and U13764 (N_13764,N_13500,N_13480);
nand U13765 (N_13765,N_13563,N_13419);
nand U13766 (N_13766,N_13482,N_13480);
or U13767 (N_13767,N_13544,N_13439);
or U13768 (N_13768,N_13427,N_13530);
xor U13769 (N_13769,N_13568,N_13500);
nor U13770 (N_13770,N_13510,N_13548);
or U13771 (N_13771,N_13451,N_13418);
nor U13772 (N_13772,N_13428,N_13442);
nand U13773 (N_13773,N_13583,N_13526);
and U13774 (N_13774,N_13448,N_13491);
and U13775 (N_13775,N_13418,N_13488);
and U13776 (N_13776,N_13478,N_13430);
or U13777 (N_13777,N_13551,N_13569);
or U13778 (N_13778,N_13554,N_13443);
or U13779 (N_13779,N_13539,N_13561);
xor U13780 (N_13780,N_13571,N_13478);
nand U13781 (N_13781,N_13436,N_13521);
and U13782 (N_13782,N_13550,N_13567);
xor U13783 (N_13783,N_13460,N_13490);
xnor U13784 (N_13784,N_13474,N_13491);
nor U13785 (N_13785,N_13441,N_13499);
and U13786 (N_13786,N_13433,N_13546);
nor U13787 (N_13787,N_13444,N_13438);
nor U13788 (N_13788,N_13569,N_13555);
and U13789 (N_13789,N_13452,N_13588);
or U13790 (N_13790,N_13476,N_13407);
nand U13791 (N_13791,N_13575,N_13553);
xnor U13792 (N_13792,N_13463,N_13406);
nor U13793 (N_13793,N_13405,N_13487);
xor U13794 (N_13794,N_13489,N_13444);
xnor U13795 (N_13795,N_13470,N_13544);
or U13796 (N_13796,N_13519,N_13401);
xor U13797 (N_13797,N_13576,N_13556);
or U13798 (N_13798,N_13407,N_13502);
xnor U13799 (N_13799,N_13472,N_13593);
and U13800 (N_13800,N_13703,N_13790);
nor U13801 (N_13801,N_13695,N_13651);
and U13802 (N_13802,N_13764,N_13637);
xnor U13803 (N_13803,N_13794,N_13609);
nand U13804 (N_13804,N_13795,N_13740);
nand U13805 (N_13805,N_13675,N_13636);
nor U13806 (N_13806,N_13697,N_13706);
or U13807 (N_13807,N_13661,N_13618);
and U13808 (N_13808,N_13632,N_13656);
or U13809 (N_13809,N_13640,N_13648);
or U13810 (N_13810,N_13620,N_13777);
and U13811 (N_13811,N_13773,N_13670);
or U13812 (N_13812,N_13678,N_13603);
and U13813 (N_13813,N_13626,N_13638);
nor U13814 (N_13814,N_13754,N_13733);
or U13815 (N_13815,N_13724,N_13787);
nand U13816 (N_13816,N_13685,N_13792);
or U13817 (N_13817,N_13753,N_13728);
nand U13818 (N_13818,N_13729,N_13709);
and U13819 (N_13819,N_13743,N_13713);
nand U13820 (N_13820,N_13652,N_13750);
xor U13821 (N_13821,N_13704,N_13759);
or U13822 (N_13822,N_13708,N_13681);
or U13823 (N_13823,N_13757,N_13747);
nor U13824 (N_13824,N_13601,N_13745);
nand U13825 (N_13825,N_13606,N_13705);
and U13826 (N_13826,N_13614,N_13723);
nand U13827 (N_13827,N_13727,N_13692);
nor U13828 (N_13828,N_13650,N_13720);
nand U13829 (N_13829,N_13749,N_13798);
nor U13830 (N_13830,N_13744,N_13639);
nor U13831 (N_13831,N_13671,N_13687);
nand U13832 (N_13832,N_13732,N_13746);
nand U13833 (N_13833,N_13761,N_13756);
nor U13834 (N_13834,N_13734,N_13748);
xnor U13835 (N_13835,N_13717,N_13633);
nor U13836 (N_13836,N_13645,N_13643);
nor U13837 (N_13837,N_13742,N_13629);
nor U13838 (N_13838,N_13625,N_13783);
nand U13839 (N_13839,N_13760,N_13621);
or U13840 (N_13840,N_13763,N_13765);
nor U13841 (N_13841,N_13722,N_13668);
nor U13842 (N_13842,N_13775,N_13657);
or U13843 (N_13843,N_13774,N_13715);
and U13844 (N_13844,N_13776,N_13780);
xor U13845 (N_13845,N_13644,N_13769);
nor U13846 (N_13846,N_13721,N_13786);
xnor U13847 (N_13847,N_13781,N_13793);
or U13848 (N_13848,N_13688,N_13613);
nand U13849 (N_13849,N_13731,N_13762);
and U13850 (N_13850,N_13738,N_13653);
nand U13851 (N_13851,N_13667,N_13770);
xnor U13852 (N_13852,N_13736,N_13767);
nand U13853 (N_13853,N_13752,N_13666);
nor U13854 (N_13854,N_13689,N_13683);
or U13855 (N_13855,N_13610,N_13772);
and U13856 (N_13856,N_13710,N_13607);
nand U13857 (N_13857,N_13696,N_13663);
or U13858 (N_13858,N_13628,N_13701);
xor U13859 (N_13859,N_13766,N_13642);
and U13860 (N_13860,N_13686,N_13741);
and U13861 (N_13861,N_13615,N_13699);
xor U13862 (N_13862,N_13647,N_13739);
or U13863 (N_13863,N_13711,N_13634);
and U13864 (N_13864,N_13684,N_13617);
xnor U13865 (N_13865,N_13600,N_13797);
xnor U13866 (N_13866,N_13694,N_13700);
and U13867 (N_13867,N_13604,N_13782);
nand U13868 (N_13868,N_13630,N_13735);
and U13869 (N_13869,N_13771,N_13680);
or U13870 (N_13870,N_13612,N_13737);
and U13871 (N_13871,N_13646,N_13758);
nand U13872 (N_13872,N_13785,N_13677);
or U13873 (N_13873,N_13608,N_13673);
and U13874 (N_13874,N_13658,N_13791);
or U13875 (N_13875,N_13751,N_13691);
nand U13876 (N_13876,N_13796,N_13712);
nand U13877 (N_13877,N_13662,N_13789);
nor U13878 (N_13878,N_13693,N_13660);
or U13879 (N_13879,N_13602,N_13755);
nor U13880 (N_13880,N_13611,N_13635);
nor U13881 (N_13881,N_13627,N_13768);
and U13882 (N_13882,N_13665,N_13730);
nand U13883 (N_13883,N_13664,N_13659);
and U13884 (N_13884,N_13698,N_13779);
and U13885 (N_13885,N_13725,N_13719);
or U13886 (N_13886,N_13682,N_13669);
and U13887 (N_13887,N_13674,N_13623);
and U13888 (N_13888,N_13707,N_13655);
nor U13889 (N_13889,N_13624,N_13631);
or U13890 (N_13890,N_13616,N_13649);
nor U13891 (N_13891,N_13605,N_13622);
and U13892 (N_13892,N_13718,N_13690);
nor U13893 (N_13893,N_13788,N_13716);
nand U13894 (N_13894,N_13641,N_13679);
or U13895 (N_13895,N_13619,N_13784);
and U13896 (N_13896,N_13676,N_13654);
or U13897 (N_13897,N_13726,N_13714);
or U13898 (N_13898,N_13672,N_13799);
and U13899 (N_13899,N_13702,N_13778);
or U13900 (N_13900,N_13669,N_13713);
xor U13901 (N_13901,N_13700,N_13655);
xnor U13902 (N_13902,N_13628,N_13615);
nor U13903 (N_13903,N_13795,N_13704);
xor U13904 (N_13904,N_13776,N_13766);
xor U13905 (N_13905,N_13609,N_13780);
nand U13906 (N_13906,N_13686,N_13692);
xor U13907 (N_13907,N_13750,N_13775);
nand U13908 (N_13908,N_13628,N_13660);
and U13909 (N_13909,N_13653,N_13662);
and U13910 (N_13910,N_13692,N_13797);
xnor U13911 (N_13911,N_13635,N_13723);
nand U13912 (N_13912,N_13742,N_13716);
xor U13913 (N_13913,N_13792,N_13665);
nand U13914 (N_13914,N_13684,N_13692);
nand U13915 (N_13915,N_13787,N_13720);
nor U13916 (N_13916,N_13762,N_13681);
nand U13917 (N_13917,N_13792,N_13686);
nand U13918 (N_13918,N_13750,N_13624);
nor U13919 (N_13919,N_13697,N_13640);
xor U13920 (N_13920,N_13733,N_13729);
nand U13921 (N_13921,N_13669,N_13722);
and U13922 (N_13922,N_13618,N_13773);
or U13923 (N_13923,N_13614,N_13753);
nor U13924 (N_13924,N_13705,N_13711);
nor U13925 (N_13925,N_13767,N_13761);
nand U13926 (N_13926,N_13781,N_13691);
nor U13927 (N_13927,N_13655,N_13702);
nand U13928 (N_13928,N_13649,N_13652);
and U13929 (N_13929,N_13690,N_13716);
xor U13930 (N_13930,N_13756,N_13653);
or U13931 (N_13931,N_13690,N_13759);
or U13932 (N_13932,N_13711,N_13690);
and U13933 (N_13933,N_13730,N_13683);
nor U13934 (N_13934,N_13744,N_13611);
nor U13935 (N_13935,N_13635,N_13658);
and U13936 (N_13936,N_13794,N_13769);
or U13937 (N_13937,N_13663,N_13602);
xor U13938 (N_13938,N_13717,N_13793);
xnor U13939 (N_13939,N_13618,N_13735);
and U13940 (N_13940,N_13615,N_13669);
or U13941 (N_13941,N_13649,N_13780);
and U13942 (N_13942,N_13741,N_13651);
nor U13943 (N_13943,N_13715,N_13736);
nor U13944 (N_13944,N_13683,N_13781);
nor U13945 (N_13945,N_13732,N_13781);
and U13946 (N_13946,N_13749,N_13773);
and U13947 (N_13947,N_13676,N_13701);
nor U13948 (N_13948,N_13730,N_13612);
nor U13949 (N_13949,N_13656,N_13688);
nand U13950 (N_13950,N_13691,N_13735);
nor U13951 (N_13951,N_13690,N_13612);
nor U13952 (N_13952,N_13670,N_13629);
xnor U13953 (N_13953,N_13632,N_13717);
or U13954 (N_13954,N_13671,N_13781);
and U13955 (N_13955,N_13797,N_13687);
nor U13956 (N_13956,N_13643,N_13660);
xor U13957 (N_13957,N_13779,N_13701);
nand U13958 (N_13958,N_13706,N_13686);
nor U13959 (N_13959,N_13756,N_13798);
nor U13960 (N_13960,N_13695,N_13675);
nor U13961 (N_13961,N_13609,N_13734);
nor U13962 (N_13962,N_13615,N_13607);
xnor U13963 (N_13963,N_13646,N_13613);
and U13964 (N_13964,N_13729,N_13639);
xnor U13965 (N_13965,N_13718,N_13658);
and U13966 (N_13966,N_13714,N_13741);
or U13967 (N_13967,N_13752,N_13626);
nand U13968 (N_13968,N_13712,N_13738);
xor U13969 (N_13969,N_13683,N_13770);
or U13970 (N_13970,N_13609,N_13720);
nor U13971 (N_13971,N_13671,N_13759);
or U13972 (N_13972,N_13743,N_13763);
and U13973 (N_13973,N_13790,N_13601);
nor U13974 (N_13974,N_13791,N_13602);
nand U13975 (N_13975,N_13773,N_13710);
nor U13976 (N_13976,N_13737,N_13658);
or U13977 (N_13977,N_13674,N_13724);
nand U13978 (N_13978,N_13769,N_13721);
xor U13979 (N_13979,N_13633,N_13675);
nand U13980 (N_13980,N_13694,N_13723);
nor U13981 (N_13981,N_13620,N_13642);
and U13982 (N_13982,N_13749,N_13613);
nor U13983 (N_13983,N_13621,N_13704);
or U13984 (N_13984,N_13761,N_13793);
xnor U13985 (N_13985,N_13675,N_13672);
and U13986 (N_13986,N_13631,N_13619);
or U13987 (N_13987,N_13718,N_13623);
and U13988 (N_13988,N_13722,N_13704);
nand U13989 (N_13989,N_13766,N_13795);
or U13990 (N_13990,N_13765,N_13611);
nor U13991 (N_13991,N_13739,N_13714);
or U13992 (N_13992,N_13602,N_13758);
nor U13993 (N_13993,N_13633,N_13727);
nor U13994 (N_13994,N_13615,N_13612);
xnor U13995 (N_13995,N_13741,N_13613);
or U13996 (N_13996,N_13785,N_13762);
nor U13997 (N_13997,N_13621,N_13787);
xor U13998 (N_13998,N_13669,N_13665);
and U13999 (N_13999,N_13633,N_13629);
or U14000 (N_14000,N_13938,N_13907);
or U14001 (N_14001,N_13914,N_13803);
xor U14002 (N_14002,N_13875,N_13926);
and U14003 (N_14003,N_13877,N_13922);
or U14004 (N_14004,N_13954,N_13944);
nand U14005 (N_14005,N_13884,N_13928);
or U14006 (N_14006,N_13949,N_13859);
nor U14007 (N_14007,N_13996,N_13992);
xor U14008 (N_14008,N_13882,N_13902);
nor U14009 (N_14009,N_13873,N_13931);
or U14010 (N_14010,N_13961,N_13836);
xnor U14011 (N_14011,N_13981,N_13853);
nand U14012 (N_14012,N_13971,N_13878);
nor U14013 (N_14013,N_13821,N_13960);
and U14014 (N_14014,N_13917,N_13876);
nand U14015 (N_14015,N_13872,N_13924);
or U14016 (N_14016,N_13871,N_13935);
nor U14017 (N_14017,N_13955,N_13813);
xnor U14018 (N_14018,N_13833,N_13987);
or U14019 (N_14019,N_13899,N_13934);
xor U14020 (N_14020,N_13831,N_13844);
and U14021 (N_14021,N_13915,N_13863);
nand U14022 (N_14022,N_13905,N_13834);
nand U14023 (N_14023,N_13950,N_13898);
xor U14024 (N_14024,N_13812,N_13823);
nand U14025 (N_14025,N_13858,N_13886);
or U14026 (N_14026,N_13945,N_13866);
and U14027 (N_14027,N_13930,N_13837);
or U14028 (N_14028,N_13976,N_13849);
or U14029 (N_14029,N_13982,N_13895);
nand U14030 (N_14030,N_13865,N_13838);
and U14031 (N_14031,N_13929,N_13840);
xnor U14032 (N_14032,N_13921,N_13941);
or U14033 (N_14033,N_13850,N_13901);
xor U14034 (N_14034,N_13942,N_13986);
and U14035 (N_14035,N_13968,N_13818);
nor U14036 (N_14036,N_13868,N_13842);
and U14037 (N_14037,N_13879,N_13825);
xor U14038 (N_14038,N_13993,N_13851);
xnor U14039 (N_14039,N_13835,N_13841);
nor U14040 (N_14040,N_13810,N_13888);
and U14041 (N_14041,N_13947,N_13966);
xnor U14042 (N_14042,N_13965,N_13903);
or U14043 (N_14043,N_13811,N_13827);
and U14044 (N_14044,N_13932,N_13867);
nor U14045 (N_14045,N_13925,N_13998);
nand U14046 (N_14046,N_13860,N_13862);
xor U14047 (N_14047,N_13889,N_13874);
or U14048 (N_14048,N_13852,N_13896);
xor U14049 (N_14049,N_13906,N_13956);
or U14050 (N_14050,N_13824,N_13820);
nand U14051 (N_14051,N_13943,N_13819);
nor U14052 (N_14052,N_13978,N_13848);
xor U14053 (N_14053,N_13885,N_13995);
xnor U14054 (N_14054,N_13809,N_13937);
and U14055 (N_14055,N_13946,N_13883);
nand U14056 (N_14056,N_13897,N_13843);
nor U14057 (N_14057,N_13985,N_13999);
nor U14058 (N_14058,N_13890,N_13984);
nor U14059 (N_14059,N_13967,N_13940);
or U14060 (N_14060,N_13904,N_13958);
and U14061 (N_14061,N_13972,N_13856);
nand U14062 (N_14062,N_13894,N_13962);
and U14063 (N_14063,N_13948,N_13991);
nand U14064 (N_14064,N_13887,N_13912);
nor U14065 (N_14065,N_13814,N_13861);
nor U14066 (N_14066,N_13919,N_13893);
and U14067 (N_14067,N_13936,N_13970);
and U14068 (N_14068,N_13913,N_13845);
nor U14069 (N_14069,N_13951,N_13920);
nand U14070 (N_14070,N_13892,N_13846);
or U14071 (N_14071,N_13963,N_13805);
nand U14072 (N_14072,N_13854,N_13828);
and U14073 (N_14073,N_13979,N_13801);
nand U14074 (N_14074,N_13880,N_13909);
nor U14075 (N_14075,N_13826,N_13959);
and U14076 (N_14076,N_13857,N_13832);
or U14077 (N_14077,N_13933,N_13989);
and U14078 (N_14078,N_13808,N_13870);
nor U14079 (N_14079,N_13807,N_13900);
and U14080 (N_14080,N_13997,N_13911);
or U14081 (N_14081,N_13973,N_13800);
nand U14082 (N_14082,N_13939,N_13975);
or U14083 (N_14083,N_13977,N_13869);
nand U14084 (N_14084,N_13839,N_13829);
or U14085 (N_14085,N_13990,N_13855);
nand U14086 (N_14086,N_13817,N_13988);
and U14087 (N_14087,N_13891,N_13952);
and U14088 (N_14088,N_13881,N_13806);
nand U14089 (N_14089,N_13816,N_13918);
and U14090 (N_14090,N_13802,N_13980);
or U14091 (N_14091,N_13957,N_13815);
or U14092 (N_14092,N_13927,N_13974);
and U14093 (N_14093,N_13910,N_13830);
nand U14094 (N_14094,N_13983,N_13916);
nor U14095 (N_14095,N_13969,N_13822);
or U14096 (N_14096,N_13847,N_13864);
xnor U14097 (N_14097,N_13994,N_13923);
and U14098 (N_14098,N_13953,N_13908);
or U14099 (N_14099,N_13804,N_13964);
xnor U14100 (N_14100,N_13902,N_13800);
and U14101 (N_14101,N_13996,N_13865);
nor U14102 (N_14102,N_13814,N_13993);
and U14103 (N_14103,N_13910,N_13851);
or U14104 (N_14104,N_13911,N_13866);
nand U14105 (N_14105,N_13894,N_13849);
nor U14106 (N_14106,N_13847,N_13971);
xnor U14107 (N_14107,N_13960,N_13984);
xnor U14108 (N_14108,N_13882,N_13823);
nand U14109 (N_14109,N_13925,N_13900);
and U14110 (N_14110,N_13963,N_13959);
or U14111 (N_14111,N_13920,N_13949);
or U14112 (N_14112,N_13909,N_13990);
or U14113 (N_14113,N_13900,N_13838);
nor U14114 (N_14114,N_13968,N_13848);
or U14115 (N_14115,N_13812,N_13920);
nor U14116 (N_14116,N_13992,N_13824);
nor U14117 (N_14117,N_13808,N_13991);
and U14118 (N_14118,N_13944,N_13959);
nor U14119 (N_14119,N_13842,N_13879);
nor U14120 (N_14120,N_13848,N_13901);
or U14121 (N_14121,N_13850,N_13959);
nor U14122 (N_14122,N_13940,N_13932);
nor U14123 (N_14123,N_13831,N_13864);
and U14124 (N_14124,N_13978,N_13830);
xnor U14125 (N_14125,N_13812,N_13916);
and U14126 (N_14126,N_13838,N_13982);
xnor U14127 (N_14127,N_13952,N_13967);
nand U14128 (N_14128,N_13983,N_13850);
and U14129 (N_14129,N_13997,N_13929);
nand U14130 (N_14130,N_13954,N_13900);
nand U14131 (N_14131,N_13922,N_13993);
nand U14132 (N_14132,N_13855,N_13906);
xnor U14133 (N_14133,N_13850,N_13996);
or U14134 (N_14134,N_13872,N_13937);
nand U14135 (N_14135,N_13906,N_13848);
nand U14136 (N_14136,N_13898,N_13840);
and U14137 (N_14137,N_13949,N_13869);
nor U14138 (N_14138,N_13936,N_13861);
and U14139 (N_14139,N_13956,N_13819);
or U14140 (N_14140,N_13989,N_13813);
xor U14141 (N_14141,N_13936,N_13940);
and U14142 (N_14142,N_13872,N_13829);
xor U14143 (N_14143,N_13818,N_13993);
or U14144 (N_14144,N_13994,N_13958);
or U14145 (N_14145,N_13957,N_13816);
or U14146 (N_14146,N_13957,N_13804);
nand U14147 (N_14147,N_13970,N_13859);
nand U14148 (N_14148,N_13977,N_13834);
or U14149 (N_14149,N_13807,N_13995);
nand U14150 (N_14150,N_13892,N_13806);
and U14151 (N_14151,N_13828,N_13885);
xor U14152 (N_14152,N_13993,N_13881);
nor U14153 (N_14153,N_13937,N_13884);
or U14154 (N_14154,N_13906,N_13820);
xnor U14155 (N_14155,N_13944,N_13997);
and U14156 (N_14156,N_13806,N_13948);
and U14157 (N_14157,N_13928,N_13940);
and U14158 (N_14158,N_13908,N_13926);
nor U14159 (N_14159,N_13894,N_13986);
xnor U14160 (N_14160,N_13909,N_13895);
or U14161 (N_14161,N_13952,N_13849);
nor U14162 (N_14162,N_13898,N_13945);
or U14163 (N_14163,N_13994,N_13972);
nor U14164 (N_14164,N_13831,N_13896);
xor U14165 (N_14165,N_13872,N_13900);
xor U14166 (N_14166,N_13979,N_13983);
or U14167 (N_14167,N_13872,N_13857);
nor U14168 (N_14168,N_13946,N_13865);
and U14169 (N_14169,N_13935,N_13846);
nand U14170 (N_14170,N_13889,N_13876);
xor U14171 (N_14171,N_13988,N_13981);
or U14172 (N_14172,N_13913,N_13995);
and U14173 (N_14173,N_13868,N_13850);
nor U14174 (N_14174,N_13940,N_13991);
or U14175 (N_14175,N_13905,N_13984);
xnor U14176 (N_14176,N_13935,N_13840);
and U14177 (N_14177,N_13855,N_13889);
or U14178 (N_14178,N_13831,N_13983);
nand U14179 (N_14179,N_13881,N_13971);
nand U14180 (N_14180,N_13808,N_13809);
and U14181 (N_14181,N_13859,N_13997);
or U14182 (N_14182,N_13995,N_13945);
and U14183 (N_14183,N_13820,N_13980);
and U14184 (N_14184,N_13876,N_13924);
xnor U14185 (N_14185,N_13925,N_13936);
or U14186 (N_14186,N_13819,N_13995);
and U14187 (N_14187,N_13968,N_13838);
or U14188 (N_14188,N_13830,N_13863);
nand U14189 (N_14189,N_13961,N_13872);
xor U14190 (N_14190,N_13829,N_13813);
or U14191 (N_14191,N_13986,N_13969);
xnor U14192 (N_14192,N_13847,N_13979);
or U14193 (N_14193,N_13988,N_13959);
or U14194 (N_14194,N_13989,N_13906);
or U14195 (N_14195,N_13978,N_13806);
xnor U14196 (N_14196,N_13963,N_13985);
xor U14197 (N_14197,N_13935,N_13834);
xor U14198 (N_14198,N_13974,N_13829);
xor U14199 (N_14199,N_13846,N_13854);
nor U14200 (N_14200,N_14195,N_14182);
and U14201 (N_14201,N_14197,N_14146);
or U14202 (N_14202,N_14173,N_14000);
nor U14203 (N_14203,N_14069,N_14123);
xnor U14204 (N_14204,N_14142,N_14044);
or U14205 (N_14205,N_14127,N_14003);
or U14206 (N_14206,N_14138,N_14095);
nand U14207 (N_14207,N_14009,N_14167);
nand U14208 (N_14208,N_14007,N_14184);
or U14209 (N_14209,N_14178,N_14040);
nand U14210 (N_14210,N_14104,N_14109);
nor U14211 (N_14211,N_14191,N_14059);
xor U14212 (N_14212,N_14168,N_14068);
or U14213 (N_14213,N_14198,N_14090);
nand U14214 (N_14214,N_14033,N_14015);
and U14215 (N_14215,N_14112,N_14042);
nand U14216 (N_14216,N_14154,N_14099);
nand U14217 (N_14217,N_14058,N_14190);
or U14218 (N_14218,N_14005,N_14031);
nor U14219 (N_14219,N_14083,N_14077);
nor U14220 (N_14220,N_14103,N_14027);
nor U14221 (N_14221,N_14110,N_14125);
or U14222 (N_14222,N_14091,N_14049);
or U14223 (N_14223,N_14194,N_14171);
or U14224 (N_14224,N_14081,N_14012);
nand U14225 (N_14225,N_14126,N_14183);
nor U14226 (N_14226,N_14078,N_14010);
and U14227 (N_14227,N_14017,N_14115);
xor U14228 (N_14228,N_14124,N_14045);
and U14229 (N_14229,N_14075,N_14021);
nor U14230 (N_14230,N_14151,N_14163);
nor U14231 (N_14231,N_14016,N_14144);
nor U14232 (N_14232,N_14051,N_14067);
xor U14233 (N_14233,N_14189,N_14092);
xnor U14234 (N_14234,N_14047,N_14166);
nor U14235 (N_14235,N_14065,N_14120);
xor U14236 (N_14236,N_14041,N_14032);
xnor U14237 (N_14237,N_14038,N_14175);
or U14238 (N_14238,N_14094,N_14176);
nor U14239 (N_14239,N_14193,N_14076);
nor U14240 (N_14240,N_14004,N_14122);
and U14241 (N_14241,N_14172,N_14119);
nand U14242 (N_14242,N_14048,N_14139);
nand U14243 (N_14243,N_14085,N_14035);
and U14244 (N_14244,N_14088,N_14046);
nand U14245 (N_14245,N_14006,N_14147);
and U14246 (N_14246,N_14158,N_14188);
nor U14247 (N_14247,N_14159,N_14150);
nand U14248 (N_14248,N_14155,N_14029);
and U14249 (N_14249,N_14162,N_14179);
xnor U14250 (N_14250,N_14084,N_14072);
xnor U14251 (N_14251,N_14026,N_14028);
xor U14252 (N_14252,N_14101,N_14140);
or U14253 (N_14253,N_14199,N_14066);
nor U14254 (N_14254,N_14060,N_14023);
nor U14255 (N_14255,N_14100,N_14114);
or U14256 (N_14256,N_14131,N_14113);
or U14257 (N_14257,N_14054,N_14050);
nand U14258 (N_14258,N_14071,N_14129);
or U14259 (N_14259,N_14011,N_14108);
nand U14260 (N_14260,N_14022,N_14160);
nand U14261 (N_14261,N_14014,N_14082);
nand U14262 (N_14262,N_14153,N_14096);
xor U14263 (N_14263,N_14061,N_14079);
xnor U14264 (N_14264,N_14008,N_14118);
and U14265 (N_14265,N_14148,N_14002);
or U14266 (N_14266,N_14052,N_14025);
nor U14267 (N_14267,N_14106,N_14013);
nand U14268 (N_14268,N_14143,N_14020);
nor U14269 (N_14269,N_14098,N_14001);
and U14270 (N_14270,N_14161,N_14117);
xnor U14271 (N_14271,N_14057,N_14039);
xnor U14272 (N_14272,N_14174,N_14141);
xnor U14273 (N_14273,N_14064,N_14185);
xnor U14274 (N_14274,N_14105,N_14024);
nand U14275 (N_14275,N_14102,N_14133);
nor U14276 (N_14276,N_14137,N_14177);
or U14277 (N_14277,N_14107,N_14055);
and U14278 (N_14278,N_14130,N_14019);
or U14279 (N_14279,N_14097,N_14121);
or U14280 (N_14280,N_14063,N_14053);
nor U14281 (N_14281,N_14156,N_14132);
and U14282 (N_14282,N_14186,N_14111);
and U14283 (N_14283,N_14056,N_14116);
nand U14284 (N_14284,N_14062,N_14145);
xnor U14285 (N_14285,N_14037,N_14165);
and U14286 (N_14286,N_14170,N_14187);
nand U14287 (N_14287,N_14074,N_14086);
nand U14288 (N_14288,N_14087,N_14036);
xnor U14289 (N_14289,N_14030,N_14135);
nor U14290 (N_14290,N_14070,N_14169);
and U14291 (N_14291,N_14136,N_14073);
nor U14292 (N_14292,N_14134,N_14080);
and U14293 (N_14293,N_14149,N_14164);
or U14294 (N_14294,N_14043,N_14196);
and U14295 (N_14295,N_14181,N_14192);
or U14296 (N_14296,N_14180,N_14157);
nor U14297 (N_14297,N_14034,N_14018);
nor U14298 (N_14298,N_14152,N_14089);
nand U14299 (N_14299,N_14128,N_14093);
or U14300 (N_14300,N_14033,N_14128);
xor U14301 (N_14301,N_14166,N_14096);
or U14302 (N_14302,N_14141,N_14099);
nand U14303 (N_14303,N_14193,N_14114);
and U14304 (N_14304,N_14049,N_14143);
or U14305 (N_14305,N_14066,N_14036);
or U14306 (N_14306,N_14019,N_14119);
and U14307 (N_14307,N_14106,N_14170);
xor U14308 (N_14308,N_14078,N_14077);
and U14309 (N_14309,N_14011,N_14107);
or U14310 (N_14310,N_14092,N_14136);
nand U14311 (N_14311,N_14107,N_14057);
nand U14312 (N_14312,N_14023,N_14128);
xnor U14313 (N_14313,N_14075,N_14195);
and U14314 (N_14314,N_14198,N_14087);
or U14315 (N_14315,N_14130,N_14151);
xnor U14316 (N_14316,N_14096,N_14065);
or U14317 (N_14317,N_14002,N_14059);
and U14318 (N_14318,N_14153,N_14026);
xor U14319 (N_14319,N_14141,N_14170);
and U14320 (N_14320,N_14183,N_14051);
and U14321 (N_14321,N_14087,N_14150);
or U14322 (N_14322,N_14004,N_14078);
nand U14323 (N_14323,N_14154,N_14062);
xnor U14324 (N_14324,N_14146,N_14046);
nand U14325 (N_14325,N_14007,N_14157);
or U14326 (N_14326,N_14109,N_14023);
or U14327 (N_14327,N_14191,N_14025);
xor U14328 (N_14328,N_14196,N_14004);
and U14329 (N_14329,N_14039,N_14139);
xnor U14330 (N_14330,N_14038,N_14018);
nand U14331 (N_14331,N_14131,N_14041);
or U14332 (N_14332,N_14003,N_14107);
xnor U14333 (N_14333,N_14104,N_14118);
xnor U14334 (N_14334,N_14162,N_14139);
nand U14335 (N_14335,N_14194,N_14169);
nor U14336 (N_14336,N_14071,N_14036);
or U14337 (N_14337,N_14125,N_14173);
nand U14338 (N_14338,N_14156,N_14136);
and U14339 (N_14339,N_14136,N_14077);
nand U14340 (N_14340,N_14133,N_14192);
or U14341 (N_14341,N_14174,N_14199);
or U14342 (N_14342,N_14155,N_14095);
xor U14343 (N_14343,N_14012,N_14120);
nand U14344 (N_14344,N_14041,N_14079);
nand U14345 (N_14345,N_14010,N_14023);
nand U14346 (N_14346,N_14109,N_14021);
or U14347 (N_14347,N_14078,N_14000);
nor U14348 (N_14348,N_14151,N_14093);
xor U14349 (N_14349,N_14070,N_14073);
or U14350 (N_14350,N_14165,N_14098);
or U14351 (N_14351,N_14126,N_14007);
nand U14352 (N_14352,N_14178,N_14165);
nor U14353 (N_14353,N_14151,N_14196);
and U14354 (N_14354,N_14025,N_14185);
and U14355 (N_14355,N_14106,N_14178);
nor U14356 (N_14356,N_14178,N_14037);
xor U14357 (N_14357,N_14102,N_14063);
nor U14358 (N_14358,N_14105,N_14134);
xor U14359 (N_14359,N_14186,N_14080);
and U14360 (N_14360,N_14178,N_14060);
or U14361 (N_14361,N_14000,N_14135);
xnor U14362 (N_14362,N_14049,N_14040);
and U14363 (N_14363,N_14078,N_14132);
nor U14364 (N_14364,N_14024,N_14030);
nand U14365 (N_14365,N_14133,N_14054);
nor U14366 (N_14366,N_14115,N_14135);
and U14367 (N_14367,N_14018,N_14157);
and U14368 (N_14368,N_14185,N_14015);
xnor U14369 (N_14369,N_14056,N_14194);
or U14370 (N_14370,N_14122,N_14104);
xnor U14371 (N_14371,N_14091,N_14060);
nor U14372 (N_14372,N_14038,N_14002);
xor U14373 (N_14373,N_14117,N_14085);
nor U14374 (N_14374,N_14155,N_14017);
xnor U14375 (N_14375,N_14183,N_14114);
nor U14376 (N_14376,N_14169,N_14178);
nor U14377 (N_14377,N_14074,N_14009);
nand U14378 (N_14378,N_14016,N_14155);
nand U14379 (N_14379,N_14159,N_14108);
nand U14380 (N_14380,N_14138,N_14058);
xor U14381 (N_14381,N_14114,N_14142);
xnor U14382 (N_14382,N_14192,N_14198);
xnor U14383 (N_14383,N_14015,N_14197);
nor U14384 (N_14384,N_14096,N_14191);
and U14385 (N_14385,N_14152,N_14003);
xnor U14386 (N_14386,N_14078,N_14199);
and U14387 (N_14387,N_14016,N_14105);
nor U14388 (N_14388,N_14017,N_14143);
or U14389 (N_14389,N_14065,N_14070);
nor U14390 (N_14390,N_14035,N_14115);
xor U14391 (N_14391,N_14050,N_14039);
xnor U14392 (N_14392,N_14186,N_14183);
xnor U14393 (N_14393,N_14037,N_14010);
nand U14394 (N_14394,N_14126,N_14176);
nand U14395 (N_14395,N_14198,N_14114);
nor U14396 (N_14396,N_14177,N_14034);
xor U14397 (N_14397,N_14139,N_14115);
or U14398 (N_14398,N_14183,N_14028);
or U14399 (N_14399,N_14167,N_14078);
xor U14400 (N_14400,N_14296,N_14209);
nor U14401 (N_14401,N_14364,N_14263);
and U14402 (N_14402,N_14337,N_14267);
and U14403 (N_14403,N_14285,N_14268);
or U14404 (N_14404,N_14336,N_14358);
xnor U14405 (N_14405,N_14314,N_14353);
nor U14406 (N_14406,N_14228,N_14241);
nor U14407 (N_14407,N_14207,N_14389);
or U14408 (N_14408,N_14231,N_14261);
and U14409 (N_14409,N_14227,N_14375);
xnor U14410 (N_14410,N_14213,N_14303);
or U14411 (N_14411,N_14334,N_14351);
or U14412 (N_14412,N_14275,N_14370);
nand U14413 (N_14413,N_14210,N_14352);
or U14414 (N_14414,N_14206,N_14244);
xnor U14415 (N_14415,N_14248,N_14317);
nand U14416 (N_14416,N_14309,N_14297);
and U14417 (N_14417,N_14237,N_14324);
and U14418 (N_14418,N_14325,N_14392);
or U14419 (N_14419,N_14327,N_14279);
xor U14420 (N_14420,N_14382,N_14270);
and U14421 (N_14421,N_14239,N_14251);
or U14422 (N_14422,N_14211,N_14347);
nand U14423 (N_14423,N_14362,N_14259);
nor U14424 (N_14424,N_14319,N_14283);
nand U14425 (N_14425,N_14288,N_14242);
or U14426 (N_14426,N_14376,N_14346);
nand U14427 (N_14427,N_14258,N_14233);
and U14428 (N_14428,N_14315,N_14274);
or U14429 (N_14429,N_14257,N_14374);
xnor U14430 (N_14430,N_14255,N_14322);
and U14431 (N_14431,N_14373,N_14371);
nor U14432 (N_14432,N_14215,N_14217);
xnor U14433 (N_14433,N_14218,N_14264);
or U14434 (N_14434,N_14365,N_14243);
or U14435 (N_14435,N_14273,N_14342);
nand U14436 (N_14436,N_14338,N_14304);
or U14437 (N_14437,N_14223,N_14333);
and U14438 (N_14438,N_14311,N_14294);
or U14439 (N_14439,N_14398,N_14286);
nor U14440 (N_14440,N_14205,N_14356);
or U14441 (N_14441,N_14256,N_14219);
or U14442 (N_14442,N_14203,N_14368);
xor U14443 (N_14443,N_14226,N_14341);
and U14444 (N_14444,N_14230,N_14277);
and U14445 (N_14445,N_14282,N_14320);
xor U14446 (N_14446,N_14299,N_14369);
and U14447 (N_14447,N_14378,N_14349);
and U14448 (N_14448,N_14202,N_14235);
nand U14449 (N_14449,N_14381,N_14220);
xnor U14450 (N_14450,N_14359,N_14212);
xnor U14451 (N_14451,N_14348,N_14271);
xor U14452 (N_14452,N_14272,N_14387);
nand U14453 (N_14453,N_14312,N_14329);
xor U14454 (N_14454,N_14254,N_14379);
nor U14455 (N_14455,N_14276,N_14383);
nand U14456 (N_14456,N_14253,N_14236);
xnor U14457 (N_14457,N_14344,N_14224);
nor U14458 (N_14458,N_14214,N_14308);
nand U14459 (N_14459,N_14372,N_14302);
xnor U14460 (N_14460,N_14245,N_14395);
nand U14461 (N_14461,N_14350,N_14246);
or U14462 (N_14462,N_14307,N_14295);
nand U14463 (N_14463,N_14269,N_14366);
nor U14464 (N_14464,N_14355,N_14291);
nand U14465 (N_14465,N_14247,N_14396);
and U14466 (N_14466,N_14225,N_14326);
or U14467 (N_14467,N_14284,N_14301);
or U14468 (N_14468,N_14280,N_14332);
and U14469 (N_14469,N_14345,N_14377);
and U14470 (N_14470,N_14361,N_14232);
nand U14471 (N_14471,N_14278,N_14208);
xor U14472 (N_14472,N_14204,N_14363);
or U14473 (N_14473,N_14354,N_14250);
xor U14474 (N_14474,N_14229,N_14399);
and U14475 (N_14475,N_14343,N_14265);
or U14476 (N_14476,N_14384,N_14238);
and U14477 (N_14477,N_14281,N_14260);
nor U14478 (N_14478,N_14252,N_14249);
nor U14479 (N_14479,N_14201,N_14390);
or U14480 (N_14480,N_14330,N_14318);
and U14481 (N_14481,N_14290,N_14298);
and U14482 (N_14482,N_14340,N_14339);
and U14483 (N_14483,N_14310,N_14300);
xor U14484 (N_14484,N_14240,N_14380);
xnor U14485 (N_14485,N_14287,N_14385);
nor U14486 (N_14486,N_14234,N_14313);
nand U14487 (N_14487,N_14357,N_14391);
nand U14488 (N_14488,N_14321,N_14360);
nand U14489 (N_14489,N_14305,N_14293);
or U14490 (N_14490,N_14222,N_14262);
xnor U14491 (N_14491,N_14335,N_14323);
and U14492 (N_14492,N_14328,N_14292);
nand U14493 (N_14493,N_14367,N_14216);
xnor U14494 (N_14494,N_14394,N_14331);
xnor U14495 (N_14495,N_14316,N_14388);
or U14496 (N_14496,N_14289,N_14266);
xnor U14497 (N_14497,N_14200,N_14393);
nand U14498 (N_14498,N_14386,N_14306);
and U14499 (N_14499,N_14397,N_14221);
or U14500 (N_14500,N_14219,N_14245);
and U14501 (N_14501,N_14275,N_14204);
nand U14502 (N_14502,N_14367,N_14289);
nand U14503 (N_14503,N_14371,N_14384);
nand U14504 (N_14504,N_14246,N_14268);
and U14505 (N_14505,N_14397,N_14207);
xor U14506 (N_14506,N_14284,N_14371);
nand U14507 (N_14507,N_14370,N_14378);
nand U14508 (N_14508,N_14356,N_14287);
xor U14509 (N_14509,N_14376,N_14219);
nand U14510 (N_14510,N_14378,N_14245);
nor U14511 (N_14511,N_14322,N_14222);
nand U14512 (N_14512,N_14296,N_14360);
xor U14513 (N_14513,N_14216,N_14312);
nand U14514 (N_14514,N_14386,N_14344);
and U14515 (N_14515,N_14304,N_14221);
or U14516 (N_14516,N_14353,N_14334);
or U14517 (N_14517,N_14282,N_14233);
xor U14518 (N_14518,N_14210,N_14304);
and U14519 (N_14519,N_14380,N_14333);
and U14520 (N_14520,N_14336,N_14369);
and U14521 (N_14521,N_14393,N_14270);
or U14522 (N_14522,N_14362,N_14274);
and U14523 (N_14523,N_14325,N_14234);
and U14524 (N_14524,N_14319,N_14201);
nor U14525 (N_14525,N_14272,N_14374);
nor U14526 (N_14526,N_14232,N_14230);
nand U14527 (N_14527,N_14250,N_14252);
nor U14528 (N_14528,N_14205,N_14233);
and U14529 (N_14529,N_14377,N_14251);
nor U14530 (N_14530,N_14356,N_14243);
xor U14531 (N_14531,N_14259,N_14395);
nor U14532 (N_14532,N_14305,N_14336);
and U14533 (N_14533,N_14210,N_14263);
nand U14534 (N_14534,N_14239,N_14309);
xnor U14535 (N_14535,N_14228,N_14385);
nand U14536 (N_14536,N_14397,N_14272);
nor U14537 (N_14537,N_14373,N_14352);
or U14538 (N_14538,N_14362,N_14267);
xnor U14539 (N_14539,N_14223,N_14317);
nor U14540 (N_14540,N_14226,N_14357);
nor U14541 (N_14541,N_14213,N_14308);
and U14542 (N_14542,N_14267,N_14221);
or U14543 (N_14543,N_14203,N_14284);
nand U14544 (N_14544,N_14359,N_14345);
nand U14545 (N_14545,N_14312,N_14301);
nand U14546 (N_14546,N_14204,N_14289);
and U14547 (N_14547,N_14385,N_14227);
nand U14548 (N_14548,N_14326,N_14361);
nand U14549 (N_14549,N_14373,N_14334);
nand U14550 (N_14550,N_14226,N_14306);
or U14551 (N_14551,N_14363,N_14371);
nor U14552 (N_14552,N_14391,N_14377);
xor U14553 (N_14553,N_14238,N_14381);
and U14554 (N_14554,N_14384,N_14301);
and U14555 (N_14555,N_14376,N_14356);
or U14556 (N_14556,N_14318,N_14289);
and U14557 (N_14557,N_14311,N_14234);
nand U14558 (N_14558,N_14308,N_14356);
or U14559 (N_14559,N_14243,N_14207);
nand U14560 (N_14560,N_14281,N_14206);
or U14561 (N_14561,N_14321,N_14233);
xnor U14562 (N_14562,N_14278,N_14251);
nor U14563 (N_14563,N_14265,N_14283);
nor U14564 (N_14564,N_14211,N_14362);
and U14565 (N_14565,N_14238,N_14318);
nand U14566 (N_14566,N_14290,N_14254);
nand U14567 (N_14567,N_14306,N_14219);
or U14568 (N_14568,N_14211,N_14226);
and U14569 (N_14569,N_14354,N_14398);
nand U14570 (N_14570,N_14213,N_14320);
xor U14571 (N_14571,N_14308,N_14390);
nor U14572 (N_14572,N_14201,N_14250);
nor U14573 (N_14573,N_14387,N_14217);
nand U14574 (N_14574,N_14305,N_14227);
xnor U14575 (N_14575,N_14224,N_14299);
nand U14576 (N_14576,N_14318,N_14309);
nor U14577 (N_14577,N_14293,N_14232);
or U14578 (N_14578,N_14224,N_14372);
xor U14579 (N_14579,N_14332,N_14352);
nor U14580 (N_14580,N_14376,N_14238);
xor U14581 (N_14581,N_14353,N_14326);
and U14582 (N_14582,N_14226,N_14354);
nand U14583 (N_14583,N_14275,N_14229);
nand U14584 (N_14584,N_14265,N_14379);
xnor U14585 (N_14585,N_14399,N_14344);
xnor U14586 (N_14586,N_14396,N_14286);
nand U14587 (N_14587,N_14296,N_14254);
or U14588 (N_14588,N_14344,N_14357);
and U14589 (N_14589,N_14330,N_14297);
xor U14590 (N_14590,N_14298,N_14378);
or U14591 (N_14591,N_14205,N_14308);
and U14592 (N_14592,N_14387,N_14201);
nand U14593 (N_14593,N_14353,N_14229);
xor U14594 (N_14594,N_14260,N_14216);
nor U14595 (N_14595,N_14383,N_14351);
nand U14596 (N_14596,N_14362,N_14308);
xor U14597 (N_14597,N_14256,N_14358);
and U14598 (N_14598,N_14320,N_14338);
and U14599 (N_14599,N_14399,N_14222);
or U14600 (N_14600,N_14556,N_14406);
and U14601 (N_14601,N_14416,N_14410);
nand U14602 (N_14602,N_14471,N_14475);
nor U14603 (N_14603,N_14530,N_14512);
and U14604 (N_14604,N_14505,N_14426);
nand U14605 (N_14605,N_14496,N_14460);
or U14606 (N_14606,N_14465,N_14545);
nand U14607 (N_14607,N_14594,N_14578);
nand U14608 (N_14608,N_14534,N_14543);
or U14609 (N_14609,N_14504,N_14486);
or U14610 (N_14610,N_14470,N_14519);
nand U14611 (N_14611,N_14569,N_14559);
nand U14612 (N_14612,N_14516,N_14452);
xor U14613 (N_14613,N_14518,N_14520);
nor U14614 (N_14614,N_14405,N_14571);
or U14615 (N_14615,N_14595,N_14531);
nor U14616 (N_14616,N_14541,N_14501);
xnor U14617 (N_14617,N_14533,N_14549);
nor U14618 (N_14618,N_14523,N_14548);
nand U14619 (N_14619,N_14438,N_14529);
nand U14620 (N_14620,N_14437,N_14482);
and U14621 (N_14621,N_14420,N_14575);
xor U14622 (N_14622,N_14400,N_14440);
xor U14623 (N_14623,N_14444,N_14478);
or U14624 (N_14624,N_14493,N_14542);
nor U14625 (N_14625,N_14461,N_14506);
xnor U14626 (N_14626,N_14587,N_14536);
nor U14627 (N_14627,N_14586,N_14490);
xor U14628 (N_14628,N_14417,N_14443);
xor U14629 (N_14629,N_14450,N_14430);
nor U14630 (N_14630,N_14418,N_14407);
or U14631 (N_14631,N_14579,N_14561);
nor U14632 (N_14632,N_14599,N_14422);
xor U14633 (N_14633,N_14458,N_14421);
xor U14634 (N_14634,N_14435,N_14564);
nor U14635 (N_14635,N_14546,N_14597);
or U14636 (N_14636,N_14509,N_14591);
nand U14637 (N_14637,N_14483,N_14466);
xor U14638 (N_14638,N_14585,N_14442);
or U14639 (N_14639,N_14491,N_14557);
and U14640 (N_14640,N_14596,N_14484);
nand U14641 (N_14641,N_14558,N_14473);
nor U14642 (N_14642,N_14551,N_14414);
xor U14643 (N_14643,N_14547,N_14429);
nor U14644 (N_14644,N_14412,N_14521);
or U14645 (N_14645,N_14485,N_14565);
or U14646 (N_14646,N_14574,N_14580);
or U14647 (N_14647,N_14581,N_14446);
xnor U14648 (N_14648,N_14495,N_14507);
xor U14649 (N_14649,N_14566,N_14497);
nor U14650 (N_14650,N_14572,N_14488);
and U14651 (N_14651,N_14477,N_14514);
xor U14652 (N_14652,N_14456,N_14563);
nor U14653 (N_14653,N_14423,N_14502);
or U14654 (N_14654,N_14498,N_14472);
and U14655 (N_14655,N_14553,N_14582);
xor U14656 (N_14656,N_14489,N_14526);
nand U14657 (N_14657,N_14481,N_14469);
nand U14658 (N_14658,N_14439,N_14499);
nor U14659 (N_14659,N_14448,N_14419);
xor U14660 (N_14660,N_14589,N_14570);
and U14661 (N_14661,N_14455,N_14451);
nor U14662 (N_14662,N_14598,N_14508);
xnor U14663 (N_14663,N_14517,N_14464);
and U14664 (N_14664,N_14434,N_14590);
and U14665 (N_14665,N_14402,N_14428);
and U14666 (N_14666,N_14528,N_14513);
or U14667 (N_14667,N_14447,N_14568);
xor U14668 (N_14668,N_14463,N_14424);
xor U14669 (N_14669,N_14515,N_14411);
nor U14670 (N_14670,N_14593,N_14492);
xor U14671 (N_14671,N_14583,N_14474);
and U14672 (N_14672,N_14560,N_14449);
and U14673 (N_14673,N_14433,N_14487);
nor U14674 (N_14674,N_14436,N_14408);
nor U14675 (N_14675,N_14540,N_14539);
nor U14676 (N_14676,N_14432,N_14404);
and U14677 (N_14677,N_14401,N_14550);
and U14678 (N_14678,N_14573,N_14544);
nor U14679 (N_14679,N_14476,N_14552);
or U14680 (N_14680,N_14535,N_14441);
xor U14681 (N_14681,N_14527,N_14524);
nor U14682 (N_14682,N_14522,N_14500);
and U14683 (N_14683,N_14588,N_14413);
xor U14684 (N_14684,N_14457,N_14494);
and U14685 (N_14685,N_14525,N_14425);
and U14686 (N_14686,N_14453,N_14567);
and U14687 (N_14687,N_14576,N_14467);
and U14688 (N_14688,N_14415,N_14468);
xnor U14689 (N_14689,N_14409,N_14592);
or U14690 (N_14690,N_14445,N_14510);
nand U14691 (N_14691,N_14479,N_14537);
nor U14692 (N_14692,N_14554,N_14511);
xor U14693 (N_14693,N_14459,N_14454);
xor U14694 (N_14694,N_14503,N_14584);
xor U14695 (N_14695,N_14427,N_14555);
and U14696 (N_14696,N_14532,N_14431);
and U14697 (N_14697,N_14577,N_14562);
xnor U14698 (N_14698,N_14462,N_14538);
xnor U14699 (N_14699,N_14480,N_14403);
nand U14700 (N_14700,N_14526,N_14577);
or U14701 (N_14701,N_14513,N_14453);
xor U14702 (N_14702,N_14460,N_14401);
xnor U14703 (N_14703,N_14585,N_14577);
or U14704 (N_14704,N_14491,N_14532);
nand U14705 (N_14705,N_14428,N_14466);
xnor U14706 (N_14706,N_14591,N_14563);
or U14707 (N_14707,N_14478,N_14570);
nand U14708 (N_14708,N_14457,N_14418);
or U14709 (N_14709,N_14472,N_14509);
nor U14710 (N_14710,N_14574,N_14569);
or U14711 (N_14711,N_14514,N_14492);
and U14712 (N_14712,N_14454,N_14478);
nand U14713 (N_14713,N_14406,N_14509);
and U14714 (N_14714,N_14415,N_14472);
and U14715 (N_14715,N_14539,N_14489);
nor U14716 (N_14716,N_14531,N_14496);
or U14717 (N_14717,N_14427,N_14497);
xnor U14718 (N_14718,N_14494,N_14445);
nor U14719 (N_14719,N_14549,N_14564);
and U14720 (N_14720,N_14579,N_14529);
xnor U14721 (N_14721,N_14458,N_14413);
and U14722 (N_14722,N_14529,N_14402);
or U14723 (N_14723,N_14463,N_14539);
or U14724 (N_14724,N_14480,N_14593);
nand U14725 (N_14725,N_14534,N_14549);
and U14726 (N_14726,N_14451,N_14545);
and U14727 (N_14727,N_14587,N_14463);
xor U14728 (N_14728,N_14487,N_14486);
or U14729 (N_14729,N_14425,N_14567);
and U14730 (N_14730,N_14409,N_14407);
or U14731 (N_14731,N_14501,N_14586);
and U14732 (N_14732,N_14484,N_14472);
or U14733 (N_14733,N_14499,N_14534);
nand U14734 (N_14734,N_14407,N_14585);
nor U14735 (N_14735,N_14497,N_14507);
nor U14736 (N_14736,N_14570,N_14501);
xor U14737 (N_14737,N_14520,N_14492);
xor U14738 (N_14738,N_14475,N_14489);
nand U14739 (N_14739,N_14590,N_14562);
and U14740 (N_14740,N_14411,N_14427);
nand U14741 (N_14741,N_14442,N_14418);
xnor U14742 (N_14742,N_14593,N_14442);
nor U14743 (N_14743,N_14526,N_14500);
and U14744 (N_14744,N_14551,N_14474);
xor U14745 (N_14745,N_14532,N_14449);
xnor U14746 (N_14746,N_14598,N_14491);
nor U14747 (N_14747,N_14471,N_14444);
xor U14748 (N_14748,N_14423,N_14476);
and U14749 (N_14749,N_14556,N_14430);
xnor U14750 (N_14750,N_14594,N_14479);
nor U14751 (N_14751,N_14439,N_14473);
nand U14752 (N_14752,N_14433,N_14515);
xor U14753 (N_14753,N_14568,N_14440);
nand U14754 (N_14754,N_14471,N_14585);
and U14755 (N_14755,N_14425,N_14472);
xnor U14756 (N_14756,N_14487,N_14568);
xor U14757 (N_14757,N_14481,N_14443);
xnor U14758 (N_14758,N_14590,N_14405);
or U14759 (N_14759,N_14497,N_14406);
or U14760 (N_14760,N_14564,N_14480);
nand U14761 (N_14761,N_14512,N_14583);
xor U14762 (N_14762,N_14558,N_14405);
nor U14763 (N_14763,N_14482,N_14549);
nand U14764 (N_14764,N_14450,N_14592);
or U14765 (N_14765,N_14464,N_14470);
and U14766 (N_14766,N_14572,N_14523);
xnor U14767 (N_14767,N_14426,N_14532);
and U14768 (N_14768,N_14484,N_14586);
and U14769 (N_14769,N_14414,N_14493);
nand U14770 (N_14770,N_14541,N_14498);
xor U14771 (N_14771,N_14400,N_14599);
and U14772 (N_14772,N_14487,N_14494);
or U14773 (N_14773,N_14571,N_14552);
nor U14774 (N_14774,N_14427,N_14570);
and U14775 (N_14775,N_14545,N_14565);
and U14776 (N_14776,N_14513,N_14462);
nor U14777 (N_14777,N_14530,N_14505);
or U14778 (N_14778,N_14593,N_14471);
nor U14779 (N_14779,N_14417,N_14457);
nor U14780 (N_14780,N_14594,N_14589);
xor U14781 (N_14781,N_14476,N_14569);
nor U14782 (N_14782,N_14533,N_14420);
or U14783 (N_14783,N_14518,N_14461);
or U14784 (N_14784,N_14469,N_14529);
nand U14785 (N_14785,N_14543,N_14563);
nand U14786 (N_14786,N_14521,N_14519);
xor U14787 (N_14787,N_14501,N_14412);
nor U14788 (N_14788,N_14452,N_14524);
nor U14789 (N_14789,N_14495,N_14436);
nor U14790 (N_14790,N_14422,N_14481);
or U14791 (N_14791,N_14425,N_14530);
and U14792 (N_14792,N_14469,N_14435);
nand U14793 (N_14793,N_14547,N_14418);
nand U14794 (N_14794,N_14524,N_14424);
xnor U14795 (N_14795,N_14565,N_14481);
nor U14796 (N_14796,N_14580,N_14516);
nor U14797 (N_14797,N_14477,N_14413);
nor U14798 (N_14798,N_14462,N_14470);
nor U14799 (N_14799,N_14598,N_14558);
nor U14800 (N_14800,N_14647,N_14605);
and U14801 (N_14801,N_14735,N_14793);
and U14802 (N_14802,N_14616,N_14785);
xor U14803 (N_14803,N_14798,N_14671);
nor U14804 (N_14804,N_14757,N_14713);
nor U14805 (N_14805,N_14767,N_14670);
or U14806 (N_14806,N_14669,N_14617);
nor U14807 (N_14807,N_14772,N_14646);
xor U14808 (N_14808,N_14784,N_14660);
xnor U14809 (N_14809,N_14756,N_14708);
or U14810 (N_14810,N_14737,N_14792);
nor U14811 (N_14811,N_14672,N_14739);
nor U14812 (N_14812,N_14736,N_14751);
nand U14813 (N_14813,N_14642,N_14602);
nor U14814 (N_14814,N_14618,N_14782);
nand U14815 (N_14815,N_14733,N_14667);
nand U14816 (N_14816,N_14611,N_14781);
or U14817 (N_14817,N_14765,N_14604);
nor U14818 (N_14818,N_14743,N_14759);
nand U14819 (N_14819,N_14752,N_14710);
and U14820 (N_14820,N_14693,N_14740);
xnor U14821 (N_14821,N_14658,N_14675);
nor U14822 (N_14822,N_14741,N_14609);
nand U14823 (N_14823,N_14632,N_14777);
xor U14824 (N_14824,N_14746,N_14625);
and U14825 (N_14825,N_14721,N_14705);
or U14826 (N_14826,N_14629,N_14718);
nor U14827 (N_14827,N_14698,N_14657);
nor U14828 (N_14828,N_14600,N_14788);
nor U14829 (N_14829,N_14786,N_14783);
or U14830 (N_14830,N_14628,N_14795);
nand U14831 (N_14831,N_14731,N_14796);
or U14832 (N_14832,N_14758,N_14747);
and U14833 (N_14833,N_14653,N_14714);
and U14834 (N_14834,N_14701,N_14779);
xnor U14835 (N_14835,N_14665,N_14794);
nor U14836 (N_14836,N_14601,N_14627);
nor U14837 (N_14837,N_14706,N_14717);
or U14838 (N_14838,N_14734,N_14728);
or U14839 (N_14839,N_14761,N_14732);
nor U14840 (N_14840,N_14656,N_14754);
nor U14841 (N_14841,N_14755,N_14654);
and U14842 (N_14842,N_14711,N_14662);
xor U14843 (N_14843,N_14615,N_14633);
and U14844 (N_14844,N_14787,N_14622);
or U14845 (N_14845,N_14676,N_14624);
xor U14846 (N_14846,N_14635,N_14715);
nor U14847 (N_14847,N_14690,N_14770);
or U14848 (N_14848,N_14655,N_14606);
and U14849 (N_14849,N_14621,N_14695);
or U14850 (N_14850,N_14749,N_14694);
nand U14851 (N_14851,N_14724,N_14607);
xnor U14852 (N_14852,N_14666,N_14688);
xnor U14853 (N_14853,N_14723,N_14742);
or U14854 (N_14854,N_14769,N_14645);
or U14855 (N_14855,N_14610,N_14679);
xnor U14856 (N_14856,N_14644,N_14744);
xor U14857 (N_14857,N_14649,N_14730);
nor U14858 (N_14858,N_14699,N_14614);
and U14859 (N_14859,N_14650,N_14750);
and U14860 (N_14860,N_14683,N_14661);
nand U14861 (N_14861,N_14674,N_14613);
nor U14862 (N_14862,N_14630,N_14641);
and U14863 (N_14863,N_14720,N_14697);
nand U14864 (N_14864,N_14722,N_14678);
nand U14865 (N_14865,N_14764,N_14689);
nand U14866 (N_14866,N_14738,N_14789);
nor U14867 (N_14867,N_14760,N_14775);
or U14868 (N_14868,N_14664,N_14637);
xor U14869 (N_14869,N_14659,N_14780);
xor U14870 (N_14870,N_14640,N_14691);
and U14871 (N_14871,N_14729,N_14677);
nand U14872 (N_14872,N_14623,N_14626);
and U14873 (N_14873,N_14612,N_14725);
nor U14874 (N_14874,N_14643,N_14639);
or U14875 (N_14875,N_14776,N_14703);
nand U14876 (N_14876,N_14763,N_14799);
nand U14877 (N_14877,N_14712,N_14719);
xnor U14878 (N_14878,N_14762,N_14687);
nor U14879 (N_14879,N_14668,N_14636);
or U14880 (N_14880,N_14692,N_14726);
or U14881 (N_14881,N_14704,N_14791);
or U14882 (N_14882,N_14631,N_14709);
and U14883 (N_14883,N_14790,N_14686);
and U14884 (N_14884,N_14608,N_14707);
or U14885 (N_14885,N_14638,N_14745);
nand U14886 (N_14886,N_14652,N_14700);
nor U14887 (N_14887,N_14685,N_14663);
and U14888 (N_14888,N_14603,N_14771);
and U14889 (N_14889,N_14619,N_14684);
and U14890 (N_14890,N_14620,N_14773);
xnor U14891 (N_14891,N_14778,N_14648);
or U14892 (N_14892,N_14702,N_14774);
xnor U14893 (N_14893,N_14716,N_14696);
nand U14894 (N_14894,N_14797,N_14673);
xnor U14895 (N_14895,N_14634,N_14682);
nand U14896 (N_14896,N_14768,N_14766);
nand U14897 (N_14897,N_14680,N_14681);
and U14898 (N_14898,N_14753,N_14651);
nand U14899 (N_14899,N_14727,N_14748);
nor U14900 (N_14900,N_14709,N_14618);
nor U14901 (N_14901,N_14688,N_14684);
xnor U14902 (N_14902,N_14627,N_14747);
xor U14903 (N_14903,N_14796,N_14631);
and U14904 (N_14904,N_14779,N_14736);
nand U14905 (N_14905,N_14653,N_14637);
nand U14906 (N_14906,N_14703,N_14660);
nor U14907 (N_14907,N_14732,N_14649);
nor U14908 (N_14908,N_14718,N_14645);
nor U14909 (N_14909,N_14637,N_14706);
and U14910 (N_14910,N_14715,N_14664);
nor U14911 (N_14911,N_14763,N_14632);
or U14912 (N_14912,N_14788,N_14682);
or U14913 (N_14913,N_14736,N_14628);
or U14914 (N_14914,N_14620,N_14704);
nor U14915 (N_14915,N_14769,N_14787);
nor U14916 (N_14916,N_14692,N_14732);
nand U14917 (N_14917,N_14699,N_14602);
nor U14918 (N_14918,N_14644,N_14787);
nand U14919 (N_14919,N_14615,N_14792);
and U14920 (N_14920,N_14792,N_14748);
and U14921 (N_14921,N_14670,N_14733);
nor U14922 (N_14922,N_14737,N_14783);
or U14923 (N_14923,N_14786,N_14760);
nor U14924 (N_14924,N_14691,N_14604);
nand U14925 (N_14925,N_14725,N_14657);
xnor U14926 (N_14926,N_14738,N_14782);
and U14927 (N_14927,N_14713,N_14633);
nand U14928 (N_14928,N_14773,N_14675);
xnor U14929 (N_14929,N_14707,N_14725);
xor U14930 (N_14930,N_14629,N_14685);
xor U14931 (N_14931,N_14726,N_14729);
and U14932 (N_14932,N_14717,N_14643);
xnor U14933 (N_14933,N_14634,N_14692);
nor U14934 (N_14934,N_14789,N_14731);
xor U14935 (N_14935,N_14796,N_14798);
nand U14936 (N_14936,N_14605,N_14690);
nand U14937 (N_14937,N_14627,N_14671);
or U14938 (N_14938,N_14601,N_14765);
xnor U14939 (N_14939,N_14654,N_14674);
nor U14940 (N_14940,N_14671,N_14649);
and U14941 (N_14941,N_14679,N_14714);
nand U14942 (N_14942,N_14760,N_14674);
nand U14943 (N_14943,N_14612,N_14681);
or U14944 (N_14944,N_14734,N_14752);
nor U14945 (N_14945,N_14737,N_14604);
and U14946 (N_14946,N_14746,N_14761);
and U14947 (N_14947,N_14786,N_14799);
or U14948 (N_14948,N_14710,N_14604);
nand U14949 (N_14949,N_14766,N_14634);
nor U14950 (N_14950,N_14600,N_14701);
nand U14951 (N_14951,N_14611,N_14799);
xnor U14952 (N_14952,N_14707,N_14613);
and U14953 (N_14953,N_14777,N_14606);
nand U14954 (N_14954,N_14676,N_14747);
nor U14955 (N_14955,N_14675,N_14781);
nor U14956 (N_14956,N_14603,N_14693);
or U14957 (N_14957,N_14610,N_14790);
xor U14958 (N_14958,N_14602,N_14777);
xor U14959 (N_14959,N_14678,N_14721);
nand U14960 (N_14960,N_14763,N_14635);
or U14961 (N_14961,N_14733,N_14606);
and U14962 (N_14962,N_14739,N_14783);
xor U14963 (N_14963,N_14667,N_14680);
xnor U14964 (N_14964,N_14688,N_14752);
or U14965 (N_14965,N_14697,N_14785);
xor U14966 (N_14966,N_14799,N_14713);
or U14967 (N_14967,N_14604,N_14718);
nor U14968 (N_14968,N_14766,N_14696);
and U14969 (N_14969,N_14631,N_14777);
xnor U14970 (N_14970,N_14602,N_14679);
xor U14971 (N_14971,N_14749,N_14678);
or U14972 (N_14972,N_14782,N_14656);
or U14973 (N_14973,N_14719,N_14645);
and U14974 (N_14974,N_14620,N_14769);
or U14975 (N_14975,N_14788,N_14649);
nor U14976 (N_14976,N_14742,N_14710);
nand U14977 (N_14977,N_14786,N_14759);
nand U14978 (N_14978,N_14648,N_14784);
and U14979 (N_14979,N_14673,N_14732);
or U14980 (N_14980,N_14723,N_14638);
nand U14981 (N_14981,N_14678,N_14635);
nand U14982 (N_14982,N_14777,N_14692);
and U14983 (N_14983,N_14600,N_14666);
xnor U14984 (N_14984,N_14765,N_14794);
nor U14985 (N_14985,N_14674,N_14605);
or U14986 (N_14986,N_14672,N_14728);
nand U14987 (N_14987,N_14622,N_14779);
nand U14988 (N_14988,N_14648,N_14689);
nand U14989 (N_14989,N_14631,N_14714);
xor U14990 (N_14990,N_14698,N_14717);
or U14991 (N_14991,N_14736,N_14682);
xnor U14992 (N_14992,N_14685,N_14683);
nand U14993 (N_14993,N_14639,N_14615);
nor U14994 (N_14994,N_14641,N_14779);
nand U14995 (N_14995,N_14736,N_14610);
and U14996 (N_14996,N_14743,N_14688);
and U14997 (N_14997,N_14735,N_14684);
nor U14998 (N_14998,N_14678,N_14650);
and U14999 (N_14999,N_14614,N_14698);
and U15000 (N_15000,N_14815,N_14857);
xnor U15001 (N_15001,N_14985,N_14922);
and U15002 (N_15002,N_14990,N_14976);
or U15003 (N_15003,N_14882,N_14996);
nand U15004 (N_15004,N_14884,N_14819);
and U15005 (N_15005,N_14860,N_14868);
or U15006 (N_15006,N_14864,N_14944);
nand U15007 (N_15007,N_14973,N_14850);
nor U15008 (N_15008,N_14945,N_14871);
and U15009 (N_15009,N_14911,N_14998);
and U15010 (N_15010,N_14852,N_14994);
or U15011 (N_15011,N_14873,N_14942);
or U15012 (N_15012,N_14925,N_14967);
nand U15013 (N_15013,N_14977,N_14935);
or U15014 (N_15014,N_14965,N_14903);
or U15015 (N_15015,N_14889,N_14997);
and U15016 (N_15016,N_14824,N_14934);
and U15017 (N_15017,N_14837,N_14877);
nand U15018 (N_15018,N_14825,N_14827);
nor U15019 (N_15019,N_14964,N_14806);
nor U15020 (N_15020,N_14839,N_14954);
and U15021 (N_15021,N_14817,N_14905);
nor U15022 (N_15022,N_14875,N_14854);
and U15023 (N_15023,N_14890,N_14895);
xor U15024 (N_15024,N_14855,N_14993);
xor U15025 (N_15025,N_14948,N_14943);
or U15026 (N_15026,N_14972,N_14823);
and U15027 (N_15027,N_14816,N_14874);
or U15028 (N_15028,N_14955,N_14908);
or U15029 (N_15029,N_14926,N_14931);
or U15030 (N_15030,N_14963,N_14933);
or U15031 (N_15031,N_14856,N_14947);
and U15032 (N_15032,N_14863,N_14888);
nand U15033 (N_15033,N_14891,N_14941);
or U15034 (N_15034,N_14983,N_14896);
nor U15035 (N_15035,N_14961,N_14845);
nand U15036 (N_15036,N_14840,N_14807);
and U15037 (N_15037,N_14921,N_14865);
nor U15038 (N_15038,N_14986,N_14966);
nand U15039 (N_15039,N_14880,N_14887);
nand U15040 (N_15040,N_14894,N_14907);
or U15041 (N_15041,N_14915,N_14960);
nor U15042 (N_15042,N_14851,N_14987);
and U15043 (N_15043,N_14927,N_14870);
and U15044 (N_15044,N_14917,N_14821);
nor U15045 (N_15045,N_14900,N_14812);
or U15046 (N_15046,N_14968,N_14971);
or U15047 (N_15047,N_14952,N_14876);
nand U15048 (N_15048,N_14958,N_14918);
and U15049 (N_15049,N_14978,N_14841);
nand U15050 (N_15050,N_14909,N_14859);
and U15051 (N_15051,N_14835,N_14809);
nand U15052 (N_15052,N_14975,N_14910);
and U15053 (N_15053,N_14897,N_14881);
or U15054 (N_15054,N_14829,N_14898);
and U15055 (N_15055,N_14962,N_14867);
nor U15056 (N_15056,N_14847,N_14802);
nor U15057 (N_15057,N_14879,N_14801);
and U15058 (N_15058,N_14886,N_14979);
or U15059 (N_15059,N_14995,N_14937);
and U15060 (N_15060,N_14842,N_14822);
nand U15061 (N_15061,N_14813,N_14901);
xor U15062 (N_15062,N_14970,N_14981);
or U15063 (N_15063,N_14833,N_14883);
nor U15064 (N_15064,N_14949,N_14866);
nand U15065 (N_15065,N_14808,N_14902);
xnor U15066 (N_15066,N_14853,N_14928);
xnor U15067 (N_15067,N_14938,N_14916);
xnor U15068 (N_15068,N_14930,N_14820);
nor U15069 (N_15069,N_14858,N_14885);
nand U15070 (N_15070,N_14923,N_14913);
nand U15071 (N_15071,N_14939,N_14929);
and U15072 (N_15072,N_14834,N_14956);
nor U15073 (N_15073,N_14988,N_14951);
and U15074 (N_15074,N_14924,N_14869);
nor U15075 (N_15075,N_14849,N_14861);
xor U15076 (N_15076,N_14982,N_14936);
nor U15077 (N_15077,N_14862,N_14838);
and U15078 (N_15078,N_14992,N_14974);
nor U15079 (N_15079,N_14920,N_14940);
and U15080 (N_15080,N_14800,N_14832);
and U15081 (N_15081,N_14919,N_14989);
nand U15082 (N_15082,N_14810,N_14826);
nor U15083 (N_15083,N_14844,N_14946);
or U15084 (N_15084,N_14811,N_14980);
or U15085 (N_15085,N_14818,N_14848);
and U15086 (N_15086,N_14912,N_14893);
or U15087 (N_15087,N_14906,N_14814);
or U15088 (N_15088,N_14804,N_14999);
xor U15089 (N_15089,N_14984,N_14969);
nor U15090 (N_15090,N_14932,N_14831);
nand U15091 (N_15091,N_14950,N_14953);
or U15092 (N_15092,N_14805,N_14803);
nor U15093 (N_15093,N_14899,N_14836);
nand U15094 (N_15094,N_14904,N_14846);
or U15095 (N_15095,N_14872,N_14843);
nor U15096 (N_15096,N_14959,N_14878);
nor U15097 (N_15097,N_14991,N_14828);
nand U15098 (N_15098,N_14892,N_14957);
or U15099 (N_15099,N_14830,N_14914);
nand U15100 (N_15100,N_14810,N_14995);
nand U15101 (N_15101,N_14852,N_14822);
xnor U15102 (N_15102,N_14980,N_14955);
and U15103 (N_15103,N_14819,N_14919);
and U15104 (N_15104,N_14857,N_14909);
or U15105 (N_15105,N_14816,N_14866);
nand U15106 (N_15106,N_14836,N_14885);
or U15107 (N_15107,N_14899,N_14943);
nand U15108 (N_15108,N_14948,N_14873);
and U15109 (N_15109,N_14970,N_14847);
nand U15110 (N_15110,N_14883,N_14936);
or U15111 (N_15111,N_14931,N_14969);
nor U15112 (N_15112,N_14869,N_14891);
xor U15113 (N_15113,N_14812,N_14835);
nand U15114 (N_15114,N_14921,N_14920);
nor U15115 (N_15115,N_14837,N_14999);
nor U15116 (N_15116,N_14946,N_14907);
and U15117 (N_15117,N_14938,N_14963);
or U15118 (N_15118,N_14901,N_14975);
xor U15119 (N_15119,N_14826,N_14904);
and U15120 (N_15120,N_14809,N_14914);
or U15121 (N_15121,N_14985,N_14969);
and U15122 (N_15122,N_14864,N_14898);
nand U15123 (N_15123,N_14971,N_14942);
xor U15124 (N_15124,N_14821,N_14982);
xnor U15125 (N_15125,N_14824,N_14804);
xor U15126 (N_15126,N_14855,N_14841);
and U15127 (N_15127,N_14856,N_14841);
nand U15128 (N_15128,N_14873,N_14800);
nor U15129 (N_15129,N_14865,N_14846);
and U15130 (N_15130,N_14935,N_14864);
or U15131 (N_15131,N_14991,N_14913);
or U15132 (N_15132,N_14823,N_14971);
xor U15133 (N_15133,N_14931,N_14976);
or U15134 (N_15134,N_14818,N_14804);
or U15135 (N_15135,N_14994,N_14827);
or U15136 (N_15136,N_14906,N_14946);
nor U15137 (N_15137,N_14893,N_14996);
nor U15138 (N_15138,N_14847,N_14870);
nor U15139 (N_15139,N_14916,N_14836);
and U15140 (N_15140,N_14842,N_14968);
nand U15141 (N_15141,N_14932,N_14956);
nand U15142 (N_15142,N_14808,N_14867);
nand U15143 (N_15143,N_14861,N_14829);
and U15144 (N_15144,N_14982,N_14857);
nor U15145 (N_15145,N_14820,N_14939);
nand U15146 (N_15146,N_14875,N_14860);
nor U15147 (N_15147,N_14887,N_14886);
xor U15148 (N_15148,N_14831,N_14870);
or U15149 (N_15149,N_14949,N_14875);
and U15150 (N_15150,N_14865,N_14858);
nand U15151 (N_15151,N_14999,N_14972);
nor U15152 (N_15152,N_14829,N_14800);
nor U15153 (N_15153,N_14816,N_14941);
xnor U15154 (N_15154,N_14920,N_14827);
nand U15155 (N_15155,N_14899,N_14852);
nand U15156 (N_15156,N_14876,N_14919);
or U15157 (N_15157,N_14993,N_14872);
xor U15158 (N_15158,N_14826,N_14816);
nor U15159 (N_15159,N_14869,N_14973);
or U15160 (N_15160,N_14883,N_14869);
and U15161 (N_15161,N_14805,N_14837);
or U15162 (N_15162,N_14807,N_14906);
and U15163 (N_15163,N_14969,N_14964);
or U15164 (N_15164,N_14837,N_14817);
xor U15165 (N_15165,N_14898,N_14971);
nand U15166 (N_15166,N_14940,N_14903);
or U15167 (N_15167,N_14857,N_14997);
nor U15168 (N_15168,N_14962,N_14912);
xnor U15169 (N_15169,N_14891,N_14837);
and U15170 (N_15170,N_14909,N_14907);
nand U15171 (N_15171,N_14850,N_14913);
xor U15172 (N_15172,N_14899,N_14807);
xnor U15173 (N_15173,N_14929,N_14947);
nor U15174 (N_15174,N_14953,N_14928);
xnor U15175 (N_15175,N_14909,N_14994);
or U15176 (N_15176,N_14993,N_14971);
and U15177 (N_15177,N_14855,N_14907);
nand U15178 (N_15178,N_14900,N_14958);
nor U15179 (N_15179,N_14896,N_14806);
nand U15180 (N_15180,N_14946,N_14905);
and U15181 (N_15181,N_14997,N_14974);
or U15182 (N_15182,N_14905,N_14829);
xor U15183 (N_15183,N_14975,N_14825);
nand U15184 (N_15184,N_14856,N_14995);
or U15185 (N_15185,N_14988,N_14810);
nor U15186 (N_15186,N_14808,N_14920);
nand U15187 (N_15187,N_14991,N_14870);
nor U15188 (N_15188,N_14886,N_14855);
nor U15189 (N_15189,N_14877,N_14926);
nor U15190 (N_15190,N_14969,N_14812);
or U15191 (N_15191,N_14999,N_14818);
or U15192 (N_15192,N_14950,N_14999);
nor U15193 (N_15193,N_14866,N_14920);
or U15194 (N_15194,N_14888,N_14980);
xnor U15195 (N_15195,N_14949,N_14932);
or U15196 (N_15196,N_14803,N_14942);
and U15197 (N_15197,N_14853,N_14992);
and U15198 (N_15198,N_14972,N_14953);
nand U15199 (N_15199,N_14956,N_14909);
nor U15200 (N_15200,N_15059,N_15157);
and U15201 (N_15201,N_15171,N_15077);
nor U15202 (N_15202,N_15195,N_15045);
nor U15203 (N_15203,N_15075,N_15127);
and U15204 (N_15204,N_15181,N_15074);
and U15205 (N_15205,N_15010,N_15011);
and U15206 (N_15206,N_15009,N_15123);
and U15207 (N_15207,N_15156,N_15065);
or U15208 (N_15208,N_15076,N_15064);
nor U15209 (N_15209,N_15160,N_15174);
nand U15210 (N_15210,N_15113,N_15017);
xnor U15211 (N_15211,N_15090,N_15020);
and U15212 (N_15212,N_15040,N_15197);
or U15213 (N_15213,N_15177,N_15120);
and U15214 (N_15214,N_15111,N_15046);
nand U15215 (N_15215,N_15167,N_15005);
nor U15216 (N_15216,N_15097,N_15173);
nor U15217 (N_15217,N_15116,N_15187);
or U15218 (N_15218,N_15152,N_15028);
xor U15219 (N_15219,N_15122,N_15096);
or U15220 (N_15220,N_15133,N_15034);
nor U15221 (N_15221,N_15159,N_15030);
nand U15222 (N_15222,N_15110,N_15108);
xnor U15223 (N_15223,N_15062,N_15142);
nand U15224 (N_15224,N_15119,N_15183);
nor U15225 (N_15225,N_15025,N_15124);
xnor U15226 (N_15226,N_15199,N_15088);
or U15227 (N_15227,N_15188,N_15115);
nor U15228 (N_15228,N_15042,N_15193);
or U15229 (N_15229,N_15155,N_15130);
or U15230 (N_15230,N_15033,N_15175);
nand U15231 (N_15231,N_15112,N_15036);
xor U15232 (N_15232,N_15024,N_15139);
and U15233 (N_15233,N_15098,N_15041);
nor U15234 (N_15234,N_15180,N_15095);
and U15235 (N_15235,N_15068,N_15163);
and U15236 (N_15236,N_15056,N_15050);
nand U15237 (N_15237,N_15189,N_15066);
nand U15238 (N_15238,N_15178,N_15136);
or U15239 (N_15239,N_15054,N_15186);
xnor U15240 (N_15240,N_15162,N_15100);
nand U15241 (N_15241,N_15140,N_15037);
or U15242 (N_15242,N_15007,N_15170);
xnor U15243 (N_15243,N_15104,N_15169);
nand U15244 (N_15244,N_15089,N_15151);
xnor U15245 (N_15245,N_15125,N_15158);
xnor U15246 (N_15246,N_15093,N_15013);
nand U15247 (N_15247,N_15029,N_15079);
nor U15248 (N_15248,N_15053,N_15000);
nor U15249 (N_15249,N_15145,N_15055);
or U15250 (N_15250,N_15144,N_15132);
xnor U15251 (N_15251,N_15149,N_15191);
xnor U15252 (N_15252,N_15080,N_15032);
nor U15253 (N_15253,N_15094,N_15052);
nand U15254 (N_15254,N_15057,N_15015);
or U15255 (N_15255,N_15179,N_15103);
nand U15256 (N_15256,N_15038,N_15154);
or U15257 (N_15257,N_15099,N_15109);
and U15258 (N_15258,N_15018,N_15084);
or U15259 (N_15259,N_15004,N_15190);
nor U15260 (N_15260,N_15150,N_15083);
or U15261 (N_15261,N_15166,N_15168);
nor U15262 (N_15262,N_15129,N_15134);
nor U15263 (N_15263,N_15114,N_15138);
nor U15264 (N_15264,N_15107,N_15001);
nand U15265 (N_15265,N_15184,N_15137);
or U15266 (N_15266,N_15087,N_15182);
nor U15267 (N_15267,N_15078,N_15086);
xnor U15268 (N_15268,N_15101,N_15161);
nor U15269 (N_15269,N_15026,N_15049);
and U15270 (N_15270,N_15121,N_15105);
or U15271 (N_15271,N_15039,N_15006);
xnor U15272 (N_15272,N_15148,N_15131);
nor U15273 (N_15273,N_15063,N_15070);
and U15274 (N_15274,N_15146,N_15023);
nand U15275 (N_15275,N_15196,N_15003);
xor U15276 (N_15276,N_15198,N_15147);
nor U15277 (N_15277,N_15027,N_15126);
and U15278 (N_15278,N_15008,N_15128);
or U15279 (N_15279,N_15021,N_15071);
xor U15280 (N_15280,N_15143,N_15102);
and U15281 (N_15281,N_15069,N_15016);
and U15282 (N_15282,N_15194,N_15092);
nor U15283 (N_15283,N_15073,N_15153);
xor U15284 (N_15284,N_15067,N_15031);
nand U15285 (N_15285,N_15035,N_15118);
nand U15286 (N_15286,N_15082,N_15047);
xor U15287 (N_15287,N_15192,N_15164);
or U15288 (N_15288,N_15044,N_15022);
or U15289 (N_15289,N_15165,N_15106);
nor U15290 (N_15290,N_15014,N_15081);
xor U15291 (N_15291,N_15012,N_15141);
xor U15292 (N_15292,N_15117,N_15002);
xnor U15293 (N_15293,N_15048,N_15051);
nand U15294 (N_15294,N_15061,N_15019);
and U15295 (N_15295,N_15091,N_15058);
and U15296 (N_15296,N_15085,N_15172);
or U15297 (N_15297,N_15135,N_15176);
nor U15298 (N_15298,N_15060,N_15185);
xnor U15299 (N_15299,N_15072,N_15043);
or U15300 (N_15300,N_15080,N_15181);
or U15301 (N_15301,N_15125,N_15188);
and U15302 (N_15302,N_15144,N_15156);
nand U15303 (N_15303,N_15174,N_15102);
nand U15304 (N_15304,N_15008,N_15024);
and U15305 (N_15305,N_15190,N_15115);
xor U15306 (N_15306,N_15111,N_15120);
or U15307 (N_15307,N_15002,N_15141);
xnor U15308 (N_15308,N_15052,N_15073);
nand U15309 (N_15309,N_15048,N_15160);
nor U15310 (N_15310,N_15067,N_15180);
xor U15311 (N_15311,N_15194,N_15144);
xor U15312 (N_15312,N_15151,N_15068);
xnor U15313 (N_15313,N_15117,N_15067);
xnor U15314 (N_15314,N_15148,N_15032);
nor U15315 (N_15315,N_15143,N_15128);
xnor U15316 (N_15316,N_15048,N_15161);
or U15317 (N_15317,N_15052,N_15158);
nand U15318 (N_15318,N_15143,N_15118);
and U15319 (N_15319,N_15156,N_15053);
or U15320 (N_15320,N_15082,N_15050);
and U15321 (N_15321,N_15113,N_15105);
and U15322 (N_15322,N_15138,N_15151);
or U15323 (N_15323,N_15001,N_15035);
and U15324 (N_15324,N_15041,N_15019);
nand U15325 (N_15325,N_15133,N_15007);
nor U15326 (N_15326,N_15148,N_15078);
nand U15327 (N_15327,N_15005,N_15087);
nand U15328 (N_15328,N_15085,N_15012);
xnor U15329 (N_15329,N_15162,N_15156);
xnor U15330 (N_15330,N_15178,N_15155);
xnor U15331 (N_15331,N_15168,N_15109);
nand U15332 (N_15332,N_15015,N_15162);
or U15333 (N_15333,N_15002,N_15120);
nand U15334 (N_15334,N_15056,N_15032);
nor U15335 (N_15335,N_15092,N_15101);
nand U15336 (N_15336,N_15038,N_15135);
nand U15337 (N_15337,N_15027,N_15108);
xor U15338 (N_15338,N_15074,N_15135);
and U15339 (N_15339,N_15111,N_15090);
nor U15340 (N_15340,N_15159,N_15114);
nor U15341 (N_15341,N_15097,N_15185);
xnor U15342 (N_15342,N_15039,N_15147);
nor U15343 (N_15343,N_15124,N_15135);
xor U15344 (N_15344,N_15178,N_15111);
or U15345 (N_15345,N_15066,N_15040);
nand U15346 (N_15346,N_15128,N_15176);
nor U15347 (N_15347,N_15002,N_15130);
nand U15348 (N_15348,N_15121,N_15051);
nand U15349 (N_15349,N_15007,N_15141);
or U15350 (N_15350,N_15060,N_15178);
or U15351 (N_15351,N_15189,N_15179);
nand U15352 (N_15352,N_15129,N_15010);
xor U15353 (N_15353,N_15009,N_15149);
nand U15354 (N_15354,N_15132,N_15122);
nor U15355 (N_15355,N_15158,N_15196);
nor U15356 (N_15356,N_15004,N_15106);
xnor U15357 (N_15357,N_15171,N_15181);
nor U15358 (N_15358,N_15199,N_15081);
and U15359 (N_15359,N_15112,N_15015);
and U15360 (N_15360,N_15139,N_15159);
nor U15361 (N_15361,N_15037,N_15170);
or U15362 (N_15362,N_15132,N_15063);
nand U15363 (N_15363,N_15197,N_15110);
or U15364 (N_15364,N_15099,N_15171);
or U15365 (N_15365,N_15198,N_15001);
and U15366 (N_15366,N_15121,N_15094);
xor U15367 (N_15367,N_15075,N_15065);
xor U15368 (N_15368,N_15029,N_15123);
and U15369 (N_15369,N_15059,N_15020);
xor U15370 (N_15370,N_15099,N_15076);
nand U15371 (N_15371,N_15162,N_15069);
and U15372 (N_15372,N_15038,N_15176);
or U15373 (N_15373,N_15121,N_15049);
xor U15374 (N_15374,N_15091,N_15117);
xnor U15375 (N_15375,N_15100,N_15191);
nor U15376 (N_15376,N_15138,N_15046);
or U15377 (N_15377,N_15191,N_15032);
nor U15378 (N_15378,N_15122,N_15045);
and U15379 (N_15379,N_15097,N_15060);
nand U15380 (N_15380,N_15195,N_15011);
xnor U15381 (N_15381,N_15107,N_15094);
or U15382 (N_15382,N_15181,N_15090);
xnor U15383 (N_15383,N_15120,N_15113);
and U15384 (N_15384,N_15191,N_15105);
or U15385 (N_15385,N_15174,N_15014);
nor U15386 (N_15386,N_15149,N_15060);
and U15387 (N_15387,N_15014,N_15186);
nand U15388 (N_15388,N_15077,N_15124);
nor U15389 (N_15389,N_15119,N_15030);
or U15390 (N_15390,N_15105,N_15084);
nor U15391 (N_15391,N_15170,N_15146);
nor U15392 (N_15392,N_15184,N_15177);
or U15393 (N_15393,N_15002,N_15041);
and U15394 (N_15394,N_15095,N_15133);
xnor U15395 (N_15395,N_15111,N_15142);
or U15396 (N_15396,N_15109,N_15136);
nor U15397 (N_15397,N_15093,N_15122);
and U15398 (N_15398,N_15079,N_15162);
or U15399 (N_15399,N_15173,N_15053);
nor U15400 (N_15400,N_15349,N_15217);
nand U15401 (N_15401,N_15203,N_15306);
nor U15402 (N_15402,N_15251,N_15343);
or U15403 (N_15403,N_15348,N_15366);
or U15404 (N_15404,N_15278,N_15252);
nor U15405 (N_15405,N_15248,N_15223);
xor U15406 (N_15406,N_15299,N_15293);
xnor U15407 (N_15407,N_15326,N_15398);
and U15408 (N_15408,N_15334,N_15201);
and U15409 (N_15409,N_15250,N_15368);
nand U15410 (N_15410,N_15328,N_15303);
xor U15411 (N_15411,N_15387,N_15282);
nor U15412 (N_15412,N_15382,N_15233);
nand U15413 (N_15413,N_15311,N_15381);
nor U15414 (N_15414,N_15283,N_15200);
nor U15415 (N_15415,N_15389,N_15263);
or U15416 (N_15416,N_15377,N_15327);
xnor U15417 (N_15417,N_15209,N_15245);
xor U15418 (N_15418,N_15253,N_15374);
xor U15419 (N_15419,N_15359,N_15222);
and U15420 (N_15420,N_15344,N_15386);
xnor U15421 (N_15421,N_15331,N_15224);
or U15422 (N_15422,N_15287,N_15315);
nand U15423 (N_15423,N_15260,N_15211);
or U15424 (N_15424,N_15259,N_15296);
and U15425 (N_15425,N_15330,N_15391);
and U15426 (N_15426,N_15212,N_15290);
and U15427 (N_15427,N_15305,N_15355);
nor U15428 (N_15428,N_15205,N_15225);
nand U15429 (N_15429,N_15304,N_15323);
xor U15430 (N_15430,N_15345,N_15370);
nand U15431 (N_15431,N_15347,N_15365);
nand U15432 (N_15432,N_15332,N_15291);
and U15433 (N_15433,N_15244,N_15228);
and U15434 (N_15434,N_15238,N_15231);
nor U15435 (N_15435,N_15310,N_15254);
xor U15436 (N_15436,N_15322,N_15346);
or U15437 (N_15437,N_15277,N_15392);
xor U15438 (N_15438,N_15294,N_15236);
xor U15439 (N_15439,N_15383,N_15394);
nor U15440 (N_15440,N_15246,N_15362);
or U15441 (N_15441,N_15393,N_15369);
or U15442 (N_15442,N_15308,N_15397);
or U15443 (N_15443,N_15337,N_15339);
xnor U15444 (N_15444,N_15247,N_15358);
and U15445 (N_15445,N_15227,N_15329);
xnor U15446 (N_15446,N_15206,N_15342);
xnor U15447 (N_15447,N_15367,N_15276);
or U15448 (N_15448,N_15354,N_15265);
and U15449 (N_15449,N_15333,N_15312);
and U15450 (N_15450,N_15388,N_15364);
nand U15451 (N_15451,N_15219,N_15271);
nand U15452 (N_15452,N_15241,N_15218);
or U15453 (N_15453,N_15202,N_15385);
and U15454 (N_15454,N_15360,N_15268);
nor U15455 (N_15455,N_15261,N_15313);
xnor U15456 (N_15456,N_15340,N_15270);
and U15457 (N_15457,N_15372,N_15280);
xor U15458 (N_15458,N_15318,N_15262);
nor U15459 (N_15459,N_15338,N_15350);
nor U15460 (N_15460,N_15237,N_15256);
nor U15461 (N_15461,N_15279,N_15357);
or U15462 (N_15462,N_15267,N_15274);
nand U15463 (N_15463,N_15320,N_15235);
and U15464 (N_15464,N_15275,N_15284);
xor U15465 (N_15465,N_15361,N_15242);
xor U15466 (N_15466,N_15309,N_15243);
nor U15467 (N_15467,N_15214,N_15379);
nor U15468 (N_15468,N_15371,N_15335);
and U15469 (N_15469,N_15395,N_15324);
nor U15470 (N_15470,N_15351,N_15399);
xor U15471 (N_15471,N_15302,N_15356);
nor U15472 (N_15472,N_15234,N_15316);
xor U15473 (N_15473,N_15336,N_15226);
or U15474 (N_15474,N_15239,N_15380);
nor U15475 (N_15475,N_15301,N_15289);
and U15476 (N_15476,N_15321,N_15300);
nor U15477 (N_15477,N_15230,N_15297);
nor U15478 (N_15478,N_15375,N_15376);
nand U15479 (N_15479,N_15295,N_15373);
or U15480 (N_15480,N_15363,N_15269);
or U15481 (N_15481,N_15288,N_15314);
or U15482 (N_15482,N_15286,N_15255);
and U15483 (N_15483,N_15264,N_15232);
nor U15484 (N_15484,N_15221,N_15258);
or U15485 (N_15485,N_15249,N_15298);
and U15486 (N_15486,N_15378,N_15207);
xnor U15487 (N_15487,N_15292,N_15240);
and U15488 (N_15488,N_15220,N_15319);
xor U15489 (N_15489,N_15384,N_15266);
nor U15490 (N_15490,N_15281,N_15215);
nand U15491 (N_15491,N_15216,N_15353);
nor U15492 (N_15492,N_15272,N_15341);
nand U15493 (N_15493,N_15204,N_15210);
or U15494 (N_15494,N_15307,N_15396);
xor U15495 (N_15495,N_15208,N_15285);
nor U15496 (N_15496,N_15325,N_15273);
nor U15497 (N_15497,N_15317,N_15390);
nand U15498 (N_15498,N_15213,N_15229);
nor U15499 (N_15499,N_15352,N_15257);
nor U15500 (N_15500,N_15393,N_15349);
or U15501 (N_15501,N_15354,N_15238);
or U15502 (N_15502,N_15250,N_15346);
xor U15503 (N_15503,N_15289,N_15382);
and U15504 (N_15504,N_15280,N_15264);
nor U15505 (N_15505,N_15278,N_15395);
nor U15506 (N_15506,N_15335,N_15338);
xor U15507 (N_15507,N_15232,N_15200);
nor U15508 (N_15508,N_15218,N_15214);
and U15509 (N_15509,N_15363,N_15310);
nand U15510 (N_15510,N_15297,N_15379);
and U15511 (N_15511,N_15296,N_15382);
and U15512 (N_15512,N_15283,N_15207);
or U15513 (N_15513,N_15229,N_15264);
nor U15514 (N_15514,N_15360,N_15359);
nand U15515 (N_15515,N_15262,N_15225);
or U15516 (N_15516,N_15247,N_15327);
xor U15517 (N_15517,N_15227,N_15229);
nand U15518 (N_15518,N_15216,N_15343);
nand U15519 (N_15519,N_15268,N_15260);
nand U15520 (N_15520,N_15231,N_15269);
or U15521 (N_15521,N_15397,N_15372);
nand U15522 (N_15522,N_15257,N_15225);
or U15523 (N_15523,N_15336,N_15218);
and U15524 (N_15524,N_15360,N_15213);
or U15525 (N_15525,N_15287,N_15341);
nand U15526 (N_15526,N_15218,N_15332);
or U15527 (N_15527,N_15342,N_15351);
nand U15528 (N_15528,N_15390,N_15351);
nand U15529 (N_15529,N_15368,N_15383);
or U15530 (N_15530,N_15363,N_15352);
nor U15531 (N_15531,N_15353,N_15375);
nor U15532 (N_15532,N_15358,N_15309);
or U15533 (N_15533,N_15236,N_15282);
and U15534 (N_15534,N_15297,N_15366);
and U15535 (N_15535,N_15323,N_15233);
xor U15536 (N_15536,N_15230,N_15396);
nor U15537 (N_15537,N_15360,N_15271);
or U15538 (N_15538,N_15224,N_15237);
nor U15539 (N_15539,N_15372,N_15282);
xor U15540 (N_15540,N_15350,N_15302);
or U15541 (N_15541,N_15332,N_15313);
xnor U15542 (N_15542,N_15358,N_15392);
nor U15543 (N_15543,N_15225,N_15387);
xnor U15544 (N_15544,N_15381,N_15276);
nor U15545 (N_15545,N_15239,N_15221);
or U15546 (N_15546,N_15365,N_15245);
or U15547 (N_15547,N_15220,N_15377);
nor U15548 (N_15548,N_15310,N_15265);
xor U15549 (N_15549,N_15301,N_15317);
and U15550 (N_15550,N_15208,N_15378);
nand U15551 (N_15551,N_15296,N_15354);
nor U15552 (N_15552,N_15357,N_15205);
and U15553 (N_15553,N_15228,N_15226);
xnor U15554 (N_15554,N_15361,N_15357);
nor U15555 (N_15555,N_15263,N_15236);
nor U15556 (N_15556,N_15389,N_15381);
and U15557 (N_15557,N_15332,N_15229);
nor U15558 (N_15558,N_15324,N_15274);
nand U15559 (N_15559,N_15240,N_15276);
nand U15560 (N_15560,N_15388,N_15217);
or U15561 (N_15561,N_15365,N_15392);
and U15562 (N_15562,N_15206,N_15392);
and U15563 (N_15563,N_15388,N_15332);
nand U15564 (N_15564,N_15218,N_15328);
xor U15565 (N_15565,N_15301,N_15351);
or U15566 (N_15566,N_15244,N_15339);
and U15567 (N_15567,N_15227,N_15206);
nor U15568 (N_15568,N_15297,N_15286);
and U15569 (N_15569,N_15242,N_15282);
nor U15570 (N_15570,N_15307,N_15301);
or U15571 (N_15571,N_15265,N_15220);
and U15572 (N_15572,N_15278,N_15352);
nand U15573 (N_15573,N_15237,N_15258);
xor U15574 (N_15574,N_15398,N_15243);
or U15575 (N_15575,N_15267,N_15269);
and U15576 (N_15576,N_15342,N_15270);
nor U15577 (N_15577,N_15316,N_15345);
and U15578 (N_15578,N_15289,N_15322);
xor U15579 (N_15579,N_15282,N_15366);
and U15580 (N_15580,N_15299,N_15214);
xnor U15581 (N_15581,N_15260,N_15205);
and U15582 (N_15582,N_15357,N_15319);
nand U15583 (N_15583,N_15204,N_15329);
xnor U15584 (N_15584,N_15268,N_15375);
and U15585 (N_15585,N_15251,N_15340);
xor U15586 (N_15586,N_15389,N_15219);
nand U15587 (N_15587,N_15360,N_15334);
nor U15588 (N_15588,N_15323,N_15314);
xnor U15589 (N_15589,N_15388,N_15207);
and U15590 (N_15590,N_15226,N_15345);
and U15591 (N_15591,N_15238,N_15213);
or U15592 (N_15592,N_15206,N_15268);
and U15593 (N_15593,N_15307,N_15350);
and U15594 (N_15594,N_15312,N_15300);
and U15595 (N_15595,N_15249,N_15238);
and U15596 (N_15596,N_15290,N_15359);
nand U15597 (N_15597,N_15389,N_15270);
xnor U15598 (N_15598,N_15200,N_15204);
xnor U15599 (N_15599,N_15237,N_15204);
and U15600 (N_15600,N_15415,N_15541);
nor U15601 (N_15601,N_15430,N_15432);
xor U15602 (N_15602,N_15450,N_15413);
nor U15603 (N_15603,N_15510,N_15427);
nor U15604 (N_15604,N_15491,N_15436);
nand U15605 (N_15605,N_15406,N_15424);
nand U15606 (N_15606,N_15443,N_15565);
nand U15607 (N_15607,N_15405,N_15417);
nand U15608 (N_15608,N_15463,N_15429);
nor U15609 (N_15609,N_15512,N_15576);
nand U15610 (N_15610,N_15515,N_15409);
nand U15611 (N_15611,N_15469,N_15435);
nor U15612 (N_15612,N_15455,N_15407);
xnor U15613 (N_15613,N_15559,N_15412);
and U15614 (N_15614,N_15503,N_15571);
xor U15615 (N_15615,N_15434,N_15552);
xnor U15616 (N_15616,N_15585,N_15421);
and U15617 (N_15617,N_15489,N_15550);
xnor U15618 (N_15618,N_15534,N_15403);
or U15619 (N_15619,N_15582,N_15459);
nor U15620 (N_15620,N_15579,N_15560);
and U15621 (N_15621,N_15589,N_15465);
xor U15622 (N_15622,N_15451,N_15522);
nor U15623 (N_15623,N_15468,N_15461);
nand U15624 (N_15624,N_15423,N_15454);
xor U15625 (N_15625,N_15476,N_15470);
nand U15626 (N_15626,N_15493,N_15481);
nor U15627 (N_15627,N_15447,N_15437);
and U15628 (N_15628,N_15477,N_15547);
nor U15629 (N_15629,N_15537,N_15453);
and U15630 (N_15630,N_15572,N_15482);
nor U15631 (N_15631,N_15528,N_15478);
and U15632 (N_15632,N_15519,N_15597);
nor U15633 (N_15633,N_15414,N_15595);
nor U15634 (N_15634,N_15456,N_15555);
or U15635 (N_15635,N_15480,N_15543);
nand U15636 (N_15636,N_15533,N_15591);
and U15637 (N_15637,N_15535,N_15483);
and U15638 (N_15638,N_15484,N_15462);
nor U15639 (N_15639,N_15587,N_15580);
or U15640 (N_15640,N_15410,N_15488);
xnor U15641 (N_15641,N_15594,N_15408);
or U15642 (N_15642,N_15556,N_15509);
xnor U15643 (N_15643,N_15506,N_15425);
xnor U15644 (N_15644,N_15561,N_15592);
nor U15645 (N_15645,N_15577,N_15438);
nor U15646 (N_15646,N_15420,N_15497);
nand U15647 (N_15647,N_15418,N_15567);
xor U15648 (N_15648,N_15449,N_15524);
nor U15649 (N_15649,N_15558,N_15445);
and U15650 (N_15650,N_15460,N_15440);
or U15651 (N_15651,N_15507,N_15471);
nor U15652 (N_15652,N_15578,N_15596);
nor U15653 (N_15653,N_15568,N_15544);
and U15654 (N_15654,N_15426,N_15411);
nor U15655 (N_15655,N_15563,N_15516);
nor U15656 (N_15656,N_15439,N_15566);
xnor U15657 (N_15657,N_15538,N_15526);
xor U15658 (N_15658,N_15400,N_15573);
xor U15659 (N_15659,N_15564,N_15498);
or U15660 (N_15660,N_15574,N_15401);
or U15661 (N_15661,N_15402,N_15475);
nor U15662 (N_15662,N_15513,N_15499);
or U15663 (N_15663,N_15508,N_15546);
nand U15664 (N_15664,N_15530,N_15518);
or U15665 (N_15665,N_15495,N_15540);
nand U15666 (N_15666,N_15487,N_15464);
nand U15667 (N_15667,N_15557,N_15473);
xnor U15668 (N_15668,N_15444,N_15520);
xor U15669 (N_15669,N_15404,N_15457);
and U15670 (N_15670,N_15441,N_15569);
xnor U15671 (N_15671,N_15586,N_15501);
nor U15672 (N_15672,N_15446,N_15433);
nand U15673 (N_15673,N_15428,N_15479);
xnor U15674 (N_15674,N_15583,N_15486);
and U15675 (N_15675,N_15554,N_15474);
xor U15676 (N_15676,N_15458,N_15545);
nand U15677 (N_15677,N_15514,N_15532);
nand U15678 (N_15678,N_15505,N_15523);
xnor U15679 (N_15679,N_15504,N_15431);
or U15680 (N_15680,N_15599,N_15551);
nand U15681 (N_15681,N_15419,N_15452);
or U15682 (N_15682,N_15472,N_15466);
nand U15683 (N_15683,N_15562,N_15485);
or U15684 (N_15684,N_15575,N_15529);
xor U15685 (N_15685,N_15590,N_15598);
nand U15686 (N_15686,N_15517,N_15525);
nor U15687 (N_15687,N_15536,N_15539);
or U15688 (N_15688,N_15422,N_15496);
xor U15689 (N_15689,N_15494,N_15581);
or U15690 (N_15690,N_15588,N_15502);
or U15691 (N_15691,N_15570,N_15527);
and U15692 (N_15692,N_15548,N_15467);
xor U15693 (N_15693,N_15542,N_15448);
or U15694 (N_15694,N_15500,N_15553);
xnor U15695 (N_15695,N_15531,N_15442);
nand U15696 (N_15696,N_15549,N_15511);
nor U15697 (N_15697,N_15492,N_15521);
xor U15698 (N_15698,N_15593,N_15584);
nand U15699 (N_15699,N_15416,N_15490);
nand U15700 (N_15700,N_15527,N_15493);
nand U15701 (N_15701,N_15473,N_15460);
or U15702 (N_15702,N_15463,N_15522);
nand U15703 (N_15703,N_15431,N_15418);
xor U15704 (N_15704,N_15444,N_15599);
xor U15705 (N_15705,N_15583,N_15484);
nand U15706 (N_15706,N_15471,N_15527);
xor U15707 (N_15707,N_15584,N_15581);
or U15708 (N_15708,N_15549,N_15546);
xor U15709 (N_15709,N_15419,N_15400);
nor U15710 (N_15710,N_15550,N_15428);
or U15711 (N_15711,N_15527,N_15512);
and U15712 (N_15712,N_15442,N_15418);
xnor U15713 (N_15713,N_15411,N_15416);
and U15714 (N_15714,N_15422,N_15541);
xnor U15715 (N_15715,N_15583,N_15561);
xor U15716 (N_15716,N_15509,N_15435);
xor U15717 (N_15717,N_15553,N_15519);
or U15718 (N_15718,N_15586,N_15542);
nand U15719 (N_15719,N_15550,N_15461);
xnor U15720 (N_15720,N_15454,N_15592);
nor U15721 (N_15721,N_15424,N_15457);
xor U15722 (N_15722,N_15438,N_15572);
nand U15723 (N_15723,N_15478,N_15537);
or U15724 (N_15724,N_15523,N_15470);
nand U15725 (N_15725,N_15583,N_15557);
nor U15726 (N_15726,N_15538,N_15428);
nand U15727 (N_15727,N_15451,N_15550);
or U15728 (N_15728,N_15510,N_15544);
nand U15729 (N_15729,N_15432,N_15519);
xnor U15730 (N_15730,N_15408,N_15452);
xor U15731 (N_15731,N_15502,N_15515);
nand U15732 (N_15732,N_15479,N_15582);
and U15733 (N_15733,N_15522,N_15466);
xor U15734 (N_15734,N_15423,N_15597);
xnor U15735 (N_15735,N_15487,N_15418);
xnor U15736 (N_15736,N_15454,N_15467);
nand U15737 (N_15737,N_15418,N_15561);
and U15738 (N_15738,N_15513,N_15434);
or U15739 (N_15739,N_15500,N_15564);
nand U15740 (N_15740,N_15408,N_15553);
nor U15741 (N_15741,N_15551,N_15550);
nand U15742 (N_15742,N_15458,N_15544);
xor U15743 (N_15743,N_15484,N_15430);
or U15744 (N_15744,N_15496,N_15564);
xor U15745 (N_15745,N_15563,N_15423);
nand U15746 (N_15746,N_15468,N_15534);
and U15747 (N_15747,N_15452,N_15481);
nand U15748 (N_15748,N_15482,N_15486);
nor U15749 (N_15749,N_15485,N_15452);
nor U15750 (N_15750,N_15440,N_15498);
xnor U15751 (N_15751,N_15407,N_15417);
or U15752 (N_15752,N_15541,N_15567);
nand U15753 (N_15753,N_15483,N_15547);
and U15754 (N_15754,N_15539,N_15583);
or U15755 (N_15755,N_15482,N_15513);
xnor U15756 (N_15756,N_15541,N_15593);
xor U15757 (N_15757,N_15404,N_15531);
nor U15758 (N_15758,N_15527,N_15571);
nor U15759 (N_15759,N_15527,N_15542);
xnor U15760 (N_15760,N_15438,N_15524);
nor U15761 (N_15761,N_15431,N_15559);
nand U15762 (N_15762,N_15527,N_15452);
or U15763 (N_15763,N_15484,N_15569);
xnor U15764 (N_15764,N_15577,N_15403);
nor U15765 (N_15765,N_15521,N_15596);
nor U15766 (N_15766,N_15446,N_15484);
nand U15767 (N_15767,N_15596,N_15558);
nor U15768 (N_15768,N_15571,N_15597);
xor U15769 (N_15769,N_15468,N_15553);
nor U15770 (N_15770,N_15564,N_15597);
or U15771 (N_15771,N_15464,N_15599);
and U15772 (N_15772,N_15463,N_15505);
and U15773 (N_15773,N_15423,N_15428);
xnor U15774 (N_15774,N_15564,N_15490);
nand U15775 (N_15775,N_15494,N_15433);
or U15776 (N_15776,N_15528,N_15408);
nand U15777 (N_15777,N_15417,N_15422);
xor U15778 (N_15778,N_15403,N_15517);
xnor U15779 (N_15779,N_15599,N_15461);
or U15780 (N_15780,N_15494,N_15404);
or U15781 (N_15781,N_15477,N_15411);
nor U15782 (N_15782,N_15425,N_15461);
xnor U15783 (N_15783,N_15479,N_15471);
and U15784 (N_15784,N_15441,N_15496);
nand U15785 (N_15785,N_15581,N_15403);
xor U15786 (N_15786,N_15544,N_15488);
and U15787 (N_15787,N_15446,N_15599);
xor U15788 (N_15788,N_15537,N_15548);
nand U15789 (N_15789,N_15511,N_15539);
nand U15790 (N_15790,N_15472,N_15570);
xnor U15791 (N_15791,N_15506,N_15593);
or U15792 (N_15792,N_15579,N_15546);
and U15793 (N_15793,N_15585,N_15450);
or U15794 (N_15794,N_15516,N_15476);
nand U15795 (N_15795,N_15483,N_15599);
nand U15796 (N_15796,N_15505,N_15575);
or U15797 (N_15797,N_15497,N_15426);
and U15798 (N_15798,N_15564,N_15581);
nand U15799 (N_15799,N_15557,N_15543);
xor U15800 (N_15800,N_15700,N_15637);
xnor U15801 (N_15801,N_15606,N_15770);
or U15802 (N_15802,N_15603,N_15717);
and U15803 (N_15803,N_15741,N_15605);
nor U15804 (N_15804,N_15651,N_15638);
nor U15805 (N_15805,N_15654,N_15691);
and U15806 (N_15806,N_15608,N_15615);
and U15807 (N_15807,N_15668,N_15627);
xor U15808 (N_15808,N_15708,N_15645);
nand U15809 (N_15809,N_15626,N_15713);
or U15810 (N_15810,N_15686,N_15611);
nand U15811 (N_15811,N_15723,N_15765);
nor U15812 (N_15812,N_15702,N_15728);
xnor U15813 (N_15813,N_15612,N_15624);
xor U15814 (N_15814,N_15640,N_15704);
nor U15815 (N_15815,N_15720,N_15772);
xnor U15816 (N_15816,N_15773,N_15791);
or U15817 (N_15817,N_15672,N_15657);
xnor U15818 (N_15818,N_15744,N_15776);
xor U15819 (N_15819,N_15629,N_15737);
and U15820 (N_15820,N_15639,N_15683);
nand U15821 (N_15821,N_15752,N_15707);
nor U15822 (N_15822,N_15601,N_15695);
or U15823 (N_15823,N_15790,N_15738);
nand U15824 (N_15824,N_15729,N_15732);
and U15825 (N_15825,N_15623,N_15722);
or U15826 (N_15826,N_15602,N_15649);
xnor U15827 (N_15827,N_15782,N_15775);
xnor U15828 (N_15828,N_15662,N_15671);
xor U15829 (N_15829,N_15721,N_15784);
or U15830 (N_15830,N_15618,N_15785);
nand U15831 (N_15831,N_15745,N_15698);
nand U15832 (N_15832,N_15788,N_15619);
or U15833 (N_15833,N_15792,N_15616);
and U15834 (N_15834,N_15669,N_15685);
and U15835 (N_15835,N_15769,N_15631);
and U15836 (N_15836,N_15724,N_15680);
xor U15837 (N_15837,N_15706,N_15794);
and U15838 (N_15838,N_15742,N_15628);
and U15839 (N_15839,N_15653,N_15674);
nor U15840 (N_15840,N_15793,N_15763);
xor U15841 (N_15841,N_15675,N_15757);
nor U15842 (N_15842,N_15771,N_15799);
or U15843 (N_15843,N_15610,N_15740);
xor U15844 (N_15844,N_15607,N_15625);
xor U15845 (N_15845,N_15762,N_15652);
xor U15846 (N_15846,N_15719,N_15664);
xnor U15847 (N_15847,N_15622,N_15697);
nor U15848 (N_15848,N_15656,N_15716);
and U15849 (N_15849,N_15635,N_15600);
or U15850 (N_15850,N_15710,N_15750);
nand U15851 (N_15851,N_15679,N_15659);
and U15852 (N_15852,N_15712,N_15767);
xor U15853 (N_15853,N_15617,N_15797);
and U15854 (N_15854,N_15758,N_15759);
nand U15855 (N_15855,N_15658,N_15768);
nand U15856 (N_15856,N_15783,N_15725);
and U15857 (N_15857,N_15687,N_15764);
xnor U15858 (N_15858,N_15621,N_15777);
and U15859 (N_15859,N_15667,N_15614);
and U15860 (N_15860,N_15647,N_15693);
xor U15861 (N_15861,N_15703,N_15778);
or U15862 (N_15862,N_15754,N_15761);
and U15863 (N_15863,N_15735,N_15796);
and U15864 (N_15864,N_15604,N_15774);
nand U15865 (N_15865,N_15753,N_15746);
nor U15866 (N_15866,N_15696,N_15779);
xnor U15867 (N_15867,N_15690,N_15756);
nor U15868 (N_15868,N_15634,N_15726);
and U15869 (N_15869,N_15666,N_15692);
and U15870 (N_15870,N_15641,N_15682);
nor U15871 (N_15871,N_15665,N_15689);
nor U15872 (N_15872,N_15630,N_15648);
or U15873 (N_15873,N_15646,N_15655);
and U15874 (N_15874,N_15676,N_15644);
nand U15875 (N_15875,N_15787,N_15633);
nand U15876 (N_15876,N_15673,N_15727);
or U15877 (N_15877,N_15620,N_15705);
nand U15878 (N_15878,N_15798,N_15609);
nand U15879 (N_15879,N_15694,N_15789);
or U15880 (N_15880,N_15715,N_15748);
xor U15881 (N_15881,N_15677,N_15751);
nand U15882 (N_15882,N_15660,N_15670);
xnor U15883 (N_15883,N_15642,N_15636);
and U15884 (N_15884,N_15739,N_15699);
and U15885 (N_15885,N_15688,N_15781);
or U15886 (N_15886,N_15733,N_15743);
nand U15887 (N_15887,N_15795,N_15663);
and U15888 (N_15888,N_15632,N_15734);
xnor U15889 (N_15889,N_15678,N_15711);
and U15890 (N_15890,N_15643,N_15650);
nor U15891 (N_15891,N_15760,N_15730);
xor U15892 (N_15892,N_15786,N_15736);
xnor U15893 (N_15893,N_15701,N_15747);
nor U15894 (N_15894,N_15718,N_15661);
nor U15895 (N_15895,N_15684,N_15681);
xnor U15896 (N_15896,N_15709,N_15613);
nor U15897 (N_15897,N_15766,N_15714);
xor U15898 (N_15898,N_15780,N_15731);
xor U15899 (N_15899,N_15749,N_15755);
xnor U15900 (N_15900,N_15654,N_15604);
or U15901 (N_15901,N_15757,N_15667);
nand U15902 (N_15902,N_15786,N_15685);
nor U15903 (N_15903,N_15780,N_15673);
nor U15904 (N_15904,N_15798,N_15764);
and U15905 (N_15905,N_15698,N_15794);
or U15906 (N_15906,N_15730,N_15631);
and U15907 (N_15907,N_15713,N_15714);
nand U15908 (N_15908,N_15717,N_15716);
and U15909 (N_15909,N_15738,N_15662);
nor U15910 (N_15910,N_15685,N_15721);
xor U15911 (N_15911,N_15743,N_15649);
and U15912 (N_15912,N_15670,N_15735);
or U15913 (N_15913,N_15763,N_15707);
nor U15914 (N_15914,N_15756,N_15626);
or U15915 (N_15915,N_15732,N_15682);
or U15916 (N_15916,N_15675,N_15601);
nor U15917 (N_15917,N_15647,N_15730);
xnor U15918 (N_15918,N_15673,N_15627);
nor U15919 (N_15919,N_15754,N_15748);
xnor U15920 (N_15920,N_15799,N_15637);
or U15921 (N_15921,N_15758,N_15636);
and U15922 (N_15922,N_15616,N_15606);
nand U15923 (N_15923,N_15692,N_15634);
xnor U15924 (N_15924,N_15619,N_15679);
nor U15925 (N_15925,N_15651,N_15672);
nor U15926 (N_15926,N_15783,N_15608);
or U15927 (N_15927,N_15627,N_15762);
and U15928 (N_15928,N_15779,N_15796);
nand U15929 (N_15929,N_15615,N_15635);
or U15930 (N_15930,N_15621,N_15628);
nand U15931 (N_15931,N_15616,N_15644);
xor U15932 (N_15932,N_15662,N_15620);
nor U15933 (N_15933,N_15743,N_15762);
nand U15934 (N_15934,N_15615,N_15676);
xor U15935 (N_15935,N_15792,N_15711);
xnor U15936 (N_15936,N_15607,N_15660);
or U15937 (N_15937,N_15659,N_15701);
nand U15938 (N_15938,N_15699,N_15775);
nand U15939 (N_15939,N_15736,N_15632);
and U15940 (N_15940,N_15729,N_15723);
nor U15941 (N_15941,N_15644,N_15745);
nor U15942 (N_15942,N_15696,N_15739);
and U15943 (N_15943,N_15739,N_15652);
nand U15944 (N_15944,N_15735,N_15667);
nand U15945 (N_15945,N_15707,N_15747);
nand U15946 (N_15946,N_15799,N_15626);
and U15947 (N_15947,N_15626,N_15613);
or U15948 (N_15948,N_15711,N_15670);
and U15949 (N_15949,N_15643,N_15698);
xnor U15950 (N_15950,N_15614,N_15697);
or U15951 (N_15951,N_15757,N_15795);
xnor U15952 (N_15952,N_15707,N_15673);
nor U15953 (N_15953,N_15693,N_15789);
nor U15954 (N_15954,N_15652,N_15728);
nand U15955 (N_15955,N_15736,N_15691);
xnor U15956 (N_15956,N_15797,N_15618);
nand U15957 (N_15957,N_15755,N_15660);
xnor U15958 (N_15958,N_15735,N_15663);
xnor U15959 (N_15959,N_15712,N_15781);
or U15960 (N_15960,N_15792,N_15699);
and U15961 (N_15961,N_15642,N_15653);
xor U15962 (N_15962,N_15626,N_15761);
nor U15963 (N_15963,N_15730,N_15652);
or U15964 (N_15964,N_15635,N_15704);
nand U15965 (N_15965,N_15753,N_15693);
and U15966 (N_15966,N_15730,N_15656);
nor U15967 (N_15967,N_15629,N_15751);
and U15968 (N_15968,N_15686,N_15628);
or U15969 (N_15969,N_15613,N_15739);
or U15970 (N_15970,N_15604,N_15686);
and U15971 (N_15971,N_15767,N_15689);
nor U15972 (N_15972,N_15707,N_15648);
nand U15973 (N_15973,N_15799,N_15727);
xnor U15974 (N_15974,N_15799,N_15710);
nor U15975 (N_15975,N_15728,N_15677);
nor U15976 (N_15976,N_15724,N_15688);
nor U15977 (N_15977,N_15608,N_15654);
nor U15978 (N_15978,N_15699,N_15648);
and U15979 (N_15979,N_15682,N_15769);
nand U15980 (N_15980,N_15775,N_15760);
nor U15981 (N_15981,N_15774,N_15707);
and U15982 (N_15982,N_15698,N_15663);
and U15983 (N_15983,N_15737,N_15701);
and U15984 (N_15984,N_15684,N_15683);
and U15985 (N_15985,N_15645,N_15661);
nand U15986 (N_15986,N_15757,N_15673);
or U15987 (N_15987,N_15703,N_15735);
xor U15988 (N_15988,N_15715,N_15672);
and U15989 (N_15989,N_15726,N_15608);
nor U15990 (N_15990,N_15700,N_15776);
or U15991 (N_15991,N_15689,N_15703);
nor U15992 (N_15992,N_15713,N_15669);
and U15993 (N_15993,N_15755,N_15721);
nand U15994 (N_15994,N_15641,N_15731);
xnor U15995 (N_15995,N_15627,N_15790);
nor U15996 (N_15996,N_15752,N_15788);
or U15997 (N_15997,N_15663,N_15688);
nor U15998 (N_15998,N_15608,N_15736);
and U15999 (N_15999,N_15699,N_15777);
nand U16000 (N_16000,N_15826,N_15956);
or U16001 (N_16001,N_15886,N_15811);
nor U16002 (N_16002,N_15829,N_15902);
xor U16003 (N_16003,N_15821,N_15859);
and U16004 (N_16004,N_15999,N_15893);
and U16005 (N_16005,N_15994,N_15898);
or U16006 (N_16006,N_15962,N_15970);
nand U16007 (N_16007,N_15949,N_15824);
xor U16008 (N_16008,N_15885,N_15895);
nand U16009 (N_16009,N_15883,N_15959);
nand U16010 (N_16010,N_15965,N_15920);
nor U16011 (N_16011,N_15825,N_15888);
nand U16012 (N_16012,N_15917,N_15990);
nor U16013 (N_16013,N_15918,N_15843);
or U16014 (N_16014,N_15980,N_15948);
and U16015 (N_16015,N_15838,N_15813);
and U16016 (N_16016,N_15926,N_15889);
and U16017 (N_16017,N_15985,N_15951);
nand U16018 (N_16018,N_15946,N_15900);
and U16019 (N_16019,N_15870,N_15992);
and U16020 (N_16020,N_15805,N_15927);
nand U16021 (N_16021,N_15868,N_15933);
or U16022 (N_16022,N_15878,N_15861);
and U16023 (N_16023,N_15906,N_15986);
or U16024 (N_16024,N_15876,N_15851);
nand U16025 (N_16025,N_15847,N_15942);
and U16026 (N_16026,N_15802,N_15973);
or U16027 (N_16027,N_15993,N_15833);
xor U16028 (N_16028,N_15880,N_15940);
nand U16029 (N_16029,N_15931,N_15874);
xnor U16030 (N_16030,N_15862,N_15896);
nor U16031 (N_16031,N_15977,N_15855);
and U16032 (N_16032,N_15822,N_15803);
and U16033 (N_16033,N_15935,N_15913);
and U16034 (N_16034,N_15807,N_15804);
or U16035 (N_16035,N_15881,N_15966);
or U16036 (N_16036,N_15976,N_15869);
and U16037 (N_16037,N_15995,N_15967);
nand U16038 (N_16038,N_15988,N_15969);
xor U16039 (N_16039,N_15939,N_15835);
xnor U16040 (N_16040,N_15879,N_15809);
nand U16041 (N_16041,N_15800,N_15844);
xor U16042 (N_16042,N_15839,N_15836);
and U16043 (N_16043,N_15950,N_15936);
or U16044 (N_16044,N_15972,N_15842);
nand U16045 (N_16045,N_15832,N_15823);
nand U16046 (N_16046,N_15963,N_15998);
xor U16047 (N_16047,N_15850,N_15932);
xnor U16048 (N_16048,N_15905,N_15974);
or U16049 (N_16049,N_15830,N_15820);
or U16050 (N_16050,N_15915,N_15984);
nor U16051 (N_16051,N_15971,N_15907);
and U16052 (N_16052,N_15846,N_15947);
and U16053 (N_16053,N_15877,N_15852);
and U16054 (N_16054,N_15923,N_15866);
nand U16055 (N_16055,N_15854,N_15922);
nor U16056 (N_16056,N_15996,N_15858);
xor U16057 (N_16057,N_15801,N_15867);
nor U16058 (N_16058,N_15892,N_15916);
and U16059 (N_16059,N_15882,N_15814);
nand U16060 (N_16060,N_15938,N_15964);
or U16061 (N_16061,N_15944,N_15989);
xnor U16062 (N_16062,N_15997,N_15914);
and U16063 (N_16063,N_15899,N_15827);
and U16064 (N_16064,N_15828,N_15860);
or U16065 (N_16065,N_15991,N_15887);
and U16066 (N_16066,N_15812,N_15853);
nor U16067 (N_16067,N_15911,N_15958);
or U16068 (N_16068,N_15982,N_15817);
xnor U16069 (N_16069,N_15894,N_15841);
xnor U16070 (N_16070,N_15981,N_15840);
nor U16071 (N_16071,N_15810,N_15924);
nor U16072 (N_16072,N_15831,N_15960);
xnor U16073 (N_16073,N_15945,N_15904);
xor U16074 (N_16074,N_15864,N_15806);
xor U16075 (N_16075,N_15819,N_15908);
nor U16076 (N_16076,N_15909,N_15983);
nand U16077 (N_16077,N_15925,N_15897);
nand U16078 (N_16078,N_15901,N_15979);
nand U16079 (N_16079,N_15837,N_15808);
or U16080 (N_16080,N_15961,N_15953);
and U16081 (N_16081,N_15955,N_15957);
and U16082 (N_16082,N_15815,N_15875);
xnor U16083 (N_16083,N_15930,N_15968);
nor U16084 (N_16084,N_15934,N_15818);
or U16085 (N_16085,N_15872,N_15871);
nor U16086 (N_16086,N_15928,N_15941);
nor U16087 (N_16087,N_15856,N_15863);
and U16088 (N_16088,N_15929,N_15834);
nand U16089 (N_16089,N_15978,N_15884);
nor U16090 (N_16090,N_15919,N_15857);
xnor U16091 (N_16091,N_15937,N_15910);
or U16092 (N_16092,N_15890,N_15987);
xor U16093 (N_16093,N_15845,N_15849);
nor U16094 (N_16094,N_15873,N_15975);
nor U16095 (N_16095,N_15848,N_15943);
nor U16096 (N_16096,N_15952,N_15865);
nand U16097 (N_16097,N_15891,N_15954);
xnor U16098 (N_16098,N_15921,N_15816);
or U16099 (N_16099,N_15903,N_15912);
and U16100 (N_16100,N_15944,N_15997);
nand U16101 (N_16101,N_15962,N_15850);
or U16102 (N_16102,N_15854,N_15933);
xnor U16103 (N_16103,N_15874,N_15962);
nor U16104 (N_16104,N_15827,N_15975);
nand U16105 (N_16105,N_15823,N_15868);
nor U16106 (N_16106,N_15819,N_15920);
xor U16107 (N_16107,N_15906,N_15854);
nand U16108 (N_16108,N_15943,N_15948);
xnor U16109 (N_16109,N_15914,N_15880);
xor U16110 (N_16110,N_15807,N_15930);
nor U16111 (N_16111,N_15918,N_15864);
nor U16112 (N_16112,N_15868,N_15806);
nor U16113 (N_16113,N_15973,N_15873);
and U16114 (N_16114,N_15827,N_15878);
nor U16115 (N_16115,N_15838,N_15945);
xnor U16116 (N_16116,N_15833,N_15959);
or U16117 (N_16117,N_15856,N_15989);
and U16118 (N_16118,N_15931,N_15925);
nor U16119 (N_16119,N_15855,N_15858);
or U16120 (N_16120,N_15910,N_15892);
nor U16121 (N_16121,N_15981,N_15939);
and U16122 (N_16122,N_15850,N_15924);
and U16123 (N_16123,N_15882,N_15973);
nand U16124 (N_16124,N_15974,N_15887);
xor U16125 (N_16125,N_15885,N_15927);
nand U16126 (N_16126,N_15943,N_15813);
nor U16127 (N_16127,N_15948,N_15903);
nand U16128 (N_16128,N_15992,N_15839);
or U16129 (N_16129,N_15906,N_15964);
or U16130 (N_16130,N_15934,N_15937);
nor U16131 (N_16131,N_15897,N_15890);
or U16132 (N_16132,N_15807,N_15968);
and U16133 (N_16133,N_15886,N_15885);
and U16134 (N_16134,N_15884,N_15824);
nand U16135 (N_16135,N_15946,N_15872);
xor U16136 (N_16136,N_15987,N_15901);
and U16137 (N_16137,N_15970,N_15965);
or U16138 (N_16138,N_15930,N_15909);
and U16139 (N_16139,N_15817,N_15986);
nand U16140 (N_16140,N_15956,N_15909);
or U16141 (N_16141,N_15939,N_15982);
nor U16142 (N_16142,N_15824,N_15801);
nand U16143 (N_16143,N_15967,N_15905);
and U16144 (N_16144,N_15971,N_15875);
nand U16145 (N_16145,N_15832,N_15967);
and U16146 (N_16146,N_15800,N_15996);
xnor U16147 (N_16147,N_15811,N_15961);
nand U16148 (N_16148,N_15887,N_15914);
and U16149 (N_16149,N_15973,N_15916);
and U16150 (N_16150,N_15817,N_15812);
xnor U16151 (N_16151,N_15837,N_15948);
nor U16152 (N_16152,N_15922,N_15875);
nand U16153 (N_16153,N_15955,N_15800);
nor U16154 (N_16154,N_15826,N_15928);
and U16155 (N_16155,N_15846,N_15902);
and U16156 (N_16156,N_15891,N_15803);
and U16157 (N_16157,N_15985,N_15977);
xor U16158 (N_16158,N_15874,N_15908);
and U16159 (N_16159,N_15802,N_15995);
xor U16160 (N_16160,N_15988,N_15822);
nand U16161 (N_16161,N_15969,N_15939);
nand U16162 (N_16162,N_15814,N_15948);
nor U16163 (N_16163,N_15880,N_15912);
xor U16164 (N_16164,N_15905,N_15801);
and U16165 (N_16165,N_15867,N_15822);
nand U16166 (N_16166,N_15917,N_15815);
nand U16167 (N_16167,N_15884,N_15982);
and U16168 (N_16168,N_15972,N_15910);
nor U16169 (N_16169,N_15971,N_15883);
or U16170 (N_16170,N_15827,N_15969);
and U16171 (N_16171,N_15855,N_15823);
and U16172 (N_16172,N_15905,N_15868);
nand U16173 (N_16173,N_15906,N_15861);
nor U16174 (N_16174,N_15883,N_15811);
nor U16175 (N_16175,N_15878,N_15880);
and U16176 (N_16176,N_15979,N_15984);
nor U16177 (N_16177,N_15814,N_15847);
xor U16178 (N_16178,N_15868,N_15818);
or U16179 (N_16179,N_15940,N_15965);
nand U16180 (N_16180,N_15981,N_15883);
nand U16181 (N_16181,N_15877,N_15987);
or U16182 (N_16182,N_15876,N_15869);
nand U16183 (N_16183,N_15950,N_15992);
nor U16184 (N_16184,N_15984,N_15865);
nand U16185 (N_16185,N_15985,N_15873);
nor U16186 (N_16186,N_15805,N_15832);
xor U16187 (N_16187,N_15868,N_15901);
xor U16188 (N_16188,N_15860,N_15987);
xor U16189 (N_16189,N_15802,N_15877);
and U16190 (N_16190,N_15945,N_15975);
xor U16191 (N_16191,N_15978,N_15865);
or U16192 (N_16192,N_15839,N_15991);
nand U16193 (N_16193,N_15946,N_15832);
and U16194 (N_16194,N_15997,N_15825);
and U16195 (N_16195,N_15882,N_15888);
nand U16196 (N_16196,N_15867,N_15846);
and U16197 (N_16197,N_15950,N_15880);
nor U16198 (N_16198,N_15979,N_15821);
nor U16199 (N_16199,N_15820,N_15959);
nand U16200 (N_16200,N_16137,N_16150);
and U16201 (N_16201,N_16113,N_16091);
nor U16202 (N_16202,N_16136,N_16140);
nand U16203 (N_16203,N_16186,N_16104);
nand U16204 (N_16204,N_16081,N_16171);
nand U16205 (N_16205,N_16048,N_16120);
xor U16206 (N_16206,N_16138,N_16192);
nor U16207 (N_16207,N_16191,N_16036);
or U16208 (N_16208,N_16108,N_16094);
nor U16209 (N_16209,N_16143,N_16029);
nand U16210 (N_16210,N_16178,N_16039);
nand U16211 (N_16211,N_16055,N_16072);
and U16212 (N_16212,N_16043,N_16033);
and U16213 (N_16213,N_16118,N_16063);
nand U16214 (N_16214,N_16093,N_16031);
or U16215 (N_16215,N_16159,N_16044);
and U16216 (N_16216,N_16125,N_16129);
xor U16217 (N_16217,N_16126,N_16097);
nor U16218 (N_16218,N_16195,N_16042);
or U16219 (N_16219,N_16183,N_16080);
or U16220 (N_16220,N_16182,N_16088);
nand U16221 (N_16221,N_16051,N_16100);
nand U16222 (N_16222,N_16010,N_16151);
nand U16223 (N_16223,N_16034,N_16035);
nand U16224 (N_16224,N_16001,N_16181);
nand U16225 (N_16225,N_16199,N_16050);
and U16226 (N_16226,N_16180,N_16024);
nand U16227 (N_16227,N_16121,N_16185);
nand U16228 (N_16228,N_16076,N_16116);
nor U16229 (N_16229,N_16198,N_16047);
xor U16230 (N_16230,N_16066,N_16067);
or U16231 (N_16231,N_16015,N_16166);
xor U16232 (N_16232,N_16078,N_16188);
nor U16233 (N_16233,N_16065,N_16038);
or U16234 (N_16234,N_16197,N_16144);
nand U16235 (N_16235,N_16172,N_16148);
nand U16236 (N_16236,N_16106,N_16109);
nor U16237 (N_16237,N_16084,N_16013);
xnor U16238 (N_16238,N_16141,N_16187);
nor U16239 (N_16239,N_16053,N_16092);
nor U16240 (N_16240,N_16165,N_16134);
or U16241 (N_16241,N_16114,N_16023);
xnor U16242 (N_16242,N_16032,N_16018);
xnor U16243 (N_16243,N_16176,N_16160);
nor U16244 (N_16244,N_16008,N_16158);
and U16245 (N_16245,N_16028,N_16105);
and U16246 (N_16246,N_16027,N_16083);
or U16247 (N_16247,N_16014,N_16128);
or U16248 (N_16248,N_16194,N_16167);
nand U16249 (N_16249,N_16154,N_16095);
or U16250 (N_16250,N_16135,N_16087);
nor U16251 (N_16251,N_16006,N_16089);
nand U16252 (N_16252,N_16073,N_16062);
nor U16253 (N_16253,N_16085,N_16169);
and U16254 (N_16254,N_16012,N_16030);
nand U16255 (N_16255,N_16133,N_16068);
nor U16256 (N_16256,N_16102,N_16101);
or U16257 (N_16257,N_16082,N_16112);
or U16258 (N_16258,N_16170,N_16058);
and U16259 (N_16259,N_16161,N_16054);
nor U16260 (N_16260,N_16060,N_16079);
nand U16261 (N_16261,N_16074,N_16017);
xnor U16262 (N_16262,N_16179,N_16156);
or U16263 (N_16263,N_16070,N_16069);
nor U16264 (N_16264,N_16064,N_16146);
and U16265 (N_16265,N_16016,N_16174);
and U16266 (N_16266,N_16177,N_16077);
xor U16267 (N_16267,N_16004,N_16111);
and U16268 (N_16268,N_16021,N_16124);
nor U16269 (N_16269,N_16041,N_16020);
nand U16270 (N_16270,N_16196,N_16164);
xnor U16271 (N_16271,N_16071,N_16152);
or U16272 (N_16272,N_16184,N_16007);
nand U16273 (N_16273,N_16009,N_16190);
nor U16274 (N_16274,N_16022,N_16145);
nor U16275 (N_16275,N_16107,N_16149);
nor U16276 (N_16276,N_16189,N_16061);
nand U16277 (N_16277,N_16040,N_16011);
xor U16278 (N_16278,N_16163,N_16127);
or U16279 (N_16279,N_16115,N_16046);
nor U16280 (N_16280,N_16059,N_16086);
or U16281 (N_16281,N_16162,N_16131);
and U16282 (N_16282,N_16052,N_16110);
or U16283 (N_16283,N_16096,N_16056);
or U16284 (N_16284,N_16173,N_16005);
nand U16285 (N_16285,N_16142,N_16168);
or U16286 (N_16286,N_16119,N_16139);
nand U16287 (N_16287,N_16098,N_16099);
or U16288 (N_16288,N_16026,N_16132);
or U16289 (N_16289,N_16090,N_16123);
or U16290 (N_16290,N_16155,N_16075);
nor U16291 (N_16291,N_16057,N_16000);
and U16292 (N_16292,N_16019,N_16003);
xor U16293 (N_16293,N_16103,N_16193);
xor U16294 (N_16294,N_16045,N_16117);
xor U16295 (N_16295,N_16153,N_16049);
and U16296 (N_16296,N_16002,N_16147);
and U16297 (N_16297,N_16037,N_16130);
nor U16298 (N_16298,N_16157,N_16025);
nor U16299 (N_16299,N_16122,N_16175);
nor U16300 (N_16300,N_16165,N_16060);
nand U16301 (N_16301,N_16117,N_16110);
nor U16302 (N_16302,N_16192,N_16159);
nor U16303 (N_16303,N_16160,N_16068);
nor U16304 (N_16304,N_16039,N_16067);
xor U16305 (N_16305,N_16055,N_16147);
nand U16306 (N_16306,N_16152,N_16144);
xor U16307 (N_16307,N_16053,N_16082);
and U16308 (N_16308,N_16062,N_16150);
nor U16309 (N_16309,N_16075,N_16190);
nand U16310 (N_16310,N_16018,N_16105);
or U16311 (N_16311,N_16006,N_16199);
and U16312 (N_16312,N_16108,N_16115);
xnor U16313 (N_16313,N_16089,N_16037);
or U16314 (N_16314,N_16127,N_16181);
nor U16315 (N_16315,N_16160,N_16078);
nor U16316 (N_16316,N_16019,N_16022);
nor U16317 (N_16317,N_16092,N_16008);
or U16318 (N_16318,N_16187,N_16172);
xor U16319 (N_16319,N_16112,N_16015);
xor U16320 (N_16320,N_16072,N_16078);
nand U16321 (N_16321,N_16019,N_16163);
xor U16322 (N_16322,N_16036,N_16112);
nand U16323 (N_16323,N_16070,N_16122);
and U16324 (N_16324,N_16196,N_16070);
or U16325 (N_16325,N_16130,N_16034);
or U16326 (N_16326,N_16040,N_16073);
nor U16327 (N_16327,N_16064,N_16176);
or U16328 (N_16328,N_16109,N_16061);
xor U16329 (N_16329,N_16125,N_16081);
and U16330 (N_16330,N_16174,N_16112);
or U16331 (N_16331,N_16045,N_16107);
and U16332 (N_16332,N_16012,N_16112);
nor U16333 (N_16333,N_16077,N_16086);
nor U16334 (N_16334,N_16171,N_16197);
and U16335 (N_16335,N_16180,N_16001);
or U16336 (N_16336,N_16177,N_16135);
and U16337 (N_16337,N_16006,N_16039);
xnor U16338 (N_16338,N_16049,N_16074);
nand U16339 (N_16339,N_16085,N_16010);
or U16340 (N_16340,N_16025,N_16083);
or U16341 (N_16341,N_16081,N_16040);
nor U16342 (N_16342,N_16127,N_16166);
nor U16343 (N_16343,N_16022,N_16165);
xor U16344 (N_16344,N_16029,N_16002);
xor U16345 (N_16345,N_16035,N_16069);
xnor U16346 (N_16346,N_16078,N_16135);
nor U16347 (N_16347,N_16153,N_16087);
nor U16348 (N_16348,N_16007,N_16075);
or U16349 (N_16349,N_16071,N_16004);
and U16350 (N_16350,N_16152,N_16098);
or U16351 (N_16351,N_16113,N_16117);
and U16352 (N_16352,N_16011,N_16037);
or U16353 (N_16353,N_16066,N_16136);
nand U16354 (N_16354,N_16198,N_16094);
or U16355 (N_16355,N_16079,N_16180);
and U16356 (N_16356,N_16010,N_16144);
or U16357 (N_16357,N_16019,N_16160);
and U16358 (N_16358,N_16142,N_16028);
and U16359 (N_16359,N_16173,N_16054);
and U16360 (N_16360,N_16018,N_16046);
nand U16361 (N_16361,N_16166,N_16005);
nand U16362 (N_16362,N_16008,N_16053);
and U16363 (N_16363,N_16190,N_16140);
xor U16364 (N_16364,N_16098,N_16117);
nor U16365 (N_16365,N_16142,N_16071);
xnor U16366 (N_16366,N_16109,N_16003);
nor U16367 (N_16367,N_16082,N_16195);
nand U16368 (N_16368,N_16075,N_16188);
and U16369 (N_16369,N_16135,N_16006);
or U16370 (N_16370,N_16054,N_16163);
nand U16371 (N_16371,N_16116,N_16012);
or U16372 (N_16372,N_16125,N_16159);
or U16373 (N_16373,N_16184,N_16176);
or U16374 (N_16374,N_16082,N_16001);
nor U16375 (N_16375,N_16060,N_16091);
nor U16376 (N_16376,N_16072,N_16029);
and U16377 (N_16377,N_16124,N_16169);
and U16378 (N_16378,N_16098,N_16161);
nor U16379 (N_16379,N_16160,N_16076);
nand U16380 (N_16380,N_16044,N_16171);
nor U16381 (N_16381,N_16117,N_16154);
nor U16382 (N_16382,N_16055,N_16084);
or U16383 (N_16383,N_16178,N_16158);
or U16384 (N_16384,N_16134,N_16092);
nor U16385 (N_16385,N_16167,N_16098);
nand U16386 (N_16386,N_16039,N_16118);
or U16387 (N_16387,N_16146,N_16150);
nor U16388 (N_16388,N_16168,N_16061);
and U16389 (N_16389,N_16025,N_16146);
xnor U16390 (N_16390,N_16022,N_16060);
xor U16391 (N_16391,N_16101,N_16181);
or U16392 (N_16392,N_16096,N_16158);
nor U16393 (N_16393,N_16053,N_16170);
and U16394 (N_16394,N_16087,N_16170);
nor U16395 (N_16395,N_16195,N_16158);
and U16396 (N_16396,N_16181,N_16008);
nor U16397 (N_16397,N_16035,N_16027);
nand U16398 (N_16398,N_16126,N_16143);
nor U16399 (N_16399,N_16129,N_16040);
or U16400 (N_16400,N_16378,N_16237);
and U16401 (N_16401,N_16329,N_16294);
and U16402 (N_16402,N_16203,N_16296);
and U16403 (N_16403,N_16261,N_16395);
nor U16404 (N_16404,N_16327,N_16274);
nand U16405 (N_16405,N_16252,N_16390);
and U16406 (N_16406,N_16357,N_16368);
nand U16407 (N_16407,N_16371,N_16381);
or U16408 (N_16408,N_16302,N_16260);
nor U16409 (N_16409,N_16334,N_16212);
xor U16410 (N_16410,N_16267,N_16376);
nand U16411 (N_16411,N_16293,N_16306);
nand U16412 (N_16412,N_16385,N_16312);
and U16413 (N_16413,N_16367,N_16200);
or U16414 (N_16414,N_16298,N_16289);
nor U16415 (N_16415,N_16372,N_16325);
nand U16416 (N_16416,N_16382,N_16311);
and U16417 (N_16417,N_16251,N_16255);
or U16418 (N_16418,N_16288,N_16351);
nand U16419 (N_16419,N_16316,N_16309);
nand U16420 (N_16420,N_16343,N_16208);
xnor U16421 (N_16421,N_16389,N_16304);
nor U16422 (N_16422,N_16330,N_16340);
nor U16423 (N_16423,N_16213,N_16308);
and U16424 (N_16424,N_16265,N_16322);
nor U16425 (N_16425,N_16332,N_16204);
and U16426 (N_16426,N_16232,N_16290);
xor U16427 (N_16427,N_16380,N_16249);
and U16428 (N_16428,N_16353,N_16242);
and U16429 (N_16429,N_16276,N_16336);
nand U16430 (N_16430,N_16250,N_16226);
nand U16431 (N_16431,N_16373,N_16315);
xnor U16432 (N_16432,N_16358,N_16313);
or U16433 (N_16433,N_16225,N_16331);
nor U16434 (N_16434,N_16337,N_16346);
or U16435 (N_16435,N_16211,N_16361);
nand U16436 (N_16436,N_16206,N_16247);
nand U16437 (N_16437,N_16280,N_16391);
xnor U16438 (N_16438,N_16259,N_16349);
nor U16439 (N_16439,N_16301,N_16221);
or U16440 (N_16440,N_16374,N_16317);
nand U16441 (N_16441,N_16362,N_16207);
nor U16442 (N_16442,N_16239,N_16297);
nand U16443 (N_16443,N_16364,N_16269);
nor U16444 (N_16444,N_16366,N_16360);
or U16445 (N_16445,N_16256,N_16314);
and U16446 (N_16446,N_16214,N_16227);
xor U16447 (N_16447,N_16359,N_16278);
xor U16448 (N_16448,N_16338,N_16347);
xnor U16449 (N_16449,N_16348,N_16219);
or U16450 (N_16450,N_16216,N_16234);
nor U16451 (N_16451,N_16210,N_16393);
xor U16452 (N_16452,N_16396,N_16285);
and U16453 (N_16453,N_16377,N_16277);
nor U16454 (N_16454,N_16248,N_16272);
or U16455 (N_16455,N_16355,N_16310);
and U16456 (N_16456,N_16392,N_16258);
xor U16457 (N_16457,N_16339,N_16320);
or U16458 (N_16458,N_16354,N_16209);
and U16459 (N_16459,N_16292,N_16341);
and U16460 (N_16460,N_16246,N_16344);
and U16461 (N_16461,N_16370,N_16375);
or U16462 (N_16462,N_16387,N_16223);
or U16463 (N_16463,N_16397,N_16202);
nor U16464 (N_16464,N_16238,N_16275);
nor U16465 (N_16465,N_16319,N_16240);
xnor U16466 (N_16466,N_16384,N_16201);
nor U16467 (N_16467,N_16318,N_16222);
xor U16468 (N_16468,N_16388,N_16352);
nand U16469 (N_16469,N_16263,N_16271);
nand U16470 (N_16470,N_16399,N_16365);
xor U16471 (N_16471,N_16287,N_16386);
or U16472 (N_16472,N_16253,N_16335);
nand U16473 (N_16473,N_16229,N_16282);
nand U16474 (N_16474,N_16262,N_16363);
nor U16475 (N_16475,N_16205,N_16398);
nor U16476 (N_16476,N_16286,N_16270);
xor U16477 (N_16477,N_16356,N_16300);
xor U16478 (N_16478,N_16228,N_16236);
and U16479 (N_16479,N_16273,N_16235);
and U16480 (N_16480,N_16283,N_16350);
or U16481 (N_16481,N_16254,N_16379);
nor U16482 (N_16482,N_16243,N_16326);
xor U16483 (N_16483,N_16279,N_16342);
xnor U16484 (N_16484,N_16217,N_16244);
xor U16485 (N_16485,N_16224,N_16215);
xnor U16486 (N_16486,N_16284,N_16369);
nor U16487 (N_16487,N_16333,N_16257);
or U16488 (N_16488,N_16307,N_16266);
nand U16489 (N_16489,N_16321,N_16305);
or U16490 (N_16490,N_16264,N_16323);
xnor U16491 (N_16491,N_16383,N_16345);
nand U16492 (N_16492,N_16268,N_16241);
xnor U16493 (N_16493,N_16233,N_16245);
xnor U16494 (N_16494,N_16394,N_16281);
or U16495 (N_16495,N_16295,N_16324);
nand U16496 (N_16496,N_16220,N_16218);
nand U16497 (N_16497,N_16291,N_16299);
and U16498 (N_16498,N_16303,N_16231);
or U16499 (N_16499,N_16328,N_16230);
xor U16500 (N_16500,N_16211,N_16278);
xnor U16501 (N_16501,N_16378,N_16208);
xnor U16502 (N_16502,N_16243,N_16319);
nand U16503 (N_16503,N_16225,N_16349);
xnor U16504 (N_16504,N_16306,N_16397);
nand U16505 (N_16505,N_16240,N_16330);
or U16506 (N_16506,N_16347,N_16344);
nor U16507 (N_16507,N_16368,N_16242);
nand U16508 (N_16508,N_16260,N_16317);
nand U16509 (N_16509,N_16255,N_16204);
nand U16510 (N_16510,N_16378,N_16373);
xor U16511 (N_16511,N_16301,N_16277);
xnor U16512 (N_16512,N_16357,N_16249);
and U16513 (N_16513,N_16346,N_16252);
and U16514 (N_16514,N_16331,N_16297);
and U16515 (N_16515,N_16339,N_16227);
and U16516 (N_16516,N_16341,N_16200);
nand U16517 (N_16517,N_16304,N_16328);
nand U16518 (N_16518,N_16204,N_16358);
nand U16519 (N_16519,N_16370,N_16206);
and U16520 (N_16520,N_16292,N_16296);
nor U16521 (N_16521,N_16271,N_16315);
nand U16522 (N_16522,N_16237,N_16218);
or U16523 (N_16523,N_16287,N_16344);
or U16524 (N_16524,N_16245,N_16372);
xnor U16525 (N_16525,N_16214,N_16272);
nor U16526 (N_16526,N_16394,N_16384);
xor U16527 (N_16527,N_16300,N_16293);
xor U16528 (N_16528,N_16294,N_16269);
nor U16529 (N_16529,N_16317,N_16346);
nor U16530 (N_16530,N_16294,N_16277);
nand U16531 (N_16531,N_16229,N_16270);
nor U16532 (N_16532,N_16242,N_16323);
or U16533 (N_16533,N_16380,N_16245);
xnor U16534 (N_16534,N_16282,N_16291);
nor U16535 (N_16535,N_16279,N_16386);
and U16536 (N_16536,N_16245,N_16293);
nand U16537 (N_16537,N_16391,N_16378);
or U16538 (N_16538,N_16296,N_16367);
and U16539 (N_16539,N_16263,N_16241);
nor U16540 (N_16540,N_16285,N_16258);
nand U16541 (N_16541,N_16231,N_16315);
xnor U16542 (N_16542,N_16211,N_16349);
and U16543 (N_16543,N_16200,N_16252);
and U16544 (N_16544,N_16260,N_16323);
or U16545 (N_16545,N_16322,N_16201);
or U16546 (N_16546,N_16299,N_16218);
xor U16547 (N_16547,N_16326,N_16307);
nor U16548 (N_16548,N_16201,N_16205);
nand U16549 (N_16549,N_16387,N_16339);
xnor U16550 (N_16550,N_16211,N_16228);
xnor U16551 (N_16551,N_16334,N_16209);
xnor U16552 (N_16552,N_16329,N_16228);
nand U16553 (N_16553,N_16383,N_16232);
nor U16554 (N_16554,N_16230,N_16204);
or U16555 (N_16555,N_16200,N_16259);
or U16556 (N_16556,N_16366,N_16248);
nor U16557 (N_16557,N_16227,N_16219);
nor U16558 (N_16558,N_16266,N_16210);
and U16559 (N_16559,N_16268,N_16210);
or U16560 (N_16560,N_16307,N_16380);
xor U16561 (N_16561,N_16256,N_16223);
nand U16562 (N_16562,N_16346,N_16233);
and U16563 (N_16563,N_16252,N_16332);
and U16564 (N_16564,N_16388,N_16316);
xnor U16565 (N_16565,N_16313,N_16210);
nor U16566 (N_16566,N_16211,N_16219);
or U16567 (N_16567,N_16394,N_16218);
nand U16568 (N_16568,N_16270,N_16365);
nand U16569 (N_16569,N_16341,N_16317);
and U16570 (N_16570,N_16377,N_16282);
xor U16571 (N_16571,N_16336,N_16258);
nor U16572 (N_16572,N_16340,N_16262);
nor U16573 (N_16573,N_16275,N_16333);
or U16574 (N_16574,N_16251,N_16315);
nand U16575 (N_16575,N_16341,N_16395);
and U16576 (N_16576,N_16269,N_16389);
or U16577 (N_16577,N_16330,N_16304);
nand U16578 (N_16578,N_16397,N_16388);
or U16579 (N_16579,N_16310,N_16242);
or U16580 (N_16580,N_16325,N_16364);
or U16581 (N_16581,N_16206,N_16268);
and U16582 (N_16582,N_16201,N_16364);
and U16583 (N_16583,N_16308,N_16236);
xor U16584 (N_16584,N_16293,N_16307);
and U16585 (N_16585,N_16205,N_16257);
nand U16586 (N_16586,N_16296,N_16210);
xnor U16587 (N_16587,N_16381,N_16220);
or U16588 (N_16588,N_16352,N_16258);
xor U16589 (N_16589,N_16288,N_16298);
nor U16590 (N_16590,N_16230,N_16248);
and U16591 (N_16591,N_16338,N_16342);
xnor U16592 (N_16592,N_16224,N_16330);
nor U16593 (N_16593,N_16215,N_16298);
xnor U16594 (N_16594,N_16223,N_16309);
or U16595 (N_16595,N_16381,N_16321);
or U16596 (N_16596,N_16285,N_16200);
nor U16597 (N_16597,N_16279,N_16206);
nand U16598 (N_16598,N_16262,N_16304);
xor U16599 (N_16599,N_16355,N_16369);
or U16600 (N_16600,N_16537,N_16492);
nor U16601 (N_16601,N_16437,N_16496);
and U16602 (N_16602,N_16412,N_16490);
xnor U16603 (N_16603,N_16548,N_16536);
and U16604 (N_16604,N_16572,N_16554);
nor U16605 (N_16605,N_16481,N_16567);
nor U16606 (N_16606,N_16491,N_16578);
xor U16607 (N_16607,N_16580,N_16558);
nand U16608 (N_16608,N_16555,N_16478);
and U16609 (N_16609,N_16411,N_16522);
nor U16610 (N_16610,N_16458,N_16594);
or U16611 (N_16611,N_16533,N_16428);
nor U16612 (N_16612,N_16585,N_16447);
nor U16613 (N_16613,N_16520,N_16511);
or U16614 (N_16614,N_16429,N_16579);
nand U16615 (N_16615,N_16484,N_16436);
nor U16616 (N_16616,N_16507,N_16530);
xor U16617 (N_16617,N_16434,N_16472);
xor U16618 (N_16618,N_16591,N_16423);
nand U16619 (N_16619,N_16486,N_16430);
or U16620 (N_16620,N_16444,N_16476);
xor U16621 (N_16621,N_16512,N_16577);
and U16622 (N_16622,N_16466,N_16535);
nand U16623 (N_16623,N_16420,N_16559);
and U16624 (N_16624,N_16531,N_16457);
nand U16625 (N_16625,N_16564,N_16431);
nand U16626 (N_16626,N_16575,N_16570);
or U16627 (N_16627,N_16583,N_16584);
nand U16628 (N_16628,N_16422,N_16549);
and U16629 (N_16629,N_16506,N_16401);
and U16630 (N_16630,N_16552,N_16526);
xor U16631 (N_16631,N_16442,N_16596);
xor U16632 (N_16632,N_16427,N_16510);
nor U16633 (N_16633,N_16569,N_16474);
nand U16634 (N_16634,N_16438,N_16505);
and U16635 (N_16635,N_16471,N_16545);
or U16636 (N_16636,N_16400,N_16519);
nor U16637 (N_16637,N_16404,N_16456);
nor U16638 (N_16638,N_16599,N_16460);
or U16639 (N_16639,N_16413,N_16573);
and U16640 (N_16640,N_16527,N_16433);
or U16641 (N_16641,N_16547,N_16403);
and U16642 (N_16642,N_16516,N_16419);
nor U16643 (N_16643,N_16452,N_16406);
nand U16644 (N_16644,N_16528,N_16565);
xnor U16645 (N_16645,N_16539,N_16508);
nand U16646 (N_16646,N_16502,N_16524);
or U16647 (N_16647,N_16482,N_16415);
xor U16648 (N_16648,N_16475,N_16513);
xnor U16649 (N_16649,N_16521,N_16538);
or U16650 (N_16650,N_16414,N_16529);
nand U16651 (N_16651,N_16409,N_16473);
nand U16652 (N_16652,N_16553,N_16421);
nor U16653 (N_16653,N_16542,N_16417);
nand U16654 (N_16654,N_16590,N_16501);
nor U16655 (N_16655,N_16546,N_16557);
nor U16656 (N_16656,N_16525,N_16418);
or U16657 (N_16657,N_16509,N_16532);
nand U16658 (N_16658,N_16461,N_16445);
and U16659 (N_16659,N_16487,N_16483);
xnor U16660 (N_16660,N_16534,N_16504);
nand U16661 (N_16661,N_16551,N_16459);
xor U16662 (N_16662,N_16435,N_16440);
or U16663 (N_16663,N_16499,N_16402);
nor U16664 (N_16664,N_16497,N_16463);
nand U16665 (N_16665,N_16550,N_16480);
or U16666 (N_16666,N_16518,N_16470);
nor U16667 (N_16667,N_16540,N_16592);
nor U16668 (N_16668,N_16581,N_16448);
or U16669 (N_16669,N_16468,N_16465);
xor U16670 (N_16670,N_16439,N_16543);
xnor U16671 (N_16671,N_16494,N_16561);
and U16672 (N_16672,N_16574,N_16449);
or U16673 (N_16673,N_16597,N_16443);
nand U16674 (N_16674,N_16563,N_16562);
nand U16675 (N_16675,N_16560,N_16598);
nand U16676 (N_16676,N_16489,N_16582);
and U16677 (N_16677,N_16407,N_16462);
or U16678 (N_16678,N_16451,N_16593);
or U16679 (N_16679,N_16450,N_16405);
or U16680 (N_16680,N_16587,N_16424);
xor U16681 (N_16681,N_16576,N_16426);
or U16682 (N_16682,N_16541,N_16477);
and U16683 (N_16683,N_16453,N_16514);
and U16684 (N_16684,N_16515,N_16568);
and U16685 (N_16685,N_16454,N_16523);
and U16686 (N_16686,N_16467,N_16469);
nor U16687 (N_16687,N_16455,N_16408);
or U16688 (N_16688,N_16432,N_16446);
nand U16689 (N_16689,N_16416,N_16488);
xor U16690 (N_16690,N_16479,N_16464);
or U16691 (N_16691,N_16589,N_16498);
and U16692 (N_16692,N_16425,N_16500);
and U16693 (N_16693,N_16571,N_16556);
nor U16694 (N_16694,N_16517,N_16566);
and U16695 (N_16695,N_16588,N_16441);
and U16696 (N_16696,N_16586,N_16595);
or U16697 (N_16697,N_16485,N_16493);
and U16698 (N_16698,N_16503,N_16410);
xor U16699 (N_16699,N_16495,N_16544);
nor U16700 (N_16700,N_16478,N_16406);
nor U16701 (N_16701,N_16585,N_16471);
nor U16702 (N_16702,N_16516,N_16532);
nor U16703 (N_16703,N_16487,N_16572);
or U16704 (N_16704,N_16428,N_16410);
or U16705 (N_16705,N_16470,N_16431);
or U16706 (N_16706,N_16531,N_16420);
nor U16707 (N_16707,N_16455,N_16517);
or U16708 (N_16708,N_16555,N_16498);
and U16709 (N_16709,N_16421,N_16520);
xnor U16710 (N_16710,N_16510,N_16506);
or U16711 (N_16711,N_16496,N_16526);
or U16712 (N_16712,N_16592,N_16432);
or U16713 (N_16713,N_16551,N_16597);
or U16714 (N_16714,N_16488,N_16539);
nor U16715 (N_16715,N_16574,N_16466);
nor U16716 (N_16716,N_16581,N_16522);
nand U16717 (N_16717,N_16406,N_16403);
and U16718 (N_16718,N_16548,N_16410);
nor U16719 (N_16719,N_16504,N_16583);
nor U16720 (N_16720,N_16420,N_16410);
nor U16721 (N_16721,N_16555,N_16458);
and U16722 (N_16722,N_16418,N_16483);
nor U16723 (N_16723,N_16513,N_16533);
and U16724 (N_16724,N_16516,N_16400);
nand U16725 (N_16725,N_16496,N_16459);
and U16726 (N_16726,N_16565,N_16487);
nor U16727 (N_16727,N_16454,N_16411);
and U16728 (N_16728,N_16551,N_16596);
or U16729 (N_16729,N_16474,N_16544);
or U16730 (N_16730,N_16411,N_16563);
nand U16731 (N_16731,N_16403,N_16553);
nor U16732 (N_16732,N_16589,N_16501);
or U16733 (N_16733,N_16471,N_16432);
and U16734 (N_16734,N_16509,N_16468);
nor U16735 (N_16735,N_16497,N_16534);
nand U16736 (N_16736,N_16543,N_16552);
nor U16737 (N_16737,N_16467,N_16495);
nand U16738 (N_16738,N_16496,N_16539);
xor U16739 (N_16739,N_16441,N_16568);
or U16740 (N_16740,N_16470,N_16591);
nand U16741 (N_16741,N_16430,N_16488);
and U16742 (N_16742,N_16559,N_16479);
nor U16743 (N_16743,N_16532,N_16429);
and U16744 (N_16744,N_16480,N_16584);
xor U16745 (N_16745,N_16409,N_16493);
nand U16746 (N_16746,N_16540,N_16522);
nand U16747 (N_16747,N_16587,N_16527);
nor U16748 (N_16748,N_16569,N_16463);
or U16749 (N_16749,N_16556,N_16409);
and U16750 (N_16750,N_16404,N_16485);
nor U16751 (N_16751,N_16449,N_16542);
or U16752 (N_16752,N_16530,N_16430);
or U16753 (N_16753,N_16484,N_16497);
nor U16754 (N_16754,N_16530,N_16553);
xnor U16755 (N_16755,N_16487,N_16535);
xor U16756 (N_16756,N_16474,N_16461);
and U16757 (N_16757,N_16447,N_16475);
nor U16758 (N_16758,N_16426,N_16584);
nor U16759 (N_16759,N_16409,N_16454);
xor U16760 (N_16760,N_16550,N_16502);
nand U16761 (N_16761,N_16465,N_16409);
or U16762 (N_16762,N_16497,N_16574);
nor U16763 (N_16763,N_16524,N_16586);
nand U16764 (N_16764,N_16487,N_16449);
and U16765 (N_16765,N_16570,N_16549);
xnor U16766 (N_16766,N_16477,N_16418);
xnor U16767 (N_16767,N_16436,N_16576);
nor U16768 (N_16768,N_16424,N_16536);
xor U16769 (N_16769,N_16463,N_16570);
and U16770 (N_16770,N_16540,N_16586);
or U16771 (N_16771,N_16598,N_16456);
nand U16772 (N_16772,N_16564,N_16414);
nand U16773 (N_16773,N_16500,N_16449);
or U16774 (N_16774,N_16410,N_16485);
and U16775 (N_16775,N_16539,N_16500);
nor U16776 (N_16776,N_16414,N_16496);
or U16777 (N_16777,N_16427,N_16553);
nor U16778 (N_16778,N_16570,N_16578);
or U16779 (N_16779,N_16488,N_16424);
xnor U16780 (N_16780,N_16447,N_16501);
nor U16781 (N_16781,N_16597,N_16528);
nand U16782 (N_16782,N_16500,N_16590);
nand U16783 (N_16783,N_16484,N_16590);
nor U16784 (N_16784,N_16510,N_16527);
nand U16785 (N_16785,N_16594,N_16439);
and U16786 (N_16786,N_16498,N_16426);
or U16787 (N_16787,N_16530,N_16417);
nor U16788 (N_16788,N_16405,N_16475);
or U16789 (N_16789,N_16451,N_16468);
nand U16790 (N_16790,N_16559,N_16489);
nor U16791 (N_16791,N_16403,N_16539);
nand U16792 (N_16792,N_16591,N_16560);
nor U16793 (N_16793,N_16529,N_16503);
or U16794 (N_16794,N_16427,N_16538);
nor U16795 (N_16795,N_16569,N_16496);
and U16796 (N_16796,N_16576,N_16465);
or U16797 (N_16797,N_16459,N_16476);
or U16798 (N_16798,N_16400,N_16574);
and U16799 (N_16799,N_16461,N_16451);
xnor U16800 (N_16800,N_16637,N_16731);
and U16801 (N_16801,N_16641,N_16600);
nor U16802 (N_16802,N_16693,N_16691);
and U16803 (N_16803,N_16700,N_16710);
or U16804 (N_16804,N_16790,N_16771);
or U16805 (N_16805,N_16758,N_16772);
or U16806 (N_16806,N_16698,N_16602);
nor U16807 (N_16807,N_16669,N_16682);
nand U16808 (N_16808,N_16715,N_16639);
xnor U16809 (N_16809,N_16777,N_16621);
nor U16810 (N_16810,N_16774,N_16782);
nand U16811 (N_16811,N_16615,N_16714);
or U16812 (N_16812,N_16666,N_16634);
nor U16813 (N_16813,N_16694,N_16651);
xor U16814 (N_16814,N_16762,N_16675);
nor U16815 (N_16815,N_16661,N_16635);
and U16816 (N_16816,N_16649,N_16724);
and U16817 (N_16817,N_16722,N_16644);
nand U16818 (N_16818,N_16659,N_16619);
nand U16819 (N_16819,N_16748,N_16640);
or U16820 (N_16820,N_16629,N_16791);
nor U16821 (N_16821,N_16753,N_16618);
xnor U16822 (N_16822,N_16628,N_16674);
nand U16823 (N_16823,N_16797,N_16717);
xor U16824 (N_16824,N_16787,N_16750);
nor U16825 (N_16825,N_16609,N_16733);
xnor U16826 (N_16826,N_16789,N_16729);
and U16827 (N_16827,N_16712,N_16792);
nor U16828 (N_16828,N_16743,N_16799);
and U16829 (N_16829,N_16763,N_16678);
or U16830 (N_16830,N_16650,N_16784);
or U16831 (N_16831,N_16677,N_16760);
xnor U16832 (N_16832,N_16648,N_16670);
or U16833 (N_16833,N_16721,N_16645);
and U16834 (N_16834,N_16632,N_16720);
xnor U16835 (N_16835,N_16690,N_16657);
and U16836 (N_16836,N_16739,N_16770);
nand U16837 (N_16837,N_16779,N_16627);
nor U16838 (N_16838,N_16668,N_16671);
nand U16839 (N_16839,N_16686,N_16741);
nor U16840 (N_16840,N_16667,N_16624);
nor U16841 (N_16841,N_16613,N_16765);
nor U16842 (N_16842,N_16601,N_16630);
or U16843 (N_16843,N_16692,N_16764);
xor U16844 (N_16844,N_16633,N_16704);
and U16845 (N_16845,N_16785,N_16728);
nor U16846 (N_16846,N_16681,N_16747);
nand U16847 (N_16847,N_16798,N_16773);
xor U16848 (N_16848,N_16688,N_16620);
xor U16849 (N_16849,N_16673,N_16737);
or U16850 (N_16850,N_16796,N_16746);
and U16851 (N_16851,N_16638,N_16723);
or U16852 (N_16852,N_16608,N_16756);
nand U16853 (N_16853,N_16636,N_16744);
nor U16854 (N_16854,N_16749,N_16709);
xnor U16855 (N_16855,N_16658,N_16734);
nand U16856 (N_16856,N_16718,N_16625);
and U16857 (N_16857,N_16769,N_16663);
or U16858 (N_16858,N_16786,N_16727);
nand U16859 (N_16859,N_16738,N_16626);
or U16860 (N_16860,N_16730,N_16684);
nor U16861 (N_16861,N_16788,N_16654);
xnor U16862 (N_16862,N_16755,N_16612);
nor U16863 (N_16863,N_16719,N_16604);
xor U16864 (N_16864,N_16754,N_16707);
xnor U16865 (N_16865,N_16696,N_16680);
xnor U16866 (N_16866,N_16685,N_16713);
xnor U16867 (N_16867,N_16793,N_16795);
nor U16868 (N_16868,N_16701,N_16664);
and U16869 (N_16869,N_16776,N_16647);
xor U16870 (N_16870,N_16605,N_16736);
nor U16871 (N_16871,N_16726,N_16652);
nor U16872 (N_16872,N_16706,N_16689);
or U16873 (N_16873,N_16665,N_16606);
or U16874 (N_16874,N_16614,N_16643);
nor U16875 (N_16875,N_16607,N_16646);
xnor U16876 (N_16876,N_16617,N_16603);
nor U16877 (N_16877,N_16716,N_16699);
and U16878 (N_16878,N_16768,N_16757);
or U16879 (N_16879,N_16705,N_16759);
or U16880 (N_16880,N_16735,N_16611);
xnor U16881 (N_16881,N_16778,N_16697);
nand U16882 (N_16882,N_16631,N_16708);
xor U16883 (N_16883,N_16655,N_16662);
or U16884 (N_16884,N_16687,N_16745);
nor U16885 (N_16885,N_16725,N_16767);
and U16886 (N_16886,N_16642,N_16653);
or U16887 (N_16887,N_16683,N_16775);
nor U16888 (N_16888,N_16740,N_16623);
nand U16889 (N_16889,N_16660,N_16766);
nor U16890 (N_16890,N_16742,N_16679);
nand U16891 (N_16891,N_16711,N_16794);
nand U16892 (N_16892,N_16751,N_16676);
and U16893 (N_16893,N_16781,N_16622);
nor U16894 (N_16894,N_16695,N_16672);
and U16895 (N_16895,N_16656,N_16780);
and U16896 (N_16896,N_16752,N_16702);
xnor U16897 (N_16897,N_16616,N_16703);
nor U16898 (N_16898,N_16732,N_16783);
or U16899 (N_16899,N_16610,N_16761);
nand U16900 (N_16900,N_16791,N_16656);
xnor U16901 (N_16901,N_16727,N_16746);
xor U16902 (N_16902,N_16766,N_16633);
nand U16903 (N_16903,N_16768,N_16711);
or U16904 (N_16904,N_16633,N_16728);
nor U16905 (N_16905,N_16653,N_16661);
or U16906 (N_16906,N_16732,N_16640);
nand U16907 (N_16907,N_16604,N_16773);
and U16908 (N_16908,N_16664,N_16705);
nor U16909 (N_16909,N_16766,N_16787);
or U16910 (N_16910,N_16640,N_16633);
xnor U16911 (N_16911,N_16703,N_16639);
or U16912 (N_16912,N_16742,N_16797);
xnor U16913 (N_16913,N_16678,N_16648);
nand U16914 (N_16914,N_16681,N_16632);
nand U16915 (N_16915,N_16655,N_16637);
xnor U16916 (N_16916,N_16634,N_16639);
xnor U16917 (N_16917,N_16665,N_16702);
or U16918 (N_16918,N_16624,N_16619);
xor U16919 (N_16919,N_16627,N_16687);
or U16920 (N_16920,N_16779,N_16689);
nor U16921 (N_16921,N_16797,N_16671);
or U16922 (N_16922,N_16664,N_16656);
nor U16923 (N_16923,N_16741,N_16647);
nand U16924 (N_16924,N_16607,N_16624);
or U16925 (N_16925,N_16756,N_16795);
nor U16926 (N_16926,N_16657,N_16653);
nand U16927 (N_16927,N_16609,N_16765);
nor U16928 (N_16928,N_16706,N_16779);
nand U16929 (N_16929,N_16738,N_16755);
xnor U16930 (N_16930,N_16650,N_16627);
and U16931 (N_16931,N_16670,N_16626);
nor U16932 (N_16932,N_16766,N_16750);
nor U16933 (N_16933,N_16627,N_16787);
or U16934 (N_16934,N_16609,N_16707);
or U16935 (N_16935,N_16701,N_16692);
and U16936 (N_16936,N_16604,N_16778);
nor U16937 (N_16937,N_16687,N_16689);
nor U16938 (N_16938,N_16627,N_16781);
or U16939 (N_16939,N_16712,N_16716);
xnor U16940 (N_16940,N_16684,N_16690);
nor U16941 (N_16941,N_16700,N_16660);
nor U16942 (N_16942,N_16704,N_16722);
and U16943 (N_16943,N_16669,N_16665);
nor U16944 (N_16944,N_16714,N_16782);
nor U16945 (N_16945,N_16607,N_16681);
or U16946 (N_16946,N_16733,N_16672);
xnor U16947 (N_16947,N_16625,N_16787);
nor U16948 (N_16948,N_16748,N_16661);
xnor U16949 (N_16949,N_16772,N_16694);
or U16950 (N_16950,N_16707,N_16652);
nor U16951 (N_16951,N_16744,N_16773);
xnor U16952 (N_16952,N_16716,N_16612);
nand U16953 (N_16953,N_16784,N_16756);
or U16954 (N_16954,N_16694,N_16734);
nor U16955 (N_16955,N_16727,N_16709);
and U16956 (N_16956,N_16749,N_16613);
nand U16957 (N_16957,N_16716,N_16606);
or U16958 (N_16958,N_16681,N_16623);
xor U16959 (N_16959,N_16771,N_16696);
xnor U16960 (N_16960,N_16638,N_16745);
nor U16961 (N_16961,N_16730,N_16621);
nor U16962 (N_16962,N_16605,N_16676);
nor U16963 (N_16963,N_16605,N_16794);
nand U16964 (N_16964,N_16752,N_16759);
or U16965 (N_16965,N_16636,N_16709);
xor U16966 (N_16966,N_16705,N_16706);
nor U16967 (N_16967,N_16609,N_16708);
nor U16968 (N_16968,N_16772,N_16689);
or U16969 (N_16969,N_16723,N_16776);
or U16970 (N_16970,N_16672,N_16603);
nand U16971 (N_16971,N_16762,N_16622);
and U16972 (N_16972,N_16661,N_16698);
nand U16973 (N_16973,N_16632,N_16612);
nand U16974 (N_16974,N_16633,N_16606);
xor U16975 (N_16975,N_16690,N_16770);
nor U16976 (N_16976,N_16776,N_16645);
or U16977 (N_16977,N_16639,N_16767);
nor U16978 (N_16978,N_16761,N_16650);
and U16979 (N_16979,N_16681,N_16612);
or U16980 (N_16980,N_16737,N_16690);
nor U16981 (N_16981,N_16795,N_16767);
and U16982 (N_16982,N_16723,N_16655);
nor U16983 (N_16983,N_16729,N_16643);
nor U16984 (N_16984,N_16686,N_16743);
xor U16985 (N_16985,N_16691,N_16787);
and U16986 (N_16986,N_16795,N_16615);
or U16987 (N_16987,N_16753,N_16679);
xnor U16988 (N_16988,N_16665,N_16773);
xnor U16989 (N_16989,N_16674,N_16786);
xor U16990 (N_16990,N_16642,N_16772);
or U16991 (N_16991,N_16620,N_16788);
nor U16992 (N_16992,N_16681,N_16663);
nand U16993 (N_16993,N_16618,N_16653);
nor U16994 (N_16994,N_16723,N_16793);
or U16995 (N_16995,N_16616,N_16744);
and U16996 (N_16996,N_16706,N_16692);
or U16997 (N_16997,N_16659,N_16626);
or U16998 (N_16998,N_16721,N_16703);
or U16999 (N_16999,N_16722,N_16677);
nor U17000 (N_17000,N_16909,N_16838);
and U17001 (N_17001,N_16976,N_16898);
nor U17002 (N_17002,N_16982,N_16888);
xor U17003 (N_17003,N_16843,N_16808);
or U17004 (N_17004,N_16887,N_16827);
nor U17005 (N_17005,N_16980,N_16880);
nand U17006 (N_17006,N_16992,N_16983);
or U17007 (N_17007,N_16846,N_16943);
and U17008 (N_17008,N_16938,N_16975);
nand U17009 (N_17009,N_16879,N_16963);
xor U17010 (N_17010,N_16860,N_16806);
nor U17011 (N_17011,N_16886,N_16930);
nor U17012 (N_17012,N_16825,N_16807);
nor U17013 (N_17013,N_16834,N_16997);
nand U17014 (N_17014,N_16826,N_16899);
nor U17015 (N_17015,N_16922,N_16839);
and U17016 (N_17016,N_16931,N_16881);
nor U17017 (N_17017,N_16958,N_16856);
xor U17018 (N_17018,N_16837,N_16999);
and U17019 (N_17019,N_16893,N_16845);
and U17020 (N_17020,N_16900,N_16944);
xor U17021 (N_17021,N_16853,N_16818);
nor U17022 (N_17022,N_16965,N_16923);
and U17023 (N_17023,N_16959,N_16863);
or U17024 (N_17024,N_16800,N_16932);
nor U17025 (N_17025,N_16934,N_16957);
nor U17026 (N_17026,N_16941,N_16830);
and U17027 (N_17027,N_16949,N_16950);
xnor U17028 (N_17028,N_16815,N_16872);
or U17029 (N_17029,N_16862,N_16884);
xnor U17030 (N_17030,N_16969,N_16882);
nor U17031 (N_17031,N_16803,N_16964);
or U17032 (N_17032,N_16935,N_16876);
or U17033 (N_17033,N_16877,N_16927);
nand U17034 (N_17034,N_16924,N_16849);
or U17035 (N_17035,N_16991,N_16841);
nand U17036 (N_17036,N_16988,N_16937);
or U17037 (N_17037,N_16809,N_16821);
nand U17038 (N_17038,N_16817,N_16867);
nand U17039 (N_17039,N_16891,N_16955);
and U17040 (N_17040,N_16917,N_16870);
and U17041 (N_17041,N_16933,N_16953);
or U17042 (N_17042,N_16996,N_16858);
and U17043 (N_17043,N_16844,N_16819);
nor U17044 (N_17044,N_16993,N_16961);
nor U17045 (N_17045,N_16812,N_16972);
nor U17046 (N_17046,N_16810,N_16901);
nand U17047 (N_17047,N_16904,N_16866);
and U17048 (N_17048,N_16912,N_16948);
or U17049 (N_17049,N_16921,N_16820);
xor U17050 (N_17050,N_16851,N_16928);
nand U17051 (N_17051,N_16929,N_16805);
or U17052 (N_17052,N_16977,N_16801);
or U17053 (N_17053,N_16926,N_16911);
xor U17054 (N_17054,N_16962,N_16871);
and U17055 (N_17055,N_16954,N_16908);
xnor U17056 (N_17056,N_16855,N_16873);
and U17057 (N_17057,N_16865,N_16889);
or U17058 (N_17058,N_16836,N_16915);
and U17059 (N_17059,N_16916,N_16864);
xor U17060 (N_17060,N_16918,N_16968);
xor U17061 (N_17061,N_16885,N_16914);
and U17062 (N_17062,N_16895,N_16985);
or U17063 (N_17063,N_16990,N_16994);
nand U17064 (N_17064,N_16804,N_16894);
and U17065 (N_17065,N_16945,N_16906);
xnor U17066 (N_17066,N_16811,N_16905);
nor U17067 (N_17067,N_16890,N_16824);
xnor U17068 (N_17068,N_16946,N_16852);
nand U17069 (N_17069,N_16816,N_16832);
or U17070 (N_17070,N_16925,N_16868);
or U17071 (N_17071,N_16907,N_16981);
nand U17072 (N_17072,N_16978,N_16897);
nor U17073 (N_17073,N_16939,N_16875);
nor U17074 (N_17074,N_16854,N_16942);
nor U17075 (N_17075,N_16878,N_16952);
or U17076 (N_17076,N_16971,N_16974);
nand U17077 (N_17077,N_16828,N_16987);
or U17078 (N_17078,N_16857,N_16951);
xnor U17079 (N_17079,N_16823,N_16995);
xor U17080 (N_17080,N_16940,N_16896);
nor U17081 (N_17081,N_16869,N_16861);
and U17082 (N_17082,N_16984,N_16920);
or U17083 (N_17083,N_16829,N_16913);
xor U17084 (N_17084,N_16903,N_16835);
xor U17085 (N_17085,N_16967,N_16910);
nand U17086 (N_17086,N_16989,N_16947);
and U17087 (N_17087,N_16833,N_16966);
or U17088 (N_17088,N_16822,N_16960);
nor U17089 (N_17089,N_16956,N_16892);
or U17090 (N_17090,N_16842,N_16883);
nand U17091 (N_17091,N_16813,N_16814);
nor U17092 (N_17092,N_16936,N_16802);
xnor U17093 (N_17093,N_16998,N_16850);
nor U17094 (N_17094,N_16986,N_16973);
nand U17095 (N_17095,N_16831,N_16848);
or U17096 (N_17096,N_16902,N_16859);
or U17097 (N_17097,N_16979,N_16970);
or U17098 (N_17098,N_16847,N_16840);
xnor U17099 (N_17099,N_16874,N_16919);
and U17100 (N_17100,N_16812,N_16927);
and U17101 (N_17101,N_16871,N_16850);
and U17102 (N_17102,N_16920,N_16843);
nor U17103 (N_17103,N_16910,N_16897);
nand U17104 (N_17104,N_16975,N_16949);
and U17105 (N_17105,N_16929,N_16967);
or U17106 (N_17106,N_16914,N_16900);
nand U17107 (N_17107,N_16901,N_16876);
and U17108 (N_17108,N_16894,N_16841);
nand U17109 (N_17109,N_16855,N_16814);
and U17110 (N_17110,N_16957,N_16972);
xnor U17111 (N_17111,N_16874,N_16966);
or U17112 (N_17112,N_16816,N_16837);
nand U17113 (N_17113,N_16889,N_16819);
nor U17114 (N_17114,N_16938,N_16870);
and U17115 (N_17115,N_16971,N_16941);
or U17116 (N_17116,N_16847,N_16959);
and U17117 (N_17117,N_16846,N_16810);
nand U17118 (N_17118,N_16910,N_16832);
xor U17119 (N_17119,N_16898,N_16824);
or U17120 (N_17120,N_16825,N_16885);
nand U17121 (N_17121,N_16824,N_16869);
xor U17122 (N_17122,N_16884,N_16923);
nand U17123 (N_17123,N_16849,N_16886);
xnor U17124 (N_17124,N_16842,N_16948);
nand U17125 (N_17125,N_16911,N_16933);
or U17126 (N_17126,N_16924,N_16875);
nand U17127 (N_17127,N_16858,N_16805);
or U17128 (N_17128,N_16839,N_16893);
or U17129 (N_17129,N_16906,N_16807);
or U17130 (N_17130,N_16841,N_16947);
or U17131 (N_17131,N_16994,N_16932);
xnor U17132 (N_17132,N_16803,N_16933);
nor U17133 (N_17133,N_16900,N_16874);
and U17134 (N_17134,N_16836,N_16916);
or U17135 (N_17135,N_16821,N_16844);
and U17136 (N_17136,N_16929,N_16905);
nand U17137 (N_17137,N_16853,N_16875);
xor U17138 (N_17138,N_16860,N_16865);
and U17139 (N_17139,N_16869,N_16834);
nand U17140 (N_17140,N_16812,N_16933);
or U17141 (N_17141,N_16913,N_16948);
and U17142 (N_17142,N_16828,N_16811);
or U17143 (N_17143,N_16962,N_16844);
nor U17144 (N_17144,N_16990,N_16898);
nand U17145 (N_17145,N_16878,N_16825);
xnor U17146 (N_17146,N_16804,N_16912);
or U17147 (N_17147,N_16867,N_16861);
nand U17148 (N_17148,N_16892,N_16975);
nand U17149 (N_17149,N_16917,N_16886);
and U17150 (N_17150,N_16843,N_16971);
and U17151 (N_17151,N_16920,N_16818);
or U17152 (N_17152,N_16979,N_16902);
or U17153 (N_17153,N_16892,N_16883);
nand U17154 (N_17154,N_16927,N_16865);
and U17155 (N_17155,N_16809,N_16985);
xnor U17156 (N_17156,N_16923,N_16953);
nand U17157 (N_17157,N_16870,N_16983);
xnor U17158 (N_17158,N_16968,N_16915);
xnor U17159 (N_17159,N_16843,N_16829);
nor U17160 (N_17160,N_16815,N_16945);
nand U17161 (N_17161,N_16942,N_16977);
xor U17162 (N_17162,N_16893,N_16882);
or U17163 (N_17163,N_16829,N_16976);
and U17164 (N_17164,N_16948,N_16996);
or U17165 (N_17165,N_16962,N_16926);
or U17166 (N_17166,N_16875,N_16864);
and U17167 (N_17167,N_16866,N_16931);
and U17168 (N_17168,N_16952,N_16887);
and U17169 (N_17169,N_16991,N_16978);
nand U17170 (N_17170,N_16826,N_16898);
nor U17171 (N_17171,N_16977,N_16986);
nand U17172 (N_17172,N_16976,N_16987);
xor U17173 (N_17173,N_16839,N_16986);
nand U17174 (N_17174,N_16992,N_16847);
nor U17175 (N_17175,N_16802,N_16901);
nor U17176 (N_17176,N_16924,N_16813);
xor U17177 (N_17177,N_16966,N_16819);
and U17178 (N_17178,N_16861,N_16839);
nor U17179 (N_17179,N_16807,N_16892);
or U17180 (N_17180,N_16980,N_16869);
nor U17181 (N_17181,N_16996,N_16860);
and U17182 (N_17182,N_16953,N_16880);
or U17183 (N_17183,N_16830,N_16835);
xnor U17184 (N_17184,N_16867,N_16897);
or U17185 (N_17185,N_16926,N_16861);
xnor U17186 (N_17186,N_16920,N_16838);
xor U17187 (N_17187,N_16918,N_16809);
nand U17188 (N_17188,N_16951,N_16835);
nor U17189 (N_17189,N_16813,N_16949);
nor U17190 (N_17190,N_16857,N_16942);
or U17191 (N_17191,N_16822,N_16843);
xnor U17192 (N_17192,N_16802,N_16863);
nand U17193 (N_17193,N_16811,N_16825);
or U17194 (N_17194,N_16985,N_16830);
xor U17195 (N_17195,N_16998,N_16989);
xor U17196 (N_17196,N_16810,N_16866);
xor U17197 (N_17197,N_16910,N_16930);
xor U17198 (N_17198,N_16852,N_16942);
nor U17199 (N_17199,N_16807,N_16861);
and U17200 (N_17200,N_17068,N_17119);
nand U17201 (N_17201,N_17025,N_17121);
nand U17202 (N_17202,N_17080,N_17183);
xor U17203 (N_17203,N_17047,N_17150);
or U17204 (N_17204,N_17178,N_17075);
nor U17205 (N_17205,N_17139,N_17006);
xnor U17206 (N_17206,N_17198,N_17014);
or U17207 (N_17207,N_17083,N_17032);
and U17208 (N_17208,N_17074,N_17180);
or U17209 (N_17209,N_17060,N_17194);
nor U17210 (N_17210,N_17158,N_17107);
and U17211 (N_17211,N_17067,N_17157);
nor U17212 (N_17212,N_17069,N_17169);
nand U17213 (N_17213,N_17120,N_17004);
and U17214 (N_17214,N_17009,N_17000);
xnor U17215 (N_17215,N_17043,N_17170);
or U17216 (N_17216,N_17087,N_17077);
or U17217 (N_17217,N_17095,N_17058);
nand U17218 (N_17218,N_17114,N_17151);
and U17219 (N_17219,N_17176,N_17024);
and U17220 (N_17220,N_17090,N_17097);
and U17221 (N_17221,N_17076,N_17137);
and U17222 (N_17222,N_17131,N_17030);
nand U17223 (N_17223,N_17084,N_17044);
nor U17224 (N_17224,N_17051,N_17152);
or U17225 (N_17225,N_17191,N_17126);
or U17226 (N_17226,N_17066,N_17093);
nand U17227 (N_17227,N_17070,N_17101);
xor U17228 (N_17228,N_17181,N_17042);
xor U17229 (N_17229,N_17094,N_17096);
xnor U17230 (N_17230,N_17112,N_17011);
and U17231 (N_17231,N_17039,N_17188);
nor U17232 (N_17232,N_17111,N_17145);
xor U17233 (N_17233,N_17197,N_17018);
nand U17234 (N_17234,N_17088,N_17162);
or U17235 (N_17235,N_17186,N_17023);
or U17236 (N_17236,N_17135,N_17089);
nand U17237 (N_17237,N_17125,N_17082);
nor U17238 (N_17238,N_17050,N_17003);
nor U17239 (N_17239,N_17038,N_17061);
or U17240 (N_17240,N_17122,N_17046);
xnor U17241 (N_17241,N_17182,N_17029);
nor U17242 (N_17242,N_17179,N_17128);
nor U17243 (N_17243,N_17031,N_17173);
and U17244 (N_17244,N_17063,N_17085);
or U17245 (N_17245,N_17054,N_17037);
nand U17246 (N_17246,N_17106,N_17059);
or U17247 (N_17247,N_17146,N_17005);
or U17248 (N_17248,N_17099,N_17109);
or U17249 (N_17249,N_17091,N_17149);
or U17250 (N_17250,N_17104,N_17155);
xnor U17251 (N_17251,N_17081,N_17168);
nor U17252 (N_17252,N_17195,N_17140);
nand U17253 (N_17253,N_17098,N_17020);
nor U17254 (N_17254,N_17102,N_17172);
xor U17255 (N_17255,N_17045,N_17078);
or U17256 (N_17256,N_17123,N_17163);
xnor U17257 (N_17257,N_17138,N_17161);
nor U17258 (N_17258,N_17013,N_17144);
xor U17259 (N_17259,N_17022,N_17064);
xnor U17260 (N_17260,N_17192,N_17117);
xor U17261 (N_17261,N_17190,N_17133);
xnor U17262 (N_17262,N_17196,N_17115);
nor U17263 (N_17263,N_17164,N_17166);
nand U17264 (N_17264,N_17154,N_17021);
or U17265 (N_17265,N_17103,N_17079);
xor U17266 (N_17266,N_17015,N_17041);
and U17267 (N_17267,N_17142,N_17033);
nor U17268 (N_17268,N_17062,N_17100);
xnor U17269 (N_17269,N_17127,N_17108);
nand U17270 (N_17270,N_17027,N_17113);
nor U17271 (N_17271,N_17184,N_17086);
and U17272 (N_17272,N_17160,N_17053);
nand U17273 (N_17273,N_17028,N_17010);
xnor U17274 (N_17274,N_17136,N_17052);
xor U17275 (N_17275,N_17019,N_17057);
nand U17276 (N_17276,N_17055,N_17072);
xnor U17277 (N_17277,N_17110,N_17141);
nand U17278 (N_17278,N_17012,N_17134);
nor U17279 (N_17279,N_17049,N_17185);
nor U17280 (N_17280,N_17156,N_17092);
xnor U17281 (N_17281,N_17026,N_17171);
and U17282 (N_17282,N_17147,N_17177);
or U17283 (N_17283,N_17073,N_17153);
and U17284 (N_17284,N_17167,N_17065);
nand U17285 (N_17285,N_17199,N_17159);
nor U17286 (N_17286,N_17130,N_17189);
or U17287 (N_17287,N_17035,N_17040);
nor U17288 (N_17288,N_17034,N_17017);
nor U17289 (N_17289,N_17001,N_17132);
xnor U17290 (N_17290,N_17187,N_17129);
nand U17291 (N_17291,N_17036,N_17175);
and U17292 (N_17292,N_17193,N_17048);
or U17293 (N_17293,N_17071,N_17116);
or U17294 (N_17294,N_17016,N_17124);
nor U17295 (N_17295,N_17174,N_17118);
or U17296 (N_17296,N_17056,N_17008);
nand U17297 (N_17297,N_17007,N_17143);
or U17298 (N_17298,N_17105,N_17148);
xnor U17299 (N_17299,N_17165,N_17002);
or U17300 (N_17300,N_17197,N_17030);
xor U17301 (N_17301,N_17050,N_17042);
nand U17302 (N_17302,N_17148,N_17181);
xor U17303 (N_17303,N_17085,N_17049);
nand U17304 (N_17304,N_17019,N_17039);
nand U17305 (N_17305,N_17103,N_17194);
or U17306 (N_17306,N_17186,N_17195);
and U17307 (N_17307,N_17177,N_17115);
and U17308 (N_17308,N_17124,N_17129);
and U17309 (N_17309,N_17028,N_17123);
xor U17310 (N_17310,N_17175,N_17017);
and U17311 (N_17311,N_17113,N_17054);
nor U17312 (N_17312,N_17027,N_17017);
nand U17313 (N_17313,N_17107,N_17103);
xnor U17314 (N_17314,N_17128,N_17090);
and U17315 (N_17315,N_17071,N_17144);
xor U17316 (N_17316,N_17160,N_17039);
xnor U17317 (N_17317,N_17084,N_17186);
or U17318 (N_17318,N_17081,N_17042);
or U17319 (N_17319,N_17194,N_17170);
nand U17320 (N_17320,N_17028,N_17040);
and U17321 (N_17321,N_17056,N_17134);
xor U17322 (N_17322,N_17114,N_17047);
or U17323 (N_17323,N_17045,N_17049);
xor U17324 (N_17324,N_17107,N_17017);
and U17325 (N_17325,N_17199,N_17039);
nand U17326 (N_17326,N_17149,N_17147);
xor U17327 (N_17327,N_17039,N_17044);
xnor U17328 (N_17328,N_17195,N_17104);
or U17329 (N_17329,N_17021,N_17188);
nand U17330 (N_17330,N_17076,N_17029);
nor U17331 (N_17331,N_17147,N_17173);
and U17332 (N_17332,N_17177,N_17016);
xor U17333 (N_17333,N_17181,N_17150);
or U17334 (N_17334,N_17148,N_17053);
nand U17335 (N_17335,N_17191,N_17038);
nor U17336 (N_17336,N_17125,N_17002);
nor U17337 (N_17337,N_17058,N_17020);
nand U17338 (N_17338,N_17102,N_17107);
xnor U17339 (N_17339,N_17181,N_17097);
or U17340 (N_17340,N_17149,N_17141);
nor U17341 (N_17341,N_17026,N_17000);
nor U17342 (N_17342,N_17106,N_17130);
and U17343 (N_17343,N_17163,N_17025);
nand U17344 (N_17344,N_17192,N_17150);
nand U17345 (N_17345,N_17038,N_17025);
nand U17346 (N_17346,N_17090,N_17141);
or U17347 (N_17347,N_17191,N_17170);
xnor U17348 (N_17348,N_17126,N_17063);
and U17349 (N_17349,N_17021,N_17016);
nand U17350 (N_17350,N_17125,N_17142);
xor U17351 (N_17351,N_17064,N_17163);
and U17352 (N_17352,N_17149,N_17155);
nor U17353 (N_17353,N_17059,N_17129);
xnor U17354 (N_17354,N_17111,N_17123);
xor U17355 (N_17355,N_17007,N_17128);
and U17356 (N_17356,N_17132,N_17047);
and U17357 (N_17357,N_17131,N_17011);
xor U17358 (N_17358,N_17158,N_17070);
nand U17359 (N_17359,N_17005,N_17034);
or U17360 (N_17360,N_17042,N_17182);
xor U17361 (N_17361,N_17197,N_17147);
and U17362 (N_17362,N_17102,N_17034);
nand U17363 (N_17363,N_17072,N_17196);
and U17364 (N_17364,N_17063,N_17049);
or U17365 (N_17365,N_17163,N_17091);
and U17366 (N_17366,N_17103,N_17055);
nand U17367 (N_17367,N_17143,N_17064);
or U17368 (N_17368,N_17120,N_17193);
nand U17369 (N_17369,N_17024,N_17057);
nand U17370 (N_17370,N_17082,N_17173);
or U17371 (N_17371,N_17029,N_17192);
nand U17372 (N_17372,N_17121,N_17007);
nand U17373 (N_17373,N_17165,N_17071);
nor U17374 (N_17374,N_17033,N_17079);
nand U17375 (N_17375,N_17132,N_17006);
nand U17376 (N_17376,N_17115,N_17133);
or U17377 (N_17377,N_17070,N_17163);
or U17378 (N_17378,N_17132,N_17184);
nand U17379 (N_17379,N_17143,N_17029);
nand U17380 (N_17380,N_17017,N_17161);
or U17381 (N_17381,N_17112,N_17034);
xnor U17382 (N_17382,N_17045,N_17150);
or U17383 (N_17383,N_17188,N_17054);
xnor U17384 (N_17384,N_17194,N_17001);
nand U17385 (N_17385,N_17045,N_17118);
nor U17386 (N_17386,N_17020,N_17186);
xnor U17387 (N_17387,N_17085,N_17071);
or U17388 (N_17388,N_17015,N_17153);
xor U17389 (N_17389,N_17007,N_17131);
xnor U17390 (N_17390,N_17119,N_17171);
and U17391 (N_17391,N_17022,N_17152);
or U17392 (N_17392,N_17186,N_17160);
nor U17393 (N_17393,N_17044,N_17041);
or U17394 (N_17394,N_17183,N_17109);
xor U17395 (N_17395,N_17144,N_17079);
or U17396 (N_17396,N_17037,N_17044);
nor U17397 (N_17397,N_17090,N_17123);
and U17398 (N_17398,N_17145,N_17074);
nor U17399 (N_17399,N_17112,N_17115);
and U17400 (N_17400,N_17249,N_17274);
or U17401 (N_17401,N_17360,N_17394);
nand U17402 (N_17402,N_17257,N_17339);
xor U17403 (N_17403,N_17324,N_17327);
or U17404 (N_17404,N_17223,N_17292);
nand U17405 (N_17405,N_17233,N_17263);
xnor U17406 (N_17406,N_17241,N_17298);
nand U17407 (N_17407,N_17396,N_17310);
or U17408 (N_17408,N_17328,N_17382);
or U17409 (N_17409,N_17281,N_17242);
nor U17410 (N_17410,N_17212,N_17359);
nor U17411 (N_17411,N_17288,N_17377);
and U17412 (N_17412,N_17334,N_17203);
and U17413 (N_17413,N_17220,N_17269);
nand U17414 (N_17414,N_17368,N_17349);
xnor U17415 (N_17415,N_17306,N_17236);
xor U17416 (N_17416,N_17286,N_17283);
or U17417 (N_17417,N_17336,N_17398);
nor U17418 (N_17418,N_17227,N_17246);
nand U17419 (N_17419,N_17393,N_17322);
nor U17420 (N_17420,N_17376,N_17320);
nand U17421 (N_17421,N_17289,N_17307);
xor U17422 (N_17422,N_17399,N_17348);
xor U17423 (N_17423,N_17300,N_17226);
xnor U17424 (N_17424,N_17332,N_17346);
and U17425 (N_17425,N_17204,N_17378);
xor U17426 (N_17426,N_17273,N_17205);
nor U17427 (N_17427,N_17271,N_17369);
nand U17428 (N_17428,N_17285,N_17211);
xor U17429 (N_17429,N_17287,N_17312);
nor U17430 (N_17430,N_17279,N_17276);
nor U17431 (N_17431,N_17237,N_17352);
and U17432 (N_17432,N_17303,N_17337);
nand U17433 (N_17433,N_17383,N_17391);
and U17434 (N_17434,N_17221,N_17308);
xnor U17435 (N_17435,N_17270,N_17299);
xor U17436 (N_17436,N_17370,N_17268);
or U17437 (N_17437,N_17304,N_17341);
or U17438 (N_17438,N_17240,N_17244);
or U17439 (N_17439,N_17367,N_17228);
nand U17440 (N_17440,N_17243,N_17375);
or U17441 (N_17441,N_17296,N_17350);
and U17442 (N_17442,N_17275,N_17231);
nand U17443 (N_17443,N_17260,N_17395);
xor U17444 (N_17444,N_17372,N_17326);
xor U17445 (N_17445,N_17208,N_17254);
or U17446 (N_17446,N_17250,N_17389);
xnor U17447 (N_17447,N_17361,N_17363);
xor U17448 (N_17448,N_17305,N_17261);
or U17449 (N_17449,N_17329,N_17293);
xor U17450 (N_17450,N_17245,N_17338);
nor U17451 (N_17451,N_17239,N_17319);
nor U17452 (N_17452,N_17309,N_17219);
xor U17453 (N_17453,N_17282,N_17222);
or U17454 (N_17454,N_17247,N_17225);
nand U17455 (N_17455,N_17330,N_17371);
nand U17456 (N_17456,N_17272,N_17277);
nand U17457 (N_17457,N_17294,N_17355);
nor U17458 (N_17458,N_17387,N_17342);
xnor U17459 (N_17459,N_17267,N_17258);
and U17460 (N_17460,N_17278,N_17366);
nand U17461 (N_17461,N_17206,N_17200);
nor U17462 (N_17462,N_17214,N_17333);
and U17463 (N_17463,N_17207,N_17262);
xor U17464 (N_17464,N_17216,N_17215);
nor U17465 (N_17465,N_17290,N_17256);
or U17466 (N_17466,N_17253,N_17344);
and U17467 (N_17467,N_17291,N_17255);
nand U17468 (N_17468,N_17316,N_17248);
or U17469 (N_17469,N_17362,N_17374);
nand U17470 (N_17470,N_17259,N_17357);
or U17471 (N_17471,N_17210,N_17252);
or U17472 (N_17472,N_17284,N_17392);
nand U17473 (N_17473,N_17217,N_17295);
nand U17474 (N_17474,N_17354,N_17345);
nor U17475 (N_17475,N_17302,N_17384);
nor U17476 (N_17476,N_17358,N_17265);
nor U17477 (N_17477,N_17238,N_17314);
nor U17478 (N_17478,N_17325,N_17317);
xnor U17479 (N_17479,N_17251,N_17340);
xor U17480 (N_17480,N_17380,N_17311);
nor U17481 (N_17481,N_17335,N_17356);
nand U17482 (N_17482,N_17202,N_17321);
nand U17483 (N_17483,N_17385,N_17213);
or U17484 (N_17484,N_17364,N_17315);
nor U17485 (N_17485,N_17301,N_17201);
and U17486 (N_17486,N_17234,N_17230);
or U17487 (N_17487,N_17229,N_17343);
xnor U17488 (N_17488,N_17351,N_17347);
nor U17489 (N_17489,N_17390,N_17224);
or U17490 (N_17490,N_17381,N_17397);
nand U17491 (N_17491,N_17388,N_17297);
or U17492 (N_17492,N_17353,N_17264);
or U17493 (N_17493,N_17266,N_17318);
and U17494 (N_17494,N_17232,N_17331);
or U17495 (N_17495,N_17209,N_17313);
or U17496 (N_17496,N_17379,N_17373);
nand U17497 (N_17497,N_17280,N_17365);
xor U17498 (N_17498,N_17235,N_17218);
or U17499 (N_17499,N_17386,N_17323);
or U17500 (N_17500,N_17207,N_17274);
or U17501 (N_17501,N_17331,N_17297);
xnor U17502 (N_17502,N_17268,N_17382);
nand U17503 (N_17503,N_17319,N_17225);
nor U17504 (N_17504,N_17361,N_17358);
nor U17505 (N_17505,N_17381,N_17263);
nor U17506 (N_17506,N_17232,N_17286);
or U17507 (N_17507,N_17390,N_17288);
nand U17508 (N_17508,N_17348,N_17397);
xnor U17509 (N_17509,N_17353,N_17218);
nand U17510 (N_17510,N_17285,N_17392);
nand U17511 (N_17511,N_17212,N_17343);
or U17512 (N_17512,N_17264,N_17388);
nand U17513 (N_17513,N_17310,N_17329);
nand U17514 (N_17514,N_17381,N_17313);
xnor U17515 (N_17515,N_17284,N_17215);
and U17516 (N_17516,N_17387,N_17222);
nand U17517 (N_17517,N_17393,N_17268);
and U17518 (N_17518,N_17394,N_17236);
nor U17519 (N_17519,N_17309,N_17209);
xor U17520 (N_17520,N_17286,N_17260);
and U17521 (N_17521,N_17323,N_17279);
nor U17522 (N_17522,N_17249,N_17202);
xor U17523 (N_17523,N_17292,N_17262);
or U17524 (N_17524,N_17344,N_17349);
or U17525 (N_17525,N_17362,N_17355);
nand U17526 (N_17526,N_17389,N_17281);
or U17527 (N_17527,N_17352,N_17335);
or U17528 (N_17528,N_17228,N_17284);
or U17529 (N_17529,N_17226,N_17249);
and U17530 (N_17530,N_17283,N_17333);
nand U17531 (N_17531,N_17239,N_17292);
nor U17532 (N_17532,N_17397,N_17242);
nand U17533 (N_17533,N_17200,N_17341);
or U17534 (N_17534,N_17313,N_17330);
and U17535 (N_17535,N_17279,N_17268);
or U17536 (N_17536,N_17328,N_17248);
nand U17537 (N_17537,N_17237,N_17362);
nand U17538 (N_17538,N_17269,N_17305);
nor U17539 (N_17539,N_17360,N_17270);
nand U17540 (N_17540,N_17271,N_17220);
xnor U17541 (N_17541,N_17368,N_17219);
xnor U17542 (N_17542,N_17399,N_17381);
and U17543 (N_17543,N_17261,N_17257);
nor U17544 (N_17544,N_17338,N_17351);
xor U17545 (N_17545,N_17222,N_17326);
xnor U17546 (N_17546,N_17236,N_17224);
or U17547 (N_17547,N_17371,N_17290);
or U17548 (N_17548,N_17398,N_17312);
and U17549 (N_17549,N_17393,N_17360);
xor U17550 (N_17550,N_17340,N_17372);
nor U17551 (N_17551,N_17284,N_17240);
nand U17552 (N_17552,N_17356,N_17310);
xor U17553 (N_17553,N_17210,N_17373);
and U17554 (N_17554,N_17247,N_17220);
xor U17555 (N_17555,N_17384,N_17376);
or U17556 (N_17556,N_17340,N_17222);
xnor U17557 (N_17557,N_17384,N_17252);
and U17558 (N_17558,N_17271,N_17371);
nand U17559 (N_17559,N_17311,N_17367);
nor U17560 (N_17560,N_17368,N_17318);
and U17561 (N_17561,N_17374,N_17223);
nand U17562 (N_17562,N_17318,N_17200);
and U17563 (N_17563,N_17256,N_17303);
or U17564 (N_17564,N_17388,N_17344);
nand U17565 (N_17565,N_17320,N_17253);
xor U17566 (N_17566,N_17274,N_17359);
or U17567 (N_17567,N_17278,N_17334);
nor U17568 (N_17568,N_17397,N_17340);
xor U17569 (N_17569,N_17272,N_17343);
nand U17570 (N_17570,N_17395,N_17380);
and U17571 (N_17571,N_17296,N_17258);
or U17572 (N_17572,N_17276,N_17345);
and U17573 (N_17573,N_17357,N_17339);
nor U17574 (N_17574,N_17266,N_17295);
and U17575 (N_17575,N_17251,N_17342);
nand U17576 (N_17576,N_17350,N_17309);
and U17577 (N_17577,N_17360,N_17233);
and U17578 (N_17578,N_17361,N_17353);
nor U17579 (N_17579,N_17387,N_17376);
nand U17580 (N_17580,N_17270,N_17366);
or U17581 (N_17581,N_17361,N_17327);
nor U17582 (N_17582,N_17349,N_17379);
xnor U17583 (N_17583,N_17246,N_17387);
or U17584 (N_17584,N_17216,N_17232);
or U17585 (N_17585,N_17264,N_17375);
nand U17586 (N_17586,N_17297,N_17360);
and U17587 (N_17587,N_17337,N_17383);
and U17588 (N_17588,N_17279,N_17240);
nand U17589 (N_17589,N_17325,N_17212);
nand U17590 (N_17590,N_17200,N_17399);
or U17591 (N_17591,N_17223,N_17313);
or U17592 (N_17592,N_17258,N_17298);
and U17593 (N_17593,N_17255,N_17298);
xnor U17594 (N_17594,N_17241,N_17234);
or U17595 (N_17595,N_17249,N_17304);
xor U17596 (N_17596,N_17288,N_17336);
or U17597 (N_17597,N_17301,N_17292);
or U17598 (N_17598,N_17392,N_17247);
nor U17599 (N_17599,N_17232,N_17246);
and U17600 (N_17600,N_17577,N_17512);
and U17601 (N_17601,N_17539,N_17593);
or U17602 (N_17602,N_17400,N_17487);
nand U17603 (N_17603,N_17588,N_17420);
nand U17604 (N_17604,N_17482,N_17538);
or U17605 (N_17605,N_17528,N_17424);
xor U17606 (N_17606,N_17573,N_17566);
or U17607 (N_17607,N_17550,N_17432);
or U17608 (N_17608,N_17513,N_17497);
nand U17609 (N_17609,N_17584,N_17509);
xor U17610 (N_17610,N_17471,N_17439);
xnor U17611 (N_17611,N_17426,N_17418);
nor U17612 (N_17612,N_17403,N_17430);
nor U17613 (N_17613,N_17543,N_17540);
xnor U17614 (N_17614,N_17570,N_17425);
or U17615 (N_17615,N_17536,N_17559);
and U17616 (N_17616,N_17500,N_17477);
nand U17617 (N_17617,N_17555,N_17459);
nand U17618 (N_17618,N_17547,N_17561);
xor U17619 (N_17619,N_17575,N_17467);
nand U17620 (N_17620,N_17413,N_17484);
and U17621 (N_17621,N_17414,N_17522);
or U17622 (N_17622,N_17526,N_17438);
and U17623 (N_17623,N_17565,N_17409);
nor U17624 (N_17624,N_17450,N_17502);
nand U17625 (N_17625,N_17456,N_17419);
and U17626 (N_17626,N_17521,N_17533);
and U17627 (N_17627,N_17589,N_17415);
or U17628 (N_17628,N_17595,N_17537);
nor U17629 (N_17629,N_17583,N_17520);
or U17630 (N_17630,N_17435,N_17428);
xnor U17631 (N_17631,N_17407,N_17597);
or U17632 (N_17632,N_17452,N_17529);
nand U17633 (N_17633,N_17591,N_17581);
nor U17634 (N_17634,N_17544,N_17569);
xnor U17635 (N_17635,N_17493,N_17551);
or U17636 (N_17636,N_17486,N_17571);
nand U17637 (N_17637,N_17451,N_17574);
xnor U17638 (N_17638,N_17417,N_17401);
nand U17639 (N_17639,N_17485,N_17492);
or U17640 (N_17640,N_17563,N_17423);
and U17641 (N_17641,N_17434,N_17542);
or U17642 (N_17642,N_17444,N_17476);
nand U17643 (N_17643,N_17554,N_17576);
xor U17644 (N_17644,N_17488,N_17516);
xnor U17645 (N_17645,N_17599,N_17412);
xnor U17646 (N_17646,N_17578,N_17436);
and U17647 (N_17647,N_17553,N_17532);
and U17648 (N_17648,N_17556,N_17515);
nor U17649 (N_17649,N_17530,N_17442);
nor U17650 (N_17650,N_17489,N_17470);
nand U17651 (N_17651,N_17525,N_17534);
nand U17652 (N_17652,N_17552,N_17511);
xor U17653 (N_17653,N_17504,N_17546);
nor U17654 (N_17654,N_17572,N_17491);
and U17655 (N_17655,N_17545,N_17455);
xor U17656 (N_17656,N_17466,N_17524);
nor U17657 (N_17657,N_17454,N_17498);
xor U17658 (N_17658,N_17568,N_17519);
or U17659 (N_17659,N_17445,N_17411);
or U17660 (N_17660,N_17427,N_17523);
xnor U17661 (N_17661,N_17429,N_17587);
or U17662 (N_17662,N_17469,N_17505);
or U17663 (N_17663,N_17480,N_17433);
and U17664 (N_17664,N_17478,N_17517);
or U17665 (N_17665,N_17594,N_17503);
xor U17666 (N_17666,N_17507,N_17541);
xor U17667 (N_17667,N_17453,N_17490);
nand U17668 (N_17668,N_17531,N_17585);
and U17669 (N_17669,N_17548,N_17592);
and U17670 (N_17670,N_17441,N_17475);
or U17671 (N_17671,N_17481,N_17580);
and U17672 (N_17672,N_17549,N_17458);
or U17673 (N_17673,N_17447,N_17464);
and U17674 (N_17674,N_17495,N_17405);
xnor U17675 (N_17675,N_17461,N_17462);
xor U17676 (N_17676,N_17416,N_17527);
nor U17677 (N_17677,N_17590,N_17518);
xor U17678 (N_17678,N_17479,N_17473);
and U17679 (N_17679,N_17472,N_17474);
and U17680 (N_17680,N_17586,N_17510);
xor U17681 (N_17681,N_17449,N_17567);
nor U17682 (N_17682,N_17494,N_17468);
xnor U17683 (N_17683,N_17562,N_17483);
nor U17684 (N_17684,N_17460,N_17506);
or U17685 (N_17685,N_17446,N_17579);
nor U17686 (N_17686,N_17422,N_17501);
and U17687 (N_17687,N_17402,N_17421);
and U17688 (N_17688,N_17465,N_17437);
or U17689 (N_17689,N_17560,N_17404);
xnor U17690 (N_17690,N_17557,N_17596);
nor U17691 (N_17691,N_17496,N_17406);
nor U17692 (N_17692,N_17463,N_17410);
xnor U17693 (N_17693,N_17408,N_17448);
xor U17694 (N_17694,N_17558,N_17440);
nor U17695 (N_17695,N_17443,N_17431);
nor U17696 (N_17696,N_17514,N_17535);
nor U17697 (N_17697,N_17582,N_17499);
or U17698 (N_17698,N_17564,N_17598);
and U17699 (N_17699,N_17457,N_17508);
nand U17700 (N_17700,N_17484,N_17456);
or U17701 (N_17701,N_17550,N_17584);
nor U17702 (N_17702,N_17472,N_17521);
xor U17703 (N_17703,N_17513,N_17485);
xnor U17704 (N_17704,N_17418,N_17590);
nand U17705 (N_17705,N_17438,N_17518);
xor U17706 (N_17706,N_17539,N_17512);
nand U17707 (N_17707,N_17546,N_17473);
nand U17708 (N_17708,N_17517,N_17432);
and U17709 (N_17709,N_17523,N_17503);
and U17710 (N_17710,N_17483,N_17444);
xor U17711 (N_17711,N_17491,N_17593);
xnor U17712 (N_17712,N_17591,N_17505);
nor U17713 (N_17713,N_17439,N_17464);
nor U17714 (N_17714,N_17417,N_17434);
and U17715 (N_17715,N_17430,N_17528);
and U17716 (N_17716,N_17445,N_17478);
or U17717 (N_17717,N_17511,N_17582);
xnor U17718 (N_17718,N_17474,N_17535);
nor U17719 (N_17719,N_17448,N_17543);
nor U17720 (N_17720,N_17467,N_17587);
xnor U17721 (N_17721,N_17484,N_17538);
nor U17722 (N_17722,N_17582,N_17589);
nand U17723 (N_17723,N_17493,N_17499);
and U17724 (N_17724,N_17531,N_17509);
nand U17725 (N_17725,N_17526,N_17571);
or U17726 (N_17726,N_17497,N_17401);
or U17727 (N_17727,N_17477,N_17486);
nand U17728 (N_17728,N_17404,N_17555);
or U17729 (N_17729,N_17552,N_17483);
or U17730 (N_17730,N_17535,N_17575);
xnor U17731 (N_17731,N_17598,N_17463);
xnor U17732 (N_17732,N_17518,N_17406);
and U17733 (N_17733,N_17400,N_17545);
nor U17734 (N_17734,N_17496,N_17586);
nor U17735 (N_17735,N_17402,N_17526);
and U17736 (N_17736,N_17492,N_17574);
or U17737 (N_17737,N_17440,N_17529);
and U17738 (N_17738,N_17525,N_17449);
or U17739 (N_17739,N_17572,N_17518);
and U17740 (N_17740,N_17543,N_17441);
nand U17741 (N_17741,N_17567,N_17566);
nor U17742 (N_17742,N_17464,N_17413);
or U17743 (N_17743,N_17487,N_17419);
xor U17744 (N_17744,N_17598,N_17556);
nor U17745 (N_17745,N_17510,N_17450);
xnor U17746 (N_17746,N_17540,N_17574);
nand U17747 (N_17747,N_17574,N_17482);
or U17748 (N_17748,N_17558,N_17414);
xnor U17749 (N_17749,N_17408,N_17595);
nor U17750 (N_17750,N_17528,N_17519);
or U17751 (N_17751,N_17588,N_17419);
nor U17752 (N_17752,N_17409,N_17547);
xnor U17753 (N_17753,N_17407,N_17564);
or U17754 (N_17754,N_17411,N_17487);
nand U17755 (N_17755,N_17472,N_17452);
nor U17756 (N_17756,N_17532,N_17507);
nor U17757 (N_17757,N_17510,N_17568);
nand U17758 (N_17758,N_17442,N_17419);
xnor U17759 (N_17759,N_17488,N_17458);
xor U17760 (N_17760,N_17557,N_17476);
xnor U17761 (N_17761,N_17549,N_17597);
and U17762 (N_17762,N_17464,N_17404);
nand U17763 (N_17763,N_17423,N_17446);
nor U17764 (N_17764,N_17592,N_17482);
nand U17765 (N_17765,N_17447,N_17480);
and U17766 (N_17766,N_17470,N_17590);
xor U17767 (N_17767,N_17464,N_17528);
nand U17768 (N_17768,N_17436,N_17588);
or U17769 (N_17769,N_17436,N_17521);
nand U17770 (N_17770,N_17535,N_17479);
or U17771 (N_17771,N_17500,N_17434);
and U17772 (N_17772,N_17592,N_17479);
xnor U17773 (N_17773,N_17556,N_17444);
nor U17774 (N_17774,N_17565,N_17576);
or U17775 (N_17775,N_17457,N_17431);
or U17776 (N_17776,N_17455,N_17449);
nand U17777 (N_17777,N_17504,N_17521);
nand U17778 (N_17778,N_17559,N_17586);
or U17779 (N_17779,N_17462,N_17558);
nor U17780 (N_17780,N_17416,N_17589);
nor U17781 (N_17781,N_17484,N_17501);
xnor U17782 (N_17782,N_17552,N_17453);
nand U17783 (N_17783,N_17443,N_17471);
nor U17784 (N_17784,N_17500,N_17528);
nor U17785 (N_17785,N_17466,N_17510);
xor U17786 (N_17786,N_17466,N_17548);
and U17787 (N_17787,N_17553,N_17531);
or U17788 (N_17788,N_17419,N_17413);
nand U17789 (N_17789,N_17509,N_17523);
and U17790 (N_17790,N_17413,N_17449);
xor U17791 (N_17791,N_17484,N_17553);
nand U17792 (N_17792,N_17402,N_17472);
or U17793 (N_17793,N_17426,N_17513);
nor U17794 (N_17794,N_17568,N_17515);
nand U17795 (N_17795,N_17543,N_17425);
xor U17796 (N_17796,N_17421,N_17478);
or U17797 (N_17797,N_17415,N_17437);
xnor U17798 (N_17798,N_17565,N_17411);
nor U17799 (N_17799,N_17580,N_17414);
nor U17800 (N_17800,N_17717,N_17751);
or U17801 (N_17801,N_17694,N_17681);
and U17802 (N_17802,N_17711,N_17773);
xor U17803 (N_17803,N_17658,N_17649);
and U17804 (N_17804,N_17612,N_17767);
and U17805 (N_17805,N_17660,N_17616);
or U17806 (N_17806,N_17732,N_17781);
and U17807 (N_17807,N_17666,N_17742);
and U17808 (N_17808,N_17684,N_17662);
nand U17809 (N_17809,N_17644,N_17623);
xor U17810 (N_17810,N_17776,N_17606);
xnor U17811 (N_17811,N_17611,N_17796);
and U17812 (N_17812,N_17746,N_17687);
and U17813 (N_17813,N_17697,N_17638);
nand U17814 (N_17814,N_17688,N_17772);
nand U17815 (N_17815,N_17693,N_17710);
or U17816 (N_17816,N_17620,N_17603);
nor U17817 (N_17817,N_17700,N_17625);
nor U17818 (N_17818,N_17723,N_17769);
xnor U17819 (N_17819,N_17613,N_17738);
nand U17820 (N_17820,N_17601,N_17736);
nor U17821 (N_17821,N_17709,N_17741);
and U17822 (N_17822,N_17698,N_17793);
xnor U17823 (N_17823,N_17798,N_17701);
or U17824 (N_17824,N_17725,N_17626);
or U17825 (N_17825,N_17654,N_17784);
nand U17826 (N_17826,N_17756,N_17750);
nand U17827 (N_17827,N_17627,N_17682);
or U17828 (N_17828,N_17633,N_17743);
nor U17829 (N_17829,N_17788,N_17739);
or U17830 (N_17830,N_17735,N_17777);
and U17831 (N_17831,N_17770,N_17721);
or U17832 (N_17832,N_17669,N_17640);
xor U17833 (N_17833,N_17631,N_17624);
nor U17834 (N_17834,N_17794,N_17636);
xor U17835 (N_17835,N_17643,N_17671);
and U17836 (N_17836,N_17729,N_17650);
nor U17837 (N_17837,N_17705,N_17622);
nand U17838 (N_17838,N_17747,N_17665);
or U17839 (N_17839,N_17653,N_17674);
nor U17840 (N_17840,N_17608,N_17761);
and U17841 (N_17841,N_17706,N_17628);
and U17842 (N_17842,N_17621,N_17629);
nand U17843 (N_17843,N_17605,N_17791);
nand U17844 (N_17844,N_17672,N_17648);
or U17845 (N_17845,N_17778,N_17785);
nand U17846 (N_17846,N_17749,N_17673);
xor U17847 (N_17847,N_17779,N_17600);
or U17848 (N_17848,N_17783,N_17617);
or U17849 (N_17849,N_17782,N_17632);
nor U17850 (N_17850,N_17766,N_17609);
or U17851 (N_17851,N_17753,N_17795);
or U17852 (N_17852,N_17680,N_17716);
and U17853 (N_17853,N_17760,N_17696);
or U17854 (N_17854,N_17790,N_17733);
or U17855 (N_17855,N_17659,N_17663);
nand U17856 (N_17856,N_17708,N_17651);
xnor U17857 (N_17857,N_17780,N_17762);
xnor U17858 (N_17858,N_17685,N_17792);
xor U17859 (N_17859,N_17731,N_17752);
xnor U17860 (N_17860,N_17754,N_17763);
or U17861 (N_17861,N_17677,N_17724);
nand U17862 (N_17862,N_17690,N_17695);
or U17863 (N_17863,N_17657,N_17703);
and U17864 (N_17864,N_17730,N_17775);
nand U17865 (N_17865,N_17789,N_17728);
nor U17866 (N_17866,N_17699,N_17758);
and U17867 (N_17867,N_17635,N_17604);
and U17868 (N_17868,N_17734,N_17757);
nor U17869 (N_17869,N_17718,N_17707);
xnor U17870 (N_17870,N_17615,N_17704);
nor U17871 (N_17871,N_17737,N_17686);
xor U17872 (N_17872,N_17661,N_17676);
nor U17873 (N_17873,N_17712,N_17655);
nor U17874 (N_17874,N_17765,N_17774);
nand U17875 (N_17875,N_17637,N_17713);
or U17876 (N_17876,N_17646,N_17744);
or U17877 (N_17877,N_17664,N_17759);
and U17878 (N_17878,N_17787,N_17797);
nor U17879 (N_17879,N_17642,N_17726);
or U17880 (N_17880,N_17748,N_17667);
nand U17881 (N_17881,N_17675,N_17764);
or U17882 (N_17882,N_17740,N_17692);
nor U17883 (N_17883,N_17745,N_17645);
or U17884 (N_17884,N_17727,N_17607);
xnor U17885 (N_17885,N_17602,N_17639);
nand U17886 (N_17886,N_17768,N_17668);
nand U17887 (N_17887,N_17610,N_17619);
nand U17888 (N_17888,N_17715,N_17634);
and U17889 (N_17889,N_17618,N_17630);
nand U17890 (N_17890,N_17786,N_17683);
and U17891 (N_17891,N_17678,N_17652);
xor U17892 (N_17892,N_17720,N_17719);
nand U17893 (N_17893,N_17722,N_17691);
xnor U17894 (N_17894,N_17647,N_17641);
and U17895 (N_17895,N_17656,N_17670);
and U17896 (N_17896,N_17799,N_17689);
xor U17897 (N_17897,N_17755,N_17614);
and U17898 (N_17898,N_17679,N_17714);
nor U17899 (N_17899,N_17771,N_17702);
xor U17900 (N_17900,N_17754,N_17665);
and U17901 (N_17901,N_17628,N_17605);
nor U17902 (N_17902,N_17638,N_17643);
or U17903 (N_17903,N_17655,N_17745);
and U17904 (N_17904,N_17713,N_17658);
and U17905 (N_17905,N_17659,N_17613);
and U17906 (N_17906,N_17624,N_17745);
or U17907 (N_17907,N_17609,N_17781);
and U17908 (N_17908,N_17650,N_17618);
or U17909 (N_17909,N_17775,N_17683);
nand U17910 (N_17910,N_17703,N_17740);
or U17911 (N_17911,N_17607,N_17745);
nor U17912 (N_17912,N_17633,N_17754);
nor U17913 (N_17913,N_17793,N_17663);
nand U17914 (N_17914,N_17766,N_17791);
nor U17915 (N_17915,N_17791,N_17684);
nand U17916 (N_17916,N_17772,N_17639);
nand U17917 (N_17917,N_17780,N_17794);
nor U17918 (N_17918,N_17706,N_17666);
or U17919 (N_17919,N_17629,N_17608);
xor U17920 (N_17920,N_17663,N_17788);
or U17921 (N_17921,N_17717,N_17655);
nand U17922 (N_17922,N_17604,N_17752);
and U17923 (N_17923,N_17681,N_17658);
xnor U17924 (N_17924,N_17741,N_17785);
xnor U17925 (N_17925,N_17624,N_17795);
xnor U17926 (N_17926,N_17778,N_17678);
nor U17927 (N_17927,N_17618,N_17778);
and U17928 (N_17928,N_17623,N_17742);
xor U17929 (N_17929,N_17706,N_17774);
nand U17930 (N_17930,N_17792,N_17626);
and U17931 (N_17931,N_17662,N_17638);
and U17932 (N_17932,N_17761,N_17726);
xnor U17933 (N_17933,N_17616,N_17780);
nand U17934 (N_17934,N_17678,N_17659);
and U17935 (N_17935,N_17725,N_17622);
xor U17936 (N_17936,N_17650,N_17737);
xnor U17937 (N_17937,N_17769,N_17782);
and U17938 (N_17938,N_17695,N_17622);
nand U17939 (N_17939,N_17654,N_17645);
and U17940 (N_17940,N_17791,N_17721);
or U17941 (N_17941,N_17632,N_17735);
or U17942 (N_17942,N_17614,N_17729);
nand U17943 (N_17943,N_17660,N_17745);
nor U17944 (N_17944,N_17697,N_17618);
xor U17945 (N_17945,N_17685,N_17656);
nor U17946 (N_17946,N_17750,N_17698);
nand U17947 (N_17947,N_17773,N_17658);
xnor U17948 (N_17948,N_17796,N_17786);
and U17949 (N_17949,N_17733,N_17722);
xnor U17950 (N_17950,N_17648,N_17608);
xor U17951 (N_17951,N_17675,N_17622);
and U17952 (N_17952,N_17639,N_17744);
xnor U17953 (N_17953,N_17652,N_17619);
and U17954 (N_17954,N_17780,N_17680);
nor U17955 (N_17955,N_17721,N_17753);
and U17956 (N_17956,N_17721,N_17754);
or U17957 (N_17957,N_17676,N_17614);
and U17958 (N_17958,N_17651,N_17791);
or U17959 (N_17959,N_17607,N_17660);
and U17960 (N_17960,N_17670,N_17761);
and U17961 (N_17961,N_17671,N_17672);
xnor U17962 (N_17962,N_17631,N_17792);
nand U17963 (N_17963,N_17695,N_17777);
nor U17964 (N_17964,N_17730,N_17788);
nor U17965 (N_17965,N_17639,N_17664);
xor U17966 (N_17966,N_17696,N_17759);
nand U17967 (N_17967,N_17658,N_17745);
xor U17968 (N_17968,N_17655,N_17635);
nand U17969 (N_17969,N_17718,N_17763);
nand U17970 (N_17970,N_17794,N_17765);
xnor U17971 (N_17971,N_17618,N_17684);
xor U17972 (N_17972,N_17686,N_17740);
or U17973 (N_17973,N_17673,N_17674);
and U17974 (N_17974,N_17605,N_17633);
nand U17975 (N_17975,N_17773,N_17707);
xor U17976 (N_17976,N_17614,N_17638);
nor U17977 (N_17977,N_17639,N_17661);
or U17978 (N_17978,N_17630,N_17666);
nand U17979 (N_17979,N_17720,N_17737);
or U17980 (N_17980,N_17739,N_17640);
or U17981 (N_17981,N_17627,N_17671);
nand U17982 (N_17982,N_17741,N_17664);
nand U17983 (N_17983,N_17635,N_17725);
and U17984 (N_17984,N_17649,N_17777);
nand U17985 (N_17985,N_17736,N_17798);
xnor U17986 (N_17986,N_17649,N_17783);
nand U17987 (N_17987,N_17750,N_17727);
xnor U17988 (N_17988,N_17630,N_17726);
nor U17989 (N_17989,N_17773,N_17751);
nor U17990 (N_17990,N_17729,N_17682);
and U17991 (N_17991,N_17740,N_17603);
nand U17992 (N_17992,N_17781,N_17731);
xor U17993 (N_17993,N_17606,N_17670);
and U17994 (N_17994,N_17744,N_17608);
nor U17995 (N_17995,N_17752,N_17602);
nand U17996 (N_17996,N_17769,N_17736);
xnor U17997 (N_17997,N_17731,N_17612);
or U17998 (N_17998,N_17636,N_17708);
nor U17999 (N_17999,N_17632,N_17655);
nand U18000 (N_18000,N_17869,N_17854);
nand U18001 (N_18001,N_17977,N_17898);
and U18002 (N_18002,N_17983,N_17973);
nand U18003 (N_18003,N_17816,N_17950);
and U18004 (N_18004,N_17890,N_17953);
xnor U18005 (N_18005,N_17864,N_17955);
nand U18006 (N_18006,N_17928,N_17995);
nor U18007 (N_18007,N_17989,N_17954);
nor U18008 (N_18008,N_17951,N_17982);
nand U18009 (N_18009,N_17978,N_17812);
xnor U18010 (N_18010,N_17968,N_17979);
nor U18011 (N_18011,N_17847,N_17845);
and U18012 (N_18012,N_17827,N_17932);
and U18013 (N_18013,N_17834,N_17937);
xnor U18014 (N_18014,N_17856,N_17859);
and U18015 (N_18015,N_17824,N_17835);
xnor U18016 (N_18016,N_17842,N_17878);
or U18017 (N_18017,N_17942,N_17922);
nor U18018 (N_18018,N_17974,N_17930);
nor U18019 (N_18019,N_17870,N_17844);
xnor U18020 (N_18020,N_17855,N_17881);
nor U18021 (N_18021,N_17993,N_17825);
nor U18022 (N_18022,N_17829,N_17908);
or U18023 (N_18023,N_17944,N_17947);
nor U18024 (N_18024,N_17998,N_17970);
xnor U18025 (N_18025,N_17868,N_17963);
xor U18026 (N_18026,N_17888,N_17893);
or U18027 (N_18027,N_17985,N_17902);
or U18028 (N_18028,N_17894,N_17860);
and U18029 (N_18029,N_17988,N_17931);
or U18030 (N_18030,N_17990,N_17965);
and U18031 (N_18031,N_17806,N_17866);
and U18032 (N_18032,N_17895,N_17933);
xnor U18033 (N_18033,N_17921,N_17846);
xnor U18034 (N_18034,N_17850,N_17882);
xnor U18035 (N_18035,N_17958,N_17927);
and U18036 (N_18036,N_17873,N_17964);
and U18037 (N_18037,N_17828,N_17897);
and U18038 (N_18038,N_17929,N_17956);
and U18039 (N_18039,N_17826,N_17948);
and U18040 (N_18040,N_17971,N_17906);
nor U18041 (N_18041,N_17991,N_17848);
and U18042 (N_18042,N_17841,N_17858);
nand U18043 (N_18043,N_17884,N_17849);
nand U18044 (N_18044,N_17838,N_17885);
xnor U18045 (N_18045,N_17853,N_17851);
xor U18046 (N_18046,N_17913,N_17810);
nand U18047 (N_18047,N_17821,N_17960);
and U18048 (N_18048,N_17814,N_17802);
nand U18049 (N_18049,N_17889,N_17915);
nor U18050 (N_18050,N_17803,N_17938);
nand U18051 (N_18051,N_17952,N_17962);
nand U18052 (N_18052,N_17975,N_17904);
and U18053 (N_18053,N_17926,N_17874);
nor U18054 (N_18054,N_17986,N_17976);
nor U18055 (N_18055,N_17905,N_17833);
or U18056 (N_18056,N_17839,N_17832);
or U18057 (N_18057,N_17949,N_17867);
nand U18058 (N_18058,N_17823,N_17901);
and U18059 (N_18059,N_17923,N_17910);
nand U18060 (N_18060,N_17843,N_17831);
and U18061 (N_18061,N_17883,N_17992);
nand U18062 (N_18062,N_17903,N_17822);
or U18063 (N_18063,N_17801,N_17875);
and U18064 (N_18064,N_17877,N_17961);
or U18065 (N_18065,N_17994,N_17946);
and U18066 (N_18066,N_17813,N_17861);
nor U18067 (N_18067,N_17836,N_17886);
or U18068 (N_18068,N_17916,N_17857);
or U18069 (N_18069,N_17809,N_17997);
xnor U18070 (N_18070,N_17969,N_17815);
xor U18071 (N_18071,N_17917,N_17872);
nor U18072 (N_18072,N_17880,N_17966);
xor U18073 (N_18073,N_17805,N_17936);
and U18074 (N_18074,N_17911,N_17876);
xnor U18075 (N_18075,N_17808,N_17943);
and U18076 (N_18076,N_17879,N_17818);
and U18077 (N_18077,N_17996,N_17924);
nor U18078 (N_18078,N_17934,N_17941);
and U18079 (N_18079,N_17800,N_17837);
and U18080 (N_18080,N_17984,N_17980);
and U18081 (N_18081,N_17811,N_17900);
or U18082 (N_18082,N_17840,N_17871);
nand U18083 (N_18083,N_17999,N_17957);
and U18084 (N_18084,N_17891,N_17887);
or U18085 (N_18085,N_17967,N_17863);
nor U18086 (N_18086,N_17804,N_17945);
and U18087 (N_18087,N_17959,N_17865);
xor U18088 (N_18088,N_17892,N_17939);
or U18089 (N_18089,N_17920,N_17817);
nor U18090 (N_18090,N_17909,N_17918);
or U18091 (N_18091,N_17940,N_17935);
nor U18092 (N_18092,N_17896,N_17830);
or U18093 (N_18093,N_17972,N_17919);
or U18094 (N_18094,N_17987,N_17899);
nand U18095 (N_18095,N_17907,N_17981);
or U18096 (N_18096,N_17925,N_17914);
nand U18097 (N_18097,N_17862,N_17852);
or U18098 (N_18098,N_17820,N_17807);
nor U18099 (N_18099,N_17912,N_17819);
nor U18100 (N_18100,N_17891,N_17883);
and U18101 (N_18101,N_17970,N_17950);
nor U18102 (N_18102,N_17883,N_17994);
xnor U18103 (N_18103,N_17842,N_17800);
xor U18104 (N_18104,N_17975,N_17955);
and U18105 (N_18105,N_17925,N_17800);
xnor U18106 (N_18106,N_17892,N_17910);
nor U18107 (N_18107,N_17842,N_17860);
or U18108 (N_18108,N_17834,N_17855);
nand U18109 (N_18109,N_17833,N_17880);
nand U18110 (N_18110,N_17978,N_17863);
or U18111 (N_18111,N_17887,N_17801);
and U18112 (N_18112,N_17908,N_17904);
xor U18113 (N_18113,N_17987,N_17974);
or U18114 (N_18114,N_17890,N_17934);
and U18115 (N_18115,N_17932,N_17829);
or U18116 (N_18116,N_17976,N_17980);
nand U18117 (N_18117,N_17873,N_17972);
and U18118 (N_18118,N_17967,N_17903);
and U18119 (N_18119,N_17994,N_17817);
nand U18120 (N_18120,N_17828,N_17810);
nor U18121 (N_18121,N_17821,N_17938);
nor U18122 (N_18122,N_17986,N_17910);
and U18123 (N_18123,N_17976,N_17909);
xor U18124 (N_18124,N_17878,N_17920);
nor U18125 (N_18125,N_17812,N_17864);
and U18126 (N_18126,N_17811,N_17974);
nor U18127 (N_18127,N_17963,N_17920);
nor U18128 (N_18128,N_17855,N_17941);
and U18129 (N_18129,N_17903,N_17858);
and U18130 (N_18130,N_17904,N_17866);
and U18131 (N_18131,N_17993,N_17941);
or U18132 (N_18132,N_17840,N_17933);
or U18133 (N_18133,N_17850,N_17915);
or U18134 (N_18134,N_17872,N_17959);
xor U18135 (N_18135,N_17962,N_17991);
and U18136 (N_18136,N_17856,N_17814);
and U18137 (N_18137,N_17827,N_17951);
and U18138 (N_18138,N_17937,N_17800);
and U18139 (N_18139,N_17907,N_17997);
or U18140 (N_18140,N_17830,N_17883);
nor U18141 (N_18141,N_17924,N_17975);
nand U18142 (N_18142,N_17990,N_17812);
nand U18143 (N_18143,N_17908,N_17857);
nand U18144 (N_18144,N_17988,N_17997);
xnor U18145 (N_18145,N_17833,N_17853);
and U18146 (N_18146,N_17983,N_17862);
and U18147 (N_18147,N_17871,N_17983);
or U18148 (N_18148,N_17967,N_17977);
and U18149 (N_18149,N_17955,N_17821);
and U18150 (N_18150,N_17927,N_17961);
xor U18151 (N_18151,N_17841,N_17953);
nand U18152 (N_18152,N_17853,N_17940);
or U18153 (N_18153,N_17815,N_17950);
and U18154 (N_18154,N_17825,N_17815);
xnor U18155 (N_18155,N_17979,N_17929);
or U18156 (N_18156,N_17933,N_17871);
nor U18157 (N_18157,N_17844,N_17929);
nor U18158 (N_18158,N_17979,N_17881);
nor U18159 (N_18159,N_17866,N_17849);
xor U18160 (N_18160,N_17966,N_17816);
xnor U18161 (N_18161,N_17932,N_17870);
nand U18162 (N_18162,N_17877,N_17825);
nand U18163 (N_18163,N_17952,N_17989);
nor U18164 (N_18164,N_17836,N_17965);
nor U18165 (N_18165,N_17983,N_17971);
nor U18166 (N_18166,N_17811,N_17822);
and U18167 (N_18167,N_17911,N_17990);
nor U18168 (N_18168,N_17982,N_17808);
xnor U18169 (N_18169,N_17884,N_17839);
nand U18170 (N_18170,N_17814,N_17837);
or U18171 (N_18171,N_17833,N_17887);
and U18172 (N_18172,N_17832,N_17910);
nand U18173 (N_18173,N_17854,N_17800);
or U18174 (N_18174,N_17964,N_17891);
nand U18175 (N_18175,N_17971,N_17995);
nand U18176 (N_18176,N_17824,N_17954);
or U18177 (N_18177,N_17884,N_17840);
xor U18178 (N_18178,N_17877,N_17933);
nand U18179 (N_18179,N_17823,N_17889);
xnor U18180 (N_18180,N_17860,N_17890);
xor U18181 (N_18181,N_17823,N_17860);
and U18182 (N_18182,N_17856,N_17958);
or U18183 (N_18183,N_17930,N_17889);
nor U18184 (N_18184,N_17834,N_17800);
xor U18185 (N_18185,N_17838,N_17859);
nand U18186 (N_18186,N_17945,N_17864);
nand U18187 (N_18187,N_17871,N_17884);
nor U18188 (N_18188,N_17891,N_17936);
or U18189 (N_18189,N_17840,N_17804);
or U18190 (N_18190,N_17923,N_17913);
nand U18191 (N_18191,N_17894,N_17832);
xor U18192 (N_18192,N_17888,N_17981);
and U18193 (N_18193,N_17882,N_17941);
or U18194 (N_18194,N_17894,N_17939);
xor U18195 (N_18195,N_17805,N_17835);
and U18196 (N_18196,N_17978,N_17840);
and U18197 (N_18197,N_17853,N_17845);
nor U18198 (N_18198,N_17939,N_17958);
xor U18199 (N_18199,N_17838,N_17867);
and U18200 (N_18200,N_18162,N_18019);
nor U18201 (N_18201,N_18006,N_18059);
or U18202 (N_18202,N_18137,N_18150);
nand U18203 (N_18203,N_18144,N_18194);
and U18204 (N_18204,N_18106,N_18133);
and U18205 (N_18205,N_18062,N_18053);
nand U18206 (N_18206,N_18061,N_18085);
nand U18207 (N_18207,N_18088,N_18078);
or U18208 (N_18208,N_18154,N_18192);
nor U18209 (N_18209,N_18158,N_18185);
xnor U18210 (N_18210,N_18069,N_18096);
or U18211 (N_18211,N_18091,N_18083);
nor U18212 (N_18212,N_18094,N_18122);
xor U18213 (N_18213,N_18152,N_18020);
nand U18214 (N_18214,N_18128,N_18125);
and U18215 (N_18215,N_18012,N_18063);
and U18216 (N_18216,N_18140,N_18171);
or U18217 (N_18217,N_18101,N_18027);
nor U18218 (N_18218,N_18195,N_18161);
nand U18219 (N_18219,N_18017,N_18193);
or U18220 (N_18220,N_18198,N_18180);
nand U18221 (N_18221,N_18084,N_18108);
xor U18222 (N_18222,N_18025,N_18037);
xor U18223 (N_18223,N_18112,N_18100);
or U18224 (N_18224,N_18040,N_18132);
xor U18225 (N_18225,N_18015,N_18079);
xnor U18226 (N_18226,N_18159,N_18119);
nand U18227 (N_18227,N_18157,N_18107);
nor U18228 (N_18228,N_18076,N_18110);
and U18229 (N_18229,N_18102,N_18167);
nand U18230 (N_18230,N_18064,N_18072);
and U18231 (N_18231,N_18135,N_18087);
nand U18232 (N_18232,N_18034,N_18190);
nand U18233 (N_18233,N_18138,N_18127);
or U18234 (N_18234,N_18098,N_18036);
nand U18235 (N_18235,N_18163,N_18058);
or U18236 (N_18236,N_18000,N_18042);
and U18237 (N_18237,N_18104,N_18074);
or U18238 (N_18238,N_18177,N_18024);
xor U18239 (N_18239,N_18089,N_18156);
xor U18240 (N_18240,N_18183,N_18035);
and U18241 (N_18241,N_18187,N_18052);
nor U18242 (N_18242,N_18188,N_18067);
nor U18243 (N_18243,N_18124,N_18103);
or U18244 (N_18244,N_18115,N_18048);
nand U18245 (N_18245,N_18046,N_18005);
and U18246 (N_18246,N_18118,N_18149);
xor U18247 (N_18247,N_18120,N_18197);
xor U18248 (N_18248,N_18174,N_18050);
nor U18249 (N_18249,N_18142,N_18029);
nor U18250 (N_18250,N_18105,N_18054);
and U18251 (N_18251,N_18051,N_18033);
nand U18252 (N_18252,N_18070,N_18126);
nand U18253 (N_18253,N_18099,N_18186);
or U18254 (N_18254,N_18191,N_18155);
and U18255 (N_18255,N_18014,N_18049);
or U18256 (N_18256,N_18129,N_18093);
xnor U18257 (N_18257,N_18116,N_18199);
or U18258 (N_18258,N_18179,N_18032);
or U18259 (N_18259,N_18045,N_18153);
and U18260 (N_18260,N_18090,N_18009);
or U18261 (N_18261,N_18041,N_18131);
or U18262 (N_18262,N_18022,N_18139);
and U18263 (N_18263,N_18189,N_18008);
nand U18264 (N_18264,N_18134,N_18143);
and U18265 (N_18265,N_18007,N_18055);
or U18266 (N_18266,N_18111,N_18003);
xnor U18267 (N_18267,N_18172,N_18146);
xnor U18268 (N_18268,N_18184,N_18011);
nor U18269 (N_18269,N_18175,N_18018);
nand U18270 (N_18270,N_18038,N_18165);
or U18271 (N_18271,N_18056,N_18130);
nor U18272 (N_18272,N_18004,N_18182);
or U18273 (N_18273,N_18031,N_18021);
and U18274 (N_18274,N_18023,N_18114);
or U18275 (N_18275,N_18121,N_18071);
and U18276 (N_18276,N_18044,N_18097);
nor U18277 (N_18277,N_18145,N_18082);
and U18278 (N_18278,N_18136,N_18010);
or U18279 (N_18279,N_18039,N_18043);
or U18280 (N_18280,N_18123,N_18095);
nor U18281 (N_18281,N_18168,N_18147);
or U18282 (N_18282,N_18001,N_18170);
and U18283 (N_18283,N_18113,N_18117);
nor U18284 (N_18284,N_18151,N_18173);
and U18285 (N_18285,N_18178,N_18077);
xnor U18286 (N_18286,N_18057,N_18016);
nand U18287 (N_18287,N_18075,N_18164);
xnor U18288 (N_18288,N_18109,N_18081);
or U18289 (N_18289,N_18030,N_18013);
or U18290 (N_18290,N_18196,N_18028);
and U18291 (N_18291,N_18002,N_18148);
or U18292 (N_18292,N_18181,N_18066);
nor U18293 (N_18293,N_18047,N_18065);
and U18294 (N_18294,N_18086,N_18160);
xor U18295 (N_18295,N_18068,N_18073);
and U18296 (N_18296,N_18141,N_18176);
nand U18297 (N_18297,N_18166,N_18092);
and U18298 (N_18298,N_18026,N_18080);
nor U18299 (N_18299,N_18169,N_18060);
nand U18300 (N_18300,N_18133,N_18104);
or U18301 (N_18301,N_18118,N_18133);
xor U18302 (N_18302,N_18070,N_18018);
or U18303 (N_18303,N_18003,N_18002);
and U18304 (N_18304,N_18071,N_18110);
or U18305 (N_18305,N_18141,N_18199);
or U18306 (N_18306,N_18007,N_18194);
or U18307 (N_18307,N_18161,N_18115);
and U18308 (N_18308,N_18133,N_18066);
and U18309 (N_18309,N_18153,N_18051);
nand U18310 (N_18310,N_18082,N_18099);
xnor U18311 (N_18311,N_18143,N_18054);
or U18312 (N_18312,N_18070,N_18151);
xor U18313 (N_18313,N_18004,N_18144);
nand U18314 (N_18314,N_18049,N_18161);
and U18315 (N_18315,N_18069,N_18050);
nand U18316 (N_18316,N_18191,N_18183);
nand U18317 (N_18317,N_18008,N_18111);
xnor U18318 (N_18318,N_18180,N_18095);
and U18319 (N_18319,N_18146,N_18009);
and U18320 (N_18320,N_18053,N_18061);
xor U18321 (N_18321,N_18170,N_18092);
nor U18322 (N_18322,N_18087,N_18076);
and U18323 (N_18323,N_18124,N_18051);
and U18324 (N_18324,N_18140,N_18001);
xnor U18325 (N_18325,N_18122,N_18049);
or U18326 (N_18326,N_18118,N_18181);
and U18327 (N_18327,N_18161,N_18144);
xor U18328 (N_18328,N_18171,N_18134);
xnor U18329 (N_18329,N_18115,N_18019);
xor U18330 (N_18330,N_18182,N_18190);
nor U18331 (N_18331,N_18175,N_18172);
nand U18332 (N_18332,N_18015,N_18084);
nand U18333 (N_18333,N_18108,N_18100);
nor U18334 (N_18334,N_18034,N_18037);
nand U18335 (N_18335,N_18174,N_18082);
nor U18336 (N_18336,N_18151,N_18134);
or U18337 (N_18337,N_18001,N_18167);
or U18338 (N_18338,N_18172,N_18124);
nand U18339 (N_18339,N_18049,N_18145);
nor U18340 (N_18340,N_18157,N_18106);
or U18341 (N_18341,N_18111,N_18104);
nor U18342 (N_18342,N_18040,N_18092);
and U18343 (N_18343,N_18028,N_18167);
or U18344 (N_18344,N_18125,N_18000);
or U18345 (N_18345,N_18118,N_18155);
or U18346 (N_18346,N_18062,N_18090);
xnor U18347 (N_18347,N_18116,N_18066);
nand U18348 (N_18348,N_18157,N_18139);
nand U18349 (N_18349,N_18014,N_18064);
xnor U18350 (N_18350,N_18181,N_18088);
xor U18351 (N_18351,N_18004,N_18195);
or U18352 (N_18352,N_18029,N_18109);
xnor U18353 (N_18353,N_18150,N_18104);
or U18354 (N_18354,N_18086,N_18116);
and U18355 (N_18355,N_18149,N_18003);
xor U18356 (N_18356,N_18098,N_18019);
nand U18357 (N_18357,N_18057,N_18102);
and U18358 (N_18358,N_18188,N_18127);
xnor U18359 (N_18359,N_18094,N_18086);
or U18360 (N_18360,N_18103,N_18002);
nor U18361 (N_18361,N_18055,N_18041);
and U18362 (N_18362,N_18114,N_18039);
nor U18363 (N_18363,N_18133,N_18127);
xnor U18364 (N_18364,N_18189,N_18064);
xor U18365 (N_18365,N_18111,N_18108);
nor U18366 (N_18366,N_18011,N_18126);
and U18367 (N_18367,N_18003,N_18185);
nor U18368 (N_18368,N_18101,N_18173);
nand U18369 (N_18369,N_18009,N_18021);
and U18370 (N_18370,N_18137,N_18159);
and U18371 (N_18371,N_18198,N_18124);
nor U18372 (N_18372,N_18049,N_18100);
or U18373 (N_18373,N_18078,N_18027);
nand U18374 (N_18374,N_18194,N_18155);
and U18375 (N_18375,N_18061,N_18115);
xnor U18376 (N_18376,N_18149,N_18085);
nor U18377 (N_18377,N_18031,N_18136);
or U18378 (N_18378,N_18021,N_18073);
nor U18379 (N_18379,N_18179,N_18107);
nor U18380 (N_18380,N_18112,N_18049);
or U18381 (N_18381,N_18195,N_18125);
or U18382 (N_18382,N_18124,N_18046);
or U18383 (N_18383,N_18060,N_18078);
xor U18384 (N_18384,N_18029,N_18051);
nand U18385 (N_18385,N_18011,N_18032);
and U18386 (N_18386,N_18191,N_18197);
or U18387 (N_18387,N_18098,N_18154);
and U18388 (N_18388,N_18056,N_18093);
xor U18389 (N_18389,N_18174,N_18077);
nand U18390 (N_18390,N_18050,N_18022);
nor U18391 (N_18391,N_18069,N_18028);
nand U18392 (N_18392,N_18060,N_18014);
nand U18393 (N_18393,N_18043,N_18120);
or U18394 (N_18394,N_18110,N_18127);
xor U18395 (N_18395,N_18157,N_18164);
or U18396 (N_18396,N_18019,N_18064);
nor U18397 (N_18397,N_18123,N_18016);
nand U18398 (N_18398,N_18144,N_18183);
xnor U18399 (N_18399,N_18163,N_18165);
or U18400 (N_18400,N_18294,N_18391);
and U18401 (N_18401,N_18330,N_18210);
nand U18402 (N_18402,N_18336,N_18309);
or U18403 (N_18403,N_18381,N_18252);
nor U18404 (N_18404,N_18350,N_18259);
or U18405 (N_18405,N_18378,N_18370);
nor U18406 (N_18406,N_18207,N_18367);
xnor U18407 (N_18407,N_18329,N_18316);
nor U18408 (N_18408,N_18244,N_18254);
or U18409 (N_18409,N_18303,N_18343);
nor U18410 (N_18410,N_18286,N_18392);
nor U18411 (N_18411,N_18268,N_18200);
or U18412 (N_18412,N_18393,N_18347);
and U18413 (N_18413,N_18293,N_18237);
nor U18414 (N_18414,N_18364,N_18306);
nor U18415 (N_18415,N_18365,N_18340);
xor U18416 (N_18416,N_18319,N_18265);
nor U18417 (N_18417,N_18250,N_18387);
nor U18418 (N_18418,N_18235,N_18284);
or U18419 (N_18419,N_18221,N_18380);
xnor U18420 (N_18420,N_18247,N_18264);
nor U18421 (N_18421,N_18311,N_18389);
nand U18422 (N_18422,N_18262,N_18217);
and U18423 (N_18423,N_18332,N_18351);
nor U18424 (N_18424,N_18338,N_18339);
or U18425 (N_18425,N_18271,N_18276);
and U18426 (N_18426,N_18395,N_18223);
xnor U18427 (N_18427,N_18201,N_18206);
nand U18428 (N_18428,N_18325,N_18398);
or U18429 (N_18429,N_18241,N_18372);
xnor U18430 (N_18430,N_18234,N_18256);
or U18431 (N_18431,N_18238,N_18231);
nor U18432 (N_18432,N_18226,N_18305);
nand U18433 (N_18433,N_18356,N_18292);
or U18434 (N_18434,N_18317,N_18242);
nor U18435 (N_18435,N_18344,N_18353);
nand U18436 (N_18436,N_18310,N_18354);
nor U18437 (N_18437,N_18366,N_18346);
nor U18438 (N_18438,N_18218,N_18272);
xor U18439 (N_18439,N_18248,N_18215);
and U18440 (N_18440,N_18204,N_18257);
nand U18441 (N_18441,N_18359,N_18283);
nor U18442 (N_18442,N_18225,N_18361);
and U18443 (N_18443,N_18342,N_18261);
nor U18444 (N_18444,N_18296,N_18239);
and U18445 (N_18445,N_18287,N_18321);
xnor U18446 (N_18446,N_18358,N_18349);
or U18447 (N_18447,N_18320,N_18270);
or U18448 (N_18448,N_18281,N_18352);
and U18449 (N_18449,N_18327,N_18299);
xnor U18450 (N_18450,N_18212,N_18377);
nand U18451 (N_18451,N_18363,N_18369);
nor U18452 (N_18452,N_18253,N_18341);
nand U18453 (N_18453,N_18355,N_18297);
xor U18454 (N_18454,N_18373,N_18227);
nand U18455 (N_18455,N_18232,N_18295);
and U18456 (N_18456,N_18384,N_18382);
xor U18457 (N_18457,N_18345,N_18279);
and U18458 (N_18458,N_18229,N_18277);
and U18459 (N_18459,N_18209,N_18326);
nor U18460 (N_18460,N_18360,N_18396);
or U18461 (N_18461,N_18333,N_18394);
nand U18462 (N_18462,N_18203,N_18285);
nand U18463 (N_18463,N_18278,N_18267);
nand U18464 (N_18464,N_18307,N_18216);
xor U18465 (N_18465,N_18385,N_18202);
nor U18466 (N_18466,N_18314,N_18245);
and U18467 (N_18467,N_18255,N_18375);
or U18468 (N_18468,N_18280,N_18258);
or U18469 (N_18469,N_18390,N_18362);
and U18470 (N_18470,N_18328,N_18266);
xor U18471 (N_18471,N_18224,N_18301);
or U18472 (N_18472,N_18230,N_18282);
nand U18473 (N_18473,N_18376,N_18291);
nor U18474 (N_18474,N_18368,N_18318);
and U18475 (N_18475,N_18397,N_18348);
or U18476 (N_18476,N_18379,N_18304);
or U18477 (N_18477,N_18249,N_18313);
nand U18478 (N_18478,N_18334,N_18308);
nor U18479 (N_18479,N_18208,N_18288);
and U18480 (N_18480,N_18246,N_18240);
or U18481 (N_18481,N_18399,N_18275);
nor U18482 (N_18482,N_18219,N_18236);
or U18483 (N_18483,N_18323,N_18322);
nor U18484 (N_18484,N_18233,N_18386);
nand U18485 (N_18485,N_18383,N_18371);
nand U18486 (N_18486,N_18220,N_18300);
and U18487 (N_18487,N_18211,N_18324);
or U18488 (N_18488,N_18331,N_18205);
nor U18489 (N_18489,N_18243,N_18315);
or U18490 (N_18490,N_18289,N_18312);
nand U18491 (N_18491,N_18263,N_18337);
nand U18492 (N_18492,N_18298,N_18213);
nand U18493 (N_18493,N_18260,N_18222);
xor U18494 (N_18494,N_18269,N_18274);
and U18495 (N_18495,N_18357,N_18214);
or U18496 (N_18496,N_18388,N_18273);
and U18497 (N_18497,N_18228,N_18335);
or U18498 (N_18498,N_18290,N_18302);
xnor U18499 (N_18499,N_18374,N_18251);
or U18500 (N_18500,N_18294,N_18283);
nand U18501 (N_18501,N_18297,N_18317);
nor U18502 (N_18502,N_18218,N_18219);
nand U18503 (N_18503,N_18228,N_18292);
or U18504 (N_18504,N_18240,N_18255);
nand U18505 (N_18505,N_18369,N_18221);
nand U18506 (N_18506,N_18212,N_18293);
and U18507 (N_18507,N_18281,N_18372);
xnor U18508 (N_18508,N_18373,N_18253);
xnor U18509 (N_18509,N_18296,N_18275);
or U18510 (N_18510,N_18201,N_18274);
nand U18511 (N_18511,N_18222,N_18317);
and U18512 (N_18512,N_18300,N_18235);
and U18513 (N_18513,N_18248,N_18329);
or U18514 (N_18514,N_18228,N_18246);
nor U18515 (N_18515,N_18317,N_18271);
nor U18516 (N_18516,N_18370,N_18350);
or U18517 (N_18517,N_18293,N_18386);
or U18518 (N_18518,N_18213,N_18362);
xor U18519 (N_18519,N_18309,N_18265);
and U18520 (N_18520,N_18286,N_18271);
nand U18521 (N_18521,N_18357,N_18332);
xor U18522 (N_18522,N_18285,N_18234);
or U18523 (N_18523,N_18222,N_18384);
nand U18524 (N_18524,N_18243,N_18232);
or U18525 (N_18525,N_18288,N_18365);
nand U18526 (N_18526,N_18382,N_18377);
or U18527 (N_18527,N_18314,N_18229);
xor U18528 (N_18528,N_18247,N_18219);
nand U18529 (N_18529,N_18252,N_18245);
xnor U18530 (N_18530,N_18317,N_18341);
nand U18531 (N_18531,N_18278,N_18328);
and U18532 (N_18532,N_18365,N_18233);
nand U18533 (N_18533,N_18277,N_18390);
nor U18534 (N_18534,N_18235,N_18309);
xnor U18535 (N_18535,N_18218,N_18201);
nand U18536 (N_18536,N_18394,N_18224);
xor U18537 (N_18537,N_18278,N_18341);
and U18538 (N_18538,N_18385,N_18274);
or U18539 (N_18539,N_18280,N_18374);
nand U18540 (N_18540,N_18339,N_18275);
nor U18541 (N_18541,N_18251,N_18354);
nor U18542 (N_18542,N_18351,N_18213);
and U18543 (N_18543,N_18372,N_18303);
or U18544 (N_18544,N_18301,N_18393);
or U18545 (N_18545,N_18308,N_18390);
and U18546 (N_18546,N_18298,N_18290);
xnor U18547 (N_18547,N_18272,N_18352);
xnor U18548 (N_18548,N_18255,N_18386);
xnor U18549 (N_18549,N_18320,N_18302);
and U18550 (N_18550,N_18216,N_18364);
xnor U18551 (N_18551,N_18203,N_18216);
nand U18552 (N_18552,N_18245,N_18238);
and U18553 (N_18553,N_18266,N_18234);
xor U18554 (N_18554,N_18319,N_18365);
xor U18555 (N_18555,N_18344,N_18311);
nor U18556 (N_18556,N_18382,N_18365);
nor U18557 (N_18557,N_18325,N_18379);
or U18558 (N_18558,N_18335,N_18214);
xor U18559 (N_18559,N_18314,N_18304);
xor U18560 (N_18560,N_18340,N_18344);
nand U18561 (N_18561,N_18307,N_18251);
and U18562 (N_18562,N_18232,N_18360);
and U18563 (N_18563,N_18278,N_18327);
nor U18564 (N_18564,N_18341,N_18304);
and U18565 (N_18565,N_18280,N_18279);
nand U18566 (N_18566,N_18220,N_18229);
or U18567 (N_18567,N_18365,N_18216);
or U18568 (N_18568,N_18396,N_18361);
nor U18569 (N_18569,N_18342,N_18251);
and U18570 (N_18570,N_18311,N_18296);
nand U18571 (N_18571,N_18331,N_18226);
and U18572 (N_18572,N_18217,N_18351);
and U18573 (N_18573,N_18327,N_18306);
xor U18574 (N_18574,N_18396,N_18390);
and U18575 (N_18575,N_18375,N_18239);
or U18576 (N_18576,N_18282,N_18382);
nor U18577 (N_18577,N_18311,N_18348);
nor U18578 (N_18578,N_18310,N_18281);
nand U18579 (N_18579,N_18317,N_18345);
nand U18580 (N_18580,N_18385,N_18240);
and U18581 (N_18581,N_18323,N_18203);
nand U18582 (N_18582,N_18298,N_18226);
nor U18583 (N_18583,N_18267,N_18399);
or U18584 (N_18584,N_18316,N_18388);
nor U18585 (N_18585,N_18356,N_18231);
nor U18586 (N_18586,N_18343,N_18270);
nand U18587 (N_18587,N_18305,N_18343);
or U18588 (N_18588,N_18267,N_18313);
or U18589 (N_18589,N_18238,N_18298);
nor U18590 (N_18590,N_18256,N_18203);
nor U18591 (N_18591,N_18354,N_18229);
nand U18592 (N_18592,N_18291,N_18377);
nor U18593 (N_18593,N_18336,N_18296);
or U18594 (N_18594,N_18269,N_18254);
xor U18595 (N_18595,N_18298,N_18202);
nand U18596 (N_18596,N_18359,N_18394);
or U18597 (N_18597,N_18304,N_18203);
xor U18598 (N_18598,N_18258,N_18344);
and U18599 (N_18599,N_18285,N_18353);
or U18600 (N_18600,N_18478,N_18566);
or U18601 (N_18601,N_18570,N_18511);
nand U18602 (N_18602,N_18464,N_18580);
nand U18603 (N_18603,N_18448,N_18443);
nor U18604 (N_18604,N_18479,N_18585);
or U18605 (N_18605,N_18568,N_18544);
and U18606 (N_18606,N_18595,N_18537);
xor U18607 (N_18607,N_18527,N_18551);
or U18608 (N_18608,N_18477,N_18427);
and U18609 (N_18609,N_18574,N_18416);
and U18610 (N_18610,N_18526,N_18539);
or U18611 (N_18611,N_18474,N_18453);
nand U18612 (N_18612,N_18409,N_18548);
and U18613 (N_18613,N_18457,N_18414);
and U18614 (N_18614,N_18475,N_18470);
or U18615 (N_18615,N_18488,N_18456);
nor U18616 (N_18616,N_18410,N_18515);
nand U18617 (N_18617,N_18493,N_18408);
xnor U18618 (N_18618,N_18460,N_18517);
and U18619 (N_18619,N_18507,N_18582);
nand U18620 (N_18620,N_18500,N_18461);
nand U18621 (N_18621,N_18411,N_18407);
xor U18622 (N_18622,N_18417,N_18576);
nor U18623 (N_18623,N_18520,N_18487);
nor U18624 (N_18624,N_18578,N_18424);
nor U18625 (N_18625,N_18543,N_18429);
xnor U18626 (N_18626,N_18529,N_18405);
or U18627 (N_18627,N_18432,N_18450);
xnor U18628 (N_18628,N_18528,N_18555);
and U18629 (N_18629,N_18597,N_18506);
and U18630 (N_18630,N_18495,N_18445);
or U18631 (N_18631,N_18403,N_18471);
or U18632 (N_18632,N_18412,N_18567);
nor U18633 (N_18633,N_18430,N_18490);
or U18634 (N_18634,N_18459,N_18489);
and U18635 (N_18635,N_18428,N_18547);
and U18636 (N_18636,N_18501,N_18590);
nor U18637 (N_18637,N_18458,N_18485);
nand U18638 (N_18638,N_18513,N_18550);
nor U18639 (N_18639,N_18404,N_18447);
and U18640 (N_18640,N_18522,N_18473);
and U18641 (N_18641,N_18451,N_18402);
or U18642 (N_18642,N_18524,N_18521);
nand U18643 (N_18643,N_18554,N_18491);
xnor U18644 (N_18644,N_18469,N_18433);
nor U18645 (N_18645,N_18577,N_18545);
nand U18646 (N_18646,N_18426,N_18497);
nand U18647 (N_18647,N_18540,N_18423);
xor U18648 (N_18648,N_18465,N_18421);
or U18649 (N_18649,N_18535,N_18468);
and U18650 (N_18650,N_18594,N_18444);
xnor U18651 (N_18651,N_18466,N_18599);
nor U18652 (N_18652,N_18519,N_18586);
and U18653 (N_18653,N_18542,N_18439);
nand U18654 (N_18654,N_18549,N_18484);
nand U18655 (N_18655,N_18492,N_18467);
nor U18656 (N_18656,N_18588,N_18502);
and U18657 (N_18657,N_18406,N_18565);
nor U18658 (N_18658,N_18591,N_18514);
or U18659 (N_18659,N_18573,N_18505);
or U18660 (N_18660,N_18532,N_18481);
nor U18661 (N_18661,N_18476,N_18592);
nor U18662 (N_18662,N_18418,N_18431);
nand U18663 (N_18663,N_18496,N_18499);
xnor U18664 (N_18664,N_18498,N_18569);
and U18665 (N_18665,N_18446,N_18516);
nand U18666 (N_18666,N_18572,N_18434);
or U18667 (N_18667,N_18531,N_18454);
and U18668 (N_18668,N_18449,N_18546);
nand U18669 (N_18669,N_18509,N_18503);
and U18670 (N_18670,N_18441,N_18419);
xor U18671 (N_18671,N_18557,N_18425);
nor U18672 (N_18672,N_18536,N_18579);
nand U18673 (N_18673,N_18512,N_18518);
or U18674 (N_18674,N_18401,N_18523);
or U18675 (N_18675,N_18435,N_18482);
or U18676 (N_18676,N_18583,N_18472);
xnor U18677 (N_18677,N_18462,N_18400);
and U18678 (N_18678,N_18589,N_18571);
nor U18679 (N_18679,N_18525,N_18508);
or U18680 (N_18680,N_18538,N_18564);
nand U18681 (N_18681,N_18556,N_18413);
nand U18682 (N_18682,N_18442,N_18530);
and U18683 (N_18683,N_18598,N_18552);
nor U18684 (N_18684,N_18510,N_18581);
or U18685 (N_18685,N_18480,N_18438);
or U18686 (N_18686,N_18463,N_18560);
nand U18687 (N_18687,N_18436,N_18440);
or U18688 (N_18688,N_18420,N_18452);
nor U18689 (N_18689,N_18563,N_18533);
nor U18690 (N_18690,N_18486,N_18561);
and U18691 (N_18691,N_18575,N_18422);
nand U18692 (N_18692,N_18455,N_18559);
nand U18693 (N_18693,N_18483,N_18584);
nor U18694 (N_18694,N_18541,N_18593);
xnor U18695 (N_18695,N_18596,N_18504);
xor U18696 (N_18696,N_18534,N_18437);
nor U18697 (N_18697,N_18553,N_18558);
and U18698 (N_18698,N_18587,N_18415);
and U18699 (N_18699,N_18562,N_18494);
xor U18700 (N_18700,N_18461,N_18492);
xnor U18701 (N_18701,N_18505,N_18517);
or U18702 (N_18702,N_18479,N_18452);
xnor U18703 (N_18703,N_18437,N_18564);
xor U18704 (N_18704,N_18548,N_18494);
nor U18705 (N_18705,N_18493,N_18432);
nand U18706 (N_18706,N_18521,N_18548);
xnor U18707 (N_18707,N_18575,N_18446);
or U18708 (N_18708,N_18550,N_18479);
xor U18709 (N_18709,N_18560,N_18429);
or U18710 (N_18710,N_18494,N_18413);
xnor U18711 (N_18711,N_18486,N_18405);
nand U18712 (N_18712,N_18546,N_18475);
nand U18713 (N_18713,N_18431,N_18439);
nor U18714 (N_18714,N_18535,N_18517);
nand U18715 (N_18715,N_18500,N_18592);
xnor U18716 (N_18716,N_18428,N_18433);
nand U18717 (N_18717,N_18423,N_18518);
and U18718 (N_18718,N_18539,N_18428);
and U18719 (N_18719,N_18419,N_18488);
or U18720 (N_18720,N_18453,N_18546);
xnor U18721 (N_18721,N_18485,N_18546);
nor U18722 (N_18722,N_18455,N_18581);
nand U18723 (N_18723,N_18451,N_18442);
xnor U18724 (N_18724,N_18452,N_18579);
xor U18725 (N_18725,N_18545,N_18594);
xnor U18726 (N_18726,N_18542,N_18458);
nand U18727 (N_18727,N_18538,N_18569);
or U18728 (N_18728,N_18513,N_18462);
or U18729 (N_18729,N_18544,N_18417);
or U18730 (N_18730,N_18506,N_18554);
and U18731 (N_18731,N_18568,N_18593);
or U18732 (N_18732,N_18405,N_18400);
xnor U18733 (N_18733,N_18467,N_18594);
xnor U18734 (N_18734,N_18493,N_18589);
xnor U18735 (N_18735,N_18556,N_18554);
nor U18736 (N_18736,N_18421,N_18589);
nor U18737 (N_18737,N_18597,N_18534);
nor U18738 (N_18738,N_18593,N_18454);
or U18739 (N_18739,N_18512,N_18543);
and U18740 (N_18740,N_18453,N_18547);
nor U18741 (N_18741,N_18493,N_18557);
nor U18742 (N_18742,N_18466,N_18427);
nor U18743 (N_18743,N_18572,N_18490);
nand U18744 (N_18744,N_18578,N_18503);
or U18745 (N_18745,N_18488,N_18445);
nand U18746 (N_18746,N_18504,N_18483);
and U18747 (N_18747,N_18469,N_18526);
and U18748 (N_18748,N_18595,N_18428);
nor U18749 (N_18749,N_18527,N_18535);
and U18750 (N_18750,N_18422,N_18558);
and U18751 (N_18751,N_18525,N_18584);
nand U18752 (N_18752,N_18439,N_18451);
nor U18753 (N_18753,N_18504,N_18414);
xnor U18754 (N_18754,N_18555,N_18443);
or U18755 (N_18755,N_18419,N_18460);
xnor U18756 (N_18756,N_18461,N_18534);
or U18757 (N_18757,N_18505,N_18523);
xor U18758 (N_18758,N_18475,N_18455);
or U18759 (N_18759,N_18569,N_18506);
xnor U18760 (N_18760,N_18465,N_18459);
nor U18761 (N_18761,N_18582,N_18530);
xor U18762 (N_18762,N_18442,N_18598);
and U18763 (N_18763,N_18412,N_18497);
or U18764 (N_18764,N_18495,N_18551);
nor U18765 (N_18765,N_18488,N_18482);
nor U18766 (N_18766,N_18414,N_18580);
nand U18767 (N_18767,N_18576,N_18455);
and U18768 (N_18768,N_18422,N_18421);
and U18769 (N_18769,N_18572,N_18488);
or U18770 (N_18770,N_18475,N_18405);
nand U18771 (N_18771,N_18400,N_18420);
and U18772 (N_18772,N_18553,N_18444);
and U18773 (N_18773,N_18537,N_18436);
and U18774 (N_18774,N_18532,N_18447);
nand U18775 (N_18775,N_18593,N_18576);
or U18776 (N_18776,N_18472,N_18480);
and U18777 (N_18777,N_18497,N_18523);
nand U18778 (N_18778,N_18476,N_18491);
and U18779 (N_18779,N_18495,N_18518);
or U18780 (N_18780,N_18579,N_18518);
nand U18781 (N_18781,N_18579,N_18526);
xor U18782 (N_18782,N_18456,N_18432);
and U18783 (N_18783,N_18437,N_18505);
or U18784 (N_18784,N_18443,N_18449);
and U18785 (N_18785,N_18471,N_18543);
nor U18786 (N_18786,N_18409,N_18514);
nand U18787 (N_18787,N_18415,N_18502);
or U18788 (N_18788,N_18571,N_18524);
and U18789 (N_18789,N_18559,N_18451);
and U18790 (N_18790,N_18520,N_18536);
nor U18791 (N_18791,N_18497,N_18473);
and U18792 (N_18792,N_18570,N_18503);
nor U18793 (N_18793,N_18593,N_18467);
nor U18794 (N_18794,N_18415,N_18599);
xnor U18795 (N_18795,N_18442,N_18548);
or U18796 (N_18796,N_18446,N_18564);
or U18797 (N_18797,N_18592,N_18583);
nand U18798 (N_18798,N_18490,N_18451);
or U18799 (N_18799,N_18485,N_18445);
xor U18800 (N_18800,N_18610,N_18688);
or U18801 (N_18801,N_18602,N_18726);
nand U18802 (N_18802,N_18677,N_18727);
nor U18803 (N_18803,N_18614,N_18748);
or U18804 (N_18804,N_18762,N_18739);
or U18805 (N_18805,N_18655,N_18734);
and U18806 (N_18806,N_18669,N_18797);
or U18807 (N_18807,N_18722,N_18659);
xnor U18808 (N_18808,N_18755,N_18786);
and U18809 (N_18809,N_18766,N_18784);
and U18810 (N_18810,N_18643,N_18617);
and U18811 (N_18811,N_18639,N_18710);
xnor U18812 (N_18812,N_18737,N_18666);
xnor U18813 (N_18813,N_18633,N_18663);
or U18814 (N_18814,N_18767,N_18683);
nor U18815 (N_18815,N_18648,N_18746);
or U18816 (N_18816,N_18751,N_18763);
nor U18817 (N_18817,N_18634,N_18758);
xnor U18818 (N_18818,N_18676,N_18785);
nand U18819 (N_18819,N_18724,N_18750);
nand U18820 (N_18820,N_18601,N_18795);
nor U18821 (N_18821,N_18613,N_18628);
or U18822 (N_18822,N_18696,N_18778);
nor U18823 (N_18823,N_18749,N_18753);
and U18824 (N_18824,N_18627,N_18760);
xor U18825 (N_18825,N_18708,N_18703);
or U18826 (N_18826,N_18793,N_18773);
or U18827 (N_18827,N_18681,N_18651);
nand U18828 (N_18828,N_18667,N_18754);
xor U18829 (N_18829,N_18612,N_18671);
nand U18830 (N_18830,N_18641,N_18698);
or U18831 (N_18831,N_18656,N_18764);
and U18832 (N_18832,N_18680,N_18711);
nand U18833 (N_18833,N_18789,N_18745);
nor U18834 (N_18834,N_18777,N_18787);
or U18835 (N_18835,N_18661,N_18650);
nand U18836 (N_18836,N_18788,N_18713);
and U18837 (N_18837,N_18603,N_18660);
nand U18838 (N_18838,N_18619,N_18728);
and U18839 (N_18839,N_18640,N_18790);
nand U18840 (N_18840,N_18684,N_18717);
nor U18841 (N_18841,N_18630,N_18735);
nand U18842 (N_18842,N_18709,N_18765);
nand U18843 (N_18843,N_18647,N_18705);
and U18844 (N_18844,N_18772,N_18674);
nor U18845 (N_18845,N_18649,N_18692);
nand U18846 (N_18846,N_18798,N_18794);
nand U18847 (N_18847,N_18700,N_18679);
or U18848 (N_18848,N_18740,N_18620);
nand U18849 (N_18849,N_18637,N_18622);
nor U18850 (N_18850,N_18757,N_18704);
and U18851 (N_18851,N_18729,N_18699);
xnor U18852 (N_18852,N_18668,N_18686);
or U18853 (N_18853,N_18662,N_18621);
nand U18854 (N_18854,N_18744,N_18670);
xor U18855 (N_18855,N_18731,N_18780);
nor U18856 (N_18856,N_18720,N_18657);
nor U18857 (N_18857,N_18609,N_18629);
or U18858 (N_18858,N_18730,N_18687);
and U18859 (N_18859,N_18605,N_18646);
nand U18860 (N_18860,N_18636,N_18615);
nor U18861 (N_18861,N_18623,N_18685);
nor U18862 (N_18862,N_18718,N_18616);
and U18863 (N_18863,N_18626,N_18695);
nand U18864 (N_18864,N_18606,N_18691);
nor U18865 (N_18865,N_18768,N_18638);
xor U18866 (N_18866,N_18665,N_18721);
xnor U18867 (N_18867,N_18776,N_18752);
xor U18868 (N_18868,N_18608,N_18715);
nor U18869 (N_18869,N_18782,N_18658);
and U18870 (N_18870,N_18697,N_18631);
nor U18871 (N_18871,N_18642,N_18747);
or U18872 (N_18872,N_18652,N_18781);
nor U18873 (N_18873,N_18618,N_18733);
xor U18874 (N_18874,N_18664,N_18611);
nand U18875 (N_18875,N_18742,N_18672);
xnor U18876 (N_18876,N_18644,N_18792);
nor U18877 (N_18877,N_18723,N_18635);
and U18878 (N_18878,N_18796,N_18771);
or U18879 (N_18879,N_18707,N_18690);
or U18880 (N_18880,N_18654,N_18738);
nand U18881 (N_18881,N_18625,N_18719);
or U18882 (N_18882,N_18706,N_18743);
xor U18883 (N_18883,N_18600,N_18607);
nor U18884 (N_18884,N_18632,N_18736);
nand U18885 (N_18885,N_18783,N_18682);
nand U18886 (N_18886,N_18759,N_18689);
nor U18887 (N_18887,N_18714,N_18702);
xor U18888 (N_18888,N_18624,N_18774);
and U18889 (N_18889,N_18712,N_18673);
nand U18890 (N_18890,N_18675,N_18716);
and U18891 (N_18891,N_18779,N_18645);
xnor U18892 (N_18892,N_18791,N_18741);
nand U18893 (N_18893,N_18678,N_18604);
or U18894 (N_18894,N_18756,N_18769);
nand U18895 (N_18895,N_18732,N_18701);
nand U18896 (N_18896,N_18770,N_18653);
nor U18897 (N_18897,N_18694,N_18775);
nor U18898 (N_18898,N_18725,N_18761);
nor U18899 (N_18899,N_18799,N_18693);
and U18900 (N_18900,N_18771,N_18645);
and U18901 (N_18901,N_18741,N_18662);
nor U18902 (N_18902,N_18612,N_18738);
xnor U18903 (N_18903,N_18702,N_18690);
nand U18904 (N_18904,N_18702,N_18680);
or U18905 (N_18905,N_18749,N_18678);
and U18906 (N_18906,N_18765,N_18652);
and U18907 (N_18907,N_18783,N_18748);
nor U18908 (N_18908,N_18607,N_18734);
xor U18909 (N_18909,N_18667,N_18678);
nor U18910 (N_18910,N_18618,N_18760);
or U18911 (N_18911,N_18701,N_18683);
and U18912 (N_18912,N_18653,N_18799);
and U18913 (N_18913,N_18791,N_18665);
nor U18914 (N_18914,N_18678,N_18659);
and U18915 (N_18915,N_18707,N_18696);
and U18916 (N_18916,N_18696,N_18659);
or U18917 (N_18917,N_18735,N_18785);
nand U18918 (N_18918,N_18714,N_18671);
and U18919 (N_18919,N_18617,N_18739);
and U18920 (N_18920,N_18796,N_18751);
xor U18921 (N_18921,N_18795,N_18653);
nor U18922 (N_18922,N_18777,N_18723);
nand U18923 (N_18923,N_18784,N_18792);
and U18924 (N_18924,N_18729,N_18743);
nand U18925 (N_18925,N_18726,N_18724);
nand U18926 (N_18926,N_18638,N_18674);
xor U18927 (N_18927,N_18783,N_18605);
nand U18928 (N_18928,N_18714,N_18650);
nor U18929 (N_18929,N_18706,N_18758);
or U18930 (N_18930,N_18710,N_18617);
and U18931 (N_18931,N_18650,N_18726);
nand U18932 (N_18932,N_18668,N_18719);
nand U18933 (N_18933,N_18638,N_18647);
and U18934 (N_18934,N_18656,N_18671);
nor U18935 (N_18935,N_18799,N_18684);
or U18936 (N_18936,N_18750,N_18605);
xnor U18937 (N_18937,N_18674,N_18733);
and U18938 (N_18938,N_18744,N_18657);
xnor U18939 (N_18939,N_18729,N_18636);
nor U18940 (N_18940,N_18726,N_18729);
nand U18941 (N_18941,N_18695,N_18765);
nand U18942 (N_18942,N_18679,N_18716);
and U18943 (N_18943,N_18704,N_18700);
nand U18944 (N_18944,N_18725,N_18705);
nand U18945 (N_18945,N_18765,N_18677);
xnor U18946 (N_18946,N_18745,N_18608);
nand U18947 (N_18947,N_18767,N_18645);
xnor U18948 (N_18948,N_18652,N_18795);
nor U18949 (N_18949,N_18784,N_18684);
nor U18950 (N_18950,N_18770,N_18761);
nand U18951 (N_18951,N_18776,N_18654);
and U18952 (N_18952,N_18704,N_18753);
nor U18953 (N_18953,N_18605,N_18630);
nand U18954 (N_18954,N_18700,N_18780);
and U18955 (N_18955,N_18736,N_18680);
nor U18956 (N_18956,N_18676,N_18684);
or U18957 (N_18957,N_18650,N_18730);
nand U18958 (N_18958,N_18703,N_18698);
xnor U18959 (N_18959,N_18622,N_18702);
nor U18960 (N_18960,N_18671,N_18672);
and U18961 (N_18961,N_18703,N_18619);
and U18962 (N_18962,N_18682,N_18709);
and U18963 (N_18963,N_18619,N_18652);
or U18964 (N_18964,N_18674,N_18684);
nor U18965 (N_18965,N_18611,N_18769);
and U18966 (N_18966,N_18701,N_18687);
or U18967 (N_18967,N_18630,N_18662);
xnor U18968 (N_18968,N_18639,N_18635);
nor U18969 (N_18969,N_18777,N_18739);
nand U18970 (N_18970,N_18687,N_18639);
nor U18971 (N_18971,N_18788,N_18771);
or U18972 (N_18972,N_18794,N_18739);
nor U18973 (N_18973,N_18636,N_18721);
xor U18974 (N_18974,N_18767,N_18636);
xor U18975 (N_18975,N_18639,N_18670);
or U18976 (N_18976,N_18716,N_18614);
or U18977 (N_18977,N_18717,N_18782);
and U18978 (N_18978,N_18621,N_18695);
nor U18979 (N_18979,N_18715,N_18770);
nor U18980 (N_18980,N_18612,N_18713);
nor U18981 (N_18981,N_18657,N_18683);
nand U18982 (N_18982,N_18630,N_18637);
nand U18983 (N_18983,N_18653,N_18759);
nand U18984 (N_18984,N_18664,N_18721);
or U18985 (N_18985,N_18724,N_18713);
nand U18986 (N_18986,N_18658,N_18634);
nand U18987 (N_18987,N_18656,N_18795);
and U18988 (N_18988,N_18754,N_18710);
or U18989 (N_18989,N_18702,N_18788);
nand U18990 (N_18990,N_18663,N_18699);
and U18991 (N_18991,N_18680,N_18694);
nand U18992 (N_18992,N_18739,N_18635);
or U18993 (N_18993,N_18749,N_18717);
or U18994 (N_18994,N_18790,N_18780);
or U18995 (N_18995,N_18600,N_18736);
and U18996 (N_18996,N_18791,N_18763);
xor U18997 (N_18997,N_18642,N_18714);
or U18998 (N_18998,N_18745,N_18754);
nor U18999 (N_18999,N_18651,N_18702);
or U19000 (N_19000,N_18864,N_18815);
xnor U19001 (N_19001,N_18909,N_18904);
or U19002 (N_19002,N_18944,N_18835);
and U19003 (N_19003,N_18968,N_18932);
xor U19004 (N_19004,N_18905,N_18858);
xor U19005 (N_19005,N_18908,N_18841);
nand U19006 (N_19006,N_18804,N_18906);
xnor U19007 (N_19007,N_18827,N_18868);
nor U19008 (N_19008,N_18936,N_18977);
nor U19009 (N_19009,N_18852,N_18990);
and U19010 (N_19010,N_18913,N_18998);
and U19011 (N_19011,N_18945,N_18888);
nor U19012 (N_19012,N_18927,N_18928);
nor U19013 (N_19013,N_18878,N_18991);
nor U19014 (N_19014,N_18870,N_18832);
and U19015 (N_19015,N_18987,N_18829);
xor U19016 (N_19016,N_18893,N_18846);
xor U19017 (N_19017,N_18853,N_18891);
nor U19018 (N_19018,N_18857,N_18881);
and U19019 (N_19019,N_18813,N_18923);
nand U19020 (N_19020,N_18890,N_18889);
nor U19021 (N_19021,N_18876,N_18942);
or U19022 (N_19022,N_18989,N_18924);
and U19023 (N_19023,N_18847,N_18951);
and U19024 (N_19024,N_18866,N_18974);
nor U19025 (N_19025,N_18988,N_18865);
or U19026 (N_19026,N_18900,N_18921);
nor U19027 (N_19027,N_18896,N_18976);
or U19028 (N_19028,N_18996,N_18872);
or U19029 (N_19029,N_18912,N_18862);
and U19030 (N_19030,N_18838,N_18980);
or U19031 (N_19031,N_18802,N_18933);
or U19032 (N_19032,N_18947,N_18837);
nor U19033 (N_19033,N_18819,N_18986);
and U19034 (N_19034,N_18810,N_18972);
and U19035 (N_19035,N_18825,N_18843);
nor U19036 (N_19036,N_18871,N_18885);
xnor U19037 (N_19037,N_18993,N_18950);
and U19038 (N_19038,N_18812,N_18879);
xnor U19039 (N_19039,N_18894,N_18946);
nor U19040 (N_19040,N_18961,N_18994);
or U19041 (N_19041,N_18897,N_18940);
and U19042 (N_19042,N_18823,N_18964);
xor U19043 (N_19043,N_18960,N_18820);
xor U19044 (N_19044,N_18954,N_18875);
and U19045 (N_19045,N_18939,N_18800);
nand U19046 (N_19046,N_18957,N_18929);
xor U19047 (N_19047,N_18886,N_18975);
or U19048 (N_19048,N_18952,N_18999);
nor U19049 (N_19049,N_18925,N_18930);
nor U19050 (N_19050,N_18839,N_18836);
and U19051 (N_19051,N_18801,N_18850);
nor U19052 (N_19052,N_18873,N_18808);
nor U19053 (N_19053,N_18816,N_18911);
and U19054 (N_19054,N_18874,N_18992);
xnor U19055 (N_19055,N_18822,N_18969);
or U19056 (N_19056,N_18985,N_18824);
and U19057 (N_19057,N_18867,N_18984);
and U19058 (N_19058,N_18895,N_18971);
xor U19059 (N_19059,N_18861,N_18811);
nand U19060 (N_19060,N_18883,N_18803);
xor U19061 (N_19061,N_18914,N_18834);
or U19062 (N_19062,N_18849,N_18915);
and U19063 (N_19063,N_18973,N_18920);
nand U19064 (N_19064,N_18860,N_18848);
xnor U19065 (N_19065,N_18807,N_18937);
nor U19066 (N_19066,N_18943,N_18809);
nand U19067 (N_19067,N_18917,N_18981);
xor U19068 (N_19068,N_18880,N_18863);
or U19069 (N_19069,N_18877,N_18855);
and U19070 (N_19070,N_18995,N_18997);
and U19071 (N_19071,N_18902,N_18959);
nor U19072 (N_19072,N_18931,N_18830);
or U19073 (N_19073,N_18826,N_18926);
or U19074 (N_19074,N_18948,N_18955);
nor U19075 (N_19075,N_18840,N_18956);
and U19076 (N_19076,N_18898,N_18983);
nor U19077 (N_19077,N_18935,N_18842);
or U19078 (N_19078,N_18982,N_18851);
xor U19079 (N_19079,N_18967,N_18949);
nor U19080 (N_19080,N_18910,N_18978);
nor U19081 (N_19081,N_18922,N_18806);
nand U19082 (N_19082,N_18884,N_18903);
and U19083 (N_19083,N_18882,N_18869);
nand U19084 (N_19084,N_18953,N_18833);
nor U19085 (N_19085,N_18965,N_18817);
xor U19086 (N_19086,N_18899,N_18963);
and U19087 (N_19087,N_18916,N_18979);
xnor U19088 (N_19088,N_18828,N_18887);
xor U19089 (N_19089,N_18831,N_18845);
nor U19090 (N_19090,N_18907,N_18814);
or U19091 (N_19091,N_18966,N_18854);
and U19092 (N_19092,N_18941,N_18856);
or U19093 (N_19093,N_18934,N_18901);
xor U19094 (N_19094,N_18962,N_18958);
nand U19095 (N_19095,N_18892,N_18821);
nand U19096 (N_19096,N_18919,N_18970);
and U19097 (N_19097,N_18805,N_18938);
nor U19098 (N_19098,N_18859,N_18918);
and U19099 (N_19099,N_18818,N_18844);
or U19100 (N_19100,N_18871,N_18914);
nor U19101 (N_19101,N_18896,N_18883);
nand U19102 (N_19102,N_18960,N_18832);
xor U19103 (N_19103,N_18869,N_18871);
or U19104 (N_19104,N_18882,N_18870);
and U19105 (N_19105,N_18860,N_18851);
xor U19106 (N_19106,N_18905,N_18918);
xnor U19107 (N_19107,N_18892,N_18990);
nand U19108 (N_19108,N_18951,N_18868);
xor U19109 (N_19109,N_18931,N_18917);
nor U19110 (N_19110,N_18805,N_18856);
nand U19111 (N_19111,N_18843,N_18918);
nor U19112 (N_19112,N_18930,N_18978);
nor U19113 (N_19113,N_18871,N_18889);
and U19114 (N_19114,N_18946,N_18961);
or U19115 (N_19115,N_18825,N_18928);
nand U19116 (N_19116,N_18979,N_18885);
xnor U19117 (N_19117,N_18986,N_18814);
xor U19118 (N_19118,N_18970,N_18991);
nor U19119 (N_19119,N_18880,N_18954);
or U19120 (N_19120,N_18996,N_18840);
and U19121 (N_19121,N_18957,N_18816);
and U19122 (N_19122,N_18817,N_18993);
and U19123 (N_19123,N_18931,N_18934);
or U19124 (N_19124,N_18903,N_18928);
nor U19125 (N_19125,N_18859,N_18882);
or U19126 (N_19126,N_18985,N_18860);
or U19127 (N_19127,N_18980,N_18869);
nor U19128 (N_19128,N_18961,N_18851);
xnor U19129 (N_19129,N_18925,N_18893);
or U19130 (N_19130,N_18872,N_18903);
xnor U19131 (N_19131,N_18867,N_18872);
or U19132 (N_19132,N_18945,N_18882);
nand U19133 (N_19133,N_18900,N_18872);
xnor U19134 (N_19134,N_18847,N_18905);
xnor U19135 (N_19135,N_18842,N_18985);
xor U19136 (N_19136,N_18863,N_18867);
and U19137 (N_19137,N_18904,N_18920);
and U19138 (N_19138,N_18852,N_18986);
nor U19139 (N_19139,N_18954,N_18902);
nor U19140 (N_19140,N_18979,N_18960);
nand U19141 (N_19141,N_18852,N_18805);
or U19142 (N_19142,N_18839,N_18808);
nand U19143 (N_19143,N_18948,N_18828);
nand U19144 (N_19144,N_18845,N_18804);
or U19145 (N_19145,N_18818,N_18952);
nand U19146 (N_19146,N_18903,N_18834);
and U19147 (N_19147,N_18897,N_18800);
and U19148 (N_19148,N_18816,N_18817);
and U19149 (N_19149,N_18980,N_18951);
nor U19150 (N_19150,N_18928,N_18916);
and U19151 (N_19151,N_18844,N_18906);
xnor U19152 (N_19152,N_18807,N_18883);
and U19153 (N_19153,N_18845,N_18963);
xnor U19154 (N_19154,N_18807,N_18829);
and U19155 (N_19155,N_18872,N_18889);
nand U19156 (N_19156,N_18954,N_18944);
nand U19157 (N_19157,N_18833,N_18851);
xnor U19158 (N_19158,N_18907,N_18826);
nor U19159 (N_19159,N_18911,N_18938);
or U19160 (N_19160,N_18922,N_18867);
nor U19161 (N_19161,N_18974,N_18939);
nand U19162 (N_19162,N_18809,N_18970);
and U19163 (N_19163,N_18832,N_18853);
nand U19164 (N_19164,N_18947,N_18840);
nand U19165 (N_19165,N_18875,N_18934);
or U19166 (N_19166,N_18816,N_18964);
or U19167 (N_19167,N_18889,N_18930);
nand U19168 (N_19168,N_18853,N_18958);
xnor U19169 (N_19169,N_18969,N_18872);
nand U19170 (N_19170,N_18906,N_18940);
xnor U19171 (N_19171,N_18871,N_18965);
nand U19172 (N_19172,N_18945,N_18877);
nand U19173 (N_19173,N_18839,N_18898);
xnor U19174 (N_19174,N_18872,N_18815);
nor U19175 (N_19175,N_18889,N_18905);
xnor U19176 (N_19176,N_18916,N_18900);
xor U19177 (N_19177,N_18909,N_18934);
or U19178 (N_19178,N_18994,N_18885);
xnor U19179 (N_19179,N_18964,N_18993);
nand U19180 (N_19180,N_18933,N_18854);
or U19181 (N_19181,N_18983,N_18904);
and U19182 (N_19182,N_18869,N_18959);
nor U19183 (N_19183,N_18907,N_18810);
xor U19184 (N_19184,N_18998,N_18853);
xnor U19185 (N_19185,N_18810,N_18870);
xor U19186 (N_19186,N_18956,N_18940);
nor U19187 (N_19187,N_18855,N_18806);
xor U19188 (N_19188,N_18891,N_18970);
nor U19189 (N_19189,N_18888,N_18866);
xor U19190 (N_19190,N_18800,N_18929);
xnor U19191 (N_19191,N_18999,N_18843);
xor U19192 (N_19192,N_18841,N_18988);
xnor U19193 (N_19193,N_18981,N_18865);
or U19194 (N_19194,N_18906,N_18854);
nor U19195 (N_19195,N_18939,N_18984);
xnor U19196 (N_19196,N_18837,N_18818);
nand U19197 (N_19197,N_18989,N_18804);
xor U19198 (N_19198,N_18984,N_18952);
or U19199 (N_19199,N_18911,N_18989);
or U19200 (N_19200,N_19193,N_19136);
and U19201 (N_19201,N_19013,N_19190);
nor U19202 (N_19202,N_19102,N_19081);
or U19203 (N_19203,N_19047,N_19056);
or U19204 (N_19204,N_19140,N_19128);
and U19205 (N_19205,N_19116,N_19018);
and U19206 (N_19206,N_19088,N_19164);
xnor U19207 (N_19207,N_19194,N_19113);
nor U19208 (N_19208,N_19134,N_19009);
xor U19209 (N_19209,N_19050,N_19185);
nor U19210 (N_19210,N_19179,N_19192);
and U19211 (N_19211,N_19044,N_19065);
and U19212 (N_19212,N_19106,N_19020);
and U19213 (N_19213,N_19072,N_19076);
or U19214 (N_19214,N_19145,N_19098);
or U19215 (N_19215,N_19173,N_19167);
or U19216 (N_19216,N_19135,N_19086);
xnor U19217 (N_19217,N_19114,N_19057);
xnor U19218 (N_19218,N_19168,N_19191);
and U19219 (N_19219,N_19046,N_19023);
nor U19220 (N_19220,N_19016,N_19012);
or U19221 (N_19221,N_19174,N_19127);
or U19222 (N_19222,N_19042,N_19077);
xnor U19223 (N_19223,N_19144,N_19015);
nand U19224 (N_19224,N_19131,N_19107);
and U19225 (N_19225,N_19039,N_19069);
and U19226 (N_19226,N_19026,N_19126);
xnor U19227 (N_19227,N_19125,N_19158);
and U19228 (N_19228,N_19100,N_19011);
or U19229 (N_19229,N_19138,N_19027);
nand U19230 (N_19230,N_19079,N_19051);
or U19231 (N_19231,N_19177,N_19034);
and U19232 (N_19232,N_19181,N_19119);
xor U19233 (N_19233,N_19176,N_19189);
nand U19234 (N_19234,N_19070,N_19137);
or U19235 (N_19235,N_19115,N_19172);
or U19236 (N_19236,N_19166,N_19058);
and U19237 (N_19237,N_19085,N_19175);
or U19238 (N_19238,N_19182,N_19035);
and U19239 (N_19239,N_19180,N_19092);
nand U19240 (N_19240,N_19161,N_19037);
xnor U19241 (N_19241,N_19075,N_19148);
nor U19242 (N_19242,N_19055,N_19066);
and U19243 (N_19243,N_19154,N_19087);
or U19244 (N_19244,N_19111,N_19082);
nand U19245 (N_19245,N_19094,N_19199);
or U19246 (N_19246,N_19063,N_19029);
nand U19247 (N_19247,N_19002,N_19089);
xor U19248 (N_19248,N_19053,N_19078);
and U19249 (N_19249,N_19083,N_19157);
nand U19250 (N_19250,N_19162,N_19061);
nand U19251 (N_19251,N_19062,N_19043);
nor U19252 (N_19252,N_19097,N_19188);
nand U19253 (N_19253,N_19093,N_19084);
nand U19254 (N_19254,N_19052,N_19030);
or U19255 (N_19255,N_19096,N_19007);
and U19256 (N_19256,N_19123,N_19187);
and U19257 (N_19257,N_19130,N_19095);
nor U19258 (N_19258,N_19198,N_19003);
xnor U19259 (N_19259,N_19155,N_19091);
xnor U19260 (N_19260,N_19129,N_19184);
xor U19261 (N_19261,N_19153,N_19197);
xor U19262 (N_19262,N_19060,N_19152);
xnor U19263 (N_19263,N_19170,N_19028);
nor U19264 (N_19264,N_19186,N_19151);
and U19265 (N_19265,N_19146,N_19143);
and U19266 (N_19266,N_19104,N_19171);
nand U19267 (N_19267,N_19169,N_19165);
nor U19268 (N_19268,N_19067,N_19159);
nand U19269 (N_19269,N_19118,N_19045);
xnor U19270 (N_19270,N_19054,N_19049);
or U19271 (N_19271,N_19059,N_19019);
nand U19272 (N_19272,N_19132,N_19041);
xnor U19273 (N_19273,N_19099,N_19147);
xnor U19274 (N_19274,N_19103,N_19001);
nor U19275 (N_19275,N_19110,N_19105);
and U19276 (N_19276,N_19160,N_19024);
nor U19277 (N_19277,N_19080,N_19101);
and U19278 (N_19278,N_19178,N_19149);
nand U19279 (N_19279,N_19010,N_19006);
nand U19280 (N_19280,N_19073,N_19040);
nand U19281 (N_19281,N_19150,N_19196);
xor U19282 (N_19282,N_19090,N_19031);
and U19283 (N_19283,N_19124,N_19033);
nor U19284 (N_19284,N_19195,N_19156);
xor U19285 (N_19285,N_19121,N_19000);
and U19286 (N_19286,N_19139,N_19133);
xnor U19287 (N_19287,N_19122,N_19109);
nand U19288 (N_19288,N_19141,N_19163);
nand U19289 (N_19289,N_19032,N_19183);
nand U19290 (N_19290,N_19142,N_19064);
nor U19291 (N_19291,N_19008,N_19038);
nor U19292 (N_19292,N_19005,N_19036);
nor U19293 (N_19293,N_19068,N_19112);
or U19294 (N_19294,N_19074,N_19022);
and U19295 (N_19295,N_19014,N_19108);
or U19296 (N_19296,N_19004,N_19017);
nor U19297 (N_19297,N_19048,N_19120);
nand U19298 (N_19298,N_19025,N_19117);
or U19299 (N_19299,N_19021,N_19071);
or U19300 (N_19300,N_19111,N_19038);
or U19301 (N_19301,N_19016,N_19092);
nand U19302 (N_19302,N_19107,N_19135);
xnor U19303 (N_19303,N_19154,N_19066);
nor U19304 (N_19304,N_19098,N_19009);
and U19305 (N_19305,N_19168,N_19197);
xnor U19306 (N_19306,N_19063,N_19026);
nand U19307 (N_19307,N_19177,N_19180);
and U19308 (N_19308,N_19132,N_19027);
and U19309 (N_19309,N_19008,N_19006);
nor U19310 (N_19310,N_19134,N_19071);
nor U19311 (N_19311,N_19075,N_19085);
nor U19312 (N_19312,N_19078,N_19036);
nand U19313 (N_19313,N_19194,N_19109);
or U19314 (N_19314,N_19131,N_19084);
nor U19315 (N_19315,N_19013,N_19082);
nand U19316 (N_19316,N_19087,N_19139);
and U19317 (N_19317,N_19004,N_19143);
and U19318 (N_19318,N_19033,N_19110);
or U19319 (N_19319,N_19055,N_19053);
or U19320 (N_19320,N_19076,N_19014);
and U19321 (N_19321,N_19061,N_19049);
or U19322 (N_19322,N_19095,N_19188);
and U19323 (N_19323,N_19109,N_19188);
nand U19324 (N_19324,N_19179,N_19067);
or U19325 (N_19325,N_19027,N_19079);
and U19326 (N_19326,N_19166,N_19044);
xnor U19327 (N_19327,N_19006,N_19197);
or U19328 (N_19328,N_19094,N_19108);
or U19329 (N_19329,N_19070,N_19068);
nor U19330 (N_19330,N_19013,N_19110);
nor U19331 (N_19331,N_19080,N_19171);
nor U19332 (N_19332,N_19187,N_19032);
or U19333 (N_19333,N_19047,N_19149);
nor U19334 (N_19334,N_19174,N_19034);
or U19335 (N_19335,N_19017,N_19016);
nand U19336 (N_19336,N_19174,N_19184);
or U19337 (N_19337,N_19119,N_19172);
xnor U19338 (N_19338,N_19101,N_19162);
and U19339 (N_19339,N_19162,N_19154);
and U19340 (N_19340,N_19047,N_19070);
nand U19341 (N_19341,N_19176,N_19005);
nor U19342 (N_19342,N_19018,N_19110);
xnor U19343 (N_19343,N_19097,N_19071);
nand U19344 (N_19344,N_19108,N_19033);
nand U19345 (N_19345,N_19087,N_19190);
nor U19346 (N_19346,N_19138,N_19024);
nand U19347 (N_19347,N_19145,N_19031);
or U19348 (N_19348,N_19184,N_19100);
xnor U19349 (N_19349,N_19101,N_19037);
or U19350 (N_19350,N_19070,N_19185);
xnor U19351 (N_19351,N_19152,N_19025);
xor U19352 (N_19352,N_19117,N_19156);
xor U19353 (N_19353,N_19198,N_19161);
nor U19354 (N_19354,N_19108,N_19158);
or U19355 (N_19355,N_19080,N_19134);
or U19356 (N_19356,N_19156,N_19102);
xnor U19357 (N_19357,N_19021,N_19042);
and U19358 (N_19358,N_19005,N_19142);
or U19359 (N_19359,N_19072,N_19155);
or U19360 (N_19360,N_19198,N_19073);
or U19361 (N_19361,N_19120,N_19135);
nand U19362 (N_19362,N_19126,N_19162);
xor U19363 (N_19363,N_19144,N_19180);
and U19364 (N_19364,N_19178,N_19179);
and U19365 (N_19365,N_19136,N_19199);
xor U19366 (N_19366,N_19062,N_19003);
nor U19367 (N_19367,N_19000,N_19185);
nor U19368 (N_19368,N_19140,N_19105);
nor U19369 (N_19369,N_19131,N_19046);
nor U19370 (N_19370,N_19117,N_19181);
nand U19371 (N_19371,N_19011,N_19111);
nand U19372 (N_19372,N_19193,N_19022);
and U19373 (N_19373,N_19083,N_19148);
and U19374 (N_19374,N_19128,N_19064);
xor U19375 (N_19375,N_19150,N_19031);
xor U19376 (N_19376,N_19186,N_19164);
or U19377 (N_19377,N_19151,N_19124);
and U19378 (N_19378,N_19149,N_19122);
nor U19379 (N_19379,N_19098,N_19194);
nand U19380 (N_19380,N_19121,N_19027);
nor U19381 (N_19381,N_19026,N_19080);
and U19382 (N_19382,N_19013,N_19023);
or U19383 (N_19383,N_19090,N_19124);
xor U19384 (N_19384,N_19071,N_19054);
nor U19385 (N_19385,N_19114,N_19059);
and U19386 (N_19386,N_19104,N_19023);
and U19387 (N_19387,N_19043,N_19042);
or U19388 (N_19388,N_19076,N_19031);
nand U19389 (N_19389,N_19153,N_19150);
xor U19390 (N_19390,N_19067,N_19117);
nor U19391 (N_19391,N_19014,N_19145);
nor U19392 (N_19392,N_19183,N_19157);
nor U19393 (N_19393,N_19126,N_19119);
or U19394 (N_19394,N_19067,N_19138);
xor U19395 (N_19395,N_19114,N_19098);
or U19396 (N_19396,N_19046,N_19077);
nor U19397 (N_19397,N_19030,N_19105);
nor U19398 (N_19398,N_19190,N_19044);
xor U19399 (N_19399,N_19114,N_19152);
nor U19400 (N_19400,N_19279,N_19350);
or U19401 (N_19401,N_19242,N_19268);
xnor U19402 (N_19402,N_19314,N_19271);
nand U19403 (N_19403,N_19281,N_19393);
and U19404 (N_19404,N_19259,N_19267);
xnor U19405 (N_19405,N_19331,N_19349);
or U19406 (N_19406,N_19395,N_19365);
nand U19407 (N_19407,N_19252,N_19347);
nor U19408 (N_19408,N_19231,N_19298);
nor U19409 (N_19409,N_19262,N_19381);
or U19410 (N_19410,N_19233,N_19261);
or U19411 (N_19411,N_19212,N_19317);
nor U19412 (N_19412,N_19200,N_19299);
and U19413 (N_19413,N_19228,N_19217);
xnor U19414 (N_19414,N_19239,N_19265);
xnor U19415 (N_19415,N_19370,N_19323);
xnor U19416 (N_19416,N_19294,N_19390);
or U19417 (N_19417,N_19332,N_19351);
nor U19418 (N_19418,N_19302,N_19247);
and U19419 (N_19419,N_19398,N_19205);
nand U19420 (N_19420,N_19328,N_19333);
xor U19421 (N_19421,N_19316,N_19293);
and U19422 (N_19422,N_19241,N_19288);
nand U19423 (N_19423,N_19270,N_19245);
xor U19424 (N_19424,N_19209,N_19218);
nor U19425 (N_19425,N_19246,N_19216);
nor U19426 (N_19426,N_19389,N_19287);
xor U19427 (N_19427,N_19263,N_19213);
or U19428 (N_19428,N_19321,N_19366);
or U19429 (N_19429,N_19301,N_19243);
xor U19430 (N_19430,N_19300,N_19324);
or U19431 (N_19431,N_19325,N_19282);
and U19432 (N_19432,N_19214,N_19318);
or U19433 (N_19433,N_19260,N_19235);
nor U19434 (N_19434,N_19211,N_19286);
xor U19435 (N_19435,N_19306,N_19221);
nand U19436 (N_19436,N_19319,N_19254);
or U19437 (N_19437,N_19358,N_19227);
and U19438 (N_19438,N_19308,N_19348);
xnor U19439 (N_19439,N_19326,N_19269);
or U19440 (N_19440,N_19232,N_19225);
xor U19441 (N_19441,N_19354,N_19355);
and U19442 (N_19442,N_19207,N_19344);
or U19443 (N_19443,N_19215,N_19255);
nand U19444 (N_19444,N_19357,N_19234);
or U19445 (N_19445,N_19334,N_19329);
or U19446 (N_19446,N_19368,N_19250);
or U19447 (N_19447,N_19285,N_19201);
nor U19448 (N_19448,N_19237,N_19304);
nand U19449 (N_19449,N_19283,N_19387);
and U19450 (N_19450,N_19210,N_19367);
or U19451 (N_19451,N_19361,N_19278);
nand U19452 (N_19452,N_19384,N_19284);
or U19453 (N_19453,N_19337,N_19330);
and U19454 (N_19454,N_19315,N_19388);
xnor U19455 (N_19455,N_19297,N_19391);
nor U19456 (N_19456,N_19343,N_19291);
nand U19457 (N_19457,N_19369,N_19360);
nand U19458 (N_19458,N_19296,N_19327);
or U19459 (N_19459,N_19258,N_19311);
xor U19460 (N_19460,N_19257,N_19379);
and U19461 (N_19461,N_19295,N_19399);
xor U19462 (N_19462,N_19394,N_19248);
and U19463 (N_19463,N_19385,N_19274);
nand U19464 (N_19464,N_19377,N_19386);
nand U19465 (N_19465,N_19292,N_19277);
xor U19466 (N_19466,N_19222,N_19346);
and U19467 (N_19467,N_19373,N_19356);
xnor U19468 (N_19468,N_19345,N_19249);
xor U19469 (N_19469,N_19396,N_19380);
nand U19470 (N_19470,N_19264,N_19305);
nand U19471 (N_19471,N_19338,N_19256);
nor U19472 (N_19472,N_19364,N_19303);
or U19473 (N_19473,N_19310,N_19378);
xnor U19474 (N_19474,N_19230,N_19266);
or U19475 (N_19475,N_19236,N_19289);
and U19476 (N_19476,N_19371,N_19203);
and U19477 (N_19477,N_19290,N_19353);
and U19478 (N_19478,N_19307,N_19280);
or U19479 (N_19479,N_19375,N_19229);
or U19480 (N_19480,N_19339,N_19224);
or U19481 (N_19481,N_19352,N_19275);
xnor U19482 (N_19482,N_19219,N_19340);
nor U19483 (N_19483,N_19240,N_19397);
nand U19484 (N_19484,N_19376,N_19251);
xnor U19485 (N_19485,N_19313,N_19382);
xnor U19486 (N_19486,N_19312,N_19206);
or U19487 (N_19487,N_19244,N_19363);
or U19488 (N_19488,N_19253,N_19208);
xnor U19489 (N_19489,N_19223,N_19204);
nand U19490 (N_19490,N_19362,N_19272);
or U19491 (N_19491,N_19273,N_19335);
nor U19492 (N_19492,N_19392,N_19359);
nand U19493 (N_19493,N_19202,N_19341);
and U19494 (N_19494,N_19372,N_19374);
nor U19495 (N_19495,N_19238,N_19226);
xor U19496 (N_19496,N_19220,N_19320);
nand U19497 (N_19497,N_19276,N_19383);
nand U19498 (N_19498,N_19342,N_19336);
nor U19499 (N_19499,N_19309,N_19322);
and U19500 (N_19500,N_19271,N_19359);
xnor U19501 (N_19501,N_19369,N_19371);
nand U19502 (N_19502,N_19398,N_19203);
and U19503 (N_19503,N_19394,N_19242);
and U19504 (N_19504,N_19287,N_19375);
or U19505 (N_19505,N_19229,N_19201);
xor U19506 (N_19506,N_19279,N_19207);
xnor U19507 (N_19507,N_19254,N_19305);
or U19508 (N_19508,N_19237,N_19256);
nor U19509 (N_19509,N_19222,N_19306);
xnor U19510 (N_19510,N_19296,N_19319);
xnor U19511 (N_19511,N_19235,N_19274);
or U19512 (N_19512,N_19338,N_19388);
or U19513 (N_19513,N_19372,N_19214);
or U19514 (N_19514,N_19294,N_19233);
or U19515 (N_19515,N_19222,N_19345);
nor U19516 (N_19516,N_19356,N_19371);
and U19517 (N_19517,N_19374,N_19268);
or U19518 (N_19518,N_19240,N_19309);
nand U19519 (N_19519,N_19283,N_19257);
and U19520 (N_19520,N_19389,N_19285);
nor U19521 (N_19521,N_19206,N_19243);
nor U19522 (N_19522,N_19229,N_19232);
xor U19523 (N_19523,N_19336,N_19349);
or U19524 (N_19524,N_19357,N_19388);
nand U19525 (N_19525,N_19383,N_19252);
xnor U19526 (N_19526,N_19393,N_19358);
or U19527 (N_19527,N_19356,N_19323);
nand U19528 (N_19528,N_19374,N_19210);
xnor U19529 (N_19529,N_19231,N_19316);
nor U19530 (N_19530,N_19293,N_19388);
nand U19531 (N_19531,N_19396,N_19312);
nor U19532 (N_19532,N_19232,N_19367);
nor U19533 (N_19533,N_19325,N_19284);
nor U19534 (N_19534,N_19298,N_19334);
or U19535 (N_19535,N_19291,N_19387);
and U19536 (N_19536,N_19279,N_19201);
nand U19537 (N_19537,N_19210,N_19387);
xnor U19538 (N_19538,N_19325,N_19341);
nor U19539 (N_19539,N_19390,N_19323);
nor U19540 (N_19540,N_19278,N_19399);
and U19541 (N_19541,N_19312,N_19330);
nand U19542 (N_19542,N_19316,N_19278);
or U19543 (N_19543,N_19283,N_19332);
and U19544 (N_19544,N_19202,N_19228);
and U19545 (N_19545,N_19343,N_19275);
or U19546 (N_19546,N_19362,N_19277);
nand U19547 (N_19547,N_19379,N_19286);
and U19548 (N_19548,N_19251,N_19345);
xor U19549 (N_19549,N_19359,N_19288);
and U19550 (N_19550,N_19203,N_19229);
nor U19551 (N_19551,N_19248,N_19301);
nand U19552 (N_19552,N_19267,N_19380);
or U19553 (N_19553,N_19327,N_19344);
nand U19554 (N_19554,N_19364,N_19361);
and U19555 (N_19555,N_19211,N_19222);
or U19556 (N_19556,N_19237,N_19263);
and U19557 (N_19557,N_19335,N_19345);
xnor U19558 (N_19558,N_19349,N_19372);
and U19559 (N_19559,N_19233,N_19205);
nand U19560 (N_19560,N_19217,N_19333);
and U19561 (N_19561,N_19310,N_19201);
xor U19562 (N_19562,N_19313,N_19357);
and U19563 (N_19563,N_19278,N_19328);
or U19564 (N_19564,N_19359,N_19280);
or U19565 (N_19565,N_19265,N_19205);
and U19566 (N_19566,N_19217,N_19237);
nand U19567 (N_19567,N_19368,N_19208);
or U19568 (N_19568,N_19248,N_19212);
or U19569 (N_19569,N_19241,N_19246);
and U19570 (N_19570,N_19306,N_19309);
nor U19571 (N_19571,N_19360,N_19213);
or U19572 (N_19572,N_19376,N_19249);
xnor U19573 (N_19573,N_19203,N_19238);
nand U19574 (N_19574,N_19266,N_19379);
xor U19575 (N_19575,N_19255,N_19380);
and U19576 (N_19576,N_19267,N_19367);
nand U19577 (N_19577,N_19260,N_19233);
nor U19578 (N_19578,N_19276,N_19363);
or U19579 (N_19579,N_19207,N_19218);
nor U19580 (N_19580,N_19317,N_19300);
nand U19581 (N_19581,N_19214,N_19347);
and U19582 (N_19582,N_19302,N_19281);
xor U19583 (N_19583,N_19383,N_19267);
xnor U19584 (N_19584,N_19384,N_19389);
or U19585 (N_19585,N_19341,N_19384);
nand U19586 (N_19586,N_19343,N_19356);
nand U19587 (N_19587,N_19393,N_19294);
xnor U19588 (N_19588,N_19378,N_19297);
nor U19589 (N_19589,N_19316,N_19374);
and U19590 (N_19590,N_19360,N_19362);
nand U19591 (N_19591,N_19338,N_19348);
nor U19592 (N_19592,N_19264,N_19221);
and U19593 (N_19593,N_19352,N_19345);
nand U19594 (N_19594,N_19395,N_19371);
nand U19595 (N_19595,N_19330,N_19245);
nor U19596 (N_19596,N_19327,N_19285);
xor U19597 (N_19597,N_19208,N_19248);
and U19598 (N_19598,N_19250,N_19243);
nor U19599 (N_19599,N_19326,N_19399);
or U19600 (N_19600,N_19575,N_19411);
nor U19601 (N_19601,N_19538,N_19406);
or U19602 (N_19602,N_19519,N_19467);
or U19603 (N_19603,N_19529,N_19469);
nor U19604 (N_19604,N_19487,N_19522);
or U19605 (N_19605,N_19426,N_19493);
or U19606 (N_19606,N_19562,N_19449);
nor U19607 (N_19607,N_19404,N_19596);
nand U19608 (N_19608,N_19581,N_19516);
nand U19609 (N_19609,N_19554,N_19434);
xnor U19610 (N_19610,N_19412,N_19503);
or U19611 (N_19611,N_19507,N_19428);
xor U19612 (N_19612,N_19501,N_19505);
or U19613 (N_19613,N_19565,N_19413);
xor U19614 (N_19614,N_19448,N_19474);
or U19615 (N_19615,N_19485,N_19541);
or U19616 (N_19616,N_19441,N_19588);
and U19617 (N_19617,N_19424,N_19436);
nor U19618 (N_19618,N_19417,N_19468);
or U19619 (N_19619,N_19542,N_19402);
xor U19620 (N_19620,N_19590,N_19582);
nor U19621 (N_19621,N_19400,N_19544);
or U19622 (N_19622,N_19460,N_19499);
nand U19623 (N_19623,N_19577,N_19466);
nand U19624 (N_19624,N_19414,N_19571);
xor U19625 (N_19625,N_19446,N_19586);
xnor U19626 (N_19626,N_19583,N_19452);
or U19627 (N_19627,N_19543,N_19504);
or U19628 (N_19628,N_19564,N_19464);
or U19629 (N_19629,N_19570,N_19478);
nand U19630 (N_19630,N_19534,N_19420);
and U19631 (N_19631,N_19584,N_19526);
nand U19632 (N_19632,N_19445,N_19476);
nand U19633 (N_19633,N_19563,N_19566);
or U19634 (N_19634,N_19473,N_19589);
nand U19635 (N_19635,N_19567,N_19451);
or U19636 (N_19636,N_19560,N_19568);
and U19637 (N_19637,N_19416,N_19592);
and U19638 (N_19638,N_19410,N_19421);
nand U19639 (N_19639,N_19457,N_19523);
and U19640 (N_19640,N_19438,N_19553);
nand U19641 (N_19641,N_19407,N_19486);
nor U19642 (N_19642,N_19491,N_19472);
or U19643 (N_19643,N_19511,N_19479);
nor U19644 (N_19644,N_19513,N_19450);
or U19645 (N_19645,N_19490,N_19540);
nor U19646 (N_19646,N_19520,N_19498);
nand U19647 (N_19647,N_19492,N_19548);
nor U19648 (N_19648,N_19524,N_19459);
and U19649 (N_19649,N_19593,N_19550);
or U19650 (N_19650,N_19477,N_19442);
nand U19651 (N_19651,N_19509,N_19495);
nor U19652 (N_19652,N_19515,N_19433);
xnor U19653 (N_19653,N_19578,N_19458);
and U19654 (N_19654,N_19431,N_19423);
and U19655 (N_19655,N_19539,N_19585);
xor U19656 (N_19656,N_19465,N_19595);
or U19657 (N_19657,N_19530,N_19470);
nor U19658 (N_19658,N_19535,N_19537);
and U19659 (N_19659,N_19521,N_19552);
xnor U19660 (N_19660,N_19455,N_19525);
nor U19661 (N_19661,N_19546,N_19444);
or U19662 (N_19662,N_19497,N_19528);
and U19663 (N_19663,N_19531,N_19555);
and U19664 (N_19664,N_19481,N_19432);
nor U19665 (N_19665,N_19599,N_19573);
and U19666 (N_19666,N_19430,N_19591);
xor U19667 (N_19667,N_19594,N_19512);
and U19668 (N_19668,N_19405,N_19463);
xor U19669 (N_19669,N_19514,N_19453);
or U19670 (N_19670,N_19574,N_19415);
xor U19671 (N_19671,N_19561,N_19429);
xor U19672 (N_19672,N_19572,N_19569);
xnor U19673 (N_19673,N_19422,N_19427);
xor U19674 (N_19674,N_19482,N_19527);
xnor U19675 (N_19675,N_19556,N_19425);
nor U19676 (N_19676,N_19454,N_19461);
or U19677 (N_19677,N_19435,N_19579);
nor U19678 (N_19678,N_19532,N_19456);
or U19679 (N_19679,N_19462,N_19484);
xnor U19680 (N_19680,N_19518,N_19506);
nor U19681 (N_19681,N_19483,N_19557);
xnor U19682 (N_19682,N_19418,N_19408);
or U19683 (N_19683,N_19559,N_19403);
and U19684 (N_19684,N_19510,N_19447);
xnor U19685 (N_19685,N_19533,N_19443);
nor U19686 (N_19686,N_19488,N_19587);
nand U19687 (N_19687,N_19437,N_19480);
or U19688 (N_19688,N_19401,N_19489);
xnor U19689 (N_19689,N_19500,N_19496);
and U19690 (N_19690,N_19409,N_19576);
nor U19691 (N_19691,N_19597,N_19508);
xor U19692 (N_19692,N_19502,N_19580);
nor U19693 (N_19693,N_19475,N_19598);
nand U19694 (N_19694,N_19536,N_19440);
and U19695 (N_19695,N_19558,N_19549);
and U19696 (N_19696,N_19471,N_19551);
and U19697 (N_19697,N_19545,N_19517);
or U19698 (N_19698,N_19547,N_19494);
nand U19699 (N_19699,N_19439,N_19419);
xnor U19700 (N_19700,N_19446,N_19559);
nor U19701 (N_19701,N_19588,N_19471);
xor U19702 (N_19702,N_19559,N_19414);
nand U19703 (N_19703,N_19463,N_19591);
and U19704 (N_19704,N_19561,N_19423);
and U19705 (N_19705,N_19444,N_19564);
xor U19706 (N_19706,N_19515,N_19535);
and U19707 (N_19707,N_19566,N_19554);
and U19708 (N_19708,N_19542,N_19463);
and U19709 (N_19709,N_19419,N_19471);
and U19710 (N_19710,N_19592,N_19587);
and U19711 (N_19711,N_19549,N_19489);
xor U19712 (N_19712,N_19514,N_19447);
xnor U19713 (N_19713,N_19445,N_19414);
nor U19714 (N_19714,N_19411,N_19563);
nand U19715 (N_19715,N_19529,N_19589);
xnor U19716 (N_19716,N_19578,N_19476);
and U19717 (N_19717,N_19417,N_19423);
nand U19718 (N_19718,N_19402,N_19416);
nor U19719 (N_19719,N_19471,N_19478);
or U19720 (N_19720,N_19550,N_19451);
xor U19721 (N_19721,N_19539,N_19424);
or U19722 (N_19722,N_19586,N_19565);
nor U19723 (N_19723,N_19515,N_19494);
or U19724 (N_19724,N_19565,N_19553);
or U19725 (N_19725,N_19514,N_19437);
xnor U19726 (N_19726,N_19467,N_19500);
xor U19727 (N_19727,N_19484,N_19548);
and U19728 (N_19728,N_19550,N_19598);
nand U19729 (N_19729,N_19440,N_19554);
nand U19730 (N_19730,N_19527,N_19471);
or U19731 (N_19731,N_19481,N_19419);
nor U19732 (N_19732,N_19472,N_19444);
and U19733 (N_19733,N_19528,N_19562);
xnor U19734 (N_19734,N_19474,N_19586);
and U19735 (N_19735,N_19453,N_19558);
nor U19736 (N_19736,N_19596,N_19541);
xnor U19737 (N_19737,N_19507,N_19448);
nor U19738 (N_19738,N_19442,N_19429);
nand U19739 (N_19739,N_19450,N_19444);
nor U19740 (N_19740,N_19485,N_19425);
or U19741 (N_19741,N_19480,N_19421);
and U19742 (N_19742,N_19420,N_19463);
or U19743 (N_19743,N_19592,N_19511);
nor U19744 (N_19744,N_19541,N_19416);
nor U19745 (N_19745,N_19477,N_19505);
nor U19746 (N_19746,N_19514,N_19402);
nor U19747 (N_19747,N_19593,N_19432);
and U19748 (N_19748,N_19589,N_19584);
or U19749 (N_19749,N_19462,N_19565);
nand U19750 (N_19750,N_19411,N_19587);
nor U19751 (N_19751,N_19441,N_19595);
or U19752 (N_19752,N_19545,N_19419);
or U19753 (N_19753,N_19524,N_19549);
xor U19754 (N_19754,N_19419,N_19445);
nand U19755 (N_19755,N_19418,N_19546);
and U19756 (N_19756,N_19413,N_19561);
and U19757 (N_19757,N_19507,N_19548);
xnor U19758 (N_19758,N_19524,N_19485);
nand U19759 (N_19759,N_19413,N_19556);
nor U19760 (N_19760,N_19529,N_19544);
or U19761 (N_19761,N_19469,N_19487);
nor U19762 (N_19762,N_19589,N_19568);
nor U19763 (N_19763,N_19450,N_19586);
or U19764 (N_19764,N_19469,N_19468);
and U19765 (N_19765,N_19507,N_19458);
and U19766 (N_19766,N_19599,N_19477);
or U19767 (N_19767,N_19556,N_19460);
xor U19768 (N_19768,N_19409,N_19418);
and U19769 (N_19769,N_19481,N_19479);
nand U19770 (N_19770,N_19595,N_19566);
or U19771 (N_19771,N_19549,N_19468);
or U19772 (N_19772,N_19482,N_19444);
or U19773 (N_19773,N_19461,N_19563);
or U19774 (N_19774,N_19526,N_19446);
and U19775 (N_19775,N_19562,N_19555);
xnor U19776 (N_19776,N_19410,N_19560);
or U19777 (N_19777,N_19458,N_19430);
nor U19778 (N_19778,N_19507,N_19533);
xnor U19779 (N_19779,N_19597,N_19515);
nand U19780 (N_19780,N_19562,N_19416);
xnor U19781 (N_19781,N_19410,N_19514);
and U19782 (N_19782,N_19431,N_19469);
nand U19783 (N_19783,N_19558,N_19482);
or U19784 (N_19784,N_19475,N_19599);
xnor U19785 (N_19785,N_19478,N_19550);
or U19786 (N_19786,N_19408,N_19412);
and U19787 (N_19787,N_19402,N_19512);
nand U19788 (N_19788,N_19562,N_19496);
or U19789 (N_19789,N_19457,N_19404);
nand U19790 (N_19790,N_19526,N_19457);
xnor U19791 (N_19791,N_19572,N_19594);
nand U19792 (N_19792,N_19562,N_19594);
or U19793 (N_19793,N_19503,N_19583);
xnor U19794 (N_19794,N_19436,N_19548);
nand U19795 (N_19795,N_19453,N_19461);
nor U19796 (N_19796,N_19594,N_19519);
and U19797 (N_19797,N_19588,N_19578);
and U19798 (N_19798,N_19558,N_19468);
or U19799 (N_19799,N_19593,N_19412);
nand U19800 (N_19800,N_19638,N_19746);
and U19801 (N_19801,N_19753,N_19668);
and U19802 (N_19802,N_19773,N_19780);
and U19803 (N_19803,N_19777,N_19616);
nor U19804 (N_19804,N_19692,N_19664);
nand U19805 (N_19805,N_19715,N_19767);
or U19806 (N_19806,N_19645,N_19614);
and U19807 (N_19807,N_19649,N_19755);
xnor U19808 (N_19808,N_19737,N_19627);
or U19809 (N_19809,N_19681,N_19740);
xor U19810 (N_19810,N_19702,N_19685);
nor U19811 (N_19811,N_19726,N_19640);
and U19812 (N_19812,N_19723,N_19717);
or U19813 (N_19813,N_19673,N_19701);
or U19814 (N_19814,N_19760,N_19724);
nor U19815 (N_19815,N_19678,N_19743);
and U19816 (N_19816,N_19725,N_19789);
nand U19817 (N_19817,N_19675,N_19629);
nor U19818 (N_19818,N_19601,N_19646);
nand U19819 (N_19819,N_19669,N_19766);
or U19820 (N_19820,N_19759,N_19618);
nand U19821 (N_19821,N_19720,N_19697);
nand U19822 (N_19822,N_19729,N_19703);
and U19823 (N_19823,N_19748,N_19710);
nor U19824 (N_19824,N_19632,N_19796);
nor U19825 (N_19825,N_19736,N_19786);
and U19826 (N_19826,N_19612,N_19644);
xnor U19827 (N_19827,N_19744,N_19642);
nor U19828 (N_19828,N_19651,N_19750);
nor U19829 (N_19829,N_19713,N_19624);
nand U19830 (N_19830,N_19648,N_19738);
xnor U19831 (N_19831,N_19747,N_19658);
xnor U19832 (N_19832,N_19680,N_19781);
and U19833 (N_19833,N_19667,N_19652);
xor U19834 (N_19834,N_19636,N_19719);
and U19835 (N_19835,N_19783,N_19609);
or U19836 (N_19836,N_19765,N_19660);
nand U19837 (N_19837,N_19635,N_19634);
or U19838 (N_19838,N_19730,N_19684);
and U19839 (N_19839,N_19734,N_19615);
or U19840 (N_19840,N_19787,N_19788);
and U19841 (N_19841,N_19798,N_19631);
xnor U19842 (N_19842,N_19661,N_19745);
or U19843 (N_19843,N_19700,N_19792);
nand U19844 (N_19844,N_19695,N_19683);
xnor U19845 (N_19845,N_19693,N_19791);
xnor U19846 (N_19846,N_19769,N_19778);
xor U19847 (N_19847,N_19672,N_19705);
or U19848 (N_19848,N_19727,N_19770);
xnor U19849 (N_19849,N_19604,N_19785);
or U19850 (N_19850,N_19714,N_19757);
and U19851 (N_19851,N_19756,N_19674);
xor U19852 (N_19852,N_19718,N_19690);
nor U19853 (N_19853,N_19763,N_19602);
and U19854 (N_19854,N_19613,N_19768);
xor U19855 (N_19855,N_19622,N_19682);
nand U19856 (N_19856,N_19775,N_19784);
or U19857 (N_19857,N_19731,N_19637);
or U19858 (N_19858,N_19607,N_19626);
or U19859 (N_19859,N_19721,N_19709);
or U19860 (N_19860,N_19790,N_19732);
nand U19861 (N_19861,N_19691,N_19774);
nand U19862 (N_19862,N_19625,N_19694);
nand U19863 (N_19863,N_19620,N_19610);
nand U19864 (N_19864,N_19733,N_19686);
nor U19865 (N_19865,N_19706,N_19716);
or U19866 (N_19866,N_19742,N_19799);
or U19867 (N_19867,N_19647,N_19679);
and U19868 (N_19868,N_19722,N_19741);
nand U19869 (N_19869,N_19671,N_19657);
and U19870 (N_19870,N_19762,N_19670);
or U19871 (N_19871,N_19689,N_19643);
xnor U19872 (N_19872,N_19779,N_19603);
nor U19873 (N_19873,N_19782,N_19655);
nor U19874 (N_19874,N_19608,N_19739);
nor U19875 (N_19875,N_19630,N_19628);
and U19876 (N_19876,N_19621,N_19605);
or U19877 (N_19877,N_19617,N_19600);
nor U19878 (N_19878,N_19707,N_19676);
or U19879 (N_19879,N_19711,N_19653);
xnor U19880 (N_19880,N_19797,N_19698);
nand U19881 (N_19881,N_19662,N_19654);
nor U19882 (N_19882,N_19656,N_19639);
and U19883 (N_19883,N_19665,N_19699);
and U19884 (N_19884,N_19677,N_19696);
nand U19885 (N_19885,N_19751,N_19761);
nor U19886 (N_19886,N_19633,N_19772);
nand U19887 (N_19887,N_19793,N_19666);
and U19888 (N_19888,N_19735,N_19764);
or U19889 (N_19889,N_19619,N_19728);
xor U19890 (N_19890,N_19611,N_19758);
nand U19891 (N_19891,N_19687,N_19795);
or U19892 (N_19892,N_19704,N_19776);
nand U19893 (N_19893,N_19663,N_19794);
nor U19894 (N_19894,N_19623,N_19771);
nor U19895 (N_19895,N_19752,N_19659);
xnor U19896 (N_19896,N_19688,N_19606);
and U19897 (N_19897,N_19754,N_19749);
nor U19898 (N_19898,N_19712,N_19641);
and U19899 (N_19899,N_19650,N_19708);
or U19900 (N_19900,N_19617,N_19669);
nor U19901 (N_19901,N_19671,N_19686);
nor U19902 (N_19902,N_19675,N_19710);
xor U19903 (N_19903,N_19713,N_19777);
and U19904 (N_19904,N_19774,N_19636);
or U19905 (N_19905,N_19774,N_19662);
and U19906 (N_19906,N_19736,N_19793);
or U19907 (N_19907,N_19736,N_19711);
and U19908 (N_19908,N_19664,N_19694);
nor U19909 (N_19909,N_19641,N_19646);
or U19910 (N_19910,N_19752,N_19704);
or U19911 (N_19911,N_19666,N_19763);
xnor U19912 (N_19912,N_19753,N_19655);
nand U19913 (N_19913,N_19645,N_19693);
and U19914 (N_19914,N_19736,N_19762);
nand U19915 (N_19915,N_19701,N_19601);
nor U19916 (N_19916,N_19764,N_19775);
and U19917 (N_19917,N_19783,N_19664);
nand U19918 (N_19918,N_19606,N_19660);
xnor U19919 (N_19919,N_19648,N_19673);
xor U19920 (N_19920,N_19751,N_19679);
xor U19921 (N_19921,N_19744,N_19673);
nor U19922 (N_19922,N_19622,N_19747);
nor U19923 (N_19923,N_19672,N_19655);
xor U19924 (N_19924,N_19646,N_19621);
nor U19925 (N_19925,N_19656,N_19676);
nand U19926 (N_19926,N_19712,N_19770);
or U19927 (N_19927,N_19726,N_19670);
nor U19928 (N_19928,N_19635,N_19626);
nand U19929 (N_19929,N_19609,N_19666);
and U19930 (N_19930,N_19635,N_19723);
nand U19931 (N_19931,N_19745,N_19711);
xnor U19932 (N_19932,N_19691,N_19619);
xnor U19933 (N_19933,N_19654,N_19616);
or U19934 (N_19934,N_19784,N_19680);
or U19935 (N_19935,N_19705,N_19670);
and U19936 (N_19936,N_19719,N_19664);
nor U19937 (N_19937,N_19688,N_19737);
nor U19938 (N_19938,N_19789,N_19620);
and U19939 (N_19939,N_19731,N_19675);
nor U19940 (N_19940,N_19787,N_19647);
nor U19941 (N_19941,N_19728,N_19713);
or U19942 (N_19942,N_19792,N_19693);
nand U19943 (N_19943,N_19638,N_19647);
xnor U19944 (N_19944,N_19770,N_19741);
or U19945 (N_19945,N_19652,N_19706);
nand U19946 (N_19946,N_19762,N_19763);
nor U19947 (N_19947,N_19684,N_19617);
nand U19948 (N_19948,N_19682,N_19651);
and U19949 (N_19949,N_19624,N_19616);
nand U19950 (N_19950,N_19741,N_19736);
xor U19951 (N_19951,N_19621,N_19780);
or U19952 (N_19952,N_19779,N_19793);
xor U19953 (N_19953,N_19778,N_19688);
nand U19954 (N_19954,N_19672,N_19636);
and U19955 (N_19955,N_19781,N_19704);
and U19956 (N_19956,N_19647,N_19674);
and U19957 (N_19957,N_19679,N_19716);
nor U19958 (N_19958,N_19716,N_19695);
xor U19959 (N_19959,N_19730,N_19708);
xnor U19960 (N_19960,N_19648,N_19751);
xor U19961 (N_19961,N_19757,N_19608);
nand U19962 (N_19962,N_19668,N_19734);
and U19963 (N_19963,N_19630,N_19712);
or U19964 (N_19964,N_19639,N_19777);
and U19965 (N_19965,N_19714,N_19652);
or U19966 (N_19966,N_19632,N_19669);
nor U19967 (N_19967,N_19601,N_19763);
nand U19968 (N_19968,N_19783,N_19733);
and U19969 (N_19969,N_19675,N_19681);
and U19970 (N_19970,N_19673,N_19776);
or U19971 (N_19971,N_19690,N_19717);
or U19972 (N_19972,N_19748,N_19609);
xor U19973 (N_19973,N_19673,N_19740);
nand U19974 (N_19974,N_19683,N_19747);
and U19975 (N_19975,N_19760,N_19669);
and U19976 (N_19976,N_19780,N_19748);
or U19977 (N_19977,N_19701,N_19631);
nor U19978 (N_19978,N_19791,N_19644);
xnor U19979 (N_19979,N_19650,N_19795);
nand U19980 (N_19980,N_19628,N_19663);
and U19981 (N_19981,N_19638,N_19653);
and U19982 (N_19982,N_19712,N_19797);
nand U19983 (N_19983,N_19606,N_19690);
nand U19984 (N_19984,N_19769,N_19691);
or U19985 (N_19985,N_19696,N_19685);
nor U19986 (N_19986,N_19681,N_19625);
or U19987 (N_19987,N_19693,N_19673);
xor U19988 (N_19988,N_19740,N_19662);
and U19989 (N_19989,N_19746,N_19680);
nand U19990 (N_19990,N_19612,N_19618);
and U19991 (N_19991,N_19672,N_19676);
nor U19992 (N_19992,N_19639,N_19754);
and U19993 (N_19993,N_19681,N_19786);
nand U19994 (N_19994,N_19745,N_19682);
nand U19995 (N_19995,N_19745,N_19724);
nand U19996 (N_19996,N_19681,N_19622);
or U19997 (N_19997,N_19707,N_19614);
or U19998 (N_19998,N_19773,N_19646);
nor U19999 (N_19999,N_19682,N_19722);
or U20000 (N_20000,N_19933,N_19935);
or U20001 (N_20001,N_19838,N_19904);
xor U20002 (N_20002,N_19816,N_19824);
nand U20003 (N_20003,N_19869,N_19919);
xor U20004 (N_20004,N_19993,N_19922);
xor U20005 (N_20005,N_19975,N_19952);
nand U20006 (N_20006,N_19971,N_19827);
and U20007 (N_20007,N_19887,N_19808);
and U20008 (N_20008,N_19804,N_19830);
nand U20009 (N_20009,N_19999,N_19888);
and U20010 (N_20010,N_19940,N_19985);
and U20011 (N_20011,N_19848,N_19944);
nand U20012 (N_20012,N_19981,N_19989);
and U20013 (N_20013,N_19906,N_19964);
or U20014 (N_20014,N_19883,N_19941);
nand U20015 (N_20015,N_19959,N_19942);
nor U20016 (N_20016,N_19949,N_19937);
and U20017 (N_20017,N_19801,N_19862);
nor U20018 (N_20018,N_19832,N_19965);
or U20019 (N_20019,N_19820,N_19884);
nor U20020 (N_20020,N_19834,N_19910);
nor U20021 (N_20021,N_19846,N_19899);
nor U20022 (N_20022,N_19903,N_19923);
or U20023 (N_20023,N_19995,N_19998);
or U20024 (N_20024,N_19802,N_19874);
or U20025 (N_20025,N_19864,N_19877);
or U20026 (N_20026,N_19889,N_19875);
nor U20027 (N_20027,N_19852,N_19870);
nor U20028 (N_20028,N_19882,N_19853);
nand U20029 (N_20029,N_19980,N_19977);
nor U20030 (N_20030,N_19924,N_19831);
xor U20031 (N_20031,N_19990,N_19991);
nand U20032 (N_20032,N_19909,N_19894);
and U20033 (N_20033,N_19900,N_19913);
and U20034 (N_20034,N_19920,N_19974);
xnor U20035 (N_20035,N_19876,N_19836);
xnor U20036 (N_20036,N_19898,N_19847);
and U20037 (N_20037,N_19982,N_19945);
nand U20038 (N_20038,N_19851,N_19837);
xnor U20039 (N_20039,N_19955,N_19916);
xnor U20040 (N_20040,N_19936,N_19907);
and U20041 (N_20041,N_19918,N_19973);
nor U20042 (N_20042,N_19967,N_19994);
nand U20043 (N_20043,N_19806,N_19826);
xor U20044 (N_20044,N_19809,N_19871);
and U20045 (N_20045,N_19868,N_19925);
nand U20046 (N_20046,N_19844,N_19934);
nand U20047 (N_20047,N_19835,N_19926);
xnor U20048 (N_20048,N_19842,N_19885);
nor U20049 (N_20049,N_19823,N_19912);
or U20050 (N_20050,N_19893,N_19954);
and U20051 (N_20051,N_19992,N_19976);
or U20052 (N_20052,N_19839,N_19818);
xor U20053 (N_20053,N_19896,N_19908);
xnor U20054 (N_20054,N_19891,N_19927);
xor U20055 (N_20055,N_19921,N_19931);
or U20056 (N_20056,N_19911,N_19929);
xor U20057 (N_20057,N_19962,N_19895);
nor U20058 (N_20058,N_19857,N_19860);
and U20059 (N_20059,N_19953,N_19939);
nand U20060 (N_20060,N_19960,N_19833);
xnor U20061 (N_20061,N_19829,N_19983);
or U20062 (N_20062,N_19886,N_19880);
and U20063 (N_20063,N_19805,N_19812);
nor U20064 (N_20064,N_19822,N_19890);
or U20065 (N_20065,N_19845,N_19956);
xor U20066 (N_20066,N_19996,N_19803);
xnor U20067 (N_20067,N_19873,N_19854);
xnor U20068 (N_20068,N_19800,N_19849);
nand U20069 (N_20069,N_19969,N_19855);
nand U20070 (N_20070,N_19810,N_19872);
or U20071 (N_20071,N_19950,N_19859);
or U20072 (N_20072,N_19958,N_19867);
or U20073 (N_20073,N_19951,N_19963);
or U20074 (N_20074,N_19861,N_19914);
and U20075 (N_20075,N_19879,N_19984);
and U20076 (N_20076,N_19828,N_19881);
and U20077 (N_20077,N_19817,N_19856);
and U20078 (N_20078,N_19815,N_19957);
xor U20079 (N_20079,N_19972,N_19840);
nor U20080 (N_20080,N_19970,N_19947);
xnor U20081 (N_20081,N_19821,N_19930);
and U20082 (N_20082,N_19814,N_19988);
or U20083 (N_20083,N_19902,N_19915);
or U20084 (N_20084,N_19946,N_19978);
and U20085 (N_20085,N_19948,N_19938);
nor U20086 (N_20086,N_19850,N_19905);
and U20087 (N_20087,N_19997,N_19863);
nor U20088 (N_20088,N_19917,N_19901);
or U20089 (N_20089,N_19807,N_19858);
and U20090 (N_20090,N_19966,N_19841);
or U20091 (N_20091,N_19811,N_19813);
and U20092 (N_20092,N_19843,N_19892);
nor U20093 (N_20093,N_19819,N_19897);
xnor U20094 (N_20094,N_19932,N_19987);
and U20095 (N_20095,N_19825,N_19866);
nand U20096 (N_20096,N_19968,N_19979);
nand U20097 (N_20097,N_19943,N_19865);
or U20098 (N_20098,N_19986,N_19928);
nand U20099 (N_20099,N_19961,N_19878);
nor U20100 (N_20100,N_19872,N_19827);
nand U20101 (N_20101,N_19916,N_19875);
xor U20102 (N_20102,N_19821,N_19938);
and U20103 (N_20103,N_19867,N_19911);
or U20104 (N_20104,N_19996,N_19928);
or U20105 (N_20105,N_19925,N_19824);
nor U20106 (N_20106,N_19911,N_19992);
and U20107 (N_20107,N_19970,N_19889);
nor U20108 (N_20108,N_19967,N_19804);
nand U20109 (N_20109,N_19963,N_19897);
and U20110 (N_20110,N_19902,N_19886);
and U20111 (N_20111,N_19905,N_19887);
nand U20112 (N_20112,N_19822,N_19895);
nand U20113 (N_20113,N_19852,N_19869);
xnor U20114 (N_20114,N_19984,N_19913);
xnor U20115 (N_20115,N_19939,N_19856);
and U20116 (N_20116,N_19910,N_19829);
nor U20117 (N_20117,N_19811,N_19844);
nand U20118 (N_20118,N_19897,N_19875);
or U20119 (N_20119,N_19902,N_19866);
xnor U20120 (N_20120,N_19845,N_19911);
nor U20121 (N_20121,N_19864,N_19894);
xnor U20122 (N_20122,N_19873,N_19830);
nor U20123 (N_20123,N_19906,N_19983);
nor U20124 (N_20124,N_19939,N_19834);
and U20125 (N_20125,N_19902,N_19867);
nor U20126 (N_20126,N_19874,N_19840);
and U20127 (N_20127,N_19987,N_19973);
or U20128 (N_20128,N_19883,N_19927);
or U20129 (N_20129,N_19803,N_19868);
and U20130 (N_20130,N_19939,N_19882);
xor U20131 (N_20131,N_19981,N_19886);
or U20132 (N_20132,N_19871,N_19936);
nor U20133 (N_20133,N_19861,N_19875);
nor U20134 (N_20134,N_19866,N_19820);
nor U20135 (N_20135,N_19964,N_19978);
xor U20136 (N_20136,N_19854,N_19897);
xnor U20137 (N_20137,N_19904,N_19923);
nand U20138 (N_20138,N_19880,N_19970);
xnor U20139 (N_20139,N_19927,N_19893);
nor U20140 (N_20140,N_19812,N_19928);
nand U20141 (N_20141,N_19974,N_19924);
nand U20142 (N_20142,N_19849,N_19975);
nand U20143 (N_20143,N_19810,N_19992);
and U20144 (N_20144,N_19873,N_19898);
or U20145 (N_20145,N_19863,N_19964);
xnor U20146 (N_20146,N_19988,N_19885);
nand U20147 (N_20147,N_19920,N_19851);
and U20148 (N_20148,N_19897,N_19879);
xnor U20149 (N_20149,N_19809,N_19999);
nor U20150 (N_20150,N_19826,N_19973);
nand U20151 (N_20151,N_19874,N_19940);
or U20152 (N_20152,N_19810,N_19842);
or U20153 (N_20153,N_19818,N_19813);
and U20154 (N_20154,N_19847,N_19950);
and U20155 (N_20155,N_19867,N_19907);
and U20156 (N_20156,N_19987,N_19902);
xnor U20157 (N_20157,N_19959,N_19860);
and U20158 (N_20158,N_19898,N_19964);
or U20159 (N_20159,N_19872,N_19966);
nor U20160 (N_20160,N_19926,N_19932);
or U20161 (N_20161,N_19879,N_19927);
nor U20162 (N_20162,N_19915,N_19850);
and U20163 (N_20163,N_19990,N_19829);
nor U20164 (N_20164,N_19959,N_19940);
xor U20165 (N_20165,N_19906,N_19939);
nand U20166 (N_20166,N_19819,N_19999);
and U20167 (N_20167,N_19929,N_19875);
or U20168 (N_20168,N_19933,N_19874);
and U20169 (N_20169,N_19870,N_19987);
xor U20170 (N_20170,N_19927,N_19860);
and U20171 (N_20171,N_19816,N_19976);
and U20172 (N_20172,N_19944,N_19809);
nor U20173 (N_20173,N_19905,N_19875);
and U20174 (N_20174,N_19807,N_19801);
and U20175 (N_20175,N_19948,N_19929);
nand U20176 (N_20176,N_19823,N_19859);
nand U20177 (N_20177,N_19808,N_19998);
nand U20178 (N_20178,N_19862,N_19833);
xor U20179 (N_20179,N_19846,N_19814);
and U20180 (N_20180,N_19907,N_19926);
and U20181 (N_20181,N_19949,N_19955);
and U20182 (N_20182,N_19891,N_19803);
nor U20183 (N_20183,N_19824,N_19836);
xor U20184 (N_20184,N_19829,N_19988);
or U20185 (N_20185,N_19851,N_19830);
nor U20186 (N_20186,N_19864,N_19911);
xnor U20187 (N_20187,N_19974,N_19933);
or U20188 (N_20188,N_19891,N_19882);
or U20189 (N_20189,N_19920,N_19838);
or U20190 (N_20190,N_19845,N_19995);
xnor U20191 (N_20191,N_19873,N_19872);
and U20192 (N_20192,N_19933,N_19924);
xnor U20193 (N_20193,N_19868,N_19995);
xor U20194 (N_20194,N_19899,N_19858);
and U20195 (N_20195,N_19973,N_19959);
xnor U20196 (N_20196,N_19901,N_19891);
xnor U20197 (N_20197,N_19843,N_19820);
xor U20198 (N_20198,N_19911,N_19922);
nor U20199 (N_20199,N_19835,N_19986);
xor U20200 (N_20200,N_20174,N_20061);
nor U20201 (N_20201,N_20084,N_20197);
and U20202 (N_20202,N_20079,N_20078);
and U20203 (N_20203,N_20111,N_20124);
or U20204 (N_20204,N_20037,N_20004);
nand U20205 (N_20205,N_20170,N_20137);
xor U20206 (N_20206,N_20067,N_20009);
or U20207 (N_20207,N_20114,N_20194);
nor U20208 (N_20208,N_20085,N_20002);
nand U20209 (N_20209,N_20158,N_20049);
nor U20210 (N_20210,N_20048,N_20044);
xor U20211 (N_20211,N_20108,N_20083);
xor U20212 (N_20212,N_20028,N_20157);
nor U20213 (N_20213,N_20077,N_20099);
or U20214 (N_20214,N_20155,N_20125);
nor U20215 (N_20215,N_20035,N_20193);
and U20216 (N_20216,N_20101,N_20154);
and U20217 (N_20217,N_20071,N_20039);
nand U20218 (N_20218,N_20090,N_20107);
xnor U20219 (N_20219,N_20014,N_20102);
nand U20220 (N_20220,N_20054,N_20179);
nor U20221 (N_20221,N_20198,N_20142);
and U20222 (N_20222,N_20092,N_20056);
xor U20223 (N_20223,N_20177,N_20057);
or U20224 (N_20224,N_20116,N_20168);
xnor U20225 (N_20225,N_20191,N_20171);
and U20226 (N_20226,N_20058,N_20143);
xor U20227 (N_20227,N_20165,N_20173);
xnor U20228 (N_20228,N_20105,N_20086);
nand U20229 (N_20229,N_20192,N_20022);
and U20230 (N_20230,N_20074,N_20120);
xnor U20231 (N_20231,N_20066,N_20118);
nor U20232 (N_20232,N_20189,N_20036);
or U20233 (N_20233,N_20127,N_20095);
nor U20234 (N_20234,N_20041,N_20182);
nor U20235 (N_20235,N_20091,N_20152);
and U20236 (N_20236,N_20115,N_20062);
or U20237 (N_20237,N_20199,N_20013);
xor U20238 (N_20238,N_20073,N_20075);
and U20239 (N_20239,N_20126,N_20010);
xor U20240 (N_20240,N_20055,N_20060);
xnor U20241 (N_20241,N_20052,N_20151);
and U20242 (N_20242,N_20025,N_20065);
nand U20243 (N_20243,N_20141,N_20008);
nand U20244 (N_20244,N_20130,N_20007);
and U20245 (N_20245,N_20129,N_20017);
xnor U20246 (N_20246,N_20006,N_20001);
nor U20247 (N_20247,N_20185,N_20082);
or U20248 (N_20248,N_20160,N_20123);
xor U20249 (N_20249,N_20087,N_20138);
or U20250 (N_20250,N_20180,N_20181);
nand U20251 (N_20251,N_20100,N_20146);
xnor U20252 (N_20252,N_20163,N_20104);
nor U20253 (N_20253,N_20021,N_20110);
nor U20254 (N_20254,N_20148,N_20106);
nand U20255 (N_20255,N_20183,N_20135);
and U20256 (N_20256,N_20196,N_20068);
or U20257 (N_20257,N_20038,N_20018);
nand U20258 (N_20258,N_20005,N_20015);
and U20259 (N_20259,N_20011,N_20136);
and U20260 (N_20260,N_20169,N_20132);
and U20261 (N_20261,N_20081,N_20093);
or U20262 (N_20262,N_20033,N_20139);
xor U20263 (N_20263,N_20166,N_20023);
or U20264 (N_20264,N_20153,N_20134);
or U20265 (N_20265,N_20051,N_20190);
and U20266 (N_20266,N_20053,N_20150);
xor U20267 (N_20267,N_20043,N_20156);
nand U20268 (N_20268,N_20031,N_20059);
nor U20269 (N_20269,N_20050,N_20188);
nor U20270 (N_20270,N_20167,N_20186);
xnor U20271 (N_20271,N_20128,N_20072);
nand U20272 (N_20272,N_20133,N_20187);
and U20273 (N_20273,N_20076,N_20119);
or U20274 (N_20274,N_20042,N_20089);
nor U20275 (N_20275,N_20145,N_20103);
and U20276 (N_20276,N_20029,N_20000);
xor U20277 (N_20277,N_20027,N_20034);
nor U20278 (N_20278,N_20140,N_20178);
or U20279 (N_20279,N_20024,N_20117);
nand U20280 (N_20280,N_20080,N_20047);
nand U20281 (N_20281,N_20063,N_20122);
and U20282 (N_20282,N_20069,N_20159);
or U20283 (N_20283,N_20112,N_20045);
xnor U20284 (N_20284,N_20070,N_20184);
xor U20285 (N_20285,N_20149,N_20088);
and U20286 (N_20286,N_20176,N_20162);
nor U20287 (N_20287,N_20109,N_20161);
or U20288 (N_20288,N_20164,N_20003);
nand U20289 (N_20289,N_20030,N_20121);
nand U20290 (N_20290,N_20131,N_20113);
nand U20291 (N_20291,N_20147,N_20026);
nor U20292 (N_20292,N_20064,N_20144);
nor U20293 (N_20293,N_20020,N_20016);
nor U20294 (N_20294,N_20040,N_20097);
and U20295 (N_20295,N_20175,N_20172);
nand U20296 (N_20296,N_20012,N_20046);
and U20297 (N_20297,N_20096,N_20094);
or U20298 (N_20298,N_20195,N_20019);
xnor U20299 (N_20299,N_20032,N_20098);
xnor U20300 (N_20300,N_20097,N_20157);
xor U20301 (N_20301,N_20120,N_20141);
xnor U20302 (N_20302,N_20099,N_20149);
nor U20303 (N_20303,N_20133,N_20059);
and U20304 (N_20304,N_20171,N_20126);
nand U20305 (N_20305,N_20044,N_20196);
nand U20306 (N_20306,N_20198,N_20003);
or U20307 (N_20307,N_20046,N_20166);
xnor U20308 (N_20308,N_20124,N_20168);
xnor U20309 (N_20309,N_20107,N_20161);
or U20310 (N_20310,N_20029,N_20005);
and U20311 (N_20311,N_20172,N_20180);
and U20312 (N_20312,N_20099,N_20052);
nand U20313 (N_20313,N_20028,N_20061);
nand U20314 (N_20314,N_20023,N_20177);
nor U20315 (N_20315,N_20133,N_20065);
and U20316 (N_20316,N_20075,N_20030);
or U20317 (N_20317,N_20132,N_20190);
xnor U20318 (N_20318,N_20057,N_20001);
or U20319 (N_20319,N_20069,N_20043);
or U20320 (N_20320,N_20012,N_20111);
nand U20321 (N_20321,N_20056,N_20148);
nand U20322 (N_20322,N_20140,N_20032);
nor U20323 (N_20323,N_20031,N_20052);
nand U20324 (N_20324,N_20006,N_20061);
or U20325 (N_20325,N_20091,N_20121);
xor U20326 (N_20326,N_20183,N_20176);
nand U20327 (N_20327,N_20161,N_20146);
nand U20328 (N_20328,N_20073,N_20171);
and U20329 (N_20329,N_20162,N_20037);
or U20330 (N_20330,N_20174,N_20049);
or U20331 (N_20331,N_20082,N_20005);
nand U20332 (N_20332,N_20176,N_20170);
nand U20333 (N_20333,N_20016,N_20031);
and U20334 (N_20334,N_20065,N_20000);
nor U20335 (N_20335,N_20066,N_20133);
nand U20336 (N_20336,N_20127,N_20155);
or U20337 (N_20337,N_20056,N_20137);
or U20338 (N_20338,N_20169,N_20186);
xnor U20339 (N_20339,N_20121,N_20146);
nor U20340 (N_20340,N_20056,N_20118);
nor U20341 (N_20341,N_20140,N_20017);
nor U20342 (N_20342,N_20177,N_20106);
nor U20343 (N_20343,N_20144,N_20192);
nand U20344 (N_20344,N_20169,N_20124);
or U20345 (N_20345,N_20118,N_20188);
or U20346 (N_20346,N_20005,N_20076);
nor U20347 (N_20347,N_20057,N_20098);
or U20348 (N_20348,N_20129,N_20187);
nand U20349 (N_20349,N_20158,N_20003);
nand U20350 (N_20350,N_20023,N_20100);
xor U20351 (N_20351,N_20116,N_20120);
and U20352 (N_20352,N_20108,N_20127);
nor U20353 (N_20353,N_20190,N_20112);
nor U20354 (N_20354,N_20001,N_20003);
nor U20355 (N_20355,N_20003,N_20056);
and U20356 (N_20356,N_20002,N_20176);
nand U20357 (N_20357,N_20166,N_20106);
xor U20358 (N_20358,N_20059,N_20044);
xnor U20359 (N_20359,N_20055,N_20160);
nand U20360 (N_20360,N_20132,N_20069);
nor U20361 (N_20361,N_20142,N_20104);
xor U20362 (N_20362,N_20196,N_20129);
nor U20363 (N_20363,N_20151,N_20002);
and U20364 (N_20364,N_20123,N_20135);
xnor U20365 (N_20365,N_20134,N_20035);
xor U20366 (N_20366,N_20133,N_20167);
xnor U20367 (N_20367,N_20142,N_20160);
nand U20368 (N_20368,N_20174,N_20051);
and U20369 (N_20369,N_20093,N_20083);
nor U20370 (N_20370,N_20190,N_20184);
and U20371 (N_20371,N_20053,N_20170);
xor U20372 (N_20372,N_20149,N_20043);
or U20373 (N_20373,N_20089,N_20198);
nand U20374 (N_20374,N_20179,N_20163);
or U20375 (N_20375,N_20165,N_20100);
nor U20376 (N_20376,N_20051,N_20189);
and U20377 (N_20377,N_20041,N_20158);
nor U20378 (N_20378,N_20113,N_20118);
and U20379 (N_20379,N_20043,N_20044);
xnor U20380 (N_20380,N_20110,N_20134);
and U20381 (N_20381,N_20148,N_20190);
nand U20382 (N_20382,N_20048,N_20141);
and U20383 (N_20383,N_20159,N_20134);
or U20384 (N_20384,N_20159,N_20139);
xor U20385 (N_20385,N_20006,N_20165);
nor U20386 (N_20386,N_20022,N_20182);
or U20387 (N_20387,N_20024,N_20066);
nand U20388 (N_20388,N_20190,N_20140);
or U20389 (N_20389,N_20084,N_20024);
nor U20390 (N_20390,N_20020,N_20156);
and U20391 (N_20391,N_20141,N_20137);
and U20392 (N_20392,N_20045,N_20144);
nand U20393 (N_20393,N_20002,N_20070);
xor U20394 (N_20394,N_20124,N_20146);
xnor U20395 (N_20395,N_20163,N_20170);
and U20396 (N_20396,N_20019,N_20013);
or U20397 (N_20397,N_20058,N_20189);
nand U20398 (N_20398,N_20011,N_20156);
xor U20399 (N_20399,N_20131,N_20193);
nor U20400 (N_20400,N_20282,N_20320);
xor U20401 (N_20401,N_20363,N_20350);
nand U20402 (N_20402,N_20237,N_20367);
xnor U20403 (N_20403,N_20287,N_20269);
nor U20404 (N_20404,N_20370,N_20289);
nor U20405 (N_20405,N_20330,N_20217);
nand U20406 (N_20406,N_20364,N_20303);
xor U20407 (N_20407,N_20257,N_20292);
and U20408 (N_20408,N_20377,N_20207);
nor U20409 (N_20409,N_20225,N_20349);
xor U20410 (N_20410,N_20371,N_20329);
xnor U20411 (N_20411,N_20241,N_20391);
nor U20412 (N_20412,N_20239,N_20252);
and U20413 (N_20413,N_20378,N_20212);
nor U20414 (N_20414,N_20375,N_20325);
xor U20415 (N_20415,N_20384,N_20307);
xor U20416 (N_20416,N_20392,N_20305);
xnor U20417 (N_20417,N_20357,N_20281);
nor U20418 (N_20418,N_20213,N_20343);
or U20419 (N_20419,N_20210,N_20390);
nand U20420 (N_20420,N_20273,N_20328);
xor U20421 (N_20421,N_20333,N_20355);
xnor U20422 (N_20422,N_20279,N_20206);
nand U20423 (N_20423,N_20297,N_20319);
nand U20424 (N_20424,N_20353,N_20271);
and U20425 (N_20425,N_20227,N_20288);
xnor U20426 (N_20426,N_20233,N_20242);
and U20427 (N_20427,N_20261,N_20290);
nand U20428 (N_20428,N_20395,N_20299);
and U20429 (N_20429,N_20345,N_20286);
or U20430 (N_20430,N_20321,N_20285);
xor U20431 (N_20431,N_20314,N_20276);
nor U20432 (N_20432,N_20250,N_20260);
nand U20433 (N_20433,N_20296,N_20379);
or U20434 (N_20434,N_20341,N_20201);
nand U20435 (N_20435,N_20385,N_20270);
nor U20436 (N_20436,N_20302,N_20202);
or U20437 (N_20437,N_20322,N_20246);
xor U20438 (N_20438,N_20263,N_20308);
xnor U20439 (N_20439,N_20339,N_20315);
or U20440 (N_20440,N_20300,N_20362);
nor U20441 (N_20441,N_20310,N_20266);
and U20442 (N_20442,N_20253,N_20203);
and U20443 (N_20443,N_20388,N_20389);
nand U20444 (N_20444,N_20268,N_20332);
and U20445 (N_20445,N_20346,N_20223);
nand U20446 (N_20446,N_20398,N_20244);
xor U20447 (N_20447,N_20348,N_20380);
xnor U20448 (N_20448,N_20317,N_20274);
nand U20449 (N_20449,N_20278,N_20369);
xnor U20450 (N_20450,N_20366,N_20265);
nor U20451 (N_20451,N_20262,N_20323);
or U20452 (N_20452,N_20226,N_20230);
xor U20453 (N_20453,N_20326,N_20200);
nor U20454 (N_20454,N_20272,N_20243);
and U20455 (N_20455,N_20372,N_20309);
and U20456 (N_20456,N_20208,N_20338);
and U20457 (N_20457,N_20386,N_20209);
nor U20458 (N_20458,N_20336,N_20324);
or U20459 (N_20459,N_20331,N_20373);
nand U20460 (N_20460,N_20275,N_20215);
or U20461 (N_20461,N_20220,N_20219);
nand U20462 (N_20462,N_20235,N_20354);
nor U20463 (N_20463,N_20383,N_20356);
and U20464 (N_20464,N_20259,N_20283);
nor U20465 (N_20465,N_20304,N_20358);
and U20466 (N_20466,N_20318,N_20258);
nand U20467 (N_20467,N_20365,N_20254);
or U20468 (N_20468,N_20231,N_20224);
or U20469 (N_20469,N_20337,N_20312);
xnor U20470 (N_20470,N_20236,N_20218);
nand U20471 (N_20471,N_20264,N_20301);
nand U20472 (N_20472,N_20229,N_20284);
nand U20473 (N_20473,N_20399,N_20280);
xor U20474 (N_20474,N_20311,N_20316);
nor U20475 (N_20475,N_20387,N_20238);
xor U20476 (N_20476,N_20211,N_20397);
nand U20477 (N_20477,N_20360,N_20396);
or U20478 (N_20478,N_20298,N_20361);
or U20479 (N_20479,N_20335,N_20294);
or U20480 (N_20480,N_20214,N_20327);
nand U20481 (N_20481,N_20295,N_20240);
nand U20482 (N_20482,N_20277,N_20376);
nor U20483 (N_20483,N_20313,N_20267);
or U20484 (N_20484,N_20245,N_20293);
nand U20485 (N_20485,N_20352,N_20381);
and U20486 (N_20486,N_20344,N_20234);
and U20487 (N_20487,N_20255,N_20216);
xor U20488 (N_20488,N_20205,N_20248);
or U20489 (N_20489,N_20394,N_20347);
and U20490 (N_20490,N_20306,N_20247);
xnor U20491 (N_20491,N_20204,N_20232);
or U20492 (N_20492,N_20374,N_20249);
nand U20493 (N_20493,N_20256,N_20368);
nor U20494 (N_20494,N_20382,N_20340);
or U20495 (N_20495,N_20334,N_20342);
nor U20496 (N_20496,N_20222,N_20393);
and U20497 (N_20497,N_20291,N_20228);
xor U20498 (N_20498,N_20351,N_20359);
or U20499 (N_20499,N_20251,N_20221);
nor U20500 (N_20500,N_20387,N_20209);
or U20501 (N_20501,N_20269,N_20212);
nand U20502 (N_20502,N_20361,N_20299);
nand U20503 (N_20503,N_20315,N_20341);
and U20504 (N_20504,N_20211,N_20303);
nand U20505 (N_20505,N_20365,N_20273);
nor U20506 (N_20506,N_20297,N_20396);
xor U20507 (N_20507,N_20270,N_20358);
nor U20508 (N_20508,N_20273,N_20378);
or U20509 (N_20509,N_20392,N_20273);
nand U20510 (N_20510,N_20221,N_20266);
or U20511 (N_20511,N_20207,N_20211);
nand U20512 (N_20512,N_20323,N_20305);
nor U20513 (N_20513,N_20272,N_20370);
and U20514 (N_20514,N_20238,N_20282);
nand U20515 (N_20515,N_20351,N_20312);
xor U20516 (N_20516,N_20280,N_20332);
nor U20517 (N_20517,N_20366,N_20393);
or U20518 (N_20518,N_20284,N_20375);
xor U20519 (N_20519,N_20309,N_20213);
nand U20520 (N_20520,N_20267,N_20394);
xnor U20521 (N_20521,N_20216,N_20231);
nor U20522 (N_20522,N_20359,N_20366);
or U20523 (N_20523,N_20282,N_20388);
nand U20524 (N_20524,N_20252,N_20287);
and U20525 (N_20525,N_20268,N_20245);
nand U20526 (N_20526,N_20332,N_20279);
nand U20527 (N_20527,N_20386,N_20255);
nor U20528 (N_20528,N_20209,N_20314);
nor U20529 (N_20529,N_20302,N_20282);
nand U20530 (N_20530,N_20365,N_20392);
xnor U20531 (N_20531,N_20334,N_20228);
and U20532 (N_20532,N_20347,N_20333);
and U20533 (N_20533,N_20398,N_20201);
nand U20534 (N_20534,N_20242,N_20298);
nor U20535 (N_20535,N_20276,N_20227);
or U20536 (N_20536,N_20384,N_20262);
nand U20537 (N_20537,N_20246,N_20235);
nor U20538 (N_20538,N_20246,N_20394);
nor U20539 (N_20539,N_20306,N_20339);
nor U20540 (N_20540,N_20284,N_20296);
nand U20541 (N_20541,N_20320,N_20387);
or U20542 (N_20542,N_20263,N_20271);
or U20543 (N_20543,N_20260,N_20366);
xnor U20544 (N_20544,N_20398,N_20203);
xnor U20545 (N_20545,N_20334,N_20268);
nor U20546 (N_20546,N_20372,N_20363);
or U20547 (N_20547,N_20268,N_20281);
nand U20548 (N_20548,N_20230,N_20235);
nand U20549 (N_20549,N_20221,N_20368);
and U20550 (N_20550,N_20337,N_20347);
xnor U20551 (N_20551,N_20204,N_20243);
and U20552 (N_20552,N_20201,N_20239);
xor U20553 (N_20553,N_20355,N_20272);
xor U20554 (N_20554,N_20346,N_20212);
xor U20555 (N_20555,N_20366,N_20271);
nand U20556 (N_20556,N_20298,N_20388);
xor U20557 (N_20557,N_20248,N_20204);
xnor U20558 (N_20558,N_20372,N_20376);
or U20559 (N_20559,N_20329,N_20324);
or U20560 (N_20560,N_20212,N_20372);
or U20561 (N_20561,N_20354,N_20205);
or U20562 (N_20562,N_20356,N_20367);
and U20563 (N_20563,N_20238,N_20350);
xnor U20564 (N_20564,N_20285,N_20318);
or U20565 (N_20565,N_20377,N_20361);
nor U20566 (N_20566,N_20322,N_20361);
and U20567 (N_20567,N_20254,N_20383);
and U20568 (N_20568,N_20241,N_20393);
and U20569 (N_20569,N_20266,N_20241);
and U20570 (N_20570,N_20292,N_20270);
and U20571 (N_20571,N_20340,N_20356);
or U20572 (N_20572,N_20267,N_20266);
and U20573 (N_20573,N_20273,N_20274);
nor U20574 (N_20574,N_20342,N_20208);
and U20575 (N_20575,N_20244,N_20363);
nor U20576 (N_20576,N_20375,N_20265);
and U20577 (N_20577,N_20342,N_20201);
and U20578 (N_20578,N_20376,N_20364);
nand U20579 (N_20579,N_20355,N_20349);
and U20580 (N_20580,N_20254,N_20208);
nand U20581 (N_20581,N_20237,N_20296);
nor U20582 (N_20582,N_20240,N_20330);
nor U20583 (N_20583,N_20334,N_20251);
or U20584 (N_20584,N_20305,N_20390);
or U20585 (N_20585,N_20342,N_20264);
nor U20586 (N_20586,N_20231,N_20291);
or U20587 (N_20587,N_20330,N_20250);
nor U20588 (N_20588,N_20395,N_20289);
or U20589 (N_20589,N_20277,N_20399);
xnor U20590 (N_20590,N_20297,N_20258);
or U20591 (N_20591,N_20221,N_20300);
xnor U20592 (N_20592,N_20327,N_20302);
or U20593 (N_20593,N_20200,N_20243);
or U20594 (N_20594,N_20327,N_20218);
xnor U20595 (N_20595,N_20222,N_20311);
nor U20596 (N_20596,N_20209,N_20352);
nor U20597 (N_20597,N_20254,N_20319);
nand U20598 (N_20598,N_20366,N_20334);
nor U20599 (N_20599,N_20375,N_20324);
nor U20600 (N_20600,N_20589,N_20433);
nor U20601 (N_20601,N_20499,N_20459);
nor U20602 (N_20602,N_20502,N_20507);
or U20603 (N_20603,N_20508,N_20463);
xnor U20604 (N_20604,N_20552,N_20521);
and U20605 (N_20605,N_20434,N_20597);
nand U20606 (N_20606,N_20549,N_20545);
nor U20607 (N_20607,N_20450,N_20412);
or U20608 (N_20608,N_20586,N_20556);
xnor U20609 (N_20609,N_20415,N_20538);
xor U20610 (N_20610,N_20573,N_20474);
or U20611 (N_20611,N_20500,N_20461);
or U20612 (N_20612,N_20567,N_20587);
nor U20613 (N_20613,N_20446,N_20443);
or U20614 (N_20614,N_20419,N_20458);
xor U20615 (N_20615,N_20490,N_20471);
nand U20616 (N_20616,N_20553,N_20493);
or U20617 (N_20617,N_20515,N_20531);
and U20618 (N_20618,N_20579,N_20451);
or U20619 (N_20619,N_20491,N_20470);
nand U20620 (N_20620,N_20519,N_20505);
nand U20621 (N_20621,N_20486,N_20488);
nand U20622 (N_20622,N_20475,N_20422);
and U20623 (N_20623,N_20598,N_20527);
and U20624 (N_20624,N_20543,N_20539);
nand U20625 (N_20625,N_20467,N_20420);
nand U20626 (N_20626,N_20423,N_20456);
xnor U20627 (N_20627,N_20535,N_20481);
xor U20628 (N_20628,N_20557,N_20516);
xnor U20629 (N_20629,N_20476,N_20438);
xnor U20630 (N_20630,N_20453,N_20501);
nand U20631 (N_20631,N_20593,N_20489);
nor U20632 (N_20632,N_20546,N_20568);
xnor U20633 (N_20633,N_20492,N_20574);
nand U20634 (N_20634,N_20599,N_20506);
or U20635 (N_20635,N_20540,N_20444);
nand U20636 (N_20636,N_20482,N_20437);
or U20637 (N_20637,N_20594,N_20407);
nand U20638 (N_20638,N_20401,N_20426);
nand U20639 (N_20639,N_20427,N_20429);
or U20640 (N_20640,N_20485,N_20517);
nand U20641 (N_20641,N_20581,N_20509);
nand U20642 (N_20642,N_20569,N_20484);
or U20643 (N_20643,N_20590,N_20542);
nor U20644 (N_20644,N_20466,N_20550);
and U20645 (N_20645,N_20409,N_20523);
nand U20646 (N_20646,N_20462,N_20582);
nand U20647 (N_20647,N_20465,N_20411);
nand U20648 (N_20648,N_20580,N_20400);
nand U20649 (N_20649,N_20551,N_20410);
or U20650 (N_20650,N_20406,N_20478);
or U20651 (N_20651,N_20530,N_20532);
or U20652 (N_20652,N_20548,N_20421);
and U20653 (N_20653,N_20588,N_20578);
nor U20654 (N_20654,N_20522,N_20591);
nor U20655 (N_20655,N_20439,N_20554);
nand U20656 (N_20656,N_20479,N_20469);
or U20657 (N_20657,N_20562,N_20457);
nor U20658 (N_20658,N_20503,N_20577);
nand U20659 (N_20659,N_20536,N_20565);
nand U20660 (N_20660,N_20441,N_20436);
xor U20661 (N_20661,N_20583,N_20404);
or U20662 (N_20662,N_20529,N_20408);
and U20663 (N_20663,N_20480,N_20430);
and U20664 (N_20664,N_20566,N_20520);
or U20665 (N_20665,N_20468,N_20526);
nand U20666 (N_20666,N_20555,N_20416);
nand U20667 (N_20667,N_20559,N_20428);
nor U20668 (N_20668,N_20431,N_20448);
xnor U20669 (N_20669,N_20564,N_20524);
nor U20670 (N_20670,N_20454,N_20447);
or U20671 (N_20671,N_20405,N_20442);
and U20672 (N_20672,N_20494,N_20514);
nor U20673 (N_20673,N_20544,N_20413);
or U20674 (N_20674,N_20497,N_20495);
nand U20675 (N_20675,N_20528,N_20473);
xnor U20676 (N_20676,N_20472,N_20402);
or U20677 (N_20677,N_20575,N_20518);
nor U20678 (N_20678,N_20424,N_20432);
nor U20679 (N_20679,N_20585,N_20455);
and U20680 (N_20680,N_20592,N_20418);
and U20681 (N_20681,N_20435,N_20417);
or U20682 (N_20682,N_20561,N_20571);
and U20683 (N_20683,N_20512,N_20533);
nand U20684 (N_20684,N_20477,N_20425);
and U20685 (N_20685,N_20496,N_20525);
or U20686 (N_20686,N_20596,N_20572);
xor U20687 (N_20687,N_20513,N_20563);
xnor U20688 (N_20688,N_20547,N_20534);
nand U20689 (N_20689,N_20541,N_20403);
xor U20690 (N_20690,N_20414,N_20452);
xor U20691 (N_20691,N_20595,N_20449);
and U20692 (N_20692,N_20460,N_20487);
and U20693 (N_20693,N_20510,N_20560);
or U20694 (N_20694,N_20504,N_20570);
or U20695 (N_20695,N_20483,N_20537);
or U20696 (N_20696,N_20558,N_20498);
nand U20697 (N_20697,N_20584,N_20464);
nand U20698 (N_20698,N_20576,N_20440);
or U20699 (N_20699,N_20445,N_20511);
and U20700 (N_20700,N_20562,N_20578);
xnor U20701 (N_20701,N_20461,N_20451);
or U20702 (N_20702,N_20513,N_20573);
nor U20703 (N_20703,N_20533,N_20521);
nand U20704 (N_20704,N_20445,N_20405);
nand U20705 (N_20705,N_20545,N_20488);
xnor U20706 (N_20706,N_20552,N_20433);
nand U20707 (N_20707,N_20592,N_20557);
xor U20708 (N_20708,N_20528,N_20589);
nor U20709 (N_20709,N_20407,N_20538);
nand U20710 (N_20710,N_20558,N_20563);
and U20711 (N_20711,N_20464,N_20503);
xor U20712 (N_20712,N_20443,N_20465);
nor U20713 (N_20713,N_20425,N_20492);
nor U20714 (N_20714,N_20416,N_20564);
and U20715 (N_20715,N_20459,N_20471);
xor U20716 (N_20716,N_20549,N_20481);
nor U20717 (N_20717,N_20406,N_20492);
nand U20718 (N_20718,N_20440,N_20538);
and U20719 (N_20719,N_20571,N_20556);
xnor U20720 (N_20720,N_20477,N_20538);
and U20721 (N_20721,N_20546,N_20515);
nor U20722 (N_20722,N_20504,N_20467);
or U20723 (N_20723,N_20509,N_20529);
or U20724 (N_20724,N_20507,N_20465);
xor U20725 (N_20725,N_20540,N_20528);
nor U20726 (N_20726,N_20500,N_20429);
xnor U20727 (N_20727,N_20584,N_20549);
nand U20728 (N_20728,N_20433,N_20438);
and U20729 (N_20729,N_20514,N_20489);
nand U20730 (N_20730,N_20556,N_20436);
or U20731 (N_20731,N_20522,N_20480);
and U20732 (N_20732,N_20407,N_20508);
nor U20733 (N_20733,N_20559,N_20475);
and U20734 (N_20734,N_20551,N_20574);
and U20735 (N_20735,N_20505,N_20534);
nand U20736 (N_20736,N_20500,N_20565);
nand U20737 (N_20737,N_20566,N_20453);
xor U20738 (N_20738,N_20420,N_20458);
or U20739 (N_20739,N_20508,N_20456);
or U20740 (N_20740,N_20514,N_20460);
or U20741 (N_20741,N_20538,N_20531);
nand U20742 (N_20742,N_20586,N_20544);
and U20743 (N_20743,N_20530,N_20422);
or U20744 (N_20744,N_20457,N_20482);
nor U20745 (N_20745,N_20556,N_20588);
and U20746 (N_20746,N_20456,N_20479);
nand U20747 (N_20747,N_20582,N_20512);
or U20748 (N_20748,N_20597,N_20480);
or U20749 (N_20749,N_20490,N_20580);
or U20750 (N_20750,N_20493,N_20513);
xnor U20751 (N_20751,N_20521,N_20432);
and U20752 (N_20752,N_20403,N_20405);
nand U20753 (N_20753,N_20496,N_20484);
xor U20754 (N_20754,N_20431,N_20553);
and U20755 (N_20755,N_20492,N_20474);
or U20756 (N_20756,N_20447,N_20535);
nand U20757 (N_20757,N_20512,N_20592);
nand U20758 (N_20758,N_20410,N_20587);
nor U20759 (N_20759,N_20587,N_20462);
nor U20760 (N_20760,N_20590,N_20577);
nand U20761 (N_20761,N_20532,N_20512);
xnor U20762 (N_20762,N_20448,N_20476);
and U20763 (N_20763,N_20507,N_20535);
and U20764 (N_20764,N_20531,N_20509);
and U20765 (N_20765,N_20487,N_20592);
and U20766 (N_20766,N_20509,N_20477);
nor U20767 (N_20767,N_20442,N_20457);
nand U20768 (N_20768,N_20554,N_20531);
and U20769 (N_20769,N_20458,N_20543);
xnor U20770 (N_20770,N_20490,N_20564);
xnor U20771 (N_20771,N_20509,N_20546);
xnor U20772 (N_20772,N_20468,N_20546);
or U20773 (N_20773,N_20542,N_20404);
nand U20774 (N_20774,N_20410,N_20585);
and U20775 (N_20775,N_20567,N_20401);
and U20776 (N_20776,N_20505,N_20593);
nor U20777 (N_20777,N_20583,N_20599);
xnor U20778 (N_20778,N_20482,N_20529);
or U20779 (N_20779,N_20432,N_20445);
and U20780 (N_20780,N_20446,N_20448);
xnor U20781 (N_20781,N_20531,N_20542);
nand U20782 (N_20782,N_20485,N_20440);
xor U20783 (N_20783,N_20495,N_20500);
nand U20784 (N_20784,N_20434,N_20419);
nor U20785 (N_20785,N_20507,N_20554);
and U20786 (N_20786,N_20489,N_20522);
or U20787 (N_20787,N_20581,N_20592);
or U20788 (N_20788,N_20451,N_20406);
and U20789 (N_20789,N_20478,N_20413);
and U20790 (N_20790,N_20443,N_20489);
nand U20791 (N_20791,N_20532,N_20511);
or U20792 (N_20792,N_20445,N_20561);
and U20793 (N_20793,N_20444,N_20479);
nand U20794 (N_20794,N_20410,N_20553);
or U20795 (N_20795,N_20567,N_20576);
nor U20796 (N_20796,N_20464,N_20590);
and U20797 (N_20797,N_20526,N_20595);
and U20798 (N_20798,N_20432,N_20429);
xnor U20799 (N_20799,N_20453,N_20429);
nor U20800 (N_20800,N_20623,N_20632);
and U20801 (N_20801,N_20731,N_20780);
xnor U20802 (N_20802,N_20601,N_20696);
and U20803 (N_20803,N_20771,N_20667);
and U20804 (N_20804,N_20676,N_20759);
or U20805 (N_20805,N_20796,N_20652);
nor U20806 (N_20806,N_20778,N_20747);
or U20807 (N_20807,N_20608,N_20713);
xor U20808 (N_20808,N_20664,N_20784);
or U20809 (N_20809,N_20774,N_20790);
and U20810 (N_20810,N_20793,N_20628);
nand U20811 (N_20811,N_20721,N_20706);
xnor U20812 (N_20812,N_20723,N_20733);
and U20813 (N_20813,N_20714,N_20712);
nand U20814 (N_20814,N_20702,N_20647);
nor U20815 (N_20815,N_20604,N_20799);
nor U20816 (N_20816,N_20772,N_20665);
nor U20817 (N_20817,N_20743,N_20677);
nand U20818 (N_20818,N_20616,N_20657);
xnor U20819 (N_20819,N_20697,N_20719);
nand U20820 (N_20820,N_20787,N_20736);
nand U20821 (N_20821,N_20624,N_20678);
nor U20822 (N_20822,N_20634,N_20625);
and U20823 (N_20823,N_20795,N_20755);
or U20824 (N_20824,N_20646,N_20607);
nand U20825 (N_20825,N_20658,N_20749);
nor U20826 (N_20826,N_20727,N_20758);
and U20827 (N_20827,N_20668,N_20732);
and U20828 (N_20828,N_20783,N_20698);
xnor U20829 (N_20829,N_20726,N_20602);
nor U20830 (N_20830,N_20770,N_20687);
and U20831 (N_20831,N_20710,N_20617);
and U20832 (N_20832,N_20656,N_20785);
nor U20833 (N_20833,N_20773,N_20720);
xor U20834 (N_20834,N_20782,N_20729);
or U20835 (N_20835,N_20798,N_20661);
nand U20836 (N_20836,N_20612,N_20666);
and U20837 (N_20837,N_20748,N_20688);
or U20838 (N_20838,N_20606,N_20769);
nand U20839 (N_20839,N_20672,N_20674);
nor U20840 (N_20840,N_20752,N_20767);
and U20841 (N_20841,N_20662,N_20750);
and U20842 (N_20842,N_20707,N_20671);
nor U20843 (N_20843,N_20663,N_20762);
and U20844 (N_20844,N_20627,N_20722);
and U20845 (N_20845,N_20600,N_20768);
nor U20846 (N_20846,N_20635,N_20610);
and U20847 (N_20847,N_20630,N_20746);
nor U20848 (N_20848,N_20645,N_20739);
and U20849 (N_20849,N_20682,N_20766);
or U20850 (N_20850,N_20649,N_20614);
and U20851 (N_20851,N_20695,N_20611);
xnor U20852 (N_20852,N_20692,N_20648);
nand U20853 (N_20853,N_20705,N_20659);
nand U20854 (N_20854,N_20641,N_20615);
or U20855 (N_20855,N_20741,N_20763);
or U20856 (N_20856,N_20684,N_20788);
and U20857 (N_20857,N_20637,N_20699);
nor U20858 (N_20858,N_20613,N_20753);
nand U20859 (N_20859,N_20751,N_20670);
nor U20860 (N_20860,N_20740,N_20711);
nor U20861 (N_20861,N_20689,N_20734);
nand U20862 (N_20862,N_20760,N_20685);
xnor U20863 (N_20863,N_20715,N_20756);
and U20864 (N_20864,N_20728,N_20777);
xnor U20865 (N_20865,N_20683,N_20764);
and U20866 (N_20866,N_20738,N_20701);
nand U20867 (N_20867,N_20603,N_20620);
nor U20868 (N_20868,N_20754,N_20791);
and U20869 (N_20869,N_20631,N_20626);
xor U20870 (N_20870,N_20690,N_20651);
nand U20871 (N_20871,N_20724,N_20673);
nand U20872 (N_20872,N_20633,N_20638);
or U20873 (N_20873,N_20716,N_20618);
or U20874 (N_20874,N_20704,N_20789);
or U20875 (N_20875,N_20644,N_20745);
nor U20876 (N_20876,N_20686,N_20757);
xnor U20877 (N_20877,N_20642,N_20742);
xnor U20878 (N_20878,N_20775,N_20639);
xnor U20879 (N_20879,N_20680,N_20737);
or U20880 (N_20880,N_20669,N_20797);
xnor U20881 (N_20881,N_20640,N_20694);
nand U20882 (N_20882,N_20643,N_20655);
or U20883 (N_20883,N_20700,N_20725);
or U20884 (N_20884,N_20650,N_20781);
or U20885 (N_20885,N_20636,N_20693);
xor U20886 (N_20886,N_20605,N_20765);
xnor U20887 (N_20887,N_20621,N_20792);
nand U20888 (N_20888,N_20709,N_20629);
xor U20889 (N_20889,N_20718,N_20703);
nand U20890 (N_20890,N_20691,N_20660);
nor U20891 (N_20891,N_20779,N_20654);
and U20892 (N_20892,N_20619,N_20776);
nor U20893 (N_20893,N_20794,N_20679);
nand U20894 (N_20894,N_20675,N_20735);
and U20895 (N_20895,N_20717,N_20681);
or U20896 (N_20896,N_20786,N_20761);
or U20897 (N_20897,N_20744,N_20609);
or U20898 (N_20898,N_20653,N_20708);
nand U20899 (N_20899,N_20730,N_20622);
xnor U20900 (N_20900,N_20760,N_20747);
nand U20901 (N_20901,N_20657,N_20729);
and U20902 (N_20902,N_20674,N_20769);
and U20903 (N_20903,N_20622,N_20637);
xnor U20904 (N_20904,N_20600,N_20674);
or U20905 (N_20905,N_20673,N_20652);
nor U20906 (N_20906,N_20792,N_20764);
nand U20907 (N_20907,N_20655,N_20647);
and U20908 (N_20908,N_20634,N_20749);
nand U20909 (N_20909,N_20645,N_20763);
and U20910 (N_20910,N_20796,N_20752);
and U20911 (N_20911,N_20641,N_20776);
nor U20912 (N_20912,N_20723,N_20748);
xor U20913 (N_20913,N_20719,N_20774);
or U20914 (N_20914,N_20780,N_20645);
and U20915 (N_20915,N_20604,N_20704);
and U20916 (N_20916,N_20763,N_20796);
nand U20917 (N_20917,N_20651,N_20640);
xor U20918 (N_20918,N_20725,N_20778);
nor U20919 (N_20919,N_20670,N_20674);
nand U20920 (N_20920,N_20707,N_20714);
xor U20921 (N_20921,N_20737,N_20624);
nand U20922 (N_20922,N_20677,N_20660);
or U20923 (N_20923,N_20631,N_20617);
xnor U20924 (N_20924,N_20686,N_20668);
and U20925 (N_20925,N_20762,N_20793);
xor U20926 (N_20926,N_20723,N_20790);
nor U20927 (N_20927,N_20761,N_20701);
xor U20928 (N_20928,N_20660,N_20784);
nand U20929 (N_20929,N_20668,N_20710);
nand U20930 (N_20930,N_20626,N_20718);
xor U20931 (N_20931,N_20647,N_20799);
nand U20932 (N_20932,N_20624,N_20736);
nand U20933 (N_20933,N_20711,N_20667);
and U20934 (N_20934,N_20773,N_20705);
xor U20935 (N_20935,N_20694,N_20758);
or U20936 (N_20936,N_20758,N_20790);
nor U20937 (N_20937,N_20696,N_20710);
nor U20938 (N_20938,N_20741,N_20786);
and U20939 (N_20939,N_20777,N_20668);
nor U20940 (N_20940,N_20795,N_20754);
and U20941 (N_20941,N_20716,N_20677);
or U20942 (N_20942,N_20634,N_20637);
xnor U20943 (N_20943,N_20612,N_20722);
xnor U20944 (N_20944,N_20616,N_20710);
or U20945 (N_20945,N_20777,N_20674);
or U20946 (N_20946,N_20786,N_20758);
nand U20947 (N_20947,N_20784,N_20755);
or U20948 (N_20948,N_20616,N_20652);
or U20949 (N_20949,N_20783,N_20695);
nand U20950 (N_20950,N_20650,N_20672);
xnor U20951 (N_20951,N_20650,N_20627);
xnor U20952 (N_20952,N_20765,N_20778);
xor U20953 (N_20953,N_20749,N_20766);
nor U20954 (N_20954,N_20706,N_20796);
nand U20955 (N_20955,N_20727,N_20780);
nand U20956 (N_20956,N_20742,N_20681);
and U20957 (N_20957,N_20611,N_20683);
nor U20958 (N_20958,N_20649,N_20618);
and U20959 (N_20959,N_20630,N_20658);
or U20960 (N_20960,N_20727,N_20684);
and U20961 (N_20961,N_20792,N_20691);
nand U20962 (N_20962,N_20770,N_20783);
nor U20963 (N_20963,N_20772,N_20680);
and U20964 (N_20964,N_20673,N_20756);
nand U20965 (N_20965,N_20726,N_20757);
and U20966 (N_20966,N_20660,N_20751);
xnor U20967 (N_20967,N_20683,N_20728);
xnor U20968 (N_20968,N_20673,N_20763);
or U20969 (N_20969,N_20770,N_20757);
xnor U20970 (N_20970,N_20618,N_20757);
and U20971 (N_20971,N_20788,N_20787);
nor U20972 (N_20972,N_20669,N_20788);
nor U20973 (N_20973,N_20791,N_20667);
nand U20974 (N_20974,N_20604,N_20764);
or U20975 (N_20975,N_20646,N_20684);
and U20976 (N_20976,N_20714,N_20786);
or U20977 (N_20977,N_20619,N_20626);
nand U20978 (N_20978,N_20640,N_20725);
nand U20979 (N_20979,N_20788,N_20797);
and U20980 (N_20980,N_20722,N_20761);
or U20981 (N_20981,N_20618,N_20710);
xnor U20982 (N_20982,N_20761,N_20715);
nor U20983 (N_20983,N_20776,N_20740);
and U20984 (N_20984,N_20778,N_20709);
and U20985 (N_20985,N_20640,N_20619);
and U20986 (N_20986,N_20690,N_20720);
and U20987 (N_20987,N_20720,N_20711);
nand U20988 (N_20988,N_20733,N_20629);
nor U20989 (N_20989,N_20749,N_20675);
xnor U20990 (N_20990,N_20626,N_20668);
nor U20991 (N_20991,N_20733,N_20627);
xor U20992 (N_20992,N_20757,N_20749);
and U20993 (N_20993,N_20783,N_20704);
and U20994 (N_20994,N_20731,N_20744);
and U20995 (N_20995,N_20737,N_20673);
and U20996 (N_20996,N_20627,N_20775);
or U20997 (N_20997,N_20779,N_20767);
nand U20998 (N_20998,N_20697,N_20755);
nand U20999 (N_20999,N_20670,N_20617);
or U21000 (N_21000,N_20862,N_20956);
nand U21001 (N_21001,N_20835,N_20897);
xor U21002 (N_21002,N_20802,N_20925);
nor U21003 (N_21003,N_20983,N_20931);
nand U21004 (N_21004,N_20974,N_20946);
nor U21005 (N_21005,N_20883,N_20866);
nor U21006 (N_21006,N_20998,N_20807);
xor U21007 (N_21007,N_20858,N_20818);
nor U21008 (N_21008,N_20895,N_20877);
xnor U21009 (N_21009,N_20841,N_20923);
nor U21010 (N_21010,N_20806,N_20943);
xnor U21011 (N_21011,N_20881,N_20864);
and U21012 (N_21012,N_20810,N_20838);
nor U21013 (N_21013,N_20947,N_20855);
and U21014 (N_21014,N_20813,N_20850);
nor U21015 (N_21015,N_20856,N_20913);
nand U21016 (N_21016,N_20859,N_20996);
nor U21017 (N_21017,N_20955,N_20990);
nand U21018 (N_21018,N_20819,N_20971);
xnor U21019 (N_21019,N_20900,N_20961);
and U21020 (N_21020,N_20888,N_20811);
xnor U21021 (N_21021,N_20800,N_20889);
or U21022 (N_21022,N_20975,N_20911);
xor U21023 (N_21023,N_20977,N_20814);
xnor U21024 (N_21024,N_20853,N_20816);
or U21025 (N_21025,N_20884,N_20849);
and U21026 (N_21026,N_20916,N_20939);
nor U21027 (N_21027,N_20832,N_20936);
or U21028 (N_21028,N_20976,N_20903);
nor U21029 (N_21029,N_20969,N_20929);
or U21030 (N_21030,N_20804,N_20890);
xor U21031 (N_21031,N_20979,N_20970);
xor U21032 (N_21032,N_20840,N_20886);
xnor U21033 (N_21033,N_20966,N_20869);
nor U21034 (N_21034,N_20885,N_20892);
or U21035 (N_21035,N_20826,N_20863);
or U21036 (N_21036,N_20952,N_20847);
xor U21037 (N_21037,N_20910,N_20896);
and U21038 (N_21038,N_20972,N_20879);
or U21039 (N_21039,N_20941,N_20868);
or U21040 (N_21040,N_20940,N_20872);
or U21041 (N_21041,N_20882,N_20934);
and U21042 (N_21042,N_20991,N_20928);
xor U21043 (N_21043,N_20948,N_20857);
or U21044 (N_21044,N_20957,N_20978);
and U21045 (N_21045,N_20875,N_20824);
nor U21046 (N_21046,N_20980,N_20950);
xor U21047 (N_21047,N_20917,N_20815);
xnor U21048 (N_21048,N_20878,N_20909);
nand U21049 (N_21049,N_20839,N_20962);
nor U21050 (N_21050,N_20921,N_20907);
xor U21051 (N_21051,N_20965,N_20844);
xnor U21052 (N_21052,N_20876,N_20904);
or U21053 (N_21053,N_20959,N_20820);
and U21054 (N_21054,N_20932,N_20993);
or U21055 (N_21055,N_20836,N_20845);
xnor U21056 (N_21056,N_20831,N_20842);
nand U21057 (N_21057,N_20809,N_20898);
and U21058 (N_21058,N_20828,N_20801);
nor U21059 (N_21059,N_20914,N_20987);
nor U21060 (N_21060,N_20860,N_20817);
and U21061 (N_21061,N_20964,N_20905);
nor U21062 (N_21062,N_20981,N_20803);
nand U21063 (N_21063,N_20949,N_20927);
nand U21064 (N_21064,N_20837,N_20852);
nand U21065 (N_21065,N_20861,N_20899);
or U21066 (N_21066,N_20937,N_20989);
and U21067 (N_21067,N_20843,N_20999);
nand U21068 (N_21068,N_20958,N_20973);
nand U21069 (N_21069,N_20871,N_20846);
nor U21070 (N_21070,N_20865,N_20933);
nor U21071 (N_21071,N_20854,N_20912);
and U21072 (N_21072,N_20902,N_20920);
or U21073 (N_21073,N_20825,N_20919);
or U21074 (N_21074,N_20924,N_20848);
nor U21075 (N_21075,N_20985,N_20867);
nor U21076 (N_21076,N_20822,N_20880);
and U21077 (N_21077,N_20874,N_20894);
xnor U21078 (N_21078,N_20805,N_20930);
and U21079 (N_21079,N_20935,N_20906);
nand U21080 (N_21080,N_20938,N_20942);
nor U21081 (N_21081,N_20984,N_20908);
nand U21082 (N_21082,N_20968,N_20873);
and U21083 (N_21083,N_20945,N_20823);
nor U21084 (N_21084,N_20997,N_20833);
and U21085 (N_21085,N_20986,N_20960);
nor U21086 (N_21086,N_20870,N_20992);
or U21087 (N_21087,N_20915,N_20851);
xnor U21088 (N_21088,N_20982,N_20988);
and U21089 (N_21089,N_20967,N_20954);
xnor U21090 (N_21090,N_20821,N_20829);
or U21091 (N_21091,N_20951,N_20953);
or U21092 (N_21092,N_20922,N_20995);
nand U21093 (N_21093,N_20893,N_20944);
or U21094 (N_21094,N_20834,N_20808);
nand U21095 (N_21095,N_20827,N_20830);
xor U21096 (N_21096,N_20812,N_20918);
or U21097 (N_21097,N_20887,N_20994);
xnor U21098 (N_21098,N_20901,N_20891);
nor U21099 (N_21099,N_20926,N_20963);
xor U21100 (N_21100,N_20849,N_20844);
or U21101 (N_21101,N_20971,N_20975);
or U21102 (N_21102,N_20805,N_20925);
and U21103 (N_21103,N_20871,N_20893);
nor U21104 (N_21104,N_20961,N_20933);
or U21105 (N_21105,N_20881,N_20909);
xnor U21106 (N_21106,N_20941,N_20999);
xor U21107 (N_21107,N_20815,N_20874);
nand U21108 (N_21108,N_20962,N_20849);
nand U21109 (N_21109,N_20850,N_20817);
or U21110 (N_21110,N_20805,N_20801);
nand U21111 (N_21111,N_20811,N_20825);
and U21112 (N_21112,N_20913,N_20822);
nand U21113 (N_21113,N_20855,N_20832);
or U21114 (N_21114,N_20925,N_20938);
nand U21115 (N_21115,N_20900,N_20992);
and U21116 (N_21116,N_20938,N_20977);
xnor U21117 (N_21117,N_20936,N_20820);
or U21118 (N_21118,N_20845,N_20869);
nand U21119 (N_21119,N_20864,N_20876);
nor U21120 (N_21120,N_20973,N_20886);
and U21121 (N_21121,N_20988,N_20927);
nand U21122 (N_21122,N_20816,N_20993);
and U21123 (N_21123,N_20889,N_20999);
and U21124 (N_21124,N_20869,N_20929);
nand U21125 (N_21125,N_20829,N_20845);
or U21126 (N_21126,N_20844,N_20880);
xor U21127 (N_21127,N_20849,N_20932);
and U21128 (N_21128,N_20913,N_20834);
nor U21129 (N_21129,N_20803,N_20824);
and U21130 (N_21130,N_20958,N_20826);
and U21131 (N_21131,N_20932,N_20934);
nor U21132 (N_21132,N_20856,N_20833);
xnor U21133 (N_21133,N_20912,N_20940);
xnor U21134 (N_21134,N_20849,N_20800);
and U21135 (N_21135,N_20891,N_20807);
xor U21136 (N_21136,N_20854,N_20933);
xnor U21137 (N_21137,N_20893,N_20829);
xor U21138 (N_21138,N_20858,N_20967);
xnor U21139 (N_21139,N_20955,N_20928);
xnor U21140 (N_21140,N_20996,N_20879);
nand U21141 (N_21141,N_20837,N_20820);
or U21142 (N_21142,N_20820,N_20822);
nand U21143 (N_21143,N_20840,N_20990);
xnor U21144 (N_21144,N_20854,N_20825);
nand U21145 (N_21145,N_20891,N_20940);
and U21146 (N_21146,N_20989,N_20980);
xor U21147 (N_21147,N_20889,N_20803);
xor U21148 (N_21148,N_20899,N_20916);
or U21149 (N_21149,N_20843,N_20917);
nor U21150 (N_21150,N_20979,N_20905);
nor U21151 (N_21151,N_20971,N_20969);
xor U21152 (N_21152,N_20986,N_20899);
xor U21153 (N_21153,N_20991,N_20886);
nand U21154 (N_21154,N_20963,N_20911);
xor U21155 (N_21155,N_20991,N_20819);
nand U21156 (N_21156,N_20951,N_20998);
nand U21157 (N_21157,N_20898,N_20855);
nor U21158 (N_21158,N_20961,N_20994);
nor U21159 (N_21159,N_20803,N_20983);
nor U21160 (N_21160,N_20806,N_20890);
nand U21161 (N_21161,N_20898,N_20955);
nor U21162 (N_21162,N_20858,N_20874);
nor U21163 (N_21163,N_20986,N_20885);
xnor U21164 (N_21164,N_20837,N_20915);
or U21165 (N_21165,N_20875,N_20803);
xnor U21166 (N_21166,N_20836,N_20875);
xnor U21167 (N_21167,N_20848,N_20905);
nand U21168 (N_21168,N_20906,N_20821);
xnor U21169 (N_21169,N_20935,N_20850);
nand U21170 (N_21170,N_20853,N_20960);
xnor U21171 (N_21171,N_20862,N_20822);
xor U21172 (N_21172,N_20903,N_20812);
or U21173 (N_21173,N_20882,N_20840);
nand U21174 (N_21174,N_20938,N_20984);
xor U21175 (N_21175,N_20855,N_20890);
and U21176 (N_21176,N_20969,N_20803);
xnor U21177 (N_21177,N_20891,N_20979);
nor U21178 (N_21178,N_20849,N_20930);
or U21179 (N_21179,N_20842,N_20880);
nor U21180 (N_21180,N_20955,N_20859);
or U21181 (N_21181,N_20977,N_20833);
nor U21182 (N_21182,N_20824,N_20947);
and U21183 (N_21183,N_20802,N_20974);
xnor U21184 (N_21184,N_20804,N_20918);
nand U21185 (N_21185,N_20836,N_20955);
xor U21186 (N_21186,N_20927,N_20966);
nor U21187 (N_21187,N_20928,N_20919);
or U21188 (N_21188,N_20979,N_20981);
nor U21189 (N_21189,N_20807,N_20811);
xor U21190 (N_21190,N_20966,N_20826);
nor U21191 (N_21191,N_20897,N_20869);
xor U21192 (N_21192,N_20878,N_20822);
nand U21193 (N_21193,N_20874,N_20990);
nor U21194 (N_21194,N_20896,N_20826);
xnor U21195 (N_21195,N_20926,N_20820);
or U21196 (N_21196,N_20922,N_20974);
or U21197 (N_21197,N_20999,N_20837);
nand U21198 (N_21198,N_20837,N_20949);
nor U21199 (N_21199,N_20880,N_20833);
or U21200 (N_21200,N_21090,N_21014);
nor U21201 (N_21201,N_21170,N_21094);
nand U21202 (N_21202,N_21144,N_21158);
and U21203 (N_21203,N_21065,N_21056);
xor U21204 (N_21204,N_21103,N_21044);
or U21205 (N_21205,N_21022,N_21082);
and U21206 (N_21206,N_21162,N_21174);
and U21207 (N_21207,N_21123,N_21182);
nand U21208 (N_21208,N_21122,N_21084);
and U21209 (N_21209,N_21010,N_21039);
or U21210 (N_21210,N_21095,N_21161);
or U21211 (N_21211,N_21115,N_21047);
nor U21212 (N_21212,N_21129,N_21043);
and U21213 (N_21213,N_21165,N_21079);
nand U21214 (N_21214,N_21197,N_21004);
or U21215 (N_21215,N_21118,N_21192);
and U21216 (N_21216,N_21042,N_21074);
nor U21217 (N_21217,N_21052,N_21134);
xor U21218 (N_21218,N_21113,N_21181);
nor U21219 (N_21219,N_21175,N_21183);
nand U21220 (N_21220,N_21085,N_21001);
or U21221 (N_21221,N_21119,N_21045);
nand U21222 (N_21222,N_21066,N_21109);
or U21223 (N_21223,N_21126,N_21127);
nand U21224 (N_21224,N_21027,N_21147);
xor U21225 (N_21225,N_21121,N_21153);
nand U21226 (N_21226,N_21169,N_21193);
or U21227 (N_21227,N_21072,N_21196);
xnor U21228 (N_21228,N_21083,N_21033);
and U21229 (N_21229,N_21116,N_21024);
and U21230 (N_21230,N_21178,N_21008);
xor U21231 (N_21231,N_21187,N_21054);
nor U21232 (N_21232,N_21075,N_21015);
and U21233 (N_21233,N_21003,N_21117);
nand U21234 (N_21234,N_21070,N_21110);
xor U21235 (N_21235,N_21111,N_21006);
nand U21236 (N_21236,N_21159,N_21191);
or U21237 (N_21237,N_21061,N_21104);
nor U21238 (N_21238,N_21125,N_21068);
xor U21239 (N_21239,N_21057,N_21138);
and U21240 (N_21240,N_21180,N_21098);
or U21241 (N_21241,N_21102,N_21114);
nor U21242 (N_21242,N_21150,N_21011);
or U21243 (N_21243,N_21137,N_21131);
xnor U21244 (N_21244,N_21189,N_21031);
and U21245 (N_21245,N_21160,N_21023);
xnor U21246 (N_21246,N_21176,N_21053);
nor U21247 (N_21247,N_21021,N_21164);
nand U21248 (N_21248,N_21186,N_21096);
or U21249 (N_21249,N_21002,N_21173);
or U21250 (N_21250,N_21076,N_21124);
xor U21251 (N_21251,N_21194,N_21152);
or U21252 (N_21252,N_21157,N_21067);
nand U21253 (N_21253,N_21025,N_21133);
nand U21254 (N_21254,N_21064,N_21167);
or U21255 (N_21255,N_21060,N_21005);
or U21256 (N_21256,N_21046,N_21041);
xor U21257 (N_21257,N_21107,N_21097);
nand U21258 (N_21258,N_21035,N_21059);
and U21259 (N_21259,N_21156,N_21130);
or U21260 (N_21260,N_21088,N_21093);
nand U21261 (N_21261,N_21199,N_21168);
nand U21262 (N_21262,N_21012,N_21058);
nand U21263 (N_21263,N_21149,N_21143);
nand U21264 (N_21264,N_21040,N_21092);
xnor U21265 (N_21265,N_21049,N_21034);
xor U21266 (N_21266,N_21029,N_21185);
or U21267 (N_21267,N_21018,N_21177);
or U21268 (N_21268,N_21087,N_21184);
xor U21269 (N_21269,N_21032,N_21081);
xor U21270 (N_21270,N_21062,N_21148);
and U21271 (N_21271,N_21100,N_21020);
nor U21272 (N_21272,N_21142,N_21089);
nor U21273 (N_21273,N_21195,N_21080);
nor U21274 (N_21274,N_21141,N_21112);
nor U21275 (N_21275,N_21108,N_21140);
or U21276 (N_21276,N_21077,N_21050);
and U21277 (N_21277,N_21139,N_21128);
and U21278 (N_21278,N_21030,N_21071);
and U21279 (N_21279,N_21188,N_21055);
xor U21280 (N_21280,N_21163,N_21000);
and U21281 (N_21281,N_21078,N_21135);
nand U21282 (N_21282,N_21154,N_21091);
nor U21283 (N_21283,N_21166,N_21105);
and U21284 (N_21284,N_21013,N_21038);
or U21285 (N_21285,N_21019,N_21017);
nand U21286 (N_21286,N_21120,N_21099);
xor U21287 (N_21287,N_21145,N_21101);
nand U21288 (N_21288,N_21155,N_21136);
nor U21289 (N_21289,N_21037,N_21172);
nand U21290 (N_21290,N_21179,N_21069);
xnor U21291 (N_21291,N_21063,N_21048);
nand U21292 (N_21292,N_21190,N_21009);
xnor U21293 (N_21293,N_21016,N_21036);
xor U21294 (N_21294,N_21028,N_21151);
nor U21295 (N_21295,N_21073,N_21051);
and U21296 (N_21296,N_21026,N_21007);
nor U21297 (N_21297,N_21171,N_21106);
and U21298 (N_21298,N_21086,N_21132);
and U21299 (N_21299,N_21146,N_21198);
xor U21300 (N_21300,N_21071,N_21093);
nand U21301 (N_21301,N_21067,N_21074);
or U21302 (N_21302,N_21032,N_21004);
nor U21303 (N_21303,N_21164,N_21054);
and U21304 (N_21304,N_21102,N_21176);
and U21305 (N_21305,N_21001,N_21011);
or U21306 (N_21306,N_21030,N_21053);
and U21307 (N_21307,N_21104,N_21025);
nand U21308 (N_21308,N_21188,N_21171);
nor U21309 (N_21309,N_21193,N_21052);
and U21310 (N_21310,N_21003,N_21080);
nor U21311 (N_21311,N_21070,N_21164);
nor U21312 (N_21312,N_21175,N_21167);
nand U21313 (N_21313,N_21172,N_21001);
nor U21314 (N_21314,N_21078,N_21067);
nand U21315 (N_21315,N_21152,N_21010);
xnor U21316 (N_21316,N_21175,N_21078);
or U21317 (N_21317,N_21106,N_21077);
nand U21318 (N_21318,N_21124,N_21035);
xor U21319 (N_21319,N_21160,N_21150);
nor U21320 (N_21320,N_21015,N_21001);
or U21321 (N_21321,N_21029,N_21114);
nor U21322 (N_21322,N_21072,N_21181);
or U21323 (N_21323,N_21029,N_21061);
or U21324 (N_21324,N_21064,N_21111);
nor U21325 (N_21325,N_21192,N_21119);
nand U21326 (N_21326,N_21154,N_21193);
or U21327 (N_21327,N_21093,N_21045);
and U21328 (N_21328,N_21184,N_21003);
or U21329 (N_21329,N_21123,N_21071);
nor U21330 (N_21330,N_21191,N_21036);
xnor U21331 (N_21331,N_21043,N_21041);
xor U21332 (N_21332,N_21109,N_21060);
or U21333 (N_21333,N_21153,N_21093);
nor U21334 (N_21334,N_21051,N_21085);
or U21335 (N_21335,N_21150,N_21124);
nor U21336 (N_21336,N_21100,N_21155);
nor U21337 (N_21337,N_21109,N_21102);
nor U21338 (N_21338,N_21094,N_21151);
and U21339 (N_21339,N_21074,N_21072);
xnor U21340 (N_21340,N_21046,N_21091);
nor U21341 (N_21341,N_21072,N_21012);
nand U21342 (N_21342,N_21155,N_21035);
xnor U21343 (N_21343,N_21177,N_21089);
or U21344 (N_21344,N_21001,N_21108);
nand U21345 (N_21345,N_21188,N_21027);
nor U21346 (N_21346,N_21027,N_21167);
and U21347 (N_21347,N_21112,N_21108);
xnor U21348 (N_21348,N_21118,N_21198);
or U21349 (N_21349,N_21068,N_21095);
xor U21350 (N_21350,N_21088,N_21083);
nor U21351 (N_21351,N_21098,N_21020);
xor U21352 (N_21352,N_21198,N_21045);
xnor U21353 (N_21353,N_21180,N_21025);
xnor U21354 (N_21354,N_21136,N_21105);
and U21355 (N_21355,N_21133,N_21026);
and U21356 (N_21356,N_21091,N_21165);
nand U21357 (N_21357,N_21183,N_21014);
nor U21358 (N_21358,N_21008,N_21132);
or U21359 (N_21359,N_21105,N_21066);
and U21360 (N_21360,N_21156,N_21161);
xor U21361 (N_21361,N_21034,N_21150);
and U21362 (N_21362,N_21019,N_21037);
xor U21363 (N_21363,N_21172,N_21005);
nor U21364 (N_21364,N_21109,N_21075);
and U21365 (N_21365,N_21027,N_21134);
nand U21366 (N_21366,N_21086,N_21181);
xnor U21367 (N_21367,N_21030,N_21000);
nand U21368 (N_21368,N_21143,N_21158);
nor U21369 (N_21369,N_21065,N_21018);
nor U21370 (N_21370,N_21046,N_21116);
and U21371 (N_21371,N_21025,N_21046);
nor U21372 (N_21372,N_21007,N_21117);
nor U21373 (N_21373,N_21043,N_21001);
and U21374 (N_21374,N_21116,N_21066);
and U21375 (N_21375,N_21146,N_21164);
xnor U21376 (N_21376,N_21064,N_21140);
and U21377 (N_21377,N_21024,N_21135);
and U21378 (N_21378,N_21193,N_21018);
or U21379 (N_21379,N_21041,N_21010);
xnor U21380 (N_21380,N_21061,N_21003);
and U21381 (N_21381,N_21137,N_21164);
xor U21382 (N_21382,N_21081,N_21087);
or U21383 (N_21383,N_21180,N_21164);
nor U21384 (N_21384,N_21165,N_21124);
nor U21385 (N_21385,N_21021,N_21160);
xor U21386 (N_21386,N_21150,N_21174);
xor U21387 (N_21387,N_21067,N_21119);
nand U21388 (N_21388,N_21138,N_21131);
nor U21389 (N_21389,N_21153,N_21036);
and U21390 (N_21390,N_21186,N_21071);
xnor U21391 (N_21391,N_21080,N_21097);
or U21392 (N_21392,N_21128,N_21108);
xnor U21393 (N_21393,N_21156,N_21154);
xnor U21394 (N_21394,N_21070,N_21169);
nor U21395 (N_21395,N_21199,N_21151);
or U21396 (N_21396,N_21108,N_21157);
and U21397 (N_21397,N_21130,N_21006);
or U21398 (N_21398,N_21164,N_21065);
and U21399 (N_21399,N_21092,N_21146);
nand U21400 (N_21400,N_21213,N_21390);
xnor U21401 (N_21401,N_21313,N_21300);
nor U21402 (N_21402,N_21255,N_21377);
nand U21403 (N_21403,N_21305,N_21200);
and U21404 (N_21404,N_21309,N_21207);
nor U21405 (N_21405,N_21279,N_21219);
nor U21406 (N_21406,N_21239,N_21346);
nand U21407 (N_21407,N_21392,N_21383);
nand U21408 (N_21408,N_21316,N_21218);
and U21409 (N_21409,N_21368,N_21324);
nor U21410 (N_21410,N_21250,N_21273);
nor U21411 (N_21411,N_21275,N_21290);
and U21412 (N_21412,N_21292,N_21358);
nor U21413 (N_21413,N_21240,N_21366);
nor U21414 (N_21414,N_21281,N_21204);
nand U21415 (N_21415,N_21257,N_21256);
nand U21416 (N_21416,N_21352,N_21301);
nand U21417 (N_21417,N_21360,N_21399);
and U21418 (N_21418,N_21342,N_21388);
xnor U21419 (N_21419,N_21303,N_21282);
or U21420 (N_21420,N_21337,N_21336);
nor U21421 (N_21421,N_21386,N_21341);
xor U21422 (N_21422,N_21372,N_21272);
and U21423 (N_21423,N_21306,N_21381);
nor U21424 (N_21424,N_21398,N_21259);
or U21425 (N_21425,N_21252,N_21329);
nor U21426 (N_21426,N_21326,N_21216);
and U21427 (N_21427,N_21293,N_21232);
or U21428 (N_21428,N_21349,N_21243);
nor U21429 (N_21429,N_21288,N_21371);
xnor U21430 (N_21430,N_21268,N_21314);
and U21431 (N_21431,N_21362,N_21354);
nor U21432 (N_21432,N_21345,N_21344);
or U21433 (N_21433,N_21319,N_21353);
or U21434 (N_21434,N_21247,N_21340);
nand U21435 (N_21435,N_21327,N_21389);
xnor U21436 (N_21436,N_21221,N_21287);
nor U21437 (N_21437,N_21269,N_21376);
nand U21438 (N_21438,N_21276,N_21330);
xnor U21439 (N_21439,N_21311,N_21203);
nand U21440 (N_21440,N_21251,N_21334);
and U21441 (N_21441,N_21222,N_21244);
and U21442 (N_21442,N_21363,N_21270);
nor U21443 (N_21443,N_21226,N_21210);
nand U21444 (N_21444,N_21361,N_21231);
nand U21445 (N_21445,N_21223,N_21387);
or U21446 (N_21446,N_21289,N_21318);
nand U21447 (N_21447,N_21205,N_21249);
and U21448 (N_21448,N_21237,N_21350);
nor U21449 (N_21449,N_21320,N_21295);
xor U21450 (N_21450,N_21339,N_21261);
or U21451 (N_21451,N_21296,N_21315);
xnor U21452 (N_21452,N_21291,N_21234);
xor U21453 (N_21453,N_21307,N_21338);
xnor U21454 (N_21454,N_21263,N_21278);
xnor U21455 (N_21455,N_21245,N_21393);
nor U21456 (N_21456,N_21343,N_21317);
nor U21457 (N_21457,N_21285,N_21328);
or U21458 (N_21458,N_21214,N_21298);
nor U21459 (N_21459,N_21308,N_21379);
xnor U21460 (N_21460,N_21322,N_21374);
nand U21461 (N_21461,N_21373,N_21202);
nand U21462 (N_21462,N_21331,N_21236);
and U21463 (N_21463,N_21370,N_21229);
or U21464 (N_21464,N_21384,N_21233);
and U21465 (N_21465,N_21323,N_21378);
or U21466 (N_21466,N_21271,N_21211);
nor U21467 (N_21467,N_21242,N_21356);
and U21468 (N_21468,N_21206,N_21321);
nand U21469 (N_21469,N_21286,N_21304);
and U21470 (N_21470,N_21230,N_21359);
nand U21471 (N_21471,N_21325,N_21227);
xor U21472 (N_21472,N_21208,N_21333);
and U21473 (N_21473,N_21209,N_21264);
or U21474 (N_21474,N_21260,N_21375);
or U21475 (N_21475,N_21225,N_21395);
or U21476 (N_21476,N_21253,N_21365);
nand U21477 (N_21477,N_21246,N_21201);
xor U21478 (N_21478,N_21382,N_21332);
nor U21479 (N_21479,N_21235,N_21258);
or U21480 (N_21480,N_21280,N_21283);
xnor U21481 (N_21481,N_21294,N_21396);
nand U21482 (N_21482,N_21335,N_21364);
and U21483 (N_21483,N_21262,N_21394);
nor U21484 (N_21484,N_21265,N_21380);
nor U21485 (N_21485,N_21357,N_21224);
and U21486 (N_21486,N_21220,N_21312);
or U21487 (N_21487,N_21248,N_21391);
nand U21488 (N_21488,N_21369,N_21277);
xnor U21489 (N_21489,N_21355,N_21348);
xor U21490 (N_21490,N_21297,N_21347);
xor U21491 (N_21491,N_21310,N_21274);
nor U21492 (N_21492,N_21228,N_21284);
and U21493 (N_21493,N_21302,N_21267);
xnor U21494 (N_21494,N_21397,N_21367);
nor U21495 (N_21495,N_21385,N_21238);
and U21496 (N_21496,N_21215,N_21241);
and U21497 (N_21497,N_21299,N_21351);
or U21498 (N_21498,N_21212,N_21254);
xor U21499 (N_21499,N_21217,N_21266);
nor U21500 (N_21500,N_21311,N_21375);
and U21501 (N_21501,N_21259,N_21269);
and U21502 (N_21502,N_21399,N_21315);
and U21503 (N_21503,N_21221,N_21262);
nor U21504 (N_21504,N_21252,N_21381);
xnor U21505 (N_21505,N_21326,N_21213);
nor U21506 (N_21506,N_21378,N_21296);
or U21507 (N_21507,N_21368,N_21278);
nor U21508 (N_21508,N_21266,N_21368);
or U21509 (N_21509,N_21312,N_21287);
xor U21510 (N_21510,N_21392,N_21296);
or U21511 (N_21511,N_21251,N_21341);
and U21512 (N_21512,N_21372,N_21257);
xor U21513 (N_21513,N_21383,N_21314);
nand U21514 (N_21514,N_21369,N_21318);
xor U21515 (N_21515,N_21203,N_21392);
or U21516 (N_21516,N_21276,N_21391);
and U21517 (N_21517,N_21281,N_21304);
nand U21518 (N_21518,N_21360,N_21216);
xor U21519 (N_21519,N_21342,N_21210);
nand U21520 (N_21520,N_21254,N_21209);
or U21521 (N_21521,N_21207,N_21211);
or U21522 (N_21522,N_21355,N_21370);
nor U21523 (N_21523,N_21242,N_21290);
xor U21524 (N_21524,N_21241,N_21261);
or U21525 (N_21525,N_21283,N_21338);
xor U21526 (N_21526,N_21356,N_21390);
nor U21527 (N_21527,N_21212,N_21384);
or U21528 (N_21528,N_21211,N_21301);
and U21529 (N_21529,N_21257,N_21332);
or U21530 (N_21530,N_21274,N_21239);
nand U21531 (N_21531,N_21307,N_21248);
or U21532 (N_21532,N_21255,N_21303);
and U21533 (N_21533,N_21271,N_21285);
or U21534 (N_21534,N_21220,N_21214);
nand U21535 (N_21535,N_21375,N_21347);
xnor U21536 (N_21536,N_21261,N_21316);
or U21537 (N_21537,N_21360,N_21317);
nand U21538 (N_21538,N_21252,N_21376);
xnor U21539 (N_21539,N_21304,N_21253);
nand U21540 (N_21540,N_21344,N_21380);
nand U21541 (N_21541,N_21386,N_21323);
xor U21542 (N_21542,N_21381,N_21303);
nor U21543 (N_21543,N_21305,N_21298);
nor U21544 (N_21544,N_21206,N_21312);
or U21545 (N_21545,N_21218,N_21330);
xor U21546 (N_21546,N_21303,N_21326);
nand U21547 (N_21547,N_21288,N_21294);
and U21548 (N_21548,N_21212,N_21371);
xnor U21549 (N_21549,N_21230,N_21210);
nand U21550 (N_21550,N_21376,N_21272);
or U21551 (N_21551,N_21251,N_21350);
and U21552 (N_21552,N_21276,N_21224);
xnor U21553 (N_21553,N_21267,N_21218);
or U21554 (N_21554,N_21270,N_21223);
nor U21555 (N_21555,N_21297,N_21233);
nand U21556 (N_21556,N_21275,N_21330);
xor U21557 (N_21557,N_21221,N_21271);
nor U21558 (N_21558,N_21382,N_21368);
xnor U21559 (N_21559,N_21240,N_21279);
xnor U21560 (N_21560,N_21301,N_21246);
xor U21561 (N_21561,N_21240,N_21208);
xor U21562 (N_21562,N_21332,N_21221);
or U21563 (N_21563,N_21315,N_21214);
nand U21564 (N_21564,N_21209,N_21349);
xnor U21565 (N_21565,N_21218,N_21369);
nand U21566 (N_21566,N_21278,N_21347);
and U21567 (N_21567,N_21353,N_21266);
nor U21568 (N_21568,N_21225,N_21289);
and U21569 (N_21569,N_21222,N_21289);
or U21570 (N_21570,N_21391,N_21200);
xor U21571 (N_21571,N_21212,N_21336);
xnor U21572 (N_21572,N_21322,N_21399);
and U21573 (N_21573,N_21225,N_21318);
or U21574 (N_21574,N_21363,N_21279);
and U21575 (N_21575,N_21232,N_21306);
and U21576 (N_21576,N_21251,N_21388);
nand U21577 (N_21577,N_21338,N_21382);
xnor U21578 (N_21578,N_21353,N_21237);
and U21579 (N_21579,N_21221,N_21362);
and U21580 (N_21580,N_21284,N_21386);
and U21581 (N_21581,N_21366,N_21238);
or U21582 (N_21582,N_21382,N_21391);
xor U21583 (N_21583,N_21389,N_21256);
xor U21584 (N_21584,N_21314,N_21320);
xor U21585 (N_21585,N_21305,N_21241);
nor U21586 (N_21586,N_21391,N_21263);
nor U21587 (N_21587,N_21389,N_21329);
or U21588 (N_21588,N_21317,N_21307);
xnor U21589 (N_21589,N_21395,N_21355);
and U21590 (N_21590,N_21234,N_21221);
nor U21591 (N_21591,N_21309,N_21332);
and U21592 (N_21592,N_21213,N_21372);
nand U21593 (N_21593,N_21286,N_21292);
nor U21594 (N_21594,N_21267,N_21321);
nand U21595 (N_21595,N_21268,N_21313);
and U21596 (N_21596,N_21289,N_21294);
and U21597 (N_21597,N_21203,N_21279);
and U21598 (N_21598,N_21313,N_21224);
nand U21599 (N_21599,N_21332,N_21239);
and U21600 (N_21600,N_21568,N_21493);
xor U21601 (N_21601,N_21559,N_21509);
nand U21602 (N_21602,N_21585,N_21439);
or U21603 (N_21603,N_21553,N_21534);
or U21604 (N_21604,N_21544,N_21520);
xor U21605 (N_21605,N_21483,N_21480);
nor U21606 (N_21606,N_21589,N_21442);
and U21607 (N_21607,N_21584,N_21418);
nor U21608 (N_21608,N_21550,N_21528);
or U21609 (N_21609,N_21431,N_21463);
nand U21610 (N_21610,N_21576,N_21467);
and U21611 (N_21611,N_21411,N_21437);
xnor U21612 (N_21612,N_21432,N_21443);
and U21613 (N_21613,N_21557,N_21512);
and U21614 (N_21614,N_21539,N_21413);
xor U21615 (N_21615,N_21583,N_21598);
and U21616 (N_21616,N_21489,N_21501);
nand U21617 (N_21617,N_21516,N_21447);
or U21618 (N_21618,N_21476,N_21594);
nor U21619 (N_21619,N_21569,N_21420);
nor U21620 (N_21620,N_21435,N_21421);
or U21621 (N_21621,N_21491,N_21457);
and U21622 (N_21622,N_21441,N_21451);
and U21623 (N_21623,N_21454,N_21535);
xnor U21624 (N_21624,N_21473,N_21474);
nand U21625 (N_21625,N_21548,N_21571);
and U21626 (N_21626,N_21470,N_21472);
nor U21627 (N_21627,N_21580,N_21555);
or U21628 (N_21628,N_21401,N_21500);
and U21629 (N_21629,N_21551,N_21565);
nor U21630 (N_21630,N_21582,N_21475);
and U21631 (N_21631,N_21487,N_21547);
and U21632 (N_21632,N_21578,N_21517);
and U21633 (N_21633,N_21462,N_21567);
and U21634 (N_21634,N_21453,N_21426);
or U21635 (N_21635,N_21440,N_21566);
nand U21636 (N_21636,N_21450,N_21422);
or U21637 (N_21637,N_21419,N_21486);
nand U21638 (N_21638,N_21523,N_21504);
xor U21639 (N_21639,N_21506,N_21525);
nor U21640 (N_21640,N_21403,N_21558);
nor U21641 (N_21641,N_21524,N_21505);
nor U21642 (N_21642,N_21479,N_21529);
nor U21643 (N_21643,N_21514,N_21423);
or U21644 (N_21644,N_21495,N_21560);
or U21645 (N_21645,N_21405,N_21540);
xnor U21646 (N_21646,N_21577,N_21438);
or U21647 (N_21647,N_21446,N_21452);
and U21648 (N_21648,N_21507,N_21537);
xnor U21649 (N_21649,N_21597,N_21590);
nand U21650 (N_21650,N_21592,N_21518);
xnor U21651 (N_21651,N_21595,N_21428);
xor U21652 (N_21652,N_21496,N_21542);
xor U21653 (N_21653,N_21445,N_21427);
and U21654 (N_21654,N_21459,N_21471);
nor U21655 (N_21655,N_21564,N_21492);
xor U21656 (N_21656,N_21400,N_21466);
or U21657 (N_21657,N_21494,N_21574);
xnor U21658 (N_21658,N_21541,N_21587);
and U21659 (N_21659,N_21510,N_21490);
and U21660 (N_21660,N_21586,N_21469);
xnor U21661 (N_21661,N_21468,N_21543);
and U21662 (N_21662,N_21521,N_21465);
xnor U21663 (N_21663,N_21536,N_21460);
xor U21664 (N_21664,N_21549,N_21531);
or U21665 (N_21665,N_21407,N_21519);
nor U21666 (N_21666,N_21481,N_21449);
xnor U21667 (N_21667,N_21409,N_21458);
xnor U21668 (N_21668,N_21538,N_21497);
or U21669 (N_21669,N_21588,N_21554);
or U21670 (N_21670,N_21562,N_21570);
xor U21671 (N_21671,N_21515,N_21572);
nand U21672 (N_21672,N_21556,N_21532);
and U21673 (N_21673,N_21581,N_21415);
xnor U21674 (N_21674,N_21508,N_21546);
or U21675 (N_21675,N_21561,N_21408);
nor U21676 (N_21676,N_21436,N_21526);
nand U21677 (N_21677,N_21424,N_21429);
nor U21678 (N_21678,N_21522,N_21573);
and U21679 (N_21679,N_21414,N_21545);
nand U21680 (N_21680,N_21464,N_21513);
and U21681 (N_21681,N_21402,N_21485);
xnor U21682 (N_21682,N_21499,N_21530);
or U21683 (N_21683,N_21591,N_21579);
or U21684 (N_21684,N_21599,N_21575);
nand U21685 (N_21685,N_21593,N_21425);
xor U21686 (N_21686,N_21482,N_21448);
nor U21687 (N_21687,N_21416,N_21456);
or U21688 (N_21688,N_21478,N_21433);
nand U21689 (N_21689,N_21434,N_21498);
xor U21690 (N_21690,N_21406,N_21502);
or U21691 (N_21691,N_21484,N_21417);
nor U21692 (N_21692,N_21477,N_21527);
xnor U21693 (N_21693,N_21511,N_21410);
nand U21694 (N_21694,N_21430,N_21533);
nand U21695 (N_21695,N_21596,N_21461);
or U21696 (N_21696,N_21412,N_21455);
nor U21697 (N_21697,N_21552,N_21563);
xor U21698 (N_21698,N_21488,N_21444);
nand U21699 (N_21699,N_21503,N_21404);
and U21700 (N_21700,N_21587,N_21403);
nand U21701 (N_21701,N_21559,N_21443);
nor U21702 (N_21702,N_21541,N_21403);
xnor U21703 (N_21703,N_21407,N_21484);
xnor U21704 (N_21704,N_21445,N_21509);
or U21705 (N_21705,N_21586,N_21598);
and U21706 (N_21706,N_21450,N_21439);
xnor U21707 (N_21707,N_21527,N_21545);
xnor U21708 (N_21708,N_21443,N_21551);
nor U21709 (N_21709,N_21422,N_21426);
xnor U21710 (N_21710,N_21498,N_21541);
nand U21711 (N_21711,N_21552,N_21586);
nand U21712 (N_21712,N_21418,N_21437);
nand U21713 (N_21713,N_21429,N_21462);
nor U21714 (N_21714,N_21475,N_21497);
and U21715 (N_21715,N_21426,N_21563);
and U21716 (N_21716,N_21544,N_21555);
nor U21717 (N_21717,N_21541,N_21532);
xnor U21718 (N_21718,N_21446,N_21590);
xor U21719 (N_21719,N_21484,N_21564);
nor U21720 (N_21720,N_21430,N_21519);
xor U21721 (N_21721,N_21555,N_21436);
or U21722 (N_21722,N_21588,N_21403);
nor U21723 (N_21723,N_21562,N_21439);
xnor U21724 (N_21724,N_21599,N_21416);
xnor U21725 (N_21725,N_21442,N_21581);
nor U21726 (N_21726,N_21426,N_21502);
nand U21727 (N_21727,N_21416,N_21555);
nor U21728 (N_21728,N_21482,N_21476);
or U21729 (N_21729,N_21444,N_21443);
or U21730 (N_21730,N_21425,N_21472);
nor U21731 (N_21731,N_21559,N_21427);
xor U21732 (N_21732,N_21401,N_21451);
nor U21733 (N_21733,N_21533,N_21515);
xor U21734 (N_21734,N_21461,N_21425);
nor U21735 (N_21735,N_21429,N_21546);
or U21736 (N_21736,N_21468,N_21508);
xnor U21737 (N_21737,N_21516,N_21465);
or U21738 (N_21738,N_21486,N_21544);
or U21739 (N_21739,N_21412,N_21444);
or U21740 (N_21740,N_21447,N_21476);
xor U21741 (N_21741,N_21480,N_21545);
xnor U21742 (N_21742,N_21468,N_21536);
and U21743 (N_21743,N_21512,N_21545);
and U21744 (N_21744,N_21528,N_21446);
and U21745 (N_21745,N_21400,N_21539);
or U21746 (N_21746,N_21400,N_21583);
nand U21747 (N_21747,N_21448,N_21461);
nand U21748 (N_21748,N_21515,N_21548);
xnor U21749 (N_21749,N_21557,N_21516);
or U21750 (N_21750,N_21467,N_21520);
xnor U21751 (N_21751,N_21405,N_21452);
nand U21752 (N_21752,N_21527,N_21488);
or U21753 (N_21753,N_21437,N_21441);
and U21754 (N_21754,N_21487,N_21453);
nor U21755 (N_21755,N_21494,N_21507);
or U21756 (N_21756,N_21539,N_21432);
and U21757 (N_21757,N_21490,N_21579);
nand U21758 (N_21758,N_21556,N_21461);
nand U21759 (N_21759,N_21410,N_21459);
xor U21760 (N_21760,N_21587,N_21429);
nand U21761 (N_21761,N_21444,N_21420);
and U21762 (N_21762,N_21524,N_21414);
and U21763 (N_21763,N_21567,N_21427);
xnor U21764 (N_21764,N_21422,N_21538);
xor U21765 (N_21765,N_21566,N_21558);
and U21766 (N_21766,N_21443,N_21584);
nor U21767 (N_21767,N_21511,N_21506);
and U21768 (N_21768,N_21470,N_21415);
or U21769 (N_21769,N_21497,N_21535);
or U21770 (N_21770,N_21596,N_21444);
or U21771 (N_21771,N_21560,N_21526);
nor U21772 (N_21772,N_21577,N_21491);
and U21773 (N_21773,N_21497,N_21594);
nor U21774 (N_21774,N_21488,N_21514);
or U21775 (N_21775,N_21479,N_21516);
or U21776 (N_21776,N_21451,N_21440);
nand U21777 (N_21777,N_21501,N_21491);
nor U21778 (N_21778,N_21536,N_21458);
nand U21779 (N_21779,N_21512,N_21495);
xor U21780 (N_21780,N_21496,N_21481);
xnor U21781 (N_21781,N_21575,N_21570);
or U21782 (N_21782,N_21451,N_21448);
and U21783 (N_21783,N_21538,N_21443);
nor U21784 (N_21784,N_21464,N_21517);
nor U21785 (N_21785,N_21534,N_21456);
nand U21786 (N_21786,N_21430,N_21458);
xnor U21787 (N_21787,N_21488,N_21544);
xor U21788 (N_21788,N_21495,N_21493);
and U21789 (N_21789,N_21458,N_21564);
and U21790 (N_21790,N_21573,N_21475);
or U21791 (N_21791,N_21418,N_21449);
xor U21792 (N_21792,N_21564,N_21595);
nand U21793 (N_21793,N_21470,N_21596);
nor U21794 (N_21794,N_21463,N_21481);
nand U21795 (N_21795,N_21598,N_21454);
or U21796 (N_21796,N_21435,N_21416);
nand U21797 (N_21797,N_21527,N_21569);
nor U21798 (N_21798,N_21565,N_21423);
nand U21799 (N_21799,N_21449,N_21487);
and U21800 (N_21800,N_21619,N_21637);
nor U21801 (N_21801,N_21726,N_21663);
or U21802 (N_21802,N_21626,N_21750);
or U21803 (N_21803,N_21778,N_21790);
nor U21804 (N_21804,N_21765,N_21748);
xor U21805 (N_21805,N_21611,N_21634);
and U21806 (N_21806,N_21694,N_21719);
and U21807 (N_21807,N_21775,N_21666);
nand U21808 (N_21808,N_21799,N_21785);
nand U21809 (N_21809,N_21733,N_21728);
nand U21810 (N_21810,N_21624,N_21673);
nand U21811 (N_21811,N_21758,N_21668);
and U21812 (N_21812,N_21695,N_21732);
nor U21813 (N_21813,N_21630,N_21772);
nor U21814 (N_21814,N_21740,N_21621);
and U21815 (N_21815,N_21690,N_21780);
and U21816 (N_21816,N_21771,N_21784);
and U21817 (N_21817,N_21704,N_21777);
and U21818 (N_21818,N_21672,N_21706);
and U21819 (N_21819,N_21741,N_21703);
xor U21820 (N_21820,N_21607,N_21769);
or U21821 (N_21821,N_21757,N_21752);
nand U21822 (N_21822,N_21656,N_21720);
xnor U21823 (N_21823,N_21646,N_21761);
nor U21824 (N_21824,N_21675,N_21691);
nand U21825 (N_21825,N_21718,N_21699);
or U21826 (N_21826,N_21682,N_21725);
or U21827 (N_21827,N_21601,N_21749);
or U21828 (N_21828,N_21796,N_21755);
or U21829 (N_21829,N_21709,N_21665);
nor U21830 (N_21830,N_21716,N_21684);
and U21831 (N_21831,N_21677,N_21683);
or U21832 (N_21832,N_21746,N_21667);
xnor U21833 (N_21833,N_21658,N_21625);
nor U21834 (N_21834,N_21620,N_21734);
or U21835 (N_21835,N_21711,N_21707);
nor U21836 (N_21836,N_21710,N_21743);
and U21837 (N_21837,N_21693,N_21680);
nand U21838 (N_21838,N_21788,N_21617);
and U21839 (N_21839,N_21652,N_21739);
or U21840 (N_21840,N_21708,N_21701);
or U21841 (N_21841,N_21687,N_21659);
xnor U21842 (N_21842,N_21615,N_21633);
and U21843 (N_21843,N_21787,N_21635);
and U21844 (N_21844,N_21618,N_21688);
nor U21845 (N_21845,N_21730,N_21721);
or U21846 (N_21846,N_21797,N_21767);
nand U21847 (N_21847,N_21671,N_21770);
or U21848 (N_21848,N_21763,N_21715);
and U21849 (N_21849,N_21766,N_21760);
nor U21850 (N_21850,N_21674,N_21657);
nand U21851 (N_21851,N_21696,N_21794);
xnor U21852 (N_21852,N_21622,N_21664);
nor U21853 (N_21853,N_21782,N_21705);
xor U21854 (N_21854,N_21735,N_21698);
nor U21855 (N_21855,N_21616,N_21722);
nand U21856 (N_21856,N_21729,N_21639);
or U21857 (N_21857,N_21774,N_21650);
nor U21858 (N_21858,N_21603,N_21713);
nor U21859 (N_21859,N_21742,N_21795);
xnor U21860 (N_21860,N_21655,N_21638);
nand U21861 (N_21861,N_21662,N_21712);
or U21862 (N_21862,N_21644,N_21613);
nor U21863 (N_21863,N_21737,N_21793);
and U21864 (N_21864,N_21602,N_21627);
and U21865 (N_21865,N_21679,N_21681);
nand U21866 (N_21866,N_21643,N_21689);
nor U21867 (N_21867,N_21653,N_21632);
and U21868 (N_21868,N_21628,N_21600);
or U21869 (N_21869,N_21764,N_21636);
xnor U21870 (N_21870,N_21669,N_21744);
nor U21871 (N_21871,N_21731,N_21647);
xor U21872 (N_21872,N_21605,N_21612);
or U21873 (N_21873,N_21651,N_21609);
xor U21874 (N_21874,N_21783,N_21623);
or U21875 (N_21875,N_21727,N_21745);
and U21876 (N_21876,N_21686,N_21645);
and U21877 (N_21877,N_21604,N_21676);
nor U21878 (N_21878,N_21702,N_21738);
or U21879 (N_21879,N_21660,N_21762);
and U21880 (N_21880,N_21786,N_21700);
or U21881 (N_21881,N_21779,N_21792);
nand U21882 (N_21882,N_21606,N_21723);
and U21883 (N_21883,N_21717,N_21631);
xor U21884 (N_21884,N_21751,N_21798);
and U21885 (N_21885,N_21754,N_21608);
nor U21886 (N_21886,N_21648,N_21642);
nor U21887 (N_21887,N_21649,N_21789);
nand U21888 (N_21888,N_21753,N_21697);
or U21889 (N_21889,N_21614,N_21610);
and U21890 (N_21890,N_21692,N_21781);
xor U21891 (N_21891,N_21654,N_21629);
nand U21892 (N_21892,N_21776,N_21736);
and U21893 (N_21893,N_21773,N_21641);
or U21894 (N_21894,N_21724,N_21670);
nand U21895 (N_21895,N_21747,N_21791);
and U21896 (N_21896,N_21661,N_21759);
or U21897 (N_21897,N_21640,N_21685);
and U21898 (N_21898,N_21714,N_21756);
xnor U21899 (N_21899,N_21768,N_21678);
and U21900 (N_21900,N_21722,N_21675);
nand U21901 (N_21901,N_21613,N_21702);
and U21902 (N_21902,N_21683,N_21601);
xor U21903 (N_21903,N_21742,N_21663);
and U21904 (N_21904,N_21631,N_21694);
and U21905 (N_21905,N_21691,N_21604);
xnor U21906 (N_21906,N_21606,N_21731);
or U21907 (N_21907,N_21737,N_21786);
or U21908 (N_21908,N_21730,N_21619);
and U21909 (N_21909,N_21685,N_21730);
nand U21910 (N_21910,N_21747,N_21671);
or U21911 (N_21911,N_21716,N_21650);
and U21912 (N_21912,N_21608,N_21679);
and U21913 (N_21913,N_21635,N_21753);
nand U21914 (N_21914,N_21728,N_21707);
and U21915 (N_21915,N_21675,N_21679);
or U21916 (N_21916,N_21634,N_21665);
or U21917 (N_21917,N_21745,N_21746);
xnor U21918 (N_21918,N_21699,N_21750);
nand U21919 (N_21919,N_21773,N_21697);
or U21920 (N_21920,N_21647,N_21712);
xnor U21921 (N_21921,N_21731,N_21611);
nand U21922 (N_21922,N_21736,N_21752);
or U21923 (N_21923,N_21723,N_21650);
nand U21924 (N_21924,N_21667,N_21668);
and U21925 (N_21925,N_21626,N_21735);
and U21926 (N_21926,N_21629,N_21796);
and U21927 (N_21927,N_21695,N_21701);
or U21928 (N_21928,N_21658,N_21768);
nand U21929 (N_21929,N_21743,N_21671);
nor U21930 (N_21930,N_21699,N_21667);
nor U21931 (N_21931,N_21693,N_21731);
and U21932 (N_21932,N_21695,N_21739);
and U21933 (N_21933,N_21711,N_21605);
or U21934 (N_21934,N_21665,N_21763);
or U21935 (N_21935,N_21644,N_21715);
xor U21936 (N_21936,N_21746,N_21729);
xor U21937 (N_21937,N_21684,N_21679);
nor U21938 (N_21938,N_21772,N_21782);
nand U21939 (N_21939,N_21693,N_21647);
nor U21940 (N_21940,N_21673,N_21733);
nand U21941 (N_21941,N_21710,N_21629);
nor U21942 (N_21942,N_21629,N_21760);
or U21943 (N_21943,N_21666,N_21679);
nor U21944 (N_21944,N_21606,N_21798);
and U21945 (N_21945,N_21653,N_21670);
nand U21946 (N_21946,N_21784,N_21742);
or U21947 (N_21947,N_21601,N_21615);
or U21948 (N_21948,N_21731,N_21745);
nand U21949 (N_21949,N_21649,N_21625);
or U21950 (N_21950,N_21720,N_21689);
and U21951 (N_21951,N_21766,N_21790);
nand U21952 (N_21952,N_21605,N_21626);
nand U21953 (N_21953,N_21626,N_21718);
xor U21954 (N_21954,N_21664,N_21653);
xor U21955 (N_21955,N_21786,N_21649);
or U21956 (N_21956,N_21633,N_21674);
or U21957 (N_21957,N_21682,N_21786);
or U21958 (N_21958,N_21657,N_21715);
or U21959 (N_21959,N_21627,N_21767);
nand U21960 (N_21960,N_21654,N_21743);
nand U21961 (N_21961,N_21680,N_21753);
nor U21962 (N_21962,N_21733,N_21616);
xor U21963 (N_21963,N_21667,N_21634);
xor U21964 (N_21964,N_21650,N_21771);
xor U21965 (N_21965,N_21690,N_21683);
and U21966 (N_21966,N_21735,N_21614);
nand U21967 (N_21967,N_21739,N_21740);
xor U21968 (N_21968,N_21667,N_21665);
or U21969 (N_21969,N_21769,N_21707);
xor U21970 (N_21970,N_21704,N_21628);
or U21971 (N_21971,N_21746,N_21734);
nor U21972 (N_21972,N_21663,N_21756);
nor U21973 (N_21973,N_21648,N_21678);
and U21974 (N_21974,N_21704,N_21720);
and U21975 (N_21975,N_21733,N_21678);
nand U21976 (N_21976,N_21774,N_21667);
or U21977 (N_21977,N_21748,N_21681);
nor U21978 (N_21978,N_21751,N_21709);
xnor U21979 (N_21979,N_21655,N_21615);
and U21980 (N_21980,N_21630,N_21729);
xor U21981 (N_21981,N_21692,N_21667);
or U21982 (N_21982,N_21628,N_21725);
nand U21983 (N_21983,N_21601,N_21719);
or U21984 (N_21984,N_21728,N_21702);
or U21985 (N_21985,N_21644,N_21659);
or U21986 (N_21986,N_21760,N_21707);
and U21987 (N_21987,N_21685,N_21710);
xor U21988 (N_21988,N_21617,N_21757);
nor U21989 (N_21989,N_21627,N_21649);
or U21990 (N_21990,N_21659,N_21764);
nand U21991 (N_21991,N_21759,N_21788);
or U21992 (N_21992,N_21622,N_21641);
xor U21993 (N_21993,N_21696,N_21634);
nor U21994 (N_21994,N_21627,N_21714);
or U21995 (N_21995,N_21613,N_21655);
or U21996 (N_21996,N_21706,N_21754);
and U21997 (N_21997,N_21744,N_21619);
and U21998 (N_21998,N_21785,N_21719);
nand U21999 (N_21999,N_21724,N_21690);
or U22000 (N_22000,N_21969,N_21864);
xnor U22001 (N_22001,N_21824,N_21987);
nand U22002 (N_22002,N_21833,N_21996);
nand U22003 (N_22003,N_21809,N_21863);
or U22004 (N_22004,N_21953,N_21975);
nor U22005 (N_22005,N_21949,N_21837);
or U22006 (N_22006,N_21925,N_21828);
or U22007 (N_22007,N_21961,N_21872);
xnor U22008 (N_22008,N_21825,N_21859);
and U22009 (N_22009,N_21867,N_21808);
nor U22010 (N_22010,N_21955,N_21951);
nand U22011 (N_22011,N_21906,N_21998);
and U22012 (N_22012,N_21973,N_21899);
xor U22013 (N_22013,N_21964,N_21818);
nor U22014 (N_22014,N_21845,N_21986);
xnor U22015 (N_22015,N_21822,N_21880);
nor U22016 (N_22016,N_21983,N_21991);
and U22017 (N_22017,N_21963,N_21815);
xor U22018 (N_22018,N_21958,N_21908);
xnor U22019 (N_22019,N_21870,N_21854);
nor U22020 (N_22020,N_21890,N_21976);
or U22021 (N_22021,N_21971,N_21993);
nor U22022 (N_22022,N_21974,N_21873);
nor U22023 (N_22023,N_21928,N_21915);
nor U22024 (N_22024,N_21930,N_21823);
and U22025 (N_22025,N_21940,N_21924);
and U22026 (N_22026,N_21840,N_21947);
xnor U22027 (N_22027,N_21935,N_21972);
or U22028 (N_22028,N_21826,N_21843);
xnor U22029 (N_22029,N_21865,N_21851);
and U22030 (N_22030,N_21838,N_21813);
nand U22031 (N_22031,N_21876,N_21897);
xnor U22032 (N_22032,N_21909,N_21978);
nand U22033 (N_22033,N_21831,N_21962);
and U22034 (N_22034,N_21861,N_21920);
xnor U22035 (N_22035,N_21927,N_21904);
and U22036 (N_22036,N_21878,N_21835);
and U22037 (N_22037,N_21802,N_21800);
and U22038 (N_22038,N_21913,N_21981);
or U22039 (N_22039,N_21919,N_21979);
xor U22040 (N_22040,N_21892,N_21852);
nor U22041 (N_22041,N_21807,N_21803);
and U22042 (N_22042,N_21887,N_21966);
xor U22043 (N_22043,N_21944,N_21846);
and U22044 (N_22044,N_21860,N_21844);
nor U22045 (N_22045,N_21805,N_21967);
xnor U22046 (N_22046,N_21894,N_21985);
xor U22047 (N_22047,N_21888,N_21942);
and U22048 (N_22048,N_21862,N_21934);
xor U22049 (N_22049,N_21801,N_21938);
nor U22050 (N_22050,N_21885,N_21902);
nand U22051 (N_22051,N_21914,N_21917);
nor U22052 (N_22052,N_21907,N_21893);
nand U22053 (N_22053,N_21817,N_21901);
xor U22054 (N_22054,N_21950,N_21946);
or U22055 (N_22055,N_21956,N_21900);
nand U22056 (N_22056,N_21933,N_21857);
or U22057 (N_22057,N_21877,N_21905);
nand U22058 (N_22058,N_21980,N_21999);
nor U22059 (N_22059,N_21995,N_21994);
or U22060 (N_22060,N_21959,N_21882);
and U22061 (N_22061,N_21891,N_21936);
nor U22062 (N_22062,N_21960,N_21937);
nand U22063 (N_22063,N_21977,N_21957);
nand U22064 (N_22064,N_21886,N_21952);
nand U22065 (N_22065,N_21889,N_21911);
nor U22066 (N_22066,N_21821,N_21839);
xnor U22067 (N_22067,N_21879,N_21997);
and U22068 (N_22068,N_21820,N_21847);
and U22069 (N_22069,N_21984,N_21881);
nand U22070 (N_22070,N_21834,N_21939);
nor U22071 (N_22071,N_21806,N_21968);
and U22072 (N_22072,N_21829,N_21856);
nand U22073 (N_22073,N_21912,N_21812);
nand U22074 (N_22074,N_21884,N_21842);
or U22075 (N_22075,N_21903,N_21875);
nand U22076 (N_22076,N_21868,N_21841);
xnor U22077 (N_22077,N_21954,N_21988);
nand U22078 (N_22078,N_21895,N_21943);
and U22079 (N_22079,N_21921,N_21910);
nand U22080 (N_22080,N_21926,N_21932);
or U22081 (N_22081,N_21811,N_21853);
nand U22082 (N_22082,N_21970,N_21896);
and U22083 (N_22083,N_21830,N_21836);
xnor U22084 (N_22084,N_21858,N_21827);
xnor U22085 (N_22085,N_21990,N_21814);
or U22086 (N_22086,N_21850,N_21810);
xnor U22087 (N_22087,N_21869,N_21931);
nand U22088 (N_22088,N_21832,N_21923);
nor U22089 (N_22089,N_21918,N_21922);
and U22090 (N_22090,N_21916,N_21992);
or U22091 (N_22091,N_21945,N_21804);
nand U22092 (N_22092,N_21819,N_21929);
nor U22093 (N_22093,N_21874,N_21849);
nand U22094 (N_22094,N_21866,N_21871);
xor U22095 (N_22095,N_21989,N_21855);
nand U22096 (N_22096,N_21982,N_21941);
nand U22097 (N_22097,N_21948,N_21848);
nand U22098 (N_22098,N_21965,N_21898);
xor U22099 (N_22099,N_21816,N_21883);
or U22100 (N_22100,N_21856,N_21830);
nand U22101 (N_22101,N_21960,N_21991);
xor U22102 (N_22102,N_21875,N_21987);
nand U22103 (N_22103,N_21982,N_21997);
nand U22104 (N_22104,N_21925,N_21829);
nand U22105 (N_22105,N_21819,N_21956);
nor U22106 (N_22106,N_21955,N_21898);
xnor U22107 (N_22107,N_21932,N_21987);
nand U22108 (N_22108,N_21838,N_21967);
nand U22109 (N_22109,N_21982,N_21939);
nor U22110 (N_22110,N_21903,N_21979);
nand U22111 (N_22111,N_21850,N_21987);
xnor U22112 (N_22112,N_21841,N_21940);
and U22113 (N_22113,N_21983,N_21990);
xor U22114 (N_22114,N_21883,N_21948);
and U22115 (N_22115,N_21826,N_21960);
xor U22116 (N_22116,N_21966,N_21932);
xor U22117 (N_22117,N_21992,N_21900);
or U22118 (N_22118,N_21841,N_21873);
nand U22119 (N_22119,N_21916,N_21898);
nand U22120 (N_22120,N_21847,N_21874);
nand U22121 (N_22121,N_21994,N_21931);
and U22122 (N_22122,N_21930,N_21962);
and U22123 (N_22123,N_21976,N_21809);
and U22124 (N_22124,N_21870,N_21820);
xnor U22125 (N_22125,N_21869,N_21897);
nand U22126 (N_22126,N_21892,N_21936);
or U22127 (N_22127,N_21977,N_21867);
and U22128 (N_22128,N_21924,N_21927);
nand U22129 (N_22129,N_21949,N_21981);
nor U22130 (N_22130,N_21937,N_21905);
nand U22131 (N_22131,N_21975,N_21851);
nor U22132 (N_22132,N_21869,N_21915);
or U22133 (N_22133,N_21876,N_21906);
and U22134 (N_22134,N_21978,N_21870);
nor U22135 (N_22135,N_21813,N_21847);
nand U22136 (N_22136,N_21893,N_21814);
nor U22137 (N_22137,N_21846,N_21982);
or U22138 (N_22138,N_21922,N_21906);
xnor U22139 (N_22139,N_21810,N_21895);
xor U22140 (N_22140,N_21868,N_21854);
xor U22141 (N_22141,N_21821,N_21892);
nor U22142 (N_22142,N_21952,N_21945);
or U22143 (N_22143,N_21856,N_21827);
nand U22144 (N_22144,N_21946,N_21999);
xnor U22145 (N_22145,N_21861,N_21889);
nor U22146 (N_22146,N_21899,N_21894);
or U22147 (N_22147,N_21905,N_21942);
xor U22148 (N_22148,N_21953,N_21853);
nor U22149 (N_22149,N_21967,N_21941);
xnor U22150 (N_22150,N_21927,N_21996);
nor U22151 (N_22151,N_21840,N_21845);
and U22152 (N_22152,N_21949,N_21982);
nand U22153 (N_22153,N_21953,N_21814);
and U22154 (N_22154,N_21986,N_21959);
nand U22155 (N_22155,N_21834,N_21994);
xor U22156 (N_22156,N_21991,N_21998);
xor U22157 (N_22157,N_21828,N_21958);
or U22158 (N_22158,N_21929,N_21817);
xnor U22159 (N_22159,N_21822,N_21998);
and U22160 (N_22160,N_21933,N_21831);
or U22161 (N_22161,N_21984,N_21945);
nor U22162 (N_22162,N_21884,N_21902);
xnor U22163 (N_22163,N_21910,N_21889);
nor U22164 (N_22164,N_21993,N_21997);
xor U22165 (N_22165,N_21846,N_21905);
xor U22166 (N_22166,N_21938,N_21841);
nand U22167 (N_22167,N_21830,N_21945);
and U22168 (N_22168,N_21811,N_21837);
or U22169 (N_22169,N_21825,N_21919);
nand U22170 (N_22170,N_21845,N_21966);
xor U22171 (N_22171,N_21816,N_21935);
nand U22172 (N_22172,N_21832,N_21825);
and U22173 (N_22173,N_21961,N_21847);
xor U22174 (N_22174,N_21848,N_21895);
or U22175 (N_22175,N_21851,N_21906);
and U22176 (N_22176,N_21963,N_21938);
xor U22177 (N_22177,N_21826,N_21870);
nand U22178 (N_22178,N_21943,N_21874);
xor U22179 (N_22179,N_21971,N_21981);
or U22180 (N_22180,N_21874,N_21833);
or U22181 (N_22181,N_21939,N_21956);
nor U22182 (N_22182,N_21877,N_21837);
and U22183 (N_22183,N_21898,N_21921);
nor U22184 (N_22184,N_21918,N_21936);
xnor U22185 (N_22185,N_21826,N_21941);
xnor U22186 (N_22186,N_21903,N_21916);
nand U22187 (N_22187,N_21940,N_21926);
nand U22188 (N_22188,N_21883,N_21934);
xor U22189 (N_22189,N_21877,N_21835);
xor U22190 (N_22190,N_21863,N_21942);
or U22191 (N_22191,N_21989,N_21839);
or U22192 (N_22192,N_21873,N_21803);
nand U22193 (N_22193,N_21904,N_21962);
and U22194 (N_22194,N_21935,N_21907);
xnor U22195 (N_22195,N_21833,N_21987);
nand U22196 (N_22196,N_21992,N_21847);
and U22197 (N_22197,N_21815,N_21834);
nand U22198 (N_22198,N_21850,N_21960);
xnor U22199 (N_22199,N_21961,N_21838);
or U22200 (N_22200,N_22068,N_22045);
nand U22201 (N_22201,N_22098,N_22016);
or U22202 (N_22202,N_22177,N_22165);
nand U22203 (N_22203,N_22151,N_22019);
nor U22204 (N_22204,N_22195,N_22064);
and U22205 (N_22205,N_22182,N_22010);
and U22206 (N_22206,N_22158,N_22100);
nand U22207 (N_22207,N_22198,N_22154);
and U22208 (N_22208,N_22136,N_22172);
xor U22209 (N_22209,N_22189,N_22128);
nand U22210 (N_22210,N_22022,N_22051);
nor U22211 (N_22211,N_22117,N_22109);
and U22212 (N_22212,N_22017,N_22197);
or U22213 (N_22213,N_22075,N_22078);
nor U22214 (N_22214,N_22114,N_22112);
xor U22215 (N_22215,N_22031,N_22148);
or U22216 (N_22216,N_22169,N_22080);
xnor U22217 (N_22217,N_22036,N_22027);
nor U22218 (N_22218,N_22171,N_22183);
or U22219 (N_22219,N_22086,N_22059);
and U22220 (N_22220,N_22181,N_22192);
nor U22221 (N_22221,N_22155,N_22140);
and U22222 (N_22222,N_22186,N_22161);
xor U22223 (N_22223,N_22138,N_22089);
nor U22224 (N_22224,N_22105,N_22190);
and U22225 (N_22225,N_22118,N_22162);
nand U22226 (N_22226,N_22091,N_22127);
nand U22227 (N_22227,N_22099,N_22054);
nor U22228 (N_22228,N_22006,N_22170);
or U22229 (N_22229,N_22005,N_22048);
nand U22230 (N_22230,N_22053,N_22133);
or U22231 (N_22231,N_22088,N_22057);
nand U22232 (N_22232,N_22095,N_22050);
or U22233 (N_22233,N_22084,N_22153);
or U22234 (N_22234,N_22168,N_22087);
xnor U22235 (N_22235,N_22119,N_22063);
and U22236 (N_22236,N_22156,N_22163);
nand U22237 (N_22237,N_22038,N_22061);
and U22238 (N_22238,N_22055,N_22145);
nor U22239 (N_22239,N_22094,N_22188);
or U22240 (N_22240,N_22160,N_22101);
and U22241 (N_22241,N_22003,N_22150);
and U22242 (N_22242,N_22026,N_22139);
nand U22243 (N_22243,N_22009,N_22049);
xor U22244 (N_22244,N_22060,N_22073);
or U22245 (N_22245,N_22129,N_22015);
and U22246 (N_22246,N_22137,N_22144);
nand U22247 (N_22247,N_22028,N_22146);
and U22248 (N_22248,N_22074,N_22108);
nand U22249 (N_22249,N_22130,N_22135);
nor U22250 (N_22250,N_22093,N_22012);
nand U22251 (N_22251,N_22167,N_22187);
nand U22252 (N_22252,N_22029,N_22081);
xor U22253 (N_22253,N_22030,N_22143);
or U22254 (N_22254,N_22041,N_22040);
nand U22255 (N_22255,N_22157,N_22024);
nand U22256 (N_22256,N_22076,N_22196);
nor U22257 (N_22257,N_22120,N_22107);
xor U22258 (N_22258,N_22032,N_22152);
nor U22259 (N_22259,N_22072,N_22065);
nand U22260 (N_22260,N_22037,N_22001);
or U22261 (N_22261,N_22132,N_22007);
and U22262 (N_22262,N_22176,N_22142);
xor U22263 (N_22263,N_22173,N_22193);
nor U22264 (N_22264,N_22166,N_22020);
nor U22265 (N_22265,N_22033,N_22077);
and U22266 (N_22266,N_22069,N_22046);
or U22267 (N_22267,N_22175,N_22134);
nor U22268 (N_22268,N_22199,N_22115);
nand U22269 (N_22269,N_22110,N_22062);
xor U22270 (N_22270,N_22083,N_22131);
or U22271 (N_22271,N_22071,N_22174);
xnor U22272 (N_22272,N_22004,N_22021);
and U22273 (N_22273,N_22124,N_22122);
nand U22274 (N_22274,N_22191,N_22066);
or U22275 (N_22275,N_22178,N_22116);
nor U22276 (N_22276,N_22000,N_22149);
nor U22277 (N_22277,N_22018,N_22070);
and U22278 (N_22278,N_22097,N_22103);
nor U22279 (N_22279,N_22047,N_22104);
nand U22280 (N_22280,N_22023,N_22025);
xor U22281 (N_22281,N_22008,N_22002);
nor U22282 (N_22282,N_22111,N_22164);
xnor U22283 (N_22283,N_22052,N_22147);
or U22284 (N_22284,N_22014,N_22184);
nand U22285 (N_22285,N_22067,N_22044);
and U22286 (N_22286,N_22042,N_22125);
or U22287 (N_22287,N_22096,N_22058);
xor U22288 (N_22288,N_22113,N_22034);
xor U22289 (N_22289,N_22092,N_22043);
nor U22290 (N_22290,N_22123,N_22102);
nor U22291 (N_22291,N_22179,N_22194);
xnor U22292 (N_22292,N_22121,N_22013);
xor U22293 (N_22293,N_22090,N_22011);
or U22294 (N_22294,N_22126,N_22180);
nand U22295 (N_22295,N_22185,N_22085);
and U22296 (N_22296,N_22039,N_22056);
xor U22297 (N_22297,N_22106,N_22079);
xor U22298 (N_22298,N_22141,N_22159);
nor U22299 (N_22299,N_22035,N_22082);
or U22300 (N_22300,N_22138,N_22158);
xor U22301 (N_22301,N_22112,N_22125);
and U22302 (N_22302,N_22136,N_22063);
xnor U22303 (N_22303,N_22002,N_22144);
or U22304 (N_22304,N_22152,N_22039);
or U22305 (N_22305,N_22181,N_22153);
or U22306 (N_22306,N_22167,N_22184);
nor U22307 (N_22307,N_22051,N_22126);
and U22308 (N_22308,N_22180,N_22140);
nand U22309 (N_22309,N_22029,N_22091);
and U22310 (N_22310,N_22063,N_22188);
or U22311 (N_22311,N_22016,N_22133);
nand U22312 (N_22312,N_22138,N_22174);
nand U22313 (N_22313,N_22100,N_22148);
xor U22314 (N_22314,N_22110,N_22026);
nor U22315 (N_22315,N_22065,N_22133);
or U22316 (N_22316,N_22107,N_22179);
xnor U22317 (N_22317,N_22061,N_22174);
nand U22318 (N_22318,N_22179,N_22121);
and U22319 (N_22319,N_22027,N_22196);
and U22320 (N_22320,N_22129,N_22152);
nor U22321 (N_22321,N_22090,N_22032);
or U22322 (N_22322,N_22172,N_22022);
xor U22323 (N_22323,N_22059,N_22166);
nand U22324 (N_22324,N_22158,N_22140);
nor U22325 (N_22325,N_22126,N_22056);
nor U22326 (N_22326,N_22154,N_22087);
nand U22327 (N_22327,N_22028,N_22033);
and U22328 (N_22328,N_22021,N_22162);
and U22329 (N_22329,N_22146,N_22150);
nand U22330 (N_22330,N_22176,N_22084);
and U22331 (N_22331,N_22156,N_22127);
nand U22332 (N_22332,N_22194,N_22020);
xnor U22333 (N_22333,N_22129,N_22130);
xor U22334 (N_22334,N_22091,N_22156);
or U22335 (N_22335,N_22138,N_22098);
nand U22336 (N_22336,N_22147,N_22025);
and U22337 (N_22337,N_22179,N_22061);
nor U22338 (N_22338,N_22020,N_22183);
or U22339 (N_22339,N_22100,N_22080);
nor U22340 (N_22340,N_22065,N_22002);
nor U22341 (N_22341,N_22178,N_22017);
and U22342 (N_22342,N_22072,N_22195);
nand U22343 (N_22343,N_22088,N_22087);
or U22344 (N_22344,N_22046,N_22012);
xnor U22345 (N_22345,N_22065,N_22131);
xor U22346 (N_22346,N_22111,N_22187);
and U22347 (N_22347,N_22164,N_22046);
and U22348 (N_22348,N_22080,N_22182);
xor U22349 (N_22349,N_22114,N_22124);
nor U22350 (N_22350,N_22063,N_22083);
xor U22351 (N_22351,N_22093,N_22057);
nor U22352 (N_22352,N_22026,N_22089);
nand U22353 (N_22353,N_22127,N_22089);
or U22354 (N_22354,N_22199,N_22077);
nand U22355 (N_22355,N_22191,N_22196);
xnor U22356 (N_22356,N_22119,N_22074);
or U22357 (N_22357,N_22060,N_22129);
and U22358 (N_22358,N_22192,N_22021);
nor U22359 (N_22359,N_22124,N_22164);
xor U22360 (N_22360,N_22022,N_22156);
nor U22361 (N_22361,N_22183,N_22074);
nor U22362 (N_22362,N_22195,N_22061);
nor U22363 (N_22363,N_22111,N_22087);
nor U22364 (N_22364,N_22047,N_22116);
nor U22365 (N_22365,N_22006,N_22145);
or U22366 (N_22366,N_22024,N_22137);
and U22367 (N_22367,N_22079,N_22160);
nand U22368 (N_22368,N_22021,N_22026);
nand U22369 (N_22369,N_22191,N_22033);
nor U22370 (N_22370,N_22072,N_22114);
and U22371 (N_22371,N_22035,N_22020);
nor U22372 (N_22372,N_22009,N_22138);
or U22373 (N_22373,N_22162,N_22166);
nand U22374 (N_22374,N_22093,N_22067);
and U22375 (N_22375,N_22047,N_22024);
xor U22376 (N_22376,N_22038,N_22022);
nand U22377 (N_22377,N_22030,N_22127);
nand U22378 (N_22378,N_22114,N_22037);
xor U22379 (N_22379,N_22111,N_22015);
and U22380 (N_22380,N_22137,N_22187);
and U22381 (N_22381,N_22128,N_22155);
nor U22382 (N_22382,N_22043,N_22135);
xnor U22383 (N_22383,N_22160,N_22170);
nor U22384 (N_22384,N_22143,N_22087);
xor U22385 (N_22385,N_22105,N_22065);
xor U22386 (N_22386,N_22167,N_22174);
xnor U22387 (N_22387,N_22006,N_22077);
xor U22388 (N_22388,N_22116,N_22191);
nand U22389 (N_22389,N_22037,N_22121);
nor U22390 (N_22390,N_22084,N_22104);
or U22391 (N_22391,N_22117,N_22042);
and U22392 (N_22392,N_22013,N_22103);
nand U22393 (N_22393,N_22026,N_22187);
nor U22394 (N_22394,N_22027,N_22163);
or U22395 (N_22395,N_22079,N_22168);
or U22396 (N_22396,N_22062,N_22127);
and U22397 (N_22397,N_22028,N_22067);
nor U22398 (N_22398,N_22184,N_22030);
or U22399 (N_22399,N_22184,N_22013);
nand U22400 (N_22400,N_22201,N_22285);
nor U22401 (N_22401,N_22355,N_22324);
nand U22402 (N_22402,N_22340,N_22257);
xor U22403 (N_22403,N_22336,N_22327);
xnor U22404 (N_22404,N_22305,N_22227);
or U22405 (N_22405,N_22319,N_22322);
nand U22406 (N_22406,N_22398,N_22291);
nor U22407 (N_22407,N_22213,N_22241);
or U22408 (N_22408,N_22205,N_22343);
nand U22409 (N_22409,N_22278,N_22234);
xor U22410 (N_22410,N_22335,N_22240);
or U22411 (N_22411,N_22255,N_22202);
or U22412 (N_22412,N_22269,N_22390);
or U22413 (N_22413,N_22308,N_22245);
nor U22414 (N_22414,N_22207,N_22215);
nor U22415 (N_22415,N_22366,N_22273);
and U22416 (N_22416,N_22365,N_22231);
nor U22417 (N_22417,N_22353,N_22381);
or U22418 (N_22418,N_22356,N_22393);
xor U22419 (N_22419,N_22362,N_22239);
and U22420 (N_22420,N_22237,N_22375);
and U22421 (N_22421,N_22272,N_22345);
or U22422 (N_22422,N_22391,N_22303);
or U22423 (N_22423,N_22317,N_22320);
nand U22424 (N_22424,N_22251,N_22265);
nand U22425 (N_22425,N_22312,N_22352);
or U22426 (N_22426,N_22395,N_22211);
nand U22427 (N_22427,N_22309,N_22318);
nand U22428 (N_22428,N_22329,N_22293);
or U22429 (N_22429,N_22268,N_22388);
nand U22430 (N_22430,N_22330,N_22263);
or U22431 (N_22431,N_22208,N_22337);
and U22432 (N_22432,N_22292,N_22382);
xor U22433 (N_22433,N_22229,N_22399);
and U22434 (N_22434,N_22321,N_22304);
or U22435 (N_22435,N_22252,N_22367);
nor U22436 (N_22436,N_22221,N_22378);
or U22437 (N_22437,N_22235,N_22346);
xnor U22438 (N_22438,N_22228,N_22332);
nor U22439 (N_22439,N_22282,N_22220);
nand U22440 (N_22440,N_22383,N_22357);
xor U22441 (N_22441,N_22219,N_22225);
xnor U22442 (N_22442,N_22204,N_22253);
xnor U22443 (N_22443,N_22328,N_22379);
and U22444 (N_22444,N_22325,N_22230);
nand U22445 (N_22445,N_22250,N_22364);
or U22446 (N_22446,N_22358,N_22350);
nand U22447 (N_22447,N_22370,N_22311);
nand U22448 (N_22448,N_22259,N_22316);
and U22449 (N_22449,N_22323,N_22396);
nor U22450 (N_22450,N_22274,N_22386);
nor U22451 (N_22451,N_22217,N_22286);
or U22452 (N_22452,N_22310,N_22315);
and U22453 (N_22453,N_22348,N_22384);
nor U22454 (N_22454,N_22376,N_22244);
and U22455 (N_22455,N_22294,N_22218);
nor U22456 (N_22456,N_22203,N_22333);
and U22457 (N_22457,N_22387,N_22279);
nand U22458 (N_22458,N_22214,N_22296);
or U22459 (N_22459,N_22372,N_22297);
nor U22460 (N_22460,N_22361,N_22385);
and U22461 (N_22461,N_22209,N_22280);
nor U22462 (N_22462,N_22363,N_22397);
and U22463 (N_22463,N_22249,N_22306);
xnor U22464 (N_22464,N_22256,N_22258);
and U22465 (N_22465,N_22264,N_22314);
or U22466 (N_22466,N_22206,N_22301);
or U22467 (N_22467,N_22248,N_22283);
nand U22468 (N_22468,N_22226,N_22359);
nor U22469 (N_22469,N_22254,N_22392);
nor U22470 (N_22470,N_22289,N_22295);
and U22471 (N_22471,N_22290,N_22284);
or U22472 (N_22472,N_22373,N_22300);
or U22473 (N_22473,N_22313,N_22270);
nor U22474 (N_22474,N_22281,N_22267);
or U22475 (N_22475,N_22339,N_22354);
and U22476 (N_22476,N_22371,N_22334);
or U22477 (N_22477,N_22238,N_22298);
and U22478 (N_22478,N_22380,N_22275);
and U22479 (N_22479,N_22351,N_22266);
and U22480 (N_22480,N_22224,N_22277);
nor U22481 (N_22481,N_22342,N_22338);
or U22482 (N_22482,N_22242,N_22246);
xor U22483 (N_22483,N_22276,N_22223);
xor U22484 (N_22484,N_22271,N_22377);
nor U22485 (N_22485,N_22233,N_22216);
or U22486 (N_22486,N_22307,N_22287);
nand U22487 (N_22487,N_22299,N_22200);
and U22488 (N_22488,N_22344,N_22261);
and U22489 (N_22489,N_22262,N_22302);
xor U22490 (N_22490,N_22260,N_22247);
or U22491 (N_22491,N_22394,N_22232);
or U22492 (N_22492,N_22389,N_22369);
xor U22493 (N_22493,N_22236,N_22341);
or U22494 (N_22494,N_22326,N_22212);
xnor U22495 (N_22495,N_22210,N_22347);
or U22496 (N_22496,N_22288,N_22349);
nor U22497 (N_22497,N_22374,N_22368);
nor U22498 (N_22498,N_22331,N_22222);
nor U22499 (N_22499,N_22243,N_22360);
nor U22500 (N_22500,N_22313,N_22332);
and U22501 (N_22501,N_22284,N_22208);
nor U22502 (N_22502,N_22218,N_22372);
nand U22503 (N_22503,N_22358,N_22347);
or U22504 (N_22504,N_22211,N_22203);
and U22505 (N_22505,N_22270,N_22348);
or U22506 (N_22506,N_22275,N_22298);
nand U22507 (N_22507,N_22300,N_22397);
and U22508 (N_22508,N_22242,N_22308);
nor U22509 (N_22509,N_22384,N_22388);
xor U22510 (N_22510,N_22251,N_22206);
nor U22511 (N_22511,N_22221,N_22280);
nand U22512 (N_22512,N_22313,N_22316);
xnor U22513 (N_22513,N_22376,N_22334);
or U22514 (N_22514,N_22237,N_22320);
xor U22515 (N_22515,N_22208,N_22299);
nor U22516 (N_22516,N_22393,N_22305);
or U22517 (N_22517,N_22291,N_22375);
xor U22518 (N_22518,N_22349,N_22242);
nor U22519 (N_22519,N_22307,N_22221);
xnor U22520 (N_22520,N_22274,N_22318);
nand U22521 (N_22521,N_22348,N_22353);
and U22522 (N_22522,N_22318,N_22254);
xor U22523 (N_22523,N_22291,N_22294);
nor U22524 (N_22524,N_22373,N_22348);
or U22525 (N_22525,N_22329,N_22328);
nor U22526 (N_22526,N_22202,N_22219);
and U22527 (N_22527,N_22307,N_22262);
nor U22528 (N_22528,N_22228,N_22277);
and U22529 (N_22529,N_22362,N_22368);
nand U22530 (N_22530,N_22230,N_22362);
nor U22531 (N_22531,N_22229,N_22306);
nand U22532 (N_22532,N_22383,N_22253);
or U22533 (N_22533,N_22336,N_22204);
xor U22534 (N_22534,N_22282,N_22322);
or U22535 (N_22535,N_22222,N_22232);
nand U22536 (N_22536,N_22236,N_22366);
xnor U22537 (N_22537,N_22208,N_22372);
xnor U22538 (N_22538,N_22326,N_22256);
or U22539 (N_22539,N_22200,N_22317);
xor U22540 (N_22540,N_22329,N_22279);
or U22541 (N_22541,N_22334,N_22323);
xor U22542 (N_22542,N_22281,N_22243);
or U22543 (N_22543,N_22302,N_22377);
nor U22544 (N_22544,N_22297,N_22321);
or U22545 (N_22545,N_22277,N_22360);
and U22546 (N_22546,N_22373,N_22260);
or U22547 (N_22547,N_22378,N_22365);
nand U22548 (N_22548,N_22201,N_22391);
nand U22549 (N_22549,N_22298,N_22288);
and U22550 (N_22550,N_22383,N_22298);
nand U22551 (N_22551,N_22333,N_22367);
xnor U22552 (N_22552,N_22290,N_22364);
nand U22553 (N_22553,N_22349,N_22304);
nand U22554 (N_22554,N_22339,N_22246);
nor U22555 (N_22555,N_22296,N_22377);
nand U22556 (N_22556,N_22278,N_22297);
xor U22557 (N_22557,N_22356,N_22357);
and U22558 (N_22558,N_22251,N_22275);
nor U22559 (N_22559,N_22340,N_22216);
nor U22560 (N_22560,N_22378,N_22206);
and U22561 (N_22561,N_22301,N_22394);
nor U22562 (N_22562,N_22221,N_22354);
nor U22563 (N_22563,N_22202,N_22226);
nand U22564 (N_22564,N_22226,N_22221);
nor U22565 (N_22565,N_22270,N_22356);
nor U22566 (N_22566,N_22385,N_22274);
nand U22567 (N_22567,N_22387,N_22334);
nor U22568 (N_22568,N_22385,N_22266);
nand U22569 (N_22569,N_22293,N_22309);
xnor U22570 (N_22570,N_22316,N_22324);
and U22571 (N_22571,N_22212,N_22276);
or U22572 (N_22572,N_22395,N_22335);
and U22573 (N_22573,N_22252,N_22246);
nor U22574 (N_22574,N_22344,N_22275);
nand U22575 (N_22575,N_22389,N_22315);
or U22576 (N_22576,N_22214,N_22375);
and U22577 (N_22577,N_22270,N_22364);
xor U22578 (N_22578,N_22350,N_22328);
nor U22579 (N_22579,N_22336,N_22273);
nor U22580 (N_22580,N_22331,N_22233);
nand U22581 (N_22581,N_22337,N_22295);
xnor U22582 (N_22582,N_22222,N_22272);
and U22583 (N_22583,N_22277,N_22333);
nor U22584 (N_22584,N_22330,N_22304);
xnor U22585 (N_22585,N_22266,N_22229);
xor U22586 (N_22586,N_22278,N_22240);
nor U22587 (N_22587,N_22338,N_22230);
xor U22588 (N_22588,N_22370,N_22350);
nand U22589 (N_22589,N_22357,N_22271);
or U22590 (N_22590,N_22277,N_22318);
nand U22591 (N_22591,N_22277,N_22227);
xor U22592 (N_22592,N_22348,N_22241);
nand U22593 (N_22593,N_22379,N_22281);
xnor U22594 (N_22594,N_22258,N_22288);
nand U22595 (N_22595,N_22364,N_22238);
nor U22596 (N_22596,N_22202,N_22261);
and U22597 (N_22597,N_22286,N_22296);
and U22598 (N_22598,N_22266,N_22364);
and U22599 (N_22599,N_22271,N_22296);
and U22600 (N_22600,N_22460,N_22438);
nand U22601 (N_22601,N_22409,N_22401);
xnor U22602 (N_22602,N_22442,N_22462);
and U22603 (N_22603,N_22465,N_22546);
nor U22604 (N_22604,N_22530,N_22564);
nor U22605 (N_22605,N_22585,N_22524);
nand U22606 (N_22606,N_22556,N_22533);
and U22607 (N_22607,N_22563,N_22466);
and U22608 (N_22608,N_22547,N_22405);
and U22609 (N_22609,N_22505,N_22554);
xor U22610 (N_22610,N_22486,N_22481);
xnor U22611 (N_22611,N_22436,N_22592);
and U22612 (N_22612,N_22537,N_22518);
or U22613 (N_22613,N_22421,N_22484);
nand U22614 (N_22614,N_22557,N_22503);
and U22615 (N_22615,N_22569,N_22539);
nand U22616 (N_22616,N_22572,N_22425);
or U22617 (N_22617,N_22440,N_22517);
and U22618 (N_22618,N_22415,N_22595);
and U22619 (N_22619,N_22534,N_22561);
or U22620 (N_22620,N_22548,N_22587);
xor U22621 (N_22621,N_22452,N_22558);
or U22622 (N_22622,N_22568,N_22454);
nand U22623 (N_22623,N_22506,N_22448);
and U22624 (N_22624,N_22566,N_22528);
and U22625 (N_22625,N_22471,N_22497);
and U22626 (N_22626,N_22535,N_22426);
nor U22627 (N_22627,N_22428,N_22514);
or U22628 (N_22628,N_22461,N_22458);
and U22629 (N_22629,N_22437,N_22483);
or U22630 (N_22630,N_22487,N_22589);
and U22631 (N_22631,N_22499,N_22498);
nor U22632 (N_22632,N_22420,N_22526);
xor U22633 (N_22633,N_22555,N_22473);
nand U22634 (N_22634,N_22532,N_22418);
xor U22635 (N_22635,N_22404,N_22495);
xor U22636 (N_22636,N_22504,N_22485);
xnor U22637 (N_22637,N_22540,N_22450);
xor U22638 (N_22638,N_22411,N_22463);
nor U22639 (N_22639,N_22449,N_22576);
or U22640 (N_22640,N_22553,N_22480);
nor U22641 (N_22641,N_22477,N_22416);
nand U22642 (N_22642,N_22523,N_22599);
nor U22643 (N_22643,N_22493,N_22408);
nor U22644 (N_22644,N_22544,N_22451);
xnor U22645 (N_22645,N_22542,N_22446);
or U22646 (N_22646,N_22527,N_22422);
or U22647 (N_22647,N_22513,N_22406);
xor U22648 (N_22648,N_22434,N_22522);
and U22649 (N_22649,N_22444,N_22489);
or U22650 (N_22650,N_22536,N_22476);
xnor U22651 (N_22651,N_22464,N_22516);
xor U22652 (N_22652,N_22457,N_22580);
nor U22653 (N_22653,N_22431,N_22511);
nor U22654 (N_22654,N_22562,N_22570);
nand U22655 (N_22655,N_22492,N_22456);
nor U22656 (N_22656,N_22445,N_22551);
or U22657 (N_22657,N_22591,N_22560);
nand U22658 (N_22658,N_22565,N_22413);
xnor U22659 (N_22659,N_22575,N_22496);
nor U22660 (N_22660,N_22494,N_22472);
nand U22661 (N_22661,N_22597,N_22470);
and U22662 (N_22662,N_22482,N_22593);
xor U22663 (N_22663,N_22598,N_22543);
xor U22664 (N_22664,N_22531,N_22468);
and U22665 (N_22665,N_22419,N_22478);
nand U22666 (N_22666,N_22512,N_22501);
xor U22667 (N_22667,N_22400,N_22578);
xor U22668 (N_22668,N_22529,N_22509);
xor U22669 (N_22669,N_22594,N_22402);
and U22670 (N_22670,N_22525,N_22521);
and U22671 (N_22671,N_22488,N_22520);
and U22672 (N_22672,N_22441,N_22459);
or U22673 (N_22673,N_22475,N_22577);
nor U22674 (N_22674,N_22549,N_22574);
or U22675 (N_22675,N_22455,N_22467);
or U22676 (N_22676,N_22586,N_22453);
xnor U22677 (N_22677,N_22507,N_22491);
xor U22678 (N_22678,N_22510,N_22469);
nand U22679 (N_22679,N_22545,N_22559);
nor U22680 (N_22680,N_22582,N_22579);
xnor U22681 (N_22681,N_22412,N_22417);
xnor U22682 (N_22682,N_22541,N_22474);
xor U22683 (N_22683,N_22439,N_22519);
or U22684 (N_22684,N_22430,N_22424);
nand U22685 (N_22685,N_22573,N_22410);
or U22686 (N_22686,N_22414,N_22584);
or U22687 (N_22687,N_22588,N_22552);
and U22688 (N_22688,N_22407,N_22508);
xor U22689 (N_22689,N_22567,N_22429);
nand U22690 (N_22690,N_22479,N_22500);
nand U22691 (N_22691,N_22432,N_22423);
nand U22692 (N_22692,N_22427,N_22581);
or U22693 (N_22693,N_22490,N_22590);
nor U22694 (N_22694,N_22550,N_22502);
nand U22695 (N_22695,N_22538,N_22443);
xnor U22696 (N_22696,N_22433,N_22447);
nand U22697 (N_22697,N_22583,N_22403);
and U22698 (N_22698,N_22571,N_22435);
nand U22699 (N_22699,N_22596,N_22515);
and U22700 (N_22700,N_22433,N_22506);
and U22701 (N_22701,N_22474,N_22531);
nor U22702 (N_22702,N_22597,N_22531);
and U22703 (N_22703,N_22588,N_22487);
nor U22704 (N_22704,N_22586,N_22441);
nand U22705 (N_22705,N_22570,N_22587);
xnor U22706 (N_22706,N_22506,N_22522);
and U22707 (N_22707,N_22406,N_22565);
nand U22708 (N_22708,N_22481,N_22580);
and U22709 (N_22709,N_22517,N_22454);
and U22710 (N_22710,N_22486,N_22432);
and U22711 (N_22711,N_22525,N_22454);
and U22712 (N_22712,N_22584,N_22514);
nand U22713 (N_22713,N_22500,N_22416);
nand U22714 (N_22714,N_22546,N_22489);
nand U22715 (N_22715,N_22468,N_22503);
or U22716 (N_22716,N_22591,N_22542);
nor U22717 (N_22717,N_22554,N_22475);
nand U22718 (N_22718,N_22460,N_22472);
nand U22719 (N_22719,N_22472,N_22456);
nand U22720 (N_22720,N_22575,N_22415);
nor U22721 (N_22721,N_22483,N_22541);
or U22722 (N_22722,N_22507,N_22404);
xor U22723 (N_22723,N_22525,N_22506);
and U22724 (N_22724,N_22480,N_22589);
nor U22725 (N_22725,N_22485,N_22511);
xor U22726 (N_22726,N_22419,N_22405);
nand U22727 (N_22727,N_22457,N_22419);
xnor U22728 (N_22728,N_22430,N_22403);
xor U22729 (N_22729,N_22578,N_22540);
and U22730 (N_22730,N_22550,N_22533);
xnor U22731 (N_22731,N_22559,N_22590);
and U22732 (N_22732,N_22424,N_22487);
nor U22733 (N_22733,N_22558,N_22518);
and U22734 (N_22734,N_22462,N_22407);
xor U22735 (N_22735,N_22489,N_22434);
nand U22736 (N_22736,N_22528,N_22555);
and U22737 (N_22737,N_22523,N_22475);
xor U22738 (N_22738,N_22546,N_22432);
nand U22739 (N_22739,N_22492,N_22573);
or U22740 (N_22740,N_22433,N_22408);
or U22741 (N_22741,N_22518,N_22493);
nor U22742 (N_22742,N_22525,N_22529);
xnor U22743 (N_22743,N_22453,N_22430);
or U22744 (N_22744,N_22460,N_22544);
nand U22745 (N_22745,N_22544,N_22582);
and U22746 (N_22746,N_22491,N_22479);
and U22747 (N_22747,N_22569,N_22517);
nor U22748 (N_22748,N_22557,N_22581);
nor U22749 (N_22749,N_22487,N_22437);
nand U22750 (N_22750,N_22488,N_22455);
nor U22751 (N_22751,N_22453,N_22428);
or U22752 (N_22752,N_22410,N_22539);
and U22753 (N_22753,N_22594,N_22581);
and U22754 (N_22754,N_22490,N_22466);
nor U22755 (N_22755,N_22420,N_22466);
nor U22756 (N_22756,N_22447,N_22554);
and U22757 (N_22757,N_22464,N_22420);
nor U22758 (N_22758,N_22477,N_22438);
and U22759 (N_22759,N_22445,N_22466);
nand U22760 (N_22760,N_22565,N_22522);
nand U22761 (N_22761,N_22589,N_22427);
or U22762 (N_22762,N_22592,N_22504);
and U22763 (N_22763,N_22455,N_22578);
nor U22764 (N_22764,N_22595,N_22561);
or U22765 (N_22765,N_22478,N_22524);
or U22766 (N_22766,N_22574,N_22474);
xnor U22767 (N_22767,N_22509,N_22533);
nor U22768 (N_22768,N_22557,N_22586);
nor U22769 (N_22769,N_22482,N_22477);
or U22770 (N_22770,N_22515,N_22439);
xnor U22771 (N_22771,N_22484,N_22467);
or U22772 (N_22772,N_22441,N_22571);
or U22773 (N_22773,N_22428,N_22468);
or U22774 (N_22774,N_22419,N_22431);
nand U22775 (N_22775,N_22492,N_22560);
nand U22776 (N_22776,N_22553,N_22565);
and U22777 (N_22777,N_22469,N_22464);
xor U22778 (N_22778,N_22472,N_22544);
or U22779 (N_22779,N_22537,N_22569);
nor U22780 (N_22780,N_22438,N_22587);
nand U22781 (N_22781,N_22528,N_22456);
nand U22782 (N_22782,N_22504,N_22560);
or U22783 (N_22783,N_22408,N_22402);
xnor U22784 (N_22784,N_22435,N_22590);
nand U22785 (N_22785,N_22507,N_22550);
nand U22786 (N_22786,N_22414,N_22456);
or U22787 (N_22787,N_22543,N_22564);
and U22788 (N_22788,N_22483,N_22596);
or U22789 (N_22789,N_22560,N_22417);
or U22790 (N_22790,N_22590,N_22521);
nor U22791 (N_22791,N_22566,N_22450);
nor U22792 (N_22792,N_22492,N_22433);
nand U22793 (N_22793,N_22504,N_22487);
nand U22794 (N_22794,N_22488,N_22538);
or U22795 (N_22795,N_22448,N_22485);
and U22796 (N_22796,N_22496,N_22566);
or U22797 (N_22797,N_22433,N_22457);
and U22798 (N_22798,N_22495,N_22420);
and U22799 (N_22799,N_22570,N_22402);
or U22800 (N_22800,N_22653,N_22770);
xor U22801 (N_22801,N_22796,N_22722);
xnor U22802 (N_22802,N_22740,N_22704);
nand U22803 (N_22803,N_22714,N_22658);
xnor U22804 (N_22804,N_22792,N_22616);
and U22805 (N_22805,N_22764,N_22759);
and U22806 (N_22806,N_22647,N_22628);
or U22807 (N_22807,N_22638,N_22679);
nand U22808 (N_22808,N_22600,N_22717);
nand U22809 (N_22809,N_22785,N_22729);
and U22810 (N_22810,N_22701,N_22753);
xor U22811 (N_22811,N_22716,N_22705);
nor U22812 (N_22812,N_22604,N_22786);
nand U22813 (N_22813,N_22718,N_22681);
and U22814 (N_22814,N_22707,N_22766);
and U22815 (N_22815,N_22648,N_22755);
xnor U22816 (N_22816,N_22745,N_22635);
and U22817 (N_22817,N_22685,N_22692);
or U22818 (N_22818,N_22769,N_22708);
or U22819 (N_22819,N_22735,N_22671);
and U22820 (N_22820,N_22631,N_22694);
or U22821 (N_22821,N_22683,N_22746);
nor U22822 (N_22822,N_22656,N_22602);
nand U22823 (N_22823,N_22737,N_22601);
xnor U22824 (N_22824,N_22742,N_22646);
xor U22825 (N_22825,N_22621,N_22787);
and U22826 (N_22826,N_22605,N_22726);
nand U22827 (N_22827,N_22623,N_22669);
and U22828 (N_22828,N_22762,N_22613);
or U22829 (N_22829,N_22733,N_22677);
nor U22830 (N_22830,N_22629,N_22676);
or U22831 (N_22831,N_22696,N_22715);
and U22832 (N_22832,N_22781,N_22667);
and U22833 (N_22833,N_22773,N_22614);
and U22834 (N_22834,N_22761,N_22754);
nand U22835 (N_22835,N_22727,N_22642);
and U22836 (N_22836,N_22651,N_22657);
and U22837 (N_22837,N_22712,N_22702);
nand U22838 (N_22838,N_22695,N_22663);
or U22839 (N_22839,N_22797,N_22768);
xnor U22840 (N_22840,N_22636,N_22720);
nor U22841 (N_22841,N_22672,N_22641);
and U22842 (N_22842,N_22738,N_22661);
nor U22843 (N_22843,N_22783,N_22778);
nand U22844 (N_22844,N_22721,N_22609);
and U22845 (N_22845,N_22758,N_22739);
xor U22846 (N_22846,N_22619,N_22650);
and U22847 (N_22847,N_22706,N_22782);
nand U22848 (N_22848,N_22674,N_22730);
nand U22849 (N_22849,N_22625,N_22713);
xnor U22850 (N_22850,N_22666,N_22637);
xnor U22851 (N_22851,N_22734,N_22678);
xnor U22852 (N_22852,N_22607,N_22662);
nand U22853 (N_22853,N_22618,N_22644);
xor U22854 (N_22854,N_22624,N_22699);
and U22855 (N_22855,N_22675,N_22691);
or U22856 (N_22856,N_22728,N_22686);
or U22857 (N_22857,N_22756,N_22794);
nor U22858 (N_22858,N_22767,N_22789);
nor U22859 (N_22859,N_22795,N_22757);
nor U22860 (N_22860,N_22649,N_22788);
xnor U22861 (N_22861,N_22611,N_22670);
or U22862 (N_22862,N_22682,N_22655);
or U22863 (N_22863,N_22645,N_22765);
nor U22864 (N_22864,N_22747,N_22774);
xnor U22865 (N_22865,N_22640,N_22689);
nor U22866 (N_22866,N_22606,N_22731);
xnor U22867 (N_22867,N_22603,N_22622);
and U22868 (N_22868,N_22700,N_22608);
or U22869 (N_22869,N_22684,N_22724);
and U22870 (N_22870,N_22643,N_22634);
and U22871 (N_22871,N_22620,N_22749);
and U22872 (N_22872,N_22752,N_22710);
or U22873 (N_22873,N_22776,N_22617);
or U22874 (N_22874,N_22741,N_22652);
or U22875 (N_22875,N_22772,N_22748);
nand U22876 (N_22876,N_22784,N_22698);
and U22877 (N_22877,N_22743,N_22630);
or U22878 (N_22878,N_22751,N_22639);
xor U22879 (N_22879,N_22690,N_22771);
nor U22880 (N_22880,N_22687,N_22711);
or U22881 (N_22881,N_22668,N_22632);
nor U22882 (N_22882,N_22719,N_22779);
xnor U22883 (N_22883,N_22732,N_22610);
nor U22884 (N_22884,N_22697,N_22760);
nor U22885 (N_22885,N_22703,N_22709);
and U22886 (N_22886,N_22780,N_22664);
nor U22887 (N_22887,N_22723,N_22799);
and U22888 (N_22888,N_22654,N_22660);
nor U22889 (N_22889,N_22633,N_22612);
or U22890 (N_22890,N_22688,N_22673);
xor U22891 (N_22891,N_22626,N_22790);
nor U22892 (N_22892,N_22763,N_22750);
nor U22893 (N_22893,N_22736,N_22680);
nor U22894 (N_22894,N_22793,N_22659);
xnor U22895 (N_22895,N_22775,N_22665);
nor U22896 (N_22896,N_22725,N_22777);
nand U22897 (N_22897,N_22693,N_22791);
nor U22898 (N_22898,N_22798,N_22744);
and U22899 (N_22899,N_22615,N_22627);
xor U22900 (N_22900,N_22627,N_22665);
nand U22901 (N_22901,N_22647,N_22722);
nand U22902 (N_22902,N_22718,N_22743);
nand U22903 (N_22903,N_22620,N_22698);
or U22904 (N_22904,N_22792,N_22663);
nand U22905 (N_22905,N_22700,N_22740);
xnor U22906 (N_22906,N_22665,N_22684);
and U22907 (N_22907,N_22643,N_22703);
xnor U22908 (N_22908,N_22755,N_22708);
or U22909 (N_22909,N_22777,N_22748);
nor U22910 (N_22910,N_22602,N_22725);
and U22911 (N_22911,N_22666,N_22784);
and U22912 (N_22912,N_22612,N_22724);
xor U22913 (N_22913,N_22654,N_22793);
xor U22914 (N_22914,N_22708,N_22746);
nor U22915 (N_22915,N_22743,N_22784);
and U22916 (N_22916,N_22666,N_22710);
or U22917 (N_22917,N_22739,N_22680);
nor U22918 (N_22918,N_22792,N_22764);
nor U22919 (N_22919,N_22646,N_22745);
nor U22920 (N_22920,N_22733,N_22685);
xnor U22921 (N_22921,N_22629,N_22699);
nand U22922 (N_22922,N_22694,N_22664);
or U22923 (N_22923,N_22600,N_22652);
nor U22924 (N_22924,N_22685,N_22638);
or U22925 (N_22925,N_22634,N_22714);
nor U22926 (N_22926,N_22757,N_22644);
and U22927 (N_22927,N_22727,N_22610);
nor U22928 (N_22928,N_22759,N_22708);
nor U22929 (N_22929,N_22631,N_22677);
or U22930 (N_22930,N_22615,N_22748);
and U22931 (N_22931,N_22774,N_22607);
and U22932 (N_22932,N_22726,N_22610);
or U22933 (N_22933,N_22692,N_22719);
nor U22934 (N_22934,N_22711,N_22699);
xor U22935 (N_22935,N_22698,N_22628);
nand U22936 (N_22936,N_22740,N_22776);
or U22937 (N_22937,N_22668,N_22758);
and U22938 (N_22938,N_22785,N_22646);
xor U22939 (N_22939,N_22616,N_22759);
nor U22940 (N_22940,N_22645,N_22611);
or U22941 (N_22941,N_22756,N_22665);
or U22942 (N_22942,N_22641,N_22755);
nor U22943 (N_22943,N_22634,N_22604);
xnor U22944 (N_22944,N_22686,N_22616);
nand U22945 (N_22945,N_22724,N_22727);
and U22946 (N_22946,N_22662,N_22671);
or U22947 (N_22947,N_22605,N_22714);
and U22948 (N_22948,N_22792,N_22734);
and U22949 (N_22949,N_22737,N_22615);
xnor U22950 (N_22950,N_22707,N_22705);
or U22951 (N_22951,N_22727,N_22791);
or U22952 (N_22952,N_22783,N_22648);
and U22953 (N_22953,N_22726,N_22628);
nand U22954 (N_22954,N_22670,N_22675);
nand U22955 (N_22955,N_22640,N_22708);
and U22956 (N_22956,N_22621,N_22632);
or U22957 (N_22957,N_22674,N_22753);
nand U22958 (N_22958,N_22610,N_22729);
nand U22959 (N_22959,N_22644,N_22745);
and U22960 (N_22960,N_22764,N_22610);
nand U22961 (N_22961,N_22694,N_22790);
nor U22962 (N_22962,N_22602,N_22696);
or U22963 (N_22963,N_22617,N_22741);
and U22964 (N_22964,N_22606,N_22783);
xor U22965 (N_22965,N_22663,N_22607);
and U22966 (N_22966,N_22748,N_22698);
and U22967 (N_22967,N_22698,N_22683);
nor U22968 (N_22968,N_22753,N_22626);
nand U22969 (N_22969,N_22705,N_22781);
xor U22970 (N_22970,N_22728,N_22665);
nand U22971 (N_22971,N_22609,N_22723);
and U22972 (N_22972,N_22678,N_22766);
nor U22973 (N_22973,N_22718,N_22774);
xnor U22974 (N_22974,N_22730,N_22664);
or U22975 (N_22975,N_22790,N_22781);
xor U22976 (N_22976,N_22763,N_22690);
nor U22977 (N_22977,N_22742,N_22781);
nand U22978 (N_22978,N_22729,N_22741);
nor U22979 (N_22979,N_22600,N_22734);
nand U22980 (N_22980,N_22679,N_22640);
or U22981 (N_22981,N_22603,N_22743);
xnor U22982 (N_22982,N_22656,N_22724);
xor U22983 (N_22983,N_22650,N_22615);
xnor U22984 (N_22984,N_22642,N_22636);
xnor U22985 (N_22985,N_22711,N_22629);
nor U22986 (N_22986,N_22781,N_22786);
nand U22987 (N_22987,N_22752,N_22648);
nand U22988 (N_22988,N_22773,N_22630);
xnor U22989 (N_22989,N_22794,N_22730);
nor U22990 (N_22990,N_22686,N_22678);
nand U22991 (N_22991,N_22604,N_22727);
xnor U22992 (N_22992,N_22614,N_22721);
and U22993 (N_22993,N_22760,N_22734);
or U22994 (N_22994,N_22779,N_22765);
or U22995 (N_22995,N_22756,N_22644);
or U22996 (N_22996,N_22641,N_22766);
and U22997 (N_22997,N_22781,N_22798);
nand U22998 (N_22998,N_22657,N_22703);
and U22999 (N_22999,N_22738,N_22788);
xor U23000 (N_23000,N_22875,N_22961);
nor U23001 (N_23001,N_22858,N_22982);
nand U23002 (N_23002,N_22897,N_22890);
nor U23003 (N_23003,N_22811,N_22851);
xnor U23004 (N_23004,N_22817,N_22845);
nand U23005 (N_23005,N_22885,N_22848);
or U23006 (N_23006,N_22988,N_22912);
xnor U23007 (N_23007,N_22867,N_22878);
xnor U23008 (N_23008,N_22972,N_22866);
xnor U23009 (N_23009,N_22944,N_22911);
xor U23010 (N_23010,N_22828,N_22929);
xor U23011 (N_23011,N_22870,N_22913);
nor U23012 (N_23012,N_22914,N_22903);
or U23013 (N_23013,N_22987,N_22951);
and U23014 (N_23014,N_22806,N_22801);
or U23015 (N_23015,N_22985,N_22871);
nand U23016 (N_23016,N_22962,N_22927);
nor U23017 (N_23017,N_22937,N_22821);
nor U23018 (N_23018,N_22835,N_22926);
or U23019 (N_23019,N_22983,N_22833);
xor U23020 (N_23020,N_22876,N_22984);
nor U23021 (N_23021,N_22831,N_22886);
nor U23022 (N_23022,N_22933,N_22949);
and U23023 (N_23023,N_22919,N_22992);
nand U23024 (N_23024,N_22869,N_22935);
and U23025 (N_23025,N_22946,N_22888);
xor U23026 (N_23026,N_22953,N_22840);
and U23027 (N_23027,N_22896,N_22923);
or U23028 (N_23028,N_22857,N_22930);
and U23029 (N_23029,N_22938,N_22980);
or U23030 (N_23030,N_22809,N_22824);
or U23031 (N_23031,N_22884,N_22877);
and U23032 (N_23032,N_22964,N_22852);
xor U23033 (N_23033,N_22823,N_22856);
nand U23034 (N_23034,N_22808,N_22943);
and U23035 (N_23035,N_22805,N_22922);
nand U23036 (N_23036,N_22844,N_22874);
nor U23037 (N_23037,N_22853,N_22999);
xor U23038 (N_23038,N_22901,N_22873);
nor U23039 (N_23039,N_22822,N_22836);
and U23040 (N_23040,N_22918,N_22893);
xnor U23041 (N_23041,N_22803,N_22975);
xnor U23042 (N_23042,N_22861,N_22954);
nor U23043 (N_23043,N_22849,N_22994);
and U23044 (N_23044,N_22966,N_22978);
and U23045 (N_23045,N_22997,N_22963);
or U23046 (N_23046,N_22932,N_22924);
or U23047 (N_23047,N_22965,N_22991);
or U23048 (N_23048,N_22902,N_22958);
nor U23049 (N_23049,N_22925,N_22906);
nor U23050 (N_23050,N_22855,N_22812);
nand U23051 (N_23051,N_22976,N_22820);
nand U23052 (N_23052,N_22928,N_22862);
nor U23053 (N_23053,N_22940,N_22904);
nor U23054 (N_23054,N_22957,N_22860);
and U23055 (N_23055,N_22910,N_22971);
nor U23056 (N_23056,N_22981,N_22838);
nand U23057 (N_23057,N_22917,N_22825);
or U23058 (N_23058,N_22947,N_22899);
nand U23059 (N_23059,N_22883,N_22815);
and U23060 (N_23060,N_22939,N_22810);
nand U23061 (N_23061,N_22967,N_22955);
nand U23062 (N_23062,N_22892,N_22931);
and U23063 (N_23063,N_22936,N_22863);
or U23064 (N_23064,N_22916,N_22802);
and U23065 (N_23065,N_22841,N_22909);
nand U23066 (N_23066,N_22882,N_22819);
nor U23067 (N_23067,N_22830,N_22859);
or U23068 (N_23068,N_22968,N_22843);
or U23069 (N_23069,N_22813,N_22864);
nor U23070 (N_23070,N_22837,N_22887);
nand U23071 (N_23071,N_22974,N_22894);
nor U23072 (N_23072,N_22827,N_22990);
and U23073 (N_23073,N_22847,N_22832);
and U23074 (N_23074,N_22977,N_22814);
nand U23075 (N_23075,N_22986,N_22979);
nor U23076 (N_23076,N_22891,N_22872);
xor U23077 (N_23077,N_22834,N_22842);
xnor U23078 (N_23078,N_22804,N_22948);
nor U23079 (N_23079,N_22816,N_22942);
and U23080 (N_23080,N_22959,N_22895);
nor U23081 (N_23081,N_22915,N_22846);
xnor U23082 (N_23082,N_22865,N_22839);
or U23083 (N_23083,N_22970,N_22945);
nor U23084 (N_23084,N_22941,N_22969);
nor U23085 (N_23085,N_22960,N_22868);
xor U23086 (N_23086,N_22900,N_22818);
nor U23087 (N_23087,N_22934,N_22993);
nand U23088 (N_23088,N_22989,N_22998);
and U23089 (N_23089,N_22854,N_22879);
and U23090 (N_23090,N_22956,N_22905);
nor U23091 (N_23091,N_22807,N_22898);
nand U23092 (N_23092,N_22973,N_22920);
nand U23093 (N_23093,N_22921,N_22850);
or U23094 (N_23094,N_22829,N_22907);
nand U23095 (N_23095,N_22950,N_22908);
xor U23096 (N_23096,N_22881,N_22995);
nor U23097 (N_23097,N_22952,N_22880);
xnor U23098 (N_23098,N_22826,N_22800);
xor U23099 (N_23099,N_22996,N_22889);
nor U23100 (N_23100,N_22845,N_22969);
nor U23101 (N_23101,N_22972,N_22881);
or U23102 (N_23102,N_22800,N_22926);
xor U23103 (N_23103,N_22932,N_22893);
and U23104 (N_23104,N_22848,N_22836);
and U23105 (N_23105,N_22915,N_22983);
nor U23106 (N_23106,N_22809,N_22904);
or U23107 (N_23107,N_22935,N_22985);
or U23108 (N_23108,N_22843,N_22989);
and U23109 (N_23109,N_22875,N_22827);
or U23110 (N_23110,N_22962,N_22902);
xnor U23111 (N_23111,N_22992,N_22817);
or U23112 (N_23112,N_22838,N_22925);
nor U23113 (N_23113,N_22816,N_22940);
nor U23114 (N_23114,N_22850,N_22914);
and U23115 (N_23115,N_22982,N_22913);
nor U23116 (N_23116,N_22824,N_22841);
or U23117 (N_23117,N_22878,N_22917);
or U23118 (N_23118,N_22912,N_22985);
and U23119 (N_23119,N_22949,N_22881);
nor U23120 (N_23120,N_22966,N_22899);
xor U23121 (N_23121,N_22855,N_22879);
xor U23122 (N_23122,N_22895,N_22974);
nor U23123 (N_23123,N_22908,N_22865);
or U23124 (N_23124,N_22964,N_22965);
nand U23125 (N_23125,N_22852,N_22919);
or U23126 (N_23126,N_22962,N_22839);
and U23127 (N_23127,N_22981,N_22853);
nand U23128 (N_23128,N_22991,N_22828);
and U23129 (N_23129,N_22805,N_22840);
nand U23130 (N_23130,N_22855,N_22945);
xnor U23131 (N_23131,N_22976,N_22984);
and U23132 (N_23132,N_22896,N_22990);
and U23133 (N_23133,N_22859,N_22826);
and U23134 (N_23134,N_22943,N_22955);
and U23135 (N_23135,N_22974,N_22932);
nor U23136 (N_23136,N_22832,N_22841);
or U23137 (N_23137,N_22854,N_22919);
or U23138 (N_23138,N_22900,N_22809);
and U23139 (N_23139,N_22845,N_22830);
nand U23140 (N_23140,N_22976,N_22919);
nor U23141 (N_23141,N_22855,N_22971);
xnor U23142 (N_23142,N_22854,N_22909);
xor U23143 (N_23143,N_22879,N_22919);
nand U23144 (N_23144,N_22814,N_22933);
xor U23145 (N_23145,N_22894,N_22833);
nor U23146 (N_23146,N_22864,N_22892);
and U23147 (N_23147,N_22992,N_22941);
xor U23148 (N_23148,N_22834,N_22839);
nand U23149 (N_23149,N_22926,N_22878);
nor U23150 (N_23150,N_22953,N_22956);
xor U23151 (N_23151,N_22968,N_22926);
or U23152 (N_23152,N_22918,N_22842);
nor U23153 (N_23153,N_22959,N_22914);
nor U23154 (N_23154,N_22941,N_22931);
nand U23155 (N_23155,N_22875,N_22877);
xnor U23156 (N_23156,N_22966,N_22827);
nor U23157 (N_23157,N_22943,N_22917);
or U23158 (N_23158,N_22832,N_22807);
and U23159 (N_23159,N_22852,N_22829);
and U23160 (N_23160,N_22853,N_22984);
xnor U23161 (N_23161,N_22809,N_22958);
xor U23162 (N_23162,N_22876,N_22995);
or U23163 (N_23163,N_22832,N_22963);
nor U23164 (N_23164,N_22825,N_22818);
nand U23165 (N_23165,N_22949,N_22912);
or U23166 (N_23166,N_22919,N_22800);
or U23167 (N_23167,N_22842,N_22893);
or U23168 (N_23168,N_22920,N_22961);
xor U23169 (N_23169,N_22957,N_22997);
nand U23170 (N_23170,N_22968,N_22831);
and U23171 (N_23171,N_22850,N_22989);
or U23172 (N_23172,N_22910,N_22815);
or U23173 (N_23173,N_22889,N_22869);
nand U23174 (N_23174,N_22952,N_22999);
xnor U23175 (N_23175,N_22931,N_22814);
xor U23176 (N_23176,N_22918,N_22968);
nand U23177 (N_23177,N_22923,N_22846);
nand U23178 (N_23178,N_22846,N_22814);
nor U23179 (N_23179,N_22971,N_22826);
nor U23180 (N_23180,N_22835,N_22929);
or U23181 (N_23181,N_22883,N_22945);
or U23182 (N_23182,N_22847,N_22880);
and U23183 (N_23183,N_22951,N_22880);
and U23184 (N_23184,N_22921,N_22881);
nor U23185 (N_23185,N_22994,N_22800);
nor U23186 (N_23186,N_22908,N_22906);
xor U23187 (N_23187,N_22947,N_22953);
and U23188 (N_23188,N_22881,N_22887);
xor U23189 (N_23189,N_22800,N_22816);
xor U23190 (N_23190,N_22809,N_22990);
nor U23191 (N_23191,N_22950,N_22875);
nand U23192 (N_23192,N_22967,N_22924);
nand U23193 (N_23193,N_22856,N_22980);
xnor U23194 (N_23194,N_22903,N_22936);
nor U23195 (N_23195,N_22938,N_22845);
nor U23196 (N_23196,N_22873,N_22926);
xnor U23197 (N_23197,N_22820,N_22866);
nand U23198 (N_23198,N_22839,N_22919);
or U23199 (N_23199,N_22811,N_22983);
nand U23200 (N_23200,N_23018,N_23120);
nand U23201 (N_23201,N_23077,N_23092);
nor U23202 (N_23202,N_23000,N_23103);
xor U23203 (N_23203,N_23171,N_23027);
nand U23204 (N_23204,N_23163,N_23186);
and U23205 (N_23205,N_23106,N_23001);
nand U23206 (N_23206,N_23139,N_23020);
or U23207 (N_23207,N_23048,N_23060);
or U23208 (N_23208,N_23069,N_23035);
nand U23209 (N_23209,N_23182,N_23012);
xor U23210 (N_23210,N_23006,N_23108);
xnor U23211 (N_23211,N_23191,N_23063);
and U23212 (N_23212,N_23109,N_23101);
nand U23213 (N_23213,N_23011,N_23136);
xor U23214 (N_23214,N_23043,N_23189);
or U23215 (N_23215,N_23087,N_23031);
or U23216 (N_23216,N_23039,N_23073);
nand U23217 (N_23217,N_23061,N_23085);
or U23218 (N_23218,N_23026,N_23115);
nor U23219 (N_23219,N_23152,N_23003);
and U23220 (N_23220,N_23030,N_23117);
nand U23221 (N_23221,N_23095,N_23162);
nor U23222 (N_23222,N_23150,N_23118);
nor U23223 (N_23223,N_23021,N_23160);
or U23224 (N_23224,N_23185,N_23125);
nand U23225 (N_23225,N_23126,N_23164);
nand U23226 (N_23226,N_23054,N_23140);
xor U23227 (N_23227,N_23167,N_23016);
and U23228 (N_23228,N_23196,N_23119);
nand U23229 (N_23229,N_23166,N_23046);
and U23230 (N_23230,N_23015,N_23157);
and U23231 (N_23231,N_23057,N_23188);
nand U23232 (N_23232,N_23190,N_23199);
or U23233 (N_23233,N_23124,N_23195);
nand U23234 (N_23234,N_23019,N_23037);
or U23235 (N_23235,N_23170,N_23128);
or U23236 (N_23236,N_23013,N_23083);
and U23237 (N_23237,N_23187,N_23148);
and U23238 (N_23238,N_23032,N_23181);
nor U23239 (N_23239,N_23146,N_23153);
and U23240 (N_23240,N_23070,N_23014);
or U23241 (N_23241,N_23110,N_23168);
nor U23242 (N_23242,N_23068,N_23071);
and U23243 (N_23243,N_23034,N_23096);
and U23244 (N_23244,N_23050,N_23076);
and U23245 (N_23245,N_23133,N_23138);
nor U23246 (N_23246,N_23149,N_23010);
nand U23247 (N_23247,N_23135,N_23184);
and U23248 (N_23248,N_23122,N_23194);
nand U23249 (N_23249,N_23052,N_23192);
or U23250 (N_23250,N_23044,N_23066);
nor U23251 (N_23251,N_23082,N_23112);
xnor U23252 (N_23252,N_23180,N_23081);
nor U23253 (N_23253,N_23004,N_23065);
nand U23254 (N_23254,N_23058,N_23002);
and U23255 (N_23255,N_23141,N_23121);
xor U23256 (N_23256,N_23056,N_23169);
or U23257 (N_23257,N_23098,N_23172);
nor U23258 (N_23258,N_23130,N_23059);
nand U23259 (N_23259,N_23102,N_23104);
or U23260 (N_23260,N_23155,N_23045);
or U23261 (N_23261,N_23089,N_23075);
xor U23262 (N_23262,N_23023,N_23005);
nand U23263 (N_23263,N_23029,N_23161);
nor U23264 (N_23264,N_23142,N_23165);
or U23265 (N_23265,N_23129,N_23183);
and U23266 (N_23266,N_23041,N_23036);
nor U23267 (N_23267,N_23074,N_23147);
and U23268 (N_23268,N_23053,N_23088);
nand U23269 (N_23269,N_23024,N_23113);
nand U23270 (N_23270,N_23198,N_23025);
nor U23271 (N_23271,N_23079,N_23067);
xnor U23272 (N_23272,N_23144,N_23008);
xor U23273 (N_23273,N_23105,N_23062);
and U23274 (N_23274,N_23116,N_23028);
nand U23275 (N_23275,N_23137,N_23064);
nand U23276 (N_23276,N_23111,N_23114);
xnor U23277 (N_23277,N_23132,N_23078);
xor U23278 (N_23278,N_23022,N_23134);
or U23279 (N_23279,N_23055,N_23091);
nor U23280 (N_23280,N_23197,N_23178);
or U23281 (N_23281,N_23193,N_23097);
nand U23282 (N_23282,N_23143,N_23094);
and U23283 (N_23283,N_23123,N_23093);
nand U23284 (N_23284,N_23090,N_23145);
xnor U23285 (N_23285,N_23176,N_23033);
or U23286 (N_23286,N_23159,N_23179);
or U23287 (N_23287,N_23099,N_23017);
or U23288 (N_23288,N_23051,N_23038);
or U23289 (N_23289,N_23154,N_23084);
and U23290 (N_23290,N_23174,N_23177);
nand U23291 (N_23291,N_23107,N_23175);
and U23292 (N_23292,N_23173,N_23156);
xnor U23293 (N_23293,N_23072,N_23040);
nand U23294 (N_23294,N_23127,N_23007);
xor U23295 (N_23295,N_23158,N_23086);
and U23296 (N_23296,N_23131,N_23049);
xor U23297 (N_23297,N_23100,N_23042);
nand U23298 (N_23298,N_23009,N_23047);
xor U23299 (N_23299,N_23151,N_23080);
or U23300 (N_23300,N_23022,N_23109);
or U23301 (N_23301,N_23023,N_23028);
or U23302 (N_23302,N_23075,N_23065);
xnor U23303 (N_23303,N_23078,N_23107);
xor U23304 (N_23304,N_23173,N_23123);
or U23305 (N_23305,N_23033,N_23106);
or U23306 (N_23306,N_23111,N_23120);
xor U23307 (N_23307,N_23185,N_23135);
or U23308 (N_23308,N_23151,N_23128);
or U23309 (N_23309,N_23133,N_23062);
or U23310 (N_23310,N_23067,N_23016);
nand U23311 (N_23311,N_23100,N_23103);
nor U23312 (N_23312,N_23034,N_23160);
nand U23313 (N_23313,N_23084,N_23011);
nor U23314 (N_23314,N_23025,N_23157);
nand U23315 (N_23315,N_23053,N_23180);
or U23316 (N_23316,N_23186,N_23168);
and U23317 (N_23317,N_23122,N_23036);
xor U23318 (N_23318,N_23037,N_23159);
nand U23319 (N_23319,N_23019,N_23057);
xnor U23320 (N_23320,N_23155,N_23015);
nand U23321 (N_23321,N_23097,N_23017);
xor U23322 (N_23322,N_23129,N_23015);
nand U23323 (N_23323,N_23128,N_23141);
xor U23324 (N_23324,N_23099,N_23038);
and U23325 (N_23325,N_23115,N_23000);
xnor U23326 (N_23326,N_23057,N_23003);
nor U23327 (N_23327,N_23188,N_23103);
xor U23328 (N_23328,N_23065,N_23143);
or U23329 (N_23329,N_23127,N_23032);
nand U23330 (N_23330,N_23170,N_23132);
xnor U23331 (N_23331,N_23067,N_23162);
nand U23332 (N_23332,N_23136,N_23115);
xnor U23333 (N_23333,N_23174,N_23028);
and U23334 (N_23334,N_23064,N_23126);
or U23335 (N_23335,N_23025,N_23064);
xnor U23336 (N_23336,N_23137,N_23052);
and U23337 (N_23337,N_23153,N_23035);
nand U23338 (N_23338,N_23024,N_23046);
or U23339 (N_23339,N_23055,N_23099);
nand U23340 (N_23340,N_23197,N_23062);
xnor U23341 (N_23341,N_23098,N_23025);
xnor U23342 (N_23342,N_23173,N_23074);
xnor U23343 (N_23343,N_23187,N_23170);
nor U23344 (N_23344,N_23146,N_23164);
or U23345 (N_23345,N_23000,N_23065);
nor U23346 (N_23346,N_23182,N_23109);
nor U23347 (N_23347,N_23060,N_23035);
or U23348 (N_23348,N_23111,N_23189);
nor U23349 (N_23349,N_23078,N_23085);
nor U23350 (N_23350,N_23037,N_23113);
or U23351 (N_23351,N_23094,N_23018);
nand U23352 (N_23352,N_23072,N_23113);
or U23353 (N_23353,N_23003,N_23182);
xor U23354 (N_23354,N_23147,N_23093);
nand U23355 (N_23355,N_23063,N_23130);
nor U23356 (N_23356,N_23042,N_23150);
nor U23357 (N_23357,N_23000,N_23003);
and U23358 (N_23358,N_23076,N_23187);
nand U23359 (N_23359,N_23163,N_23054);
nand U23360 (N_23360,N_23196,N_23107);
or U23361 (N_23361,N_23125,N_23021);
nand U23362 (N_23362,N_23090,N_23093);
nor U23363 (N_23363,N_23154,N_23114);
nor U23364 (N_23364,N_23139,N_23180);
xor U23365 (N_23365,N_23186,N_23142);
nor U23366 (N_23366,N_23147,N_23013);
xnor U23367 (N_23367,N_23122,N_23038);
or U23368 (N_23368,N_23005,N_23178);
and U23369 (N_23369,N_23095,N_23186);
nand U23370 (N_23370,N_23022,N_23013);
and U23371 (N_23371,N_23181,N_23199);
or U23372 (N_23372,N_23171,N_23150);
nor U23373 (N_23373,N_23180,N_23019);
or U23374 (N_23374,N_23036,N_23014);
nor U23375 (N_23375,N_23114,N_23155);
and U23376 (N_23376,N_23115,N_23176);
nand U23377 (N_23377,N_23086,N_23168);
or U23378 (N_23378,N_23109,N_23157);
nand U23379 (N_23379,N_23021,N_23171);
nor U23380 (N_23380,N_23073,N_23067);
xnor U23381 (N_23381,N_23134,N_23004);
nor U23382 (N_23382,N_23102,N_23190);
nand U23383 (N_23383,N_23071,N_23124);
and U23384 (N_23384,N_23183,N_23164);
or U23385 (N_23385,N_23124,N_23012);
and U23386 (N_23386,N_23148,N_23191);
and U23387 (N_23387,N_23160,N_23004);
nor U23388 (N_23388,N_23136,N_23190);
nand U23389 (N_23389,N_23084,N_23132);
and U23390 (N_23390,N_23029,N_23105);
and U23391 (N_23391,N_23147,N_23063);
xnor U23392 (N_23392,N_23061,N_23087);
or U23393 (N_23393,N_23020,N_23036);
nand U23394 (N_23394,N_23145,N_23160);
nand U23395 (N_23395,N_23068,N_23166);
nor U23396 (N_23396,N_23057,N_23182);
nor U23397 (N_23397,N_23124,N_23064);
and U23398 (N_23398,N_23112,N_23110);
xor U23399 (N_23399,N_23083,N_23122);
or U23400 (N_23400,N_23311,N_23250);
or U23401 (N_23401,N_23276,N_23277);
or U23402 (N_23402,N_23290,N_23270);
and U23403 (N_23403,N_23285,N_23354);
xor U23404 (N_23404,N_23317,N_23300);
or U23405 (N_23405,N_23264,N_23242);
nand U23406 (N_23406,N_23353,N_23230);
nand U23407 (N_23407,N_23275,N_23372);
and U23408 (N_23408,N_23296,N_23220);
and U23409 (N_23409,N_23320,N_23328);
and U23410 (N_23410,N_23281,N_23324);
nand U23411 (N_23411,N_23278,N_23340);
nor U23412 (N_23412,N_23216,N_23326);
nor U23413 (N_23413,N_23229,N_23329);
and U23414 (N_23414,N_23393,N_23225);
or U23415 (N_23415,N_23343,N_23249);
nand U23416 (N_23416,N_23294,N_23298);
xor U23417 (N_23417,N_23215,N_23210);
or U23418 (N_23418,N_23291,N_23271);
or U23419 (N_23419,N_23364,N_23337);
or U23420 (N_23420,N_23263,N_23268);
nand U23421 (N_23421,N_23332,N_23387);
nand U23422 (N_23422,N_23279,N_23307);
nor U23423 (N_23423,N_23301,N_23391);
and U23424 (N_23424,N_23389,N_23348);
nand U23425 (N_23425,N_23233,N_23396);
and U23426 (N_23426,N_23303,N_23321);
or U23427 (N_23427,N_23357,N_23207);
xor U23428 (N_23428,N_23375,N_23382);
and U23429 (N_23429,N_23247,N_23273);
and U23430 (N_23430,N_23392,N_23206);
xnor U23431 (N_23431,N_23287,N_23218);
and U23432 (N_23432,N_23256,N_23333);
and U23433 (N_23433,N_23217,N_23361);
and U23434 (N_23434,N_23293,N_23269);
xnor U23435 (N_23435,N_23310,N_23390);
nand U23436 (N_23436,N_23238,N_23200);
nand U23437 (N_23437,N_23376,N_23367);
nor U23438 (N_23438,N_23334,N_23399);
nor U23439 (N_23439,N_23385,N_23380);
and U23440 (N_23440,N_23374,N_23235);
and U23441 (N_23441,N_23258,N_23252);
nand U23442 (N_23442,N_23331,N_23342);
nor U23443 (N_23443,N_23386,N_23255);
and U23444 (N_23444,N_23347,N_23222);
and U23445 (N_23445,N_23368,N_23373);
and U23446 (N_23446,N_23202,N_23356);
xor U23447 (N_23447,N_23221,N_23330);
xnor U23448 (N_23448,N_23350,N_23336);
nor U23449 (N_23449,N_23322,N_23286);
nor U23450 (N_23450,N_23234,N_23318);
and U23451 (N_23451,N_23371,N_23227);
nand U23452 (N_23452,N_23344,N_23240);
and U23453 (N_23453,N_23395,N_23208);
nand U23454 (N_23454,N_23369,N_23223);
xor U23455 (N_23455,N_23272,N_23341);
or U23456 (N_23456,N_23304,N_23288);
and U23457 (N_23457,N_23282,N_23248);
nand U23458 (N_23458,N_23209,N_23246);
or U23459 (N_23459,N_23299,N_23305);
nand U23460 (N_23460,N_23316,N_23383);
or U23461 (N_23461,N_23267,N_23280);
xor U23462 (N_23462,N_23253,N_23335);
and U23463 (N_23463,N_23284,N_23366);
nand U23464 (N_23464,N_23323,N_23319);
nand U23465 (N_23465,N_23346,N_23379);
or U23466 (N_23466,N_23384,N_23398);
xor U23467 (N_23467,N_23297,N_23214);
and U23468 (N_23468,N_23397,N_23338);
or U23469 (N_23469,N_23325,N_23388);
xnor U23470 (N_23470,N_23360,N_23212);
and U23471 (N_23471,N_23259,N_23274);
xnor U23472 (N_23472,N_23351,N_23262);
nand U23473 (N_23473,N_23370,N_23314);
nor U23474 (N_23474,N_23245,N_23295);
nand U23475 (N_23475,N_23306,N_23358);
or U23476 (N_23476,N_23309,N_23257);
and U23477 (N_23477,N_23219,N_23243);
nand U23478 (N_23478,N_23352,N_23224);
nor U23479 (N_23479,N_23363,N_23239);
and U23480 (N_23480,N_23237,N_23394);
or U23481 (N_23481,N_23378,N_23339);
nor U23482 (N_23482,N_23231,N_23362);
nor U23483 (N_23483,N_23241,N_23289);
or U23484 (N_23484,N_23315,N_23292);
nand U23485 (N_23485,N_23211,N_23236);
or U23486 (N_23486,N_23359,N_23302);
nand U23487 (N_23487,N_23313,N_23228);
nor U23488 (N_23488,N_23377,N_23355);
or U23489 (N_23489,N_23205,N_23312);
xor U23490 (N_23490,N_23232,N_23365);
nand U23491 (N_23491,N_23213,N_23203);
and U23492 (N_23492,N_23261,N_23283);
nor U23493 (N_23493,N_23349,N_23260);
nor U23494 (N_23494,N_23251,N_23381);
or U23495 (N_23495,N_23204,N_23226);
or U23496 (N_23496,N_23254,N_23327);
and U23497 (N_23497,N_23244,N_23265);
nand U23498 (N_23498,N_23201,N_23308);
and U23499 (N_23499,N_23345,N_23266);
and U23500 (N_23500,N_23287,N_23338);
nor U23501 (N_23501,N_23340,N_23224);
and U23502 (N_23502,N_23200,N_23252);
nand U23503 (N_23503,N_23301,N_23341);
nor U23504 (N_23504,N_23248,N_23216);
and U23505 (N_23505,N_23206,N_23321);
nor U23506 (N_23506,N_23372,N_23200);
nand U23507 (N_23507,N_23355,N_23279);
and U23508 (N_23508,N_23204,N_23239);
and U23509 (N_23509,N_23331,N_23284);
nand U23510 (N_23510,N_23341,N_23269);
nand U23511 (N_23511,N_23218,N_23267);
nor U23512 (N_23512,N_23368,N_23398);
xor U23513 (N_23513,N_23295,N_23324);
nor U23514 (N_23514,N_23249,N_23232);
or U23515 (N_23515,N_23330,N_23274);
xor U23516 (N_23516,N_23321,N_23385);
nor U23517 (N_23517,N_23320,N_23225);
nand U23518 (N_23518,N_23325,N_23373);
and U23519 (N_23519,N_23353,N_23291);
nor U23520 (N_23520,N_23368,N_23335);
nor U23521 (N_23521,N_23334,N_23295);
or U23522 (N_23522,N_23300,N_23333);
and U23523 (N_23523,N_23206,N_23214);
nand U23524 (N_23524,N_23315,N_23366);
or U23525 (N_23525,N_23219,N_23275);
xnor U23526 (N_23526,N_23224,N_23251);
nor U23527 (N_23527,N_23384,N_23290);
and U23528 (N_23528,N_23237,N_23305);
nor U23529 (N_23529,N_23390,N_23277);
and U23530 (N_23530,N_23297,N_23354);
xor U23531 (N_23531,N_23235,N_23349);
nor U23532 (N_23532,N_23333,N_23315);
nor U23533 (N_23533,N_23363,N_23202);
xor U23534 (N_23534,N_23233,N_23322);
or U23535 (N_23535,N_23361,N_23303);
nor U23536 (N_23536,N_23299,N_23233);
or U23537 (N_23537,N_23301,N_23239);
and U23538 (N_23538,N_23376,N_23316);
and U23539 (N_23539,N_23242,N_23335);
or U23540 (N_23540,N_23205,N_23252);
and U23541 (N_23541,N_23336,N_23239);
and U23542 (N_23542,N_23368,N_23341);
and U23543 (N_23543,N_23247,N_23300);
nand U23544 (N_23544,N_23253,N_23300);
nor U23545 (N_23545,N_23351,N_23334);
nor U23546 (N_23546,N_23326,N_23275);
nand U23547 (N_23547,N_23299,N_23229);
nand U23548 (N_23548,N_23286,N_23305);
nand U23549 (N_23549,N_23236,N_23227);
or U23550 (N_23550,N_23201,N_23323);
and U23551 (N_23551,N_23342,N_23289);
or U23552 (N_23552,N_23286,N_23268);
or U23553 (N_23553,N_23255,N_23396);
xnor U23554 (N_23554,N_23255,N_23220);
or U23555 (N_23555,N_23296,N_23289);
nor U23556 (N_23556,N_23254,N_23237);
xnor U23557 (N_23557,N_23310,N_23253);
nand U23558 (N_23558,N_23287,N_23263);
nor U23559 (N_23559,N_23386,N_23348);
xor U23560 (N_23560,N_23321,N_23380);
nand U23561 (N_23561,N_23296,N_23256);
nor U23562 (N_23562,N_23298,N_23209);
or U23563 (N_23563,N_23200,N_23210);
nand U23564 (N_23564,N_23248,N_23287);
and U23565 (N_23565,N_23309,N_23292);
nor U23566 (N_23566,N_23396,N_23343);
xor U23567 (N_23567,N_23388,N_23334);
xnor U23568 (N_23568,N_23340,N_23386);
nand U23569 (N_23569,N_23281,N_23345);
or U23570 (N_23570,N_23341,N_23256);
nor U23571 (N_23571,N_23306,N_23325);
or U23572 (N_23572,N_23308,N_23342);
nand U23573 (N_23573,N_23376,N_23212);
nor U23574 (N_23574,N_23229,N_23312);
and U23575 (N_23575,N_23380,N_23206);
and U23576 (N_23576,N_23293,N_23238);
xnor U23577 (N_23577,N_23216,N_23332);
and U23578 (N_23578,N_23370,N_23337);
nor U23579 (N_23579,N_23219,N_23338);
nand U23580 (N_23580,N_23319,N_23344);
nor U23581 (N_23581,N_23325,N_23300);
nor U23582 (N_23582,N_23236,N_23298);
and U23583 (N_23583,N_23338,N_23326);
nor U23584 (N_23584,N_23260,N_23332);
or U23585 (N_23585,N_23298,N_23265);
nor U23586 (N_23586,N_23281,N_23394);
and U23587 (N_23587,N_23218,N_23347);
and U23588 (N_23588,N_23321,N_23327);
or U23589 (N_23589,N_23343,N_23233);
and U23590 (N_23590,N_23343,N_23393);
nand U23591 (N_23591,N_23390,N_23228);
and U23592 (N_23592,N_23262,N_23360);
xor U23593 (N_23593,N_23291,N_23312);
nor U23594 (N_23594,N_23394,N_23348);
nor U23595 (N_23595,N_23356,N_23285);
xor U23596 (N_23596,N_23223,N_23346);
xor U23597 (N_23597,N_23313,N_23352);
nor U23598 (N_23598,N_23271,N_23305);
nor U23599 (N_23599,N_23253,N_23297);
xor U23600 (N_23600,N_23567,N_23448);
or U23601 (N_23601,N_23407,N_23503);
and U23602 (N_23602,N_23408,N_23401);
xnor U23603 (N_23603,N_23526,N_23461);
nor U23604 (N_23604,N_23539,N_23501);
nor U23605 (N_23605,N_23598,N_23558);
nand U23606 (N_23606,N_23561,N_23458);
or U23607 (N_23607,N_23568,N_23548);
nor U23608 (N_23608,N_23569,N_23484);
nor U23609 (N_23609,N_23563,N_23438);
xor U23610 (N_23610,N_23523,N_23404);
nor U23611 (N_23611,N_23544,N_23590);
and U23612 (N_23612,N_23459,N_23466);
nor U23613 (N_23613,N_23442,N_23417);
nor U23614 (N_23614,N_23493,N_23443);
or U23615 (N_23615,N_23535,N_23499);
xnor U23616 (N_23616,N_23410,N_23480);
xor U23617 (N_23617,N_23582,N_23490);
nand U23618 (N_23618,N_23586,N_23498);
and U23619 (N_23619,N_23464,N_23572);
xor U23620 (N_23620,N_23476,N_23456);
nor U23621 (N_23621,N_23428,N_23536);
or U23622 (N_23622,N_23471,N_23431);
xnor U23623 (N_23623,N_23412,N_23440);
nor U23624 (N_23624,N_23541,N_23505);
and U23625 (N_23625,N_23515,N_23468);
nand U23626 (N_23626,N_23425,N_23477);
and U23627 (N_23627,N_23423,N_23432);
or U23628 (N_23628,N_23421,N_23529);
xor U23629 (N_23629,N_23446,N_23422);
or U23630 (N_23630,N_23518,N_23414);
nor U23631 (N_23631,N_23427,N_23577);
xor U23632 (N_23632,N_23587,N_23588);
xor U23633 (N_23633,N_23565,N_23506);
and U23634 (N_23634,N_23524,N_23411);
nor U23635 (N_23635,N_23416,N_23514);
xnor U23636 (N_23636,N_23538,N_23495);
or U23637 (N_23637,N_23489,N_23452);
or U23638 (N_23638,N_23540,N_23556);
nand U23639 (N_23639,N_23553,N_23487);
xor U23640 (N_23640,N_23437,N_23547);
nor U23641 (N_23641,N_23400,N_23474);
nor U23642 (N_23642,N_23450,N_23574);
xor U23643 (N_23643,N_23444,N_23496);
or U23644 (N_23644,N_23581,N_23597);
nor U23645 (N_23645,N_23434,N_23566);
and U23646 (N_23646,N_23419,N_23549);
xor U23647 (N_23647,N_23492,N_23485);
and U23648 (N_23648,N_23509,N_23534);
and U23649 (N_23649,N_23579,N_23592);
nor U23650 (N_23650,N_23402,N_23543);
xor U23651 (N_23651,N_23578,N_23550);
xnor U23652 (N_23652,N_23455,N_23596);
nor U23653 (N_23653,N_23557,N_23551);
nand U23654 (N_23654,N_23595,N_23439);
xnor U23655 (N_23655,N_23469,N_23454);
nand U23656 (N_23656,N_23522,N_23441);
and U23657 (N_23657,N_23511,N_23502);
nor U23658 (N_23658,N_23560,N_23580);
nor U23659 (N_23659,N_23465,N_23537);
nor U23660 (N_23660,N_23429,N_23517);
nor U23661 (N_23661,N_23531,N_23500);
nor U23662 (N_23662,N_23486,N_23418);
xnor U23663 (N_23663,N_23463,N_23467);
and U23664 (N_23664,N_23591,N_23433);
nor U23665 (N_23665,N_23430,N_23409);
and U23666 (N_23666,N_23533,N_23478);
or U23667 (N_23667,N_23599,N_23472);
xor U23668 (N_23668,N_23513,N_23483);
nand U23669 (N_23669,N_23473,N_23542);
nand U23670 (N_23670,N_23497,N_23426);
xnor U23671 (N_23671,N_23462,N_23584);
xnor U23672 (N_23672,N_23564,N_23449);
nor U23673 (N_23673,N_23510,N_23573);
and U23674 (N_23674,N_23447,N_23460);
xor U23675 (N_23675,N_23575,N_23532);
or U23676 (N_23676,N_23494,N_23576);
and U23677 (N_23677,N_23520,N_23554);
or U23678 (N_23678,N_23451,N_23521);
xor U23679 (N_23679,N_23415,N_23508);
nand U23680 (N_23680,N_23527,N_23552);
and U23681 (N_23681,N_23530,N_23583);
nor U23682 (N_23682,N_23406,N_23589);
and U23683 (N_23683,N_23593,N_23570);
and U23684 (N_23684,N_23420,N_23413);
nand U23685 (N_23685,N_23424,N_23482);
or U23686 (N_23686,N_23559,N_23594);
xor U23687 (N_23687,N_23528,N_23445);
nand U23688 (N_23688,N_23488,N_23546);
xnor U23689 (N_23689,N_23491,N_23512);
nor U23690 (N_23690,N_23453,N_23545);
xnor U23691 (N_23691,N_23516,N_23519);
or U23692 (N_23692,N_23507,N_23457);
and U23693 (N_23693,N_23481,N_23435);
nand U23694 (N_23694,N_23585,N_23525);
nand U23695 (N_23695,N_23403,N_23504);
xor U23696 (N_23696,N_23405,N_23562);
and U23697 (N_23697,N_23479,N_23436);
or U23698 (N_23698,N_23475,N_23555);
and U23699 (N_23699,N_23571,N_23470);
nand U23700 (N_23700,N_23494,N_23593);
xnor U23701 (N_23701,N_23465,N_23543);
nor U23702 (N_23702,N_23450,N_23457);
nand U23703 (N_23703,N_23572,N_23548);
xor U23704 (N_23704,N_23563,N_23546);
xor U23705 (N_23705,N_23468,N_23405);
nor U23706 (N_23706,N_23589,N_23510);
xnor U23707 (N_23707,N_23594,N_23405);
and U23708 (N_23708,N_23511,N_23500);
or U23709 (N_23709,N_23448,N_23498);
or U23710 (N_23710,N_23503,N_23544);
nor U23711 (N_23711,N_23430,N_23526);
xor U23712 (N_23712,N_23462,N_23463);
or U23713 (N_23713,N_23581,N_23567);
or U23714 (N_23714,N_23587,N_23445);
or U23715 (N_23715,N_23527,N_23595);
xor U23716 (N_23716,N_23432,N_23403);
and U23717 (N_23717,N_23532,N_23410);
xnor U23718 (N_23718,N_23535,N_23563);
nand U23719 (N_23719,N_23593,N_23574);
or U23720 (N_23720,N_23570,N_23471);
or U23721 (N_23721,N_23475,N_23561);
nand U23722 (N_23722,N_23579,N_23595);
nand U23723 (N_23723,N_23448,N_23444);
nor U23724 (N_23724,N_23435,N_23431);
and U23725 (N_23725,N_23445,N_23531);
nor U23726 (N_23726,N_23487,N_23598);
and U23727 (N_23727,N_23500,N_23430);
xnor U23728 (N_23728,N_23584,N_23516);
nor U23729 (N_23729,N_23490,N_23577);
or U23730 (N_23730,N_23435,N_23430);
xor U23731 (N_23731,N_23452,N_23402);
nor U23732 (N_23732,N_23575,N_23404);
or U23733 (N_23733,N_23502,N_23536);
nor U23734 (N_23734,N_23546,N_23445);
or U23735 (N_23735,N_23487,N_23509);
nand U23736 (N_23736,N_23555,N_23551);
nor U23737 (N_23737,N_23593,N_23439);
or U23738 (N_23738,N_23557,N_23468);
nand U23739 (N_23739,N_23438,N_23510);
and U23740 (N_23740,N_23542,N_23404);
nor U23741 (N_23741,N_23454,N_23500);
xor U23742 (N_23742,N_23470,N_23550);
or U23743 (N_23743,N_23470,N_23516);
xor U23744 (N_23744,N_23420,N_23580);
and U23745 (N_23745,N_23485,N_23576);
or U23746 (N_23746,N_23511,N_23521);
xnor U23747 (N_23747,N_23576,N_23442);
nand U23748 (N_23748,N_23494,N_23566);
and U23749 (N_23749,N_23521,N_23534);
nand U23750 (N_23750,N_23587,N_23427);
nand U23751 (N_23751,N_23427,N_23422);
and U23752 (N_23752,N_23423,N_23473);
nor U23753 (N_23753,N_23518,N_23420);
nand U23754 (N_23754,N_23473,N_23493);
xnor U23755 (N_23755,N_23456,N_23495);
nand U23756 (N_23756,N_23513,N_23440);
nor U23757 (N_23757,N_23578,N_23523);
and U23758 (N_23758,N_23543,N_23476);
and U23759 (N_23759,N_23569,N_23560);
xnor U23760 (N_23760,N_23421,N_23507);
xor U23761 (N_23761,N_23592,N_23511);
xnor U23762 (N_23762,N_23526,N_23487);
nor U23763 (N_23763,N_23478,N_23495);
or U23764 (N_23764,N_23589,N_23579);
xnor U23765 (N_23765,N_23539,N_23450);
nand U23766 (N_23766,N_23497,N_23566);
and U23767 (N_23767,N_23446,N_23463);
xor U23768 (N_23768,N_23569,N_23582);
and U23769 (N_23769,N_23442,N_23555);
xnor U23770 (N_23770,N_23560,N_23525);
or U23771 (N_23771,N_23597,N_23448);
or U23772 (N_23772,N_23488,N_23460);
nor U23773 (N_23773,N_23589,N_23461);
and U23774 (N_23774,N_23545,N_23477);
and U23775 (N_23775,N_23579,N_23526);
or U23776 (N_23776,N_23472,N_23576);
and U23777 (N_23777,N_23495,N_23490);
and U23778 (N_23778,N_23548,N_23563);
nor U23779 (N_23779,N_23557,N_23519);
and U23780 (N_23780,N_23564,N_23583);
nor U23781 (N_23781,N_23545,N_23560);
xor U23782 (N_23782,N_23546,N_23441);
nand U23783 (N_23783,N_23465,N_23423);
xor U23784 (N_23784,N_23418,N_23516);
and U23785 (N_23785,N_23473,N_23540);
xnor U23786 (N_23786,N_23458,N_23492);
xnor U23787 (N_23787,N_23441,N_23555);
and U23788 (N_23788,N_23575,N_23504);
nand U23789 (N_23789,N_23412,N_23578);
or U23790 (N_23790,N_23490,N_23588);
nor U23791 (N_23791,N_23501,N_23569);
nand U23792 (N_23792,N_23476,N_23523);
nor U23793 (N_23793,N_23591,N_23469);
xnor U23794 (N_23794,N_23588,N_23425);
xor U23795 (N_23795,N_23446,N_23454);
or U23796 (N_23796,N_23434,N_23540);
or U23797 (N_23797,N_23492,N_23480);
xor U23798 (N_23798,N_23532,N_23590);
xor U23799 (N_23799,N_23552,N_23473);
nor U23800 (N_23800,N_23762,N_23668);
nand U23801 (N_23801,N_23639,N_23716);
nor U23802 (N_23802,N_23725,N_23726);
xor U23803 (N_23803,N_23663,N_23660);
xor U23804 (N_23804,N_23617,N_23623);
nand U23805 (N_23805,N_23645,N_23750);
or U23806 (N_23806,N_23677,N_23654);
nand U23807 (N_23807,N_23783,N_23734);
or U23808 (N_23808,N_23678,N_23642);
nor U23809 (N_23809,N_23683,N_23629);
xnor U23810 (N_23810,N_23755,N_23680);
or U23811 (N_23811,N_23761,N_23604);
or U23812 (N_23812,N_23703,N_23669);
xor U23813 (N_23813,N_23776,N_23619);
and U23814 (N_23814,N_23634,N_23730);
or U23815 (N_23815,N_23626,N_23717);
xnor U23816 (N_23816,N_23659,N_23690);
nand U23817 (N_23817,N_23739,N_23727);
nand U23818 (N_23818,N_23724,N_23618);
or U23819 (N_23819,N_23754,N_23666);
xor U23820 (N_23820,N_23606,N_23763);
or U23821 (N_23821,N_23700,N_23787);
and U23822 (N_23822,N_23785,N_23658);
xor U23823 (N_23823,N_23768,N_23741);
or U23824 (N_23824,N_23708,N_23740);
xor U23825 (N_23825,N_23705,N_23628);
nand U23826 (N_23826,N_23706,N_23735);
nand U23827 (N_23827,N_23751,N_23614);
nor U23828 (N_23828,N_23721,N_23601);
nor U23829 (N_23829,N_23622,N_23712);
nor U23830 (N_23830,N_23672,N_23746);
xor U23831 (N_23831,N_23607,N_23674);
xor U23832 (N_23832,N_23701,N_23760);
nand U23833 (N_23833,N_23702,N_23793);
and U23834 (N_23834,N_23777,N_23686);
xnor U23835 (N_23835,N_23764,N_23685);
or U23836 (N_23836,N_23778,N_23613);
and U23837 (N_23837,N_23633,N_23692);
nor U23838 (N_23838,N_23781,N_23632);
nand U23839 (N_23839,N_23693,N_23627);
xnor U23840 (N_23840,N_23722,N_23641);
or U23841 (N_23841,N_23711,N_23616);
or U23842 (N_23842,N_23676,N_23694);
nor U23843 (N_23843,N_23745,N_23753);
and U23844 (N_23844,N_23647,N_23644);
xnor U23845 (N_23845,N_23649,N_23707);
nand U23846 (N_23846,N_23718,N_23759);
xor U23847 (N_23847,N_23738,N_23782);
and U23848 (N_23848,N_23682,N_23748);
nor U23849 (N_23849,N_23752,N_23772);
or U23850 (N_23850,N_23684,N_23615);
or U23851 (N_23851,N_23791,N_23637);
or U23852 (N_23852,N_23709,N_23729);
nand U23853 (N_23853,N_23765,N_23671);
nor U23854 (N_23854,N_23661,N_23769);
xor U23855 (N_23855,N_23698,N_23681);
nand U23856 (N_23856,N_23797,N_23773);
or U23857 (N_23857,N_23667,N_23696);
xnor U23858 (N_23858,N_23675,N_23638);
nand U23859 (N_23859,N_23795,N_23670);
and U23860 (N_23860,N_23687,N_23742);
xnor U23861 (N_23861,N_23640,N_23788);
or U23862 (N_23862,N_23611,N_23631);
and U23863 (N_23863,N_23603,N_23710);
xnor U23864 (N_23864,N_23749,N_23662);
nor U23865 (N_23865,N_23664,N_23704);
nor U23866 (N_23866,N_23636,N_23652);
nor U23867 (N_23867,N_23605,N_23697);
nor U23868 (N_23868,N_23699,N_23635);
nand U23869 (N_23869,N_23655,N_23743);
and U23870 (N_23870,N_23796,N_23691);
nand U23871 (N_23871,N_23630,N_23602);
xor U23872 (N_23872,N_23625,N_23798);
or U23873 (N_23873,N_23775,N_23780);
or U23874 (N_23874,N_23757,N_23715);
and U23875 (N_23875,N_23784,N_23731);
or U23876 (N_23876,N_23612,N_23767);
nand U23877 (N_23877,N_23774,N_23608);
nand U23878 (N_23878,N_23723,N_23728);
nand U23879 (N_23879,N_23789,N_23747);
nand U23880 (N_23880,N_23758,N_23610);
xnor U23881 (N_23881,N_23720,N_23688);
nand U23882 (N_23882,N_23719,N_23624);
or U23883 (N_23883,N_23799,N_23732);
and U23884 (N_23884,N_23679,N_23733);
and U23885 (N_23885,N_23779,N_23643);
nor U23886 (N_23886,N_23766,N_23600);
or U23887 (N_23887,N_23657,N_23790);
nand U23888 (N_23888,N_23656,N_23665);
and U23889 (N_23889,N_23744,N_23648);
and U23890 (N_23890,N_23713,N_23736);
xnor U23891 (N_23891,N_23621,N_23794);
and U23892 (N_23892,N_23653,N_23651);
or U23893 (N_23893,N_23714,N_23650);
and U23894 (N_23894,N_23792,N_23771);
or U23895 (N_23895,N_23673,N_23695);
nand U23896 (N_23896,N_23620,N_23609);
nor U23897 (N_23897,N_23646,N_23689);
xor U23898 (N_23898,N_23786,N_23737);
or U23899 (N_23899,N_23770,N_23756);
nor U23900 (N_23900,N_23631,N_23682);
xor U23901 (N_23901,N_23728,N_23652);
xor U23902 (N_23902,N_23692,N_23608);
nand U23903 (N_23903,N_23603,N_23605);
and U23904 (N_23904,N_23798,N_23772);
nor U23905 (N_23905,N_23635,N_23760);
and U23906 (N_23906,N_23655,N_23631);
and U23907 (N_23907,N_23766,N_23641);
xnor U23908 (N_23908,N_23636,N_23689);
and U23909 (N_23909,N_23698,N_23667);
and U23910 (N_23910,N_23617,N_23663);
or U23911 (N_23911,N_23615,N_23798);
and U23912 (N_23912,N_23683,N_23635);
xnor U23913 (N_23913,N_23670,N_23713);
nand U23914 (N_23914,N_23705,N_23789);
xnor U23915 (N_23915,N_23704,N_23604);
and U23916 (N_23916,N_23650,N_23736);
and U23917 (N_23917,N_23670,N_23730);
nor U23918 (N_23918,N_23771,N_23724);
xnor U23919 (N_23919,N_23686,N_23633);
nand U23920 (N_23920,N_23740,N_23702);
xor U23921 (N_23921,N_23689,N_23784);
nand U23922 (N_23922,N_23747,N_23655);
or U23923 (N_23923,N_23649,N_23735);
xor U23924 (N_23924,N_23625,N_23647);
xor U23925 (N_23925,N_23763,N_23766);
nand U23926 (N_23926,N_23766,N_23701);
xor U23927 (N_23927,N_23655,N_23763);
xnor U23928 (N_23928,N_23789,N_23655);
xor U23929 (N_23929,N_23723,N_23640);
and U23930 (N_23930,N_23740,N_23705);
and U23931 (N_23931,N_23641,N_23675);
and U23932 (N_23932,N_23647,N_23694);
or U23933 (N_23933,N_23647,N_23750);
xor U23934 (N_23934,N_23654,N_23779);
or U23935 (N_23935,N_23649,N_23605);
nor U23936 (N_23936,N_23655,N_23614);
nor U23937 (N_23937,N_23779,N_23682);
or U23938 (N_23938,N_23761,N_23792);
nor U23939 (N_23939,N_23643,N_23676);
xnor U23940 (N_23940,N_23767,N_23621);
or U23941 (N_23941,N_23789,N_23797);
or U23942 (N_23942,N_23789,N_23764);
nor U23943 (N_23943,N_23601,N_23723);
nor U23944 (N_23944,N_23734,N_23792);
xor U23945 (N_23945,N_23784,N_23715);
nor U23946 (N_23946,N_23600,N_23711);
or U23947 (N_23947,N_23674,N_23605);
or U23948 (N_23948,N_23791,N_23710);
xnor U23949 (N_23949,N_23738,N_23768);
or U23950 (N_23950,N_23705,N_23602);
nand U23951 (N_23951,N_23654,N_23649);
xor U23952 (N_23952,N_23641,N_23761);
and U23953 (N_23953,N_23669,N_23701);
nor U23954 (N_23954,N_23750,N_23786);
nand U23955 (N_23955,N_23791,N_23783);
or U23956 (N_23956,N_23725,N_23681);
nand U23957 (N_23957,N_23794,N_23727);
nand U23958 (N_23958,N_23667,N_23786);
or U23959 (N_23959,N_23652,N_23627);
or U23960 (N_23960,N_23642,N_23672);
or U23961 (N_23961,N_23761,N_23601);
nor U23962 (N_23962,N_23735,N_23624);
or U23963 (N_23963,N_23704,N_23776);
nand U23964 (N_23964,N_23600,N_23699);
xnor U23965 (N_23965,N_23784,N_23733);
or U23966 (N_23966,N_23630,N_23799);
nand U23967 (N_23967,N_23603,N_23741);
nand U23968 (N_23968,N_23691,N_23755);
and U23969 (N_23969,N_23799,N_23675);
nor U23970 (N_23970,N_23777,N_23642);
nand U23971 (N_23971,N_23642,N_23602);
xnor U23972 (N_23972,N_23673,N_23794);
xnor U23973 (N_23973,N_23743,N_23636);
nor U23974 (N_23974,N_23626,N_23691);
xnor U23975 (N_23975,N_23781,N_23751);
nor U23976 (N_23976,N_23703,N_23704);
or U23977 (N_23977,N_23756,N_23634);
xor U23978 (N_23978,N_23698,N_23661);
and U23979 (N_23979,N_23636,N_23774);
nand U23980 (N_23980,N_23788,N_23753);
nor U23981 (N_23981,N_23664,N_23784);
nand U23982 (N_23982,N_23632,N_23642);
nor U23983 (N_23983,N_23740,N_23621);
nor U23984 (N_23984,N_23717,N_23631);
nand U23985 (N_23985,N_23713,N_23747);
xor U23986 (N_23986,N_23606,N_23612);
nand U23987 (N_23987,N_23612,N_23615);
and U23988 (N_23988,N_23728,N_23749);
or U23989 (N_23989,N_23688,N_23777);
and U23990 (N_23990,N_23793,N_23780);
or U23991 (N_23991,N_23660,N_23729);
or U23992 (N_23992,N_23645,N_23774);
xnor U23993 (N_23993,N_23601,N_23637);
and U23994 (N_23994,N_23707,N_23701);
and U23995 (N_23995,N_23723,N_23631);
and U23996 (N_23996,N_23743,N_23789);
and U23997 (N_23997,N_23645,N_23714);
and U23998 (N_23998,N_23786,N_23611);
xor U23999 (N_23999,N_23634,N_23703);
xor U24000 (N_24000,N_23872,N_23966);
or U24001 (N_24001,N_23912,N_23864);
nand U24002 (N_24002,N_23819,N_23895);
nor U24003 (N_24003,N_23985,N_23935);
nand U24004 (N_24004,N_23978,N_23811);
nand U24005 (N_24005,N_23932,N_23994);
nor U24006 (N_24006,N_23829,N_23928);
nand U24007 (N_24007,N_23996,N_23860);
and U24008 (N_24008,N_23898,N_23970);
and U24009 (N_24009,N_23965,N_23804);
and U24010 (N_24010,N_23874,N_23969);
nor U24011 (N_24011,N_23984,N_23871);
xor U24012 (N_24012,N_23990,N_23840);
and U24013 (N_24013,N_23814,N_23803);
and U24014 (N_24014,N_23875,N_23919);
nor U24015 (N_24015,N_23841,N_23940);
nand U24016 (N_24016,N_23815,N_23962);
xor U24017 (N_24017,N_23824,N_23820);
xor U24018 (N_24018,N_23936,N_23809);
nand U24019 (N_24019,N_23857,N_23891);
or U24020 (N_24020,N_23849,N_23876);
xnor U24021 (N_24021,N_23910,N_23873);
and U24022 (N_24022,N_23926,N_23883);
nor U24023 (N_24023,N_23844,N_23980);
or U24024 (N_24024,N_23823,N_23929);
xnor U24025 (N_24025,N_23905,N_23881);
nand U24026 (N_24026,N_23953,N_23900);
xor U24027 (N_24027,N_23892,N_23894);
and U24028 (N_24028,N_23950,N_23976);
and U24029 (N_24029,N_23934,N_23918);
nor U24030 (N_24030,N_23938,N_23838);
nor U24031 (N_24031,N_23947,N_23948);
nor U24032 (N_24032,N_23833,N_23813);
or U24033 (N_24033,N_23957,N_23882);
nand U24034 (N_24034,N_23827,N_23831);
and U24035 (N_24035,N_23805,N_23999);
and U24036 (N_24036,N_23862,N_23997);
xor U24037 (N_24037,N_23973,N_23992);
nor U24038 (N_24038,N_23958,N_23974);
nor U24039 (N_24039,N_23982,N_23931);
nor U24040 (N_24040,N_23865,N_23971);
xnor U24041 (N_24041,N_23925,N_23802);
and U24042 (N_24042,N_23884,N_23933);
or U24043 (N_24043,N_23806,N_23975);
or U24044 (N_24044,N_23920,N_23816);
nand U24045 (N_24045,N_23964,N_23812);
xnor U24046 (N_24046,N_23904,N_23941);
xnor U24047 (N_24047,N_23836,N_23879);
and U24048 (N_24048,N_23922,N_23993);
or U24049 (N_24049,N_23908,N_23835);
or U24050 (N_24050,N_23951,N_23955);
and U24051 (N_24051,N_23810,N_23899);
and U24052 (N_24052,N_23944,N_23909);
and U24053 (N_24053,N_23808,N_23896);
nor U24054 (N_24054,N_23956,N_23847);
nand U24055 (N_24055,N_23855,N_23942);
nand U24056 (N_24056,N_23987,N_23991);
nor U24057 (N_24057,N_23889,N_23983);
or U24058 (N_24058,N_23972,N_23930);
xnor U24059 (N_24059,N_23924,N_23952);
and U24060 (N_24060,N_23821,N_23986);
or U24061 (N_24061,N_23807,N_23901);
and U24062 (N_24062,N_23852,N_23887);
and U24063 (N_24063,N_23927,N_23917);
xnor U24064 (N_24064,N_23822,N_23863);
and U24065 (N_24065,N_23897,N_23989);
nand U24066 (N_24066,N_23902,N_23800);
nor U24067 (N_24067,N_23945,N_23949);
xnor U24068 (N_24068,N_23921,N_23886);
nor U24069 (N_24069,N_23998,N_23877);
xor U24070 (N_24070,N_23868,N_23885);
nor U24071 (N_24071,N_23915,N_23867);
xor U24072 (N_24072,N_23937,N_23977);
and U24073 (N_24073,N_23893,N_23825);
and U24074 (N_24074,N_23853,N_23880);
nor U24075 (N_24075,N_23848,N_23858);
nor U24076 (N_24076,N_23846,N_23801);
xnor U24077 (N_24077,N_23850,N_23979);
nor U24078 (N_24078,N_23961,N_23817);
xor U24079 (N_24079,N_23842,N_23870);
nand U24080 (N_24080,N_23967,N_23914);
xor U24081 (N_24081,N_23830,N_23963);
and U24082 (N_24082,N_23968,N_23832);
and U24083 (N_24083,N_23854,N_23837);
or U24084 (N_24084,N_23981,N_23995);
xor U24085 (N_24085,N_23906,N_23828);
nor U24086 (N_24086,N_23845,N_23869);
nor U24087 (N_24087,N_23834,N_23923);
nand U24088 (N_24088,N_23913,N_23911);
or U24089 (N_24089,N_23959,N_23960);
and U24090 (N_24090,N_23826,N_23843);
or U24091 (N_24091,N_23939,N_23916);
or U24092 (N_24092,N_23859,N_23943);
nand U24093 (N_24093,N_23907,N_23851);
xor U24094 (N_24094,N_23866,N_23988);
and U24095 (N_24095,N_23839,N_23878);
xor U24096 (N_24096,N_23856,N_23903);
or U24097 (N_24097,N_23946,N_23890);
nand U24098 (N_24098,N_23861,N_23888);
or U24099 (N_24099,N_23818,N_23954);
nor U24100 (N_24100,N_23881,N_23827);
or U24101 (N_24101,N_23905,N_23970);
or U24102 (N_24102,N_23874,N_23903);
and U24103 (N_24103,N_23842,N_23990);
or U24104 (N_24104,N_23872,N_23938);
and U24105 (N_24105,N_23881,N_23879);
and U24106 (N_24106,N_23939,N_23996);
xnor U24107 (N_24107,N_23902,N_23967);
and U24108 (N_24108,N_23842,N_23930);
nand U24109 (N_24109,N_23879,N_23986);
nor U24110 (N_24110,N_23869,N_23821);
nor U24111 (N_24111,N_23822,N_23983);
or U24112 (N_24112,N_23854,N_23801);
or U24113 (N_24113,N_23907,N_23828);
and U24114 (N_24114,N_23842,N_23840);
nor U24115 (N_24115,N_23838,N_23934);
nor U24116 (N_24116,N_23977,N_23893);
nor U24117 (N_24117,N_23922,N_23863);
xor U24118 (N_24118,N_23928,N_23941);
nor U24119 (N_24119,N_23854,N_23819);
nor U24120 (N_24120,N_23819,N_23830);
and U24121 (N_24121,N_23810,N_23960);
and U24122 (N_24122,N_23898,N_23866);
and U24123 (N_24123,N_23907,N_23943);
nand U24124 (N_24124,N_23999,N_23907);
nor U24125 (N_24125,N_23875,N_23806);
xnor U24126 (N_24126,N_23945,N_23818);
xnor U24127 (N_24127,N_23967,N_23931);
xor U24128 (N_24128,N_23992,N_23926);
nand U24129 (N_24129,N_23800,N_23895);
nor U24130 (N_24130,N_23948,N_23959);
nand U24131 (N_24131,N_23994,N_23936);
nor U24132 (N_24132,N_23867,N_23822);
nand U24133 (N_24133,N_23868,N_23838);
nand U24134 (N_24134,N_23899,N_23807);
nand U24135 (N_24135,N_23914,N_23805);
xor U24136 (N_24136,N_23980,N_23905);
nand U24137 (N_24137,N_23853,N_23870);
nor U24138 (N_24138,N_23946,N_23894);
and U24139 (N_24139,N_23843,N_23968);
and U24140 (N_24140,N_23882,N_23904);
nor U24141 (N_24141,N_23973,N_23882);
nor U24142 (N_24142,N_23908,N_23828);
xor U24143 (N_24143,N_23904,N_23849);
or U24144 (N_24144,N_23868,N_23958);
xnor U24145 (N_24145,N_23991,N_23880);
and U24146 (N_24146,N_23865,N_23816);
xnor U24147 (N_24147,N_23990,N_23984);
nor U24148 (N_24148,N_23962,N_23998);
nand U24149 (N_24149,N_23898,N_23892);
or U24150 (N_24150,N_23822,N_23930);
or U24151 (N_24151,N_23975,N_23850);
or U24152 (N_24152,N_23864,N_23947);
nand U24153 (N_24153,N_23908,N_23855);
xnor U24154 (N_24154,N_23979,N_23961);
or U24155 (N_24155,N_23879,N_23882);
and U24156 (N_24156,N_23996,N_23839);
nor U24157 (N_24157,N_23906,N_23843);
nor U24158 (N_24158,N_23921,N_23898);
and U24159 (N_24159,N_23914,N_23998);
and U24160 (N_24160,N_23831,N_23946);
xnor U24161 (N_24161,N_23888,N_23832);
xor U24162 (N_24162,N_23878,N_23927);
nand U24163 (N_24163,N_23818,N_23903);
nand U24164 (N_24164,N_23966,N_23996);
xor U24165 (N_24165,N_23990,N_23996);
and U24166 (N_24166,N_23834,N_23840);
or U24167 (N_24167,N_23884,N_23995);
nor U24168 (N_24168,N_23873,N_23998);
xnor U24169 (N_24169,N_23831,N_23917);
nor U24170 (N_24170,N_23946,N_23988);
nand U24171 (N_24171,N_23881,N_23973);
and U24172 (N_24172,N_23863,N_23912);
and U24173 (N_24173,N_23828,N_23843);
nand U24174 (N_24174,N_23950,N_23866);
or U24175 (N_24175,N_23861,N_23992);
xnor U24176 (N_24176,N_23982,N_23924);
xnor U24177 (N_24177,N_23999,N_23812);
or U24178 (N_24178,N_23937,N_23928);
and U24179 (N_24179,N_23837,N_23820);
xor U24180 (N_24180,N_23832,N_23893);
xnor U24181 (N_24181,N_23811,N_23922);
or U24182 (N_24182,N_23839,N_23848);
xnor U24183 (N_24183,N_23854,N_23830);
nand U24184 (N_24184,N_23894,N_23882);
nor U24185 (N_24185,N_23944,N_23868);
xnor U24186 (N_24186,N_23838,N_23818);
or U24187 (N_24187,N_23834,N_23910);
nand U24188 (N_24188,N_23998,N_23831);
and U24189 (N_24189,N_23943,N_23958);
or U24190 (N_24190,N_23910,N_23837);
xnor U24191 (N_24191,N_23913,N_23942);
nor U24192 (N_24192,N_23926,N_23815);
xnor U24193 (N_24193,N_23827,N_23900);
nand U24194 (N_24194,N_23864,N_23944);
and U24195 (N_24195,N_23921,N_23913);
and U24196 (N_24196,N_23975,N_23961);
nor U24197 (N_24197,N_23824,N_23858);
or U24198 (N_24198,N_23944,N_23856);
xnor U24199 (N_24199,N_23859,N_23879);
nand U24200 (N_24200,N_24150,N_24161);
nor U24201 (N_24201,N_24101,N_24191);
nor U24202 (N_24202,N_24030,N_24044);
or U24203 (N_24203,N_24052,N_24100);
nand U24204 (N_24204,N_24039,N_24173);
xor U24205 (N_24205,N_24187,N_24045);
and U24206 (N_24206,N_24199,N_24051);
nand U24207 (N_24207,N_24128,N_24165);
xnor U24208 (N_24208,N_24089,N_24195);
nand U24209 (N_24209,N_24167,N_24090);
and U24210 (N_24210,N_24036,N_24061);
nor U24211 (N_24211,N_24124,N_24169);
nor U24212 (N_24212,N_24086,N_24143);
nand U24213 (N_24213,N_24159,N_24157);
nand U24214 (N_24214,N_24062,N_24151);
or U24215 (N_24215,N_24164,N_24155);
xor U24216 (N_24216,N_24088,N_24171);
nor U24217 (N_24217,N_24107,N_24007);
xor U24218 (N_24218,N_24129,N_24182);
nand U24219 (N_24219,N_24015,N_24192);
or U24220 (N_24220,N_24053,N_24183);
or U24221 (N_24221,N_24131,N_24168);
nor U24222 (N_24222,N_24041,N_24175);
nand U24223 (N_24223,N_24026,N_24114);
xor U24224 (N_24224,N_24189,N_24034);
or U24225 (N_24225,N_24125,N_24081);
or U24226 (N_24226,N_24198,N_24013);
nand U24227 (N_24227,N_24120,N_24091);
nand U24228 (N_24228,N_24006,N_24003);
xnor U24229 (N_24229,N_24098,N_24064);
nand U24230 (N_24230,N_24126,N_24180);
nand U24231 (N_24231,N_24074,N_24139);
nor U24232 (N_24232,N_24134,N_24084);
xor U24233 (N_24233,N_24014,N_24141);
nand U24234 (N_24234,N_24079,N_24020);
or U24235 (N_24235,N_24033,N_24135);
nor U24236 (N_24236,N_24188,N_24035);
or U24237 (N_24237,N_24138,N_24093);
xnor U24238 (N_24238,N_24092,N_24067);
and U24239 (N_24239,N_24016,N_24179);
and U24240 (N_24240,N_24163,N_24121);
nand U24241 (N_24241,N_24184,N_24117);
xor U24242 (N_24242,N_24148,N_24075);
and U24243 (N_24243,N_24024,N_24057);
xnor U24244 (N_24244,N_24031,N_24108);
and U24245 (N_24245,N_24076,N_24038);
xor U24246 (N_24246,N_24008,N_24087);
and U24247 (N_24247,N_24160,N_24118);
nor U24248 (N_24248,N_24162,N_24028);
xnor U24249 (N_24249,N_24110,N_24021);
nand U24250 (N_24250,N_24048,N_24178);
nand U24251 (N_24251,N_24085,N_24001);
and U24252 (N_24252,N_24037,N_24097);
nand U24253 (N_24253,N_24146,N_24104);
and U24254 (N_24254,N_24166,N_24082);
nand U24255 (N_24255,N_24054,N_24002);
nand U24256 (N_24256,N_24049,N_24043);
and U24257 (N_24257,N_24042,N_24066);
and U24258 (N_24258,N_24127,N_24158);
nor U24259 (N_24259,N_24176,N_24113);
xnor U24260 (N_24260,N_24156,N_24144);
and U24261 (N_24261,N_24019,N_24046);
xor U24262 (N_24262,N_24000,N_24172);
nand U24263 (N_24263,N_24147,N_24185);
or U24264 (N_24264,N_24149,N_24077);
and U24265 (N_24265,N_24105,N_24027);
and U24266 (N_24266,N_24122,N_24071);
and U24267 (N_24267,N_24050,N_24083);
nand U24268 (N_24268,N_24196,N_24029);
nor U24269 (N_24269,N_24080,N_24130);
nor U24270 (N_24270,N_24136,N_24137);
or U24271 (N_24271,N_24186,N_24116);
nor U24272 (N_24272,N_24142,N_24004);
or U24273 (N_24273,N_24010,N_24111);
and U24274 (N_24274,N_24056,N_24023);
and U24275 (N_24275,N_24055,N_24119);
xnor U24276 (N_24276,N_24099,N_24132);
nor U24277 (N_24277,N_24068,N_24194);
nand U24278 (N_24278,N_24022,N_24005);
nand U24279 (N_24279,N_24115,N_24177);
and U24280 (N_24280,N_24154,N_24058);
xnor U24281 (N_24281,N_24190,N_24009);
nor U24282 (N_24282,N_24102,N_24047);
and U24283 (N_24283,N_24078,N_24040);
nand U24284 (N_24284,N_24152,N_24109);
nand U24285 (N_24285,N_24123,N_24181);
nor U24286 (N_24286,N_24193,N_24096);
and U24287 (N_24287,N_24059,N_24017);
nand U24288 (N_24288,N_24095,N_24025);
or U24289 (N_24289,N_24103,N_24063);
xnor U24290 (N_24290,N_24032,N_24106);
nor U24291 (N_24291,N_24073,N_24153);
and U24292 (N_24292,N_24065,N_24170);
and U24293 (N_24293,N_24069,N_24133);
nor U24294 (N_24294,N_24070,N_24112);
xor U24295 (N_24295,N_24197,N_24140);
nor U24296 (N_24296,N_24060,N_24012);
nor U24297 (N_24297,N_24072,N_24011);
nand U24298 (N_24298,N_24145,N_24094);
nor U24299 (N_24299,N_24018,N_24174);
and U24300 (N_24300,N_24175,N_24088);
and U24301 (N_24301,N_24185,N_24097);
nand U24302 (N_24302,N_24186,N_24140);
nand U24303 (N_24303,N_24100,N_24130);
nor U24304 (N_24304,N_24153,N_24026);
nand U24305 (N_24305,N_24017,N_24146);
and U24306 (N_24306,N_24121,N_24147);
xor U24307 (N_24307,N_24196,N_24057);
nand U24308 (N_24308,N_24123,N_24086);
nand U24309 (N_24309,N_24034,N_24194);
xnor U24310 (N_24310,N_24153,N_24185);
xor U24311 (N_24311,N_24108,N_24062);
or U24312 (N_24312,N_24001,N_24065);
nand U24313 (N_24313,N_24074,N_24082);
or U24314 (N_24314,N_24000,N_24188);
nor U24315 (N_24315,N_24025,N_24015);
nor U24316 (N_24316,N_24003,N_24108);
nor U24317 (N_24317,N_24018,N_24159);
nor U24318 (N_24318,N_24028,N_24076);
and U24319 (N_24319,N_24175,N_24066);
and U24320 (N_24320,N_24008,N_24042);
nor U24321 (N_24321,N_24036,N_24102);
and U24322 (N_24322,N_24138,N_24102);
xnor U24323 (N_24323,N_24061,N_24078);
xnor U24324 (N_24324,N_24147,N_24106);
nor U24325 (N_24325,N_24057,N_24108);
xnor U24326 (N_24326,N_24141,N_24096);
nand U24327 (N_24327,N_24080,N_24140);
nand U24328 (N_24328,N_24139,N_24127);
xor U24329 (N_24329,N_24090,N_24030);
nand U24330 (N_24330,N_24084,N_24025);
or U24331 (N_24331,N_24060,N_24144);
nor U24332 (N_24332,N_24178,N_24148);
or U24333 (N_24333,N_24187,N_24083);
or U24334 (N_24334,N_24098,N_24129);
or U24335 (N_24335,N_24170,N_24071);
and U24336 (N_24336,N_24067,N_24193);
or U24337 (N_24337,N_24158,N_24060);
xnor U24338 (N_24338,N_24045,N_24103);
or U24339 (N_24339,N_24042,N_24101);
nor U24340 (N_24340,N_24140,N_24130);
and U24341 (N_24341,N_24163,N_24074);
or U24342 (N_24342,N_24125,N_24194);
nand U24343 (N_24343,N_24124,N_24005);
and U24344 (N_24344,N_24181,N_24038);
and U24345 (N_24345,N_24040,N_24049);
xnor U24346 (N_24346,N_24070,N_24196);
and U24347 (N_24347,N_24094,N_24121);
nor U24348 (N_24348,N_24187,N_24167);
nand U24349 (N_24349,N_24102,N_24008);
xor U24350 (N_24350,N_24054,N_24179);
nand U24351 (N_24351,N_24031,N_24182);
nand U24352 (N_24352,N_24076,N_24140);
nor U24353 (N_24353,N_24155,N_24089);
nand U24354 (N_24354,N_24135,N_24182);
xnor U24355 (N_24355,N_24155,N_24059);
or U24356 (N_24356,N_24153,N_24031);
or U24357 (N_24357,N_24095,N_24188);
nand U24358 (N_24358,N_24178,N_24012);
and U24359 (N_24359,N_24159,N_24111);
or U24360 (N_24360,N_24057,N_24149);
and U24361 (N_24361,N_24196,N_24093);
xor U24362 (N_24362,N_24131,N_24158);
and U24363 (N_24363,N_24136,N_24075);
and U24364 (N_24364,N_24198,N_24150);
xor U24365 (N_24365,N_24028,N_24151);
and U24366 (N_24366,N_24081,N_24010);
and U24367 (N_24367,N_24143,N_24005);
nand U24368 (N_24368,N_24130,N_24102);
and U24369 (N_24369,N_24084,N_24131);
nand U24370 (N_24370,N_24091,N_24021);
nand U24371 (N_24371,N_24115,N_24119);
or U24372 (N_24372,N_24001,N_24067);
nor U24373 (N_24373,N_24087,N_24184);
nor U24374 (N_24374,N_24013,N_24020);
and U24375 (N_24375,N_24160,N_24192);
and U24376 (N_24376,N_24148,N_24131);
nand U24377 (N_24377,N_24152,N_24149);
nor U24378 (N_24378,N_24185,N_24197);
nand U24379 (N_24379,N_24187,N_24137);
and U24380 (N_24380,N_24054,N_24137);
or U24381 (N_24381,N_24072,N_24036);
nand U24382 (N_24382,N_24186,N_24081);
and U24383 (N_24383,N_24001,N_24052);
xor U24384 (N_24384,N_24107,N_24035);
nand U24385 (N_24385,N_24016,N_24062);
xnor U24386 (N_24386,N_24003,N_24027);
nor U24387 (N_24387,N_24098,N_24155);
nand U24388 (N_24388,N_24179,N_24166);
nor U24389 (N_24389,N_24181,N_24108);
or U24390 (N_24390,N_24142,N_24120);
nor U24391 (N_24391,N_24007,N_24034);
xor U24392 (N_24392,N_24185,N_24157);
and U24393 (N_24393,N_24183,N_24196);
nand U24394 (N_24394,N_24075,N_24018);
or U24395 (N_24395,N_24028,N_24173);
or U24396 (N_24396,N_24071,N_24002);
nand U24397 (N_24397,N_24069,N_24112);
nor U24398 (N_24398,N_24005,N_24090);
nand U24399 (N_24399,N_24087,N_24075);
nand U24400 (N_24400,N_24299,N_24374);
xor U24401 (N_24401,N_24208,N_24379);
nand U24402 (N_24402,N_24389,N_24238);
and U24403 (N_24403,N_24306,N_24336);
nor U24404 (N_24404,N_24248,N_24214);
nor U24405 (N_24405,N_24275,N_24337);
nand U24406 (N_24406,N_24213,N_24304);
or U24407 (N_24407,N_24329,N_24204);
nand U24408 (N_24408,N_24367,N_24294);
xnor U24409 (N_24409,N_24350,N_24313);
nor U24410 (N_24410,N_24369,N_24200);
xnor U24411 (N_24411,N_24316,N_24257);
nand U24412 (N_24412,N_24381,N_24284);
xor U24413 (N_24413,N_24289,N_24397);
and U24414 (N_24414,N_24301,N_24236);
and U24415 (N_24415,N_24395,N_24211);
nand U24416 (N_24416,N_24378,N_24258);
or U24417 (N_24417,N_24383,N_24298);
nand U24418 (N_24418,N_24382,N_24344);
or U24419 (N_24419,N_24287,N_24387);
nand U24420 (N_24420,N_24376,N_24203);
and U24421 (N_24421,N_24326,N_24283);
and U24422 (N_24422,N_24372,N_24218);
xor U24423 (N_24423,N_24239,N_24232);
and U24424 (N_24424,N_24245,N_24362);
nor U24425 (N_24425,N_24396,N_24302);
nor U24426 (N_24426,N_24278,N_24332);
nand U24427 (N_24427,N_24207,N_24343);
xor U24428 (N_24428,N_24240,N_24235);
or U24429 (N_24429,N_24386,N_24361);
nor U24430 (N_24430,N_24251,N_24360);
xor U24431 (N_24431,N_24388,N_24206);
nand U24432 (N_24432,N_24308,N_24384);
xnor U24433 (N_24433,N_24286,N_24233);
nor U24434 (N_24434,N_24249,N_24314);
xnor U24435 (N_24435,N_24255,N_24391);
xnor U24436 (N_24436,N_24228,N_24315);
and U24437 (N_24437,N_24277,N_24370);
nand U24438 (N_24438,N_24288,N_24338);
nor U24439 (N_24439,N_24323,N_24265);
nor U24440 (N_24440,N_24358,N_24312);
nor U24441 (N_24441,N_24242,N_24216);
xor U24442 (N_24442,N_24346,N_24311);
nand U24443 (N_24443,N_24296,N_24340);
nand U24444 (N_24444,N_24366,N_24223);
nor U24445 (N_24445,N_24279,N_24254);
or U24446 (N_24446,N_24303,N_24318);
and U24447 (N_24447,N_24307,N_24247);
nand U24448 (N_24448,N_24345,N_24225);
nand U24449 (N_24449,N_24230,N_24349);
nand U24450 (N_24450,N_24226,N_24359);
and U24451 (N_24451,N_24231,N_24319);
nand U24452 (N_24452,N_24244,N_24259);
nand U24453 (N_24453,N_24263,N_24300);
and U24454 (N_24454,N_24377,N_24268);
nor U24455 (N_24455,N_24357,N_24217);
nand U24456 (N_24456,N_24210,N_24321);
or U24457 (N_24457,N_24348,N_24237);
xor U24458 (N_24458,N_24260,N_24354);
and U24459 (N_24459,N_24241,N_24253);
nand U24460 (N_24460,N_24324,N_24327);
nand U24461 (N_24461,N_24272,N_24398);
or U24462 (N_24462,N_24293,N_24333);
nor U24463 (N_24463,N_24385,N_24202);
and U24464 (N_24464,N_24205,N_24262);
nand U24465 (N_24465,N_24274,N_24365);
and U24466 (N_24466,N_24291,N_24234);
nand U24467 (N_24467,N_24317,N_24276);
and U24468 (N_24468,N_24305,N_24281);
nand U24469 (N_24469,N_24285,N_24328);
or U24470 (N_24470,N_24339,N_24364);
nor U24471 (N_24471,N_24331,N_24341);
and U24472 (N_24472,N_24355,N_24243);
nor U24473 (N_24473,N_24256,N_24394);
nand U24474 (N_24474,N_24290,N_24282);
nand U24475 (N_24475,N_24371,N_24273);
and U24476 (N_24476,N_24224,N_24246);
xnor U24477 (N_24477,N_24222,N_24250);
xor U24478 (N_24478,N_24269,N_24352);
xnor U24479 (N_24479,N_24229,N_24220);
nor U24480 (N_24480,N_24330,N_24297);
and U24481 (N_24481,N_24270,N_24266);
nor U24482 (N_24482,N_24310,N_24322);
or U24483 (N_24483,N_24267,N_24252);
nor U24484 (N_24484,N_24221,N_24219);
nor U24485 (N_24485,N_24390,N_24215);
or U24486 (N_24486,N_24261,N_24201);
xnor U24487 (N_24487,N_24368,N_24271);
or U24488 (N_24488,N_24356,N_24227);
and U24489 (N_24489,N_24351,N_24373);
nand U24490 (N_24490,N_24399,N_24212);
or U24491 (N_24491,N_24209,N_24292);
and U24492 (N_24492,N_24320,N_24280);
nand U24493 (N_24493,N_24392,N_24380);
xor U24494 (N_24494,N_24353,N_24375);
or U24495 (N_24495,N_24295,N_24342);
nor U24496 (N_24496,N_24264,N_24363);
nand U24497 (N_24497,N_24309,N_24335);
or U24498 (N_24498,N_24325,N_24393);
and U24499 (N_24499,N_24347,N_24334);
and U24500 (N_24500,N_24342,N_24321);
nand U24501 (N_24501,N_24226,N_24296);
xnor U24502 (N_24502,N_24219,N_24382);
xnor U24503 (N_24503,N_24275,N_24246);
xor U24504 (N_24504,N_24286,N_24305);
and U24505 (N_24505,N_24291,N_24239);
nor U24506 (N_24506,N_24222,N_24372);
or U24507 (N_24507,N_24304,N_24230);
nand U24508 (N_24508,N_24397,N_24385);
and U24509 (N_24509,N_24378,N_24314);
nand U24510 (N_24510,N_24338,N_24376);
or U24511 (N_24511,N_24208,N_24218);
and U24512 (N_24512,N_24396,N_24307);
or U24513 (N_24513,N_24266,N_24252);
nor U24514 (N_24514,N_24327,N_24241);
nand U24515 (N_24515,N_24311,N_24264);
and U24516 (N_24516,N_24362,N_24275);
or U24517 (N_24517,N_24216,N_24390);
nor U24518 (N_24518,N_24343,N_24323);
nand U24519 (N_24519,N_24219,N_24398);
and U24520 (N_24520,N_24248,N_24279);
or U24521 (N_24521,N_24266,N_24246);
or U24522 (N_24522,N_24357,N_24320);
nor U24523 (N_24523,N_24271,N_24386);
and U24524 (N_24524,N_24374,N_24354);
nor U24525 (N_24525,N_24232,N_24235);
nand U24526 (N_24526,N_24320,N_24266);
and U24527 (N_24527,N_24327,N_24203);
and U24528 (N_24528,N_24257,N_24381);
nor U24529 (N_24529,N_24225,N_24315);
and U24530 (N_24530,N_24263,N_24248);
nor U24531 (N_24531,N_24368,N_24362);
nor U24532 (N_24532,N_24289,N_24382);
xnor U24533 (N_24533,N_24301,N_24359);
and U24534 (N_24534,N_24317,N_24354);
or U24535 (N_24535,N_24224,N_24323);
and U24536 (N_24536,N_24305,N_24227);
xor U24537 (N_24537,N_24203,N_24368);
nor U24538 (N_24538,N_24399,N_24321);
or U24539 (N_24539,N_24241,N_24296);
nand U24540 (N_24540,N_24341,N_24343);
and U24541 (N_24541,N_24248,N_24328);
and U24542 (N_24542,N_24378,N_24338);
nor U24543 (N_24543,N_24208,N_24310);
nand U24544 (N_24544,N_24324,N_24246);
nand U24545 (N_24545,N_24260,N_24307);
or U24546 (N_24546,N_24390,N_24317);
nor U24547 (N_24547,N_24329,N_24206);
or U24548 (N_24548,N_24263,N_24379);
nand U24549 (N_24549,N_24341,N_24359);
and U24550 (N_24550,N_24345,N_24260);
and U24551 (N_24551,N_24290,N_24279);
nor U24552 (N_24552,N_24297,N_24390);
nor U24553 (N_24553,N_24340,N_24323);
nor U24554 (N_24554,N_24328,N_24331);
nor U24555 (N_24555,N_24379,N_24265);
xor U24556 (N_24556,N_24393,N_24271);
or U24557 (N_24557,N_24228,N_24201);
xnor U24558 (N_24558,N_24275,N_24312);
nand U24559 (N_24559,N_24348,N_24391);
nand U24560 (N_24560,N_24261,N_24319);
xor U24561 (N_24561,N_24385,N_24264);
or U24562 (N_24562,N_24293,N_24390);
nor U24563 (N_24563,N_24361,N_24304);
xnor U24564 (N_24564,N_24245,N_24228);
xnor U24565 (N_24565,N_24294,N_24206);
or U24566 (N_24566,N_24372,N_24201);
xor U24567 (N_24567,N_24263,N_24284);
xor U24568 (N_24568,N_24369,N_24202);
or U24569 (N_24569,N_24336,N_24397);
and U24570 (N_24570,N_24340,N_24335);
and U24571 (N_24571,N_24319,N_24347);
or U24572 (N_24572,N_24328,N_24349);
or U24573 (N_24573,N_24238,N_24229);
xnor U24574 (N_24574,N_24371,N_24315);
nand U24575 (N_24575,N_24327,N_24298);
xnor U24576 (N_24576,N_24370,N_24225);
and U24577 (N_24577,N_24305,N_24275);
and U24578 (N_24578,N_24395,N_24202);
nand U24579 (N_24579,N_24209,N_24278);
xnor U24580 (N_24580,N_24389,N_24335);
and U24581 (N_24581,N_24391,N_24351);
xnor U24582 (N_24582,N_24277,N_24269);
and U24583 (N_24583,N_24248,N_24270);
nor U24584 (N_24584,N_24315,N_24295);
nand U24585 (N_24585,N_24246,N_24357);
nor U24586 (N_24586,N_24219,N_24251);
xor U24587 (N_24587,N_24212,N_24324);
and U24588 (N_24588,N_24250,N_24362);
nand U24589 (N_24589,N_24252,N_24398);
and U24590 (N_24590,N_24377,N_24312);
nor U24591 (N_24591,N_24297,N_24342);
or U24592 (N_24592,N_24399,N_24395);
xnor U24593 (N_24593,N_24281,N_24327);
nor U24594 (N_24594,N_24250,N_24300);
nor U24595 (N_24595,N_24280,N_24254);
nor U24596 (N_24596,N_24234,N_24377);
or U24597 (N_24597,N_24370,N_24226);
and U24598 (N_24598,N_24350,N_24222);
nand U24599 (N_24599,N_24385,N_24210);
xnor U24600 (N_24600,N_24439,N_24415);
and U24601 (N_24601,N_24599,N_24561);
and U24602 (N_24602,N_24466,N_24464);
or U24603 (N_24603,N_24526,N_24481);
nand U24604 (N_24604,N_24504,N_24465);
and U24605 (N_24605,N_24498,N_24545);
nand U24606 (N_24606,N_24578,N_24424);
or U24607 (N_24607,N_24570,N_24543);
xnor U24608 (N_24608,N_24403,N_24468);
xnor U24609 (N_24609,N_24477,N_24434);
nand U24610 (N_24610,N_24556,N_24420);
and U24611 (N_24611,N_24523,N_24512);
nor U24612 (N_24612,N_24432,N_24520);
or U24613 (N_24613,N_24429,N_24503);
xor U24614 (N_24614,N_24551,N_24472);
nand U24615 (N_24615,N_24544,N_24590);
nand U24616 (N_24616,N_24492,N_24531);
nor U24617 (N_24617,N_24530,N_24584);
and U24618 (N_24618,N_24427,N_24425);
and U24619 (N_24619,N_24594,N_24488);
xnor U24620 (N_24620,N_24490,N_24513);
and U24621 (N_24621,N_24564,N_24536);
nand U24622 (N_24622,N_24487,N_24474);
and U24623 (N_24623,N_24532,N_24524);
nor U24624 (N_24624,N_24446,N_24529);
nand U24625 (N_24625,N_24400,N_24593);
nand U24626 (N_24626,N_24552,N_24527);
xnor U24627 (N_24627,N_24500,N_24461);
nand U24628 (N_24628,N_24408,N_24563);
xnor U24629 (N_24629,N_24582,N_24473);
nor U24630 (N_24630,N_24486,N_24585);
nor U24631 (N_24631,N_24575,N_24452);
xnor U24632 (N_24632,N_24562,N_24489);
nor U24633 (N_24633,N_24597,N_24505);
or U24634 (N_24634,N_24588,N_24565);
and U24635 (N_24635,N_24480,N_24516);
and U24636 (N_24636,N_24550,N_24525);
and U24637 (N_24637,N_24411,N_24440);
nor U24638 (N_24638,N_24514,N_24482);
xnor U24639 (N_24639,N_24463,N_24540);
xor U24640 (N_24640,N_24412,N_24535);
and U24641 (N_24641,N_24428,N_24443);
xor U24642 (N_24642,N_24483,N_24515);
nand U24643 (N_24643,N_24426,N_24406);
xnor U24644 (N_24644,N_24438,N_24401);
nand U24645 (N_24645,N_24572,N_24542);
and U24646 (N_24646,N_24413,N_24587);
or U24647 (N_24647,N_24499,N_24559);
xnor U24648 (N_24648,N_24453,N_24435);
nor U24649 (N_24649,N_24557,N_24478);
or U24650 (N_24650,N_24580,N_24437);
nand U24651 (N_24651,N_24508,N_24475);
nand U24652 (N_24652,N_24414,N_24448);
nand U24653 (N_24653,N_24574,N_24460);
xor U24654 (N_24654,N_24433,N_24581);
xnor U24655 (N_24655,N_24534,N_24491);
xnor U24656 (N_24656,N_24471,N_24502);
or U24657 (N_24657,N_24476,N_24469);
nand U24658 (N_24658,N_24589,N_24467);
nand U24659 (N_24659,N_24571,N_24553);
or U24660 (N_24660,N_24456,N_24549);
xor U24661 (N_24661,N_24509,N_24450);
xnor U24662 (N_24662,N_24409,N_24577);
or U24663 (N_24663,N_24459,N_24410);
xor U24664 (N_24664,N_24442,N_24539);
or U24665 (N_24665,N_24555,N_24598);
nor U24666 (N_24666,N_24506,N_24449);
xor U24667 (N_24667,N_24454,N_24547);
or U24668 (N_24668,N_24576,N_24533);
or U24669 (N_24669,N_24518,N_24430);
xnor U24670 (N_24670,N_24507,N_24405);
and U24671 (N_24671,N_24591,N_24583);
nor U24672 (N_24672,N_24521,N_24519);
xnor U24673 (N_24673,N_24423,N_24541);
xnor U24674 (N_24674,N_24479,N_24485);
nand U24675 (N_24675,N_24548,N_24595);
and U24676 (N_24676,N_24447,N_24579);
and U24677 (N_24677,N_24431,N_24457);
or U24678 (N_24678,N_24455,N_24569);
nor U24679 (N_24679,N_24511,N_24497);
or U24680 (N_24680,N_24441,N_24451);
xor U24681 (N_24681,N_24493,N_24404);
nor U24682 (N_24682,N_24554,N_24596);
or U24683 (N_24683,N_24470,N_24592);
nand U24684 (N_24684,N_24402,N_24528);
xor U24685 (N_24685,N_24510,N_24501);
nor U24686 (N_24686,N_24418,N_24537);
xnor U24687 (N_24687,N_24422,N_24444);
and U24688 (N_24688,N_24560,N_24566);
or U24689 (N_24689,N_24496,N_24436);
or U24690 (N_24690,N_24407,N_24494);
or U24691 (N_24691,N_24445,N_24573);
nor U24692 (N_24692,N_24416,N_24568);
and U24693 (N_24693,N_24419,N_24517);
xnor U24694 (N_24694,N_24421,N_24417);
and U24695 (N_24695,N_24546,N_24567);
nor U24696 (N_24696,N_24484,N_24538);
nand U24697 (N_24697,N_24558,N_24462);
nand U24698 (N_24698,N_24495,N_24586);
xor U24699 (N_24699,N_24522,N_24458);
xnor U24700 (N_24700,N_24439,N_24450);
or U24701 (N_24701,N_24584,N_24564);
nor U24702 (N_24702,N_24520,N_24591);
or U24703 (N_24703,N_24491,N_24540);
xnor U24704 (N_24704,N_24413,N_24580);
nor U24705 (N_24705,N_24444,N_24409);
or U24706 (N_24706,N_24553,N_24539);
or U24707 (N_24707,N_24510,N_24476);
or U24708 (N_24708,N_24599,N_24540);
nor U24709 (N_24709,N_24404,N_24406);
and U24710 (N_24710,N_24415,N_24553);
xnor U24711 (N_24711,N_24510,N_24465);
or U24712 (N_24712,N_24401,N_24416);
nor U24713 (N_24713,N_24510,N_24401);
and U24714 (N_24714,N_24523,N_24573);
and U24715 (N_24715,N_24531,N_24470);
or U24716 (N_24716,N_24430,N_24447);
or U24717 (N_24717,N_24430,N_24469);
and U24718 (N_24718,N_24424,N_24455);
xor U24719 (N_24719,N_24573,N_24550);
nor U24720 (N_24720,N_24512,N_24578);
xnor U24721 (N_24721,N_24454,N_24432);
xnor U24722 (N_24722,N_24542,N_24460);
nor U24723 (N_24723,N_24442,N_24535);
or U24724 (N_24724,N_24401,N_24410);
nand U24725 (N_24725,N_24465,N_24411);
and U24726 (N_24726,N_24505,N_24576);
xnor U24727 (N_24727,N_24470,N_24439);
nand U24728 (N_24728,N_24495,N_24405);
or U24729 (N_24729,N_24417,N_24535);
and U24730 (N_24730,N_24471,N_24567);
or U24731 (N_24731,N_24409,N_24587);
nand U24732 (N_24732,N_24528,N_24589);
and U24733 (N_24733,N_24479,N_24421);
and U24734 (N_24734,N_24449,N_24427);
nor U24735 (N_24735,N_24467,N_24432);
xnor U24736 (N_24736,N_24461,N_24549);
and U24737 (N_24737,N_24444,N_24459);
nand U24738 (N_24738,N_24465,N_24435);
or U24739 (N_24739,N_24567,N_24474);
or U24740 (N_24740,N_24420,N_24593);
nor U24741 (N_24741,N_24408,N_24543);
or U24742 (N_24742,N_24478,N_24452);
xor U24743 (N_24743,N_24563,N_24559);
and U24744 (N_24744,N_24472,N_24448);
and U24745 (N_24745,N_24551,N_24470);
or U24746 (N_24746,N_24493,N_24583);
or U24747 (N_24747,N_24581,N_24517);
xor U24748 (N_24748,N_24524,N_24520);
nor U24749 (N_24749,N_24594,N_24412);
xnor U24750 (N_24750,N_24487,N_24421);
xor U24751 (N_24751,N_24590,N_24524);
xnor U24752 (N_24752,N_24507,N_24573);
xnor U24753 (N_24753,N_24551,N_24550);
nor U24754 (N_24754,N_24465,N_24509);
and U24755 (N_24755,N_24419,N_24495);
nor U24756 (N_24756,N_24462,N_24524);
and U24757 (N_24757,N_24512,N_24401);
or U24758 (N_24758,N_24455,N_24412);
xor U24759 (N_24759,N_24420,N_24466);
xor U24760 (N_24760,N_24511,N_24414);
nand U24761 (N_24761,N_24446,N_24441);
or U24762 (N_24762,N_24580,N_24597);
or U24763 (N_24763,N_24470,N_24505);
and U24764 (N_24764,N_24437,N_24587);
nor U24765 (N_24765,N_24578,N_24532);
nand U24766 (N_24766,N_24582,N_24442);
nor U24767 (N_24767,N_24596,N_24498);
and U24768 (N_24768,N_24539,N_24494);
or U24769 (N_24769,N_24575,N_24482);
nand U24770 (N_24770,N_24464,N_24491);
nor U24771 (N_24771,N_24554,N_24469);
nor U24772 (N_24772,N_24504,N_24500);
nand U24773 (N_24773,N_24443,N_24543);
nand U24774 (N_24774,N_24525,N_24535);
and U24775 (N_24775,N_24571,N_24584);
xnor U24776 (N_24776,N_24479,N_24517);
and U24777 (N_24777,N_24576,N_24405);
xnor U24778 (N_24778,N_24469,N_24447);
nor U24779 (N_24779,N_24410,N_24540);
nor U24780 (N_24780,N_24537,N_24406);
nand U24781 (N_24781,N_24438,N_24423);
nor U24782 (N_24782,N_24558,N_24523);
and U24783 (N_24783,N_24428,N_24472);
and U24784 (N_24784,N_24544,N_24549);
nand U24785 (N_24785,N_24587,N_24527);
nor U24786 (N_24786,N_24474,N_24566);
and U24787 (N_24787,N_24454,N_24412);
or U24788 (N_24788,N_24493,N_24487);
nor U24789 (N_24789,N_24444,N_24519);
nor U24790 (N_24790,N_24497,N_24585);
nor U24791 (N_24791,N_24425,N_24460);
and U24792 (N_24792,N_24516,N_24529);
or U24793 (N_24793,N_24402,N_24488);
and U24794 (N_24794,N_24596,N_24564);
xor U24795 (N_24795,N_24437,N_24460);
nor U24796 (N_24796,N_24403,N_24470);
or U24797 (N_24797,N_24417,N_24499);
xnor U24798 (N_24798,N_24478,N_24590);
xor U24799 (N_24799,N_24586,N_24550);
nand U24800 (N_24800,N_24676,N_24742);
and U24801 (N_24801,N_24794,N_24758);
xor U24802 (N_24802,N_24799,N_24641);
nor U24803 (N_24803,N_24660,N_24681);
or U24804 (N_24804,N_24619,N_24712);
nand U24805 (N_24805,N_24778,N_24618);
nor U24806 (N_24806,N_24646,N_24614);
nand U24807 (N_24807,N_24622,N_24751);
xnor U24808 (N_24808,N_24736,N_24702);
nor U24809 (N_24809,N_24688,N_24714);
nand U24810 (N_24810,N_24629,N_24666);
or U24811 (N_24811,N_24780,N_24635);
xor U24812 (N_24812,N_24620,N_24766);
xor U24813 (N_24813,N_24643,N_24729);
or U24814 (N_24814,N_24732,N_24683);
xor U24815 (N_24815,N_24670,N_24783);
xor U24816 (N_24816,N_24661,N_24679);
or U24817 (N_24817,N_24690,N_24717);
and U24818 (N_24818,N_24684,N_24790);
nor U24819 (N_24819,N_24750,N_24708);
nor U24820 (N_24820,N_24752,N_24611);
nor U24821 (N_24821,N_24662,N_24623);
and U24822 (N_24822,N_24687,N_24699);
xor U24823 (N_24823,N_24665,N_24686);
nor U24824 (N_24824,N_24604,N_24648);
nand U24825 (N_24825,N_24698,N_24721);
and U24826 (N_24826,N_24703,N_24671);
or U24827 (N_24827,N_24617,N_24645);
and U24828 (N_24828,N_24747,N_24682);
and U24829 (N_24829,N_24624,N_24607);
xnor U24830 (N_24830,N_24696,N_24627);
nor U24831 (N_24831,N_24743,N_24625);
xor U24832 (N_24832,N_24789,N_24773);
xnor U24833 (N_24833,N_24700,N_24785);
or U24834 (N_24834,N_24796,N_24630);
nor U24835 (N_24835,N_24720,N_24707);
xnor U24836 (N_24836,N_24608,N_24644);
and U24837 (N_24837,N_24771,N_24602);
nor U24838 (N_24838,N_24798,N_24672);
and U24839 (N_24839,N_24709,N_24774);
and U24840 (N_24840,N_24705,N_24775);
nor U24841 (N_24841,N_24695,N_24734);
nor U24842 (N_24842,N_24621,N_24718);
or U24843 (N_24843,N_24701,N_24740);
and U24844 (N_24844,N_24784,N_24727);
xnor U24845 (N_24845,N_24777,N_24652);
nand U24846 (N_24846,N_24738,N_24704);
or U24847 (N_24847,N_24741,N_24677);
nand U24848 (N_24848,N_24787,N_24763);
and U24849 (N_24849,N_24745,N_24779);
nor U24850 (N_24850,N_24719,N_24770);
nor U24851 (N_24851,N_24795,N_24768);
or U24852 (N_24852,N_24764,N_24781);
xor U24853 (N_24853,N_24706,N_24782);
and U24854 (N_24854,N_24754,N_24726);
xor U24855 (N_24855,N_24680,N_24767);
nor U24856 (N_24856,N_24694,N_24633);
and U24857 (N_24857,N_24797,N_24689);
nor U24858 (N_24858,N_24728,N_24610);
nor U24859 (N_24859,N_24631,N_24637);
nand U24860 (N_24860,N_24647,N_24668);
nor U24861 (N_24861,N_24716,N_24715);
and U24862 (N_24862,N_24786,N_24697);
nor U24863 (N_24863,N_24769,N_24761);
and U24864 (N_24864,N_24724,N_24649);
nor U24865 (N_24865,N_24659,N_24651);
nand U24866 (N_24866,N_24616,N_24710);
and U24867 (N_24867,N_24737,N_24601);
and U24868 (N_24868,N_24658,N_24691);
or U24869 (N_24869,N_24673,N_24744);
or U24870 (N_24870,N_24674,N_24626);
xor U24871 (N_24871,N_24606,N_24628);
or U24872 (N_24872,N_24739,N_24603);
nand U24873 (N_24873,N_24664,N_24632);
xnor U24874 (N_24874,N_24735,N_24713);
nor U24875 (N_24875,N_24636,N_24791);
nor U24876 (N_24876,N_24772,N_24711);
xnor U24877 (N_24877,N_24667,N_24653);
nand U24878 (N_24878,N_24650,N_24748);
or U24879 (N_24879,N_24759,N_24639);
xor U24880 (N_24880,N_24656,N_24757);
or U24881 (N_24881,N_24756,N_24640);
nor U24882 (N_24882,N_24788,N_24615);
nor U24883 (N_24883,N_24731,N_24600);
nand U24884 (N_24884,N_24793,N_24663);
nor U24885 (N_24885,N_24762,N_24638);
and U24886 (N_24886,N_24612,N_24678);
nand U24887 (N_24887,N_24609,N_24749);
nor U24888 (N_24888,N_24765,N_24605);
nand U24889 (N_24889,N_24792,N_24657);
nand U24890 (N_24890,N_24725,N_24634);
nand U24891 (N_24891,N_24669,N_24675);
nand U24892 (N_24892,N_24753,N_24692);
and U24893 (N_24893,N_24693,N_24655);
xnor U24894 (N_24894,N_24685,N_24722);
xor U24895 (N_24895,N_24613,N_24760);
and U24896 (N_24896,N_24654,N_24746);
xor U24897 (N_24897,N_24723,N_24733);
and U24898 (N_24898,N_24642,N_24776);
xor U24899 (N_24899,N_24730,N_24755);
or U24900 (N_24900,N_24757,N_24742);
nor U24901 (N_24901,N_24652,N_24614);
and U24902 (N_24902,N_24676,N_24648);
nor U24903 (N_24903,N_24763,N_24617);
nor U24904 (N_24904,N_24700,N_24744);
nor U24905 (N_24905,N_24791,N_24648);
or U24906 (N_24906,N_24644,N_24724);
nand U24907 (N_24907,N_24693,N_24737);
nand U24908 (N_24908,N_24610,N_24603);
or U24909 (N_24909,N_24781,N_24794);
nand U24910 (N_24910,N_24624,N_24700);
nor U24911 (N_24911,N_24612,N_24755);
nor U24912 (N_24912,N_24792,N_24790);
nand U24913 (N_24913,N_24765,N_24666);
and U24914 (N_24914,N_24635,N_24657);
xor U24915 (N_24915,N_24753,N_24747);
nor U24916 (N_24916,N_24707,N_24717);
nand U24917 (N_24917,N_24605,N_24628);
xor U24918 (N_24918,N_24750,N_24666);
nand U24919 (N_24919,N_24732,N_24600);
nor U24920 (N_24920,N_24657,N_24636);
nand U24921 (N_24921,N_24779,N_24781);
nand U24922 (N_24922,N_24770,N_24670);
nand U24923 (N_24923,N_24662,N_24630);
nand U24924 (N_24924,N_24690,N_24799);
nor U24925 (N_24925,N_24745,N_24716);
nand U24926 (N_24926,N_24604,N_24753);
or U24927 (N_24927,N_24722,N_24745);
xor U24928 (N_24928,N_24794,N_24689);
nand U24929 (N_24929,N_24736,N_24753);
xnor U24930 (N_24930,N_24668,N_24759);
or U24931 (N_24931,N_24730,N_24671);
xnor U24932 (N_24932,N_24766,N_24699);
and U24933 (N_24933,N_24603,N_24648);
nand U24934 (N_24934,N_24795,N_24704);
nor U24935 (N_24935,N_24604,N_24686);
nand U24936 (N_24936,N_24669,N_24786);
or U24937 (N_24937,N_24660,N_24793);
nand U24938 (N_24938,N_24723,N_24794);
or U24939 (N_24939,N_24647,N_24713);
or U24940 (N_24940,N_24615,N_24750);
or U24941 (N_24941,N_24782,N_24777);
nand U24942 (N_24942,N_24656,N_24743);
xor U24943 (N_24943,N_24705,N_24796);
or U24944 (N_24944,N_24634,N_24717);
nand U24945 (N_24945,N_24667,N_24620);
and U24946 (N_24946,N_24638,N_24765);
xnor U24947 (N_24947,N_24615,N_24695);
or U24948 (N_24948,N_24751,N_24786);
xnor U24949 (N_24949,N_24601,N_24712);
nor U24950 (N_24950,N_24676,N_24692);
nand U24951 (N_24951,N_24668,N_24627);
or U24952 (N_24952,N_24658,N_24752);
nor U24953 (N_24953,N_24661,N_24725);
and U24954 (N_24954,N_24663,N_24654);
nor U24955 (N_24955,N_24778,N_24759);
nand U24956 (N_24956,N_24727,N_24672);
or U24957 (N_24957,N_24611,N_24735);
xor U24958 (N_24958,N_24675,N_24665);
xor U24959 (N_24959,N_24740,N_24718);
nand U24960 (N_24960,N_24787,N_24656);
xor U24961 (N_24961,N_24707,N_24728);
or U24962 (N_24962,N_24661,N_24755);
xor U24963 (N_24963,N_24622,N_24615);
nor U24964 (N_24964,N_24646,N_24766);
nor U24965 (N_24965,N_24721,N_24688);
and U24966 (N_24966,N_24671,N_24624);
and U24967 (N_24967,N_24622,N_24631);
nor U24968 (N_24968,N_24653,N_24731);
and U24969 (N_24969,N_24701,N_24601);
nand U24970 (N_24970,N_24681,N_24677);
nand U24971 (N_24971,N_24799,N_24751);
and U24972 (N_24972,N_24634,N_24637);
or U24973 (N_24973,N_24605,N_24783);
xnor U24974 (N_24974,N_24796,N_24641);
and U24975 (N_24975,N_24637,N_24613);
nor U24976 (N_24976,N_24710,N_24788);
nand U24977 (N_24977,N_24649,N_24651);
or U24978 (N_24978,N_24745,N_24625);
nor U24979 (N_24979,N_24715,N_24620);
xnor U24980 (N_24980,N_24698,N_24629);
and U24981 (N_24981,N_24700,N_24644);
xnor U24982 (N_24982,N_24699,N_24659);
or U24983 (N_24983,N_24745,N_24691);
and U24984 (N_24984,N_24648,N_24744);
nand U24985 (N_24985,N_24641,N_24686);
and U24986 (N_24986,N_24666,N_24775);
nand U24987 (N_24987,N_24715,N_24726);
or U24988 (N_24988,N_24666,N_24693);
and U24989 (N_24989,N_24624,N_24694);
nor U24990 (N_24990,N_24796,N_24681);
and U24991 (N_24991,N_24695,N_24742);
and U24992 (N_24992,N_24794,N_24620);
xor U24993 (N_24993,N_24735,N_24772);
and U24994 (N_24994,N_24691,N_24652);
nand U24995 (N_24995,N_24653,N_24769);
nand U24996 (N_24996,N_24799,N_24631);
xor U24997 (N_24997,N_24661,N_24715);
or U24998 (N_24998,N_24712,N_24613);
nand U24999 (N_24999,N_24730,N_24701);
xnor UO_0 (O_0,N_24867,N_24960);
nor UO_1 (O_1,N_24938,N_24839);
or UO_2 (O_2,N_24900,N_24917);
and UO_3 (O_3,N_24950,N_24937);
or UO_4 (O_4,N_24877,N_24893);
xor UO_5 (O_5,N_24920,N_24857);
and UO_6 (O_6,N_24918,N_24818);
nor UO_7 (O_7,N_24903,N_24946);
xor UO_8 (O_8,N_24922,N_24869);
nand UO_9 (O_9,N_24998,N_24863);
nand UO_10 (O_10,N_24855,N_24913);
nor UO_11 (O_11,N_24813,N_24831);
xor UO_12 (O_12,N_24811,N_24876);
and UO_13 (O_13,N_24866,N_24981);
and UO_14 (O_14,N_24891,N_24934);
or UO_15 (O_15,N_24890,N_24964);
and UO_16 (O_16,N_24865,N_24822);
and UO_17 (O_17,N_24887,N_24993);
nand UO_18 (O_18,N_24898,N_24851);
and UO_19 (O_19,N_24814,N_24962);
nand UO_20 (O_20,N_24809,N_24988);
or UO_21 (O_21,N_24951,N_24933);
nand UO_22 (O_22,N_24910,N_24935);
nor UO_23 (O_23,N_24973,N_24824);
xor UO_24 (O_24,N_24827,N_24908);
or UO_25 (O_25,N_24845,N_24916);
and UO_26 (O_26,N_24833,N_24816);
xor UO_27 (O_27,N_24884,N_24921);
or UO_28 (O_28,N_24996,N_24911);
xnor UO_29 (O_29,N_24906,N_24820);
xnor UO_30 (O_30,N_24840,N_24987);
and UO_31 (O_31,N_24882,N_24800);
or UO_32 (O_32,N_24826,N_24856);
nand UO_33 (O_33,N_24894,N_24956);
nand UO_34 (O_34,N_24928,N_24929);
xnor UO_35 (O_35,N_24999,N_24854);
and UO_36 (O_36,N_24932,N_24807);
nor UO_37 (O_37,N_24909,N_24821);
and UO_38 (O_38,N_24815,N_24927);
nand UO_39 (O_39,N_24888,N_24853);
nand UO_40 (O_40,N_24837,N_24802);
or UO_41 (O_41,N_24850,N_24992);
or UO_42 (O_42,N_24961,N_24889);
and UO_43 (O_43,N_24883,N_24953);
nand UO_44 (O_44,N_24803,N_24819);
and UO_45 (O_45,N_24967,N_24808);
and UO_46 (O_46,N_24955,N_24868);
nand UO_47 (O_47,N_24858,N_24871);
nor UO_48 (O_48,N_24905,N_24849);
xor UO_49 (O_49,N_24968,N_24949);
and UO_50 (O_50,N_24986,N_24995);
or UO_51 (O_51,N_24940,N_24915);
nor UO_52 (O_52,N_24861,N_24944);
xor UO_53 (O_53,N_24991,N_24976);
nand UO_54 (O_54,N_24810,N_24930);
nor UO_55 (O_55,N_24957,N_24972);
or UO_56 (O_56,N_24892,N_24836);
nor UO_57 (O_57,N_24985,N_24805);
and UO_58 (O_58,N_24844,N_24959);
nor UO_59 (O_59,N_24907,N_24952);
and UO_60 (O_60,N_24848,N_24817);
nand UO_61 (O_61,N_24806,N_24901);
nor UO_62 (O_62,N_24945,N_24875);
or UO_63 (O_63,N_24895,N_24970);
nand UO_64 (O_64,N_24980,N_24847);
or UO_65 (O_65,N_24958,N_24879);
xnor UO_66 (O_66,N_24885,N_24864);
nand UO_67 (O_67,N_24830,N_24870);
or UO_68 (O_68,N_24982,N_24919);
xnor UO_69 (O_69,N_24843,N_24941);
xor UO_70 (O_70,N_24881,N_24828);
and UO_71 (O_71,N_24873,N_24880);
xnor UO_72 (O_72,N_24948,N_24966);
or UO_73 (O_73,N_24812,N_24846);
nor UO_74 (O_74,N_24804,N_24984);
or UO_75 (O_75,N_24902,N_24979);
nor UO_76 (O_76,N_24997,N_24823);
nor UO_77 (O_77,N_24965,N_24989);
and UO_78 (O_78,N_24860,N_24904);
xnor UO_79 (O_79,N_24862,N_24834);
and UO_80 (O_80,N_24974,N_24942);
nand UO_81 (O_81,N_24969,N_24936);
xnor UO_82 (O_82,N_24829,N_24943);
xnor UO_83 (O_83,N_24835,N_24939);
and UO_84 (O_84,N_24878,N_24923);
nand UO_85 (O_85,N_24954,N_24971);
and UO_86 (O_86,N_24838,N_24977);
nand UO_87 (O_87,N_24931,N_24825);
nor UO_88 (O_88,N_24874,N_24963);
and UO_89 (O_89,N_24872,N_24990);
xor UO_90 (O_90,N_24983,N_24994);
nand UO_91 (O_91,N_24896,N_24975);
or UO_92 (O_92,N_24899,N_24925);
and UO_93 (O_93,N_24852,N_24842);
nand UO_94 (O_94,N_24801,N_24859);
and UO_95 (O_95,N_24897,N_24947);
nand UO_96 (O_96,N_24926,N_24912);
or UO_97 (O_97,N_24841,N_24832);
or UO_98 (O_98,N_24886,N_24978);
nand UO_99 (O_99,N_24914,N_24924);
xor UO_100 (O_100,N_24817,N_24909);
xor UO_101 (O_101,N_24925,N_24982);
or UO_102 (O_102,N_24943,N_24852);
nand UO_103 (O_103,N_24837,N_24865);
xnor UO_104 (O_104,N_24873,N_24847);
or UO_105 (O_105,N_24924,N_24925);
and UO_106 (O_106,N_24933,N_24938);
xor UO_107 (O_107,N_24895,N_24997);
nor UO_108 (O_108,N_24947,N_24895);
nand UO_109 (O_109,N_24834,N_24819);
xor UO_110 (O_110,N_24848,N_24846);
nor UO_111 (O_111,N_24964,N_24889);
or UO_112 (O_112,N_24998,N_24853);
and UO_113 (O_113,N_24950,N_24989);
nor UO_114 (O_114,N_24921,N_24915);
or UO_115 (O_115,N_24961,N_24974);
xor UO_116 (O_116,N_24804,N_24921);
and UO_117 (O_117,N_24840,N_24819);
and UO_118 (O_118,N_24800,N_24948);
nand UO_119 (O_119,N_24852,N_24802);
and UO_120 (O_120,N_24943,N_24848);
nor UO_121 (O_121,N_24909,N_24993);
nand UO_122 (O_122,N_24833,N_24860);
nand UO_123 (O_123,N_24872,N_24913);
or UO_124 (O_124,N_24904,N_24896);
nor UO_125 (O_125,N_24919,N_24837);
nor UO_126 (O_126,N_24942,N_24989);
xor UO_127 (O_127,N_24805,N_24809);
nor UO_128 (O_128,N_24874,N_24825);
xor UO_129 (O_129,N_24877,N_24958);
and UO_130 (O_130,N_24930,N_24974);
or UO_131 (O_131,N_24942,N_24865);
nand UO_132 (O_132,N_24860,N_24971);
nor UO_133 (O_133,N_24979,N_24850);
and UO_134 (O_134,N_24937,N_24877);
or UO_135 (O_135,N_24845,N_24954);
and UO_136 (O_136,N_24958,N_24819);
and UO_137 (O_137,N_24970,N_24896);
xor UO_138 (O_138,N_24807,N_24963);
or UO_139 (O_139,N_24941,N_24927);
nand UO_140 (O_140,N_24816,N_24983);
xor UO_141 (O_141,N_24887,N_24960);
or UO_142 (O_142,N_24858,N_24910);
and UO_143 (O_143,N_24924,N_24801);
and UO_144 (O_144,N_24984,N_24835);
xor UO_145 (O_145,N_24858,N_24963);
and UO_146 (O_146,N_24911,N_24977);
nand UO_147 (O_147,N_24850,N_24970);
xor UO_148 (O_148,N_24944,N_24836);
or UO_149 (O_149,N_24992,N_24864);
nand UO_150 (O_150,N_24894,N_24911);
and UO_151 (O_151,N_24846,N_24816);
nor UO_152 (O_152,N_24930,N_24998);
xnor UO_153 (O_153,N_24980,N_24830);
nand UO_154 (O_154,N_24823,N_24866);
and UO_155 (O_155,N_24967,N_24900);
xor UO_156 (O_156,N_24910,N_24844);
and UO_157 (O_157,N_24913,N_24945);
xor UO_158 (O_158,N_24905,N_24896);
or UO_159 (O_159,N_24842,N_24940);
nor UO_160 (O_160,N_24947,N_24893);
xor UO_161 (O_161,N_24914,N_24944);
xnor UO_162 (O_162,N_24970,N_24809);
nor UO_163 (O_163,N_24942,N_24832);
nor UO_164 (O_164,N_24901,N_24838);
and UO_165 (O_165,N_24975,N_24951);
or UO_166 (O_166,N_24872,N_24901);
and UO_167 (O_167,N_24919,N_24904);
xnor UO_168 (O_168,N_24967,N_24955);
nor UO_169 (O_169,N_24996,N_24835);
nand UO_170 (O_170,N_24927,N_24841);
xnor UO_171 (O_171,N_24908,N_24974);
or UO_172 (O_172,N_24963,N_24888);
xor UO_173 (O_173,N_24979,N_24999);
or UO_174 (O_174,N_24853,N_24817);
or UO_175 (O_175,N_24802,N_24925);
and UO_176 (O_176,N_24928,N_24927);
nor UO_177 (O_177,N_24816,N_24874);
xnor UO_178 (O_178,N_24905,N_24880);
and UO_179 (O_179,N_24997,N_24964);
nand UO_180 (O_180,N_24890,N_24845);
or UO_181 (O_181,N_24871,N_24970);
and UO_182 (O_182,N_24932,N_24837);
or UO_183 (O_183,N_24903,N_24970);
nand UO_184 (O_184,N_24872,N_24845);
or UO_185 (O_185,N_24997,N_24913);
and UO_186 (O_186,N_24964,N_24966);
or UO_187 (O_187,N_24811,N_24869);
nor UO_188 (O_188,N_24846,N_24975);
nand UO_189 (O_189,N_24853,N_24897);
nor UO_190 (O_190,N_24939,N_24982);
xor UO_191 (O_191,N_24993,N_24914);
nand UO_192 (O_192,N_24970,N_24812);
nor UO_193 (O_193,N_24989,N_24812);
xor UO_194 (O_194,N_24996,N_24873);
xnor UO_195 (O_195,N_24964,N_24900);
nor UO_196 (O_196,N_24852,N_24904);
and UO_197 (O_197,N_24834,N_24878);
or UO_198 (O_198,N_24872,N_24849);
nand UO_199 (O_199,N_24876,N_24836);
and UO_200 (O_200,N_24830,N_24969);
and UO_201 (O_201,N_24832,N_24989);
xor UO_202 (O_202,N_24949,N_24858);
nor UO_203 (O_203,N_24857,N_24986);
xor UO_204 (O_204,N_24898,N_24877);
and UO_205 (O_205,N_24871,N_24981);
nor UO_206 (O_206,N_24916,N_24914);
and UO_207 (O_207,N_24854,N_24958);
and UO_208 (O_208,N_24926,N_24960);
nand UO_209 (O_209,N_24942,N_24895);
nor UO_210 (O_210,N_24938,N_24830);
and UO_211 (O_211,N_24977,N_24899);
nor UO_212 (O_212,N_24975,N_24947);
and UO_213 (O_213,N_24987,N_24915);
or UO_214 (O_214,N_24902,N_24827);
nand UO_215 (O_215,N_24892,N_24848);
and UO_216 (O_216,N_24879,N_24824);
xor UO_217 (O_217,N_24967,N_24849);
nor UO_218 (O_218,N_24800,N_24921);
xnor UO_219 (O_219,N_24933,N_24975);
xnor UO_220 (O_220,N_24817,N_24807);
and UO_221 (O_221,N_24887,N_24907);
nand UO_222 (O_222,N_24850,N_24927);
nand UO_223 (O_223,N_24927,N_24818);
or UO_224 (O_224,N_24840,N_24926);
nand UO_225 (O_225,N_24803,N_24973);
and UO_226 (O_226,N_24889,N_24830);
xor UO_227 (O_227,N_24966,N_24866);
xor UO_228 (O_228,N_24846,N_24956);
nor UO_229 (O_229,N_24882,N_24975);
nor UO_230 (O_230,N_24916,N_24843);
xnor UO_231 (O_231,N_24804,N_24947);
nor UO_232 (O_232,N_24833,N_24928);
and UO_233 (O_233,N_24918,N_24840);
nand UO_234 (O_234,N_24954,N_24914);
nor UO_235 (O_235,N_24947,N_24951);
nor UO_236 (O_236,N_24814,N_24880);
xnor UO_237 (O_237,N_24830,N_24845);
and UO_238 (O_238,N_24863,N_24803);
nor UO_239 (O_239,N_24935,N_24826);
and UO_240 (O_240,N_24809,N_24969);
nand UO_241 (O_241,N_24937,N_24878);
nand UO_242 (O_242,N_24928,N_24921);
xor UO_243 (O_243,N_24808,N_24972);
nand UO_244 (O_244,N_24933,N_24849);
nand UO_245 (O_245,N_24969,N_24928);
xor UO_246 (O_246,N_24958,N_24946);
nand UO_247 (O_247,N_24869,N_24982);
nand UO_248 (O_248,N_24931,N_24885);
nand UO_249 (O_249,N_24975,N_24903);
xnor UO_250 (O_250,N_24821,N_24864);
or UO_251 (O_251,N_24824,N_24814);
nand UO_252 (O_252,N_24942,N_24943);
nand UO_253 (O_253,N_24865,N_24958);
nor UO_254 (O_254,N_24961,N_24913);
and UO_255 (O_255,N_24987,N_24968);
or UO_256 (O_256,N_24908,N_24817);
or UO_257 (O_257,N_24941,N_24882);
or UO_258 (O_258,N_24985,N_24973);
and UO_259 (O_259,N_24946,N_24822);
and UO_260 (O_260,N_24836,N_24803);
xor UO_261 (O_261,N_24999,N_24869);
or UO_262 (O_262,N_24866,N_24967);
or UO_263 (O_263,N_24887,N_24888);
nor UO_264 (O_264,N_24858,N_24888);
nor UO_265 (O_265,N_24937,N_24858);
and UO_266 (O_266,N_24960,N_24892);
or UO_267 (O_267,N_24814,N_24914);
xor UO_268 (O_268,N_24914,N_24950);
nor UO_269 (O_269,N_24923,N_24966);
or UO_270 (O_270,N_24913,N_24943);
xor UO_271 (O_271,N_24886,N_24982);
and UO_272 (O_272,N_24893,N_24921);
and UO_273 (O_273,N_24954,N_24806);
or UO_274 (O_274,N_24879,N_24951);
and UO_275 (O_275,N_24847,N_24810);
nand UO_276 (O_276,N_24864,N_24843);
xor UO_277 (O_277,N_24805,N_24930);
and UO_278 (O_278,N_24952,N_24845);
and UO_279 (O_279,N_24892,N_24879);
or UO_280 (O_280,N_24858,N_24893);
and UO_281 (O_281,N_24820,N_24976);
or UO_282 (O_282,N_24966,N_24852);
and UO_283 (O_283,N_24825,N_24999);
xnor UO_284 (O_284,N_24805,N_24867);
xor UO_285 (O_285,N_24903,N_24824);
or UO_286 (O_286,N_24932,N_24944);
or UO_287 (O_287,N_24818,N_24982);
or UO_288 (O_288,N_24931,N_24937);
or UO_289 (O_289,N_24989,N_24839);
or UO_290 (O_290,N_24812,N_24937);
nor UO_291 (O_291,N_24979,N_24806);
nand UO_292 (O_292,N_24876,N_24801);
nor UO_293 (O_293,N_24882,N_24931);
nor UO_294 (O_294,N_24895,N_24925);
and UO_295 (O_295,N_24959,N_24853);
xor UO_296 (O_296,N_24956,N_24826);
nor UO_297 (O_297,N_24912,N_24805);
and UO_298 (O_298,N_24803,N_24852);
nand UO_299 (O_299,N_24941,N_24939);
xnor UO_300 (O_300,N_24915,N_24954);
or UO_301 (O_301,N_24940,N_24927);
xor UO_302 (O_302,N_24888,N_24974);
xor UO_303 (O_303,N_24856,N_24940);
nand UO_304 (O_304,N_24960,N_24953);
or UO_305 (O_305,N_24947,N_24838);
nand UO_306 (O_306,N_24898,N_24803);
nand UO_307 (O_307,N_24959,N_24814);
and UO_308 (O_308,N_24822,N_24834);
and UO_309 (O_309,N_24809,N_24939);
nand UO_310 (O_310,N_24956,N_24837);
nand UO_311 (O_311,N_24880,N_24817);
or UO_312 (O_312,N_24851,N_24824);
nor UO_313 (O_313,N_24937,N_24874);
or UO_314 (O_314,N_24905,N_24953);
xnor UO_315 (O_315,N_24852,N_24973);
nor UO_316 (O_316,N_24886,N_24941);
and UO_317 (O_317,N_24834,N_24818);
xor UO_318 (O_318,N_24965,N_24969);
or UO_319 (O_319,N_24860,N_24958);
or UO_320 (O_320,N_24857,N_24971);
nand UO_321 (O_321,N_24805,N_24933);
xnor UO_322 (O_322,N_24998,N_24958);
nand UO_323 (O_323,N_24814,N_24863);
nand UO_324 (O_324,N_24985,N_24948);
or UO_325 (O_325,N_24832,N_24817);
or UO_326 (O_326,N_24815,N_24986);
and UO_327 (O_327,N_24991,N_24999);
nor UO_328 (O_328,N_24810,N_24870);
and UO_329 (O_329,N_24841,N_24876);
xor UO_330 (O_330,N_24914,N_24965);
nor UO_331 (O_331,N_24925,N_24926);
and UO_332 (O_332,N_24882,N_24808);
nand UO_333 (O_333,N_24863,N_24950);
and UO_334 (O_334,N_24853,N_24863);
and UO_335 (O_335,N_24960,N_24937);
nor UO_336 (O_336,N_24994,N_24952);
or UO_337 (O_337,N_24868,N_24935);
xor UO_338 (O_338,N_24988,N_24880);
nand UO_339 (O_339,N_24880,N_24847);
or UO_340 (O_340,N_24995,N_24977);
nand UO_341 (O_341,N_24878,N_24983);
or UO_342 (O_342,N_24880,N_24888);
xor UO_343 (O_343,N_24985,N_24958);
nand UO_344 (O_344,N_24909,N_24801);
nor UO_345 (O_345,N_24934,N_24890);
nor UO_346 (O_346,N_24826,N_24947);
xnor UO_347 (O_347,N_24908,N_24880);
nor UO_348 (O_348,N_24838,N_24937);
and UO_349 (O_349,N_24867,N_24948);
nor UO_350 (O_350,N_24954,N_24961);
nand UO_351 (O_351,N_24948,N_24925);
nand UO_352 (O_352,N_24995,N_24910);
xnor UO_353 (O_353,N_24837,N_24812);
nor UO_354 (O_354,N_24973,N_24813);
and UO_355 (O_355,N_24873,N_24883);
nor UO_356 (O_356,N_24914,N_24939);
xnor UO_357 (O_357,N_24865,N_24983);
or UO_358 (O_358,N_24829,N_24865);
xor UO_359 (O_359,N_24908,N_24860);
xor UO_360 (O_360,N_24894,N_24980);
nor UO_361 (O_361,N_24928,N_24802);
or UO_362 (O_362,N_24922,N_24859);
nand UO_363 (O_363,N_24858,N_24869);
and UO_364 (O_364,N_24954,N_24903);
nand UO_365 (O_365,N_24973,N_24842);
xnor UO_366 (O_366,N_24883,N_24806);
and UO_367 (O_367,N_24871,N_24950);
or UO_368 (O_368,N_24822,N_24938);
and UO_369 (O_369,N_24928,N_24939);
xor UO_370 (O_370,N_24946,N_24806);
and UO_371 (O_371,N_24906,N_24913);
xnor UO_372 (O_372,N_24866,N_24855);
nand UO_373 (O_373,N_24816,N_24883);
xnor UO_374 (O_374,N_24988,N_24911);
xnor UO_375 (O_375,N_24991,N_24810);
xnor UO_376 (O_376,N_24925,N_24986);
nand UO_377 (O_377,N_24904,N_24917);
xor UO_378 (O_378,N_24813,N_24828);
nand UO_379 (O_379,N_24878,N_24976);
nand UO_380 (O_380,N_24819,N_24817);
xor UO_381 (O_381,N_24890,N_24973);
or UO_382 (O_382,N_24832,N_24825);
nor UO_383 (O_383,N_24828,N_24987);
or UO_384 (O_384,N_24971,N_24958);
nor UO_385 (O_385,N_24923,N_24982);
and UO_386 (O_386,N_24831,N_24907);
nor UO_387 (O_387,N_24899,N_24934);
nand UO_388 (O_388,N_24964,N_24923);
xnor UO_389 (O_389,N_24871,N_24938);
or UO_390 (O_390,N_24881,N_24906);
or UO_391 (O_391,N_24940,N_24981);
nand UO_392 (O_392,N_24945,N_24907);
nor UO_393 (O_393,N_24921,N_24960);
or UO_394 (O_394,N_24814,N_24968);
nor UO_395 (O_395,N_24848,N_24916);
nor UO_396 (O_396,N_24865,N_24948);
or UO_397 (O_397,N_24937,N_24933);
nor UO_398 (O_398,N_24936,N_24884);
and UO_399 (O_399,N_24957,N_24994);
xnor UO_400 (O_400,N_24808,N_24916);
nand UO_401 (O_401,N_24835,N_24967);
nand UO_402 (O_402,N_24901,N_24814);
nor UO_403 (O_403,N_24824,N_24931);
and UO_404 (O_404,N_24890,N_24965);
nor UO_405 (O_405,N_24935,N_24823);
and UO_406 (O_406,N_24961,N_24891);
or UO_407 (O_407,N_24880,N_24923);
xor UO_408 (O_408,N_24923,N_24895);
and UO_409 (O_409,N_24800,N_24883);
xor UO_410 (O_410,N_24894,N_24964);
xnor UO_411 (O_411,N_24871,N_24809);
and UO_412 (O_412,N_24964,N_24800);
and UO_413 (O_413,N_24989,N_24827);
xnor UO_414 (O_414,N_24949,N_24896);
and UO_415 (O_415,N_24805,N_24830);
xnor UO_416 (O_416,N_24835,N_24906);
xor UO_417 (O_417,N_24939,N_24980);
nand UO_418 (O_418,N_24873,N_24886);
nand UO_419 (O_419,N_24800,N_24829);
xor UO_420 (O_420,N_24858,N_24904);
nor UO_421 (O_421,N_24807,N_24950);
nor UO_422 (O_422,N_24885,N_24901);
nand UO_423 (O_423,N_24998,N_24978);
or UO_424 (O_424,N_24914,N_24899);
nor UO_425 (O_425,N_24841,N_24809);
nand UO_426 (O_426,N_24891,N_24967);
nor UO_427 (O_427,N_24970,N_24815);
and UO_428 (O_428,N_24984,N_24829);
nand UO_429 (O_429,N_24975,N_24875);
xor UO_430 (O_430,N_24830,N_24966);
nor UO_431 (O_431,N_24983,N_24918);
or UO_432 (O_432,N_24808,N_24840);
nand UO_433 (O_433,N_24971,N_24968);
or UO_434 (O_434,N_24959,N_24992);
nand UO_435 (O_435,N_24810,N_24883);
and UO_436 (O_436,N_24935,N_24981);
xor UO_437 (O_437,N_24862,N_24864);
and UO_438 (O_438,N_24811,N_24880);
nor UO_439 (O_439,N_24982,N_24819);
xnor UO_440 (O_440,N_24881,N_24999);
nand UO_441 (O_441,N_24921,N_24869);
and UO_442 (O_442,N_24978,N_24982);
nand UO_443 (O_443,N_24960,N_24988);
nand UO_444 (O_444,N_24859,N_24858);
nand UO_445 (O_445,N_24990,N_24825);
xor UO_446 (O_446,N_24922,N_24950);
xnor UO_447 (O_447,N_24908,N_24931);
or UO_448 (O_448,N_24830,N_24977);
nand UO_449 (O_449,N_24890,N_24944);
or UO_450 (O_450,N_24955,N_24982);
nand UO_451 (O_451,N_24972,N_24818);
nor UO_452 (O_452,N_24929,N_24805);
nor UO_453 (O_453,N_24808,N_24999);
or UO_454 (O_454,N_24987,N_24894);
or UO_455 (O_455,N_24912,N_24997);
and UO_456 (O_456,N_24800,N_24856);
xnor UO_457 (O_457,N_24915,N_24933);
nor UO_458 (O_458,N_24928,N_24856);
or UO_459 (O_459,N_24871,N_24812);
nand UO_460 (O_460,N_24931,N_24919);
nor UO_461 (O_461,N_24905,N_24976);
or UO_462 (O_462,N_24963,N_24832);
nor UO_463 (O_463,N_24956,N_24855);
and UO_464 (O_464,N_24967,N_24834);
or UO_465 (O_465,N_24970,N_24910);
and UO_466 (O_466,N_24835,N_24958);
nor UO_467 (O_467,N_24917,N_24998);
xor UO_468 (O_468,N_24882,N_24900);
xor UO_469 (O_469,N_24965,N_24995);
nor UO_470 (O_470,N_24937,N_24908);
or UO_471 (O_471,N_24845,N_24876);
and UO_472 (O_472,N_24990,N_24869);
or UO_473 (O_473,N_24928,N_24970);
or UO_474 (O_474,N_24987,N_24946);
nor UO_475 (O_475,N_24852,N_24902);
nand UO_476 (O_476,N_24908,N_24838);
and UO_477 (O_477,N_24850,N_24944);
xor UO_478 (O_478,N_24874,N_24883);
or UO_479 (O_479,N_24835,N_24855);
and UO_480 (O_480,N_24853,N_24937);
and UO_481 (O_481,N_24865,N_24915);
nand UO_482 (O_482,N_24846,N_24999);
or UO_483 (O_483,N_24867,N_24992);
and UO_484 (O_484,N_24962,N_24868);
and UO_485 (O_485,N_24990,N_24919);
or UO_486 (O_486,N_24999,N_24852);
nand UO_487 (O_487,N_24903,N_24969);
xor UO_488 (O_488,N_24886,N_24861);
nand UO_489 (O_489,N_24998,N_24913);
and UO_490 (O_490,N_24819,N_24802);
and UO_491 (O_491,N_24964,N_24929);
xnor UO_492 (O_492,N_24974,N_24911);
nor UO_493 (O_493,N_24867,N_24851);
nand UO_494 (O_494,N_24801,N_24835);
nand UO_495 (O_495,N_24851,N_24939);
nor UO_496 (O_496,N_24912,N_24987);
or UO_497 (O_497,N_24949,N_24876);
or UO_498 (O_498,N_24881,N_24998);
and UO_499 (O_499,N_24854,N_24997);
nor UO_500 (O_500,N_24888,N_24964);
nor UO_501 (O_501,N_24825,N_24963);
nand UO_502 (O_502,N_24865,N_24918);
or UO_503 (O_503,N_24953,N_24986);
and UO_504 (O_504,N_24837,N_24992);
nor UO_505 (O_505,N_24852,N_24858);
nor UO_506 (O_506,N_24996,N_24948);
nor UO_507 (O_507,N_24874,N_24951);
and UO_508 (O_508,N_24947,N_24923);
xor UO_509 (O_509,N_24970,N_24808);
or UO_510 (O_510,N_24879,N_24907);
and UO_511 (O_511,N_24946,N_24866);
nor UO_512 (O_512,N_24972,N_24951);
nor UO_513 (O_513,N_24980,N_24831);
or UO_514 (O_514,N_24948,N_24841);
nand UO_515 (O_515,N_24883,N_24951);
nand UO_516 (O_516,N_24873,N_24846);
or UO_517 (O_517,N_24884,N_24873);
nor UO_518 (O_518,N_24853,N_24924);
and UO_519 (O_519,N_24881,N_24924);
nor UO_520 (O_520,N_24897,N_24883);
nand UO_521 (O_521,N_24858,N_24867);
and UO_522 (O_522,N_24921,N_24832);
nand UO_523 (O_523,N_24850,N_24973);
nand UO_524 (O_524,N_24917,N_24922);
nor UO_525 (O_525,N_24880,N_24985);
nor UO_526 (O_526,N_24852,N_24872);
nor UO_527 (O_527,N_24987,N_24997);
and UO_528 (O_528,N_24902,N_24861);
xor UO_529 (O_529,N_24809,N_24940);
nand UO_530 (O_530,N_24810,N_24999);
nor UO_531 (O_531,N_24881,N_24870);
nand UO_532 (O_532,N_24934,N_24872);
nand UO_533 (O_533,N_24912,N_24949);
nor UO_534 (O_534,N_24946,N_24844);
xor UO_535 (O_535,N_24832,N_24801);
nor UO_536 (O_536,N_24882,N_24811);
xnor UO_537 (O_537,N_24815,N_24930);
xor UO_538 (O_538,N_24977,N_24945);
nand UO_539 (O_539,N_24932,N_24982);
xnor UO_540 (O_540,N_24838,N_24952);
or UO_541 (O_541,N_24934,N_24978);
nand UO_542 (O_542,N_24999,N_24948);
nor UO_543 (O_543,N_24876,N_24941);
nor UO_544 (O_544,N_24996,N_24923);
nor UO_545 (O_545,N_24995,N_24853);
xnor UO_546 (O_546,N_24812,N_24967);
or UO_547 (O_547,N_24800,N_24989);
nor UO_548 (O_548,N_24852,N_24971);
nand UO_549 (O_549,N_24944,N_24830);
and UO_550 (O_550,N_24956,N_24912);
or UO_551 (O_551,N_24842,N_24863);
nor UO_552 (O_552,N_24874,N_24976);
or UO_553 (O_553,N_24898,N_24869);
nand UO_554 (O_554,N_24990,N_24833);
xor UO_555 (O_555,N_24920,N_24965);
xnor UO_556 (O_556,N_24922,N_24951);
or UO_557 (O_557,N_24896,N_24943);
and UO_558 (O_558,N_24963,N_24877);
nor UO_559 (O_559,N_24829,N_24980);
nand UO_560 (O_560,N_24812,N_24819);
or UO_561 (O_561,N_24855,N_24939);
xor UO_562 (O_562,N_24916,N_24834);
and UO_563 (O_563,N_24935,N_24969);
and UO_564 (O_564,N_24823,N_24835);
or UO_565 (O_565,N_24980,N_24871);
xor UO_566 (O_566,N_24800,N_24838);
xnor UO_567 (O_567,N_24994,N_24944);
nand UO_568 (O_568,N_24868,N_24938);
xor UO_569 (O_569,N_24997,N_24903);
xnor UO_570 (O_570,N_24961,N_24827);
and UO_571 (O_571,N_24822,N_24887);
nand UO_572 (O_572,N_24843,N_24955);
xor UO_573 (O_573,N_24807,N_24826);
xor UO_574 (O_574,N_24930,N_24842);
or UO_575 (O_575,N_24865,N_24823);
xor UO_576 (O_576,N_24891,N_24902);
nor UO_577 (O_577,N_24962,N_24892);
nand UO_578 (O_578,N_24905,N_24988);
nand UO_579 (O_579,N_24870,N_24979);
and UO_580 (O_580,N_24886,N_24840);
and UO_581 (O_581,N_24803,N_24955);
nor UO_582 (O_582,N_24945,N_24899);
xor UO_583 (O_583,N_24953,N_24828);
or UO_584 (O_584,N_24964,N_24844);
or UO_585 (O_585,N_24861,N_24806);
and UO_586 (O_586,N_24842,N_24857);
nor UO_587 (O_587,N_24801,N_24936);
or UO_588 (O_588,N_24967,N_24872);
xnor UO_589 (O_589,N_24850,N_24843);
and UO_590 (O_590,N_24928,N_24895);
xnor UO_591 (O_591,N_24870,N_24922);
nor UO_592 (O_592,N_24914,N_24870);
nand UO_593 (O_593,N_24924,N_24986);
or UO_594 (O_594,N_24967,N_24991);
nor UO_595 (O_595,N_24994,N_24982);
and UO_596 (O_596,N_24914,N_24961);
xor UO_597 (O_597,N_24937,N_24965);
xor UO_598 (O_598,N_24905,N_24924);
nor UO_599 (O_599,N_24997,N_24955);
and UO_600 (O_600,N_24826,N_24958);
nand UO_601 (O_601,N_24933,N_24821);
and UO_602 (O_602,N_24800,N_24988);
nor UO_603 (O_603,N_24942,N_24970);
and UO_604 (O_604,N_24812,N_24800);
or UO_605 (O_605,N_24852,N_24982);
and UO_606 (O_606,N_24895,N_24820);
or UO_607 (O_607,N_24819,N_24995);
nand UO_608 (O_608,N_24921,N_24890);
and UO_609 (O_609,N_24978,N_24893);
nor UO_610 (O_610,N_24927,N_24901);
nand UO_611 (O_611,N_24969,N_24944);
xnor UO_612 (O_612,N_24839,N_24914);
and UO_613 (O_613,N_24924,N_24813);
or UO_614 (O_614,N_24839,N_24843);
and UO_615 (O_615,N_24888,N_24939);
nor UO_616 (O_616,N_24899,N_24820);
xor UO_617 (O_617,N_24864,N_24932);
nand UO_618 (O_618,N_24824,N_24967);
nor UO_619 (O_619,N_24894,N_24856);
nand UO_620 (O_620,N_24968,N_24863);
nor UO_621 (O_621,N_24949,N_24833);
or UO_622 (O_622,N_24807,N_24927);
or UO_623 (O_623,N_24896,N_24844);
or UO_624 (O_624,N_24991,N_24821);
nand UO_625 (O_625,N_24843,N_24963);
xnor UO_626 (O_626,N_24931,N_24987);
and UO_627 (O_627,N_24984,N_24827);
xnor UO_628 (O_628,N_24881,N_24907);
nor UO_629 (O_629,N_24935,N_24873);
nand UO_630 (O_630,N_24933,N_24850);
nor UO_631 (O_631,N_24821,N_24873);
and UO_632 (O_632,N_24916,N_24894);
and UO_633 (O_633,N_24812,N_24824);
xor UO_634 (O_634,N_24828,N_24864);
and UO_635 (O_635,N_24906,N_24849);
and UO_636 (O_636,N_24919,N_24897);
and UO_637 (O_637,N_24906,N_24837);
and UO_638 (O_638,N_24978,N_24898);
nand UO_639 (O_639,N_24938,N_24894);
nor UO_640 (O_640,N_24830,N_24957);
and UO_641 (O_641,N_24821,N_24965);
or UO_642 (O_642,N_24837,N_24896);
and UO_643 (O_643,N_24883,N_24860);
and UO_644 (O_644,N_24800,N_24885);
and UO_645 (O_645,N_24961,N_24919);
or UO_646 (O_646,N_24827,N_24877);
xnor UO_647 (O_647,N_24933,N_24998);
xor UO_648 (O_648,N_24914,N_24800);
nand UO_649 (O_649,N_24847,N_24869);
or UO_650 (O_650,N_24971,N_24949);
xor UO_651 (O_651,N_24940,N_24910);
or UO_652 (O_652,N_24965,N_24990);
xor UO_653 (O_653,N_24909,N_24882);
and UO_654 (O_654,N_24800,N_24875);
and UO_655 (O_655,N_24934,N_24915);
or UO_656 (O_656,N_24939,N_24834);
nor UO_657 (O_657,N_24965,N_24806);
nand UO_658 (O_658,N_24940,N_24872);
nor UO_659 (O_659,N_24930,N_24868);
or UO_660 (O_660,N_24989,N_24818);
nor UO_661 (O_661,N_24859,N_24827);
and UO_662 (O_662,N_24897,N_24962);
and UO_663 (O_663,N_24816,N_24991);
nand UO_664 (O_664,N_24921,N_24937);
nor UO_665 (O_665,N_24867,N_24935);
xor UO_666 (O_666,N_24946,N_24964);
xnor UO_667 (O_667,N_24864,N_24917);
xnor UO_668 (O_668,N_24831,N_24932);
and UO_669 (O_669,N_24997,N_24861);
nand UO_670 (O_670,N_24879,N_24957);
or UO_671 (O_671,N_24961,N_24902);
or UO_672 (O_672,N_24813,N_24835);
nand UO_673 (O_673,N_24988,N_24886);
and UO_674 (O_674,N_24808,N_24887);
nand UO_675 (O_675,N_24948,N_24878);
nor UO_676 (O_676,N_24953,N_24989);
and UO_677 (O_677,N_24845,N_24885);
or UO_678 (O_678,N_24878,N_24859);
nand UO_679 (O_679,N_24824,N_24929);
nand UO_680 (O_680,N_24932,N_24851);
xor UO_681 (O_681,N_24996,N_24974);
xor UO_682 (O_682,N_24954,N_24844);
nor UO_683 (O_683,N_24978,N_24952);
xnor UO_684 (O_684,N_24978,N_24806);
and UO_685 (O_685,N_24821,N_24861);
nand UO_686 (O_686,N_24895,N_24962);
nor UO_687 (O_687,N_24886,N_24998);
nor UO_688 (O_688,N_24981,N_24827);
nand UO_689 (O_689,N_24850,N_24975);
nand UO_690 (O_690,N_24867,N_24826);
nand UO_691 (O_691,N_24861,N_24942);
and UO_692 (O_692,N_24873,N_24986);
nand UO_693 (O_693,N_24838,N_24807);
nand UO_694 (O_694,N_24945,N_24904);
and UO_695 (O_695,N_24937,N_24995);
nor UO_696 (O_696,N_24923,N_24867);
nand UO_697 (O_697,N_24847,N_24966);
or UO_698 (O_698,N_24809,N_24886);
xnor UO_699 (O_699,N_24975,N_24864);
and UO_700 (O_700,N_24875,N_24866);
nand UO_701 (O_701,N_24902,N_24873);
nor UO_702 (O_702,N_24810,N_24854);
nor UO_703 (O_703,N_24890,N_24802);
or UO_704 (O_704,N_24969,N_24882);
or UO_705 (O_705,N_24917,N_24894);
xnor UO_706 (O_706,N_24906,N_24859);
or UO_707 (O_707,N_24824,N_24822);
nand UO_708 (O_708,N_24846,N_24810);
nand UO_709 (O_709,N_24925,N_24865);
and UO_710 (O_710,N_24883,N_24915);
and UO_711 (O_711,N_24995,N_24956);
nor UO_712 (O_712,N_24924,N_24958);
xnor UO_713 (O_713,N_24840,N_24967);
nand UO_714 (O_714,N_24936,N_24971);
nor UO_715 (O_715,N_24950,N_24975);
nand UO_716 (O_716,N_24956,N_24946);
or UO_717 (O_717,N_24846,N_24940);
and UO_718 (O_718,N_24987,N_24933);
nand UO_719 (O_719,N_24987,N_24852);
nor UO_720 (O_720,N_24973,N_24986);
nor UO_721 (O_721,N_24811,N_24946);
or UO_722 (O_722,N_24918,N_24932);
or UO_723 (O_723,N_24822,N_24927);
or UO_724 (O_724,N_24845,N_24802);
or UO_725 (O_725,N_24908,N_24962);
nand UO_726 (O_726,N_24973,N_24805);
xor UO_727 (O_727,N_24999,N_24824);
xnor UO_728 (O_728,N_24855,N_24905);
and UO_729 (O_729,N_24815,N_24828);
and UO_730 (O_730,N_24888,N_24896);
nor UO_731 (O_731,N_24976,N_24892);
nor UO_732 (O_732,N_24969,N_24927);
and UO_733 (O_733,N_24903,N_24923);
xor UO_734 (O_734,N_24903,N_24816);
nor UO_735 (O_735,N_24979,N_24853);
xnor UO_736 (O_736,N_24827,N_24906);
nor UO_737 (O_737,N_24879,N_24963);
and UO_738 (O_738,N_24851,N_24888);
nand UO_739 (O_739,N_24818,N_24884);
nor UO_740 (O_740,N_24838,N_24900);
and UO_741 (O_741,N_24956,N_24869);
xor UO_742 (O_742,N_24919,N_24949);
or UO_743 (O_743,N_24848,N_24861);
xor UO_744 (O_744,N_24937,N_24811);
nor UO_745 (O_745,N_24854,N_24862);
or UO_746 (O_746,N_24969,N_24976);
xnor UO_747 (O_747,N_24831,N_24950);
or UO_748 (O_748,N_24876,N_24844);
nand UO_749 (O_749,N_24869,N_24835);
or UO_750 (O_750,N_24803,N_24967);
xnor UO_751 (O_751,N_24990,N_24937);
nand UO_752 (O_752,N_24949,N_24993);
nand UO_753 (O_753,N_24854,N_24953);
xor UO_754 (O_754,N_24878,N_24902);
xor UO_755 (O_755,N_24834,N_24855);
or UO_756 (O_756,N_24969,N_24847);
and UO_757 (O_757,N_24921,N_24973);
nor UO_758 (O_758,N_24974,N_24824);
nor UO_759 (O_759,N_24979,N_24958);
nor UO_760 (O_760,N_24810,N_24804);
nand UO_761 (O_761,N_24845,N_24976);
nand UO_762 (O_762,N_24931,N_24821);
nor UO_763 (O_763,N_24855,N_24854);
nor UO_764 (O_764,N_24887,N_24903);
and UO_765 (O_765,N_24871,N_24860);
nor UO_766 (O_766,N_24925,N_24989);
nand UO_767 (O_767,N_24886,N_24858);
nand UO_768 (O_768,N_24873,N_24874);
nor UO_769 (O_769,N_24863,N_24927);
or UO_770 (O_770,N_24862,N_24850);
xnor UO_771 (O_771,N_24997,N_24935);
and UO_772 (O_772,N_24951,N_24819);
and UO_773 (O_773,N_24981,N_24992);
nand UO_774 (O_774,N_24994,N_24822);
xor UO_775 (O_775,N_24985,N_24978);
nor UO_776 (O_776,N_24878,N_24855);
nor UO_777 (O_777,N_24823,N_24948);
and UO_778 (O_778,N_24841,N_24814);
or UO_779 (O_779,N_24961,N_24872);
nand UO_780 (O_780,N_24971,N_24923);
xor UO_781 (O_781,N_24858,N_24814);
xor UO_782 (O_782,N_24834,N_24952);
xor UO_783 (O_783,N_24958,N_24896);
nor UO_784 (O_784,N_24936,N_24999);
nand UO_785 (O_785,N_24946,N_24863);
nor UO_786 (O_786,N_24835,N_24824);
xnor UO_787 (O_787,N_24994,N_24844);
or UO_788 (O_788,N_24957,N_24978);
nor UO_789 (O_789,N_24838,N_24874);
nor UO_790 (O_790,N_24850,N_24971);
xor UO_791 (O_791,N_24903,N_24935);
nor UO_792 (O_792,N_24839,N_24968);
nand UO_793 (O_793,N_24886,N_24947);
nor UO_794 (O_794,N_24877,N_24962);
xnor UO_795 (O_795,N_24867,N_24976);
and UO_796 (O_796,N_24839,N_24997);
nor UO_797 (O_797,N_24989,N_24918);
xnor UO_798 (O_798,N_24834,N_24807);
and UO_799 (O_799,N_24873,N_24829);
or UO_800 (O_800,N_24861,N_24973);
nor UO_801 (O_801,N_24924,N_24875);
nor UO_802 (O_802,N_24989,N_24901);
nor UO_803 (O_803,N_24914,N_24836);
or UO_804 (O_804,N_24937,N_24930);
and UO_805 (O_805,N_24979,N_24867);
or UO_806 (O_806,N_24976,N_24881);
nor UO_807 (O_807,N_24966,N_24986);
nand UO_808 (O_808,N_24907,N_24925);
and UO_809 (O_809,N_24822,N_24965);
or UO_810 (O_810,N_24812,N_24938);
or UO_811 (O_811,N_24823,N_24907);
xnor UO_812 (O_812,N_24978,N_24958);
nor UO_813 (O_813,N_24811,N_24870);
or UO_814 (O_814,N_24894,N_24988);
xnor UO_815 (O_815,N_24950,N_24852);
xor UO_816 (O_816,N_24894,N_24816);
or UO_817 (O_817,N_24815,N_24918);
nor UO_818 (O_818,N_24978,N_24895);
nand UO_819 (O_819,N_24988,N_24906);
or UO_820 (O_820,N_24981,N_24879);
and UO_821 (O_821,N_24833,N_24877);
nand UO_822 (O_822,N_24908,N_24911);
nor UO_823 (O_823,N_24831,N_24822);
xnor UO_824 (O_824,N_24877,N_24832);
xor UO_825 (O_825,N_24828,N_24997);
nor UO_826 (O_826,N_24961,N_24983);
and UO_827 (O_827,N_24886,N_24935);
nand UO_828 (O_828,N_24905,N_24967);
and UO_829 (O_829,N_24986,N_24931);
nor UO_830 (O_830,N_24846,N_24817);
nor UO_831 (O_831,N_24987,N_24803);
or UO_832 (O_832,N_24884,N_24922);
nor UO_833 (O_833,N_24887,N_24989);
nand UO_834 (O_834,N_24997,N_24953);
nor UO_835 (O_835,N_24821,N_24894);
or UO_836 (O_836,N_24832,N_24835);
and UO_837 (O_837,N_24807,N_24876);
nor UO_838 (O_838,N_24945,N_24893);
nand UO_839 (O_839,N_24926,N_24859);
xor UO_840 (O_840,N_24813,N_24802);
and UO_841 (O_841,N_24839,N_24928);
nor UO_842 (O_842,N_24948,N_24853);
xor UO_843 (O_843,N_24976,N_24839);
and UO_844 (O_844,N_24964,N_24867);
or UO_845 (O_845,N_24927,N_24821);
nand UO_846 (O_846,N_24869,N_24834);
nor UO_847 (O_847,N_24854,N_24893);
nand UO_848 (O_848,N_24812,N_24856);
nand UO_849 (O_849,N_24853,N_24907);
and UO_850 (O_850,N_24888,N_24885);
or UO_851 (O_851,N_24951,N_24851);
nor UO_852 (O_852,N_24878,N_24935);
xnor UO_853 (O_853,N_24836,N_24911);
and UO_854 (O_854,N_24865,N_24831);
or UO_855 (O_855,N_24894,N_24822);
or UO_856 (O_856,N_24820,N_24993);
nor UO_857 (O_857,N_24928,N_24949);
or UO_858 (O_858,N_24895,N_24800);
nor UO_859 (O_859,N_24906,N_24890);
or UO_860 (O_860,N_24952,N_24933);
xor UO_861 (O_861,N_24903,N_24886);
or UO_862 (O_862,N_24961,N_24979);
nand UO_863 (O_863,N_24902,N_24955);
or UO_864 (O_864,N_24849,N_24962);
or UO_865 (O_865,N_24876,N_24808);
or UO_866 (O_866,N_24920,N_24948);
or UO_867 (O_867,N_24905,N_24874);
xnor UO_868 (O_868,N_24985,N_24918);
nand UO_869 (O_869,N_24818,N_24855);
nand UO_870 (O_870,N_24880,N_24881);
or UO_871 (O_871,N_24970,N_24847);
nor UO_872 (O_872,N_24805,N_24883);
nor UO_873 (O_873,N_24911,N_24859);
and UO_874 (O_874,N_24847,N_24953);
nand UO_875 (O_875,N_24872,N_24802);
nand UO_876 (O_876,N_24891,N_24839);
xor UO_877 (O_877,N_24962,N_24980);
nor UO_878 (O_878,N_24871,N_24806);
and UO_879 (O_879,N_24975,N_24831);
nand UO_880 (O_880,N_24909,N_24862);
nand UO_881 (O_881,N_24841,N_24807);
and UO_882 (O_882,N_24998,N_24941);
nor UO_883 (O_883,N_24970,N_24930);
nor UO_884 (O_884,N_24816,N_24831);
xnor UO_885 (O_885,N_24929,N_24815);
or UO_886 (O_886,N_24954,N_24864);
or UO_887 (O_887,N_24908,N_24832);
xor UO_888 (O_888,N_24969,N_24820);
and UO_889 (O_889,N_24837,N_24960);
xor UO_890 (O_890,N_24869,N_24897);
nand UO_891 (O_891,N_24875,N_24978);
nor UO_892 (O_892,N_24941,N_24989);
and UO_893 (O_893,N_24860,N_24891);
nor UO_894 (O_894,N_24801,N_24882);
xor UO_895 (O_895,N_24985,N_24901);
nor UO_896 (O_896,N_24992,N_24853);
nand UO_897 (O_897,N_24859,N_24925);
nor UO_898 (O_898,N_24953,N_24860);
xor UO_899 (O_899,N_24820,N_24980);
or UO_900 (O_900,N_24842,N_24996);
nor UO_901 (O_901,N_24820,N_24852);
nand UO_902 (O_902,N_24896,N_24974);
xor UO_903 (O_903,N_24933,N_24969);
xnor UO_904 (O_904,N_24983,N_24839);
and UO_905 (O_905,N_24979,N_24845);
nor UO_906 (O_906,N_24936,N_24994);
or UO_907 (O_907,N_24984,N_24840);
nor UO_908 (O_908,N_24848,N_24922);
nand UO_909 (O_909,N_24977,N_24935);
nand UO_910 (O_910,N_24970,N_24887);
and UO_911 (O_911,N_24810,N_24844);
xor UO_912 (O_912,N_24831,N_24876);
or UO_913 (O_913,N_24930,N_24862);
and UO_914 (O_914,N_24962,N_24800);
nand UO_915 (O_915,N_24977,N_24941);
and UO_916 (O_916,N_24877,N_24906);
xnor UO_917 (O_917,N_24885,N_24918);
xor UO_918 (O_918,N_24808,N_24971);
or UO_919 (O_919,N_24831,N_24941);
nand UO_920 (O_920,N_24843,N_24814);
nor UO_921 (O_921,N_24995,N_24881);
nand UO_922 (O_922,N_24951,N_24856);
and UO_923 (O_923,N_24917,N_24851);
nand UO_924 (O_924,N_24936,N_24807);
or UO_925 (O_925,N_24887,N_24949);
and UO_926 (O_926,N_24987,N_24883);
nor UO_927 (O_927,N_24923,N_24884);
nor UO_928 (O_928,N_24849,N_24850);
or UO_929 (O_929,N_24996,N_24987);
nor UO_930 (O_930,N_24837,N_24815);
nand UO_931 (O_931,N_24834,N_24963);
or UO_932 (O_932,N_24876,N_24934);
and UO_933 (O_933,N_24900,N_24911);
and UO_934 (O_934,N_24869,N_24807);
and UO_935 (O_935,N_24957,N_24897);
nand UO_936 (O_936,N_24891,N_24898);
or UO_937 (O_937,N_24987,N_24979);
nand UO_938 (O_938,N_24974,N_24956);
nor UO_939 (O_939,N_24839,N_24880);
xnor UO_940 (O_940,N_24961,N_24949);
xnor UO_941 (O_941,N_24838,N_24916);
and UO_942 (O_942,N_24822,N_24990);
and UO_943 (O_943,N_24959,N_24801);
and UO_944 (O_944,N_24827,N_24820);
and UO_945 (O_945,N_24909,N_24913);
and UO_946 (O_946,N_24943,N_24903);
and UO_947 (O_947,N_24995,N_24870);
nand UO_948 (O_948,N_24803,N_24827);
xor UO_949 (O_949,N_24865,N_24855);
xnor UO_950 (O_950,N_24891,N_24955);
nand UO_951 (O_951,N_24892,N_24990);
nand UO_952 (O_952,N_24823,N_24943);
nand UO_953 (O_953,N_24829,N_24936);
nor UO_954 (O_954,N_24940,N_24851);
nand UO_955 (O_955,N_24934,N_24819);
nor UO_956 (O_956,N_24881,N_24927);
xnor UO_957 (O_957,N_24822,N_24839);
or UO_958 (O_958,N_24864,N_24942);
or UO_959 (O_959,N_24985,N_24944);
or UO_960 (O_960,N_24896,N_24845);
nand UO_961 (O_961,N_24943,N_24955);
or UO_962 (O_962,N_24871,N_24887);
or UO_963 (O_963,N_24966,N_24819);
xnor UO_964 (O_964,N_24915,N_24863);
xor UO_965 (O_965,N_24810,N_24834);
and UO_966 (O_966,N_24822,N_24966);
nand UO_967 (O_967,N_24966,N_24875);
nand UO_968 (O_968,N_24868,N_24915);
nor UO_969 (O_969,N_24828,N_24903);
nor UO_970 (O_970,N_24927,N_24906);
or UO_971 (O_971,N_24822,N_24910);
nand UO_972 (O_972,N_24912,N_24981);
or UO_973 (O_973,N_24845,N_24957);
or UO_974 (O_974,N_24894,N_24873);
xnor UO_975 (O_975,N_24860,N_24966);
nor UO_976 (O_976,N_24867,N_24959);
or UO_977 (O_977,N_24905,N_24968);
or UO_978 (O_978,N_24809,N_24965);
nor UO_979 (O_979,N_24814,N_24966);
xor UO_980 (O_980,N_24907,N_24821);
nor UO_981 (O_981,N_24835,N_24838);
nor UO_982 (O_982,N_24959,N_24805);
xnor UO_983 (O_983,N_24829,N_24878);
nand UO_984 (O_984,N_24931,N_24925);
nor UO_985 (O_985,N_24942,N_24874);
and UO_986 (O_986,N_24816,N_24810);
or UO_987 (O_987,N_24877,N_24965);
xor UO_988 (O_988,N_24813,N_24872);
nor UO_989 (O_989,N_24987,N_24938);
and UO_990 (O_990,N_24989,N_24848);
and UO_991 (O_991,N_24840,N_24864);
nor UO_992 (O_992,N_24972,N_24829);
xnor UO_993 (O_993,N_24980,N_24996);
or UO_994 (O_994,N_24878,N_24932);
or UO_995 (O_995,N_24873,N_24910);
nor UO_996 (O_996,N_24980,N_24834);
and UO_997 (O_997,N_24988,N_24902);
nand UO_998 (O_998,N_24946,N_24800);
nor UO_999 (O_999,N_24809,N_24834);
nor UO_1000 (O_1000,N_24950,N_24806);
nand UO_1001 (O_1001,N_24972,N_24876);
or UO_1002 (O_1002,N_24973,N_24812);
or UO_1003 (O_1003,N_24873,N_24921);
xnor UO_1004 (O_1004,N_24909,N_24979);
nor UO_1005 (O_1005,N_24850,N_24818);
nand UO_1006 (O_1006,N_24975,N_24948);
xor UO_1007 (O_1007,N_24985,N_24825);
nor UO_1008 (O_1008,N_24909,N_24899);
and UO_1009 (O_1009,N_24961,N_24924);
xor UO_1010 (O_1010,N_24828,N_24851);
or UO_1011 (O_1011,N_24972,N_24952);
and UO_1012 (O_1012,N_24821,N_24831);
nand UO_1013 (O_1013,N_24864,N_24836);
nor UO_1014 (O_1014,N_24936,N_24854);
nand UO_1015 (O_1015,N_24836,N_24908);
nor UO_1016 (O_1016,N_24832,N_24909);
or UO_1017 (O_1017,N_24967,N_24877);
nor UO_1018 (O_1018,N_24942,N_24828);
or UO_1019 (O_1019,N_24857,N_24913);
or UO_1020 (O_1020,N_24846,N_24927);
xnor UO_1021 (O_1021,N_24966,N_24962);
nand UO_1022 (O_1022,N_24968,N_24929);
xnor UO_1023 (O_1023,N_24931,N_24886);
nand UO_1024 (O_1024,N_24931,N_24927);
or UO_1025 (O_1025,N_24800,N_24959);
or UO_1026 (O_1026,N_24998,N_24962);
nand UO_1027 (O_1027,N_24870,N_24809);
nor UO_1028 (O_1028,N_24850,N_24822);
and UO_1029 (O_1029,N_24831,N_24810);
or UO_1030 (O_1030,N_24967,N_24831);
nor UO_1031 (O_1031,N_24844,N_24966);
and UO_1032 (O_1032,N_24940,N_24831);
or UO_1033 (O_1033,N_24946,N_24945);
nand UO_1034 (O_1034,N_24841,N_24894);
and UO_1035 (O_1035,N_24847,N_24818);
nand UO_1036 (O_1036,N_24876,N_24962);
xor UO_1037 (O_1037,N_24947,N_24918);
nor UO_1038 (O_1038,N_24821,N_24804);
and UO_1039 (O_1039,N_24855,N_24930);
and UO_1040 (O_1040,N_24854,N_24946);
or UO_1041 (O_1041,N_24900,N_24971);
or UO_1042 (O_1042,N_24976,N_24865);
nor UO_1043 (O_1043,N_24848,N_24824);
or UO_1044 (O_1044,N_24976,N_24956);
or UO_1045 (O_1045,N_24836,N_24852);
and UO_1046 (O_1046,N_24906,N_24955);
and UO_1047 (O_1047,N_24848,N_24857);
nand UO_1048 (O_1048,N_24819,N_24823);
nand UO_1049 (O_1049,N_24856,N_24882);
nor UO_1050 (O_1050,N_24926,N_24858);
or UO_1051 (O_1051,N_24943,N_24889);
and UO_1052 (O_1052,N_24819,N_24820);
and UO_1053 (O_1053,N_24976,N_24829);
xor UO_1054 (O_1054,N_24931,N_24819);
xor UO_1055 (O_1055,N_24866,N_24963);
and UO_1056 (O_1056,N_24989,N_24838);
and UO_1057 (O_1057,N_24867,N_24924);
xor UO_1058 (O_1058,N_24844,N_24939);
nor UO_1059 (O_1059,N_24803,N_24892);
and UO_1060 (O_1060,N_24867,N_24943);
or UO_1061 (O_1061,N_24871,N_24919);
or UO_1062 (O_1062,N_24912,N_24948);
and UO_1063 (O_1063,N_24895,N_24880);
nor UO_1064 (O_1064,N_24841,N_24871);
xor UO_1065 (O_1065,N_24959,N_24822);
or UO_1066 (O_1066,N_24956,N_24822);
or UO_1067 (O_1067,N_24906,N_24844);
xnor UO_1068 (O_1068,N_24918,N_24806);
xor UO_1069 (O_1069,N_24963,N_24945);
xnor UO_1070 (O_1070,N_24818,N_24904);
nor UO_1071 (O_1071,N_24816,N_24818);
nand UO_1072 (O_1072,N_24829,N_24811);
and UO_1073 (O_1073,N_24887,N_24807);
and UO_1074 (O_1074,N_24939,N_24821);
nand UO_1075 (O_1075,N_24951,N_24989);
nor UO_1076 (O_1076,N_24949,N_24832);
nand UO_1077 (O_1077,N_24982,N_24879);
nand UO_1078 (O_1078,N_24941,N_24853);
nor UO_1079 (O_1079,N_24909,N_24947);
xnor UO_1080 (O_1080,N_24803,N_24882);
and UO_1081 (O_1081,N_24853,N_24896);
nand UO_1082 (O_1082,N_24905,N_24828);
xnor UO_1083 (O_1083,N_24853,N_24947);
and UO_1084 (O_1084,N_24872,N_24949);
xor UO_1085 (O_1085,N_24882,N_24807);
nor UO_1086 (O_1086,N_24862,N_24878);
nand UO_1087 (O_1087,N_24904,N_24806);
nand UO_1088 (O_1088,N_24996,N_24807);
xnor UO_1089 (O_1089,N_24827,N_24911);
nand UO_1090 (O_1090,N_24850,N_24926);
nand UO_1091 (O_1091,N_24994,N_24825);
nand UO_1092 (O_1092,N_24811,N_24905);
and UO_1093 (O_1093,N_24986,N_24926);
or UO_1094 (O_1094,N_24969,N_24800);
nand UO_1095 (O_1095,N_24877,N_24969);
and UO_1096 (O_1096,N_24916,N_24897);
or UO_1097 (O_1097,N_24918,N_24970);
nor UO_1098 (O_1098,N_24854,N_24878);
nor UO_1099 (O_1099,N_24850,N_24828);
xnor UO_1100 (O_1100,N_24999,N_24967);
or UO_1101 (O_1101,N_24880,N_24921);
or UO_1102 (O_1102,N_24925,N_24881);
or UO_1103 (O_1103,N_24829,N_24957);
xor UO_1104 (O_1104,N_24885,N_24903);
and UO_1105 (O_1105,N_24880,N_24837);
nand UO_1106 (O_1106,N_24924,N_24959);
nand UO_1107 (O_1107,N_24952,N_24935);
and UO_1108 (O_1108,N_24978,N_24882);
and UO_1109 (O_1109,N_24805,N_24823);
nand UO_1110 (O_1110,N_24820,N_24822);
nor UO_1111 (O_1111,N_24923,N_24856);
nor UO_1112 (O_1112,N_24943,N_24915);
xnor UO_1113 (O_1113,N_24957,N_24801);
nor UO_1114 (O_1114,N_24820,N_24808);
xnor UO_1115 (O_1115,N_24826,N_24814);
or UO_1116 (O_1116,N_24978,N_24839);
xor UO_1117 (O_1117,N_24830,N_24988);
and UO_1118 (O_1118,N_24818,N_24870);
nand UO_1119 (O_1119,N_24871,N_24869);
and UO_1120 (O_1120,N_24946,N_24948);
and UO_1121 (O_1121,N_24837,N_24867);
nand UO_1122 (O_1122,N_24996,N_24971);
or UO_1123 (O_1123,N_24825,N_24820);
or UO_1124 (O_1124,N_24990,N_24841);
and UO_1125 (O_1125,N_24846,N_24874);
and UO_1126 (O_1126,N_24961,N_24869);
nor UO_1127 (O_1127,N_24963,N_24958);
xor UO_1128 (O_1128,N_24805,N_24811);
nor UO_1129 (O_1129,N_24978,N_24961);
or UO_1130 (O_1130,N_24936,N_24871);
xor UO_1131 (O_1131,N_24841,N_24988);
and UO_1132 (O_1132,N_24959,N_24819);
or UO_1133 (O_1133,N_24955,N_24904);
xnor UO_1134 (O_1134,N_24907,N_24808);
and UO_1135 (O_1135,N_24821,N_24954);
and UO_1136 (O_1136,N_24900,N_24944);
and UO_1137 (O_1137,N_24932,N_24850);
and UO_1138 (O_1138,N_24944,N_24971);
nor UO_1139 (O_1139,N_24911,N_24950);
nand UO_1140 (O_1140,N_24855,N_24935);
nor UO_1141 (O_1141,N_24859,N_24930);
nand UO_1142 (O_1142,N_24923,N_24976);
xor UO_1143 (O_1143,N_24953,N_24937);
or UO_1144 (O_1144,N_24848,N_24938);
or UO_1145 (O_1145,N_24805,N_24969);
xnor UO_1146 (O_1146,N_24879,N_24941);
or UO_1147 (O_1147,N_24823,N_24844);
and UO_1148 (O_1148,N_24864,N_24842);
and UO_1149 (O_1149,N_24919,N_24950);
or UO_1150 (O_1150,N_24925,N_24815);
xnor UO_1151 (O_1151,N_24806,N_24920);
nor UO_1152 (O_1152,N_24815,N_24901);
or UO_1153 (O_1153,N_24947,N_24966);
nor UO_1154 (O_1154,N_24987,N_24854);
nor UO_1155 (O_1155,N_24814,N_24816);
xor UO_1156 (O_1156,N_24891,N_24930);
nand UO_1157 (O_1157,N_24958,N_24991);
or UO_1158 (O_1158,N_24936,N_24815);
and UO_1159 (O_1159,N_24842,N_24974);
nand UO_1160 (O_1160,N_24872,N_24914);
nor UO_1161 (O_1161,N_24843,N_24804);
xor UO_1162 (O_1162,N_24825,N_24948);
nand UO_1163 (O_1163,N_24888,N_24848);
and UO_1164 (O_1164,N_24828,N_24860);
or UO_1165 (O_1165,N_24852,N_24923);
nand UO_1166 (O_1166,N_24914,N_24863);
or UO_1167 (O_1167,N_24878,N_24860);
nor UO_1168 (O_1168,N_24986,N_24876);
xor UO_1169 (O_1169,N_24986,N_24886);
nor UO_1170 (O_1170,N_24818,N_24967);
or UO_1171 (O_1171,N_24885,N_24967);
xnor UO_1172 (O_1172,N_24829,N_24930);
and UO_1173 (O_1173,N_24992,N_24984);
or UO_1174 (O_1174,N_24814,N_24909);
nand UO_1175 (O_1175,N_24922,N_24996);
and UO_1176 (O_1176,N_24959,N_24983);
nand UO_1177 (O_1177,N_24820,N_24962);
xor UO_1178 (O_1178,N_24954,N_24894);
and UO_1179 (O_1179,N_24842,N_24969);
or UO_1180 (O_1180,N_24950,N_24913);
nand UO_1181 (O_1181,N_24926,N_24830);
xnor UO_1182 (O_1182,N_24939,N_24887);
xor UO_1183 (O_1183,N_24913,N_24841);
xor UO_1184 (O_1184,N_24803,N_24835);
xor UO_1185 (O_1185,N_24802,N_24861);
xor UO_1186 (O_1186,N_24896,N_24848);
xnor UO_1187 (O_1187,N_24870,N_24980);
xor UO_1188 (O_1188,N_24868,N_24828);
and UO_1189 (O_1189,N_24903,N_24882);
or UO_1190 (O_1190,N_24921,N_24949);
xnor UO_1191 (O_1191,N_24939,N_24929);
or UO_1192 (O_1192,N_24822,N_24911);
nor UO_1193 (O_1193,N_24919,N_24810);
or UO_1194 (O_1194,N_24881,N_24952);
xor UO_1195 (O_1195,N_24825,N_24926);
xor UO_1196 (O_1196,N_24830,N_24918);
or UO_1197 (O_1197,N_24882,N_24964);
nor UO_1198 (O_1198,N_24811,N_24942);
or UO_1199 (O_1199,N_24969,N_24857);
nor UO_1200 (O_1200,N_24946,N_24942);
and UO_1201 (O_1201,N_24825,N_24808);
or UO_1202 (O_1202,N_24983,N_24889);
nor UO_1203 (O_1203,N_24890,N_24813);
nor UO_1204 (O_1204,N_24888,N_24915);
or UO_1205 (O_1205,N_24920,N_24971);
nand UO_1206 (O_1206,N_24985,N_24979);
and UO_1207 (O_1207,N_24836,N_24905);
and UO_1208 (O_1208,N_24967,N_24937);
xnor UO_1209 (O_1209,N_24853,N_24815);
nor UO_1210 (O_1210,N_24913,N_24992);
nor UO_1211 (O_1211,N_24872,N_24888);
and UO_1212 (O_1212,N_24841,N_24951);
nor UO_1213 (O_1213,N_24874,N_24828);
xnor UO_1214 (O_1214,N_24986,N_24897);
and UO_1215 (O_1215,N_24810,N_24950);
or UO_1216 (O_1216,N_24861,N_24916);
and UO_1217 (O_1217,N_24817,N_24980);
nand UO_1218 (O_1218,N_24817,N_24842);
and UO_1219 (O_1219,N_24844,N_24970);
xnor UO_1220 (O_1220,N_24850,N_24928);
nand UO_1221 (O_1221,N_24974,N_24838);
nand UO_1222 (O_1222,N_24851,N_24866);
xnor UO_1223 (O_1223,N_24921,N_24953);
nor UO_1224 (O_1224,N_24942,N_24987);
nand UO_1225 (O_1225,N_24876,N_24909);
nor UO_1226 (O_1226,N_24864,N_24849);
xnor UO_1227 (O_1227,N_24939,N_24942);
or UO_1228 (O_1228,N_24937,N_24924);
or UO_1229 (O_1229,N_24904,N_24981);
nand UO_1230 (O_1230,N_24816,N_24899);
nor UO_1231 (O_1231,N_24965,N_24882);
or UO_1232 (O_1232,N_24962,N_24940);
or UO_1233 (O_1233,N_24976,N_24924);
xnor UO_1234 (O_1234,N_24934,N_24994);
and UO_1235 (O_1235,N_24859,N_24965);
or UO_1236 (O_1236,N_24978,N_24906);
nand UO_1237 (O_1237,N_24890,N_24882);
xnor UO_1238 (O_1238,N_24951,N_24934);
nand UO_1239 (O_1239,N_24921,N_24877);
and UO_1240 (O_1240,N_24993,N_24936);
or UO_1241 (O_1241,N_24935,N_24936);
or UO_1242 (O_1242,N_24909,N_24948);
xnor UO_1243 (O_1243,N_24992,N_24828);
and UO_1244 (O_1244,N_24966,N_24821);
or UO_1245 (O_1245,N_24970,N_24803);
nor UO_1246 (O_1246,N_24848,N_24884);
xnor UO_1247 (O_1247,N_24980,N_24808);
nand UO_1248 (O_1248,N_24842,N_24925);
xor UO_1249 (O_1249,N_24855,N_24809);
nand UO_1250 (O_1250,N_24938,N_24862);
or UO_1251 (O_1251,N_24975,N_24998);
or UO_1252 (O_1252,N_24955,N_24855);
nor UO_1253 (O_1253,N_24834,N_24918);
xor UO_1254 (O_1254,N_24937,N_24976);
nand UO_1255 (O_1255,N_24920,N_24980);
nor UO_1256 (O_1256,N_24838,N_24985);
nand UO_1257 (O_1257,N_24925,N_24809);
nor UO_1258 (O_1258,N_24988,N_24975);
or UO_1259 (O_1259,N_24966,N_24934);
xnor UO_1260 (O_1260,N_24918,N_24933);
nand UO_1261 (O_1261,N_24938,N_24985);
and UO_1262 (O_1262,N_24841,N_24893);
nand UO_1263 (O_1263,N_24885,N_24961);
nand UO_1264 (O_1264,N_24910,N_24828);
nand UO_1265 (O_1265,N_24993,N_24822);
or UO_1266 (O_1266,N_24841,N_24914);
xor UO_1267 (O_1267,N_24829,N_24855);
nor UO_1268 (O_1268,N_24803,N_24808);
nor UO_1269 (O_1269,N_24883,N_24940);
nor UO_1270 (O_1270,N_24911,N_24978);
xor UO_1271 (O_1271,N_24949,N_24882);
and UO_1272 (O_1272,N_24933,N_24816);
nor UO_1273 (O_1273,N_24930,N_24881);
nand UO_1274 (O_1274,N_24835,N_24876);
and UO_1275 (O_1275,N_24821,N_24986);
nor UO_1276 (O_1276,N_24879,N_24997);
and UO_1277 (O_1277,N_24996,N_24881);
or UO_1278 (O_1278,N_24854,N_24919);
xnor UO_1279 (O_1279,N_24944,N_24902);
nand UO_1280 (O_1280,N_24948,N_24849);
nor UO_1281 (O_1281,N_24977,N_24828);
nor UO_1282 (O_1282,N_24911,N_24832);
and UO_1283 (O_1283,N_24955,N_24954);
nand UO_1284 (O_1284,N_24800,N_24869);
and UO_1285 (O_1285,N_24890,N_24935);
or UO_1286 (O_1286,N_24988,N_24963);
and UO_1287 (O_1287,N_24868,N_24830);
and UO_1288 (O_1288,N_24971,N_24952);
xor UO_1289 (O_1289,N_24954,N_24952);
and UO_1290 (O_1290,N_24831,N_24874);
or UO_1291 (O_1291,N_24913,N_24900);
or UO_1292 (O_1292,N_24934,N_24961);
nand UO_1293 (O_1293,N_24924,N_24812);
nor UO_1294 (O_1294,N_24960,N_24968);
nor UO_1295 (O_1295,N_24903,N_24832);
and UO_1296 (O_1296,N_24997,N_24883);
nand UO_1297 (O_1297,N_24834,N_24959);
nor UO_1298 (O_1298,N_24880,N_24987);
or UO_1299 (O_1299,N_24883,N_24976);
xor UO_1300 (O_1300,N_24815,N_24818);
nand UO_1301 (O_1301,N_24975,N_24842);
and UO_1302 (O_1302,N_24946,N_24969);
or UO_1303 (O_1303,N_24965,N_24843);
nand UO_1304 (O_1304,N_24990,N_24884);
xnor UO_1305 (O_1305,N_24995,N_24974);
and UO_1306 (O_1306,N_24997,N_24807);
nand UO_1307 (O_1307,N_24895,N_24813);
nand UO_1308 (O_1308,N_24943,N_24802);
xnor UO_1309 (O_1309,N_24802,N_24846);
and UO_1310 (O_1310,N_24849,N_24943);
or UO_1311 (O_1311,N_24861,N_24918);
or UO_1312 (O_1312,N_24800,N_24892);
xnor UO_1313 (O_1313,N_24877,N_24977);
xor UO_1314 (O_1314,N_24906,N_24943);
xor UO_1315 (O_1315,N_24994,N_24967);
and UO_1316 (O_1316,N_24978,N_24932);
nor UO_1317 (O_1317,N_24952,N_24897);
and UO_1318 (O_1318,N_24805,N_24919);
xnor UO_1319 (O_1319,N_24838,N_24891);
or UO_1320 (O_1320,N_24913,N_24838);
xnor UO_1321 (O_1321,N_24979,N_24911);
nor UO_1322 (O_1322,N_24884,N_24993);
and UO_1323 (O_1323,N_24913,N_24883);
xnor UO_1324 (O_1324,N_24997,N_24925);
or UO_1325 (O_1325,N_24816,N_24812);
nand UO_1326 (O_1326,N_24977,N_24852);
nor UO_1327 (O_1327,N_24904,N_24876);
nor UO_1328 (O_1328,N_24983,N_24989);
nor UO_1329 (O_1329,N_24984,N_24952);
nand UO_1330 (O_1330,N_24941,N_24877);
or UO_1331 (O_1331,N_24840,N_24952);
xor UO_1332 (O_1332,N_24885,N_24842);
nor UO_1333 (O_1333,N_24986,N_24908);
nor UO_1334 (O_1334,N_24989,N_24840);
or UO_1335 (O_1335,N_24848,N_24875);
or UO_1336 (O_1336,N_24996,N_24932);
and UO_1337 (O_1337,N_24829,N_24817);
and UO_1338 (O_1338,N_24952,N_24983);
xor UO_1339 (O_1339,N_24989,N_24844);
xor UO_1340 (O_1340,N_24944,N_24965);
nor UO_1341 (O_1341,N_24877,N_24886);
and UO_1342 (O_1342,N_24920,N_24808);
nor UO_1343 (O_1343,N_24870,N_24988);
xnor UO_1344 (O_1344,N_24959,N_24845);
or UO_1345 (O_1345,N_24910,N_24951);
and UO_1346 (O_1346,N_24947,N_24977);
xor UO_1347 (O_1347,N_24910,N_24906);
xor UO_1348 (O_1348,N_24826,N_24976);
or UO_1349 (O_1349,N_24823,N_24946);
or UO_1350 (O_1350,N_24917,N_24824);
nor UO_1351 (O_1351,N_24812,N_24827);
nor UO_1352 (O_1352,N_24952,N_24895);
or UO_1353 (O_1353,N_24993,N_24821);
nand UO_1354 (O_1354,N_24937,N_24881);
xnor UO_1355 (O_1355,N_24893,N_24962);
xor UO_1356 (O_1356,N_24900,N_24939);
or UO_1357 (O_1357,N_24830,N_24935);
nand UO_1358 (O_1358,N_24930,N_24817);
or UO_1359 (O_1359,N_24987,N_24806);
nor UO_1360 (O_1360,N_24914,N_24891);
or UO_1361 (O_1361,N_24875,N_24839);
and UO_1362 (O_1362,N_24916,N_24957);
or UO_1363 (O_1363,N_24921,N_24917);
nor UO_1364 (O_1364,N_24899,N_24991);
and UO_1365 (O_1365,N_24822,N_24855);
nor UO_1366 (O_1366,N_24889,N_24811);
and UO_1367 (O_1367,N_24863,N_24823);
nand UO_1368 (O_1368,N_24973,N_24960);
and UO_1369 (O_1369,N_24938,N_24948);
or UO_1370 (O_1370,N_24820,N_24807);
nand UO_1371 (O_1371,N_24807,N_24937);
xor UO_1372 (O_1372,N_24862,N_24925);
nand UO_1373 (O_1373,N_24955,N_24974);
and UO_1374 (O_1374,N_24989,N_24994);
or UO_1375 (O_1375,N_24871,N_24847);
or UO_1376 (O_1376,N_24814,N_24889);
or UO_1377 (O_1377,N_24850,N_24976);
nand UO_1378 (O_1378,N_24933,N_24829);
or UO_1379 (O_1379,N_24867,N_24821);
or UO_1380 (O_1380,N_24951,N_24892);
nand UO_1381 (O_1381,N_24910,N_24975);
or UO_1382 (O_1382,N_24817,N_24894);
and UO_1383 (O_1383,N_24934,N_24898);
and UO_1384 (O_1384,N_24896,N_24973);
xor UO_1385 (O_1385,N_24860,N_24819);
xnor UO_1386 (O_1386,N_24954,N_24889);
nor UO_1387 (O_1387,N_24843,N_24911);
or UO_1388 (O_1388,N_24992,N_24996);
xor UO_1389 (O_1389,N_24901,N_24849);
or UO_1390 (O_1390,N_24983,N_24999);
nor UO_1391 (O_1391,N_24903,N_24953);
nand UO_1392 (O_1392,N_24890,N_24892);
or UO_1393 (O_1393,N_24946,N_24982);
and UO_1394 (O_1394,N_24964,N_24893);
xor UO_1395 (O_1395,N_24926,N_24924);
nor UO_1396 (O_1396,N_24982,N_24858);
xnor UO_1397 (O_1397,N_24896,N_24879);
and UO_1398 (O_1398,N_24869,N_24832);
nand UO_1399 (O_1399,N_24857,N_24888);
and UO_1400 (O_1400,N_24976,N_24818);
nand UO_1401 (O_1401,N_24818,N_24978);
and UO_1402 (O_1402,N_24977,N_24940);
or UO_1403 (O_1403,N_24978,N_24940);
nor UO_1404 (O_1404,N_24802,N_24947);
xnor UO_1405 (O_1405,N_24949,N_24937);
nor UO_1406 (O_1406,N_24932,N_24830);
nand UO_1407 (O_1407,N_24982,N_24816);
or UO_1408 (O_1408,N_24830,N_24894);
xor UO_1409 (O_1409,N_24927,N_24913);
xnor UO_1410 (O_1410,N_24932,N_24954);
xnor UO_1411 (O_1411,N_24882,N_24884);
and UO_1412 (O_1412,N_24883,N_24900);
and UO_1413 (O_1413,N_24974,N_24803);
xnor UO_1414 (O_1414,N_24951,N_24936);
nand UO_1415 (O_1415,N_24943,N_24885);
nand UO_1416 (O_1416,N_24905,N_24922);
nand UO_1417 (O_1417,N_24946,N_24975);
nor UO_1418 (O_1418,N_24991,N_24900);
nor UO_1419 (O_1419,N_24968,N_24831);
nor UO_1420 (O_1420,N_24949,N_24965);
or UO_1421 (O_1421,N_24940,N_24826);
or UO_1422 (O_1422,N_24829,N_24815);
xor UO_1423 (O_1423,N_24851,N_24836);
and UO_1424 (O_1424,N_24866,N_24817);
and UO_1425 (O_1425,N_24807,N_24944);
xnor UO_1426 (O_1426,N_24998,N_24802);
nor UO_1427 (O_1427,N_24816,N_24998);
xor UO_1428 (O_1428,N_24822,N_24968);
nor UO_1429 (O_1429,N_24994,N_24912);
or UO_1430 (O_1430,N_24813,N_24841);
nand UO_1431 (O_1431,N_24810,N_24878);
nor UO_1432 (O_1432,N_24970,N_24807);
or UO_1433 (O_1433,N_24938,N_24919);
nand UO_1434 (O_1434,N_24874,N_24833);
nor UO_1435 (O_1435,N_24876,N_24993);
or UO_1436 (O_1436,N_24867,N_24945);
xnor UO_1437 (O_1437,N_24890,N_24857);
xor UO_1438 (O_1438,N_24916,N_24997);
or UO_1439 (O_1439,N_24899,N_24886);
nor UO_1440 (O_1440,N_24945,N_24972);
nand UO_1441 (O_1441,N_24925,N_24929);
nand UO_1442 (O_1442,N_24918,N_24852);
nor UO_1443 (O_1443,N_24861,N_24935);
xnor UO_1444 (O_1444,N_24820,N_24856);
nor UO_1445 (O_1445,N_24909,N_24835);
nand UO_1446 (O_1446,N_24829,N_24838);
nand UO_1447 (O_1447,N_24905,N_24992);
nor UO_1448 (O_1448,N_24937,N_24829);
and UO_1449 (O_1449,N_24801,N_24945);
nor UO_1450 (O_1450,N_24933,N_24896);
and UO_1451 (O_1451,N_24843,N_24954);
xnor UO_1452 (O_1452,N_24866,N_24870);
xnor UO_1453 (O_1453,N_24959,N_24987);
and UO_1454 (O_1454,N_24845,N_24963);
nor UO_1455 (O_1455,N_24815,N_24864);
nor UO_1456 (O_1456,N_24803,N_24998);
and UO_1457 (O_1457,N_24896,N_24995);
nor UO_1458 (O_1458,N_24909,N_24895);
and UO_1459 (O_1459,N_24907,N_24868);
or UO_1460 (O_1460,N_24836,N_24918);
and UO_1461 (O_1461,N_24826,N_24995);
nor UO_1462 (O_1462,N_24846,N_24876);
or UO_1463 (O_1463,N_24937,N_24920);
nand UO_1464 (O_1464,N_24800,N_24874);
and UO_1465 (O_1465,N_24800,N_24907);
or UO_1466 (O_1466,N_24898,N_24974);
nand UO_1467 (O_1467,N_24834,N_24847);
and UO_1468 (O_1468,N_24923,N_24954);
nand UO_1469 (O_1469,N_24928,N_24968);
nand UO_1470 (O_1470,N_24925,N_24967);
xnor UO_1471 (O_1471,N_24807,N_24856);
nor UO_1472 (O_1472,N_24938,N_24859);
or UO_1473 (O_1473,N_24907,N_24891);
nor UO_1474 (O_1474,N_24855,N_24912);
nand UO_1475 (O_1475,N_24938,N_24876);
or UO_1476 (O_1476,N_24881,N_24951);
nor UO_1477 (O_1477,N_24875,N_24824);
xor UO_1478 (O_1478,N_24820,N_24923);
xnor UO_1479 (O_1479,N_24903,N_24980);
nor UO_1480 (O_1480,N_24800,N_24881);
or UO_1481 (O_1481,N_24924,N_24934);
and UO_1482 (O_1482,N_24805,N_24820);
or UO_1483 (O_1483,N_24853,N_24973);
or UO_1484 (O_1484,N_24956,N_24992);
xnor UO_1485 (O_1485,N_24869,N_24928);
or UO_1486 (O_1486,N_24806,N_24966);
nand UO_1487 (O_1487,N_24880,N_24802);
or UO_1488 (O_1488,N_24836,N_24935);
or UO_1489 (O_1489,N_24814,N_24987);
or UO_1490 (O_1490,N_24930,N_24870);
and UO_1491 (O_1491,N_24935,N_24874);
or UO_1492 (O_1492,N_24950,N_24932);
and UO_1493 (O_1493,N_24956,N_24906);
nand UO_1494 (O_1494,N_24898,N_24879);
nand UO_1495 (O_1495,N_24844,N_24931);
and UO_1496 (O_1496,N_24930,N_24921);
xor UO_1497 (O_1497,N_24829,N_24965);
xnor UO_1498 (O_1498,N_24899,N_24807);
and UO_1499 (O_1499,N_24820,N_24944);
and UO_1500 (O_1500,N_24862,N_24892);
nand UO_1501 (O_1501,N_24969,N_24893);
or UO_1502 (O_1502,N_24984,N_24941);
nor UO_1503 (O_1503,N_24840,N_24844);
xor UO_1504 (O_1504,N_24926,N_24838);
and UO_1505 (O_1505,N_24974,N_24855);
nor UO_1506 (O_1506,N_24866,N_24945);
nand UO_1507 (O_1507,N_24971,N_24853);
and UO_1508 (O_1508,N_24860,N_24955);
nor UO_1509 (O_1509,N_24873,N_24987);
or UO_1510 (O_1510,N_24951,N_24862);
xor UO_1511 (O_1511,N_24945,N_24845);
xor UO_1512 (O_1512,N_24923,N_24847);
xnor UO_1513 (O_1513,N_24816,N_24990);
nor UO_1514 (O_1514,N_24976,N_24819);
nand UO_1515 (O_1515,N_24931,N_24984);
xor UO_1516 (O_1516,N_24996,N_24816);
and UO_1517 (O_1517,N_24972,N_24816);
nor UO_1518 (O_1518,N_24982,N_24893);
nor UO_1519 (O_1519,N_24975,N_24987);
xor UO_1520 (O_1520,N_24954,N_24926);
nor UO_1521 (O_1521,N_24853,N_24939);
nand UO_1522 (O_1522,N_24810,N_24841);
and UO_1523 (O_1523,N_24922,N_24815);
and UO_1524 (O_1524,N_24995,N_24996);
nor UO_1525 (O_1525,N_24827,N_24854);
and UO_1526 (O_1526,N_24947,N_24996);
nor UO_1527 (O_1527,N_24946,N_24851);
xor UO_1528 (O_1528,N_24843,N_24883);
and UO_1529 (O_1529,N_24924,N_24974);
or UO_1530 (O_1530,N_24832,N_24918);
and UO_1531 (O_1531,N_24947,N_24848);
and UO_1532 (O_1532,N_24860,N_24980);
and UO_1533 (O_1533,N_24862,N_24825);
nand UO_1534 (O_1534,N_24861,N_24903);
nand UO_1535 (O_1535,N_24939,N_24969);
or UO_1536 (O_1536,N_24939,N_24957);
and UO_1537 (O_1537,N_24966,N_24842);
nand UO_1538 (O_1538,N_24828,N_24941);
and UO_1539 (O_1539,N_24949,N_24863);
nand UO_1540 (O_1540,N_24857,N_24889);
nand UO_1541 (O_1541,N_24964,N_24995);
nor UO_1542 (O_1542,N_24830,N_24958);
or UO_1543 (O_1543,N_24805,N_24991);
nor UO_1544 (O_1544,N_24955,N_24966);
and UO_1545 (O_1545,N_24941,N_24858);
and UO_1546 (O_1546,N_24946,N_24875);
and UO_1547 (O_1547,N_24909,N_24897);
and UO_1548 (O_1548,N_24995,N_24992);
and UO_1549 (O_1549,N_24971,N_24943);
nand UO_1550 (O_1550,N_24917,N_24859);
and UO_1551 (O_1551,N_24923,N_24810);
nand UO_1552 (O_1552,N_24804,N_24932);
nor UO_1553 (O_1553,N_24931,N_24977);
nor UO_1554 (O_1554,N_24999,N_24880);
and UO_1555 (O_1555,N_24841,N_24938);
or UO_1556 (O_1556,N_24942,N_24893);
xor UO_1557 (O_1557,N_24866,N_24923);
nand UO_1558 (O_1558,N_24959,N_24898);
nand UO_1559 (O_1559,N_24952,N_24839);
nor UO_1560 (O_1560,N_24825,N_24993);
and UO_1561 (O_1561,N_24985,N_24959);
and UO_1562 (O_1562,N_24809,N_24838);
or UO_1563 (O_1563,N_24951,N_24896);
or UO_1564 (O_1564,N_24892,N_24834);
and UO_1565 (O_1565,N_24969,N_24807);
and UO_1566 (O_1566,N_24912,N_24811);
or UO_1567 (O_1567,N_24949,N_24903);
nand UO_1568 (O_1568,N_24964,N_24911);
and UO_1569 (O_1569,N_24900,N_24951);
nand UO_1570 (O_1570,N_24931,N_24888);
and UO_1571 (O_1571,N_24955,N_24831);
or UO_1572 (O_1572,N_24893,N_24889);
or UO_1573 (O_1573,N_24842,N_24809);
and UO_1574 (O_1574,N_24992,N_24849);
nand UO_1575 (O_1575,N_24894,N_24825);
nor UO_1576 (O_1576,N_24811,N_24845);
and UO_1577 (O_1577,N_24952,N_24855);
xor UO_1578 (O_1578,N_24935,N_24950);
and UO_1579 (O_1579,N_24859,N_24871);
nand UO_1580 (O_1580,N_24916,N_24943);
nand UO_1581 (O_1581,N_24923,N_24920);
and UO_1582 (O_1582,N_24863,N_24873);
and UO_1583 (O_1583,N_24947,N_24980);
or UO_1584 (O_1584,N_24807,N_24958);
nand UO_1585 (O_1585,N_24861,N_24896);
xor UO_1586 (O_1586,N_24980,N_24965);
xnor UO_1587 (O_1587,N_24878,N_24961);
and UO_1588 (O_1588,N_24873,N_24928);
nor UO_1589 (O_1589,N_24899,N_24933);
xnor UO_1590 (O_1590,N_24947,N_24911);
or UO_1591 (O_1591,N_24817,N_24895);
nor UO_1592 (O_1592,N_24818,N_24843);
and UO_1593 (O_1593,N_24953,N_24894);
and UO_1594 (O_1594,N_24831,N_24943);
and UO_1595 (O_1595,N_24949,N_24868);
nand UO_1596 (O_1596,N_24972,N_24994);
nand UO_1597 (O_1597,N_24847,N_24897);
or UO_1598 (O_1598,N_24910,N_24941);
nor UO_1599 (O_1599,N_24946,N_24929);
nand UO_1600 (O_1600,N_24839,N_24934);
nor UO_1601 (O_1601,N_24811,N_24901);
xor UO_1602 (O_1602,N_24981,N_24964);
xor UO_1603 (O_1603,N_24990,N_24855);
or UO_1604 (O_1604,N_24826,N_24986);
nand UO_1605 (O_1605,N_24836,N_24808);
and UO_1606 (O_1606,N_24835,N_24922);
nand UO_1607 (O_1607,N_24818,N_24963);
nand UO_1608 (O_1608,N_24837,N_24814);
xor UO_1609 (O_1609,N_24909,N_24954);
nand UO_1610 (O_1610,N_24956,N_24991);
nand UO_1611 (O_1611,N_24991,N_24806);
nor UO_1612 (O_1612,N_24929,N_24989);
nand UO_1613 (O_1613,N_24885,N_24986);
or UO_1614 (O_1614,N_24958,N_24926);
nand UO_1615 (O_1615,N_24981,N_24822);
nor UO_1616 (O_1616,N_24926,N_24975);
or UO_1617 (O_1617,N_24998,N_24835);
xor UO_1618 (O_1618,N_24984,N_24942);
nand UO_1619 (O_1619,N_24887,N_24971);
or UO_1620 (O_1620,N_24963,N_24974);
xnor UO_1621 (O_1621,N_24986,N_24902);
and UO_1622 (O_1622,N_24889,N_24890);
nand UO_1623 (O_1623,N_24995,N_24902);
nor UO_1624 (O_1624,N_24971,N_24907);
nor UO_1625 (O_1625,N_24847,N_24989);
xnor UO_1626 (O_1626,N_24803,N_24867);
or UO_1627 (O_1627,N_24956,N_24911);
or UO_1628 (O_1628,N_24835,N_24885);
nor UO_1629 (O_1629,N_24920,N_24929);
xnor UO_1630 (O_1630,N_24878,N_24896);
xnor UO_1631 (O_1631,N_24908,N_24964);
or UO_1632 (O_1632,N_24833,N_24969);
nor UO_1633 (O_1633,N_24806,N_24868);
nand UO_1634 (O_1634,N_24896,N_24920);
nand UO_1635 (O_1635,N_24987,N_24903);
and UO_1636 (O_1636,N_24807,N_24865);
nand UO_1637 (O_1637,N_24826,N_24955);
nor UO_1638 (O_1638,N_24911,N_24878);
and UO_1639 (O_1639,N_24926,N_24870);
or UO_1640 (O_1640,N_24863,N_24890);
nand UO_1641 (O_1641,N_24923,N_24800);
xor UO_1642 (O_1642,N_24885,N_24960);
or UO_1643 (O_1643,N_24972,N_24996);
or UO_1644 (O_1644,N_24960,N_24866);
or UO_1645 (O_1645,N_24948,N_24835);
nand UO_1646 (O_1646,N_24910,N_24914);
xnor UO_1647 (O_1647,N_24936,N_24866);
or UO_1648 (O_1648,N_24867,N_24901);
and UO_1649 (O_1649,N_24818,N_24919);
nand UO_1650 (O_1650,N_24819,N_24851);
nor UO_1651 (O_1651,N_24912,N_24964);
nand UO_1652 (O_1652,N_24823,N_24912);
nand UO_1653 (O_1653,N_24828,N_24960);
and UO_1654 (O_1654,N_24821,N_24917);
and UO_1655 (O_1655,N_24986,N_24900);
and UO_1656 (O_1656,N_24961,N_24937);
xnor UO_1657 (O_1657,N_24929,N_24887);
nand UO_1658 (O_1658,N_24945,N_24891);
or UO_1659 (O_1659,N_24867,N_24863);
or UO_1660 (O_1660,N_24998,N_24874);
nand UO_1661 (O_1661,N_24949,N_24875);
and UO_1662 (O_1662,N_24948,N_24812);
nand UO_1663 (O_1663,N_24820,N_24900);
nand UO_1664 (O_1664,N_24838,N_24820);
nor UO_1665 (O_1665,N_24901,N_24870);
xor UO_1666 (O_1666,N_24911,N_24912);
xor UO_1667 (O_1667,N_24895,N_24902);
nor UO_1668 (O_1668,N_24987,N_24800);
xor UO_1669 (O_1669,N_24833,N_24854);
and UO_1670 (O_1670,N_24972,N_24928);
nand UO_1671 (O_1671,N_24890,N_24818);
xor UO_1672 (O_1672,N_24853,N_24864);
and UO_1673 (O_1673,N_24898,N_24920);
or UO_1674 (O_1674,N_24940,N_24875);
xnor UO_1675 (O_1675,N_24954,N_24933);
nor UO_1676 (O_1676,N_24894,N_24903);
nand UO_1677 (O_1677,N_24881,N_24850);
xnor UO_1678 (O_1678,N_24920,N_24968);
nor UO_1679 (O_1679,N_24984,N_24965);
xor UO_1680 (O_1680,N_24813,N_24923);
nand UO_1681 (O_1681,N_24875,N_24889);
xor UO_1682 (O_1682,N_24925,N_24838);
xor UO_1683 (O_1683,N_24883,N_24990);
nor UO_1684 (O_1684,N_24831,N_24915);
xnor UO_1685 (O_1685,N_24913,N_24958);
nor UO_1686 (O_1686,N_24964,N_24922);
xnor UO_1687 (O_1687,N_24992,N_24946);
nand UO_1688 (O_1688,N_24974,N_24943);
nor UO_1689 (O_1689,N_24957,N_24949);
xor UO_1690 (O_1690,N_24853,N_24833);
and UO_1691 (O_1691,N_24938,N_24895);
nand UO_1692 (O_1692,N_24931,N_24905);
nor UO_1693 (O_1693,N_24812,N_24832);
or UO_1694 (O_1694,N_24865,N_24999);
nor UO_1695 (O_1695,N_24873,N_24866);
xor UO_1696 (O_1696,N_24896,N_24833);
or UO_1697 (O_1697,N_24923,N_24841);
and UO_1698 (O_1698,N_24994,N_24855);
nand UO_1699 (O_1699,N_24815,N_24958);
or UO_1700 (O_1700,N_24820,N_24929);
and UO_1701 (O_1701,N_24914,N_24883);
nand UO_1702 (O_1702,N_24834,N_24922);
nor UO_1703 (O_1703,N_24951,N_24848);
nand UO_1704 (O_1704,N_24878,N_24867);
and UO_1705 (O_1705,N_24881,N_24979);
nand UO_1706 (O_1706,N_24851,N_24880);
nor UO_1707 (O_1707,N_24942,N_24956);
or UO_1708 (O_1708,N_24991,N_24943);
nand UO_1709 (O_1709,N_24813,N_24809);
and UO_1710 (O_1710,N_24965,N_24991);
xor UO_1711 (O_1711,N_24863,N_24969);
xor UO_1712 (O_1712,N_24833,N_24847);
xor UO_1713 (O_1713,N_24888,N_24919);
nor UO_1714 (O_1714,N_24814,N_24907);
or UO_1715 (O_1715,N_24841,N_24858);
and UO_1716 (O_1716,N_24885,N_24841);
and UO_1717 (O_1717,N_24850,N_24803);
or UO_1718 (O_1718,N_24944,N_24950);
xnor UO_1719 (O_1719,N_24931,N_24951);
nor UO_1720 (O_1720,N_24848,N_24975);
nand UO_1721 (O_1721,N_24970,N_24982);
and UO_1722 (O_1722,N_24973,N_24990);
nor UO_1723 (O_1723,N_24862,N_24955);
nor UO_1724 (O_1724,N_24937,N_24834);
or UO_1725 (O_1725,N_24975,N_24894);
nand UO_1726 (O_1726,N_24868,N_24899);
or UO_1727 (O_1727,N_24974,N_24948);
nand UO_1728 (O_1728,N_24942,N_24906);
and UO_1729 (O_1729,N_24962,N_24853);
nor UO_1730 (O_1730,N_24858,N_24992);
and UO_1731 (O_1731,N_24881,N_24895);
nand UO_1732 (O_1732,N_24800,N_24928);
nor UO_1733 (O_1733,N_24895,N_24898);
and UO_1734 (O_1734,N_24840,N_24884);
xor UO_1735 (O_1735,N_24950,N_24981);
nor UO_1736 (O_1736,N_24906,N_24898);
xor UO_1737 (O_1737,N_24855,N_24883);
xnor UO_1738 (O_1738,N_24957,N_24993);
nor UO_1739 (O_1739,N_24942,N_24922);
xnor UO_1740 (O_1740,N_24874,N_24978);
or UO_1741 (O_1741,N_24852,N_24969);
nor UO_1742 (O_1742,N_24962,N_24923);
nand UO_1743 (O_1743,N_24857,N_24922);
xor UO_1744 (O_1744,N_24957,N_24863);
xor UO_1745 (O_1745,N_24940,N_24919);
nand UO_1746 (O_1746,N_24919,N_24980);
xnor UO_1747 (O_1747,N_24890,N_24901);
or UO_1748 (O_1748,N_24971,N_24976);
nor UO_1749 (O_1749,N_24979,N_24968);
nor UO_1750 (O_1750,N_24868,N_24835);
and UO_1751 (O_1751,N_24891,N_24846);
xor UO_1752 (O_1752,N_24983,N_24917);
xor UO_1753 (O_1753,N_24826,N_24891);
or UO_1754 (O_1754,N_24882,N_24897);
xor UO_1755 (O_1755,N_24890,N_24808);
nand UO_1756 (O_1756,N_24903,N_24971);
nor UO_1757 (O_1757,N_24800,N_24917);
nand UO_1758 (O_1758,N_24896,N_24972);
xnor UO_1759 (O_1759,N_24920,N_24824);
or UO_1760 (O_1760,N_24855,N_24807);
nand UO_1761 (O_1761,N_24984,N_24884);
xnor UO_1762 (O_1762,N_24998,N_24872);
xor UO_1763 (O_1763,N_24933,N_24862);
or UO_1764 (O_1764,N_24916,N_24889);
xnor UO_1765 (O_1765,N_24862,N_24861);
nor UO_1766 (O_1766,N_24924,N_24918);
nand UO_1767 (O_1767,N_24913,N_24882);
xor UO_1768 (O_1768,N_24894,N_24978);
xor UO_1769 (O_1769,N_24849,N_24832);
xnor UO_1770 (O_1770,N_24893,N_24840);
or UO_1771 (O_1771,N_24896,N_24889);
or UO_1772 (O_1772,N_24962,N_24861);
and UO_1773 (O_1773,N_24804,N_24944);
and UO_1774 (O_1774,N_24811,N_24841);
nand UO_1775 (O_1775,N_24851,N_24925);
nand UO_1776 (O_1776,N_24915,N_24970);
nand UO_1777 (O_1777,N_24825,N_24835);
xnor UO_1778 (O_1778,N_24876,N_24906);
xor UO_1779 (O_1779,N_24879,N_24998);
xnor UO_1780 (O_1780,N_24827,N_24863);
and UO_1781 (O_1781,N_24907,N_24948);
or UO_1782 (O_1782,N_24883,N_24861);
xnor UO_1783 (O_1783,N_24806,N_24927);
nand UO_1784 (O_1784,N_24814,N_24961);
nand UO_1785 (O_1785,N_24872,N_24883);
or UO_1786 (O_1786,N_24830,N_24865);
or UO_1787 (O_1787,N_24976,N_24895);
nor UO_1788 (O_1788,N_24823,N_24843);
or UO_1789 (O_1789,N_24993,N_24873);
nor UO_1790 (O_1790,N_24971,N_24879);
xnor UO_1791 (O_1791,N_24869,N_24946);
or UO_1792 (O_1792,N_24821,N_24929);
or UO_1793 (O_1793,N_24991,N_24930);
and UO_1794 (O_1794,N_24818,N_24837);
or UO_1795 (O_1795,N_24900,N_24973);
nor UO_1796 (O_1796,N_24829,N_24974);
or UO_1797 (O_1797,N_24828,N_24928);
and UO_1798 (O_1798,N_24959,N_24968);
xor UO_1799 (O_1799,N_24925,N_24974);
nor UO_1800 (O_1800,N_24928,N_24985);
or UO_1801 (O_1801,N_24924,N_24802);
or UO_1802 (O_1802,N_24826,N_24882);
xnor UO_1803 (O_1803,N_24931,N_24877);
nand UO_1804 (O_1804,N_24808,N_24939);
nor UO_1805 (O_1805,N_24878,N_24828);
xnor UO_1806 (O_1806,N_24974,N_24904);
or UO_1807 (O_1807,N_24923,N_24807);
and UO_1808 (O_1808,N_24902,N_24912);
or UO_1809 (O_1809,N_24969,N_24821);
and UO_1810 (O_1810,N_24976,N_24855);
and UO_1811 (O_1811,N_24820,N_24881);
and UO_1812 (O_1812,N_24914,N_24884);
or UO_1813 (O_1813,N_24803,N_24960);
nor UO_1814 (O_1814,N_24807,N_24816);
xor UO_1815 (O_1815,N_24849,N_24900);
or UO_1816 (O_1816,N_24867,N_24938);
nand UO_1817 (O_1817,N_24859,N_24994);
nand UO_1818 (O_1818,N_24973,N_24920);
nor UO_1819 (O_1819,N_24842,N_24918);
nor UO_1820 (O_1820,N_24849,N_24940);
nor UO_1821 (O_1821,N_24974,N_24890);
nor UO_1822 (O_1822,N_24949,N_24859);
nand UO_1823 (O_1823,N_24801,N_24944);
and UO_1824 (O_1824,N_24970,N_24959);
nor UO_1825 (O_1825,N_24829,N_24973);
xnor UO_1826 (O_1826,N_24818,N_24911);
nor UO_1827 (O_1827,N_24927,N_24859);
and UO_1828 (O_1828,N_24960,N_24947);
or UO_1829 (O_1829,N_24999,N_24882);
nor UO_1830 (O_1830,N_24800,N_24894);
nand UO_1831 (O_1831,N_24824,N_24951);
and UO_1832 (O_1832,N_24958,N_24934);
or UO_1833 (O_1833,N_24870,N_24865);
or UO_1834 (O_1834,N_24816,N_24853);
xnor UO_1835 (O_1835,N_24980,N_24863);
nor UO_1836 (O_1836,N_24864,N_24945);
nand UO_1837 (O_1837,N_24902,N_24853);
nor UO_1838 (O_1838,N_24997,N_24952);
and UO_1839 (O_1839,N_24996,N_24906);
or UO_1840 (O_1840,N_24909,N_24881);
and UO_1841 (O_1841,N_24963,N_24889);
or UO_1842 (O_1842,N_24810,N_24944);
or UO_1843 (O_1843,N_24923,N_24979);
nor UO_1844 (O_1844,N_24866,N_24874);
nand UO_1845 (O_1845,N_24964,N_24942);
or UO_1846 (O_1846,N_24817,N_24936);
or UO_1847 (O_1847,N_24972,N_24999);
nor UO_1848 (O_1848,N_24866,N_24890);
nand UO_1849 (O_1849,N_24856,N_24827);
xor UO_1850 (O_1850,N_24835,N_24816);
xnor UO_1851 (O_1851,N_24932,N_24823);
nand UO_1852 (O_1852,N_24982,N_24972);
nand UO_1853 (O_1853,N_24907,N_24920);
nand UO_1854 (O_1854,N_24869,N_24953);
or UO_1855 (O_1855,N_24972,N_24970);
nand UO_1856 (O_1856,N_24805,N_24857);
and UO_1857 (O_1857,N_24959,N_24856);
nor UO_1858 (O_1858,N_24862,N_24937);
and UO_1859 (O_1859,N_24920,N_24825);
xor UO_1860 (O_1860,N_24846,N_24878);
xor UO_1861 (O_1861,N_24905,N_24857);
nand UO_1862 (O_1862,N_24962,N_24883);
nand UO_1863 (O_1863,N_24978,N_24971);
or UO_1864 (O_1864,N_24868,N_24982);
nand UO_1865 (O_1865,N_24982,N_24971);
and UO_1866 (O_1866,N_24901,N_24897);
and UO_1867 (O_1867,N_24966,N_24864);
and UO_1868 (O_1868,N_24855,N_24831);
nor UO_1869 (O_1869,N_24888,N_24815);
nand UO_1870 (O_1870,N_24838,N_24833);
nand UO_1871 (O_1871,N_24968,N_24896);
nor UO_1872 (O_1872,N_24818,N_24832);
nor UO_1873 (O_1873,N_24955,N_24852);
xnor UO_1874 (O_1874,N_24921,N_24935);
and UO_1875 (O_1875,N_24937,N_24938);
and UO_1876 (O_1876,N_24820,N_24811);
and UO_1877 (O_1877,N_24888,N_24869);
nor UO_1878 (O_1878,N_24959,N_24915);
xnor UO_1879 (O_1879,N_24892,N_24893);
xnor UO_1880 (O_1880,N_24800,N_24971);
nor UO_1881 (O_1881,N_24971,N_24928);
and UO_1882 (O_1882,N_24976,N_24900);
nor UO_1883 (O_1883,N_24887,N_24806);
nand UO_1884 (O_1884,N_24902,N_24866);
nand UO_1885 (O_1885,N_24926,N_24888);
nand UO_1886 (O_1886,N_24829,N_24854);
nand UO_1887 (O_1887,N_24904,N_24811);
or UO_1888 (O_1888,N_24907,N_24892);
xnor UO_1889 (O_1889,N_24844,N_24894);
nand UO_1890 (O_1890,N_24843,N_24807);
nand UO_1891 (O_1891,N_24830,N_24866);
or UO_1892 (O_1892,N_24812,N_24869);
nand UO_1893 (O_1893,N_24834,N_24823);
xor UO_1894 (O_1894,N_24878,N_24889);
and UO_1895 (O_1895,N_24845,N_24960);
nand UO_1896 (O_1896,N_24819,N_24892);
nand UO_1897 (O_1897,N_24827,N_24893);
nor UO_1898 (O_1898,N_24806,N_24971);
nand UO_1899 (O_1899,N_24883,N_24809);
and UO_1900 (O_1900,N_24990,N_24977);
and UO_1901 (O_1901,N_24801,N_24875);
and UO_1902 (O_1902,N_24904,N_24953);
or UO_1903 (O_1903,N_24949,N_24956);
nor UO_1904 (O_1904,N_24896,N_24957);
and UO_1905 (O_1905,N_24879,N_24920);
nand UO_1906 (O_1906,N_24903,N_24843);
and UO_1907 (O_1907,N_24961,N_24841);
nand UO_1908 (O_1908,N_24939,N_24811);
xor UO_1909 (O_1909,N_24875,N_24828);
nand UO_1910 (O_1910,N_24952,N_24905);
xnor UO_1911 (O_1911,N_24988,N_24888);
or UO_1912 (O_1912,N_24849,N_24972);
nor UO_1913 (O_1913,N_24935,N_24959);
xor UO_1914 (O_1914,N_24845,N_24913);
and UO_1915 (O_1915,N_24878,N_24813);
nand UO_1916 (O_1916,N_24996,N_24986);
xnor UO_1917 (O_1917,N_24907,N_24877);
nand UO_1918 (O_1918,N_24981,N_24988);
and UO_1919 (O_1919,N_24830,N_24860);
or UO_1920 (O_1920,N_24950,N_24814);
xor UO_1921 (O_1921,N_24864,N_24875);
and UO_1922 (O_1922,N_24999,N_24834);
nor UO_1923 (O_1923,N_24800,N_24943);
xnor UO_1924 (O_1924,N_24953,N_24824);
nand UO_1925 (O_1925,N_24920,N_24850);
and UO_1926 (O_1926,N_24850,N_24817);
xnor UO_1927 (O_1927,N_24861,N_24910);
nor UO_1928 (O_1928,N_24973,N_24961);
nor UO_1929 (O_1929,N_24909,N_24812);
nor UO_1930 (O_1930,N_24858,N_24825);
nand UO_1931 (O_1931,N_24940,N_24805);
and UO_1932 (O_1932,N_24901,N_24858);
nor UO_1933 (O_1933,N_24934,N_24984);
nor UO_1934 (O_1934,N_24919,N_24812);
nor UO_1935 (O_1935,N_24849,N_24823);
or UO_1936 (O_1936,N_24899,N_24939);
nor UO_1937 (O_1937,N_24835,N_24839);
or UO_1938 (O_1938,N_24954,N_24869);
xnor UO_1939 (O_1939,N_24878,N_24946);
and UO_1940 (O_1940,N_24993,N_24946);
xor UO_1941 (O_1941,N_24825,N_24805);
or UO_1942 (O_1942,N_24918,N_24878);
nand UO_1943 (O_1943,N_24983,N_24914);
nand UO_1944 (O_1944,N_24877,N_24940);
nand UO_1945 (O_1945,N_24842,N_24845);
nand UO_1946 (O_1946,N_24823,N_24913);
and UO_1947 (O_1947,N_24914,N_24876);
or UO_1948 (O_1948,N_24919,N_24813);
xor UO_1949 (O_1949,N_24821,N_24863);
and UO_1950 (O_1950,N_24976,N_24940);
and UO_1951 (O_1951,N_24979,N_24866);
nor UO_1952 (O_1952,N_24866,N_24904);
or UO_1953 (O_1953,N_24869,N_24943);
and UO_1954 (O_1954,N_24829,N_24995);
and UO_1955 (O_1955,N_24961,N_24829);
xor UO_1956 (O_1956,N_24854,N_24955);
or UO_1957 (O_1957,N_24841,N_24983);
and UO_1958 (O_1958,N_24886,N_24836);
xor UO_1959 (O_1959,N_24931,N_24837);
or UO_1960 (O_1960,N_24847,N_24896);
and UO_1961 (O_1961,N_24848,N_24874);
xnor UO_1962 (O_1962,N_24998,N_24814);
or UO_1963 (O_1963,N_24943,N_24933);
xnor UO_1964 (O_1964,N_24825,N_24849);
or UO_1965 (O_1965,N_24914,N_24982);
nand UO_1966 (O_1966,N_24837,N_24813);
and UO_1967 (O_1967,N_24867,N_24915);
and UO_1968 (O_1968,N_24871,N_24805);
nand UO_1969 (O_1969,N_24988,N_24848);
and UO_1970 (O_1970,N_24832,N_24954);
or UO_1971 (O_1971,N_24991,N_24829);
and UO_1972 (O_1972,N_24930,N_24925);
xor UO_1973 (O_1973,N_24873,N_24983);
or UO_1974 (O_1974,N_24829,N_24981);
xor UO_1975 (O_1975,N_24854,N_24924);
nor UO_1976 (O_1976,N_24990,N_24818);
and UO_1977 (O_1977,N_24813,N_24808);
nor UO_1978 (O_1978,N_24934,N_24976);
or UO_1979 (O_1979,N_24893,N_24974);
xor UO_1980 (O_1980,N_24964,N_24917);
nand UO_1981 (O_1981,N_24991,N_24998);
nor UO_1982 (O_1982,N_24948,N_24887);
nor UO_1983 (O_1983,N_24861,N_24826);
nor UO_1984 (O_1984,N_24847,N_24911);
xor UO_1985 (O_1985,N_24987,N_24829);
nor UO_1986 (O_1986,N_24996,N_24998);
and UO_1987 (O_1987,N_24891,N_24940);
xor UO_1988 (O_1988,N_24911,N_24821);
or UO_1989 (O_1989,N_24837,N_24940);
nor UO_1990 (O_1990,N_24882,N_24955);
or UO_1991 (O_1991,N_24975,N_24859);
and UO_1992 (O_1992,N_24875,N_24912);
nand UO_1993 (O_1993,N_24824,N_24944);
and UO_1994 (O_1994,N_24969,N_24856);
xor UO_1995 (O_1995,N_24871,N_24880);
xor UO_1996 (O_1996,N_24850,N_24826);
nor UO_1997 (O_1997,N_24959,N_24998);
and UO_1998 (O_1998,N_24877,N_24997);
xor UO_1999 (O_1999,N_24897,N_24854);
xnor UO_2000 (O_2000,N_24930,N_24835);
nand UO_2001 (O_2001,N_24914,N_24906);
xnor UO_2002 (O_2002,N_24989,N_24992);
nor UO_2003 (O_2003,N_24856,N_24868);
or UO_2004 (O_2004,N_24924,N_24896);
and UO_2005 (O_2005,N_24963,N_24994);
nor UO_2006 (O_2006,N_24866,N_24836);
xor UO_2007 (O_2007,N_24989,N_24906);
or UO_2008 (O_2008,N_24946,N_24960);
xor UO_2009 (O_2009,N_24879,N_24850);
nand UO_2010 (O_2010,N_24953,N_24962);
or UO_2011 (O_2011,N_24802,N_24968);
nand UO_2012 (O_2012,N_24864,N_24923);
xnor UO_2013 (O_2013,N_24812,N_24811);
and UO_2014 (O_2014,N_24871,N_24958);
and UO_2015 (O_2015,N_24944,N_24832);
nand UO_2016 (O_2016,N_24982,N_24983);
nor UO_2017 (O_2017,N_24933,N_24846);
xor UO_2018 (O_2018,N_24933,N_24920);
and UO_2019 (O_2019,N_24898,N_24847);
and UO_2020 (O_2020,N_24837,N_24958);
nor UO_2021 (O_2021,N_24892,N_24880);
or UO_2022 (O_2022,N_24852,N_24868);
nor UO_2023 (O_2023,N_24851,N_24845);
xnor UO_2024 (O_2024,N_24808,N_24985);
nor UO_2025 (O_2025,N_24960,N_24895);
nor UO_2026 (O_2026,N_24852,N_24835);
nand UO_2027 (O_2027,N_24837,N_24847);
nand UO_2028 (O_2028,N_24837,N_24848);
nor UO_2029 (O_2029,N_24841,N_24817);
or UO_2030 (O_2030,N_24898,N_24823);
or UO_2031 (O_2031,N_24842,N_24816);
xor UO_2032 (O_2032,N_24917,N_24895);
nand UO_2033 (O_2033,N_24827,N_24831);
or UO_2034 (O_2034,N_24870,N_24956);
or UO_2035 (O_2035,N_24867,N_24950);
nand UO_2036 (O_2036,N_24912,N_24842);
nand UO_2037 (O_2037,N_24937,N_24809);
and UO_2038 (O_2038,N_24898,N_24967);
xnor UO_2039 (O_2039,N_24851,N_24897);
xor UO_2040 (O_2040,N_24811,N_24916);
nand UO_2041 (O_2041,N_24985,N_24966);
or UO_2042 (O_2042,N_24875,N_24958);
xor UO_2043 (O_2043,N_24976,N_24964);
nand UO_2044 (O_2044,N_24980,N_24969);
and UO_2045 (O_2045,N_24972,N_24987);
xnor UO_2046 (O_2046,N_24914,N_24896);
xor UO_2047 (O_2047,N_24909,N_24800);
nor UO_2048 (O_2048,N_24891,N_24808);
nor UO_2049 (O_2049,N_24902,N_24906);
nand UO_2050 (O_2050,N_24837,N_24893);
xor UO_2051 (O_2051,N_24910,N_24901);
nand UO_2052 (O_2052,N_24991,N_24872);
nor UO_2053 (O_2053,N_24838,N_24959);
and UO_2054 (O_2054,N_24830,N_24827);
xor UO_2055 (O_2055,N_24953,N_24988);
and UO_2056 (O_2056,N_24965,N_24918);
nand UO_2057 (O_2057,N_24933,N_24902);
nor UO_2058 (O_2058,N_24830,N_24891);
nand UO_2059 (O_2059,N_24926,N_24847);
nor UO_2060 (O_2060,N_24937,N_24991);
or UO_2061 (O_2061,N_24905,N_24928);
nor UO_2062 (O_2062,N_24984,N_24954);
or UO_2063 (O_2063,N_24832,N_24925);
or UO_2064 (O_2064,N_24888,N_24908);
or UO_2065 (O_2065,N_24847,N_24979);
xnor UO_2066 (O_2066,N_24857,N_24976);
or UO_2067 (O_2067,N_24893,N_24818);
and UO_2068 (O_2068,N_24892,N_24860);
nand UO_2069 (O_2069,N_24835,N_24927);
nor UO_2070 (O_2070,N_24918,N_24977);
xnor UO_2071 (O_2071,N_24847,N_24946);
nor UO_2072 (O_2072,N_24940,N_24914);
and UO_2073 (O_2073,N_24875,N_24994);
and UO_2074 (O_2074,N_24901,N_24808);
xnor UO_2075 (O_2075,N_24814,N_24912);
nand UO_2076 (O_2076,N_24921,N_24801);
xor UO_2077 (O_2077,N_24891,N_24993);
nand UO_2078 (O_2078,N_24829,N_24876);
nor UO_2079 (O_2079,N_24869,N_24865);
nor UO_2080 (O_2080,N_24892,N_24837);
nor UO_2081 (O_2081,N_24825,N_24967);
xnor UO_2082 (O_2082,N_24979,N_24935);
nor UO_2083 (O_2083,N_24920,N_24877);
xor UO_2084 (O_2084,N_24985,N_24964);
and UO_2085 (O_2085,N_24933,N_24993);
nand UO_2086 (O_2086,N_24876,N_24837);
or UO_2087 (O_2087,N_24905,N_24858);
and UO_2088 (O_2088,N_24868,N_24881);
nand UO_2089 (O_2089,N_24995,N_24953);
and UO_2090 (O_2090,N_24917,N_24820);
and UO_2091 (O_2091,N_24989,N_24957);
xnor UO_2092 (O_2092,N_24825,N_24976);
nand UO_2093 (O_2093,N_24893,N_24873);
nand UO_2094 (O_2094,N_24865,N_24805);
and UO_2095 (O_2095,N_24856,N_24991);
nand UO_2096 (O_2096,N_24986,N_24914);
and UO_2097 (O_2097,N_24810,N_24899);
nand UO_2098 (O_2098,N_24988,N_24976);
xnor UO_2099 (O_2099,N_24916,N_24977);
and UO_2100 (O_2100,N_24827,N_24921);
and UO_2101 (O_2101,N_24962,N_24963);
and UO_2102 (O_2102,N_24830,N_24878);
xnor UO_2103 (O_2103,N_24967,N_24981);
nand UO_2104 (O_2104,N_24843,N_24946);
xnor UO_2105 (O_2105,N_24875,N_24982);
or UO_2106 (O_2106,N_24934,N_24938);
nor UO_2107 (O_2107,N_24954,N_24899);
nand UO_2108 (O_2108,N_24943,N_24993);
nand UO_2109 (O_2109,N_24970,N_24953);
or UO_2110 (O_2110,N_24814,N_24941);
nor UO_2111 (O_2111,N_24914,N_24969);
xor UO_2112 (O_2112,N_24859,N_24928);
and UO_2113 (O_2113,N_24941,N_24809);
or UO_2114 (O_2114,N_24842,N_24987);
and UO_2115 (O_2115,N_24859,N_24915);
nand UO_2116 (O_2116,N_24875,N_24857);
xor UO_2117 (O_2117,N_24889,N_24939);
xor UO_2118 (O_2118,N_24987,N_24890);
nand UO_2119 (O_2119,N_24931,N_24910);
nor UO_2120 (O_2120,N_24826,N_24834);
and UO_2121 (O_2121,N_24853,N_24876);
nor UO_2122 (O_2122,N_24918,N_24996);
nand UO_2123 (O_2123,N_24964,N_24871);
nand UO_2124 (O_2124,N_24887,N_24968);
xnor UO_2125 (O_2125,N_24967,N_24841);
or UO_2126 (O_2126,N_24828,N_24862);
xor UO_2127 (O_2127,N_24827,N_24836);
and UO_2128 (O_2128,N_24982,N_24803);
nand UO_2129 (O_2129,N_24971,N_24975);
nor UO_2130 (O_2130,N_24925,N_24812);
and UO_2131 (O_2131,N_24994,N_24986);
nand UO_2132 (O_2132,N_24870,N_24911);
or UO_2133 (O_2133,N_24864,N_24835);
nor UO_2134 (O_2134,N_24931,N_24944);
or UO_2135 (O_2135,N_24917,N_24929);
and UO_2136 (O_2136,N_24907,N_24904);
nand UO_2137 (O_2137,N_24997,N_24947);
nor UO_2138 (O_2138,N_24954,N_24809);
nand UO_2139 (O_2139,N_24803,N_24905);
nor UO_2140 (O_2140,N_24844,N_24913);
nor UO_2141 (O_2141,N_24975,N_24916);
xor UO_2142 (O_2142,N_24910,N_24821);
and UO_2143 (O_2143,N_24912,N_24957);
xor UO_2144 (O_2144,N_24999,N_24992);
or UO_2145 (O_2145,N_24899,N_24921);
or UO_2146 (O_2146,N_24819,N_24883);
nor UO_2147 (O_2147,N_24810,N_24976);
and UO_2148 (O_2148,N_24849,N_24997);
nor UO_2149 (O_2149,N_24844,N_24958);
nor UO_2150 (O_2150,N_24805,N_24856);
nand UO_2151 (O_2151,N_24941,N_24991);
nor UO_2152 (O_2152,N_24944,N_24853);
xor UO_2153 (O_2153,N_24927,N_24935);
xnor UO_2154 (O_2154,N_24979,N_24897);
nand UO_2155 (O_2155,N_24962,N_24909);
and UO_2156 (O_2156,N_24839,N_24957);
xnor UO_2157 (O_2157,N_24901,N_24841);
xnor UO_2158 (O_2158,N_24874,N_24921);
and UO_2159 (O_2159,N_24866,N_24844);
xor UO_2160 (O_2160,N_24979,N_24820);
and UO_2161 (O_2161,N_24820,N_24860);
or UO_2162 (O_2162,N_24861,N_24875);
or UO_2163 (O_2163,N_24908,N_24815);
nand UO_2164 (O_2164,N_24910,N_24984);
and UO_2165 (O_2165,N_24802,N_24969);
nor UO_2166 (O_2166,N_24931,N_24812);
or UO_2167 (O_2167,N_24896,N_24849);
or UO_2168 (O_2168,N_24945,N_24993);
nor UO_2169 (O_2169,N_24903,N_24881);
nor UO_2170 (O_2170,N_24995,N_24916);
nor UO_2171 (O_2171,N_24962,N_24941);
or UO_2172 (O_2172,N_24879,N_24985);
xor UO_2173 (O_2173,N_24967,N_24880);
xnor UO_2174 (O_2174,N_24895,N_24975);
and UO_2175 (O_2175,N_24881,N_24897);
nor UO_2176 (O_2176,N_24857,N_24957);
and UO_2177 (O_2177,N_24934,N_24918);
nor UO_2178 (O_2178,N_24958,N_24833);
nand UO_2179 (O_2179,N_24875,N_24908);
xor UO_2180 (O_2180,N_24874,N_24820);
or UO_2181 (O_2181,N_24803,N_24813);
nor UO_2182 (O_2182,N_24891,N_24917);
xor UO_2183 (O_2183,N_24908,N_24805);
nand UO_2184 (O_2184,N_24913,N_24952);
nor UO_2185 (O_2185,N_24986,N_24993);
nand UO_2186 (O_2186,N_24892,N_24811);
nor UO_2187 (O_2187,N_24980,N_24864);
xnor UO_2188 (O_2188,N_24976,N_24943);
nor UO_2189 (O_2189,N_24891,N_24856);
or UO_2190 (O_2190,N_24853,N_24945);
xnor UO_2191 (O_2191,N_24922,N_24898);
xor UO_2192 (O_2192,N_24859,N_24815);
and UO_2193 (O_2193,N_24987,N_24884);
or UO_2194 (O_2194,N_24866,N_24903);
or UO_2195 (O_2195,N_24927,N_24885);
and UO_2196 (O_2196,N_24905,N_24813);
or UO_2197 (O_2197,N_24891,N_24901);
xor UO_2198 (O_2198,N_24839,N_24810);
nand UO_2199 (O_2199,N_24811,N_24944);
and UO_2200 (O_2200,N_24988,N_24854);
xnor UO_2201 (O_2201,N_24853,N_24912);
and UO_2202 (O_2202,N_24991,N_24997);
and UO_2203 (O_2203,N_24802,N_24892);
nor UO_2204 (O_2204,N_24861,N_24906);
nand UO_2205 (O_2205,N_24993,N_24920);
and UO_2206 (O_2206,N_24900,N_24861);
or UO_2207 (O_2207,N_24985,N_24865);
and UO_2208 (O_2208,N_24981,N_24801);
and UO_2209 (O_2209,N_24863,N_24928);
nand UO_2210 (O_2210,N_24832,N_24878);
nor UO_2211 (O_2211,N_24849,N_24916);
nand UO_2212 (O_2212,N_24912,N_24929);
or UO_2213 (O_2213,N_24801,N_24815);
nor UO_2214 (O_2214,N_24915,N_24955);
xnor UO_2215 (O_2215,N_24980,N_24880);
xor UO_2216 (O_2216,N_24972,N_24922);
and UO_2217 (O_2217,N_24871,N_24904);
and UO_2218 (O_2218,N_24832,N_24940);
xor UO_2219 (O_2219,N_24935,N_24833);
nor UO_2220 (O_2220,N_24923,N_24999);
xnor UO_2221 (O_2221,N_24889,N_24941);
xnor UO_2222 (O_2222,N_24915,N_24813);
or UO_2223 (O_2223,N_24922,N_24829);
nand UO_2224 (O_2224,N_24950,N_24801);
xnor UO_2225 (O_2225,N_24887,N_24955);
and UO_2226 (O_2226,N_24828,N_24836);
or UO_2227 (O_2227,N_24874,N_24858);
or UO_2228 (O_2228,N_24807,N_24918);
xnor UO_2229 (O_2229,N_24890,N_24833);
and UO_2230 (O_2230,N_24935,N_24825);
nand UO_2231 (O_2231,N_24815,N_24874);
nor UO_2232 (O_2232,N_24998,N_24891);
and UO_2233 (O_2233,N_24801,N_24910);
nor UO_2234 (O_2234,N_24823,N_24811);
or UO_2235 (O_2235,N_24910,N_24871);
xor UO_2236 (O_2236,N_24859,N_24854);
nor UO_2237 (O_2237,N_24913,N_24849);
xnor UO_2238 (O_2238,N_24816,N_24965);
nand UO_2239 (O_2239,N_24880,N_24889);
and UO_2240 (O_2240,N_24936,N_24877);
nor UO_2241 (O_2241,N_24927,N_24851);
nor UO_2242 (O_2242,N_24904,N_24984);
or UO_2243 (O_2243,N_24905,N_24802);
and UO_2244 (O_2244,N_24800,N_24957);
xor UO_2245 (O_2245,N_24999,N_24954);
nor UO_2246 (O_2246,N_24886,N_24916);
xnor UO_2247 (O_2247,N_24881,N_24944);
nor UO_2248 (O_2248,N_24859,N_24808);
nand UO_2249 (O_2249,N_24983,N_24956);
xor UO_2250 (O_2250,N_24804,N_24841);
or UO_2251 (O_2251,N_24899,N_24972);
and UO_2252 (O_2252,N_24884,N_24916);
and UO_2253 (O_2253,N_24907,N_24967);
xor UO_2254 (O_2254,N_24861,N_24991);
nor UO_2255 (O_2255,N_24811,N_24941);
and UO_2256 (O_2256,N_24819,N_24859);
and UO_2257 (O_2257,N_24936,N_24883);
nor UO_2258 (O_2258,N_24833,N_24919);
nand UO_2259 (O_2259,N_24973,N_24916);
and UO_2260 (O_2260,N_24834,N_24882);
or UO_2261 (O_2261,N_24868,N_24809);
xnor UO_2262 (O_2262,N_24902,N_24857);
nand UO_2263 (O_2263,N_24889,N_24846);
or UO_2264 (O_2264,N_24834,N_24994);
nand UO_2265 (O_2265,N_24898,N_24980);
or UO_2266 (O_2266,N_24913,N_24917);
and UO_2267 (O_2267,N_24973,N_24849);
xnor UO_2268 (O_2268,N_24854,N_24957);
and UO_2269 (O_2269,N_24883,N_24944);
nand UO_2270 (O_2270,N_24831,N_24850);
nand UO_2271 (O_2271,N_24991,N_24831);
xnor UO_2272 (O_2272,N_24832,N_24847);
or UO_2273 (O_2273,N_24978,N_24836);
nor UO_2274 (O_2274,N_24825,N_24947);
nor UO_2275 (O_2275,N_24948,N_24939);
and UO_2276 (O_2276,N_24855,N_24931);
nand UO_2277 (O_2277,N_24854,N_24880);
nor UO_2278 (O_2278,N_24859,N_24986);
nand UO_2279 (O_2279,N_24948,N_24943);
nor UO_2280 (O_2280,N_24896,N_24921);
or UO_2281 (O_2281,N_24858,N_24898);
or UO_2282 (O_2282,N_24900,N_24826);
or UO_2283 (O_2283,N_24932,N_24926);
and UO_2284 (O_2284,N_24830,N_24803);
or UO_2285 (O_2285,N_24829,N_24884);
nor UO_2286 (O_2286,N_24965,N_24852);
nand UO_2287 (O_2287,N_24887,N_24959);
or UO_2288 (O_2288,N_24974,N_24892);
xor UO_2289 (O_2289,N_24957,N_24927);
nor UO_2290 (O_2290,N_24822,N_24895);
nor UO_2291 (O_2291,N_24834,N_24885);
nand UO_2292 (O_2292,N_24974,N_24944);
nor UO_2293 (O_2293,N_24834,N_24905);
nor UO_2294 (O_2294,N_24945,N_24973);
xor UO_2295 (O_2295,N_24965,N_24888);
and UO_2296 (O_2296,N_24875,N_24868);
and UO_2297 (O_2297,N_24858,N_24989);
and UO_2298 (O_2298,N_24866,N_24856);
nand UO_2299 (O_2299,N_24934,N_24971);
or UO_2300 (O_2300,N_24903,N_24809);
xnor UO_2301 (O_2301,N_24956,N_24966);
xnor UO_2302 (O_2302,N_24894,N_24874);
and UO_2303 (O_2303,N_24828,N_24872);
nand UO_2304 (O_2304,N_24869,N_24998);
xnor UO_2305 (O_2305,N_24826,N_24909);
and UO_2306 (O_2306,N_24938,N_24912);
nor UO_2307 (O_2307,N_24967,N_24929);
xor UO_2308 (O_2308,N_24851,N_24920);
nand UO_2309 (O_2309,N_24804,N_24902);
or UO_2310 (O_2310,N_24890,N_24981);
or UO_2311 (O_2311,N_24899,N_24829);
nand UO_2312 (O_2312,N_24966,N_24869);
xor UO_2313 (O_2313,N_24925,N_24991);
or UO_2314 (O_2314,N_24892,N_24900);
nor UO_2315 (O_2315,N_24837,N_24983);
xor UO_2316 (O_2316,N_24917,N_24846);
xor UO_2317 (O_2317,N_24833,N_24914);
nor UO_2318 (O_2318,N_24834,N_24919);
or UO_2319 (O_2319,N_24911,N_24929);
and UO_2320 (O_2320,N_24827,N_24865);
or UO_2321 (O_2321,N_24807,N_24824);
or UO_2322 (O_2322,N_24967,N_24954);
and UO_2323 (O_2323,N_24968,N_24950);
xnor UO_2324 (O_2324,N_24811,N_24803);
nor UO_2325 (O_2325,N_24820,N_24815);
nor UO_2326 (O_2326,N_24971,N_24966);
nand UO_2327 (O_2327,N_24995,N_24967);
or UO_2328 (O_2328,N_24890,N_24909);
or UO_2329 (O_2329,N_24999,N_24900);
or UO_2330 (O_2330,N_24860,N_24818);
or UO_2331 (O_2331,N_24950,N_24954);
or UO_2332 (O_2332,N_24985,N_24831);
nor UO_2333 (O_2333,N_24977,N_24903);
nor UO_2334 (O_2334,N_24858,N_24933);
nand UO_2335 (O_2335,N_24823,N_24822);
xor UO_2336 (O_2336,N_24918,N_24897);
nor UO_2337 (O_2337,N_24827,N_24811);
or UO_2338 (O_2338,N_24848,N_24870);
nor UO_2339 (O_2339,N_24962,N_24843);
or UO_2340 (O_2340,N_24839,N_24979);
or UO_2341 (O_2341,N_24921,N_24984);
or UO_2342 (O_2342,N_24986,N_24840);
xnor UO_2343 (O_2343,N_24893,N_24810);
or UO_2344 (O_2344,N_24893,N_24857);
and UO_2345 (O_2345,N_24942,N_24929);
nand UO_2346 (O_2346,N_24945,N_24823);
and UO_2347 (O_2347,N_24899,N_24996);
nand UO_2348 (O_2348,N_24907,N_24963);
nor UO_2349 (O_2349,N_24845,N_24856);
xnor UO_2350 (O_2350,N_24987,N_24822);
xnor UO_2351 (O_2351,N_24913,N_24969);
nand UO_2352 (O_2352,N_24880,N_24939);
nand UO_2353 (O_2353,N_24864,N_24861);
and UO_2354 (O_2354,N_24822,N_24980);
xnor UO_2355 (O_2355,N_24866,N_24992);
nand UO_2356 (O_2356,N_24916,N_24813);
nand UO_2357 (O_2357,N_24896,N_24857);
or UO_2358 (O_2358,N_24857,N_24885);
and UO_2359 (O_2359,N_24920,N_24917);
xnor UO_2360 (O_2360,N_24849,N_24891);
xnor UO_2361 (O_2361,N_24878,N_24886);
nor UO_2362 (O_2362,N_24906,N_24979);
and UO_2363 (O_2363,N_24951,N_24864);
nor UO_2364 (O_2364,N_24997,N_24820);
and UO_2365 (O_2365,N_24901,N_24843);
nand UO_2366 (O_2366,N_24932,N_24911);
or UO_2367 (O_2367,N_24922,N_24897);
nor UO_2368 (O_2368,N_24898,N_24854);
nand UO_2369 (O_2369,N_24832,N_24886);
nor UO_2370 (O_2370,N_24855,N_24875);
xnor UO_2371 (O_2371,N_24967,N_24945);
xor UO_2372 (O_2372,N_24947,N_24830);
xnor UO_2373 (O_2373,N_24954,N_24929);
nor UO_2374 (O_2374,N_24828,N_24918);
xnor UO_2375 (O_2375,N_24855,N_24844);
nor UO_2376 (O_2376,N_24913,N_24848);
and UO_2377 (O_2377,N_24846,N_24922);
nor UO_2378 (O_2378,N_24906,N_24960);
xnor UO_2379 (O_2379,N_24853,N_24800);
nor UO_2380 (O_2380,N_24959,N_24864);
xnor UO_2381 (O_2381,N_24946,N_24991);
or UO_2382 (O_2382,N_24905,N_24842);
and UO_2383 (O_2383,N_24906,N_24832);
xor UO_2384 (O_2384,N_24900,N_24902);
nand UO_2385 (O_2385,N_24827,N_24851);
and UO_2386 (O_2386,N_24959,N_24818);
or UO_2387 (O_2387,N_24808,N_24926);
or UO_2388 (O_2388,N_24816,N_24967);
nand UO_2389 (O_2389,N_24898,N_24838);
or UO_2390 (O_2390,N_24951,N_24839);
or UO_2391 (O_2391,N_24903,N_24978);
or UO_2392 (O_2392,N_24974,N_24959);
nand UO_2393 (O_2393,N_24923,N_24931);
and UO_2394 (O_2394,N_24975,N_24891);
xnor UO_2395 (O_2395,N_24923,N_24838);
nor UO_2396 (O_2396,N_24822,N_24882);
nor UO_2397 (O_2397,N_24829,N_24904);
and UO_2398 (O_2398,N_24875,N_24841);
nand UO_2399 (O_2399,N_24926,N_24901);
xnor UO_2400 (O_2400,N_24856,N_24849);
nand UO_2401 (O_2401,N_24935,N_24940);
nor UO_2402 (O_2402,N_24859,N_24979);
and UO_2403 (O_2403,N_24867,N_24969);
or UO_2404 (O_2404,N_24928,N_24957);
nor UO_2405 (O_2405,N_24929,N_24924);
nor UO_2406 (O_2406,N_24882,N_24973);
xor UO_2407 (O_2407,N_24925,N_24876);
or UO_2408 (O_2408,N_24984,N_24802);
and UO_2409 (O_2409,N_24992,N_24919);
nor UO_2410 (O_2410,N_24843,N_24928);
nand UO_2411 (O_2411,N_24881,N_24972);
nor UO_2412 (O_2412,N_24875,N_24842);
and UO_2413 (O_2413,N_24945,N_24930);
and UO_2414 (O_2414,N_24969,N_24854);
nor UO_2415 (O_2415,N_24934,N_24849);
nand UO_2416 (O_2416,N_24876,N_24893);
or UO_2417 (O_2417,N_24935,N_24953);
xnor UO_2418 (O_2418,N_24823,N_24867);
nor UO_2419 (O_2419,N_24836,N_24934);
nor UO_2420 (O_2420,N_24975,N_24932);
or UO_2421 (O_2421,N_24912,N_24959);
or UO_2422 (O_2422,N_24828,N_24925);
xnor UO_2423 (O_2423,N_24921,N_24820);
xnor UO_2424 (O_2424,N_24970,N_24958);
nor UO_2425 (O_2425,N_24914,N_24850);
xnor UO_2426 (O_2426,N_24949,N_24852);
nor UO_2427 (O_2427,N_24902,N_24825);
nor UO_2428 (O_2428,N_24973,N_24901);
nor UO_2429 (O_2429,N_24804,N_24962);
or UO_2430 (O_2430,N_24901,N_24857);
nor UO_2431 (O_2431,N_24984,N_24845);
nor UO_2432 (O_2432,N_24838,N_24965);
nor UO_2433 (O_2433,N_24940,N_24951);
and UO_2434 (O_2434,N_24967,N_24854);
or UO_2435 (O_2435,N_24836,N_24919);
nand UO_2436 (O_2436,N_24811,N_24966);
or UO_2437 (O_2437,N_24806,N_24982);
and UO_2438 (O_2438,N_24835,N_24853);
and UO_2439 (O_2439,N_24969,N_24905);
and UO_2440 (O_2440,N_24879,N_24859);
nand UO_2441 (O_2441,N_24994,N_24801);
or UO_2442 (O_2442,N_24861,N_24857);
nand UO_2443 (O_2443,N_24939,N_24822);
xnor UO_2444 (O_2444,N_24944,N_24966);
and UO_2445 (O_2445,N_24901,N_24882);
xnor UO_2446 (O_2446,N_24800,N_24899);
xor UO_2447 (O_2447,N_24878,N_24917);
and UO_2448 (O_2448,N_24813,N_24914);
nand UO_2449 (O_2449,N_24937,N_24845);
nor UO_2450 (O_2450,N_24832,N_24962);
nor UO_2451 (O_2451,N_24949,N_24931);
xor UO_2452 (O_2452,N_24824,N_24938);
or UO_2453 (O_2453,N_24966,N_24883);
nand UO_2454 (O_2454,N_24801,N_24811);
and UO_2455 (O_2455,N_24880,N_24898);
nor UO_2456 (O_2456,N_24953,N_24851);
or UO_2457 (O_2457,N_24880,N_24902);
and UO_2458 (O_2458,N_24970,N_24879);
xor UO_2459 (O_2459,N_24907,N_24846);
and UO_2460 (O_2460,N_24923,N_24988);
nor UO_2461 (O_2461,N_24901,N_24908);
or UO_2462 (O_2462,N_24849,N_24919);
nor UO_2463 (O_2463,N_24960,N_24873);
xnor UO_2464 (O_2464,N_24867,N_24808);
xor UO_2465 (O_2465,N_24851,N_24885);
nand UO_2466 (O_2466,N_24931,N_24898);
xnor UO_2467 (O_2467,N_24910,N_24912);
or UO_2468 (O_2468,N_24837,N_24920);
and UO_2469 (O_2469,N_24944,N_24936);
nand UO_2470 (O_2470,N_24838,N_24906);
or UO_2471 (O_2471,N_24803,N_24860);
nor UO_2472 (O_2472,N_24995,N_24933);
and UO_2473 (O_2473,N_24873,N_24980);
nor UO_2474 (O_2474,N_24898,N_24829);
xor UO_2475 (O_2475,N_24838,N_24834);
or UO_2476 (O_2476,N_24877,N_24807);
and UO_2477 (O_2477,N_24843,N_24829);
nor UO_2478 (O_2478,N_24996,N_24895);
or UO_2479 (O_2479,N_24973,N_24930);
and UO_2480 (O_2480,N_24947,N_24910);
nand UO_2481 (O_2481,N_24980,N_24837);
xnor UO_2482 (O_2482,N_24986,N_24856);
nor UO_2483 (O_2483,N_24930,N_24888);
nand UO_2484 (O_2484,N_24820,N_24821);
and UO_2485 (O_2485,N_24951,N_24918);
xnor UO_2486 (O_2486,N_24800,N_24821);
and UO_2487 (O_2487,N_24890,N_24823);
or UO_2488 (O_2488,N_24978,N_24990);
or UO_2489 (O_2489,N_24892,N_24883);
and UO_2490 (O_2490,N_24828,N_24861);
nor UO_2491 (O_2491,N_24828,N_24965);
or UO_2492 (O_2492,N_24821,N_24948);
nand UO_2493 (O_2493,N_24841,N_24840);
or UO_2494 (O_2494,N_24985,N_24949);
or UO_2495 (O_2495,N_24903,N_24878);
nor UO_2496 (O_2496,N_24919,N_24957);
and UO_2497 (O_2497,N_24961,N_24873);
nor UO_2498 (O_2498,N_24817,N_24927);
nor UO_2499 (O_2499,N_24976,N_24982);
and UO_2500 (O_2500,N_24904,N_24902);
nand UO_2501 (O_2501,N_24960,N_24881);
or UO_2502 (O_2502,N_24947,N_24873);
and UO_2503 (O_2503,N_24884,N_24982);
or UO_2504 (O_2504,N_24832,N_24959);
nand UO_2505 (O_2505,N_24882,N_24810);
xor UO_2506 (O_2506,N_24923,N_24890);
and UO_2507 (O_2507,N_24901,N_24955);
nand UO_2508 (O_2508,N_24819,N_24975);
or UO_2509 (O_2509,N_24913,N_24898);
xnor UO_2510 (O_2510,N_24879,N_24962);
and UO_2511 (O_2511,N_24888,N_24942);
and UO_2512 (O_2512,N_24982,N_24890);
nand UO_2513 (O_2513,N_24931,N_24891);
nor UO_2514 (O_2514,N_24981,N_24892);
xor UO_2515 (O_2515,N_24896,N_24825);
and UO_2516 (O_2516,N_24934,N_24923);
nor UO_2517 (O_2517,N_24974,N_24919);
xnor UO_2518 (O_2518,N_24887,N_24857);
xnor UO_2519 (O_2519,N_24937,N_24969);
and UO_2520 (O_2520,N_24806,N_24929);
and UO_2521 (O_2521,N_24819,N_24990);
and UO_2522 (O_2522,N_24823,N_24855);
or UO_2523 (O_2523,N_24919,N_24856);
nand UO_2524 (O_2524,N_24829,N_24953);
nor UO_2525 (O_2525,N_24800,N_24842);
nand UO_2526 (O_2526,N_24822,N_24913);
nand UO_2527 (O_2527,N_24809,N_24998);
or UO_2528 (O_2528,N_24987,N_24825);
nor UO_2529 (O_2529,N_24844,N_24951);
xnor UO_2530 (O_2530,N_24948,N_24960);
nor UO_2531 (O_2531,N_24809,N_24964);
nor UO_2532 (O_2532,N_24974,N_24877);
xor UO_2533 (O_2533,N_24941,N_24808);
nor UO_2534 (O_2534,N_24827,N_24926);
and UO_2535 (O_2535,N_24960,N_24886);
and UO_2536 (O_2536,N_24990,N_24826);
and UO_2537 (O_2537,N_24943,N_24938);
xnor UO_2538 (O_2538,N_24906,N_24959);
nand UO_2539 (O_2539,N_24923,N_24887);
xnor UO_2540 (O_2540,N_24997,N_24928);
or UO_2541 (O_2541,N_24907,N_24976);
xnor UO_2542 (O_2542,N_24908,N_24900);
nor UO_2543 (O_2543,N_24976,N_24958);
nand UO_2544 (O_2544,N_24907,N_24807);
and UO_2545 (O_2545,N_24908,N_24954);
and UO_2546 (O_2546,N_24993,N_24987);
xor UO_2547 (O_2547,N_24978,N_24857);
nand UO_2548 (O_2548,N_24964,N_24903);
and UO_2549 (O_2549,N_24864,N_24895);
nand UO_2550 (O_2550,N_24895,N_24886);
or UO_2551 (O_2551,N_24973,N_24988);
or UO_2552 (O_2552,N_24954,N_24813);
xor UO_2553 (O_2553,N_24988,N_24872);
xor UO_2554 (O_2554,N_24887,N_24921);
nor UO_2555 (O_2555,N_24956,N_24813);
nand UO_2556 (O_2556,N_24992,N_24829);
or UO_2557 (O_2557,N_24876,N_24821);
and UO_2558 (O_2558,N_24978,N_24905);
or UO_2559 (O_2559,N_24853,N_24958);
xnor UO_2560 (O_2560,N_24955,N_24952);
or UO_2561 (O_2561,N_24819,N_24985);
or UO_2562 (O_2562,N_24902,N_24862);
xnor UO_2563 (O_2563,N_24979,N_24974);
nor UO_2564 (O_2564,N_24955,N_24972);
nand UO_2565 (O_2565,N_24836,N_24867);
nand UO_2566 (O_2566,N_24904,N_24868);
nor UO_2567 (O_2567,N_24879,N_24965);
or UO_2568 (O_2568,N_24948,N_24804);
or UO_2569 (O_2569,N_24967,N_24949);
nand UO_2570 (O_2570,N_24889,N_24930);
or UO_2571 (O_2571,N_24844,N_24948);
and UO_2572 (O_2572,N_24836,N_24856);
and UO_2573 (O_2573,N_24894,N_24936);
nor UO_2574 (O_2574,N_24982,N_24984);
xnor UO_2575 (O_2575,N_24816,N_24873);
xor UO_2576 (O_2576,N_24897,N_24848);
and UO_2577 (O_2577,N_24827,N_24873);
nand UO_2578 (O_2578,N_24834,N_24853);
or UO_2579 (O_2579,N_24913,N_24987);
nand UO_2580 (O_2580,N_24922,N_24919);
xnor UO_2581 (O_2581,N_24956,N_24803);
xnor UO_2582 (O_2582,N_24857,N_24907);
and UO_2583 (O_2583,N_24874,N_24965);
and UO_2584 (O_2584,N_24801,N_24861);
nand UO_2585 (O_2585,N_24851,N_24958);
or UO_2586 (O_2586,N_24930,N_24940);
and UO_2587 (O_2587,N_24817,N_24918);
nand UO_2588 (O_2588,N_24882,N_24820);
nand UO_2589 (O_2589,N_24876,N_24900);
xnor UO_2590 (O_2590,N_24868,N_24971);
or UO_2591 (O_2591,N_24996,N_24979);
nand UO_2592 (O_2592,N_24809,N_24826);
and UO_2593 (O_2593,N_24915,N_24984);
or UO_2594 (O_2594,N_24912,N_24898);
and UO_2595 (O_2595,N_24920,N_24994);
xnor UO_2596 (O_2596,N_24894,N_24955);
nand UO_2597 (O_2597,N_24958,N_24812);
nand UO_2598 (O_2598,N_24915,N_24836);
nor UO_2599 (O_2599,N_24804,N_24858);
or UO_2600 (O_2600,N_24869,N_24944);
or UO_2601 (O_2601,N_24875,N_24900);
xnor UO_2602 (O_2602,N_24861,N_24922);
nand UO_2603 (O_2603,N_24964,N_24968);
nor UO_2604 (O_2604,N_24920,N_24809);
or UO_2605 (O_2605,N_24926,N_24956);
and UO_2606 (O_2606,N_24918,N_24992);
nand UO_2607 (O_2607,N_24974,N_24990);
or UO_2608 (O_2608,N_24863,N_24892);
nand UO_2609 (O_2609,N_24861,N_24963);
nand UO_2610 (O_2610,N_24801,N_24961);
and UO_2611 (O_2611,N_24954,N_24942);
nor UO_2612 (O_2612,N_24804,N_24987);
nand UO_2613 (O_2613,N_24889,N_24832);
and UO_2614 (O_2614,N_24893,N_24838);
xor UO_2615 (O_2615,N_24811,N_24922);
xor UO_2616 (O_2616,N_24813,N_24879);
nand UO_2617 (O_2617,N_24951,N_24845);
nor UO_2618 (O_2618,N_24812,N_24817);
and UO_2619 (O_2619,N_24953,N_24990);
nand UO_2620 (O_2620,N_24835,N_24987);
xnor UO_2621 (O_2621,N_24935,N_24804);
nand UO_2622 (O_2622,N_24848,N_24934);
and UO_2623 (O_2623,N_24826,N_24835);
xor UO_2624 (O_2624,N_24820,N_24905);
and UO_2625 (O_2625,N_24927,N_24871);
xor UO_2626 (O_2626,N_24912,N_24860);
xnor UO_2627 (O_2627,N_24981,N_24850);
xnor UO_2628 (O_2628,N_24821,N_24840);
xnor UO_2629 (O_2629,N_24913,N_24859);
xnor UO_2630 (O_2630,N_24870,N_24819);
xnor UO_2631 (O_2631,N_24942,N_24996);
nand UO_2632 (O_2632,N_24806,N_24967);
or UO_2633 (O_2633,N_24865,N_24809);
nor UO_2634 (O_2634,N_24869,N_24942);
nand UO_2635 (O_2635,N_24956,N_24896);
nand UO_2636 (O_2636,N_24905,N_24851);
nor UO_2637 (O_2637,N_24878,N_24805);
or UO_2638 (O_2638,N_24817,N_24985);
and UO_2639 (O_2639,N_24887,N_24813);
xor UO_2640 (O_2640,N_24806,N_24816);
or UO_2641 (O_2641,N_24869,N_24963);
or UO_2642 (O_2642,N_24966,N_24823);
xnor UO_2643 (O_2643,N_24850,N_24913);
and UO_2644 (O_2644,N_24916,N_24862);
xor UO_2645 (O_2645,N_24978,N_24935);
or UO_2646 (O_2646,N_24829,N_24946);
or UO_2647 (O_2647,N_24833,N_24823);
xor UO_2648 (O_2648,N_24920,N_24839);
and UO_2649 (O_2649,N_24968,N_24914);
nand UO_2650 (O_2650,N_24982,N_24898);
and UO_2651 (O_2651,N_24824,N_24919);
nand UO_2652 (O_2652,N_24976,N_24877);
xnor UO_2653 (O_2653,N_24853,N_24997);
nand UO_2654 (O_2654,N_24935,N_24976);
nor UO_2655 (O_2655,N_24932,N_24937);
and UO_2656 (O_2656,N_24994,N_24872);
nor UO_2657 (O_2657,N_24819,N_24942);
nor UO_2658 (O_2658,N_24899,N_24860);
and UO_2659 (O_2659,N_24941,N_24850);
and UO_2660 (O_2660,N_24967,N_24987);
xor UO_2661 (O_2661,N_24985,N_24994);
nor UO_2662 (O_2662,N_24882,N_24937);
or UO_2663 (O_2663,N_24936,N_24897);
or UO_2664 (O_2664,N_24970,N_24827);
and UO_2665 (O_2665,N_24849,N_24929);
nor UO_2666 (O_2666,N_24996,N_24809);
or UO_2667 (O_2667,N_24825,N_24890);
and UO_2668 (O_2668,N_24849,N_24932);
or UO_2669 (O_2669,N_24931,N_24988);
xnor UO_2670 (O_2670,N_24889,N_24934);
xnor UO_2671 (O_2671,N_24895,N_24832);
and UO_2672 (O_2672,N_24882,N_24850);
xnor UO_2673 (O_2673,N_24810,N_24954);
xnor UO_2674 (O_2674,N_24878,N_24812);
and UO_2675 (O_2675,N_24956,N_24856);
and UO_2676 (O_2676,N_24921,N_24882);
or UO_2677 (O_2677,N_24880,N_24976);
and UO_2678 (O_2678,N_24990,N_24926);
nor UO_2679 (O_2679,N_24854,N_24840);
nand UO_2680 (O_2680,N_24895,N_24878);
and UO_2681 (O_2681,N_24898,N_24916);
nor UO_2682 (O_2682,N_24806,N_24809);
nand UO_2683 (O_2683,N_24800,N_24996);
and UO_2684 (O_2684,N_24886,N_24828);
or UO_2685 (O_2685,N_24965,N_24827);
and UO_2686 (O_2686,N_24925,N_24901);
nor UO_2687 (O_2687,N_24934,N_24862);
and UO_2688 (O_2688,N_24989,N_24976);
and UO_2689 (O_2689,N_24984,N_24961);
or UO_2690 (O_2690,N_24936,N_24989);
or UO_2691 (O_2691,N_24987,N_24908);
xor UO_2692 (O_2692,N_24815,N_24896);
xor UO_2693 (O_2693,N_24874,N_24811);
or UO_2694 (O_2694,N_24852,N_24883);
nand UO_2695 (O_2695,N_24919,N_24994);
nand UO_2696 (O_2696,N_24801,N_24948);
and UO_2697 (O_2697,N_24822,N_24933);
and UO_2698 (O_2698,N_24854,N_24940);
or UO_2699 (O_2699,N_24897,N_24818);
or UO_2700 (O_2700,N_24922,N_24952);
or UO_2701 (O_2701,N_24962,N_24837);
xnor UO_2702 (O_2702,N_24865,N_24936);
xnor UO_2703 (O_2703,N_24962,N_24933);
xnor UO_2704 (O_2704,N_24904,N_24884);
and UO_2705 (O_2705,N_24881,N_24862);
xor UO_2706 (O_2706,N_24978,N_24854);
or UO_2707 (O_2707,N_24915,N_24881);
xnor UO_2708 (O_2708,N_24986,N_24940);
nor UO_2709 (O_2709,N_24935,N_24948);
and UO_2710 (O_2710,N_24908,N_24902);
xnor UO_2711 (O_2711,N_24801,N_24929);
nor UO_2712 (O_2712,N_24890,N_24859);
xor UO_2713 (O_2713,N_24958,N_24820);
xor UO_2714 (O_2714,N_24995,N_24810);
nand UO_2715 (O_2715,N_24962,N_24936);
nor UO_2716 (O_2716,N_24827,N_24968);
nor UO_2717 (O_2717,N_24886,N_24834);
and UO_2718 (O_2718,N_24806,N_24997);
nor UO_2719 (O_2719,N_24954,N_24859);
nor UO_2720 (O_2720,N_24987,N_24809);
and UO_2721 (O_2721,N_24854,N_24858);
and UO_2722 (O_2722,N_24820,N_24967);
xnor UO_2723 (O_2723,N_24831,N_24826);
xnor UO_2724 (O_2724,N_24805,N_24832);
and UO_2725 (O_2725,N_24831,N_24887);
xnor UO_2726 (O_2726,N_24884,N_24809);
nor UO_2727 (O_2727,N_24822,N_24843);
nor UO_2728 (O_2728,N_24972,N_24989);
nand UO_2729 (O_2729,N_24813,N_24818);
nor UO_2730 (O_2730,N_24804,N_24894);
xor UO_2731 (O_2731,N_24892,N_24813);
nand UO_2732 (O_2732,N_24850,N_24848);
nand UO_2733 (O_2733,N_24835,N_24959);
xnor UO_2734 (O_2734,N_24908,N_24970);
xor UO_2735 (O_2735,N_24851,N_24910);
and UO_2736 (O_2736,N_24867,N_24813);
or UO_2737 (O_2737,N_24936,N_24910);
or UO_2738 (O_2738,N_24910,N_24823);
nand UO_2739 (O_2739,N_24958,N_24843);
nor UO_2740 (O_2740,N_24909,N_24810);
or UO_2741 (O_2741,N_24929,N_24892);
or UO_2742 (O_2742,N_24927,N_24814);
nand UO_2743 (O_2743,N_24807,N_24803);
and UO_2744 (O_2744,N_24993,N_24988);
xnor UO_2745 (O_2745,N_24846,N_24963);
and UO_2746 (O_2746,N_24935,N_24888);
and UO_2747 (O_2747,N_24955,N_24926);
nand UO_2748 (O_2748,N_24834,N_24889);
or UO_2749 (O_2749,N_24847,N_24856);
xor UO_2750 (O_2750,N_24991,N_24890);
or UO_2751 (O_2751,N_24952,N_24847);
nor UO_2752 (O_2752,N_24928,N_24916);
nor UO_2753 (O_2753,N_24998,N_24904);
nor UO_2754 (O_2754,N_24986,N_24883);
xnor UO_2755 (O_2755,N_24978,N_24853);
and UO_2756 (O_2756,N_24950,N_24898);
xor UO_2757 (O_2757,N_24844,N_24820);
and UO_2758 (O_2758,N_24928,N_24965);
nand UO_2759 (O_2759,N_24973,N_24981);
nor UO_2760 (O_2760,N_24937,N_24913);
nand UO_2761 (O_2761,N_24816,N_24855);
and UO_2762 (O_2762,N_24969,N_24862);
nand UO_2763 (O_2763,N_24859,N_24882);
xor UO_2764 (O_2764,N_24838,N_24968);
nand UO_2765 (O_2765,N_24830,N_24901);
or UO_2766 (O_2766,N_24813,N_24866);
nor UO_2767 (O_2767,N_24922,N_24978);
and UO_2768 (O_2768,N_24860,N_24843);
nor UO_2769 (O_2769,N_24861,N_24816);
or UO_2770 (O_2770,N_24877,N_24819);
xnor UO_2771 (O_2771,N_24984,N_24967);
or UO_2772 (O_2772,N_24969,N_24816);
nor UO_2773 (O_2773,N_24907,N_24869);
and UO_2774 (O_2774,N_24944,N_24845);
xnor UO_2775 (O_2775,N_24943,N_24947);
or UO_2776 (O_2776,N_24866,N_24896);
and UO_2777 (O_2777,N_24873,N_24948);
or UO_2778 (O_2778,N_24851,N_24936);
nand UO_2779 (O_2779,N_24895,N_24964);
nand UO_2780 (O_2780,N_24956,N_24872);
nor UO_2781 (O_2781,N_24974,N_24887);
nand UO_2782 (O_2782,N_24964,N_24818);
or UO_2783 (O_2783,N_24849,N_24920);
nor UO_2784 (O_2784,N_24961,N_24955);
or UO_2785 (O_2785,N_24954,N_24916);
nor UO_2786 (O_2786,N_24955,N_24925);
nand UO_2787 (O_2787,N_24969,N_24836);
xor UO_2788 (O_2788,N_24873,N_24941);
nor UO_2789 (O_2789,N_24976,N_24980);
nand UO_2790 (O_2790,N_24888,N_24994);
nor UO_2791 (O_2791,N_24916,N_24966);
xnor UO_2792 (O_2792,N_24818,N_24841);
xor UO_2793 (O_2793,N_24958,N_24910);
and UO_2794 (O_2794,N_24952,N_24959);
and UO_2795 (O_2795,N_24961,N_24994);
nor UO_2796 (O_2796,N_24863,N_24978);
xor UO_2797 (O_2797,N_24871,N_24986);
and UO_2798 (O_2798,N_24917,N_24938);
or UO_2799 (O_2799,N_24828,N_24902);
nand UO_2800 (O_2800,N_24954,N_24988);
xnor UO_2801 (O_2801,N_24864,N_24834);
xor UO_2802 (O_2802,N_24995,N_24824);
and UO_2803 (O_2803,N_24816,N_24928);
nand UO_2804 (O_2804,N_24862,N_24876);
or UO_2805 (O_2805,N_24832,N_24936);
xnor UO_2806 (O_2806,N_24955,N_24848);
or UO_2807 (O_2807,N_24801,N_24990);
or UO_2808 (O_2808,N_24911,N_24852);
or UO_2809 (O_2809,N_24875,N_24805);
nor UO_2810 (O_2810,N_24843,N_24832);
or UO_2811 (O_2811,N_24904,N_24973);
and UO_2812 (O_2812,N_24894,N_24833);
nor UO_2813 (O_2813,N_24908,N_24834);
or UO_2814 (O_2814,N_24957,N_24908);
xor UO_2815 (O_2815,N_24902,N_24920);
nand UO_2816 (O_2816,N_24841,N_24978);
nor UO_2817 (O_2817,N_24991,N_24986);
nand UO_2818 (O_2818,N_24855,N_24915);
xnor UO_2819 (O_2819,N_24953,N_24912);
nor UO_2820 (O_2820,N_24935,N_24972);
or UO_2821 (O_2821,N_24999,N_24956);
nor UO_2822 (O_2822,N_24848,N_24966);
or UO_2823 (O_2823,N_24858,N_24836);
or UO_2824 (O_2824,N_24848,N_24886);
or UO_2825 (O_2825,N_24994,N_24909);
nand UO_2826 (O_2826,N_24915,N_24923);
and UO_2827 (O_2827,N_24943,N_24898);
xnor UO_2828 (O_2828,N_24808,N_24866);
or UO_2829 (O_2829,N_24911,N_24902);
nand UO_2830 (O_2830,N_24878,N_24801);
or UO_2831 (O_2831,N_24860,N_24995);
xor UO_2832 (O_2832,N_24891,N_24962);
xnor UO_2833 (O_2833,N_24854,N_24819);
and UO_2834 (O_2834,N_24959,N_24891);
xnor UO_2835 (O_2835,N_24886,N_24985);
nand UO_2836 (O_2836,N_24918,N_24911);
and UO_2837 (O_2837,N_24857,N_24822);
and UO_2838 (O_2838,N_24808,N_24860);
xor UO_2839 (O_2839,N_24862,N_24870);
or UO_2840 (O_2840,N_24888,N_24957);
and UO_2841 (O_2841,N_24954,N_24835);
xnor UO_2842 (O_2842,N_24849,N_24941);
nor UO_2843 (O_2843,N_24854,N_24874);
or UO_2844 (O_2844,N_24944,N_24887);
nor UO_2845 (O_2845,N_24827,N_24946);
and UO_2846 (O_2846,N_24949,N_24996);
xor UO_2847 (O_2847,N_24987,N_24818);
nor UO_2848 (O_2848,N_24834,N_24888);
nor UO_2849 (O_2849,N_24827,N_24868);
xor UO_2850 (O_2850,N_24997,N_24941);
xnor UO_2851 (O_2851,N_24806,N_24805);
or UO_2852 (O_2852,N_24943,N_24963);
nor UO_2853 (O_2853,N_24886,N_24864);
nor UO_2854 (O_2854,N_24995,N_24885);
xnor UO_2855 (O_2855,N_24987,N_24969);
nor UO_2856 (O_2856,N_24978,N_24953);
nor UO_2857 (O_2857,N_24887,N_24919);
or UO_2858 (O_2858,N_24867,N_24806);
nor UO_2859 (O_2859,N_24966,N_24906);
nor UO_2860 (O_2860,N_24839,N_24932);
nand UO_2861 (O_2861,N_24966,N_24807);
nor UO_2862 (O_2862,N_24985,N_24970);
xnor UO_2863 (O_2863,N_24975,N_24976);
or UO_2864 (O_2864,N_24844,N_24845);
nand UO_2865 (O_2865,N_24932,N_24925);
and UO_2866 (O_2866,N_24974,N_24870);
and UO_2867 (O_2867,N_24931,N_24879);
nor UO_2868 (O_2868,N_24904,N_24982);
or UO_2869 (O_2869,N_24908,N_24852);
nand UO_2870 (O_2870,N_24801,N_24851);
xnor UO_2871 (O_2871,N_24952,N_24891);
or UO_2872 (O_2872,N_24832,N_24842);
or UO_2873 (O_2873,N_24867,N_24968);
and UO_2874 (O_2874,N_24894,N_24967);
or UO_2875 (O_2875,N_24850,N_24931);
xnor UO_2876 (O_2876,N_24878,N_24888);
nand UO_2877 (O_2877,N_24909,N_24927);
nand UO_2878 (O_2878,N_24999,N_24878);
and UO_2879 (O_2879,N_24996,N_24919);
or UO_2880 (O_2880,N_24975,N_24960);
and UO_2881 (O_2881,N_24871,N_24993);
nor UO_2882 (O_2882,N_24816,N_24987);
or UO_2883 (O_2883,N_24928,N_24953);
nand UO_2884 (O_2884,N_24936,N_24980);
nand UO_2885 (O_2885,N_24831,N_24925);
and UO_2886 (O_2886,N_24955,N_24992);
xor UO_2887 (O_2887,N_24845,N_24999);
nor UO_2888 (O_2888,N_24895,N_24949);
xnor UO_2889 (O_2889,N_24932,N_24989);
and UO_2890 (O_2890,N_24912,N_24961);
and UO_2891 (O_2891,N_24845,N_24882);
and UO_2892 (O_2892,N_24943,N_24990);
or UO_2893 (O_2893,N_24883,N_24848);
xnor UO_2894 (O_2894,N_24813,N_24902);
or UO_2895 (O_2895,N_24948,N_24906);
and UO_2896 (O_2896,N_24840,N_24899);
xor UO_2897 (O_2897,N_24842,N_24903);
xor UO_2898 (O_2898,N_24814,N_24872);
and UO_2899 (O_2899,N_24867,N_24912);
or UO_2900 (O_2900,N_24832,N_24800);
or UO_2901 (O_2901,N_24914,N_24852);
xnor UO_2902 (O_2902,N_24836,N_24954);
nor UO_2903 (O_2903,N_24999,N_24973);
or UO_2904 (O_2904,N_24907,N_24828);
nor UO_2905 (O_2905,N_24800,N_24967);
and UO_2906 (O_2906,N_24895,N_24900);
and UO_2907 (O_2907,N_24813,N_24941);
nor UO_2908 (O_2908,N_24872,N_24833);
nor UO_2909 (O_2909,N_24987,N_24991);
nand UO_2910 (O_2910,N_24993,N_24847);
xor UO_2911 (O_2911,N_24930,N_24846);
and UO_2912 (O_2912,N_24820,N_24951);
xnor UO_2913 (O_2913,N_24839,N_24878);
nor UO_2914 (O_2914,N_24988,N_24895);
and UO_2915 (O_2915,N_24837,N_24875);
xnor UO_2916 (O_2916,N_24933,N_24827);
and UO_2917 (O_2917,N_24945,N_24858);
nor UO_2918 (O_2918,N_24952,N_24963);
xor UO_2919 (O_2919,N_24917,N_24967);
and UO_2920 (O_2920,N_24829,N_24886);
nor UO_2921 (O_2921,N_24896,N_24883);
or UO_2922 (O_2922,N_24932,N_24992);
xor UO_2923 (O_2923,N_24974,N_24872);
nor UO_2924 (O_2924,N_24816,N_24995);
xor UO_2925 (O_2925,N_24858,N_24939);
or UO_2926 (O_2926,N_24929,N_24858);
xnor UO_2927 (O_2927,N_24887,N_24829);
xor UO_2928 (O_2928,N_24847,N_24893);
or UO_2929 (O_2929,N_24906,N_24963);
nand UO_2930 (O_2930,N_24801,N_24922);
nor UO_2931 (O_2931,N_24871,N_24828);
or UO_2932 (O_2932,N_24806,N_24857);
nor UO_2933 (O_2933,N_24988,N_24942);
nor UO_2934 (O_2934,N_24939,N_24897);
nand UO_2935 (O_2935,N_24977,N_24878);
xnor UO_2936 (O_2936,N_24867,N_24990);
nor UO_2937 (O_2937,N_24874,N_24917);
or UO_2938 (O_2938,N_24880,N_24823);
xor UO_2939 (O_2939,N_24869,N_24874);
and UO_2940 (O_2940,N_24904,N_24826);
nor UO_2941 (O_2941,N_24860,N_24812);
xor UO_2942 (O_2942,N_24908,N_24955);
xnor UO_2943 (O_2943,N_24877,N_24935);
nor UO_2944 (O_2944,N_24947,N_24949);
nor UO_2945 (O_2945,N_24951,N_24833);
xor UO_2946 (O_2946,N_24992,N_24827);
xor UO_2947 (O_2947,N_24912,N_24801);
or UO_2948 (O_2948,N_24879,N_24961);
and UO_2949 (O_2949,N_24819,N_24837);
nor UO_2950 (O_2950,N_24891,N_24948);
or UO_2951 (O_2951,N_24832,N_24976);
nor UO_2952 (O_2952,N_24950,N_24894);
xnor UO_2953 (O_2953,N_24960,N_24951);
nand UO_2954 (O_2954,N_24823,N_24942);
nor UO_2955 (O_2955,N_24843,N_24948);
and UO_2956 (O_2956,N_24852,N_24851);
or UO_2957 (O_2957,N_24902,N_24969);
nor UO_2958 (O_2958,N_24814,N_24898);
and UO_2959 (O_2959,N_24841,N_24956);
nor UO_2960 (O_2960,N_24951,N_24996);
xor UO_2961 (O_2961,N_24894,N_24867);
and UO_2962 (O_2962,N_24830,N_24982);
nor UO_2963 (O_2963,N_24838,N_24871);
or UO_2964 (O_2964,N_24955,N_24861);
or UO_2965 (O_2965,N_24993,N_24974);
nand UO_2966 (O_2966,N_24977,N_24861);
or UO_2967 (O_2967,N_24894,N_24883);
nand UO_2968 (O_2968,N_24939,N_24801);
and UO_2969 (O_2969,N_24897,N_24865);
xor UO_2970 (O_2970,N_24922,N_24824);
nor UO_2971 (O_2971,N_24918,N_24946);
xor UO_2972 (O_2972,N_24995,N_24888);
nand UO_2973 (O_2973,N_24993,N_24888);
nor UO_2974 (O_2974,N_24919,N_24874);
and UO_2975 (O_2975,N_24920,N_24999);
or UO_2976 (O_2976,N_24904,N_24886);
or UO_2977 (O_2977,N_24803,N_24833);
xnor UO_2978 (O_2978,N_24943,N_24919);
and UO_2979 (O_2979,N_24987,N_24808);
nand UO_2980 (O_2980,N_24960,N_24835);
xor UO_2981 (O_2981,N_24883,N_24857);
nand UO_2982 (O_2982,N_24929,N_24840);
nand UO_2983 (O_2983,N_24891,N_24949);
xnor UO_2984 (O_2984,N_24802,N_24946);
or UO_2985 (O_2985,N_24995,N_24959);
and UO_2986 (O_2986,N_24976,N_24919);
nor UO_2987 (O_2987,N_24960,N_24852);
and UO_2988 (O_2988,N_24883,N_24963);
nand UO_2989 (O_2989,N_24955,N_24864);
or UO_2990 (O_2990,N_24821,N_24988);
nand UO_2991 (O_2991,N_24859,N_24961);
nand UO_2992 (O_2992,N_24812,N_24889);
xor UO_2993 (O_2993,N_24868,N_24952);
xnor UO_2994 (O_2994,N_24915,N_24968);
nor UO_2995 (O_2995,N_24955,N_24931);
xnor UO_2996 (O_2996,N_24849,N_24936);
or UO_2997 (O_2997,N_24966,N_24907);
and UO_2998 (O_2998,N_24882,N_24916);
xor UO_2999 (O_2999,N_24980,N_24983);
endmodule