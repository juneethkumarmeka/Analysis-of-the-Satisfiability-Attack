module basic_2500_25000_3000_20_levels_10xor_2(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999;
xor U0 (N_0,In_1778,In_662);
xor U1 (N_1,In_2341,In_65);
nor U2 (N_2,In_1284,In_962);
nand U3 (N_3,In_1761,In_1106);
and U4 (N_4,In_1909,In_1637);
and U5 (N_5,In_1964,In_194);
or U6 (N_6,In_1129,In_355);
or U7 (N_7,In_1562,In_1880);
nand U8 (N_8,In_439,In_1628);
nor U9 (N_9,In_1704,In_2111);
and U10 (N_10,In_336,In_1591);
nand U11 (N_11,In_263,In_786);
xnor U12 (N_12,In_1169,In_1563);
nor U13 (N_13,In_867,In_935);
and U14 (N_14,In_1159,In_1400);
or U15 (N_15,In_237,In_1745);
and U16 (N_16,In_408,In_345);
or U17 (N_17,In_1448,In_1464);
nand U18 (N_18,In_1500,In_2431);
and U19 (N_19,In_1933,In_1269);
xor U20 (N_20,In_2295,In_1127);
xor U21 (N_21,In_857,In_1101);
and U22 (N_22,In_1438,In_2458);
nand U23 (N_23,In_1249,In_1221);
or U24 (N_24,In_1139,In_2224);
nor U25 (N_25,In_1904,In_24);
nor U26 (N_26,In_2070,In_520);
xor U27 (N_27,In_729,In_1777);
nor U28 (N_28,In_2119,In_1455);
or U29 (N_29,In_2232,In_290);
nor U30 (N_30,In_66,In_1007);
and U31 (N_31,In_1929,In_721);
nor U32 (N_32,In_278,In_2491);
nand U33 (N_33,In_391,In_584);
or U34 (N_34,In_1168,In_339);
xnor U35 (N_35,In_1160,In_1944);
nand U36 (N_36,In_2275,In_777);
nand U37 (N_37,In_2439,In_2195);
and U38 (N_38,In_310,In_252);
nor U39 (N_39,In_2371,In_2261);
nor U40 (N_40,In_1362,In_970);
nor U41 (N_41,In_1517,In_2221);
or U42 (N_42,In_23,In_2060);
nor U43 (N_43,In_1478,In_2114);
nor U44 (N_44,In_872,In_977);
nand U45 (N_45,In_1877,In_453);
nand U46 (N_46,In_1152,In_1112);
nor U47 (N_47,In_2397,In_576);
nor U48 (N_48,In_5,In_557);
nand U49 (N_49,In_1411,In_553);
and U50 (N_50,In_994,In_653);
and U51 (N_51,In_2100,In_80);
and U52 (N_52,In_657,In_1285);
nor U53 (N_53,In_578,In_154);
and U54 (N_54,In_812,In_2250);
nand U55 (N_55,In_1385,In_849);
nand U56 (N_56,In_1370,In_2426);
nor U57 (N_57,In_1542,In_1228);
and U58 (N_58,In_192,In_1807);
nand U59 (N_59,In_1241,In_1739);
xnor U60 (N_60,In_205,In_1670);
or U61 (N_61,In_846,In_602);
and U62 (N_62,In_100,In_146);
xor U63 (N_63,In_1075,In_990);
or U64 (N_64,In_538,In_1688);
xnor U65 (N_65,In_257,In_1884);
and U66 (N_66,In_2363,In_1656);
xnor U67 (N_67,In_987,In_363);
and U68 (N_68,In_1389,In_991);
xor U69 (N_69,In_556,In_2131);
and U70 (N_70,In_1328,In_2139);
or U71 (N_71,In_591,In_2023);
nor U72 (N_72,In_2302,In_879);
xnor U73 (N_73,In_181,In_684);
xor U74 (N_74,In_717,In_1900);
nor U75 (N_75,In_212,In_648);
or U76 (N_76,In_1133,In_1749);
or U77 (N_77,In_2018,In_546);
xnor U78 (N_78,In_905,In_384);
xnor U79 (N_79,In_1118,In_2094);
and U80 (N_80,In_601,In_2087);
nand U81 (N_81,In_1427,In_2078);
and U82 (N_82,In_796,In_81);
xnor U83 (N_83,In_534,In_2036);
nor U84 (N_84,In_1769,In_2047);
or U85 (N_85,In_829,In_1987);
and U86 (N_86,In_280,In_1374);
nand U87 (N_87,In_652,In_1816);
nand U88 (N_88,In_1108,In_1282);
nor U89 (N_89,In_389,In_1658);
or U90 (N_90,In_2409,In_2487);
nand U91 (N_91,In_2482,In_965);
nand U92 (N_92,In_90,In_417);
nand U93 (N_93,In_2488,In_288);
or U94 (N_94,In_1805,In_833);
and U95 (N_95,In_701,In_1050);
nor U96 (N_96,In_2156,In_2404);
nand U97 (N_97,In_1376,In_210);
and U98 (N_98,In_1371,In_2374);
or U99 (N_99,In_1222,In_1206);
nand U100 (N_100,In_824,In_2313);
or U101 (N_101,In_2142,In_744);
and U102 (N_102,In_929,In_455);
xnor U103 (N_103,In_1892,In_2057);
nor U104 (N_104,In_113,In_1463);
nand U105 (N_105,In_1086,In_2237);
xnor U106 (N_106,In_2218,In_2126);
and U107 (N_107,In_2005,In_513);
nor U108 (N_108,In_2138,In_2186);
xnor U109 (N_109,In_2266,In_815);
xnor U110 (N_110,In_2495,In_393);
or U111 (N_111,In_1010,In_886);
or U112 (N_112,In_1194,In_1996);
xnor U113 (N_113,In_742,In_55);
nor U114 (N_114,In_600,In_569);
xnor U115 (N_115,In_1103,In_1839);
nor U116 (N_116,In_197,In_1028);
and U117 (N_117,In_2219,In_1941);
nand U118 (N_118,In_1396,In_1035);
and U119 (N_119,In_1236,In_2205);
nor U120 (N_120,In_835,In_1496);
or U121 (N_121,In_82,In_972);
xor U122 (N_122,In_890,In_2164);
or U123 (N_123,In_1685,In_604);
nand U124 (N_124,In_826,In_172);
xor U125 (N_125,In_531,In_1617);
and U126 (N_126,In_873,In_2115);
xnor U127 (N_127,In_685,In_162);
nand U128 (N_128,In_70,In_2231);
or U129 (N_129,In_667,In_322);
and U130 (N_130,In_64,In_1943);
and U131 (N_131,In_409,In_1669);
nor U132 (N_132,In_765,In_341);
or U133 (N_133,In_1981,In_1363);
nand U134 (N_134,In_2473,In_2103);
xnor U135 (N_135,In_2107,In_2062);
xnor U136 (N_136,In_878,In_416);
and U137 (N_137,In_543,In_1758);
and U138 (N_138,In_1247,In_1196);
or U139 (N_139,In_1589,In_2441);
nor U140 (N_140,In_2498,In_1032);
xnor U141 (N_141,In_2386,In_2073);
xnor U142 (N_142,In_2067,In_1360);
xor U143 (N_143,In_1042,In_1504);
nand U144 (N_144,In_309,In_1104);
nor U145 (N_145,In_1992,In_1567);
xnor U146 (N_146,In_883,In_1163);
and U147 (N_147,In_2134,In_1862);
nand U148 (N_148,In_2181,In_992);
and U149 (N_149,In_1216,In_1110);
nor U150 (N_150,In_289,In_49);
nand U151 (N_151,In_858,In_784);
and U152 (N_152,In_974,In_319);
nand U153 (N_153,In_1131,In_1339);
or U154 (N_154,In_620,In_2273);
xor U155 (N_155,In_679,In_157);
or U156 (N_156,In_775,In_810);
and U157 (N_157,In_13,In_752);
xor U158 (N_158,In_1970,In_1458);
or U159 (N_159,In_2442,In_735);
nand U160 (N_160,In_1490,In_1969);
xnor U161 (N_161,In_2333,In_1938);
or U162 (N_162,In_267,In_1838);
xor U163 (N_163,In_549,In_1219);
nand U164 (N_164,In_759,In_2388);
or U165 (N_165,In_1314,In_1395);
nand U166 (N_166,In_1025,In_1533);
or U167 (N_167,In_1198,In_1979);
or U168 (N_168,In_1599,In_2197);
nor U169 (N_169,In_1757,In_827);
and U170 (N_170,In_2296,In_2343);
xnor U171 (N_171,In_1336,In_19);
or U172 (N_172,In_1803,In_868);
and U173 (N_173,In_1728,In_2058);
or U174 (N_174,In_2172,In_1509);
nand U175 (N_175,In_1058,In_1819);
xnor U176 (N_176,In_2497,In_1232);
and U177 (N_177,In_1326,In_351);
xnor U178 (N_178,In_1207,In_4);
nand U179 (N_179,In_1356,In_152);
nor U180 (N_180,In_1650,In_2130);
nand U181 (N_181,In_559,In_344);
nand U182 (N_182,In_2116,In_1940);
nor U183 (N_183,In_818,In_1802);
and U184 (N_184,In_140,In_2469);
nor U185 (N_185,In_733,In_921);
nand U186 (N_186,In_424,In_581);
nor U187 (N_187,In_1633,In_898);
nand U188 (N_188,In_508,In_2207);
nor U189 (N_189,In_2427,In_816);
nand U190 (N_190,In_1053,In_1796);
nor U191 (N_191,In_2064,In_2148);
or U192 (N_192,In_218,In_201);
nand U193 (N_193,In_1917,In_594);
and U194 (N_194,In_919,In_297);
xnor U195 (N_195,In_1432,In_1452);
nand U196 (N_196,In_1850,In_60);
xnor U197 (N_197,In_1782,In_1716);
nor U198 (N_198,In_605,In_2489);
nand U199 (N_199,In_2365,In_61);
xor U200 (N_200,In_1717,In_97);
xor U201 (N_201,In_422,In_2381);
nor U202 (N_202,In_515,In_799);
nand U203 (N_203,In_1597,In_2408);
nor U204 (N_204,In_564,In_1664);
nand U205 (N_205,In_2001,In_894);
nand U206 (N_206,In_798,In_33);
xor U207 (N_207,In_967,In_1864);
xnor U208 (N_208,In_133,In_516);
nor U209 (N_209,In_483,In_956);
and U210 (N_210,In_170,In_1180);
nand U211 (N_211,In_1183,In_188);
nor U212 (N_212,In_1623,In_362);
or U213 (N_213,In_320,In_1492);
xnor U214 (N_214,In_683,In_1199);
or U215 (N_215,In_2149,In_1566);
or U216 (N_216,In_1056,In_940);
nand U217 (N_217,In_907,In_1995);
nand U218 (N_218,In_7,In_2213);
and U219 (N_219,In_2081,In_1191);
and U220 (N_220,In_1896,In_1690);
and U221 (N_221,In_2271,In_1883);
and U222 (N_222,In_1378,In_2117);
or U223 (N_223,In_704,In_327);
xnor U224 (N_224,In_877,In_2453);
nand U225 (N_225,In_762,In_1308);
xor U226 (N_226,In_839,In_1188);
xor U227 (N_227,In_610,In_2288);
nor U228 (N_228,In_2285,In_817);
xor U229 (N_229,In_723,In_2272);
or U230 (N_230,In_769,In_85);
xnor U231 (N_231,In_782,In_1470);
or U232 (N_232,In_893,In_828);
nand U233 (N_233,In_423,In_1618);
nor U234 (N_234,In_1565,In_187);
nand U235 (N_235,In_388,In_880);
and U236 (N_236,In_213,In_2038);
or U237 (N_237,In_1668,In_1730);
xnor U238 (N_238,In_30,In_2318);
or U239 (N_239,In_674,In_1034);
or U240 (N_240,In_2444,In_1136);
or U241 (N_241,In_1854,In_1806);
nand U242 (N_242,In_1430,In_756);
xnor U243 (N_243,In_2118,In_2278);
nand U244 (N_244,In_533,In_1057);
nand U245 (N_245,In_1868,In_1384);
xnor U246 (N_246,In_1005,In_1123);
nand U247 (N_247,In_681,In_896);
nor U248 (N_248,In_1203,In_1972);
nor U249 (N_249,In_635,In_440);
nor U250 (N_250,In_1538,In_1172);
nand U251 (N_251,In_1751,In_242);
nor U252 (N_252,In_1810,In_1397);
nor U253 (N_253,In_270,In_2369);
nand U254 (N_254,In_902,In_323);
or U255 (N_255,In_2359,In_2144);
nand U256 (N_256,In_1093,In_1887);
and U257 (N_257,In_1238,In_1000);
or U258 (N_258,In_1218,In_2243);
or U259 (N_259,In_2021,In_778);
xnor U260 (N_260,In_670,In_156);
nand U261 (N_261,In_2088,In_63);
nor U262 (N_262,In_764,In_1606);
nor U263 (N_263,In_220,In_1765);
and U264 (N_264,In_1684,In_1324);
xor U265 (N_265,In_1155,In_56);
xor U266 (N_266,In_2464,In_224);
nand U267 (N_267,In_1079,In_2249);
or U268 (N_268,In_2112,In_1754);
and U269 (N_269,In_1310,In_595);
nand U270 (N_270,In_328,In_1318);
nand U271 (N_271,In_1347,In_2419);
nor U272 (N_272,In_2183,In_738);
nand U273 (N_273,In_1535,In_1632);
xnor U274 (N_274,In_971,In_1230);
nand U275 (N_275,In_266,In_16);
or U276 (N_276,In_228,In_2228);
or U277 (N_277,In_2289,In_1164);
or U278 (N_278,In_1487,In_1655);
nand U279 (N_279,In_1901,In_1962);
nand U280 (N_280,In_2099,In_1425);
nand U281 (N_281,In_1192,In_1069);
xnor U282 (N_282,In_656,In_1920);
and U283 (N_283,In_689,In_438);
and U284 (N_284,In_36,In_1620);
nor U285 (N_285,In_1026,In_359);
or U286 (N_286,In_273,In_1274);
or U287 (N_287,In_813,In_86);
nand U288 (N_288,In_2242,In_617);
or U289 (N_289,In_1298,In_925);
and U290 (N_290,In_748,In_2351);
or U291 (N_291,In_128,In_1726);
nor U292 (N_292,In_2493,In_2010);
xnor U293 (N_293,In_1811,In_589);
nor U294 (N_294,In_1999,In_1840);
and U295 (N_295,In_514,In_2043);
nand U296 (N_296,In_1762,In_161);
nand U297 (N_297,In_997,In_2072);
nand U298 (N_298,In_1342,In_561);
or U299 (N_299,In_2347,In_1878);
nor U300 (N_300,In_523,In_1270);
and U301 (N_301,In_135,In_2178);
or U302 (N_302,In_2483,In_2028);
xnor U303 (N_303,In_367,In_2367);
and U304 (N_304,In_1063,In_1644);
nand U305 (N_305,In_2122,In_727);
nand U306 (N_306,In_1844,In_803);
nand U307 (N_307,In_1609,In_2480);
nor U308 (N_308,In_209,In_1781);
and U309 (N_309,In_509,In_1706);
xor U310 (N_310,In_1516,In_1442);
or U311 (N_311,In_924,In_655);
or U312 (N_312,In_415,In_845);
nand U313 (N_313,In_261,In_1952);
or U314 (N_314,In_2410,In_562);
nand U315 (N_315,In_1067,In_2074);
or U316 (N_316,In_1624,In_457);
and U317 (N_317,In_2189,In_1150);
nand U318 (N_318,In_183,In_1647);
nor U319 (N_319,In_1399,In_1939);
and U320 (N_320,In_1872,In_1860);
nor U321 (N_321,In_969,In_91);
nor U322 (N_322,In_22,In_420);
nor U323 (N_323,In_1209,In_943);
and U324 (N_324,In_1404,In_214);
nand U325 (N_325,In_1636,In_163);
nor U326 (N_326,In_2354,In_195);
nor U327 (N_327,In_1794,In_691);
nand U328 (N_328,In_2214,In_1259);
and U329 (N_329,In_612,In_1189);
nor U330 (N_330,In_47,In_2332);
xnor U331 (N_331,In_258,In_2226);
nor U332 (N_332,In_2400,In_2405);
nand U333 (N_333,In_2246,In_2097);
nor U334 (N_334,In_1994,In_491);
xor U335 (N_335,In_1662,In_2436);
or U336 (N_336,In_848,In_2317);
or U337 (N_337,In_1175,In_481);
or U338 (N_338,In_521,In_2108);
or U339 (N_339,In_1649,In_1213);
and U340 (N_340,In_1916,In_1898);
and U341 (N_341,In_1935,In_148);
and U342 (N_342,In_2192,In_206);
xnor U343 (N_343,In_2206,In_216);
nor U344 (N_344,In_2314,In_716);
nor U345 (N_345,In_1531,In_1581);
xor U346 (N_346,In_805,In_1611);
xor U347 (N_347,In_1895,In_2339);
and U348 (N_348,In_732,In_1697);
nand U349 (N_349,In_2358,In_1435);
nor U350 (N_350,In_1253,In_486);
xor U351 (N_351,In_0,In_1923);
xor U352 (N_352,In_1262,In_1708);
and U353 (N_353,In_1248,In_1252);
nand U354 (N_354,In_467,In_229);
and U355 (N_355,In_1528,In_1666);
nor U356 (N_356,In_767,In_947);
nand U357 (N_357,In_2485,In_772);
and U358 (N_358,In_144,In_1294);
nor U359 (N_359,In_1381,In_1640);
xor U360 (N_360,In_301,In_11);
xor U361 (N_361,In_1526,In_1096);
or U362 (N_362,In_1109,In_314);
or U363 (N_363,In_1445,In_948);
and U364 (N_364,In_286,In_1020);
nor U365 (N_365,In_2040,In_62);
nor U366 (N_366,In_522,In_413);
nor U367 (N_367,In_2159,In_2398);
xor U368 (N_368,In_1608,In_277);
or U369 (N_369,In_1315,In_1122);
and U370 (N_370,In_2198,In_1398);
xnor U371 (N_371,In_1718,In_1922);
xor U372 (N_372,In_2075,In_1066);
nand U373 (N_373,In_882,In_2236);
nor U374 (N_374,In_390,In_136);
and U375 (N_375,In_2356,In_1379);
nand U376 (N_376,In_773,In_599);
xnor U377 (N_377,In_1468,In_1755);
nand U378 (N_378,In_386,In_809);
nand U379 (N_379,In_1855,In_1369);
and U380 (N_380,In_186,In_2287);
xnor U381 (N_381,In_532,In_1295);
and U382 (N_382,In_1515,In_302);
nand U383 (N_383,In_2168,In_139);
xor U384 (N_384,In_198,In_1804);
and U385 (N_385,In_1661,In_939);
xor U386 (N_386,In_2492,In_99);
and U387 (N_387,In_1424,In_527);
xnor U388 (N_388,In_2327,In_1539);
nor U389 (N_389,In_1202,In_215);
and U390 (N_390,In_1120,In_2412);
nand U391 (N_391,In_1217,In_2234);
or U392 (N_392,In_2022,In_2494);
nor U393 (N_393,In_2422,In_2027);
nor U394 (N_394,In_1338,In_1276);
or U395 (N_395,In_219,In_1553);
xnor U396 (N_396,In_1419,In_927);
nor U397 (N_397,In_671,In_1601);
and U398 (N_398,In_844,In_1467);
nand U399 (N_399,In_615,In_1946);
nor U400 (N_400,In_1639,In_294);
xor U401 (N_401,In_1712,In_519);
nand U402 (N_402,In_1866,In_524);
nand U403 (N_403,In_430,In_1520);
nor U404 (N_404,In_1030,In_2437);
nor U405 (N_405,In_1290,In_757);
nand U406 (N_406,In_2101,In_1186);
or U407 (N_407,In_641,In_920);
nor U408 (N_408,In_654,In_547);
nor U409 (N_409,In_118,In_1141);
and U410 (N_410,In_2190,In_1317);
nor U411 (N_411,In_986,In_1653);
xnor U412 (N_412,In_1791,In_165);
xnor U413 (N_413,In_2335,In_1821);
and U414 (N_414,In_1257,In_1142);
and U415 (N_415,In_177,In_895);
nand U416 (N_416,In_293,In_1214);
and U417 (N_417,In_903,In_495);
and U418 (N_418,In_1681,In_1388);
and U419 (N_419,In_1125,In_143);
nand U420 (N_420,In_1720,In_517);
xnor U421 (N_421,In_1078,In_1631);
and U422 (N_422,In_2415,In_851);
xnor U423 (N_423,In_1166,In_1978);
and U424 (N_424,In_565,In_381);
or U425 (N_425,In_73,In_2484);
or U426 (N_426,In_650,In_1277);
xnor U427 (N_427,In_1018,In_2257);
or U428 (N_428,In_1475,In_2110);
and U429 (N_429,In_1140,In_1557);
xor U430 (N_430,In_2269,In_1540);
nor U431 (N_431,In_260,In_292);
and U432 (N_432,In_1071,In_2476);
nor U433 (N_433,In_1393,In_499);
or U434 (N_434,In_1911,In_2037);
nor U435 (N_435,In_387,In_6);
nand U436 (N_436,In_542,In_505);
nand U437 (N_437,In_855,In_484);
or U438 (N_438,In_1431,In_477);
nand U439 (N_439,In_256,In_2032);
nor U440 (N_440,In_1503,In_837);
nand U441 (N_441,In_2392,In_665);
or U442 (N_442,In_917,In_330);
and U443 (N_443,In_1335,In_1246);
or U444 (N_444,In_586,In_1724);
or U445 (N_445,In_111,In_710);
xnor U446 (N_446,In_669,In_1088);
xnor U447 (N_447,In_2000,In_2362);
and U448 (N_448,In_489,In_347);
xnor U449 (N_449,In_1768,In_1263);
nor U450 (N_450,In_1812,In_131);
xnor U451 (N_451,In_1583,In_262);
nor U452 (N_452,In_1130,In_592);
and U453 (N_453,In_1998,In_1416);
or U454 (N_454,In_1665,In_1744);
xor U455 (N_455,In_20,In_2046);
nand U456 (N_456,In_392,In_1229);
nand U457 (N_457,In_2438,In_1537);
nand U458 (N_458,In_1085,In_1097);
xor U459 (N_459,In_1054,In_644);
xor U460 (N_460,In_1286,In_1818);
nor U461 (N_461,In_451,In_1990);
or U462 (N_462,In_2268,In_1420);
nor U463 (N_463,In_395,In_995);
nand U464 (N_464,In_245,In_1113);
nand U465 (N_465,In_418,In_1493);
and U466 (N_466,In_2233,In_2413);
or U467 (N_467,In_1340,In_1863);
nand U468 (N_468,In_2019,In_2270);
or U469 (N_469,In_1049,In_1629);
nand U470 (N_470,In_840,In_190);
xnor U471 (N_471,In_912,In_121);
nor U472 (N_472,In_1522,In_2061);
and U473 (N_473,In_50,In_87);
nand U474 (N_474,In_236,In_1719);
nor U475 (N_475,In_2034,In_380);
nor U476 (N_476,In_1283,In_472);
nor U477 (N_477,In_2490,In_988);
xor U478 (N_478,In_2127,In_1510);
and U479 (N_479,In_1171,In_1337);
xnor U480 (N_480,In_478,In_2403);
nand U481 (N_481,In_985,In_114);
xnor U482 (N_482,In_2066,In_2360);
or U483 (N_483,In_709,In_885);
nor U484 (N_484,In_1390,In_1903);
nand U485 (N_485,In_676,In_343);
nand U486 (N_486,In_1072,In_2163);
nand U487 (N_487,In_808,In_1409);
and U488 (N_488,In_2370,In_1048);
nor U489 (N_489,In_299,In_961);
nand U490 (N_490,In_2306,In_77);
nand U491 (N_491,In_2366,In_38);
xnor U492 (N_492,In_763,In_2443);
and U493 (N_493,In_1727,In_2373);
and U494 (N_494,In_1428,In_875);
or U495 (N_495,In_1856,In_1544);
or U496 (N_496,In_1482,In_2401);
nor U497 (N_497,In_2452,In_1268);
xor U498 (N_498,In_909,In_2009);
xnor U499 (N_499,In_1091,In_2026);
and U500 (N_500,In_906,In_1329);
and U501 (N_501,In_747,In_1197);
and U502 (N_502,In_2301,In_755);
nor U503 (N_503,In_1841,In_2225);
or U504 (N_504,In_1857,In_1040);
and U505 (N_505,In_1486,In_1226);
xor U506 (N_506,In_2321,In_2091);
nand U507 (N_507,In_132,In_1580);
or U508 (N_508,In_400,In_1549);
or U509 (N_509,In_1679,In_153);
xor U510 (N_510,In_1353,In_2297);
xnor U511 (N_511,In_134,In_397);
and U512 (N_512,In_1604,In_1473);
and U513 (N_513,In_1074,In_526);
and U514 (N_514,In_2399,In_1080);
xnor U515 (N_515,In_84,In_2031);
and U516 (N_516,In_1322,In_690);
xor U517 (N_517,In_1291,In_1735);
nor U518 (N_518,In_2202,In_2421);
and U519 (N_519,In_200,In_1960);
nor U520 (N_520,In_1523,In_568);
or U521 (N_521,In_1710,In_443);
xor U522 (N_522,In_271,In_843);
nand U523 (N_523,In_2463,In_1809);
or U524 (N_524,In_946,In_1835);
xnor U525 (N_525,In_1443,In_688);
xor U526 (N_526,In_2393,In_2389);
xor U527 (N_527,In_541,In_164);
and U528 (N_528,In_1352,In_1913);
xor U529 (N_529,In_1659,In_768);
or U530 (N_530,In_1833,In_558);
nand U531 (N_531,In_860,In_272);
and U532 (N_532,In_1156,In_414);
nand U533 (N_533,In_2254,In_897);
xnor U534 (N_534,In_563,In_1060);
or U535 (N_535,In_401,In_1233);
or U536 (N_536,In_166,In_1098);
nor U537 (N_537,In_469,In_936);
nor U538 (N_538,In_456,In_2194);
nor U539 (N_539,In_1351,In_325);
and U540 (N_540,In_2340,In_1223);
nor U541 (N_541,In_368,In_1736);
xnor U542 (N_542,In_1415,In_959);
nand U543 (N_543,In_1407,In_34);
nor U544 (N_544,In_54,In_1081);
or U545 (N_545,In_331,In_2033);
nor U546 (N_546,In_2220,In_444);
nand U547 (N_547,In_623,In_871);
xnor U548 (N_548,In_103,In_1930);
or U549 (N_549,In_740,In_2035);
or U550 (N_550,In_1721,In_1989);
or U551 (N_551,In_431,In_1341);
and U552 (N_552,In_199,In_2457);
nand U553 (N_553,In_2173,In_2361);
or U554 (N_554,In_15,In_2420);
nor U555 (N_555,In_1800,In_1089);
and U556 (N_556,In_758,In_625);
and U557 (N_557,In_631,In_2465);
nor U558 (N_558,In_1061,In_475);
or U559 (N_559,In_2169,In_2470);
xor U560 (N_560,In_2024,In_2008);
nor U561 (N_561,In_1579,In_1786);
xnor U562 (N_562,In_313,In_326);
nor U563 (N_563,In_2455,In_802);
and U564 (N_564,In_1545,In_470);
xor U565 (N_565,In_1480,In_10);
nand U566 (N_566,In_711,In_1083);
nand U567 (N_567,In_48,In_1111);
xnor U568 (N_568,In_2259,In_1976);
nor U569 (N_569,In_447,In_250);
nor U570 (N_570,In_1776,In_1680);
or U571 (N_571,In_2245,In_2102);
and U572 (N_572,In_957,In_2378);
xor U573 (N_573,In_448,In_296);
xnor U574 (N_574,In_2460,In_2311);
nand U575 (N_575,In_2241,In_1799);
nand U576 (N_576,In_249,In_1546);
nand U577 (N_577,In_1271,In_1831);
or U578 (N_578,In_112,In_2054);
nor U579 (N_579,In_2143,In_881);
nor U580 (N_580,In_92,In_2155);
or U581 (N_581,In_1983,In_2065);
and U582 (N_582,In_1373,In_1021);
and U583 (N_583,In_852,In_1584);
nor U584 (N_584,In_1615,In_507);
nand U585 (N_585,In_394,In_1595);
nand U586 (N_586,In_518,In_863);
and U587 (N_587,In_1084,In_2229);
and U588 (N_588,In_2004,In_1871);
nor U589 (N_589,In_2315,In_1477);
or U590 (N_590,In_1947,In_1622);
nand U591 (N_591,In_311,In_2294);
nand U592 (N_592,In_1971,In_1949);
and U593 (N_593,In_2160,In_1343);
xor U594 (N_594,In_2322,In_1099);
or U595 (N_595,In_2180,In_1323);
and U596 (N_596,In_800,In_364);
xnor U597 (N_597,In_2461,In_913);
xor U598 (N_598,In_46,In_208);
nor U599 (N_599,In_2252,In_1907);
nor U600 (N_600,In_1297,In_350);
and U601 (N_601,In_1465,In_700);
nor U602 (N_602,In_901,In_2411);
nor U603 (N_603,In_1372,In_2349);
or U604 (N_604,In_68,In_104);
xor U605 (N_605,In_193,In_1848);
and U606 (N_606,In_1627,In_1319);
nor U607 (N_607,In_2025,In_1421);
nand U608 (N_608,In_1394,In_1616);
or U609 (N_609,In_555,In_1176);
xor U610 (N_610,In_963,In_2150);
or U611 (N_611,In_1296,In_1847);
nor U612 (N_612,In_2217,In_407);
and U613 (N_613,In_1993,In_609);
or U614 (N_614,In_1723,In_2146);
nand U615 (N_615,In_1117,In_1293);
nor U616 (N_616,In_1260,In_1982);
xnor U617 (N_617,In_1621,In_2481);
xor U618 (N_618,In_2200,In_1094);
nor U619 (N_619,In_2177,In_2282);
nor U620 (N_620,In_1137,In_178);
and U621 (N_621,In_1003,In_1596);
nor U622 (N_622,In_243,In_1518);
nand U623 (N_623,In_371,In_406);
nor U624 (N_624,In_2434,In_1281);
nand U625 (N_625,In_180,In_1128);
or U626 (N_626,In_405,In_1849);
xor U627 (N_627,In_928,In_1012);
and U628 (N_628,In_71,In_1418);
nor U629 (N_629,In_1957,In_1017);
xnor U630 (N_630,In_1361,In_2384);
or U631 (N_631,In_1977,In_1532);
nor U632 (N_632,In_2093,In_25);
nand U633 (N_633,In_479,In_1912);
nor U634 (N_634,In_2423,In_705);
xor U635 (N_635,In_593,In_1750);
nand U636 (N_636,In_78,In_1185);
and U637 (N_637,In_155,In_1412);
and U638 (N_638,In_2003,In_231);
or U639 (N_639,In_836,In_340);
xnor U640 (N_640,In_1959,In_1882);
or U641 (N_641,In_582,In_955);
nand U642 (N_642,In_1991,In_1570);
nand U643 (N_643,In_766,In_365);
nor U644 (N_644,In_2331,In_360);
or U645 (N_645,In_1144,In_771);
xnor U646 (N_646,In_1143,In_1453);
and U647 (N_647,In_937,In_2290);
and U648 (N_648,In_1507,In_2262);
nand U649 (N_649,In_979,In_2334);
and U650 (N_650,In_2355,In_2133);
or U651 (N_651,In_437,In_487);
nor U652 (N_652,In_2309,In_1861);
xor U653 (N_653,In_1694,In_1648);
nand U654 (N_654,In_1024,In_295);
nand U655 (N_655,In_1359,In_1321);
nand U656 (N_656,In_1876,In_1087);
or U657 (N_657,In_1711,In_702);
or U658 (N_658,In_234,In_761);
nor U659 (N_659,In_2105,In_973);
or U660 (N_660,In_1102,In_203);
and U661 (N_661,In_1481,In_2223);
and U662 (N_662,In_1859,In_2013);
nor U663 (N_663,In_1255,In_1603);
or U664 (N_664,In_1357,In_281);
and U665 (N_665,In_1422,In_1902);
nor U666 (N_666,In_398,In_1759);
or U667 (N_667,In_1382,In_1585);
and U668 (N_668,In_1663,In_217);
or U669 (N_669,In_1908,In_1600);
nand U670 (N_670,In_58,In_1423);
nor U671 (N_671,In_184,In_101);
nor U672 (N_672,In_2050,In_1814);
or U673 (N_673,In_1588,In_2449);
nor U674 (N_674,In_1267,In_1366);
and U675 (N_675,In_2128,In_2425);
nand U676 (N_676,In_673,In_2132);
xnor U677 (N_677,In_923,In_2304);
nor U678 (N_678,In_1783,In_96);
or U679 (N_679,In_2496,In_2450);
nand U680 (N_680,In_596,In_613);
nand U681 (N_681,In_1985,In_2279);
or U682 (N_682,In_2239,In_227);
and U683 (N_683,In_473,In_2319);
xnor U684 (N_684,In_1368,In_1231);
nor U685 (N_685,In_349,In_494);
and U686 (N_686,In_749,In_823);
or U687 (N_687,In_718,In_536);
and U688 (N_688,In_1879,In_2353);
nor U689 (N_689,In_2293,In_2092);
nand U690 (N_690,In_191,In_1300);
xor U691 (N_691,In_528,In_151);
and U692 (N_692,In_1301,In_72);
nor U693 (N_693,In_2433,In_876);
or U694 (N_694,In_459,In_607);
xnor U695 (N_695,In_175,In_404);
or U696 (N_696,In_856,In_2051);
xnor U697 (N_697,In_116,In_1988);
xor U698 (N_698,In_353,In_59);
and U699 (N_699,In_1313,In_2171);
xor U700 (N_700,In_980,In_1702);
xor U701 (N_701,In_122,In_2424);
xnor U702 (N_702,In_2338,In_864);
xnor U703 (N_703,In_952,In_693);
and U704 (N_704,In_496,In_504);
or U705 (N_705,In_647,In_2260);
or U706 (N_706,In_1865,In_1251);
and U707 (N_707,In_1250,In_2187);
xor U708 (N_708,In_446,In_861);
and U709 (N_709,In_698,In_1641);
and U710 (N_710,In_1307,In_888);
nor U711 (N_711,In_960,In_1179);
nor U712 (N_712,In_914,In_1184);
nor U713 (N_713,In_316,In_452);
or U714 (N_714,In_1501,In_1476);
nand U715 (N_715,In_1502,In_780);
and U716 (N_716,In_1161,In_1278);
nand U717 (N_717,In_1485,In_306);
nand U718 (N_718,In_2258,In_730);
xor U719 (N_719,In_975,In_2055);
nand U720 (N_720,In_1002,In_539);
and U721 (N_721,In_2106,In_1541);
nand U722 (N_722,In_1417,In_1771);
and U723 (N_723,In_348,In_2182);
nor U724 (N_724,In_682,In_2044);
or U725 (N_725,In_583,In_2451);
nor U726 (N_726,In_2208,In_230);
or U727 (N_727,In_376,In_989);
nand U728 (N_728,In_1059,In_1204);
nor U729 (N_729,In_554,In_804);
xnor U730 (N_730,In_2276,In_1652);
or U731 (N_731,In_503,In_264);
nor U732 (N_732,In_1643,In_915);
or U733 (N_733,In_779,In_233);
nand U734 (N_734,In_1760,In_1076);
and U735 (N_735,In_2152,In_2161);
and U736 (N_736,In_2418,In_724);
nor U737 (N_737,In_1927,In_95);
and U738 (N_738,In_2120,In_2211);
or U739 (N_739,In_1645,In_606);
xor U740 (N_740,In_102,In_646);
and U741 (N_741,In_660,In_342);
xnor U742 (N_742,In_1692,In_659);
nand U743 (N_743,In_1592,In_1444);
and U744 (N_744,In_1016,In_1779);
nor U745 (N_745,In_2277,In_819);
or U746 (N_746,In_109,In_2174);
and U747 (N_747,In_1441,In_573);
nand U748 (N_748,In_2454,In_2298);
nor U749 (N_749,In_130,In_1832);
and U750 (N_750,In_1033,In_926);
nor U751 (N_751,In_40,In_982);
nand U752 (N_752,In_575,In_1915);
or U753 (N_753,In_1968,In_334);
or U754 (N_754,In_1019,In_944);
and U755 (N_755,In_1364,In_842);
nand U756 (N_756,In_1560,In_107);
xnor U757 (N_757,In_335,In_630);
xor U758 (N_758,In_2042,In_745);
nor U759 (N_759,In_1009,In_954);
nor U760 (N_760,In_1886,In_934);
or U761 (N_761,In_640,In_1287);
nor U762 (N_762,In_426,In_958);
and U763 (N_763,In_2080,In_1793);
or U764 (N_764,In_714,In_1852);
xnor U765 (N_765,In_1302,In_1747);
xor U766 (N_766,In_1950,In_2283);
nand U767 (N_767,In_1808,In_493);
and U768 (N_768,In_1858,In_1459);
or U769 (N_769,In_37,In_830);
nand U770 (N_770,In_1410,In_378);
nor U771 (N_771,In_501,In_548);
and U772 (N_772,In_1707,In_628);
xor U773 (N_773,In_1931,In_731);
nand U774 (N_774,In_722,In_1836);
or U775 (N_775,In_1358,In_2167);
nand U776 (N_776,In_2348,In_2336);
nand U777 (N_777,In_1715,In_1064);
or U778 (N_778,In_854,In_366);
or U779 (N_779,In_454,In_715);
nor U780 (N_780,In_324,In_2383);
nor U781 (N_781,In_1070,In_2352);
nand U782 (N_782,In_1354,In_1550);
nand U783 (N_783,In_1571,In_44);
xor U784 (N_784,In_2477,In_1200);
or U785 (N_785,In_1279,In_1461);
nor U786 (N_786,In_1521,In_1654);
nand U787 (N_787,In_1671,In_382);
nor U788 (N_788,In_2390,In_678);
xnor U789 (N_789,In_287,In_2478);
or U790 (N_790,In_1817,In_1937);
nand U791 (N_791,In_1038,In_629);
xnor U792 (N_792,In_1773,In_1827);
and U793 (N_793,In_2017,In_254);
xnor U794 (N_794,In_2402,In_385);
xnor U795 (N_795,In_1966,In_2006);
or U796 (N_796,In_1766,In_2084);
and U797 (N_797,In_2281,In_2346);
xnor U798 (N_798,In_632,In_1146);
nor U799 (N_799,In_182,In_807);
and U800 (N_800,In_399,In_1450);
and U801 (N_801,In_28,In_1312);
nand U802 (N_802,In_746,In_1311);
and U803 (N_803,In_31,In_1614);
nand U804 (N_804,In_2020,In_1548);
nor U805 (N_805,In_1440,In_1687);
xor U806 (N_806,In_699,In_916);
or U807 (N_807,In_2445,In_2391);
nand U808 (N_808,In_2337,In_791);
xnor U809 (N_809,In_703,In_1881);
xor U810 (N_810,In_1436,In_1763);
and U811 (N_811,In_1062,In_621);
xor U812 (N_812,In_1261,In_338);
xor U813 (N_813,In_307,In_1824);
or U814 (N_814,In_983,In_171);
and U815 (N_815,In_1170,In_1437);
or U816 (N_816,In_42,In_329);
nor U817 (N_817,In_106,In_308);
nor U818 (N_818,In_500,In_1672);
xor U819 (N_819,In_1823,In_677);
nand U820 (N_820,In_2466,In_734);
nor U821 (N_821,In_1258,In_1151);
nand U822 (N_822,In_1023,In_626);
or U823 (N_823,In_1846,In_502);
nor U824 (N_824,In_1494,In_787);
nand U825 (N_825,In_790,In_661);
nor U826 (N_826,In_2124,In_825);
xor U827 (N_827,In_2377,In_1790);
nor U828 (N_828,In_2153,In_1675);
nand U829 (N_829,In_1559,In_2284);
nand U830 (N_830,In_859,In_117);
nor U831 (N_831,In_1334,In_1752);
xnor U832 (N_832,In_1626,In_1787);
nor U833 (N_833,In_953,In_471);
nor U834 (N_834,In_608,In_332);
and U835 (N_835,In_1055,In_1001);
or U836 (N_836,In_2350,In_1558);
xnor U837 (N_837,In_189,In_2316);
nand U838 (N_838,In_2379,In_52);
nand U839 (N_839,In_129,In_1536);
and U840 (N_840,In_1239,In_2113);
nor U841 (N_841,In_356,In_2145);
nor U842 (N_842,In_1512,In_141);
nor U843 (N_843,In_1304,In_978);
or U844 (N_844,In_2045,In_1573);
or U845 (N_845,In_806,In_1330);
nand U846 (N_846,In_1613,In_2299);
nand U847 (N_847,In_950,In_2329);
or U848 (N_848,In_1401,In_1958);
nor U849 (N_849,In_908,In_318);
nor U850 (N_850,In_1682,In_1082);
xor U851 (N_851,In_1973,In_1316);
and U852 (N_852,In_643,In_1919);
xnor U853 (N_853,In_1162,In_540);
xor U854 (N_854,In_707,In_268);
xor U855 (N_855,In_1264,In_760);
nand U856 (N_856,In_127,In_651);
nand U857 (N_857,In_445,In_1210);
nand U858 (N_858,In_2380,In_1756);
or U859 (N_859,In_545,In_633);
xnor U860 (N_860,In_2216,In_1027);
and U861 (N_861,In_1280,In_89);
nand U862 (N_862,In_1479,In_291);
nand U863 (N_863,In_560,In_160);
and U864 (N_864,In_708,In_862);
nand U865 (N_865,In_1753,In_2429);
nor U866 (N_866,In_2049,In_2222);
or U867 (N_867,In_211,In_2328);
and U868 (N_868,In_1869,In_680);
or U869 (N_869,In_645,In_1530);
nand U870 (N_870,In_728,In_2015);
or U871 (N_871,In_1767,In_269);
nor U872 (N_872,In_372,In_1954);
nand U873 (N_873,In_770,In_1132);
or U874 (N_874,In_619,In_179);
xnor U875 (N_875,In_235,In_2385);
and U876 (N_876,In_1051,In_1158);
nand U877 (N_877,In_174,In_137);
or U878 (N_878,In_1635,In_2014);
nor U879 (N_879,In_2364,In_1568);
or U880 (N_880,In_2308,In_2479);
nand U881 (N_881,In_1205,In_1874);
or U882 (N_882,In_158,In_2375);
nor U883 (N_883,In_2086,In_1391);
xor U884 (N_884,In_1986,In_1256);
and U885 (N_885,In_2300,In_832);
or U886 (N_886,In_981,In_1234);
nand U887 (N_887,In_664,In_2154);
nand U888 (N_888,In_616,In_2292);
or U889 (N_889,In_1225,In_1875);
nor U890 (N_890,In_1426,In_1090);
nand U891 (N_891,In_1602,In_577);
xnor U892 (N_892,In_1574,In_588);
and U893 (N_893,In_2059,In_1734);
xnor U894 (N_894,In_614,In_1695);
nand U895 (N_895,In_2253,In_1543);
or U896 (N_896,In_1924,In_666);
nand U897 (N_897,In_2041,In_1215);
or U898 (N_898,In_18,In_1126);
nand U899 (N_899,In_2109,In_2396);
xnor U900 (N_900,In_1576,In_1676);
xor U901 (N_901,In_1508,In_535);
and U902 (N_902,In_1524,In_904);
and U903 (N_903,In_1918,In_1826);
nor U904 (N_904,In_1434,In_461);
and U905 (N_905,In_150,In_1497);
or U906 (N_906,In_566,In_889);
xnor U907 (N_907,In_303,In_1451);
xnor U908 (N_908,In_321,In_2459);
or U909 (N_909,In_2095,In_638);
and U910 (N_910,In_525,In_751);
nand U911 (N_911,In_1925,In_1788);
xor U912 (N_912,In_374,In_434);
nand U913 (N_913,In_1555,In_1764);
or U914 (N_914,In_2274,In_1116);
or U915 (N_915,In_2104,In_814);
xnor U916 (N_916,In_1936,In_2320);
and U917 (N_917,In_2166,In_725);
nand U918 (N_918,In_792,In_2069);
nor U919 (N_919,In_2394,In_720);
nand U920 (N_920,In_283,In_2157);
xnor U921 (N_921,In_253,In_1638);
or U922 (N_922,In_1484,In_1625);
xor U923 (N_923,In_1029,In_2083);
nor U924 (N_924,In_1022,In_373);
nor U925 (N_925,In_642,In_168);
or U926 (N_926,In_88,In_597);
and U927 (N_927,In_1044,In_1266);
nand U928 (N_928,In_1529,In_942);
nor U929 (N_929,In_1288,In_1471);
nor U930 (N_930,In_2125,In_634);
nand U931 (N_931,In_32,In_225);
or U932 (N_932,In_1041,In_2467);
and U933 (N_933,In_1506,In_774);
xnor U934 (N_934,In_53,In_510);
nor U935 (N_935,In_1273,In_145);
and U936 (N_936,In_27,In_480);
nor U937 (N_937,In_794,In_1700);
nand U938 (N_938,In_1174,In_550);
nor U939 (N_939,In_1701,In_247);
nor U940 (N_940,In_741,In_820);
nor U941 (N_941,In_255,In_918);
and U942 (N_942,In_419,In_737);
or U943 (N_943,In_1932,In_1693);
nor U944 (N_944,In_1582,In_1843);
or U945 (N_945,In_2141,In_1107);
xor U946 (N_946,In_1853,In_2310);
nand U947 (N_947,In_428,In_2303);
or U948 (N_948,In_2121,In_529);
and U949 (N_949,In_1466,In_1245);
nand U950 (N_950,In_1167,In_354);
nand U951 (N_951,In_675,In_1742);
and U952 (N_952,In_2416,In_1851);
xnor U953 (N_953,In_1586,In_1121);
and U954 (N_954,In_1134,In_2135);
nor U955 (N_955,In_425,In_126);
nor U956 (N_956,In_998,In_726);
xnor U957 (N_957,In_1746,In_999);
or U958 (N_958,In_945,In_1013);
nor U959 (N_959,In_1598,In_2071);
nor U960 (N_960,In_1722,In_1975);
or U961 (N_961,In_639,In_2089);
and U962 (N_962,In_2499,In_1914);
or U963 (N_963,In_2240,In_2199);
and U964 (N_964,In_429,In_2475);
or U965 (N_965,In_492,In_196);
or U966 (N_966,In_1227,In_2280);
or U967 (N_967,In_968,In_2440);
xnor U968 (N_968,In_1031,In_1873);
xnor U969 (N_969,In_1446,In_2417);
xnor U970 (N_970,In_2382,In_1961);
xor U971 (N_971,In_490,In_2053);
nor U972 (N_972,In_1190,In_2448);
or U973 (N_973,In_2068,In_1043);
or U974 (N_974,In_2265,In_637);
and U975 (N_975,In_511,In_1345);
and U976 (N_976,In_119,In_789);
and U977 (N_977,In_2052,In_279);
or U978 (N_978,In_1740,In_1505);
or U979 (N_979,In_26,In_1454);
or U980 (N_980,In_2255,In_435);
or U981 (N_981,In_1926,In_2342);
nand U982 (N_982,In_1383,In_123);
and U983 (N_983,In_1498,In_544);
or U984 (N_984,In_2286,In_2184);
and U985 (N_985,In_801,In_2201);
or U986 (N_986,In_697,In_69);
or U987 (N_987,In_2432,In_585);
nor U988 (N_988,In_1556,In_1047);
nor U989 (N_989,In_1333,In_2323);
and U990 (N_990,In_2048,In_1212);
nand U991 (N_991,In_176,In_1004);
or U992 (N_992,In_1825,In_1073);
and U993 (N_993,In_821,In_1965);
nand U994 (N_994,In_1240,In_2472);
and U995 (N_995,In_357,In_79);
or U996 (N_996,In_298,In_2085);
nor U997 (N_997,In_932,In_788);
or U998 (N_998,In_94,In_232);
nor U999 (N_999,In_427,In_120);
xor U1000 (N_1000,In_1489,In_1733);
and U1001 (N_1001,In_2430,In_2016);
and U1002 (N_1002,In_1377,In_1092);
and U1003 (N_1003,In_865,In_1713);
nand U1004 (N_1004,In_506,In_421);
or U1005 (N_1005,In_274,In_1036);
xor U1006 (N_1006,In_838,In_736);
or U1007 (N_1007,In_551,In_1380);
nor U1008 (N_1008,In_1725,In_1525);
nor U1009 (N_1009,In_2244,In_1173);
nand U1010 (N_1010,In_706,In_1235);
and U1011 (N_1011,In_579,In_996);
and U1012 (N_1012,In_2151,In_410);
and U1013 (N_1013,In_1554,In_466);
xnor U1014 (N_1014,In_1375,In_2140);
nand U1015 (N_1015,In_590,In_1870);
or U1016 (N_1016,In_1299,In_2251);
nand U1017 (N_1017,In_2235,In_1365);
nand U1018 (N_1018,In_39,In_1165);
nand U1019 (N_1019,In_29,In_2238);
xor U1020 (N_1020,In_1349,In_436);
and U1021 (N_1021,In_2007,In_2428);
or U1022 (N_1022,In_2193,In_1405);
xnor U1023 (N_1023,In_1138,In_169);
xnor U1024 (N_1024,In_874,In_1587);
xor U1025 (N_1025,In_1193,In_1842);
nor U1026 (N_1026,In_993,In_2090);
and U1027 (N_1027,In_1569,In_1738);
and U1028 (N_1028,In_1741,In_1456);
or U1029 (N_1029,In_1709,In_1039);
nor U1030 (N_1030,In_1955,In_1015);
or U1031 (N_1031,In_468,In_658);
and U1032 (N_1032,In_265,In_2357);
xnor U1033 (N_1033,In_2162,In_2312);
xnor U1034 (N_1034,In_1634,In_2158);
nor U1035 (N_1035,In_1303,In_831);
or U1036 (N_1036,In_922,In_138);
xnor U1037 (N_1037,In_1014,In_147);
or U1038 (N_1038,In_2462,In_1705);
nor U1039 (N_1039,In_1392,In_173);
and U1040 (N_1040,In_622,In_2324);
nand U1041 (N_1041,In_1077,In_1678);
or U1042 (N_1042,In_93,In_441);
nor U1043 (N_1043,In_1605,In_1195);
nand U1044 (N_1044,In_463,In_2185);
nor U1045 (N_1045,In_1242,In_1320);
nand U1046 (N_1046,In_474,In_1714);
or U1047 (N_1047,In_1921,In_1491);
and U1048 (N_1048,In_1474,In_1934);
xor U1049 (N_1049,In_841,In_668);
or U1050 (N_1050,In_464,In_2376);
xnor U1051 (N_1051,In_1612,In_1552);
nand U1052 (N_1052,In_1289,In_2165);
or U1053 (N_1053,In_938,In_2447);
and U1054 (N_1054,In_1795,In_1894);
nand U1055 (N_1055,In_222,In_1114);
xor U1056 (N_1056,In_1942,In_57);
xnor U1057 (N_1057,In_1100,In_377);
nand U1058 (N_1058,In_282,In_743);
xor U1059 (N_1059,In_931,In_1610);
nor U1060 (N_1060,In_1414,In_1);
xnor U1061 (N_1061,In_900,In_750);
xor U1062 (N_1062,In_1980,In_951);
xnor U1063 (N_1063,In_712,In_1775);
or U1064 (N_1064,In_1008,In_2123);
or U1065 (N_1065,In_2176,In_2098);
nor U1066 (N_1066,In_1309,In_611);
xor U1067 (N_1067,In_83,In_1148);
nor U1068 (N_1068,In_1292,In_2247);
or U1069 (N_1069,In_1737,In_1891);
or U1070 (N_1070,In_1495,In_1331);
xnor U1071 (N_1071,In_465,In_2204);
nand U1072 (N_1072,In_1945,In_1963);
xor U1073 (N_1073,In_2179,In_2456);
or U1074 (N_1074,In_1837,In_2256);
nor U1075 (N_1075,In_1037,In_403);
and U1076 (N_1076,In_663,In_2248);
or U1077 (N_1077,In_574,In_783);
nor U1078 (N_1078,In_1006,In_159);
nor U1079 (N_1079,In_1593,In_1642);
nand U1080 (N_1080,In_695,In_276);
and U1081 (N_1081,In_2147,In_618);
or U1082 (N_1082,In_1577,In_1667);
or U1083 (N_1083,In_572,In_933);
nor U1084 (N_1084,In_1732,In_910);
xnor U1085 (N_1085,In_1748,In_1065);
or U1086 (N_1086,In_1243,In_1211);
and U1087 (N_1087,In_1822,In_1572);
or U1088 (N_1088,In_75,In_1619);
nand U1089 (N_1089,In_1105,In_1439);
and U1090 (N_1090,In_1594,In_687);
xnor U1091 (N_1091,In_1406,In_2264);
or U1092 (N_1092,In_866,In_1564);
xnor U1093 (N_1093,In_251,In_2212);
or U1094 (N_1094,In_1472,In_1792);
and U1095 (N_1095,In_1177,In_482);
nand U1096 (N_1096,In_1897,In_2076);
xnor U1097 (N_1097,In_14,In_2063);
nor U1098 (N_1098,In_1772,In_793);
nand U1099 (N_1099,In_312,In_1686);
and U1100 (N_1100,In_1499,In_244);
and U1101 (N_1101,In_124,In_1829);
xnor U1102 (N_1102,In_1386,In_1327);
or U1103 (N_1103,In_1784,In_370);
or U1104 (N_1104,In_1135,In_2077);
nand U1105 (N_1105,In_512,In_1511);
nor U1106 (N_1106,In_1488,In_1068);
xnor U1107 (N_1107,In_1462,In_346);
and U1108 (N_1108,In_1153,In_333);
or U1109 (N_1109,In_275,In_2002);
nand U1110 (N_1110,In_1547,In_2325);
or U1111 (N_1111,In_811,In_1967);
nor U1112 (N_1112,In_552,In_142);
xnor U1113 (N_1113,In_1408,In_226);
nor U1114 (N_1114,In_1575,In_1906);
and U1115 (N_1115,In_1561,In_603);
nor U1116 (N_1116,In_1885,In_753);
nand U1117 (N_1117,In_1413,In_850);
xor U1118 (N_1118,In_1429,In_795);
xor U1119 (N_1119,In_1052,In_259);
nand U1120 (N_1120,In_1845,In_2395);
or U1121 (N_1121,In_1254,In_1910);
nand U1122 (N_1122,In_570,In_1674);
or U1123 (N_1123,In_361,In_1997);
nor U1124 (N_1124,In_2129,In_352);
or U1125 (N_1125,In_449,In_1984);
xor U1126 (N_1126,In_497,In_98);
nor U1127 (N_1127,In_1899,In_1534);
or U1128 (N_1128,In_1951,In_2468);
xnor U1129 (N_1129,In_822,In_248);
nor U1130 (N_1130,In_246,In_1457);
xor U1131 (N_1131,In_432,In_43);
nand U1132 (N_1132,In_2344,In_433);
nand U1133 (N_1133,In_2407,In_2406);
nand U1134 (N_1134,In_2446,In_1387);
xnor U1135 (N_1135,In_1660,In_2188);
xnor U1136 (N_1136,In_1367,In_1157);
nand U1137 (N_1137,In_396,In_1145);
and U1138 (N_1138,In_337,In_2196);
and U1139 (N_1139,In_241,In_125);
nand U1140 (N_1140,In_2305,In_713);
xnor U1141 (N_1141,In_460,In_853);
nand U1142 (N_1142,In_984,In_1220);
nor U1143 (N_1143,In_1673,In_1447);
or U1144 (N_1144,In_207,In_2368);
nand U1145 (N_1145,In_1178,In_1703);
xnor U1146 (N_1146,In_891,In_17);
nor U1147 (N_1147,In_567,In_1483);
or U1148 (N_1148,In_476,In_1514);
nor U1149 (N_1149,In_358,In_1797);
or U1150 (N_1150,In_2030,In_2191);
nor U1151 (N_1151,In_1789,In_1830);
or U1152 (N_1152,In_1449,In_1698);
or U1153 (N_1153,In_411,In_185);
nand U1154 (N_1154,In_870,In_1578);
xor U1155 (N_1155,In_74,In_1403);
and U1156 (N_1156,In_2203,In_2330);
xor U1157 (N_1157,In_649,In_636);
xnor U1158 (N_1158,In_2082,In_1689);
nor U1159 (N_1159,In_2079,In_2414);
or U1160 (N_1160,In_240,In_781);
and U1161 (N_1161,In_1785,In_1551);
nand U1162 (N_1162,In_1527,In_624);
nor U1163 (N_1163,In_1677,In_238);
or U1164 (N_1164,In_1147,In_485);
or U1165 (N_1165,In_2039,In_35);
or U1166 (N_1166,In_1888,In_1834);
and U1167 (N_1167,In_966,In_1182);
nand U1168 (N_1168,In_458,In_1974);
or U1169 (N_1169,In_941,In_1187);
and U1170 (N_1170,In_1348,In_1272);
xor U1171 (N_1171,In_2474,In_785);
nor U1172 (N_1172,In_284,In_202);
nor U1173 (N_1173,In_847,In_1867);
xor U1174 (N_1174,In_911,In_488);
nand U1175 (N_1175,In_1890,In_2136);
and U1176 (N_1176,In_2345,In_2012);
xor U1177 (N_1177,In_2011,In_76);
xor U1178 (N_1178,In_51,In_45);
and U1179 (N_1179,In_67,In_1696);
or U1180 (N_1180,In_2056,In_105);
or U1181 (N_1181,In_1953,In_1275);
nor U1182 (N_1182,In_1011,In_1154);
xnor U1183 (N_1183,In_450,In_887);
and U1184 (N_1184,In_1905,In_2372);
xnor U1185 (N_1185,In_976,In_1651);
or U1186 (N_1186,In_884,In_300);
xor U1187 (N_1187,In_149,In_3);
and U1188 (N_1188,In_776,In_2435);
and U1189 (N_1189,In_1729,In_2175);
nand U1190 (N_1190,In_1344,In_2227);
or U1191 (N_1191,In_1889,In_598);
and U1192 (N_1192,In_304,In_1045);
or U1193 (N_1193,In_1046,In_1265);
and U1194 (N_1194,In_108,In_1893);
nand U1195 (N_1195,In_1798,In_1743);
nor U1196 (N_1196,In_110,In_2387);
xor U1197 (N_1197,In_1460,In_317);
or U1198 (N_1198,In_2170,In_869);
and U1199 (N_1199,In_315,In_1346);
or U1200 (N_1200,In_1124,In_239);
nand U1201 (N_1201,In_1770,In_1774);
nand U1202 (N_1202,In_1355,In_285);
nand U1203 (N_1203,In_692,In_1513);
nor U1204 (N_1204,In_2307,In_1956);
nand U1205 (N_1205,In_686,In_442);
nand U1206 (N_1206,In_379,In_1519);
and U1207 (N_1207,In_1828,In_204);
nand U1208 (N_1208,In_1691,In_964);
xnor U1209 (N_1209,In_1657,In_412);
nand U1210 (N_1210,In_2209,In_2215);
xnor U1211 (N_1211,In_672,In_834);
xor U1212 (N_1212,In_2263,In_1181);
and U1213 (N_1213,In_41,In_1815);
nor U1214 (N_1214,In_1115,In_2210);
nor U1215 (N_1215,In_2096,In_797);
nand U1216 (N_1216,In_1433,In_2291);
nor U1217 (N_1217,In_221,In_1224);
xor U1218 (N_1218,In_537,In_115);
nand U1219 (N_1219,In_1402,In_21);
and U1220 (N_1220,In_8,In_949);
nor U1221 (N_1221,In_1630,In_1469);
or U1222 (N_1222,In_2326,In_1820);
or U1223 (N_1223,In_1119,In_1699);
nand U1224 (N_1224,In_930,In_1928);
or U1225 (N_1225,In_530,In_1948);
and U1226 (N_1226,In_739,In_1244);
or U1227 (N_1227,In_383,In_305);
nor U1228 (N_1228,In_580,In_899);
nand U1229 (N_1229,In_694,In_2137);
nand U1230 (N_1230,In_1731,In_462);
and U1231 (N_1231,In_587,In_498);
and U1232 (N_1232,In_12,In_1813);
nor U1233 (N_1233,In_375,In_892);
xor U1234 (N_1234,In_2471,In_719);
xnor U1235 (N_1235,In_571,In_754);
nand U1236 (N_1236,In_1801,In_2029);
nor U1237 (N_1237,In_1305,In_1237);
xor U1238 (N_1238,In_627,In_1332);
xor U1239 (N_1239,In_2267,In_1149);
xnor U1240 (N_1240,In_402,In_1683);
xnor U1241 (N_1241,In_1646,In_1095);
nand U1242 (N_1242,In_2230,In_1201);
nor U1243 (N_1243,In_1607,In_1590);
xor U1244 (N_1244,In_167,In_1325);
or U1245 (N_1245,In_223,In_2);
nor U1246 (N_1246,In_1306,In_9);
nor U1247 (N_1247,In_696,In_2486);
or U1248 (N_1248,In_1780,In_1208);
or U1249 (N_1249,In_369,In_1350);
and U1250 (N_1250,N_599,N_1078);
or U1251 (N_1251,N_372,N_15);
nand U1252 (N_1252,N_148,N_511);
nand U1253 (N_1253,N_262,N_170);
and U1254 (N_1254,N_42,N_211);
and U1255 (N_1255,N_753,N_1249);
and U1256 (N_1256,N_353,N_225);
and U1257 (N_1257,N_1127,N_594);
nor U1258 (N_1258,N_1081,N_556);
xor U1259 (N_1259,N_366,N_915);
nor U1260 (N_1260,N_662,N_842);
and U1261 (N_1261,N_525,N_1180);
nor U1262 (N_1262,N_215,N_1118);
nor U1263 (N_1263,N_34,N_947);
or U1264 (N_1264,N_365,N_963);
xor U1265 (N_1265,N_1073,N_780);
nor U1266 (N_1266,N_120,N_544);
or U1267 (N_1267,N_1087,N_758);
xor U1268 (N_1268,N_582,N_125);
nand U1269 (N_1269,N_958,N_1097);
nand U1270 (N_1270,N_340,N_1157);
nand U1271 (N_1271,N_218,N_520);
or U1272 (N_1272,N_943,N_906);
nand U1273 (N_1273,N_115,N_269);
and U1274 (N_1274,N_699,N_551);
nand U1275 (N_1275,N_1062,N_709);
or U1276 (N_1276,N_213,N_343);
or U1277 (N_1277,N_281,N_234);
nand U1278 (N_1278,N_100,N_476);
and U1279 (N_1279,N_109,N_253);
and U1280 (N_1280,N_394,N_1048);
and U1281 (N_1281,N_1202,N_837);
and U1282 (N_1282,N_941,N_506);
xnor U1283 (N_1283,N_223,N_85);
or U1284 (N_1284,N_152,N_67);
nor U1285 (N_1285,N_590,N_212);
and U1286 (N_1286,N_1027,N_362);
nand U1287 (N_1287,N_329,N_414);
nor U1288 (N_1288,N_332,N_279);
nand U1289 (N_1289,N_694,N_220);
nor U1290 (N_1290,N_157,N_700);
and U1291 (N_1291,N_685,N_79);
nand U1292 (N_1292,N_78,N_824);
xnor U1293 (N_1293,N_1142,N_130);
and U1294 (N_1294,N_265,N_178);
nand U1295 (N_1295,N_760,N_964);
nor U1296 (N_1296,N_49,N_1043);
nand U1297 (N_1297,N_274,N_386);
nand U1298 (N_1298,N_885,N_647);
xnor U1299 (N_1299,N_196,N_495);
nand U1300 (N_1300,N_1176,N_299);
and U1301 (N_1301,N_89,N_1195);
and U1302 (N_1302,N_859,N_376);
nand U1303 (N_1303,N_977,N_75);
nor U1304 (N_1304,N_450,N_287);
nor U1305 (N_1305,N_1045,N_987);
or U1306 (N_1306,N_992,N_490);
xnor U1307 (N_1307,N_789,N_494);
and U1308 (N_1308,N_369,N_1101);
nand U1309 (N_1309,N_676,N_384);
nor U1310 (N_1310,N_289,N_429);
xor U1311 (N_1311,N_275,N_895);
nand U1312 (N_1312,N_921,N_466);
nor U1313 (N_1313,N_349,N_45);
nor U1314 (N_1314,N_166,N_568);
or U1315 (N_1315,N_725,N_1034);
nor U1316 (N_1316,N_1134,N_887);
nor U1317 (N_1317,N_993,N_229);
xor U1318 (N_1318,N_953,N_385);
or U1319 (N_1319,N_534,N_33);
nor U1320 (N_1320,N_827,N_938);
xnor U1321 (N_1321,N_905,N_1152);
nor U1322 (N_1322,N_1058,N_889);
xnor U1323 (N_1323,N_339,N_187);
or U1324 (N_1324,N_620,N_810);
xnor U1325 (N_1325,N_893,N_409);
nand U1326 (N_1326,N_614,N_1124);
nand U1327 (N_1327,N_31,N_256);
nor U1328 (N_1328,N_184,N_712);
nor U1329 (N_1329,N_756,N_465);
nor U1330 (N_1330,N_421,N_1015);
or U1331 (N_1331,N_65,N_59);
nand U1332 (N_1332,N_999,N_801);
xnor U1333 (N_1333,N_675,N_722);
nor U1334 (N_1334,N_843,N_1190);
nor U1335 (N_1335,N_474,N_542);
and U1336 (N_1336,N_829,N_788);
xor U1337 (N_1337,N_762,N_392);
or U1338 (N_1338,N_496,N_442);
or U1339 (N_1339,N_733,N_617);
xnor U1340 (N_1340,N_127,N_577);
nor U1341 (N_1341,N_441,N_896);
and U1342 (N_1342,N_576,N_432);
nand U1343 (N_1343,N_249,N_569);
nor U1344 (N_1344,N_192,N_633);
nand U1345 (N_1345,N_347,N_565);
nor U1346 (N_1346,N_686,N_161);
xnor U1347 (N_1347,N_379,N_295);
nand U1348 (N_1348,N_47,N_62);
xnor U1349 (N_1349,N_1242,N_1244);
or U1350 (N_1350,N_149,N_139);
and U1351 (N_1351,N_361,N_69);
nor U1352 (N_1352,N_5,N_389);
nand U1353 (N_1353,N_397,N_759);
or U1354 (N_1354,N_588,N_1094);
xnor U1355 (N_1355,N_322,N_367);
or U1356 (N_1356,N_848,N_1010);
xnor U1357 (N_1357,N_1013,N_683);
nor U1358 (N_1358,N_418,N_1002);
nand U1359 (N_1359,N_479,N_557);
nor U1360 (N_1360,N_68,N_26);
nor U1361 (N_1361,N_899,N_567);
nor U1362 (N_1362,N_790,N_1133);
xor U1363 (N_1363,N_1248,N_373);
and U1364 (N_1364,N_919,N_995);
and U1365 (N_1365,N_74,N_784);
nor U1366 (N_1366,N_294,N_636);
and U1367 (N_1367,N_1056,N_165);
nor U1368 (N_1368,N_527,N_955);
nor U1369 (N_1369,N_1079,N_444);
and U1370 (N_1370,N_950,N_1074);
nand U1371 (N_1371,N_734,N_183);
xor U1372 (N_1372,N_711,N_1247);
or U1373 (N_1373,N_804,N_140);
xnor U1374 (N_1374,N_334,N_333);
nand U1375 (N_1375,N_198,N_350);
xnor U1376 (N_1376,N_110,N_822);
nor U1377 (N_1377,N_1214,N_1135);
nor U1378 (N_1378,N_598,N_847);
and U1379 (N_1379,N_293,N_570);
or U1380 (N_1380,N_737,N_1088);
or U1381 (N_1381,N_671,N_1077);
and U1382 (N_1382,N_888,N_924);
and U1383 (N_1383,N_431,N_1187);
and U1384 (N_1384,N_66,N_448);
xor U1385 (N_1385,N_1139,N_719);
or U1386 (N_1386,N_849,N_50);
xor U1387 (N_1387,N_961,N_169);
or U1388 (N_1388,N_546,N_302);
nand U1389 (N_1389,N_913,N_1229);
and U1390 (N_1390,N_1111,N_603);
xnor U1391 (N_1391,N_357,N_635);
and U1392 (N_1392,N_739,N_1119);
nor U1393 (N_1393,N_687,N_358);
and U1394 (N_1394,N_607,N_245);
or U1395 (N_1395,N_724,N_1050);
or U1396 (N_1396,N_285,N_1130);
nor U1397 (N_1397,N_862,N_1046);
xor U1398 (N_1398,N_589,N_420);
nor U1399 (N_1399,N_816,N_716);
nor U1400 (N_1400,N_738,N_718);
nor U1401 (N_1401,N_501,N_503);
and U1402 (N_1402,N_167,N_584);
xnor U1403 (N_1403,N_639,N_1047);
nand U1404 (N_1404,N_328,N_1159);
or U1405 (N_1405,N_1035,N_36);
or U1406 (N_1406,N_1167,N_710);
nand U1407 (N_1407,N_946,N_752);
nand U1408 (N_1408,N_1109,N_640);
nor U1409 (N_1409,N_1039,N_1216);
xnor U1410 (N_1410,N_1126,N_288);
and U1411 (N_1411,N_510,N_27);
and U1412 (N_1412,N_775,N_684);
nor U1413 (N_1413,N_473,N_858);
nand U1414 (N_1414,N_619,N_174);
or U1415 (N_1415,N_459,N_748);
or U1416 (N_1416,N_1061,N_255);
xnor U1417 (N_1417,N_297,N_702);
nand U1418 (N_1418,N_940,N_1240);
or U1419 (N_1419,N_925,N_1189);
nor U1420 (N_1420,N_292,N_307);
xor U1421 (N_1421,N_948,N_338);
and U1422 (N_1422,N_492,N_560);
nor U1423 (N_1423,N_536,N_855);
or U1424 (N_1424,N_935,N_203);
or U1425 (N_1425,N_882,N_949);
nand U1426 (N_1426,N_8,N_934);
xnor U1427 (N_1427,N_871,N_43);
xor U1428 (N_1428,N_704,N_116);
and U1429 (N_1429,N_715,N_439);
and U1430 (N_1430,N_830,N_615);
xor U1431 (N_1431,N_706,N_735);
xor U1432 (N_1432,N_540,N_886);
nor U1433 (N_1433,N_98,N_217);
nand U1434 (N_1434,N_809,N_1096);
and U1435 (N_1435,N_644,N_356);
and U1436 (N_1436,N_757,N_375);
nor U1437 (N_1437,N_1173,N_346);
nand U1438 (N_1438,N_82,N_656);
nand U1439 (N_1439,N_927,N_868);
and U1440 (N_1440,N_866,N_173);
and U1441 (N_1441,N_547,N_657);
nand U1442 (N_1442,N_162,N_348);
or U1443 (N_1443,N_70,N_1006);
nor U1444 (N_1444,N_1234,N_54);
xnor U1445 (N_1445,N_834,N_549);
nand U1446 (N_1446,N_1161,N_433);
nor U1447 (N_1447,N_621,N_894);
or U1448 (N_1448,N_531,N_673);
nand U1449 (N_1449,N_613,N_989);
and U1450 (N_1450,N_541,N_1009);
nor U1451 (N_1451,N_378,N_857);
nand U1452 (N_1452,N_91,N_478);
nand U1453 (N_1453,N_1076,N_108);
xor U1454 (N_1454,N_755,N_445);
nand U1455 (N_1455,N_874,N_410);
or U1456 (N_1456,N_680,N_264);
and U1457 (N_1457,N_661,N_781);
nand U1458 (N_1458,N_131,N_650);
nand U1459 (N_1459,N_425,N_766);
nand U1460 (N_1460,N_723,N_971);
or U1461 (N_1461,N_643,N_146);
nand U1462 (N_1462,N_18,N_813);
nand U1463 (N_1463,N_1224,N_1037);
nor U1464 (N_1464,N_188,N_430);
or U1465 (N_1465,N_423,N_931);
xor U1466 (N_1466,N_447,N_772);
nor U1467 (N_1467,N_483,N_802);
nor U1468 (N_1468,N_284,N_881);
nor U1469 (N_1469,N_489,N_912);
or U1470 (N_1470,N_1112,N_77);
nand U1471 (N_1471,N_721,N_193);
and U1472 (N_1472,N_29,N_150);
nand U1473 (N_1473,N_419,N_214);
xor U1474 (N_1474,N_32,N_241);
and U1475 (N_1475,N_1213,N_558);
xnor U1476 (N_1476,N_952,N_811);
and U1477 (N_1477,N_600,N_164);
or U1478 (N_1478,N_190,N_60);
nor U1479 (N_1479,N_1225,N_364);
xor U1480 (N_1480,N_1128,N_1029);
xor U1481 (N_1481,N_1206,N_261);
xor U1482 (N_1482,N_1117,N_1132);
nand U1483 (N_1483,N_259,N_387);
nor U1484 (N_1484,N_602,N_1200);
xor U1485 (N_1485,N_189,N_984);
xor U1486 (N_1486,N_454,N_325);
nand U1487 (N_1487,N_846,N_207);
nand U1488 (N_1488,N_457,N_25);
nor U1489 (N_1489,N_103,N_1071);
xor U1490 (N_1490,N_1164,N_151);
or U1491 (N_1491,N_1172,N_407);
or U1492 (N_1492,N_205,N_969);
nor U1493 (N_1493,N_1129,N_22);
nand U1494 (N_1494,N_861,N_562);
xnor U1495 (N_1495,N_1011,N_438);
and U1496 (N_1496,N_731,N_745);
or U1497 (N_1497,N_918,N_83);
or U1498 (N_1498,N_883,N_1120);
and U1499 (N_1499,N_539,N_337);
nor U1500 (N_1500,N_771,N_374);
and U1501 (N_1501,N_911,N_168);
or U1502 (N_1502,N_769,N_137);
or U1503 (N_1503,N_851,N_932);
nand U1504 (N_1504,N_30,N_626);
and U1505 (N_1505,N_76,N_276);
and U1506 (N_1506,N_1103,N_1201);
and U1507 (N_1507,N_668,N_982);
nor U1508 (N_1508,N_228,N_972);
nor U1509 (N_1509,N_331,N_561);
nand U1510 (N_1510,N_807,N_195);
or U1511 (N_1511,N_1095,N_497);
nand U1512 (N_1512,N_86,N_1204);
or U1513 (N_1513,N_996,N_452);
nand U1514 (N_1514,N_19,N_1114);
xnor U1515 (N_1515,N_232,N_114);
and U1516 (N_1516,N_238,N_1175);
nand U1517 (N_1517,N_814,N_254);
and U1518 (N_1518,N_985,N_87);
and U1519 (N_1519,N_957,N_522);
and U1520 (N_1520,N_172,N_1038);
and U1521 (N_1521,N_618,N_907);
nor U1522 (N_1522,N_697,N_1236);
nor U1523 (N_1523,N_1182,N_1162);
nand U1524 (N_1524,N_836,N_916);
nand U1525 (N_1525,N_1221,N_1057);
nand U1526 (N_1526,N_701,N_729);
and U1527 (N_1527,N_175,N_377);
nand U1528 (N_1528,N_118,N_136);
xor U1529 (N_1529,N_608,N_1105);
and U1530 (N_1530,N_1191,N_1012);
or U1531 (N_1531,N_502,N_277);
nor U1532 (N_1532,N_1147,N_625);
and U1533 (N_1533,N_341,N_825);
or U1534 (N_1534,N_646,N_649);
and U1535 (N_1535,N_965,N_268);
and U1536 (N_1536,N_1222,N_533);
xor U1537 (N_1537,N_1219,N_1155);
nor U1538 (N_1538,N_573,N_1042);
or U1539 (N_1539,N_303,N_1177);
nor U1540 (N_1540,N_708,N_840);
xor U1541 (N_1541,N_434,N_880);
xor U1542 (N_1542,N_645,N_124);
xor U1543 (N_1543,N_142,N_796);
or U1544 (N_1544,N_707,N_37);
xor U1545 (N_1545,N_320,N_652);
xor U1546 (N_1546,N_667,N_944);
or U1547 (N_1547,N_628,N_1060);
xnor U1548 (N_1548,N_314,N_691);
xnor U1549 (N_1549,N_1183,N_1123);
xor U1550 (N_1550,N_291,N_826);
xor U1551 (N_1551,N_988,N_1217);
and U1552 (N_1552,N_681,N_991);
xnor U1553 (N_1553,N_754,N_1211);
nor U1554 (N_1554,N_344,N_16);
nand U1555 (N_1555,N_867,N_583);
xor U1556 (N_1556,N_597,N_554);
and U1557 (N_1557,N_1150,N_233);
nor U1558 (N_1558,N_290,N_578);
xnor U1559 (N_1559,N_828,N_902);
nand U1560 (N_1560,N_616,N_20);
xnor U1561 (N_1561,N_327,N_491);
nand U1562 (N_1562,N_1230,N_160);
nor U1563 (N_1563,N_370,N_530);
or U1564 (N_1564,N_84,N_1000);
and U1565 (N_1565,N_1241,N_930);
nand U1566 (N_1566,N_835,N_1031);
and U1567 (N_1567,N_1110,N_1016);
nor U1568 (N_1568,N_305,N_664);
nand U1569 (N_1569,N_1089,N_1205);
nor U1570 (N_1570,N_134,N_226);
or U1571 (N_1571,N_660,N_630);
nand U1572 (N_1572,N_1068,N_795);
nor U1573 (N_1573,N_579,N_658);
and U1574 (N_1574,N_1146,N_61);
xnor U1575 (N_1575,N_180,N_21);
nand U1576 (N_1576,N_973,N_499);
and U1577 (N_1577,N_381,N_128);
nand U1578 (N_1578,N_200,N_975);
nand U1579 (N_1579,N_693,N_243);
nor U1580 (N_1580,N_498,N_622);
and U1581 (N_1581,N_761,N_316);
nand U1582 (N_1582,N_504,N_852);
or U1583 (N_1583,N_461,N_488);
nor U1584 (N_1584,N_186,N_552);
xor U1585 (N_1585,N_352,N_1207);
or U1586 (N_1586,N_396,N_877);
and U1587 (N_1587,N_390,N_898);
nand U1588 (N_1588,N_730,N_741);
nand U1589 (N_1589,N_689,N_1100);
nand U1590 (N_1590,N_513,N_1030);
xor U1591 (N_1591,N_523,N_1199);
nand U1592 (N_1592,N_1149,N_1186);
and U1593 (N_1593,N_763,N_917);
nor U1594 (N_1594,N_90,N_313);
or U1595 (N_1595,N_1102,N_508);
or U1596 (N_1596,N_1007,N_404);
and U1597 (N_1597,N_44,N_864);
nand U1598 (N_1598,N_821,N_391);
nand U1599 (N_1599,N_806,N_666);
nor U1600 (N_1600,N_1232,N_40);
or U1601 (N_1601,N_398,N_714);
nand U1602 (N_1602,N_856,N_1209);
nor U1603 (N_1603,N_873,N_6);
xnor U1604 (N_1604,N_765,N_1113);
nor U1605 (N_1605,N_1228,N_1131);
nor U1606 (N_1606,N_318,N_1020);
nand U1607 (N_1607,N_682,N_351);
or U1608 (N_1608,N_1059,N_519);
xnor U1609 (N_1609,N_1036,N_638);
nand U1610 (N_1610,N_1178,N_48);
or U1611 (N_1611,N_3,N_951);
and U1612 (N_1612,N_1165,N_592);
or U1613 (N_1613,N_382,N_1210);
nor U1614 (N_1614,N_897,N_863);
and U1615 (N_1615,N_224,N_99);
xnor U1616 (N_1616,N_642,N_555);
nor U1617 (N_1617,N_696,N_808);
nor U1618 (N_1618,N_823,N_669);
xor U1619 (N_1619,N_1054,N_403);
and U1620 (N_1620,N_272,N_321);
or U1621 (N_1621,N_210,N_93);
and U1622 (N_1622,N_1055,N_553);
or U1623 (N_1623,N_853,N_138);
and U1624 (N_1624,N_1115,N_1014);
nand U1625 (N_1625,N_920,N_770);
or U1626 (N_1626,N_891,N_440);
or U1627 (N_1627,N_901,N_1044);
and U1628 (N_1628,N_1080,N_92);
xnor U1629 (N_1629,N_1158,N_1194);
or U1630 (N_1630,N_514,N_612);
and U1631 (N_1631,N_521,N_575);
nand U1632 (N_1632,N_283,N_663);
xnor U1633 (N_1633,N_177,N_202);
nand U1634 (N_1634,N_453,N_648);
or U1635 (N_1635,N_892,N_1108);
xor U1636 (N_1636,N_580,N_749);
xnor U1637 (N_1637,N_983,N_156);
or U1638 (N_1638,N_119,N_1168);
and U1639 (N_1639,N_107,N_235);
nor U1640 (N_1640,N_155,N_435);
nor U1641 (N_1641,N_402,N_505);
nor U1642 (N_1642,N_908,N_623);
nor U1643 (N_1643,N_271,N_9);
xor U1644 (N_1644,N_71,N_323);
nor U1645 (N_1645,N_1004,N_970);
nand U1646 (N_1646,N_954,N_17);
nor U1647 (N_1647,N_1001,N_58);
and U1648 (N_1648,N_468,N_194);
xnor U1649 (N_1649,N_1092,N_1023);
or U1650 (N_1650,N_1070,N_97);
nor U1651 (N_1651,N_4,N_106);
xor U1652 (N_1652,N_311,N_1170);
or U1653 (N_1653,N_604,N_786);
and U1654 (N_1654,N_942,N_80);
or U1655 (N_1655,N_526,N_1227);
nor U1656 (N_1656,N_199,N_248);
nor U1657 (N_1657,N_923,N_803);
and U1658 (N_1658,N_415,N_1239);
nor U1659 (N_1659,N_105,N_482);
and U1660 (N_1660,N_12,N_1198);
nand U1661 (N_1661,N_395,N_1008);
nor U1662 (N_1662,N_966,N_11);
or U1663 (N_1663,N_670,N_41);
and U1664 (N_1664,N_122,N_23);
xor U1665 (N_1665,N_360,N_606);
or U1666 (N_1666,N_46,N_1238);
xnor U1667 (N_1667,N_250,N_605);
nor U1668 (N_1668,N_1,N_123);
or U1669 (N_1669,N_469,N_1085);
or U1670 (N_1670,N_679,N_791);
and U1671 (N_1671,N_981,N_767);
and U1672 (N_1672,N_28,N_1106);
nand U1673 (N_1673,N_7,N_672);
and U1674 (N_1674,N_1215,N_945);
nand U1675 (N_1675,N_572,N_315);
nand U1676 (N_1676,N_258,N_0);
nand U1677 (N_1677,N_1022,N_101);
and U1678 (N_1678,N_1193,N_884);
xnor U1679 (N_1679,N_586,N_246);
and U1680 (N_1680,N_979,N_764);
and U1681 (N_1681,N_286,N_280);
and U1682 (N_1682,N_310,N_1069);
and U1683 (N_1683,N_1138,N_484);
nor U1684 (N_1684,N_750,N_1226);
and U1685 (N_1685,N_158,N_698);
nand U1686 (N_1686,N_900,N_324);
and U1687 (N_1687,N_428,N_637);
nand U1688 (N_1688,N_1086,N_437);
nand U1689 (N_1689,N_793,N_838);
or U1690 (N_1690,N_1208,N_455);
nor U1691 (N_1691,N_929,N_470);
or U1692 (N_1692,N_222,N_216);
nand U1693 (N_1693,N_655,N_798);
nor U1694 (N_1694,N_1053,N_1174);
nor U1695 (N_1695,N_850,N_1063);
and U1696 (N_1696,N_910,N_239);
nand U1697 (N_1697,N_135,N_726);
nor U1698 (N_1698,N_133,N_417);
nor U1699 (N_1699,N_231,N_237);
and U1700 (N_1700,N_413,N_55);
and U1701 (N_1701,N_865,N_1021);
xor U1702 (N_1702,N_596,N_1140);
nand U1703 (N_1703,N_24,N_563);
and U1704 (N_1704,N_81,N_956);
and U1705 (N_1705,N_209,N_1181);
or U1706 (N_1706,N_703,N_665);
or U1707 (N_1707,N_773,N_1163);
or U1708 (N_1708,N_462,N_1125);
or U1709 (N_1709,N_463,N_879);
and U1710 (N_1710,N_1196,N_833);
or U1711 (N_1711,N_571,N_1137);
xnor U1712 (N_1712,N_456,N_227);
nor U1713 (N_1713,N_968,N_1049);
and U1714 (N_1714,N_634,N_273);
and U1715 (N_1715,N_998,N_399);
and U1716 (N_1716,N_1246,N_817);
and U1717 (N_1717,N_566,N_1003);
or U1718 (N_1718,N_854,N_779);
nor U1719 (N_1719,N_317,N_1083);
or U1720 (N_1720,N_1082,N_1116);
nand U1721 (N_1721,N_14,N_986);
nand U1722 (N_1722,N_1019,N_179);
or U1723 (N_1723,N_73,N_1156);
and U1724 (N_1724,N_1237,N_112);
and U1725 (N_1725,N_1065,N_319);
nor U1726 (N_1726,N_1185,N_538);
xor U1727 (N_1727,N_371,N_471);
and U1728 (N_1728,N_933,N_154);
nand U1729 (N_1729,N_38,N_820);
xnor U1730 (N_1730,N_1026,N_736);
and U1731 (N_1731,N_787,N_517);
or U1732 (N_1732,N_740,N_400);
nand U1733 (N_1733,N_776,N_72);
nor U1734 (N_1734,N_876,N_872);
or U1735 (N_1735,N_301,N_659);
and U1736 (N_1736,N_145,N_460);
or U1737 (N_1737,N_1144,N_422);
and U1738 (N_1738,N_939,N_1218);
xor U1739 (N_1739,N_909,N_298);
and U1740 (N_1740,N_185,N_1028);
nor U1741 (N_1741,N_959,N_336);
and U1742 (N_1742,N_805,N_744);
and U1743 (N_1743,N_487,N_230);
or U1744 (N_1744,N_936,N_601);
nand U1745 (N_1745,N_475,N_997);
and U1746 (N_1746,N_978,N_903);
nor U1747 (N_1747,N_51,N_875);
nor U1748 (N_1748,N_559,N_251);
nand U1749 (N_1749,N_52,N_629);
nor U1750 (N_1750,N_705,N_641);
nor U1751 (N_1751,N_412,N_221);
nor U1752 (N_1752,N_426,N_64);
nor U1753 (N_1753,N_727,N_800);
and U1754 (N_1754,N_326,N_244);
or U1755 (N_1755,N_631,N_1154);
nand U1756 (N_1756,N_267,N_1064);
or U1757 (N_1757,N_732,N_335);
xnor U1758 (N_1758,N_477,N_797);
nor U1759 (N_1759,N_1143,N_10);
nor U1760 (N_1760,N_57,N_485);
or U1761 (N_1761,N_368,N_928);
xor U1762 (N_1762,N_695,N_860);
xnor U1763 (N_1763,N_1220,N_1017);
or U1764 (N_1764,N_449,N_147);
or U1765 (N_1765,N_844,N_405);
and U1766 (N_1766,N_777,N_1104);
xor U1767 (N_1767,N_1098,N_545);
xnor U1768 (N_1768,N_1075,N_113);
nor U1769 (N_1769,N_39,N_624);
and U1770 (N_1770,N_88,N_144);
and U1771 (N_1771,N_1025,N_96);
nand U1772 (N_1772,N_922,N_282);
or U1773 (N_1773,N_1179,N_548);
nand U1774 (N_1774,N_509,N_792);
xnor U1775 (N_1775,N_1084,N_1145);
and U1776 (N_1776,N_518,N_1243);
and U1777 (N_1777,N_446,N_654);
nor U1778 (N_1778,N_436,N_1121);
xnor U1779 (N_1779,N_1235,N_564);
nand U1780 (N_1780,N_159,N_132);
nor U1781 (N_1781,N_815,N_746);
and U1782 (N_1782,N_1072,N_309);
nand U1783 (N_1783,N_300,N_1051);
and U1784 (N_1784,N_263,N_278);
nand U1785 (N_1785,N_537,N_890);
xnor U1786 (N_1786,N_153,N_467);
or U1787 (N_1787,N_742,N_94);
and U1788 (N_1788,N_1203,N_785);
nand U1789 (N_1789,N_574,N_260);
nand U1790 (N_1790,N_747,N_1184);
or U1791 (N_1791,N_411,N_713);
nor U1792 (N_1792,N_458,N_406);
or U1793 (N_1793,N_512,N_651);
xor U1794 (N_1794,N_143,N_242);
nor U1795 (N_1795,N_799,N_593);
or U1796 (N_1796,N_204,N_500);
nor U1797 (N_1797,N_611,N_581);
or U1798 (N_1798,N_1067,N_354);
and U1799 (N_1799,N_1018,N_926);
and U1800 (N_1800,N_312,N_743);
or U1801 (N_1801,N_247,N_768);
xnor U1802 (N_1802,N_774,N_472);
or U1803 (N_1803,N_728,N_1151);
and U1804 (N_1804,N_717,N_206);
and U1805 (N_1805,N_493,N_869);
nand U1806 (N_1806,N_345,N_63);
or U1807 (N_1807,N_240,N_480);
and U1808 (N_1808,N_270,N_56);
xnor U1809 (N_1809,N_841,N_464);
and U1810 (N_1810,N_1122,N_960);
or U1811 (N_1811,N_507,N_839);
nor U1812 (N_1812,N_308,N_832);
nor U1813 (N_1813,N_181,N_535);
and U1814 (N_1814,N_201,N_1192);
or U1815 (N_1815,N_515,N_1245);
and U1816 (N_1816,N_1197,N_812);
xor U1817 (N_1817,N_1090,N_1223);
or U1818 (N_1818,N_427,N_53);
and U1819 (N_1819,N_182,N_95);
nand U1820 (N_1820,N_632,N_543);
or U1821 (N_1821,N_141,N_401);
or U1822 (N_1822,N_126,N_424);
or U1823 (N_1823,N_677,N_1233);
or U1824 (N_1824,N_363,N_831);
or U1825 (N_1825,N_104,N_678);
and U1826 (N_1826,N_176,N_416);
and U1827 (N_1827,N_524,N_720);
xnor U1828 (N_1828,N_653,N_532);
or U1829 (N_1829,N_393,N_355);
xnor U1830 (N_1830,N_845,N_163);
nor U1831 (N_1831,N_383,N_1160);
or U1832 (N_1832,N_1033,N_1091);
xor U1833 (N_1833,N_252,N_878);
or U1834 (N_1834,N_688,N_751);
nand U1835 (N_1835,N_591,N_1136);
nor U1836 (N_1836,N_129,N_330);
nor U1837 (N_1837,N_236,N_443);
nor U1838 (N_1838,N_516,N_1041);
nand U1839 (N_1839,N_35,N_1148);
xor U1840 (N_1840,N_1171,N_306);
nand U1841 (N_1841,N_257,N_692);
xnor U1842 (N_1842,N_219,N_609);
xnor U1843 (N_1843,N_304,N_980);
nand U1844 (N_1844,N_1169,N_1107);
and U1845 (N_1845,N_818,N_342);
or U1846 (N_1846,N_296,N_191);
and U1847 (N_1847,N_690,N_388);
or U1848 (N_1848,N_870,N_486);
xor U1849 (N_1849,N_102,N_962);
or U1850 (N_1850,N_627,N_266);
xnor U1851 (N_1851,N_1005,N_121);
and U1852 (N_1852,N_1032,N_13);
or U1853 (N_1853,N_595,N_974);
nor U1854 (N_1854,N_1093,N_1166);
nand U1855 (N_1855,N_1099,N_778);
nand U1856 (N_1856,N_819,N_529);
or U1857 (N_1857,N_967,N_197);
and U1858 (N_1858,N_1024,N_1188);
or U1859 (N_1859,N_783,N_550);
nand U1860 (N_1860,N_994,N_937);
nor U1861 (N_1861,N_528,N_408);
nand U1862 (N_1862,N_208,N_585);
nand U1863 (N_1863,N_1040,N_2);
and U1864 (N_1864,N_976,N_117);
nor U1865 (N_1865,N_610,N_451);
nor U1866 (N_1866,N_1052,N_359);
nor U1867 (N_1867,N_1231,N_587);
and U1868 (N_1868,N_1153,N_794);
xor U1869 (N_1869,N_481,N_674);
and U1870 (N_1870,N_782,N_1066);
xnor U1871 (N_1871,N_380,N_914);
and U1872 (N_1872,N_1212,N_1141);
or U1873 (N_1873,N_171,N_111);
nor U1874 (N_1874,N_990,N_904);
and U1875 (N_1875,N_1176,N_778);
nor U1876 (N_1876,N_1167,N_298);
xor U1877 (N_1877,N_749,N_325);
and U1878 (N_1878,N_901,N_292);
nand U1879 (N_1879,N_630,N_100);
nor U1880 (N_1880,N_1217,N_16);
and U1881 (N_1881,N_433,N_247);
xor U1882 (N_1882,N_612,N_586);
and U1883 (N_1883,N_274,N_289);
nand U1884 (N_1884,N_811,N_985);
xor U1885 (N_1885,N_273,N_1038);
xor U1886 (N_1886,N_779,N_182);
and U1887 (N_1887,N_474,N_516);
nand U1888 (N_1888,N_1007,N_60);
xor U1889 (N_1889,N_246,N_637);
and U1890 (N_1890,N_1130,N_1104);
nand U1891 (N_1891,N_949,N_121);
nor U1892 (N_1892,N_773,N_54);
nor U1893 (N_1893,N_715,N_343);
xor U1894 (N_1894,N_527,N_168);
nor U1895 (N_1895,N_324,N_414);
nor U1896 (N_1896,N_102,N_183);
nand U1897 (N_1897,N_1095,N_592);
xor U1898 (N_1898,N_639,N_353);
nand U1899 (N_1899,N_216,N_1229);
or U1900 (N_1900,N_644,N_101);
nand U1901 (N_1901,N_997,N_1088);
nor U1902 (N_1902,N_990,N_88);
or U1903 (N_1903,N_719,N_699);
and U1904 (N_1904,N_96,N_1218);
and U1905 (N_1905,N_1074,N_116);
or U1906 (N_1906,N_720,N_1059);
nand U1907 (N_1907,N_1040,N_891);
nor U1908 (N_1908,N_868,N_680);
xnor U1909 (N_1909,N_1187,N_796);
xor U1910 (N_1910,N_115,N_641);
or U1911 (N_1911,N_775,N_1178);
xor U1912 (N_1912,N_1175,N_798);
or U1913 (N_1913,N_1100,N_691);
and U1914 (N_1914,N_26,N_1064);
and U1915 (N_1915,N_1020,N_9);
or U1916 (N_1916,N_46,N_740);
nand U1917 (N_1917,N_346,N_291);
nor U1918 (N_1918,N_1150,N_735);
or U1919 (N_1919,N_442,N_910);
and U1920 (N_1920,N_686,N_1075);
or U1921 (N_1921,N_107,N_55);
nor U1922 (N_1922,N_399,N_77);
or U1923 (N_1923,N_213,N_686);
nand U1924 (N_1924,N_23,N_689);
nand U1925 (N_1925,N_811,N_1160);
nand U1926 (N_1926,N_731,N_842);
xor U1927 (N_1927,N_571,N_1168);
nor U1928 (N_1928,N_393,N_577);
nand U1929 (N_1929,N_701,N_895);
xnor U1930 (N_1930,N_755,N_1147);
nor U1931 (N_1931,N_520,N_352);
nand U1932 (N_1932,N_277,N_328);
and U1933 (N_1933,N_412,N_1165);
xor U1934 (N_1934,N_48,N_600);
nor U1935 (N_1935,N_689,N_32);
and U1936 (N_1936,N_1146,N_928);
nor U1937 (N_1937,N_778,N_974);
and U1938 (N_1938,N_670,N_990);
xor U1939 (N_1939,N_353,N_1233);
or U1940 (N_1940,N_728,N_797);
and U1941 (N_1941,N_1050,N_95);
nand U1942 (N_1942,N_948,N_780);
nand U1943 (N_1943,N_458,N_210);
or U1944 (N_1944,N_456,N_715);
and U1945 (N_1945,N_942,N_830);
xor U1946 (N_1946,N_1108,N_1047);
nor U1947 (N_1947,N_723,N_276);
or U1948 (N_1948,N_134,N_252);
or U1949 (N_1949,N_483,N_703);
and U1950 (N_1950,N_999,N_124);
xnor U1951 (N_1951,N_53,N_1191);
xnor U1952 (N_1952,N_656,N_1219);
or U1953 (N_1953,N_1148,N_1223);
nor U1954 (N_1954,N_823,N_555);
or U1955 (N_1955,N_185,N_1035);
xnor U1956 (N_1956,N_288,N_1221);
nor U1957 (N_1957,N_413,N_424);
nand U1958 (N_1958,N_1018,N_349);
or U1959 (N_1959,N_974,N_106);
xor U1960 (N_1960,N_1193,N_435);
nor U1961 (N_1961,N_1219,N_346);
xor U1962 (N_1962,N_173,N_1063);
or U1963 (N_1963,N_884,N_906);
or U1964 (N_1964,N_550,N_627);
and U1965 (N_1965,N_814,N_46);
nor U1966 (N_1966,N_194,N_316);
and U1967 (N_1967,N_400,N_813);
nand U1968 (N_1968,N_424,N_461);
and U1969 (N_1969,N_1130,N_674);
xnor U1970 (N_1970,N_805,N_642);
and U1971 (N_1971,N_489,N_555);
xor U1972 (N_1972,N_1076,N_163);
nand U1973 (N_1973,N_1013,N_516);
nor U1974 (N_1974,N_523,N_337);
and U1975 (N_1975,N_44,N_419);
nor U1976 (N_1976,N_427,N_356);
or U1977 (N_1977,N_984,N_171);
nor U1978 (N_1978,N_916,N_1063);
or U1979 (N_1979,N_413,N_1030);
and U1980 (N_1980,N_336,N_782);
nor U1981 (N_1981,N_916,N_304);
nor U1982 (N_1982,N_481,N_604);
or U1983 (N_1983,N_43,N_1143);
nand U1984 (N_1984,N_472,N_1103);
nor U1985 (N_1985,N_121,N_1146);
and U1986 (N_1986,N_733,N_237);
nand U1987 (N_1987,N_1001,N_815);
nand U1988 (N_1988,N_925,N_809);
xor U1989 (N_1989,N_1027,N_56);
nand U1990 (N_1990,N_457,N_1018);
nor U1991 (N_1991,N_496,N_187);
or U1992 (N_1992,N_1003,N_1160);
and U1993 (N_1993,N_852,N_969);
xor U1994 (N_1994,N_424,N_875);
nor U1995 (N_1995,N_49,N_295);
nor U1996 (N_1996,N_757,N_38);
nor U1997 (N_1997,N_993,N_563);
nand U1998 (N_1998,N_923,N_681);
and U1999 (N_1999,N_292,N_597);
or U2000 (N_2000,N_251,N_957);
nand U2001 (N_2001,N_1047,N_306);
nor U2002 (N_2002,N_533,N_116);
nand U2003 (N_2003,N_263,N_484);
nand U2004 (N_2004,N_1082,N_24);
or U2005 (N_2005,N_841,N_1027);
xnor U2006 (N_2006,N_269,N_830);
or U2007 (N_2007,N_1195,N_88);
xor U2008 (N_2008,N_173,N_998);
nand U2009 (N_2009,N_285,N_663);
nand U2010 (N_2010,N_1243,N_1072);
nand U2011 (N_2011,N_747,N_264);
nor U2012 (N_2012,N_1135,N_745);
and U2013 (N_2013,N_818,N_170);
nor U2014 (N_2014,N_903,N_204);
nand U2015 (N_2015,N_966,N_122);
or U2016 (N_2016,N_554,N_334);
nor U2017 (N_2017,N_870,N_959);
nor U2018 (N_2018,N_293,N_703);
nand U2019 (N_2019,N_104,N_81);
nand U2020 (N_2020,N_142,N_188);
or U2021 (N_2021,N_753,N_1064);
nand U2022 (N_2022,N_679,N_123);
xor U2023 (N_2023,N_520,N_805);
xor U2024 (N_2024,N_801,N_1193);
nand U2025 (N_2025,N_1055,N_463);
nor U2026 (N_2026,N_987,N_79);
nand U2027 (N_2027,N_243,N_1183);
nand U2028 (N_2028,N_1244,N_861);
and U2029 (N_2029,N_185,N_568);
and U2030 (N_2030,N_225,N_736);
xnor U2031 (N_2031,N_422,N_1142);
nor U2032 (N_2032,N_47,N_531);
nand U2033 (N_2033,N_35,N_1179);
xor U2034 (N_2034,N_1240,N_346);
nand U2035 (N_2035,N_357,N_904);
xor U2036 (N_2036,N_299,N_601);
or U2037 (N_2037,N_620,N_341);
nand U2038 (N_2038,N_786,N_151);
or U2039 (N_2039,N_860,N_632);
nor U2040 (N_2040,N_568,N_494);
or U2041 (N_2041,N_1089,N_615);
nand U2042 (N_2042,N_1150,N_264);
xnor U2043 (N_2043,N_947,N_73);
or U2044 (N_2044,N_74,N_197);
xor U2045 (N_2045,N_74,N_177);
and U2046 (N_2046,N_988,N_238);
xor U2047 (N_2047,N_216,N_589);
and U2048 (N_2048,N_979,N_74);
or U2049 (N_2049,N_380,N_1164);
and U2050 (N_2050,N_908,N_873);
nand U2051 (N_2051,N_524,N_1034);
xnor U2052 (N_2052,N_729,N_609);
or U2053 (N_2053,N_1005,N_106);
or U2054 (N_2054,N_367,N_582);
or U2055 (N_2055,N_485,N_154);
nor U2056 (N_2056,N_35,N_1009);
and U2057 (N_2057,N_50,N_135);
nand U2058 (N_2058,N_1037,N_936);
or U2059 (N_2059,N_814,N_1047);
or U2060 (N_2060,N_163,N_396);
and U2061 (N_2061,N_7,N_214);
or U2062 (N_2062,N_320,N_824);
xor U2063 (N_2063,N_918,N_1153);
and U2064 (N_2064,N_636,N_119);
or U2065 (N_2065,N_931,N_379);
nor U2066 (N_2066,N_1030,N_600);
nand U2067 (N_2067,N_489,N_206);
nand U2068 (N_2068,N_1216,N_164);
nand U2069 (N_2069,N_321,N_205);
and U2070 (N_2070,N_1156,N_544);
and U2071 (N_2071,N_736,N_247);
xor U2072 (N_2072,N_240,N_1066);
or U2073 (N_2073,N_976,N_298);
xor U2074 (N_2074,N_922,N_499);
xnor U2075 (N_2075,N_659,N_1205);
or U2076 (N_2076,N_598,N_773);
nor U2077 (N_2077,N_566,N_1182);
or U2078 (N_2078,N_160,N_549);
and U2079 (N_2079,N_854,N_1188);
nand U2080 (N_2080,N_854,N_855);
and U2081 (N_2081,N_200,N_229);
and U2082 (N_2082,N_1197,N_988);
xnor U2083 (N_2083,N_99,N_265);
xor U2084 (N_2084,N_1029,N_1077);
xnor U2085 (N_2085,N_984,N_1172);
or U2086 (N_2086,N_166,N_852);
and U2087 (N_2087,N_214,N_690);
nor U2088 (N_2088,N_477,N_754);
and U2089 (N_2089,N_371,N_95);
or U2090 (N_2090,N_769,N_558);
nand U2091 (N_2091,N_1138,N_339);
and U2092 (N_2092,N_909,N_377);
xor U2093 (N_2093,N_556,N_733);
and U2094 (N_2094,N_395,N_1044);
or U2095 (N_2095,N_47,N_956);
xor U2096 (N_2096,N_1167,N_393);
and U2097 (N_2097,N_873,N_11);
nor U2098 (N_2098,N_1051,N_1049);
or U2099 (N_2099,N_854,N_424);
nor U2100 (N_2100,N_779,N_1030);
xnor U2101 (N_2101,N_779,N_164);
and U2102 (N_2102,N_790,N_526);
or U2103 (N_2103,N_437,N_980);
nand U2104 (N_2104,N_885,N_29);
or U2105 (N_2105,N_108,N_569);
nor U2106 (N_2106,N_252,N_43);
nor U2107 (N_2107,N_401,N_428);
nor U2108 (N_2108,N_551,N_908);
nor U2109 (N_2109,N_1083,N_789);
nor U2110 (N_2110,N_725,N_901);
nor U2111 (N_2111,N_883,N_716);
or U2112 (N_2112,N_998,N_294);
or U2113 (N_2113,N_82,N_1013);
nor U2114 (N_2114,N_440,N_525);
and U2115 (N_2115,N_252,N_213);
nand U2116 (N_2116,N_975,N_1248);
nor U2117 (N_2117,N_122,N_629);
xnor U2118 (N_2118,N_908,N_624);
nand U2119 (N_2119,N_826,N_1077);
xnor U2120 (N_2120,N_888,N_464);
nand U2121 (N_2121,N_1007,N_90);
nand U2122 (N_2122,N_378,N_441);
or U2123 (N_2123,N_1005,N_1152);
nor U2124 (N_2124,N_868,N_855);
and U2125 (N_2125,N_809,N_941);
nand U2126 (N_2126,N_360,N_1111);
xnor U2127 (N_2127,N_595,N_1188);
and U2128 (N_2128,N_905,N_1213);
xnor U2129 (N_2129,N_499,N_1176);
and U2130 (N_2130,N_222,N_619);
nand U2131 (N_2131,N_1152,N_14);
nand U2132 (N_2132,N_967,N_933);
nor U2133 (N_2133,N_975,N_199);
nor U2134 (N_2134,N_589,N_558);
nand U2135 (N_2135,N_589,N_291);
xnor U2136 (N_2136,N_1124,N_271);
or U2137 (N_2137,N_874,N_580);
xnor U2138 (N_2138,N_458,N_879);
nor U2139 (N_2139,N_581,N_836);
xor U2140 (N_2140,N_493,N_315);
or U2141 (N_2141,N_1120,N_199);
nand U2142 (N_2142,N_645,N_588);
nand U2143 (N_2143,N_417,N_14);
nand U2144 (N_2144,N_1070,N_1237);
and U2145 (N_2145,N_655,N_855);
nor U2146 (N_2146,N_1211,N_305);
nand U2147 (N_2147,N_805,N_722);
nor U2148 (N_2148,N_919,N_1192);
or U2149 (N_2149,N_443,N_1133);
nand U2150 (N_2150,N_980,N_270);
or U2151 (N_2151,N_867,N_351);
xor U2152 (N_2152,N_677,N_146);
nand U2153 (N_2153,N_693,N_1204);
xnor U2154 (N_2154,N_689,N_217);
nand U2155 (N_2155,N_795,N_1232);
and U2156 (N_2156,N_175,N_38);
nor U2157 (N_2157,N_922,N_834);
and U2158 (N_2158,N_666,N_478);
nand U2159 (N_2159,N_681,N_113);
nor U2160 (N_2160,N_448,N_688);
nor U2161 (N_2161,N_112,N_848);
or U2162 (N_2162,N_301,N_8);
nand U2163 (N_2163,N_228,N_46);
and U2164 (N_2164,N_890,N_736);
nand U2165 (N_2165,N_333,N_731);
nor U2166 (N_2166,N_1106,N_211);
and U2167 (N_2167,N_1197,N_1032);
and U2168 (N_2168,N_178,N_351);
nand U2169 (N_2169,N_349,N_1084);
and U2170 (N_2170,N_453,N_765);
nand U2171 (N_2171,N_417,N_356);
nor U2172 (N_2172,N_811,N_939);
nor U2173 (N_2173,N_1031,N_1180);
nor U2174 (N_2174,N_1116,N_1241);
and U2175 (N_2175,N_1144,N_1075);
and U2176 (N_2176,N_851,N_1062);
xor U2177 (N_2177,N_589,N_187);
nor U2178 (N_2178,N_642,N_418);
nor U2179 (N_2179,N_505,N_902);
nor U2180 (N_2180,N_72,N_925);
nand U2181 (N_2181,N_1070,N_1000);
nor U2182 (N_2182,N_228,N_1142);
or U2183 (N_2183,N_953,N_717);
and U2184 (N_2184,N_340,N_766);
xnor U2185 (N_2185,N_1242,N_962);
xor U2186 (N_2186,N_345,N_341);
and U2187 (N_2187,N_1173,N_135);
xnor U2188 (N_2188,N_260,N_449);
xor U2189 (N_2189,N_1248,N_1199);
nor U2190 (N_2190,N_248,N_956);
or U2191 (N_2191,N_147,N_624);
or U2192 (N_2192,N_1031,N_662);
nor U2193 (N_2193,N_591,N_220);
nor U2194 (N_2194,N_450,N_557);
xor U2195 (N_2195,N_399,N_1150);
xnor U2196 (N_2196,N_178,N_531);
xor U2197 (N_2197,N_303,N_345);
or U2198 (N_2198,N_1039,N_720);
nand U2199 (N_2199,N_554,N_1163);
and U2200 (N_2200,N_638,N_956);
or U2201 (N_2201,N_493,N_465);
or U2202 (N_2202,N_336,N_715);
and U2203 (N_2203,N_125,N_220);
or U2204 (N_2204,N_146,N_822);
xor U2205 (N_2205,N_1079,N_104);
and U2206 (N_2206,N_346,N_1249);
xor U2207 (N_2207,N_409,N_1161);
and U2208 (N_2208,N_1218,N_663);
nand U2209 (N_2209,N_969,N_698);
nand U2210 (N_2210,N_1122,N_381);
or U2211 (N_2211,N_563,N_135);
and U2212 (N_2212,N_966,N_1031);
and U2213 (N_2213,N_1007,N_367);
or U2214 (N_2214,N_215,N_166);
nor U2215 (N_2215,N_955,N_136);
or U2216 (N_2216,N_750,N_90);
nand U2217 (N_2217,N_1204,N_164);
and U2218 (N_2218,N_1187,N_591);
or U2219 (N_2219,N_837,N_1129);
xor U2220 (N_2220,N_310,N_186);
or U2221 (N_2221,N_708,N_701);
and U2222 (N_2222,N_1020,N_994);
nand U2223 (N_2223,N_347,N_222);
nor U2224 (N_2224,N_824,N_1140);
xor U2225 (N_2225,N_890,N_35);
nand U2226 (N_2226,N_571,N_118);
nand U2227 (N_2227,N_1175,N_38);
nand U2228 (N_2228,N_994,N_794);
nor U2229 (N_2229,N_1090,N_74);
nor U2230 (N_2230,N_560,N_66);
and U2231 (N_2231,N_519,N_251);
and U2232 (N_2232,N_57,N_417);
and U2233 (N_2233,N_284,N_772);
and U2234 (N_2234,N_107,N_196);
xor U2235 (N_2235,N_797,N_806);
and U2236 (N_2236,N_645,N_0);
or U2237 (N_2237,N_531,N_468);
and U2238 (N_2238,N_402,N_603);
or U2239 (N_2239,N_1060,N_21);
xnor U2240 (N_2240,N_377,N_35);
xnor U2241 (N_2241,N_1021,N_921);
nor U2242 (N_2242,N_552,N_309);
and U2243 (N_2243,N_1056,N_682);
nand U2244 (N_2244,N_1043,N_821);
and U2245 (N_2245,N_223,N_525);
nand U2246 (N_2246,N_65,N_822);
xor U2247 (N_2247,N_844,N_554);
and U2248 (N_2248,N_194,N_766);
nand U2249 (N_2249,N_72,N_729);
nor U2250 (N_2250,N_882,N_217);
or U2251 (N_2251,N_1231,N_1128);
nor U2252 (N_2252,N_1020,N_723);
xnor U2253 (N_2253,N_296,N_984);
or U2254 (N_2254,N_741,N_180);
or U2255 (N_2255,N_344,N_589);
nor U2256 (N_2256,N_315,N_217);
and U2257 (N_2257,N_1033,N_947);
nor U2258 (N_2258,N_512,N_740);
nor U2259 (N_2259,N_143,N_756);
nand U2260 (N_2260,N_514,N_1113);
nand U2261 (N_2261,N_314,N_950);
or U2262 (N_2262,N_979,N_771);
and U2263 (N_2263,N_317,N_701);
xnor U2264 (N_2264,N_892,N_39);
xor U2265 (N_2265,N_833,N_1096);
nand U2266 (N_2266,N_965,N_549);
or U2267 (N_2267,N_1162,N_682);
and U2268 (N_2268,N_1030,N_316);
or U2269 (N_2269,N_869,N_107);
and U2270 (N_2270,N_1222,N_1179);
or U2271 (N_2271,N_4,N_664);
xnor U2272 (N_2272,N_704,N_794);
and U2273 (N_2273,N_584,N_242);
nor U2274 (N_2274,N_538,N_595);
or U2275 (N_2275,N_407,N_1189);
xnor U2276 (N_2276,N_1050,N_821);
and U2277 (N_2277,N_540,N_1207);
xnor U2278 (N_2278,N_597,N_832);
and U2279 (N_2279,N_1022,N_315);
nand U2280 (N_2280,N_527,N_1235);
nor U2281 (N_2281,N_1047,N_1212);
nor U2282 (N_2282,N_371,N_531);
or U2283 (N_2283,N_215,N_209);
xor U2284 (N_2284,N_497,N_209);
and U2285 (N_2285,N_224,N_874);
and U2286 (N_2286,N_352,N_904);
nor U2287 (N_2287,N_1126,N_111);
or U2288 (N_2288,N_757,N_1237);
xnor U2289 (N_2289,N_153,N_1238);
and U2290 (N_2290,N_605,N_395);
or U2291 (N_2291,N_353,N_326);
or U2292 (N_2292,N_608,N_46);
xor U2293 (N_2293,N_1069,N_168);
nor U2294 (N_2294,N_971,N_419);
and U2295 (N_2295,N_774,N_321);
or U2296 (N_2296,N_595,N_50);
nand U2297 (N_2297,N_176,N_910);
and U2298 (N_2298,N_1064,N_1035);
or U2299 (N_2299,N_853,N_1182);
nor U2300 (N_2300,N_137,N_671);
nand U2301 (N_2301,N_326,N_889);
nor U2302 (N_2302,N_1101,N_240);
nor U2303 (N_2303,N_436,N_928);
nand U2304 (N_2304,N_1248,N_1126);
nor U2305 (N_2305,N_900,N_1210);
nand U2306 (N_2306,N_258,N_750);
xor U2307 (N_2307,N_884,N_323);
xnor U2308 (N_2308,N_80,N_615);
nand U2309 (N_2309,N_403,N_145);
nor U2310 (N_2310,N_1156,N_598);
nor U2311 (N_2311,N_1124,N_78);
nand U2312 (N_2312,N_325,N_130);
or U2313 (N_2313,N_258,N_700);
or U2314 (N_2314,N_1179,N_105);
or U2315 (N_2315,N_302,N_599);
nor U2316 (N_2316,N_1094,N_389);
xor U2317 (N_2317,N_182,N_649);
xor U2318 (N_2318,N_572,N_625);
or U2319 (N_2319,N_207,N_323);
nand U2320 (N_2320,N_532,N_1001);
or U2321 (N_2321,N_493,N_252);
xnor U2322 (N_2322,N_345,N_1000);
or U2323 (N_2323,N_1099,N_1118);
xor U2324 (N_2324,N_53,N_72);
nor U2325 (N_2325,N_707,N_131);
xor U2326 (N_2326,N_645,N_531);
nand U2327 (N_2327,N_36,N_1229);
xor U2328 (N_2328,N_313,N_790);
xor U2329 (N_2329,N_583,N_802);
xor U2330 (N_2330,N_954,N_642);
xor U2331 (N_2331,N_751,N_712);
xnor U2332 (N_2332,N_980,N_55);
or U2333 (N_2333,N_792,N_1239);
or U2334 (N_2334,N_47,N_645);
and U2335 (N_2335,N_1136,N_574);
and U2336 (N_2336,N_543,N_584);
xor U2337 (N_2337,N_962,N_140);
xor U2338 (N_2338,N_1205,N_820);
or U2339 (N_2339,N_153,N_285);
nor U2340 (N_2340,N_2,N_1058);
xor U2341 (N_2341,N_382,N_44);
nor U2342 (N_2342,N_825,N_445);
nor U2343 (N_2343,N_325,N_878);
or U2344 (N_2344,N_687,N_508);
and U2345 (N_2345,N_486,N_841);
xor U2346 (N_2346,N_47,N_949);
or U2347 (N_2347,N_971,N_295);
nand U2348 (N_2348,N_784,N_142);
or U2349 (N_2349,N_899,N_41);
xnor U2350 (N_2350,N_1191,N_938);
nand U2351 (N_2351,N_1058,N_614);
nor U2352 (N_2352,N_675,N_725);
nor U2353 (N_2353,N_444,N_1103);
and U2354 (N_2354,N_254,N_449);
or U2355 (N_2355,N_208,N_887);
or U2356 (N_2356,N_735,N_1106);
xnor U2357 (N_2357,N_69,N_114);
xnor U2358 (N_2358,N_948,N_457);
nor U2359 (N_2359,N_796,N_1140);
xnor U2360 (N_2360,N_1017,N_228);
nand U2361 (N_2361,N_889,N_118);
xnor U2362 (N_2362,N_140,N_1224);
xor U2363 (N_2363,N_163,N_51);
xor U2364 (N_2364,N_61,N_188);
and U2365 (N_2365,N_667,N_1188);
or U2366 (N_2366,N_232,N_398);
and U2367 (N_2367,N_1075,N_587);
or U2368 (N_2368,N_1097,N_127);
or U2369 (N_2369,N_494,N_318);
or U2370 (N_2370,N_1144,N_420);
nor U2371 (N_2371,N_868,N_719);
or U2372 (N_2372,N_1249,N_719);
nand U2373 (N_2373,N_1245,N_864);
and U2374 (N_2374,N_43,N_161);
xnor U2375 (N_2375,N_547,N_370);
nor U2376 (N_2376,N_913,N_302);
and U2377 (N_2377,N_554,N_673);
nand U2378 (N_2378,N_138,N_800);
and U2379 (N_2379,N_866,N_1157);
nor U2380 (N_2380,N_656,N_1067);
and U2381 (N_2381,N_1208,N_653);
and U2382 (N_2382,N_556,N_1112);
or U2383 (N_2383,N_465,N_543);
or U2384 (N_2384,N_1042,N_1059);
and U2385 (N_2385,N_1234,N_801);
xor U2386 (N_2386,N_717,N_178);
and U2387 (N_2387,N_2,N_591);
nand U2388 (N_2388,N_404,N_482);
nor U2389 (N_2389,N_1177,N_813);
nor U2390 (N_2390,N_1153,N_498);
xnor U2391 (N_2391,N_1084,N_859);
and U2392 (N_2392,N_18,N_1197);
nor U2393 (N_2393,N_372,N_743);
nor U2394 (N_2394,N_645,N_861);
and U2395 (N_2395,N_850,N_455);
xor U2396 (N_2396,N_1165,N_114);
xor U2397 (N_2397,N_504,N_673);
or U2398 (N_2398,N_231,N_429);
nand U2399 (N_2399,N_1208,N_817);
or U2400 (N_2400,N_1041,N_870);
nor U2401 (N_2401,N_341,N_655);
and U2402 (N_2402,N_1033,N_253);
xnor U2403 (N_2403,N_981,N_939);
and U2404 (N_2404,N_582,N_754);
xor U2405 (N_2405,N_440,N_184);
nor U2406 (N_2406,N_82,N_658);
nor U2407 (N_2407,N_503,N_40);
and U2408 (N_2408,N_759,N_640);
nor U2409 (N_2409,N_183,N_1168);
nor U2410 (N_2410,N_1188,N_163);
and U2411 (N_2411,N_904,N_534);
nand U2412 (N_2412,N_1249,N_648);
nor U2413 (N_2413,N_387,N_1141);
nor U2414 (N_2414,N_320,N_811);
nand U2415 (N_2415,N_348,N_339);
or U2416 (N_2416,N_238,N_251);
and U2417 (N_2417,N_707,N_307);
xnor U2418 (N_2418,N_1208,N_869);
and U2419 (N_2419,N_77,N_241);
nand U2420 (N_2420,N_813,N_452);
nand U2421 (N_2421,N_829,N_793);
nand U2422 (N_2422,N_1069,N_293);
nor U2423 (N_2423,N_247,N_309);
xor U2424 (N_2424,N_628,N_410);
and U2425 (N_2425,N_607,N_654);
xor U2426 (N_2426,N_1001,N_794);
or U2427 (N_2427,N_820,N_192);
nand U2428 (N_2428,N_492,N_1247);
nand U2429 (N_2429,N_389,N_501);
nand U2430 (N_2430,N_977,N_632);
and U2431 (N_2431,N_796,N_731);
and U2432 (N_2432,N_337,N_576);
nor U2433 (N_2433,N_1018,N_642);
and U2434 (N_2434,N_846,N_873);
nor U2435 (N_2435,N_456,N_613);
nand U2436 (N_2436,N_986,N_272);
or U2437 (N_2437,N_1192,N_1194);
or U2438 (N_2438,N_721,N_2);
and U2439 (N_2439,N_715,N_387);
xor U2440 (N_2440,N_1110,N_598);
xor U2441 (N_2441,N_305,N_480);
or U2442 (N_2442,N_827,N_545);
nor U2443 (N_2443,N_511,N_364);
xor U2444 (N_2444,N_1077,N_745);
xnor U2445 (N_2445,N_297,N_1044);
nand U2446 (N_2446,N_435,N_162);
xor U2447 (N_2447,N_963,N_1076);
or U2448 (N_2448,N_598,N_364);
or U2449 (N_2449,N_137,N_960);
xor U2450 (N_2450,N_466,N_744);
and U2451 (N_2451,N_869,N_862);
xor U2452 (N_2452,N_935,N_869);
and U2453 (N_2453,N_987,N_78);
and U2454 (N_2454,N_32,N_181);
nor U2455 (N_2455,N_850,N_602);
or U2456 (N_2456,N_946,N_876);
and U2457 (N_2457,N_1209,N_1023);
nand U2458 (N_2458,N_212,N_177);
nand U2459 (N_2459,N_868,N_42);
xor U2460 (N_2460,N_1135,N_1079);
nor U2461 (N_2461,N_1172,N_996);
nor U2462 (N_2462,N_984,N_985);
nand U2463 (N_2463,N_574,N_16);
xor U2464 (N_2464,N_428,N_465);
xor U2465 (N_2465,N_237,N_355);
and U2466 (N_2466,N_544,N_735);
nor U2467 (N_2467,N_1201,N_1014);
and U2468 (N_2468,N_149,N_338);
and U2469 (N_2469,N_545,N_389);
nand U2470 (N_2470,N_304,N_270);
nand U2471 (N_2471,N_156,N_559);
xor U2472 (N_2472,N_323,N_942);
nor U2473 (N_2473,N_739,N_805);
and U2474 (N_2474,N_940,N_1146);
or U2475 (N_2475,N_1117,N_217);
nor U2476 (N_2476,N_1038,N_369);
and U2477 (N_2477,N_1094,N_236);
xnor U2478 (N_2478,N_1176,N_43);
nor U2479 (N_2479,N_1122,N_261);
and U2480 (N_2480,N_161,N_987);
and U2481 (N_2481,N_238,N_854);
xnor U2482 (N_2482,N_284,N_352);
nand U2483 (N_2483,N_214,N_997);
xor U2484 (N_2484,N_205,N_249);
nand U2485 (N_2485,N_484,N_223);
xnor U2486 (N_2486,N_443,N_395);
or U2487 (N_2487,N_1078,N_831);
xor U2488 (N_2488,N_472,N_906);
nand U2489 (N_2489,N_210,N_76);
xor U2490 (N_2490,N_610,N_1073);
nand U2491 (N_2491,N_978,N_1159);
nand U2492 (N_2492,N_1167,N_1017);
nand U2493 (N_2493,N_874,N_566);
nand U2494 (N_2494,N_582,N_998);
or U2495 (N_2495,N_1087,N_889);
and U2496 (N_2496,N_231,N_134);
nand U2497 (N_2497,N_338,N_431);
nor U2498 (N_2498,N_733,N_1157);
and U2499 (N_2499,N_35,N_632);
and U2500 (N_2500,N_2427,N_1914);
nor U2501 (N_2501,N_1972,N_1583);
nand U2502 (N_2502,N_1523,N_2243);
nor U2503 (N_2503,N_1760,N_2137);
nor U2504 (N_2504,N_1886,N_2396);
and U2505 (N_2505,N_2343,N_1669);
and U2506 (N_2506,N_1356,N_2469);
or U2507 (N_2507,N_1711,N_1942);
xnor U2508 (N_2508,N_1517,N_1495);
nor U2509 (N_2509,N_1792,N_1395);
nand U2510 (N_2510,N_1414,N_2108);
and U2511 (N_2511,N_2371,N_2058);
nand U2512 (N_2512,N_1407,N_1773);
xor U2513 (N_2513,N_2179,N_1545);
nand U2514 (N_2514,N_2175,N_1320);
xnor U2515 (N_2515,N_2001,N_2277);
or U2516 (N_2516,N_2399,N_1489);
xor U2517 (N_2517,N_1503,N_1349);
nor U2518 (N_2518,N_1866,N_1862);
and U2519 (N_2519,N_1787,N_2235);
or U2520 (N_2520,N_1415,N_2468);
and U2521 (N_2521,N_2122,N_1393);
xnor U2522 (N_2522,N_2486,N_2173);
nand U2523 (N_2523,N_1332,N_2091);
and U2524 (N_2524,N_1507,N_1973);
nand U2525 (N_2525,N_1406,N_2376);
nand U2526 (N_2526,N_1959,N_1739);
nor U2527 (N_2527,N_2286,N_2111);
and U2528 (N_2528,N_1746,N_1893);
nor U2529 (N_2529,N_1537,N_2156);
xnor U2530 (N_2530,N_1516,N_1879);
nor U2531 (N_2531,N_1547,N_1983);
nor U2532 (N_2532,N_2219,N_1287);
nand U2533 (N_2533,N_2128,N_2464);
nor U2534 (N_2534,N_1825,N_2072);
nor U2535 (N_2535,N_2412,N_1645);
or U2536 (N_2536,N_2416,N_2272);
xnor U2537 (N_2537,N_1611,N_1586);
nor U2538 (N_2538,N_1253,N_1409);
nor U2539 (N_2539,N_1953,N_1998);
nor U2540 (N_2540,N_1670,N_2064);
nor U2541 (N_2541,N_2105,N_1770);
or U2542 (N_2542,N_1596,N_1837);
xor U2543 (N_2543,N_1333,N_2264);
and U2544 (N_2544,N_1593,N_2042);
nor U2545 (N_2545,N_1861,N_2135);
nand U2546 (N_2546,N_1634,N_2154);
nand U2547 (N_2547,N_2451,N_1389);
nand U2548 (N_2548,N_2241,N_2073);
nand U2549 (N_2549,N_1814,N_2303);
nand U2550 (N_2550,N_1548,N_2201);
and U2551 (N_2551,N_1937,N_2496);
nor U2552 (N_2552,N_1396,N_1930);
nor U2553 (N_2553,N_2395,N_2003);
xnor U2554 (N_2554,N_1328,N_2359);
nand U2555 (N_2555,N_2028,N_1813);
or U2556 (N_2556,N_1621,N_2292);
nand U2557 (N_2557,N_2127,N_1276);
nand U2558 (N_2558,N_1443,N_2239);
nor U2559 (N_2559,N_2065,N_2353);
nor U2560 (N_2560,N_1405,N_2188);
or U2561 (N_2561,N_1291,N_1599);
and U2562 (N_2562,N_1465,N_2210);
nand U2563 (N_2563,N_2483,N_1817);
nor U2564 (N_2564,N_2415,N_1591);
or U2565 (N_2565,N_1622,N_1284);
and U2566 (N_2566,N_1426,N_1851);
nand U2567 (N_2567,N_1890,N_1636);
nand U2568 (N_2568,N_1880,N_2302);
xnor U2569 (N_2569,N_2269,N_2138);
nor U2570 (N_2570,N_1564,N_2224);
nor U2571 (N_2571,N_2401,N_1934);
and U2572 (N_2572,N_2211,N_2041);
nand U2573 (N_2573,N_2083,N_2455);
or U2574 (N_2574,N_1490,N_2295);
nand U2575 (N_2575,N_1600,N_1769);
nand U2576 (N_2576,N_2390,N_2254);
or U2577 (N_2577,N_1781,N_1463);
and U2578 (N_2578,N_2139,N_2251);
nand U2579 (N_2579,N_1805,N_1265);
and U2580 (N_2580,N_1592,N_1999);
or U2581 (N_2581,N_1705,N_1318);
or U2582 (N_2582,N_2191,N_1294);
nand U2583 (N_2583,N_1910,N_1456);
xor U2584 (N_2584,N_2119,N_1860);
xor U2585 (N_2585,N_1300,N_2212);
and U2586 (N_2586,N_2310,N_1563);
nor U2587 (N_2587,N_2313,N_2015);
or U2588 (N_2588,N_2148,N_2163);
and U2589 (N_2589,N_1662,N_1888);
nand U2590 (N_2590,N_2037,N_2085);
nand U2591 (N_2591,N_1718,N_1572);
nor U2592 (N_2592,N_1703,N_1617);
nand U2593 (N_2593,N_2067,N_1602);
nand U2594 (N_2594,N_1909,N_1804);
nor U2595 (N_2595,N_2459,N_1767);
or U2596 (N_2596,N_2079,N_1285);
nor U2597 (N_2597,N_2082,N_1609);
xnor U2598 (N_2598,N_2081,N_1530);
xnor U2599 (N_2599,N_2132,N_1919);
xor U2600 (N_2600,N_1315,N_1690);
nor U2601 (N_2601,N_1714,N_2477);
or U2602 (N_2602,N_2236,N_2144);
and U2603 (N_2603,N_1819,N_1469);
nand U2604 (N_2604,N_1368,N_1709);
or U2605 (N_2605,N_2018,N_1853);
xnor U2606 (N_2606,N_1848,N_1971);
nor U2607 (N_2607,N_1689,N_1373);
and U2608 (N_2608,N_1730,N_1990);
nor U2609 (N_2609,N_2114,N_1873);
and U2610 (N_2610,N_1685,N_1768);
nand U2611 (N_2611,N_2192,N_2133);
and U2612 (N_2612,N_1657,N_2410);
nand U2613 (N_2613,N_2204,N_1965);
nor U2614 (N_2614,N_2424,N_1654);
and U2615 (N_2615,N_1411,N_1491);
nor U2616 (N_2616,N_2150,N_1963);
and U2617 (N_2617,N_1681,N_2411);
or U2618 (N_2618,N_1638,N_1740);
nand U2619 (N_2619,N_2123,N_2168);
or U2620 (N_2620,N_1394,N_1567);
nand U2621 (N_2621,N_2087,N_1736);
nand U2622 (N_2622,N_1920,N_1587);
nand U2623 (N_2623,N_2365,N_2033);
and U2624 (N_2624,N_2454,N_1450);
xnor U2625 (N_2625,N_2385,N_1708);
nor U2626 (N_2626,N_1459,N_1324);
or U2627 (N_2627,N_1721,N_2298);
nor U2628 (N_2628,N_1556,N_1453);
or U2629 (N_2629,N_2110,N_2088);
xnor U2630 (N_2630,N_1504,N_1541);
xor U2631 (N_2631,N_1342,N_2397);
or U2632 (N_2632,N_1260,N_2166);
nor U2633 (N_2633,N_2174,N_1264);
or U2634 (N_2634,N_1776,N_1785);
xor U2635 (N_2635,N_2420,N_1311);
nor U2636 (N_2636,N_1863,N_1964);
nor U2637 (N_2637,N_1488,N_1425);
or U2638 (N_2638,N_1508,N_2181);
and U2639 (N_2639,N_1925,N_1444);
and U2640 (N_2640,N_2382,N_1818);
xor U2641 (N_2641,N_2051,N_1330);
xnor U2642 (N_2642,N_1573,N_2318);
or U2643 (N_2643,N_1275,N_1782);
or U2644 (N_2644,N_1717,N_1928);
and U2645 (N_2645,N_2449,N_1506);
or U2646 (N_2646,N_1775,N_1641);
or U2647 (N_2647,N_2086,N_2271);
or U2648 (N_2648,N_1273,N_1620);
xor U2649 (N_2649,N_2267,N_2404);
xnor U2650 (N_2650,N_1500,N_1664);
and U2651 (N_2651,N_1496,N_2193);
or U2652 (N_2652,N_1337,N_1437);
and U2653 (N_2653,N_2336,N_2229);
and U2654 (N_2654,N_1571,N_2375);
and U2655 (N_2655,N_2498,N_1855);
or U2656 (N_2656,N_2268,N_2460);
and U2657 (N_2657,N_2333,N_1666);
xnor U2658 (N_2658,N_1949,N_1858);
or U2659 (N_2659,N_2326,N_1764);
nand U2660 (N_2660,N_1789,N_1754);
xor U2661 (N_2661,N_1310,N_1370);
nor U2662 (N_2662,N_2104,N_1939);
and U2663 (N_2663,N_2479,N_1955);
nor U2664 (N_2664,N_2060,N_2056);
nor U2665 (N_2665,N_1613,N_2417);
or U2666 (N_2666,N_2177,N_1250);
nor U2667 (N_2667,N_2124,N_2216);
or U2668 (N_2668,N_1974,N_1723);
xor U2669 (N_2669,N_2084,N_1724);
xnor U2670 (N_2670,N_2299,N_2031);
xor U2671 (N_2671,N_2422,N_2222);
nand U2672 (N_2672,N_2061,N_1435);
nand U2673 (N_2673,N_1369,N_1800);
or U2674 (N_2674,N_2368,N_1323);
nor U2675 (N_2675,N_2113,N_2473);
and U2676 (N_2676,N_2370,N_2226);
or U2677 (N_2677,N_2285,N_2349);
xor U2678 (N_2678,N_1277,N_2329);
nand U2679 (N_2679,N_1313,N_1604);
or U2680 (N_2680,N_2453,N_2439);
and U2681 (N_2681,N_1628,N_2355);
or U2682 (N_2682,N_2442,N_1663);
and U2683 (N_2683,N_1977,N_1757);
xnor U2684 (N_2684,N_1991,N_1297);
or U2685 (N_2685,N_2112,N_1912);
and U2686 (N_2686,N_2425,N_1468);
nand U2687 (N_2687,N_2499,N_2100);
nand U2688 (N_2688,N_1631,N_2036);
xnor U2689 (N_2689,N_2480,N_2161);
and U2690 (N_2690,N_2118,N_1319);
xor U2691 (N_2691,N_1797,N_1568);
xor U2692 (N_2692,N_1988,N_1283);
or U2693 (N_2693,N_2249,N_1554);
xnor U2694 (N_2694,N_1889,N_1845);
nor U2695 (N_2695,N_2461,N_1995);
or U2696 (N_2696,N_2392,N_1625);
and U2697 (N_2697,N_1694,N_1924);
xor U2698 (N_2698,N_1515,N_2402);
xor U2699 (N_2699,N_1915,N_1936);
or U2700 (N_2700,N_1780,N_1854);
xnor U2701 (N_2701,N_1551,N_2094);
nand U2702 (N_2702,N_2214,N_1446);
nand U2703 (N_2703,N_2441,N_1549);
nand U2704 (N_2704,N_1473,N_1966);
or U2705 (N_2705,N_2017,N_1993);
xnor U2706 (N_2706,N_2452,N_1552);
or U2707 (N_2707,N_1352,N_1533);
xor U2708 (N_2708,N_2472,N_2077);
nor U2709 (N_2709,N_1759,N_1864);
or U2710 (N_2710,N_2386,N_2430);
nand U2711 (N_2711,N_1832,N_2197);
or U2712 (N_2712,N_1826,N_2076);
or U2713 (N_2713,N_1887,N_1722);
nand U2714 (N_2714,N_1871,N_2450);
xor U2715 (N_2715,N_1668,N_2398);
and U2716 (N_2716,N_1471,N_1874);
and U2717 (N_2717,N_1379,N_1716);
xor U2718 (N_2718,N_1735,N_2075);
nor U2719 (N_2719,N_1314,N_1345);
nor U2720 (N_2720,N_1897,N_2317);
and U2721 (N_2721,N_1605,N_2080);
nand U2722 (N_2722,N_1293,N_1994);
nor U2723 (N_2723,N_2215,N_2045);
xnor U2724 (N_2724,N_2151,N_2413);
nand U2725 (N_2725,N_1558,N_2170);
xnor U2726 (N_2726,N_1702,N_1850);
and U2727 (N_2727,N_2182,N_1618);
nor U2728 (N_2728,N_1749,N_1470);
nor U2729 (N_2729,N_2301,N_2436);
nor U2730 (N_2730,N_2282,N_1510);
or U2731 (N_2731,N_1535,N_1292);
nand U2732 (N_2732,N_2002,N_2347);
xor U2733 (N_2733,N_1382,N_1286);
nand U2734 (N_2734,N_2246,N_1707);
xnor U2735 (N_2735,N_1808,N_2374);
or U2736 (N_2736,N_2059,N_2158);
and U2737 (N_2737,N_1566,N_1951);
xor U2738 (N_2738,N_1699,N_2230);
nor U2739 (N_2739,N_1859,N_2209);
nand U2740 (N_2740,N_1553,N_1891);
or U2741 (N_2741,N_1540,N_1978);
or U2742 (N_2742,N_1691,N_1720);
nor U2743 (N_2743,N_1262,N_1531);
xnor U2744 (N_2744,N_2021,N_2261);
nand U2745 (N_2745,N_1525,N_2419);
xnor U2746 (N_2746,N_1255,N_1779);
and U2747 (N_2747,N_1502,N_2155);
nor U2748 (N_2748,N_2095,N_2263);
xnor U2749 (N_2749,N_2372,N_1725);
or U2750 (N_2750,N_1546,N_1357);
nand U2751 (N_2751,N_1651,N_2495);
nand U2752 (N_2752,N_1539,N_1436);
and U2753 (N_2753,N_2055,N_2101);
nor U2754 (N_2754,N_2006,N_1472);
nor U2755 (N_2755,N_1270,N_1958);
and U2756 (N_2756,N_1499,N_2312);
nor U2757 (N_2757,N_2160,N_2225);
nand U2758 (N_2758,N_2068,N_2125);
xor U2759 (N_2759,N_1304,N_2043);
nand U2760 (N_2760,N_1267,N_2165);
nor U2761 (N_2761,N_1895,N_1671);
nor U2762 (N_2762,N_1334,N_1843);
and U2763 (N_2763,N_2297,N_1918);
and U2764 (N_2764,N_1712,N_2327);
or U2765 (N_2765,N_1557,N_1884);
nor U2766 (N_2766,N_2046,N_2432);
or U2767 (N_2767,N_1834,N_1584);
xor U2768 (N_2768,N_2324,N_1777);
nor U2769 (N_2769,N_1518,N_1698);
and U2770 (N_2770,N_2357,N_1271);
nor U2771 (N_2771,N_1649,N_1594);
and U2772 (N_2772,N_1343,N_2278);
and U2773 (N_2773,N_1807,N_2143);
xnor U2774 (N_2774,N_2322,N_2362);
and U2775 (N_2775,N_1281,N_1512);
xor U2776 (N_2776,N_1774,N_1646);
nor U2777 (N_2777,N_1896,N_2265);
xnor U2778 (N_2778,N_1660,N_2438);
and U2779 (N_2779,N_2283,N_2202);
nor U2780 (N_2780,N_1428,N_2408);
and U2781 (N_2781,N_2305,N_1756);
and U2782 (N_2782,N_1655,N_1387);
nand U2783 (N_2783,N_2050,N_1968);
nor U2784 (N_2784,N_1827,N_2234);
and U2785 (N_2785,N_2279,N_2240);
xor U2786 (N_2786,N_1947,N_2024);
and U2787 (N_2787,N_2007,N_1931);
and U2788 (N_2788,N_2338,N_2315);
nor U2789 (N_2789,N_1447,N_2435);
nor U2790 (N_2790,N_1981,N_1967);
or U2791 (N_2791,N_1360,N_1984);
xor U2792 (N_2792,N_2360,N_1745);
xor U2793 (N_2793,N_1695,N_2069);
nor U2794 (N_2794,N_2487,N_1823);
nor U2795 (N_2795,N_1667,N_1833);
xor U2796 (N_2796,N_1375,N_1569);
xor U2797 (N_2797,N_2159,N_2106);
nand U2798 (N_2798,N_2290,N_2103);
xnor U2799 (N_2799,N_2169,N_2199);
nand U2800 (N_2800,N_2273,N_1710);
or U2801 (N_2801,N_1578,N_1847);
nand U2802 (N_2802,N_1820,N_2328);
or U2803 (N_2803,N_1846,N_1344);
nand U2804 (N_2804,N_1413,N_1384);
xor U2805 (N_2805,N_2205,N_1257);
or U2806 (N_2806,N_1742,N_1766);
nand U2807 (N_2807,N_1575,N_2493);
or U2808 (N_2808,N_2281,N_1259);
nand U2809 (N_2809,N_2257,N_1643);
or U2810 (N_2810,N_1430,N_2213);
and U2811 (N_2811,N_1686,N_1454);
xnor U2812 (N_2812,N_1434,N_2004);
and U2813 (N_2813,N_2462,N_1422);
nor U2814 (N_2814,N_1585,N_1869);
nand U2815 (N_2815,N_1538,N_1418);
xnor U2816 (N_2816,N_1632,N_2146);
nor U2817 (N_2817,N_1616,N_1467);
and U2818 (N_2818,N_2049,N_2418);
nor U2819 (N_2819,N_1479,N_1753);
and U2820 (N_2820,N_1475,N_2470);
and U2821 (N_2821,N_2012,N_1728);
and U2822 (N_2822,N_1905,N_1788);
and U2823 (N_2823,N_1950,N_2389);
nor U2824 (N_2824,N_2198,N_1340);
xor U2825 (N_2825,N_1365,N_1731);
nand U2826 (N_2826,N_1582,N_1526);
xnor U2827 (N_2827,N_1316,N_1865);
or U2828 (N_2828,N_1341,N_1639);
nor U2829 (N_2829,N_2250,N_2027);
or U2830 (N_2830,N_2228,N_2008);
nand U2831 (N_2831,N_1700,N_1610);
nand U2832 (N_2832,N_1336,N_1580);
and U2833 (N_2833,N_2129,N_1378);
xor U2834 (N_2834,N_1856,N_2016);
and U2835 (N_2835,N_2307,N_2189);
or U2836 (N_2836,N_1917,N_2152);
or U2837 (N_2837,N_1524,N_2366);
nand U2838 (N_2838,N_1948,N_1926);
xor U2839 (N_2839,N_1793,N_2026);
nor U2840 (N_2840,N_1997,N_2147);
or U2841 (N_2841,N_1282,N_1417);
xor U2842 (N_2842,N_2323,N_1732);
nand U2843 (N_2843,N_1256,N_2238);
nor U2844 (N_2844,N_1902,N_2405);
xor U2845 (N_2845,N_2164,N_1626);
xor U2846 (N_2846,N_1483,N_1892);
xor U2847 (N_2847,N_1838,N_1288);
nand U2848 (N_2848,N_2369,N_1258);
nor U2849 (N_2849,N_1806,N_1400);
or U2850 (N_2850,N_2262,N_2437);
or U2851 (N_2851,N_1272,N_2245);
and U2852 (N_2852,N_1519,N_1816);
nor U2853 (N_2853,N_2218,N_1633);
nand U2854 (N_2854,N_2394,N_2497);
nand U2855 (N_2855,N_2485,N_1460);
xnor U2856 (N_2856,N_1386,N_1706);
or U2857 (N_2857,N_1493,N_1916);
nor U2858 (N_2858,N_2337,N_2288);
and U2859 (N_2859,N_2195,N_1362);
or U2860 (N_2860,N_1762,N_1822);
nand U2861 (N_2861,N_1486,N_2090);
nor U2862 (N_2862,N_1385,N_1404);
xnor U2863 (N_2863,N_1354,N_1642);
and U2864 (N_2864,N_1652,N_1726);
nand U2865 (N_2865,N_1261,N_2171);
nand U2866 (N_2866,N_2116,N_2185);
xor U2867 (N_2867,N_1831,N_1590);
nand U2868 (N_2868,N_2458,N_1363);
and U2869 (N_2869,N_2421,N_1903);
and U2870 (N_2870,N_1299,N_1883);
or U2871 (N_2871,N_2490,N_1899);
nor U2872 (N_2872,N_1906,N_2178);
xnor U2873 (N_2873,N_1747,N_1701);
nor U2874 (N_2874,N_2341,N_1715);
or U2875 (N_2875,N_2260,N_1836);
xor U2876 (N_2876,N_2289,N_1688);
xnor U2877 (N_2877,N_2053,N_1427);
xor U2878 (N_2878,N_2280,N_2443);
xnor U2879 (N_2879,N_1598,N_1957);
or U2880 (N_2880,N_2448,N_2126);
and U2881 (N_2881,N_1364,N_2221);
or U2882 (N_2882,N_2275,N_1885);
and U2883 (N_2883,N_1614,N_1629);
nand U2884 (N_2884,N_1380,N_2484);
or U2885 (N_2885,N_2423,N_1509);
xor U2886 (N_2886,N_2071,N_1280);
and U2887 (N_2887,N_1876,N_1251);
or U2888 (N_2888,N_1743,N_1680);
nor U2889 (N_2889,N_1637,N_1829);
and U2890 (N_2890,N_2057,N_1875);
nand U2891 (N_2891,N_1796,N_1624);
nor U2892 (N_2892,N_1741,N_1461);
or U2893 (N_2893,N_2089,N_1729);
nand U2894 (N_2894,N_1589,N_1570);
nor U2895 (N_2895,N_1329,N_1810);
and U2896 (N_2896,N_1347,N_1412);
or U2897 (N_2897,N_1606,N_1466);
nand U2898 (N_2898,N_1441,N_1901);
and U2899 (N_2899,N_2208,N_1755);
nor U2900 (N_2900,N_1301,N_1923);
nand U2901 (N_2901,N_1765,N_1451);
nand U2902 (N_2902,N_2078,N_2384);
and U2903 (N_2903,N_2287,N_1339);
nor U2904 (N_2904,N_1799,N_2332);
and U2905 (N_2905,N_2364,N_1317);
or U2906 (N_2906,N_2381,N_1403);
or U2907 (N_2907,N_2032,N_2463);
or U2908 (N_2908,N_1306,N_1674);
xor U2909 (N_2909,N_2120,N_1433);
and U2910 (N_2910,N_1361,N_1429);
nand U2911 (N_2911,N_1448,N_2237);
nand U2912 (N_2912,N_2340,N_1693);
nor U2913 (N_2913,N_2005,N_2200);
nand U2914 (N_2914,N_2232,N_1619);
or U2915 (N_2915,N_1868,N_2176);
nor U2916 (N_2916,N_2346,N_2184);
and U2917 (N_2917,N_1484,N_1577);
and U2918 (N_2918,N_2039,N_1894);
xnor U2919 (N_2919,N_1511,N_2010);
xor U2920 (N_2920,N_1733,N_2391);
nand U2921 (N_2921,N_1536,N_2259);
or U2922 (N_2922,N_1326,N_1439);
or U2923 (N_2923,N_1579,N_1677);
and U2924 (N_2924,N_2304,N_1772);
and U2925 (N_2925,N_1778,N_1355);
xor U2926 (N_2926,N_2321,N_1935);
nor U2927 (N_2927,N_2367,N_1274);
or U2928 (N_2928,N_1615,N_2035);
nor U2929 (N_2929,N_1737,N_1996);
and U2930 (N_2930,N_1630,N_1278);
xnor U2931 (N_2931,N_1532,N_1665);
nor U2932 (N_2932,N_1588,N_2023);
or U2933 (N_2933,N_1410,N_1878);
nor U2934 (N_2934,N_1907,N_1440);
xor U2935 (N_2935,N_1492,N_1980);
or U2936 (N_2936,N_2465,N_1644);
or U2937 (N_2937,N_2092,N_1943);
nor U2938 (N_2938,N_2247,N_1932);
nand U2939 (N_2939,N_1401,N_1559);
and U2940 (N_2940,N_1445,N_2097);
nor U2941 (N_2941,N_1481,N_1452);
xor U2942 (N_2942,N_1684,N_2489);
nor U2943 (N_2943,N_2406,N_1938);
and U2944 (N_2944,N_2203,N_1397);
and U2945 (N_2945,N_2187,N_1852);
xnor U2946 (N_2946,N_2047,N_2248);
xnor U2947 (N_2947,N_1945,N_2383);
nor U2948 (N_2948,N_1358,N_1839);
and U2949 (N_2949,N_1522,N_1719);
or U2950 (N_2950,N_2022,N_1798);
nand U2951 (N_2951,N_1713,N_2063);
or U2952 (N_2952,N_1659,N_2258);
or U2953 (N_2953,N_1480,N_1673);
or U2954 (N_2954,N_2207,N_2136);
nor U2955 (N_2955,N_1841,N_2109);
and U2956 (N_2956,N_2172,N_1607);
and U2957 (N_2957,N_1809,N_1987);
xnor U2958 (N_2958,N_2320,N_1302);
nor U2959 (N_2959,N_1758,N_1371);
nor U2960 (N_2960,N_2034,N_2093);
or U2961 (N_2961,N_1882,N_1744);
nand U2962 (N_2962,N_2481,N_2000);
and U2963 (N_2963,N_1482,N_1457);
and U2964 (N_2964,N_2345,N_2380);
nand U2965 (N_2965,N_2070,N_2276);
xor U2966 (N_2966,N_1402,N_1309);
and U2967 (N_2967,N_1565,N_2186);
or U2968 (N_2968,N_1786,N_2014);
or U2969 (N_2969,N_1252,N_2117);
and U2970 (N_2970,N_2311,N_2378);
nand U2971 (N_2971,N_2266,N_1458);
or U2972 (N_2972,N_1908,N_2431);
xnor U2973 (N_2973,N_1738,N_1367);
nor U2974 (N_2974,N_1346,N_2013);
and U2975 (N_2975,N_1954,N_1419);
nand U2976 (N_2976,N_1623,N_2447);
or U2977 (N_2977,N_1911,N_1922);
nand U2978 (N_2978,N_2040,N_2217);
nor U2979 (N_2979,N_1543,N_1672);
or U2980 (N_2980,N_2474,N_1989);
nand U2981 (N_2981,N_2457,N_1811);
or U2982 (N_2982,N_2102,N_2244);
nand U2983 (N_2983,N_1979,N_2393);
and U2984 (N_2984,N_2471,N_2325);
nand U2985 (N_2985,N_1290,N_1842);
or U2986 (N_2986,N_1696,N_1682);
and U2987 (N_2987,N_2330,N_2294);
nand U2988 (N_2988,N_2149,N_1656);
xor U2989 (N_2989,N_2130,N_1790);
xor U2990 (N_2990,N_1514,N_1462);
and U2991 (N_2991,N_1534,N_2194);
nor U2992 (N_2992,N_2253,N_2400);
xnor U2993 (N_2993,N_2140,N_2494);
nor U2994 (N_2994,N_2426,N_1877);
nand U2995 (N_2995,N_1455,N_1432);
nor U2996 (N_2996,N_1835,N_2363);
or U2997 (N_2997,N_1322,N_2153);
nand U2998 (N_2998,N_2488,N_2052);
nor U2999 (N_2999,N_1263,N_2162);
or U3000 (N_3000,N_1298,N_1986);
and U3001 (N_3001,N_1348,N_1350);
xor U3002 (N_3002,N_1771,N_1376);
or U3003 (N_3003,N_1544,N_2316);
xnor U3004 (N_3004,N_1658,N_2227);
nand U3005 (N_3005,N_1353,N_1576);
or U3006 (N_3006,N_1438,N_1487);
and U3007 (N_3007,N_1269,N_1562);
xor U3008 (N_3008,N_1431,N_1295);
nand U3009 (N_3009,N_1687,N_1849);
xnor U3010 (N_3010,N_2339,N_2456);
and U3011 (N_3011,N_2350,N_2309);
nand U3012 (N_3012,N_1254,N_1442);
xor U3013 (N_3013,N_1784,N_1550);
or U3014 (N_3014,N_1648,N_1595);
or U3015 (N_3015,N_2134,N_1727);
or U3016 (N_3016,N_1946,N_1704);
nor U3017 (N_3017,N_1927,N_2196);
or U3018 (N_3018,N_2344,N_1399);
xor U3019 (N_3019,N_1830,N_2038);
and U3020 (N_3020,N_1794,N_2142);
nor U3021 (N_3021,N_1763,N_1961);
nor U3022 (N_3022,N_2029,N_2296);
nor U3023 (N_3023,N_1359,N_2107);
or U3024 (N_3024,N_1970,N_1612);
nor U3025 (N_3025,N_1640,N_1351);
nand U3026 (N_3026,N_1982,N_1750);
xor U3027 (N_3027,N_2145,N_2231);
and U3028 (N_3028,N_2066,N_2414);
xor U3029 (N_3029,N_1321,N_1392);
and U3030 (N_3030,N_2121,N_2019);
nor U3031 (N_3031,N_1601,N_1635);
nand U3032 (N_3032,N_2096,N_2491);
nor U3033 (N_3033,N_1692,N_2183);
nor U3034 (N_3034,N_2314,N_1268);
nor U3035 (N_3035,N_1408,N_1390);
nor U3036 (N_3036,N_1307,N_1647);
and U3037 (N_3037,N_2445,N_2440);
nand U3038 (N_3038,N_2099,N_1338);
nor U3039 (N_3039,N_1372,N_2190);
nand U3040 (N_3040,N_2270,N_2115);
nand U3041 (N_3041,N_2433,N_1801);
nand U3042 (N_3042,N_1941,N_1795);
xor U3043 (N_3043,N_1900,N_2358);
and U3044 (N_3044,N_1679,N_1752);
and U3045 (N_3045,N_1944,N_1476);
or U3046 (N_3046,N_1904,N_1303);
xnor U3047 (N_3047,N_2011,N_1335);
nand U3048 (N_3048,N_1952,N_2466);
xnor U3049 (N_3049,N_1678,N_2361);
and U3050 (N_3050,N_2048,N_1783);
nand U3051 (N_3051,N_1675,N_1898);
and U3052 (N_3052,N_1962,N_1872);
nor U3053 (N_3053,N_1529,N_1734);
or U3054 (N_3054,N_2387,N_1560);
nor U3055 (N_3055,N_1992,N_1527);
nand U3056 (N_3056,N_1542,N_2098);
xor U3057 (N_3057,N_2478,N_1398);
nand U3058 (N_3058,N_2030,N_1266);
nand U3059 (N_3059,N_1921,N_1870);
xnor U3060 (N_3060,N_1697,N_1803);
nor U3061 (N_3061,N_1913,N_2141);
or U3062 (N_3062,N_2379,N_2062);
nor U3063 (N_3063,N_1423,N_2319);
or U3064 (N_3064,N_1388,N_2492);
or U3065 (N_3065,N_1296,N_1424);
nor U3066 (N_3066,N_2252,N_1597);
and U3067 (N_3067,N_1574,N_2157);
and U3068 (N_3068,N_2255,N_2131);
xor U3069 (N_3069,N_1650,N_1653);
nor U3070 (N_3070,N_1327,N_2482);
nor U3071 (N_3071,N_2074,N_2409);
xor U3072 (N_3072,N_2306,N_1498);
nand U3073 (N_3073,N_1933,N_1676);
xnor U3074 (N_3074,N_1748,N_2274);
and U3075 (N_3075,N_2467,N_1608);
nor U3076 (N_3076,N_1381,N_2434);
or U3077 (N_3077,N_2054,N_1505);
nand U3078 (N_3078,N_1940,N_1956);
and U3079 (N_3079,N_1867,N_2206);
nand U3080 (N_3080,N_1289,N_2308);
xnor U3081 (N_3081,N_1497,N_1325);
nand U3082 (N_3082,N_1960,N_2180);
or U3083 (N_3083,N_1501,N_2025);
nor U3084 (N_3084,N_1815,N_2348);
xnor U3085 (N_3085,N_1449,N_1383);
and U3086 (N_3086,N_2476,N_2009);
xor U3087 (N_3087,N_1929,N_2475);
and U3088 (N_3088,N_1969,N_1603);
nand U3089 (N_3089,N_1377,N_1521);
nand U3090 (N_3090,N_1791,N_1821);
and U3091 (N_3091,N_1312,N_1985);
nand U3092 (N_3092,N_1840,N_1416);
and U3093 (N_3093,N_1421,N_2167);
or U3094 (N_3094,N_1555,N_2242);
xnor U3095 (N_3095,N_2388,N_1374);
and U3096 (N_3096,N_2256,N_1844);
xnor U3097 (N_3097,N_2334,N_1420);
or U3098 (N_3098,N_2377,N_2407);
xnor U3099 (N_3099,N_2403,N_1881);
or U3100 (N_3100,N_1478,N_2020);
nor U3101 (N_3101,N_2331,N_2428);
nand U3102 (N_3102,N_1331,N_2291);
nor U3103 (N_3103,N_1751,N_1520);
nor U3104 (N_3104,N_1581,N_2335);
nor U3105 (N_3105,N_2352,N_2429);
and U3106 (N_3106,N_1824,N_1627);
xnor U3107 (N_3107,N_1528,N_1513);
nor U3108 (N_3108,N_1279,N_1802);
and U3109 (N_3109,N_1761,N_1477);
nor U3110 (N_3110,N_2342,N_2444);
and U3111 (N_3111,N_2373,N_2300);
and U3112 (N_3112,N_1391,N_1485);
nand U3113 (N_3113,N_1474,N_2233);
nand U3114 (N_3114,N_2284,N_1561);
nor U3115 (N_3115,N_1976,N_1812);
nor U3116 (N_3116,N_1464,N_1366);
nand U3117 (N_3117,N_1683,N_1308);
nand U3118 (N_3118,N_2220,N_1828);
nand U3119 (N_3119,N_2354,N_2351);
or U3120 (N_3120,N_2223,N_2044);
nand U3121 (N_3121,N_1305,N_1494);
nor U3122 (N_3122,N_2446,N_1975);
or U3123 (N_3123,N_1857,N_2293);
xnor U3124 (N_3124,N_1661,N_2356);
and U3125 (N_3125,N_1553,N_1713);
or U3126 (N_3126,N_1470,N_1476);
or U3127 (N_3127,N_2459,N_2480);
and U3128 (N_3128,N_2424,N_1543);
nand U3129 (N_3129,N_1715,N_2021);
nand U3130 (N_3130,N_1439,N_1309);
nor U3131 (N_3131,N_1737,N_2437);
nor U3132 (N_3132,N_2123,N_1958);
nor U3133 (N_3133,N_2044,N_2329);
or U3134 (N_3134,N_1557,N_2465);
nand U3135 (N_3135,N_1595,N_1724);
nor U3136 (N_3136,N_2201,N_2425);
xnor U3137 (N_3137,N_1718,N_2331);
nor U3138 (N_3138,N_1918,N_1308);
nor U3139 (N_3139,N_1503,N_2495);
or U3140 (N_3140,N_1971,N_1600);
and U3141 (N_3141,N_2385,N_1462);
nand U3142 (N_3142,N_1583,N_2185);
nand U3143 (N_3143,N_2456,N_1896);
or U3144 (N_3144,N_1476,N_1932);
or U3145 (N_3145,N_1699,N_1743);
or U3146 (N_3146,N_1675,N_2152);
xor U3147 (N_3147,N_1504,N_1850);
and U3148 (N_3148,N_2494,N_1587);
xor U3149 (N_3149,N_2422,N_2457);
and U3150 (N_3150,N_1784,N_1282);
nor U3151 (N_3151,N_2114,N_2111);
and U3152 (N_3152,N_1405,N_1813);
nor U3153 (N_3153,N_2452,N_1292);
or U3154 (N_3154,N_1682,N_2006);
xor U3155 (N_3155,N_2372,N_1356);
and U3156 (N_3156,N_2378,N_2054);
and U3157 (N_3157,N_2375,N_1917);
or U3158 (N_3158,N_1672,N_1929);
and U3159 (N_3159,N_1681,N_1686);
and U3160 (N_3160,N_1432,N_1481);
and U3161 (N_3161,N_2318,N_2178);
and U3162 (N_3162,N_1800,N_2470);
or U3163 (N_3163,N_1748,N_1783);
nand U3164 (N_3164,N_1360,N_1849);
or U3165 (N_3165,N_1685,N_1818);
nand U3166 (N_3166,N_1454,N_1424);
xnor U3167 (N_3167,N_1410,N_1650);
nand U3168 (N_3168,N_1452,N_1829);
nor U3169 (N_3169,N_1452,N_2103);
nand U3170 (N_3170,N_2420,N_1872);
xor U3171 (N_3171,N_1931,N_2129);
xor U3172 (N_3172,N_2464,N_1532);
nand U3173 (N_3173,N_1477,N_1528);
nor U3174 (N_3174,N_1874,N_1337);
and U3175 (N_3175,N_2170,N_1914);
nand U3176 (N_3176,N_2064,N_1657);
nor U3177 (N_3177,N_1547,N_1445);
nand U3178 (N_3178,N_2141,N_2135);
nor U3179 (N_3179,N_1658,N_1518);
or U3180 (N_3180,N_2255,N_1458);
xor U3181 (N_3181,N_1874,N_2422);
xor U3182 (N_3182,N_2152,N_1373);
xnor U3183 (N_3183,N_1660,N_1934);
xnor U3184 (N_3184,N_1582,N_1498);
or U3185 (N_3185,N_1647,N_1375);
nor U3186 (N_3186,N_1577,N_1662);
nor U3187 (N_3187,N_1340,N_2440);
or U3188 (N_3188,N_2000,N_1464);
or U3189 (N_3189,N_1375,N_1513);
or U3190 (N_3190,N_1716,N_1435);
xor U3191 (N_3191,N_1660,N_1778);
and U3192 (N_3192,N_2000,N_2178);
nor U3193 (N_3193,N_1635,N_2425);
xnor U3194 (N_3194,N_1758,N_1888);
nand U3195 (N_3195,N_2224,N_2283);
or U3196 (N_3196,N_2443,N_2233);
nor U3197 (N_3197,N_1597,N_2442);
or U3198 (N_3198,N_1633,N_1582);
or U3199 (N_3199,N_1661,N_2176);
xor U3200 (N_3200,N_2018,N_1935);
and U3201 (N_3201,N_2326,N_2087);
and U3202 (N_3202,N_1557,N_1624);
and U3203 (N_3203,N_2270,N_2147);
nor U3204 (N_3204,N_2216,N_2099);
nor U3205 (N_3205,N_1407,N_2219);
or U3206 (N_3206,N_1371,N_1816);
or U3207 (N_3207,N_2488,N_1468);
nand U3208 (N_3208,N_1445,N_1250);
and U3209 (N_3209,N_1570,N_1961);
nor U3210 (N_3210,N_2423,N_2164);
and U3211 (N_3211,N_1561,N_2041);
xor U3212 (N_3212,N_2410,N_1490);
nand U3213 (N_3213,N_1658,N_1477);
and U3214 (N_3214,N_1973,N_2126);
nor U3215 (N_3215,N_2177,N_2489);
and U3216 (N_3216,N_2127,N_1764);
nor U3217 (N_3217,N_1380,N_2485);
nor U3218 (N_3218,N_2440,N_1897);
xor U3219 (N_3219,N_1459,N_1516);
xnor U3220 (N_3220,N_1332,N_1303);
and U3221 (N_3221,N_1954,N_1747);
or U3222 (N_3222,N_1645,N_2317);
or U3223 (N_3223,N_1678,N_1771);
and U3224 (N_3224,N_2126,N_1338);
nor U3225 (N_3225,N_2392,N_2228);
or U3226 (N_3226,N_1385,N_2204);
xor U3227 (N_3227,N_1273,N_2310);
xor U3228 (N_3228,N_2439,N_2458);
xnor U3229 (N_3229,N_1320,N_1723);
xnor U3230 (N_3230,N_1742,N_1497);
and U3231 (N_3231,N_2107,N_1278);
nand U3232 (N_3232,N_1449,N_2069);
nor U3233 (N_3233,N_1747,N_2078);
or U3234 (N_3234,N_1980,N_1965);
nor U3235 (N_3235,N_1738,N_1975);
and U3236 (N_3236,N_1497,N_2164);
xnor U3237 (N_3237,N_2063,N_1522);
xnor U3238 (N_3238,N_2110,N_1797);
and U3239 (N_3239,N_2089,N_2186);
and U3240 (N_3240,N_2407,N_1871);
nand U3241 (N_3241,N_1838,N_2063);
xnor U3242 (N_3242,N_1747,N_2077);
nand U3243 (N_3243,N_2145,N_1375);
or U3244 (N_3244,N_1854,N_2402);
and U3245 (N_3245,N_1946,N_1730);
nor U3246 (N_3246,N_2085,N_2373);
nand U3247 (N_3247,N_1595,N_1422);
nand U3248 (N_3248,N_2061,N_1732);
xnor U3249 (N_3249,N_1626,N_1716);
xnor U3250 (N_3250,N_2266,N_2351);
nor U3251 (N_3251,N_1484,N_2163);
and U3252 (N_3252,N_1752,N_1629);
nand U3253 (N_3253,N_1839,N_1902);
xor U3254 (N_3254,N_2128,N_1751);
xor U3255 (N_3255,N_1673,N_1503);
xor U3256 (N_3256,N_1294,N_2168);
nor U3257 (N_3257,N_1454,N_1483);
and U3258 (N_3258,N_2171,N_1639);
and U3259 (N_3259,N_2206,N_2041);
nor U3260 (N_3260,N_2402,N_2275);
or U3261 (N_3261,N_2105,N_1480);
nand U3262 (N_3262,N_2347,N_2049);
xnor U3263 (N_3263,N_2218,N_1769);
and U3264 (N_3264,N_1587,N_1390);
or U3265 (N_3265,N_2379,N_1270);
or U3266 (N_3266,N_1846,N_1594);
nor U3267 (N_3267,N_2492,N_1891);
and U3268 (N_3268,N_1629,N_2261);
nor U3269 (N_3269,N_1459,N_2431);
and U3270 (N_3270,N_2279,N_2032);
or U3271 (N_3271,N_1351,N_1362);
nor U3272 (N_3272,N_2441,N_2230);
nor U3273 (N_3273,N_1366,N_2434);
xnor U3274 (N_3274,N_2376,N_1535);
xnor U3275 (N_3275,N_1645,N_1390);
xor U3276 (N_3276,N_1398,N_2437);
and U3277 (N_3277,N_1587,N_1671);
and U3278 (N_3278,N_1402,N_2242);
and U3279 (N_3279,N_2251,N_2095);
nand U3280 (N_3280,N_1822,N_1518);
nor U3281 (N_3281,N_1501,N_2485);
nand U3282 (N_3282,N_2144,N_2175);
and U3283 (N_3283,N_2371,N_1718);
and U3284 (N_3284,N_2473,N_1275);
nand U3285 (N_3285,N_1527,N_2492);
nor U3286 (N_3286,N_1845,N_1522);
nor U3287 (N_3287,N_1943,N_1381);
or U3288 (N_3288,N_1754,N_1532);
and U3289 (N_3289,N_2187,N_1681);
nand U3290 (N_3290,N_2480,N_2460);
and U3291 (N_3291,N_1723,N_1861);
nand U3292 (N_3292,N_1644,N_2365);
or U3293 (N_3293,N_2349,N_1937);
xor U3294 (N_3294,N_1939,N_2263);
and U3295 (N_3295,N_2315,N_2268);
and U3296 (N_3296,N_2018,N_2351);
nor U3297 (N_3297,N_2382,N_2324);
and U3298 (N_3298,N_1878,N_1456);
and U3299 (N_3299,N_2310,N_1564);
and U3300 (N_3300,N_2028,N_1491);
nand U3301 (N_3301,N_1384,N_1735);
nand U3302 (N_3302,N_1450,N_2016);
xor U3303 (N_3303,N_1900,N_2076);
xor U3304 (N_3304,N_1732,N_2056);
nor U3305 (N_3305,N_1713,N_1352);
nand U3306 (N_3306,N_1716,N_1794);
nor U3307 (N_3307,N_1562,N_2466);
and U3308 (N_3308,N_2354,N_2310);
nand U3309 (N_3309,N_2335,N_1358);
nand U3310 (N_3310,N_1391,N_2278);
xor U3311 (N_3311,N_1254,N_2460);
or U3312 (N_3312,N_1781,N_1895);
nor U3313 (N_3313,N_2444,N_1755);
or U3314 (N_3314,N_2393,N_1850);
or U3315 (N_3315,N_2231,N_2235);
and U3316 (N_3316,N_1950,N_2184);
nor U3317 (N_3317,N_1323,N_2417);
and U3318 (N_3318,N_2287,N_2207);
and U3319 (N_3319,N_1922,N_1549);
xor U3320 (N_3320,N_1608,N_1324);
or U3321 (N_3321,N_2173,N_2351);
xor U3322 (N_3322,N_1387,N_2061);
nor U3323 (N_3323,N_1365,N_1369);
and U3324 (N_3324,N_2042,N_2120);
nor U3325 (N_3325,N_2181,N_2322);
nor U3326 (N_3326,N_2238,N_2347);
nand U3327 (N_3327,N_1717,N_2319);
nor U3328 (N_3328,N_2177,N_1281);
nor U3329 (N_3329,N_2276,N_1865);
nor U3330 (N_3330,N_2212,N_2463);
or U3331 (N_3331,N_1428,N_2277);
nor U3332 (N_3332,N_2023,N_1835);
and U3333 (N_3333,N_1740,N_1484);
and U3334 (N_3334,N_2244,N_1986);
nand U3335 (N_3335,N_2024,N_1797);
nand U3336 (N_3336,N_1376,N_1667);
nor U3337 (N_3337,N_1725,N_1626);
xor U3338 (N_3338,N_1431,N_1802);
nor U3339 (N_3339,N_1357,N_1562);
or U3340 (N_3340,N_1822,N_1890);
or U3341 (N_3341,N_1887,N_2022);
nor U3342 (N_3342,N_2258,N_1302);
nand U3343 (N_3343,N_1395,N_2135);
or U3344 (N_3344,N_2492,N_2284);
nor U3345 (N_3345,N_2475,N_1919);
nand U3346 (N_3346,N_2273,N_1702);
and U3347 (N_3347,N_1310,N_1449);
xor U3348 (N_3348,N_2480,N_2004);
nor U3349 (N_3349,N_1761,N_1844);
nor U3350 (N_3350,N_2355,N_1343);
nand U3351 (N_3351,N_2465,N_1348);
nor U3352 (N_3352,N_2025,N_1731);
and U3353 (N_3353,N_2351,N_2155);
xor U3354 (N_3354,N_1671,N_2495);
xor U3355 (N_3355,N_2098,N_1787);
and U3356 (N_3356,N_2133,N_2486);
and U3357 (N_3357,N_1907,N_1863);
and U3358 (N_3358,N_2323,N_2267);
and U3359 (N_3359,N_2038,N_2272);
nand U3360 (N_3360,N_2050,N_2448);
and U3361 (N_3361,N_2384,N_1558);
and U3362 (N_3362,N_1627,N_1386);
or U3363 (N_3363,N_1803,N_1755);
xor U3364 (N_3364,N_1887,N_2319);
or U3365 (N_3365,N_2408,N_1313);
nor U3366 (N_3366,N_1985,N_2319);
and U3367 (N_3367,N_2138,N_2268);
and U3368 (N_3368,N_1727,N_1273);
nand U3369 (N_3369,N_2105,N_2129);
and U3370 (N_3370,N_2222,N_2204);
or U3371 (N_3371,N_2301,N_1439);
xnor U3372 (N_3372,N_2057,N_1695);
and U3373 (N_3373,N_2170,N_1702);
or U3374 (N_3374,N_2484,N_1430);
xnor U3375 (N_3375,N_1441,N_2482);
xnor U3376 (N_3376,N_2324,N_1456);
and U3377 (N_3377,N_1856,N_2295);
nor U3378 (N_3378,N_1770,N_1871);
and U3379 (N_3379,N_1959,N_1930);
nand U3380 (N_3380,N_1779,N_2013);
and U3381 (N_3381,N_2022,N_2214);
or U3382 (N_3382,N_1276,N_2181);
nor U3383 (N_3383,N_1725,N_2320);
nor U3384 (N_3384,N_1764,N_1747);
and U3385 (N_3385,N_1312,N_1806);
xnor U3386 (N_3386,N_1507,N_1827);
nand U3387 (N_3387,N_1508,N_1315);
and U3388 (N_3388,N_1443,N_1561);
xnor U3389 (N_3389,N_2376,N_1832);
or U3390 (N_3390,N_1894,N_1354);
xnor U3391 (N_3391,N_1935,N_1793);
nand U3392 (N_3392,N_1672,N_2351);
nor U3393 (N_3393,N_2336,N_1684);
or U3394 (N_3394,N_1879,N_2054);
xor U3395 (N_3395,N_2146,N_1712);
or U3396 (N_3396,N_1750,N_2152);
or U3397 (N_3397,N_1911,N_1267);
xor U3398 (N_3398,N_2379,N_1801);
and U3399 (N_3399,N_2063,N_1916);
xnor U3400 (N_3400,N_1744,N_2385);
and U3401 (N_3401,N_2250,N_2331);
xnor U3402 (N_3402,N_1488,N_2320);
nor U3403 (N_3403,N_1816,N_1648);
and U3404 (N_3404,N_1339,N_2377);
or U3405 (N_3405,N_1396,N_1298);
nand U3406 (N_3406,N_1701,N_1666);
and U3407 (N_3407,N_2246,N_1963);
and U3408 (N_3408,N_2340,N_1680);
or U3409 (N_3409,N_1871,N_1573);
or U3410 (N_3410,N_2055,N_1796);
xnor U3411 (N_3411,N_1308,N_1276);
or U3412 (N_3412,N_1468,N_2170);
or U3413 (N_3413,N_2047,N_2384);
and U3414 (N_3414,N_2204,N_1605);
or U3415 (N_3415,N_2217,N_1374);
and U3416 (N_3416,N_1354,N_1838);
and U3417 (N_3417,N_2255,N_1715);
or U3418 (N_3418,N_1470,N_1265);
and U3419 (N_3419,N_1665,N_2003);
or U3420 (N_3420,N_2469,N_1941);
xor U3421 (N_3421,N_2351,N_2017);
xnor U3422 (N_3422,N_2402,N_2006);
xor U3423 (N_3423,N_2314,N_1780);
nor U3424 (N_3424,N_1508,N_1697);
nand U3425 (N_3425,N_2388,N_2042);
xnor U3426 (N_3426,N_2457,N_1718);
nand U3427 (N_3427,N_1922,N_2090);
xor U3428 (N_3428,N_1564,N_2382);
xor U3429 (N_3429,N_1922,N_1512);
nand U3430 (N_3430,N_2376,N_1658);
nor U3431 (N_3431,N_1301,N_1555);
and U3432 (N_3432,N_1937,N_1475);
xnor U3433 (N_3433,N_1667,N_1711);
nor U3434 (N_3434,N_1971,N_1619);
nor U3435 (N_3435,N_2284,N_1599);
nor U3436 (N_3436,N_2221,N_1290);
xnor U3437 (N_3437,N_1438,N_2332);
xnor U3438 (N_3438,N_1349,N_1973);
and U3439 (N_3439,N_2457,N_2385);
nand U3440 (N_3440,N_2119,N_1822);
nor U3441 (N_3441,N_1990,N_2239);
nor U3442 (N_3442,N_1935,N_1398);
and U3443 (N_3443,N_2335,N_1963);
nor U3444 (N_3444,N_1716,N_2244);
and U3445 (N_3445,N_2163,N_1647);
nand U3446 (N_3446,N_1974,N_2385);
nand U3447 (N_3447,N_1997,N_2433);
nor U3448 (N_3448,N_1301,N_1887);
and U3449 (N_3449,N_1763,N_1510);
and U3450 (N_3450,N_1822,N_2174);
xor U3451 (N_3451,N_1679,N_1847);
or U3452 (N_3452,N_1369,N_2201);
and U3453 (N_3453,N_2350,N_2123);
or U3454 (N_3454,N_2211,N_1846);
and U3455 (N_3455,N_1538,N_2053);
nor U3456 (N_3456,N_1408,N_1994);
xor U3457 (N_3457,N_2099,N_1709);
xnor U3458 (N_3458,N_1665,N_2247);
or U3459 (N_3459,N_2122,N_1359);
nand U3460 (N_3460,N_2024,N_1582);
or U3461 (N_3461,N_2393,N_1908);
or U3462 (N_3462,N_1321,N_1525);
nor U3463 (N_3463,N_2201,N_1976);
nand U3464 (N_3464,N_2157,N_2358);
or U3465 (N_3465,N_2276,N_1627);
or U3466 (N_3466,N_1551,N_2400);
xor U3467 (N_3467,N_1918,N_1257);
nand U3468 (N_3468,N_1695,N_2101);
nand U3469 (N_3469,N_1795,N_1970);
and U3470 (N_3470,N_1430,N_1554);
nor U3471 (N_3471,N_2062,N_2412);
nor U3472 (N_3472,N_2204,N_2396);
or U3473 (N_3473,N_2220,N_1390);
xnor U3474 (N_3474,N_1420,N_1401);
and U3475 (N_3475,N_1692,N_2316);
or U3476 (N_3476,N_1481,N_2316);
nor U3477 (N_3477,N_1269,N_1337);
and U3478 (N_3478,N_1922,N_2397);
or U3479 (N_3479,N_1444,N_1295);
nor U3480 (N_3480,N_1455,N_2335);
nand U3481 (N_3481,N_1521,N_1862);
or U3482 (N_3482,N_2402,N_1340);
and U3483 (N_3483,N_1588,N_2353);
nor U3484 (N_3484,N_1547,N_1852);
and U3485 (N_3485,N_2026,N_1266);
nor U3486 (N_3486,N_2473,N_2022);
or U3487 (N_3487,N_1553,N_1749);
xor U3488 (N_3488,N_2292,N_2371);
xor U3489 (N_3489,N_1716,N_1873);
and U3490 (N_3490,N_1646,N_2131);
and U3491 (N_3491,N_1844,N_1911);
or U3492 (N_3492,N_1705,N_1710);
xor U3493 (N_3493,N_1797,N_1310);
and U3494 (N_3494,N_1292,N_2080);
or U3495 (N_3495,N_2079,N_1357);
xnor U3496 (N_3496,N_1879,N_2332);
or U3497 (N_3497,N_1343,N_2269);
nand U3498 (N_3498,N_2334,N_1393);
and U3499 (N_3499,N_2276,N_1687);
nor U3500 (N_3500,N_2154,N_1945);
and U3501 (N_3501,N_1734,N_2489);
nor U3502 (N_3502,N_2412,N_2240);
xnor U3503 (N_3503,N_1619,N_1808);
and U3504 (N_3504,N_1783,N_1359);
nor U3505 (N_3505,N_1356,N_2194);
nand U3506 (N_3506,N_1335,N_1309);
nand U3507 (N_3507,N_1833,N_1871);
and U3508 (N_3508,N_1993,N_1885);
and U3509 (N_3509,N_1304,N_1464);
nor U3510 (N_3510,N_1328,N_2072);
xnor U3511 (N_3511,N_1389,N_2498);
and U3512 (N_3512,N_1403,N_2198);
or U3513 (N_3513,N_1638,N_2292);
nor U3514 (N_3514,N_1787,N_2263);
xnor U3515 (N_3515,N_2418,N_1371);
nor U3516 (N_3516,N_1531,N_1380);
xnor U3517 (N_3517,N_1569,N_1551);
nand U3518 (N_3518,N_2256,N_2499);
nand U3519 (N_3519,N_2038,N_1356);
nor U3520 (N_3520,N_1627,N_1298);
xnor U3521 (N_3521,N_1493,N_1692);
nand U3522 (N_3522,N_2383,N_1433);
nand U3523 (N_3523,N_2311,N_1867);
nor U3524 (N_3524,N_1858,N_2405);
nand U3525 (N_3525,N_1797,N_2361);
nand U3526 (N_3526,N_2261,N_2387);
and U3527 (N_3527,N_1521,N_2343);
or U3528 (N_3528,N_1308,N_2159);
nor U3529 (N_3529,N_2129,N_2481);
xor U3530 (N_3530,N_2492,N_2379);
nand U3531 (N_3531,N_2426,N_1773);
nand U3532 (N_3532,N_1497,N_1845);
xor U3533 (N_3533,N_2062,N_2149);
nor U3534 (N_3534,N_1948,N_2391);
and U3535 (N_3535,N_2008,N_1852);
nor U3536 (N_3536,N_1806,N_1865);
and U3537 (N_3537,N_1330,N_1371);
nand U3538 (N_3538,N_1796,N_2290);
nand U3539 (N_3539,N_1447,N_2118);
nor U3540 (N_3540,N_1721,N_1922);
and U3541 (N_3541,N_1942,N_2145);
xnor U3542 (N_3542,N_1472,N_2139);
or U3543 (N_3543,N_1965,N_2043);
xnor U3544 (N_3544,N_2237,N_2351);
or U3545 (N_3545,N_2279,N_1863);
xnor U3546 (N_3546,N_1788,N_2022);
or U3547 (N_3547,N_1802,N_1552);
and U3548 (N_3548,N_1944,N_1460);
or U3549 (N_3549,N_2269,N_1808);
and U3550 (N_3550,N_1433,N_2173);
xnor U3551 (N_3551,N_2302,N_2367);
xnor U3552 (N_3552,N_2413,N_2255);
nand U3553 (N_3553,N_1801,N_1988);
nand U3554 (N_3554,N_1943,N_2425);
nor U3555 (N_3555,N_2372,N_1673);
xor U3556 (N_3556,N_1986,N_2116);
nor U3557 (N_3557,N_1718,N_1326);
nor U3558 (N_3558,N_2472,N_2388);
and U3559 (N_3559,N_1986,N_1415);
and U3560 (N_3560,N_1396,N_2383);
xnor U3561 (N_3561,N_2352,N_1458);
or U3562 (N_3562,N_1507,N_1615);
or U3563 (N_3563,N_1339,N_2085);
and U3564 (N_3564,N_1478,N_2204);
and U3565 (N_3565,N_1511,N_1891);
xnor U3566 (N_3566,N_1695,N_1290);
and U3567 (N_3567,N_2080,N_1460);
xor U3568 (N_3568,N_1873,N_1797);
nor U3569 (N_3569,N_2332,N_1723);
and U3570 (N_3570,N_2009,N_1683);
or U3571 (N_3571,N_1522,N_2012);
or U3572 (N_3572,N_1367,N_2479);
and U3573 (N_3573,N_2149,N_1956);
and U3574 (N_3574,N_1521,N_1945);
nand U3575 (N_3575,N_1851,N_1545);
nor U3576 (N_3576,N_2236,N_1486);
or U3577 (N_3577,N_2255,N_2132);
and U3578 (N_3578,N_2363,N_1696);
xnor U3579 (N_3579,N_1965,N_1517);
xnor U3580 (N_3580,N_2089,N_1868);
or U3581 (N_3581,N_2337,N_1339);
and U3582 (N_3582,N_1846,N_1413);
nor U3583 (N_3583,N_2354,N_1653);
nand U3584 (N_3584,N_1285,N_1485);
nand U3585 (N_3585,N_2490,N_1583);
and U3586 (N_3586,N_1976,N_1253);
and U3587 (N_3587,N_1383,N_1619);
xnor U3588 (N_3588,N_1674,N_1475);
and U3589 (N_3589,N_2415,N_2086);
and U3590 (N_3590,N_1725,N_1337);
or U3591 (N_3591,N_1534,N_1859);
or U3592 (N_3592,N_1304,N_2428);
nand U3593 (N_3593,N_2088,N_2272);
and U3594 (N_3594,N_1314,N_2151);
nand U3595 (N_3595,N_1405,N_1371);
xnor U3596 (N_3596,N_2237,N_1684);
or U3597 (N_3597,N_1790,N_2225);
or U3598 (N_3598,N_2025,N_1290);
xor U3599 (N_3599,N_1461,N_1375);
xnor U3600 (N_3600,N_1803,N_1388);
nor U3601 (N_3601,N_1525,N_2152);
and U3602 (N_3602,N_1327,N_1509);
xor U3603 (N_3603,N_2242,N_1802);
and U3604 (N_3604,N_2116,N_2160);
or U3605 (N_3605,N_1398,N_2315);
xor U3606 (N_3606,N_2438,N_2446);
nand U3607 (N_3607,N_1605,N_1788);
and U3608 (N_3608,N_1893,N_1622);
xnor U3609 (N_3609,N_2411,N_2420);
and U3610 (N_3610,N_1729,N_1870);
xnor U3611 (N_3611,N_2068,N_1734);
and U3612 (N_3612,N_1512,N_2104);
or U3613 (N_3613,N_1382,N_1352);
and U3614 (N_3614,N_1345,N_1289);
or U3615 (N_3615,N_1887,N_1586);
or U3616 (N_3616,N_2308,N_1668);
and U3617 (N_3617,N_2297,N_2366);
xor U3618 (N_3618,N_1270,N_1908);
xnor U3619 (N_3619,N_1259,N_2102);
and U3620 (N_3620,N_1781,N_1715);
xor U3621 (N_3621,N_1945,N_1992);
and U3622 (N_3622,N_1921,N_2011);
xor U3623 (N_3623,N_1387,N_2405);
or U3624 (N_3624,N_2343,N_1998);
xor U3625 (N_3625,N_2482,N_2391);
nor U3626 (N_3626,N_1318,N_2414);
nand U3627 (N_3627,N_2368,N_1455);
and U3628 (N_3628,N_1990,N_1825);
and U3629 (N_3629,N_2474,N_2186);
or U3630 (N_3630,N_2012,N_2470);
or U3631 (N_3631,N_1641,N_2411);
nor U3632 (N_3632,N_1840,N_1564);
or U3633 (N_3633,N_1554,N_2230);
and U3634 (N_3634,N_2023,N_1723);
nor U3635 (N_3635,N_2458,N_1875);
nor U3636 (N_3636,N_1858,N_2371);
nand U3637 (N_3637,N_2088,N_2095);
nor U3638 (N_3638,N_1997,N_2177);
nor U3639 (N_3639,N_2042,N_1408);
and U3640 (N_3640,N_1342,N_2491);
or U3641 (N_3641,N_1651,N_1675);
nand U3642 (N_3642,N_2186,N_1691);
and U3643 (N_3643,N_1660,N_1860);
nor U3644 (N_3644,N_2266,N_2001);
nor U3645 (N_3645,N_2063,N_1812);
or U3646 (N_3646,N_1661,N_1482);
xor U3647 (N_3647,N_1340,N_2498);
or U3648 (N_3648,N_1870,N_2262);
or U3649 (N_3649,N_2241,N_2009);
or U3650 (N_3650,N_1848,N_2306);
and U3651 (N_3651,N_1598,N_1997);
nand U3652 (N_3652,N_2285,N_2479);
or U3653 (N_3653,N_1618,N_2468);
xnor U3654 (N_3654,N_1829,N_2354);
nor U3655 (N_3655,N_1623,N_1457);
and U3656 (N_3656,N_1815,N_1823);
or U3657 (N_3657,N_2290,N_1409);
or U3658 (N_3658,N_2380,N_1874);
or U3659 (N_3659,N_1589,N_1840);
nor U3660 (N_3660,N_1789,N_2292);
nand U3661 (N_3661,N_2049,N_1312);
or U3662 (N_3662,N_1271,N_2313);
nor U3663 (N_3663,N_1372,N_2227);
and U3664 (N_3664,N_2443,N_2418);
or U3665 (N_3665,N_2040,N_1490);
or U3666 (N_3666,N_2050,N_1538);
nor U3667 (N_3667,N_1670,N_1358);
xnor U3668 (N_3668,N_1903,N_2340);
nor U3669 (N_3669,N_2182,N_1421);
xnor U3670 (N_3670,N_2214,N_1991);
xnor U3671 (N_3671,N_1896,N_1764);
or U3672 (N_3672,N_2142,N_2177);
xnor U3673 (N_3673,N_1804,N_2006);
xnor U3674 (N_3674,N_2385,N_1573);
xor U3675 (N_3675,N_1585,N_2359);
or U3676 (N_3676,N_1671,N_1433);
nor U3677 (N_3677,N_1999,N_1257);
or U3678 (N_3678,N_1807,N_1257);
nor U3679 (N_3679,N_1912,N_1748);
and U3680 (N_3680,N_2178,N_2377);
nand U3681 (N_3681,N_1856,N_2333);
xor U3682 (N_3682,N_1390,N_1536);
xor U3683 (N_3683,N_1396,N_1938);
and U3684 (N_3684,N_2301,N_1276);
nor U3685 (N_3685,N_2497,N_1737);
and U3686 (N_3686,N_1694,N_2485);
or U3687 (N_3687,N_1526,N_1945);
and U3688 (N_3688,N_1972,N_1407);
nand U3689 (N_3689,N_1964,N_2319);
nand U3690 (N_3690,N_2345,N_2110);
nand U3691 (N_3691,N_2105,N_2377);
nor U3692 (N_3692,N_2133,N_2457);
and U3693 (N_3693,N_2483,N_1934);
nand U3694 (N_3694,N_1266,N_1993);
or U3695 (N_3695,N_1412,N_1785);
nor U3696 (N_3696,N_1812,N_2013);
and U3697 (N_3697,N_1919,N_2454);
nand U3698 (N_3698,N_1803,N_1849);
xnor U3699 (N_3699,N_1485,N_2389);
and U3700 (N_3700,N_2156,N_2477);
nor U3701 (N_3701,N_1699,N_1438);
nor U3702 (N_3702,N_1937,N_1351);
nor U3703 (N_3703,N_1860,N_1328);
nand U3704 (N_3704,N_2405,N_1625);
and U3705 (N_3705,N_2138,N_1662);
and U3706 (N_3706,N_1309,N_2389);
and U3707 (N_3707,N_1483,N_1382);
xor U3708 (N_3708,N_1443,N_2416);
and U3709 (N_3709,N_2093,N_2055);
or U3710 (N_3710,N_2380,N_1462);
nand U3711 (N_3711,N_2255,N_1657);
xor U3712 (N_3712,N_1467,N_1458);
nand U3713 (N_3713,N_2358,N_2125);
and U3714 (N_3714,N_1921,N_2399);
and U3715 (N_3715,N_1253,N_1277);
nand U3716 (N_3716,N_1803,N_1896);
nor U3717 (N_3717,N_2273,N_2476);
or U3718 (N_3718,N_1414,N_2092);
or U3719 (N_3719,N_1789,N_2024);
and U3720 (N_3720,N_2457,N_1897);
xnor U3721 (N_3721,N_2408,N_2418);
and U3722 (N_3722,N_2350,N_2484);
nand U3723 (N_3723,N_1281,N_2451);
or U3724 (N_3724,N_2459,N_2083);
or U3725 (N_3725,N_1444,N_2227);
nor U3726 (N_3726,N_1552,N_1701);
nand U3727 (N_3727,N_2440,N_1704);
xor U3728 (N_3728,N_1698,N_1544);
or U3729 (N_3729,N_2413,N_2471);
xor U3730 (N_3730,N_2351,N_2071);
nor U3731 (N_3731,N_2367,N_1573);
nor U3732 (N_3732,N_1339,N_1696);
xnor U3733 (N_3733,N_1987,N_2341);
and U3734 (N_3734,N_2212,N_2472);
or U3735 (N_3735,N_2124,N_1666);
nor U3736 (N_3736,N_2148,N_2222);
or U3737 (N_3737,N_1540,N_2359);
xnor U3738 (N_3738,N_2005,N_2247);
xor U3739 (N_3739,N_2379,N_2162);
nand U3740 (N_3740,N_2188,N_1546);
or U3741 (N_3741,N_1934,N_1744);
nor U3742 (N_3742,N_1891,N_1892);
or U3743 (N_3743,N_1981,N_1677);
or U3744 (N_3744,N_2340,N_2025);
and U3745 (N_3745,N_1827,N_2460);
nor U3746 (N_3746,N_1565,N_2403);
nand U3747 (N_3747,N_1605,N_1926);
nand U3748 (N_3748,N_2267,N_1945);
nor U3749 (N_3749,N_1974,N_2242);
or U3750 (N_3750,N_3746,N_2535);
xor U3751 (N_3751,N_2915,N_3645);
xor U3752 (N_3752,N_3280,N_2798);
and U3753 (N_3753,N_3735,N_2839);
nor U3754 (N_3754,N_2613,N_2628);
xnor U3755 (N_3755,N_3344,N_3018);
nand U3756 (N_3756,N_2514,N_3202);
and U3757 (N_3757,N_3251,N_2893);
or U3758 (N_3758,N_3697,N_3462);
or U3759 (N_3759,N_3161,N_2638);
or U3760 (N_3760,N_3184,N_3654);
or U3761 (N_3761,N_2892,N_3110);
and U3762 (N_3762,N_3001,N_2978);
and U3763 (N_3763,N_2994,N_3372);
or U3764 (N_3764,N_3635,N_3207);
or U3765 (N_3765,N_3333,N_3568);
nand U3766 (N_3766,N_2552,N_2682);
xnor U3767 (N_3767,N_3565,N_3718);
or U3768 (N_3768,N_2887,N_2528);
and U3769 (N_3769,N_3504,N_2508);
nand U3770 (N_3770,N_2689,N_2672);
or U3771 (N_3771,N_3640,N_3113);
nor U3772 (N_3772,N_3237,N_2963);
or U3773 (N_3773,N_3498,N_2569);
xnor U3774 (N_3774,N_2600,N_3392);
nor U3775 (N_3775,N_2766,N_3408);
and U3776 (N_3776,N_3091,N_3115);
nor U3777 (N_3777,N_2663,N_3527);
nor U3778 (N_3778,N_3085,N_2862);
and U3779 (N_3779,N_3288,N_2803);
nor U3780 (N_3780,N_3573,N_3170);
xnor U3781 (N_3781,N_3402,N_2657);
and U3782 (N_3782,N_3013,N_3246);
or U3783 (N_3783,N_2800,N_3103);
nor U3784 (N_3784,N_3253,N_2815);
xnor U3785 (N_3785,N_3206,N_2807);
xor U3786 (N_3786,N_2639,N_3081);
xnor U3787 (N_3787,N_3519,N_2922);
nor U3788 (N_3788,N_2937,N_3379);
nand U3789 (N_3789,N_3455,N_2531);
nand U3790 (N_3790,N_3482,N_2885);
xor U3791 (N_3791,N_2617,N_3446);
nand U3792 (N_3792,N_3529,N_3588);
or U3793 (N_3793,N_3129,N_2987);
or U3794 (N_3794,N_3471,N_3658);
and U3795 (N_3795,N_2858,N_2995);
and U3796 (N_3796,N_3359,N_3003);
nor U3797 (N_3797,N_3114,N_3215);
nor U3798 (N_3798,N_3511,N_3044);
nor U3799 (N_3799,N_3581,N_2952);
nand U3800 (N_3800,N_2897,N_3647);
or U3801 (N_3801,N_3286,N_3008);
xnor U3802 (N_3802,N_2914,N_2556);
xnor U3803 (N_3803,N_2630,N_3499);
nor U3804 (N_3804,N_3712,N_3046);
or U3805 (N_3805,N_3281,N_2721);
and U3806 (N_3806,N_2704,N_3266);
nor U3807 (N_3807,N_2898,N_3643);
or U3808 (N_3808,N_3602,N_3101);
or U3809 (N_3809,N_3358,N_2966);
nor U3810 (N_3810,N_2668,N_3692);
nand U3811 (N_3811,N_3138,N_3211);
nand U3812 (N_3812,N_3421,N_3283);
nor U3813 (N_3813,N_3648,N_3316);
xnor U3814 (N_3814,N_2609,N_2890);
or U3815 (N_3815,N_2678,N_2680);
nor U3816 (N_3816,N_2601,N_2685);
nand U3817 (N_3817,N_3586,N_3739);
nand U3818 (N_3818,N_2566,N_3728);
nand U3819 (N_3819,N_3450,N_3339);
or U3820 (N_3820,N_3153,N_3135);
and U3821 (N_3821,N_3158,N_2542);
xnor U3822 (N_3822,N_2733,N_2673);
nor U3823 (N_3823,N_2716,N_2855);
and U3824 (N_3824,N_3104,N_3190);
nand U3825 (N_3825,N_3488,N_3249);
and U3826 (N_3826,N_3341,N_3652);
xor U3827 (N_3827,N_2539,N_3025);
and U3828 (N_3828,N_3078,N_2618);
nand U3829 (N_3829,N_3730,N_2957);
nand U3830 (N_3830,N_3520,N_3166);
nand U3831 (N_3831,N_2857,N_3089);
or U3832 (N_3832,N_2500,N_2517);
or U3833 (N_3833,N_3199,N_3047);
xor U3834 (N_3834,N_2582,N_2801);
xor U3835 (N_3835,N_2882,N_3328);
or U3836 (N_3836,N_3209,N_3084);
and U3837 (N_3837,N_3053,N_2510);
and U3838 (N_3838,N_2873,N_2782);
or U3839 (N_3839,N_2808,N_2547);
xor U3840 (N_3840,N_2718,N_3235);
nor U3841 (N_3841,N_3245,N_2606);
or U3842 (N_3842,N_3442,N_2503);
and U3843 (N_3843,N_2632,N_3416);
xnor U3844 (N_3844,N_3418,N_3345);
and U3845 (N_3845,N_3272,N_3304);
xnor U3846 (N_3846,N_2753,N_2841);
and U3847 (N_3847,N_3478,N_2749);
and U3848 (N_3848,N_3186,N_2777);
nand U3849 (N_3849,N_3031,N_3284);
nand U3850 (N_3850,N_2760,N_3323);
xnor U3851 (N_3851,N_2975,N_2602);
and U3852 (N_3852,N_3256,N_3381);
nand U3853 (N_3853,N_2828,N_3729);
or U3854 (N_3854,N_3632,N_3373);
or U3855 (N_3855,N_2834,N_3725);
and U3856 (N_3856,N_3733,N_2652);
nand U3857 (N_3857,N_3247,N_2959);
nor U3858 (N_3858,N_2674,N_3724);
nand U3859 (N_3859,N_3193,N_3386);
or U3860 (N_3860,N_3131,N_2852);
xnor U3861 (N_3861,N_2736,N_3100);
and U3862 (N_3862,N_3585,N_3298);
or U3863 (N_3863,N_3150,N_3234);
xnor U3864 (N_3864,N_3447,N_2844);
nand U3865 (N_3865,N_2504,N_2709);
xor U3866 (N_3866,N_3558,N_3415);
nor U3867 (N_3867,N_3465,N_2686);
nor U3868 (N_3868,N_2579,N_3065);
and U3869 (N_3869,N_3255,N_3722);
or U3870 (N_3870,N_3472,N_3659);
nand U3871 (N_3871,N_3321,N_3370);
nor U3872 (N_3872,N_3587,N_3507);
and U3873 (N_3873,N_2883,N_2905);
and U3874 (N_3874,N_3680,N_3723);
nand U3875 (N_3875,N_3136,N_3183);
xnor U3876 (N_3876,N_2856,N_3140);
xor U3877 (N_3877,N_3006,N_2512);
and U3878 (N_3878,N_3367,N_3411);
nand U3879 (N_3879,N_3142,N_3570);
nor U3880 (N_3880,N_3577,N_3603);
and U3881 (N_3881,N_3315,N_3634);
or U3882 (N_3882,N_3282,N_3483);
nand U3883 (N_3883,N_2605,N_3144);
nand U3884 (N_3884,N_2543,N_3277);
nand U3885 (N_3885,N_2977,N_2710);
xor U3886 (N_3886,N_3584,N_3137);
nor U3887 (N_3887,N_3351,N_2763);
nand U3888 (N_3888,N_3492,N_3546);
or U3889 (N_3889,N_3306,N_3525);
or U3890 (N_3890,N_3117,N_3204);
nor U3891 (N_3891,N_3530,N_3238);
nor U3892 (N_3892,N_3516,N_3571);
xor U3893 (N_3893,N_2973,N_3497);
or U3894 (N_3894,N_2776,N_3484);
and U3895 (N_3895,N_3685,N_2818);
and U3896 (N_3896,N_2967,N_3629);
or U3897 (N_3897,N_3133,N_2806);
xnor U3898 (N_3898,N_2594,N_3655);
nor U3899 (N_3899,N_2551,N_2746);
or U3900 (N_3900,N_3145,N_3096);
nor U3901 (N_3901,N_3696,N_3179);
nor U3902 (N_3902,N_2541,N_3064);
nor U3903 (N_3903,N_3703,N_3412);
or U3904 (N_3904,N_3325,N_2846);
nor U3905 (N_3905,N_3580,N_3627);
or U3906 (N_3906,N_2772,N_2854);
or U3907 (N_3907,N_2635,N_3120);
nand U3908 (N_3908,N_3661,N_2820);
or U3909 (N_3909,N_2793,N_3087);
xnor U3910 (N_3910,N_2990,N_3311);
nand U3911 (N_3911,N_3335,N_3268);
nand U3912 (N_3912,N_3678,N_2565);
or U3913 (N_3913,N_3010,N_2532);
nor U3914 (N_3914,N_3710,N_3317);
nor U3915 (N_3915,N_3363,N_2636);
and U3916 (N_3916,N_2879,N_2513);
nor U3917 (N_3917,N_3670,N_2965);
nor U3918 (N_3918,N_3664,N_2706);
nand U3919 (N_3919,N_3689,N_3644);
and U3920 (N_3920,N_3107,N_2592);
and U3921 (N_3921,N_2786,N_3254);
nor U3922 (N_3922,N_3506,N_2522);
nor U3923 (N_3923,N_3252,N_2545);
xnor U3924 (N_3924,N_2688,N_2928);
xor U3925 (N_3925,N_3210,N_2518);
nand U3926 (N_3926,N_2765,N_3320);
or U3927 (N_3927,N_3486,N_3226);
and U3928 (N_3928,N_2744,N_3657);
nor U3929 (N_3929,N_3651,N_2620);
or U3930 (N_3930,N_3364,N_3123);
or U3931 (N_3931,N_3083,N_3687);
or U3932 (N_3932,N_3174,N_2923);
and U3933 (N_3933,N_3023,N_2829);
and U3934 (N_3934,N_2822,N_3289);
nand U3935 (N_3935,N_3036,N_3308);
xor U3936 (N_3936,N_3708,N_3460);
or U3937 (N_3937,N_2720,N_3633);
and U3938 (N_3938,N_2738,N_2607);
nor U3939 (N_3939,N_2562,N_3297);
or U3940 (N_3940,N_3350,N_2864);
xor U3941 (N_3941,N_2802,N_3290);
or U3942 (N_3942,N_3613,N_2627);
nor U3943 (N_3943,N_3093,N_3334);
nand U3944 (N_3944,N_3691,N_2788);
or U3945 (N_3945,N_3265,N_2794);
nor U3946 (N_3946,N_2708,N_2727);
or U3947 (N_3947,N_2875,N_2523);
nand U3948 (N_3948,N_2906,N_3560);
nand U3949 (N_3949,N_2516,N_2701);
or U3950 (N_3950,N_3324,N_2859);
or U3951 (N_3951,N_3600,N_2830);
nor U3952 (N_3952,N_3074,N_3192);
and U3953 (N_3953,N_3720,N_2988);
xnor U3954 (N_3954,N_3239,N_3688);
nor U3955 (N_3955,N_2671,N_2976);
xor U3956 (N_3956,N_3354,N_3062);
or U3957 (N_3957,N_3075,N_3676);
nor U3958 (N_3958,N_2571,N_3141);
nand U3959 (N_3959,N_3068,N_2946);
or U3960 (N_3960,N_3342,N_3189);
or U3961 (N_3961,N_2544,N_3662);
nor U3962 (N_3962,N_2929,N_2936);
nor U3963 (N_3963,N_2889,N_3221);
and U3964 (N_3964,N_3072,N_2693);
nand U3965 (N_3965,N_2986,N_2947);
or U3966 (N_3966,N_3267,N_3737);
nand U3967 (N_3967,N_3242,N_2865);
or U3968 (N_3968,N_2527,N_2867);
and U3969 (N_3969,N_3149,N_3305);
nand U3970 (N_3970,N_3332,N_3329);
or U3971 (N_3971,N_3673,N_3452);
xnor U3972 (N_3972,N_3512,N_2519);
or U3973 (N_3973,N_3715,N_2762);
nor U3974 (N_3974,N_3213,N_2590);
nor U3975 (N_3975,N_2961,N_2904);
nand U3976 (N_3976,N_2884,N_2938);
nor U3977 (N_3977,N_2622,N_3555);
nand U3978 (N_3978,N_3212,N_3294);
or U3979 (N_3979,N_3404,N_3625);
xor U3980 (N_3980,N_3071,N_2707);
and U3981 (N_3981,N_3532,N_3377);
nor U3982 (N_3982,N_3427,N_2679);
nor U3983 (N_3983,N_3171,N_2741);
xnor U3984 (N_3984,N_2730,N_2833);
nand U3985 (N_3985,N_2623,N_2648);
or U3986 (N_3986,N_3671,N_3719);
or U3987 (N_3987,N_3606,N_2950);
nand U3988 (N_3988,N_2548,N_2717);
or U3989 (N_3989,N_3033,N_2700);
xnor U3990 (N_3990,N_2538,N_3572);
xnor U3991 (N_3991,N_3638,N_3596);
and U3992 (N_3992,N_3407,N_2814);
and U3993 (N_3993,N_3727,N_2525);
nand U3994 (N_3994,N_2868,N_3597);
and U3995 (N_3995,N_3000,N_3011);
nor U3996 (N_3996,N_3420,N_3626);
nor U3997 (N_3997,N_2759,N_3445);
or U3998 (N_3998,N_3491,N_3399);
nand U3999 (N_3999,N_2932,N_2810);
nand U4000 (N_4000,N_3086,N_2780);
or U4001 (N_4001,N_3194,N_2615);
nand U4002 (N_4002,N_3566,N_2916);
nor U4003 (N_4003,N_3463,N_3028);
xnor U4004 (N_4004,N_2956,N_3738);
nand U4005 (N_4005,N_2642,N_3535);
nor U4006 (N_4006,N_2930,N_3132);
nand U4007 (N_4007,N_3473,N_2901);
nand U4008 (N_4008,N_2939,N_2984);
or U4009 (N_4009,N_2999,N_2560);
nand U4010 (N_4010,N_2944,N_3037);
xnor U4011 (N_4011,N_3395,N_3424);
and U4012 (N_4012,N_3203,N_2764);
xnor U4013 (N_4013,N_2624,N_3610);
or U4014 (N_4014,N_3128,N_2913);
nand U4015 (N_4015,N_2831,N_3160);
nand U4016 (N_4016,N_3517,N_2921);
and U4017 (N_4017,N_3437,N_3459);
xnor U4018 (N_4018,N_2586,N_3466);
nand U4019 (N_4019,N_2752,N_3514);
nor U4020 (N_4020,N_3705,N_3742);
xnor U4021 (N_4021,N_2537,N_3551);
nor U4022 (N_4022,N_2908,N_2811);
and U4023 (N_4023,N_2506,N_3164);
nor U4024 (N_4024,N_2949,N_3076);
or U4025 (N_4025,N_3595,N_3749);
and U4026 (N_4026,N_3624,N_3225);
nand U4027 (N_4027,N_2895,N_3021);
nor U4028 (N_4028,N_3667,N_3677);
nor U4029 (N_4029,N_2821,N_2970);
and U4030 (N_4030,N_2781,N_3291);
or U4031 (N_4031,N_2964,N_2789);
and U4032 (N_4032,N_2874,N_3337);
and U4033 (N_4033,N_3059,N_3621);
nor U4034 (N_4034,N_2835,N_3605);
and U4035 (N_4035,N_2604,N_3244);
and U4036 (N_4036,N_2920,N_3102);
nand U4037 (N_4037,N_2646,N_2511);
and U4038 (N_4038,N_2665,N_2809);
and U4039 (N_4039,N_3653,N_2758);
xnor U4040 (N_4040,N_3574,N_3061);
xor U4041 (N_4041,N_3043,N_2667);
and U4042 (N_4042,N_3388,N_3554);
nand U4043 (N_4043,N_2953,N_3721);
nor U4044 (N_4044,N_3550,N_2585);
nand U4045 (N_4045,N_2583,N_2558);
or U4046 (N_4046,N_3544,N_3711);
and U4047 (N_4047,N_2747,N_3663);
xnor U4048 (N_4048,N_3400,N_3589);
and U4049 (N_4049,N_2998,N_3243);
nor U4050 (N_4050,N_3575,N_2694);
nand U4051 (N_4051,N_3200,N_3438);
nor U4052 (N_4052,N_2917,N_2722);
or U4053 (N_4053,N_3152,N_3361);
nor U4054 (N_4054,N_2783,N_2641);
and U4055 (N_4055,N_2843,N_3612);
nand U4056 (N_4056,N_3156,N_3187);
nand U4057 (N_4057,N_3429,N_2726);
xor U4058 (N_4058,N_3105,N_2825);
nor U4059 (N_4059,N_3146,N_2728);
nor U4060 (N_4060,N_3229,N_2817);
nor U4061 (N_4061,N_3642,N_3690);
nand U4062 (N_4062,N_2750,N_3155);
and U4063 (N_4063,N_2832,N_2546);
nand U4064 (N_4064,N_2725,N_3111);
nor U4065 (N_4065,N_3278,N_3414);
xnor U4066 (N_4066,N_3479,N_3646);
xor U4067 (N_4067,N_3263,N_2732);
nand U4068 (N_4068,N_2591,N_3014);
xnor U4069 (N_4069,N_3302,N_2712);
nor U4070 (N_4070,N_2982,N_3716);
nand U4071 (N_4071,N_3167,N_3134);
or U4072 (N_4072,N_3461,N_3318);
xor U4073 (N_4073,N_2666,N_3604);
nand U4074 (N_4074,N_2894,N_2971);
nor U4075 (N_4075,N_3599,N_3041);
nor U4076 (N_4076,N_2612,N_2827);
nand U4077 (N_4077,N_2756,N_3090);
or U4078 (N_4078,N_3177,N_2723);
and U4079 (N_4079,N_3173,N_3347);
and U4080 (N_4080,N_3224,N_2735);
and U4081 (N_4081,N_3116,N_2683);
nor U4082 (N_4082,N_3223,N_2691);
nand U4083 (N_4083,N_3458,N_2796);
xor U4084 (N_4084,N_3387,N_2941);
and U4085 (N_4085,N_3668,N_3564);
or U4086 (N_4086,N_2664,N_3607);
nor U4087 (N_4087,N_3172,N_3393);
or U4088 (N_4088,N_3143,N_3451);
nor U4089 (N_4089,N_2863,N_2595);
or U4090 (N_4090,N_3453,N_3269);
nand U4091 (N_4091,N_3054,N_2634);
nor U4092 (N_4092,N_3614,N_3180);
nand U4093 (N_4093,N_3509,N_3258);
xnor U4094 (N_4094,N_2838,N_3348);
nor U4095 (N_4095,N_3262,N_3410);
nand U4096 (N_4096,N_3413,N_2611);
or U4097 (N_4097,N_2849,N_3030);
and U4098 (N_4098,N_3518,N_3608);
nand U4099 (N_4099,N_3502,N_3549);
nand U4100 (N_4100,N_3618,N_3496);
nor U4101 (N_4101,N_3683,N_3057);
xnor U4102 (N_4102,N_3403,N_3489);
and U4103 (N_4103,N_2853,N_3045);
nor U4104 (N_4104,N_3169,N_3476);
and U4105 (N_4105,N_2697,N_3079);
and U4106 (N_4106,N_3139,N_3250);
nor U4107 (N_4107,N_3349,N_3524);
xor U4108 (N_4108,N_3552,N_3469);
nor U4109 (N_4109,N_3563,N_3579);
or U4110 (N_4110,N_2851,N_3362);
nor U4111 (N_4111,N_3205,N_3326);
and U4112 (N_4112,N_3679,N_2869);
xnor U4113 (N_4113,N_2935,N_3314);
nand U4114 (N_4114,N_2757,N_3039);
and U4115 (N_4115,N_3521,N_2816);
or U4116 (N_4116,N_2737,N_3396);
nor U4117 (N_4117,N_3425,N_3649);
and U4118 (N_4118,N_3456,N_2669);
nand U4119 (N_4119,N_3701,N_2633);
or U4120 (N_4120,N_2596,N_2713);
or U4121 (N_4121,N_3380,N_3576);
xnor U4122 (N_4122,N_3553,N_2909);
nand U4123 (N_4123,N_2681,N_2509);
or U4124 (N_4124,N_2872,N_3292);
nor U4125 (N_4125,N_2954,N_3300);
or U4126 (N_4126,N_3531,N_3195);
or U4127 (N_4127,N_3623,N_2677);
and U4128 (N_4128,N_2554,N_3038);
and U4129 (N_4129,N_2926,N_2589);
nor U4130 (N_4130,N_3271,N_2848);
xnor U4131 (N_4131,N_3434,N_2515);
xor U4132 (N_4132,N_3108,N_3175);
and U4133 (N_4133,N_2770,N_3055);
nor U4134 (N_4134,N_3748,N_3409);
xor U4135 (N_4135,N_3162,N_3261);
or U4136 (N_4136,N_2881,N_3285);
or U4137 (N_4137,N_3686,N_2540);
nor U4138 (N_4138,N_3422,N_3660);
or U4139 (N_4139,N_2695,N_2925);
nand U4140 (N_4140,N_3016,N_3622);
xnor U4141 (N_4141,N_3126,N_2651);
and U4142 (N_4142,N_2570,N_3371);
nor U4143 (N_4143,N_3695,N_3168);
and U4144 (N_4144,N_2751,N_3222);
nand U4145 (N_4145,N_3481,N_2563);
or U4146 (N_4146,N_3216,N_3214);
xnor U4147 (N_4147,N_2597,N_3449);
xnor U4148 (N_4148,N_2645,N_3240);
or U4149 (N_4149,N_2813,N_3248);
xnor U4150 (N_4150,N_2980,N_3009);
and U4151 (N_4151,N_2989,N_2779);
nor U4152 (N_4152,N_3656,N_3032);
nand U4153 (N_4153,N_2837,N_2880);
and U4154 (N_4154,N_3352,N_3109);
nand U4155 (N_4155,N_2711,N_3219);
and U4156 (N_4156,N_3440,N_2661);
and U4157 (N_4157,N_3547,N_2553);
and U4158 (N_4158,N_2996,N_3260);
nand U4159 (N_4159,N_3196,N_2690);
or U4160 (N_4160,N_2724,N_2577);
and U4161 (N_4161,N_3112,N_3448);
nor U4162 (N_4162,N_3034,N_3556);
or U4163 (N_4163,N_3148,N_2584);
and U4164 (N_4164,N_2945,N_3557);
or U4165 (N_4165,N_2745,N_3704);
nand U4166 (N_4166,N_3378,N_2997);
or U4167 (N_4167,N_2819,N_3060);
xor U4168 (N_4168,N_3307,N_3287);
or U4169 (N_4169,N_3376,N_2608);
nor U4170 (N_4170,N_2888,N_3313);
nor U4171 (N_4171,N_3383,N_3699);
xnor U4172 (N_4172,N_3389,N_3127);
nand U4173 (N_4173,N_3510,N_3665);
nor U4174 (N_4174,N_2911,N_2847);
nor U4175 (N_4175,N_3616,N_2771);
and U4176 (N_4176,N_2637,N_3515);
xor U4177 (N_4177,N_3233,N_2699);
nor U4178 (N_4178,N_2742,N_2769);
and U4179 (N_4179,N_3503,N_3569);
or U4180 (N_4180,N_2900,N_3220);
nor U4181 (N_4181,N_3002,N_3098);
nor U4182 (N_4182,N_3346,N_3181);
and U4183 (N_4183,N_2878,N_2974);
nor U4184 (N_4184,N_3092,N_2924);
and U4185 (N_4185,N_2629,N_3274);
or U4186 (N_4186,N_3619,N_2962);
nor U4187 (N_4187,N_2649,N_3375);
and U4188 (N_4188,N_3706,N_3147);
nor U4189 (N_4189,N_3468,N_3747);
or U4190 (N_4190,N_3609,N_3543);
nor U4191 (N_4191,N_2567,N_2983);
or U4192 (N_4192,N_3391,N_2576);
nor U4193 (N_4193,N_2580,N_2731);
xnor U4194 (N_4194,N_2631,N_3693);
and U4195 (N_4195,N_3312,N_3390);
and U4196 (N_4196,N_3188,N_2655);
or U4197 (N_4197,N_2739,N_3590);
and U4198 (N_4198,N_3495,N_3106);
nand U4199 (N_4199,N_3119,N_2530);
nor U4200 (N_4200,N_3264,N_3682);
and U4201 (N_4201,N_2703,N_3464);
or U4202 (N_4202,N_2588,N_2658);
nand U4203 (N_4203,N_3443,N_3198);
xor U4204 (N_4204,N_3004,N_3017);
and U4205 (N_4205,N_3165,N_3330);
nand U4206 (N_4206,N_3401,N_3594);
nor U4207 (N_4207,N_3500,N_2992);
nand U4208 (N_4208,N_3592,N_3508);
nand U4209 (N_4209,N_3698,N_2581);
and U4210 (N_4210,N_3217,N_3230);
nand U4211 (N_4211,N_2714,N_3441);
and U4212 (N_4212,N_2696,N_2774);
and U4213 (N_4213,N_3340,N_2871);
or U4214 (N_4214,N_3366,N_2734);
nand U4215 (N_4215,N_2670,N_2823);
nor U4216 (N_4216,N_2991,N_3731);
nand U4217 (N_4217,N_3545,N_2536);
nand U4218 (N_4218,N_3435,N_2910);
xor U4219 (N_4219,N_2931,N_3433);
nand U4220 (N_4220,N_2505,N_3601);
xnor U4221 (N_4221,N_2981,N_3365);
nor U4222 (N_4222,N_3490,N_2740);
and U4223 (N_4223,N_3331,N_3026);
nor U4224 (N_4224,N_3295,N_2549);
nand U4225 (N_4225,N_3709,N_2768);
nor U4226 (N_4226,N_3533,N_3501);
and U4227 (N_4227,N_3369,N_3431);
or U4228 (N_4228,N_3385,N_3082);
and U4229 (N_4229,N_2876,N_2919);
and U4230 (N_4230,N_3005,N_3562);
and U4231 (N_4231,N_2785,N_2861);
and U4232 (N_4232,N_3713,N_2775);
or U4233 (N_4233,N_2795,N_3430);
and U4234 (N_4234,N_3548,N_3069);
and U4235 (N_4235,N_2561,N_2948);
nand U4236 (N_4236,N_2684,N_3279);
and U4237 (N_4237,N_2529,N_2748);
and U4238 (N_4238,N_3125,N_2773);
nor U4239 (N_4239,N_3740,N_3666);
and U4240 (N_4240,N_3539,N_3232);
nor U4241 (N_4241,N_3384,N_3457);
or U4242 (N_4242,N_2870,N_3398);
and U4243 (N_4243,N_3493,N_2907);
xor U4244 (N_4244,N_3717,N_2896);
nor U4245 (N_4245,N_3675,N_2778);
nand U4246 (N_4246,N_2792,N_2598);
nand U4247 (N_4247,N_2743,N_3454);
nor U4248 (N_4248,N_3513,N_3475);
nor U4249 (N_4249,N_2521,N_3182);
and U4250 (N_4250,N_3121,N_3015);
nor U4251 (N_4251,N_3567,N_3327);
and U4252 (N_4252,N_3130,N_3428);
nand U4253 (N_4253,N_3019,N_2805);
nor U4254 (N_4254,N_3681,N_2692);
or U4255 (N_4255,N_2573,N_3736);
nor U4256 (N_4256,N_3310,N_3122);
or U4257 (N_4257,N_3058,N_3236);
and U4258 (N_4258,N_3559,N_3353);
and U4259 (N_4259,N_2836,N_3534);
and U4260 (N_4260,N_2626,N_3540);
nor U4261 (N_4261,N_2575,N_3163);
and U4262 (N_4262,N_2698,N_3227);
and U4263 (N_4263,N_2564,N_2705);
xor U4264 (N_4264,N_2812,N_2960);
xnor U4265 (N_4265,N_3480,N_3726);
or U4266 (N_4266,N_2955,N_2985);
nand U4267 (N_4267,N_3744,N_3012);
nand U4268 (N_4268,N_3745,N_3523);
and U4269 (N_4269,N_3368,N_2912);
nor U4270 (N_4270,N_3157,N_3052);
or U4271 (N_4271,N_3432,N_3088);
and U4272 (N_4272,N_3154,N_2979);
xor U4273 (N_4273,N_2934,N_3615);
nor U4274 (N_4274,N_3296,N_2616);
and U4275 (N_4275,N_3042,N_3322);
nand U4276 (N_4276,N_2969,N_3485);
or U4277 (N_4277,N_2572,N_2943);
nor U4278 (N_4278,N_3528,N_2845);
nor U4279 (N_4279,N_2647,N_3650);
and U4280 (N_4280,N_3097,N_3522);
and U4281 (N_4281,N_3357,N_2557);
nand U4282 (N_4282,N_3007,N_3593);
or U4283 (N_4283,N_2968,N_2942);
nor U4284 (N_4284,N_3035,N_3474);
xor U4285 (N_4285,N_3439,N_3694);
nand U4286 (N_4286,N_3303,N_3732);
or U4287 (N_4287,N_3270,N_3526);
and U4288 (N_4288,N_3360,N_2687);
or U4289 (N_4289,N_3259,N_3611);
nor U4290 (N_4290,N_3617,N_3201);
nand U4291 (N_4291,N_2676,N_2662);
xor U4292 (N_4292,N_2940,N_3185);
or U4293 (N_4293,N_2824,N_3707);
nand U4294 (N_4294,N_3040,N_2958);
and U4295 (N_4295,N_3309,N_3578);
nand U4296 (N_4296,N_3536,N_3095);
nor U4297 (N_4297,N_2927,N_2593);
and U4298 (N_4298,N_2993,N_2842);
and U4299 (N_4299,N_3741,N_3355);
or U4300 (N_4300,N_3056,N_3301);
and U4301 (N_4301,N_3024,N_2918);
nor U4302 (N_4302,N_2899,N_3293);
nor U4303 (N_4303,N_3641,N_2587);
nand U4304 (N_4304,N_3423,N_2650);
nand U4305 (N_4305,N_3118,N_2784);
xor U4306 (N_4306,N_3636,N_3080);
and U4307 (N_4307,N_2640,N_3620);
or U4308 (N_4308,N_2891,N_3124);
or U4309 (N_4309,N_3336,N_2599);
xor U4310 (N_4310,N_2755,N_2534);
nor U4311 (N_4311,N_3356,N_3426);
xnor U4312 (N_4312,N_3319,N_3382);
nor U4313 (N_4313,N_3505,N_2568);
nor U4314 (N_4314,N_3208,N_3702);
nand U4315 (N_4315,N_3674,N_2578);
and U4316 (N_4316,N_3338,N_2826);
xnor U4317 (N_4317,N_3094,N_2719);
and U4318 (N_4318,N_3257,N_3374);
and U4319 (N_4319,N_3178,N_3299);
or U4320 (N_4320,N_2501,N_3218);
nor U4321 (N_4321,N_3067,N_3561);
nand U4322 (N_4322,N_2654,N_2559);
nor U4323 (N_4323,N_2660,N_2866);
nand U4324 (N_4324,N_3582,N_3070);
or U4325 (N_4325,N_2502,N_3049);
xor U4326 (N_4326,N_3397,N_3477);
xor U4327 (N_4327,N_3467,N_3639);
or U4328 (N_4328,N_2550,N_3487);
xor U4329 (N_4329,N_2804,N_3050);
nor U4330 (N_4330,N_3734,N_3542);
xor U4331 (N_4331,N_3714,N_3159);
xor U4332 (N_4332,N_3176,N_3419);
or U4333 (N_4333,N_3591,N_2790);
nor U4334 (N_4334,N_2524,N_2903);
and U4335 (N_4335,N_3077,N_2675);
xnor U4336 (N_4336,N_3197,N_3541);
nand U4337 (N_4337,N_2659,N_3048);
or U4338 (N_4338,N_2610,N_3743);
or U4339 (N_4339,N_2555,N_2644);
xnor U4340 (N_4340,N_3637,N_3228);
and U4341 (N_4341,N_2621,N_3669);
nand U4342 (N_4342,N_3051,N_3598);
or U4343 (N_4343,N_3684,N_2761);
xnor U4344 (N_4344,N_2767,N_2860);
nor U4345 (N_4345,N_3066,N_2902);
nand U4346 (N_4346,N_3191,N_2643);
or U4347 (N_4347,N_2797,N_2715);
and U4348 (N_4348,N_2799,N_2614);
and U4349 (N_4349,N_2520,N_2603);
or U4350 (N_4350,N_3444,N_3275);
nor U4351 (N_4351,N_2507,N_3417);
nand U4352 (N_4352,N_3630,N_3470);
and U4353 (N_4353,N_2886,N_3406);
nand U4354 (N_4354,N_2933,N_3231);
or U4355 (N_4355,N_3628,N_2619);
nor U4356 (N_4356,N_3343,N_3241);
or U4357 (N_4357,N_3672,N_3631);
or U4358 (N_4358,N_2951,N_3073);
xnor U4359 (N_4359,N_2574,N_2533);
xor U4360 (N_4360,N_3436,N_3494);
or U4361 (N_4361,N_3099,N_3394);
nand U4362 (N_4362,N_3583,N_2791);
nor U4363 (N_4363,N_2656,N_3020);
nand U4364 (N_4364,N_2702,N_2729);
xnor U4365 (N_4365,N_2850,N_3405);
and U4366 (N_4366,N_3151,N_3022);
nor U4367 (N_4367,N_2625,N_2526);
nor U4368 (N_4368,N_2972,N_2840);
and U4369 (N_4369,N_3027,N_3029);
or U4370 (N_4370,N_3063,N_2877);
nor U4371 (N_4371,N_3276,N_3273);
nor U4372 (N_4372,N_2754,N_2787);
nor U4373 (N_4373,N_3537,N_2653);
xnor U4374 (N_4374,N_3538,N_3700);
nand U4375 (N_4375,N_2548,N_2586);
nand U4376 (N_4376,N_3726,N_3387);
or U4377 (N_4377,N_2650,N_2597);
xnor U4378 (N_4378,N_3433,N_2619);
xnor U4379 (N_4379,N_3324,N_3673);
nor U4380 (N_4380,N_2852,N_2920);
or U4381 (N_4381,N_2790,N_3123);
nor U4382 (N_4382,N_3658,N_2899);
or U4383 (N_4383,N_2884,N_3668);
and U4384 (N_4384,N_2890,N_2856);
and U4385 (N_4385,N_2594,N_2916);
nand U4386 (N_4386,N_3411,N_3208);
nand U4387 (N_4387,N_3611,N_2961);
nand U4388 (N_4388,N_3140,N_3444);
and U4389 (N_4389,N_3533,N_2956);
nand U4390 (N_4390,N_3289,N_2704);
nand U4391 (N_4391,N_2703,N_3328);
and U4392 (N_4392,N_2654,N_3146);
xnor U4393 (N_4393,N_3638,N_3438);
xnor U4394 (N_4394,N_2899,N_3546);
or U4395 (N_4395,N_3653,N_3396);
nand U4396 (N_4396,N_3484,N_2781);
nor U4397 (N_4397,N_2687,N_3544);
or U4398 (N_4398,N_3283,N_3343);
or U4399 (N_4399,N_3033,N_3706);
nand U4400 (N_4400,N_3101,N_2957);
nor U4401 (N_4401,N_2697,N_3235);
nor U4402 (N_4402,N_2607,N_3125);
xnor U4403 (N_4403,N_3593,N_2848);
nor U4404 (N_4404,N_3018,N_3135);
nor U4405 (N_4405,N_2694,N_3681);
nand U4406 (N_4406,N_3127,N_2675);
nor U4407 (N_4407,N_2623,N_3524);
nor U4408 (N_4408,N_3056,N_2578);
and U4409 (N_4409,N_2968,N_2840);
xor U4410 (N_4410,N_2566,N_3367);
nor U4411 (N_4411,N_2911,N_3558);
nor U4412 (N_4412,N_3275,N_2922);
nand U4413 (N_4413,N_2952,N_3398);
nand U4414 (N_4414,N_3242,N_3511);
nand U4415 (N_4415,N_3138,N_3418);
or U4416 (N_4416,N_3246,N_2762);
xor U4417 (N_4417,N_3490,N_2912);
and U4418 (N_4418,N_3590,N_3567);
nand U4419 (N_4419,N_2628,N_2500);
or U4420 (N_4420,N_2779,N_3083);
xor U4421 (N_4421,N_3698,N_3737);
xnor U4422 (N_4422,N_2876,N_2938);
nand U4423 (N_4423,N_3287,N_3719);
nand U4424 (N_4424,N_2938,N_2581);
or U4425 (N_4425,N_2950,N_3672);
and U4426 (N_4426,N_3325,N_3534);
or U4427 (N_4427,N_2523,N_3387);
or U4428 (N_4428,N_2882,N_3124);
and U4429 (N_4429,N_3431,N_2744);
and U4430 (N_4430,N_2876,N_2516);
nor U4431 (N_4431,N_2737,N_2769);
xnor U4432 (N_4432,N_3583,N_3603);
xor U4433 (N_4433,N_3495,N_3465);
or U4434 (N_4434,N_2708,N_3472);
or U4435 (N_4435,N_3503,N_3355);
nor U4436 (N_4436,N_2793,N_3458);
and U4437 (N_4437,N_2557,N_3484);
nor U4438 (N_4438,N_3196,N_2557);
and U4439 (N_4439,N_2820,N_3487);
nor U4440 (N_4440,N_3372,N_3613);
and U4441 (N_4441,N_2710,N_2989);
or U4442 (N_4442,N_2942,N_2851);
or U4443 (N_4443,N_2785,N_3724);
xnor U4444 (N_4444,N_2538,N_3313);
or U4445 (N_4445,N_3552,N_3182);
and U4446 (N_4446,N_3476,N_3674);
nand U4447 (N_4447,N_3458,N_3064);
and U4448 (N_4448,N_3533,N_2863);
and U4449 (N_4449,N_3405,N_2678);
nand U4450 (N_4450,N_3317,N_2653);
or U4451 (N_4451,N_3324,N_3027);
nor U4452 (N_4452,N_3046,N_2583);
nor U4453 (N_4453,N_3155,N_2515);
xor U4454 (N_4454,N_3190,N_3563);
nand U4455 (N_4455,N_3435,N_3388);
or U4456 (N_4456,N_3445,N_2651);
nand U4457 (N_4457,N_2854,N_2657);
xor U4458 (N_4458,N_2802,N_3141);
nand U4459 (N_4459,N_3674,N_2890);
nand U4460 (N_4460,N_3316,N_3481);
or U4461 (N_4461,N_3077,N_3040);
and U4462 (N_4462,N_3407,N_2839);
nand U4463 (N_4463,N_3069,N_3339);
xor U4464 (N_4464,N_3173,N_3197);
nor U4465 (N_4465,N_2989,N_3155);
and U4466 (N_4466,N_3526,N_3532);
and U4467 (N_4467,N_3658,N_3588);
or U4468 (N_4468,N_2579,N_2954);
nor U4469 (N_4469,N_3177,N_3141);
xnor U4470 (N_4470,N_3114,N_2781);
or U4471 (N_4471,N_3005,N_2515);
or U4472 (N_4472,N_2724,N_3717);
nand U4473 (N_4473,N_3148,N_3296);
xnor U4474 (N_4474,N_3541,N_3241);
xnor U4475 (N_4475,N_2796,N_2564);
and U4476 (N_4476,N_3047,N_3534);
xor U4477 (N_4477,N_2774,N_3216);
or U4478 (N_4478,N_2893,N_3346);
nand U4479 (N_4479,N_2560,N_3628);
nor U4480 (N_4480,N_3457,N_3541);
nor U4481 (N_4481,N_3353,N_3129);
nor U4482 (N_4482,N_2630,N_2672);
and U4483 (N_4483,N_3215,N_3445);
xnor U4484 (N_4484,N_3447,N_2586);
or U4485 (N_4485,N_2747,N_3474);
or U4486 (N_4486,N_2984,N_3704);
and U4487 (N_4487,N_3432,N_2791);
or U4488 (N_4488,N_2704,N_3431);
or U4489 (N_4489,N_3092,N_3051);
and U4490 (N_4490,N_3060,N_2897);
nand U4491 (N_4491,N_2979,N_2745);
nand U4492 (N_4492,N_3402,N_3187);
nor U4493 (N_4493,N_3524,N_3316);
or U4494 (N_4494,N_2523,N_3480);
nor U4495 (N_4495,N_2962,N_3123);
nand U4496 (N_4496,N_3596,N_2585);
nor U4497 (N_4497,N_2624,N_3477);
xor U4498 (N_4498,N_2971,N_2817);
nor U4499 (N_4499,N_3498,N_2763);
or U4500 (N_4500,N_3602,N_2712);
or U4501 (N_4501,N_2747,N_2674);
nand U4502 (N_4502,N_2873,N_3036);
and U4503 (N_4503,N_2660,N_2704);
nand U4504 (N_4504,N_3297,N_3560);
and U4505 (N_4505,N_3541,N_2704);
xor U4506 (N_4506,N_2585,N_2669);
xor U4507 (N_4507,N_2926,N_3680);
nor U4508 (N_4508,N_2879,N_3497);
and U4509 (N_4509,N_3483,N_2509);
or U4510 (N_4510,N_2721,N_3695);
xor U4511 (N_4511,N_2779,N_3139);
and U4512 (N_4512,N_2619,N_3672);
nand U4513 (N_4513,N_3373,N_3348);
xor U4514 (N_4514,N_2785,N_2636);
nor U4515 (N_4515,N_3225,N_3174);
and U4516 (N_4516,N_3195,N_2654);
xor U4517 (N_4517,N_3315,N_3468);
nand U4518 (N_4518,N_3273,N_3346);
xor U4519 (N_4519,N_3305,N_3282);
nor U4520 (N_4520,N_3149,N_3553);
nand U4521 (N_4521,N_2996,N_2507);
nor U4522 (N_4522,N_3094,N_2865);
nor U4523 (N_4523,N_3707,N_2636);
or U4524 (N_4524,N_3265,N_3186);
nand U4525 (N_4525,N_2578,N_3644);
nand U4526 (N_4526,N_3400,N_2767);
and U4527 (N_4527,N_2988,N_2505);
nor U4528 (N_4528,N_3515,N_3357);
and U4529 (N_4529,N_3570,N_2629);
nand U4530 (N_4530,N_2957,N_3376);
and U4531 (N_4531,N_3216,N_3115);
and U4532 (N_4532,N_2650,N_2529);
or U4533 (N_4533,N_2890,N_3052);
xnor U4534 (N_4534,N_2889,N_3371);
nor U4535 (N_4535,N_2864,N_2706);
or U4536 (N_4536,N_3619,N_2840);
and U4537 (N_4537,N_2583,N_3051);
xor U4538 (N_4538,N_2708,N_3423);
nand U4539 (N_4539,N_3100,N_3299);
nor U4540 (N_4540,N_2885,N_2833);
and U4541 (N_4541,N_2926,N_3384);
and U4542 (N_4542,N_3441,N_3316);
nand U4543 (N_4543,N_2520,N_3302);
or U4544 (N_4544,N_3170,N_3042);
and U4545 (N_4545,N_2731,N_2804);
xor U4546 (N_4546,N_3610,N_3571);
xor U4547 (N_4547,N_3240,N_2650);
nor U4548 (N_4548,N_3513,N_2557);
nand U4549 (N_4549,N_3326,N_3354);
nor U4550 (N_4550,N_2901,N_2662);
and U4551 (N_4551,N_3708,N_2739);
nand U4552 (N_4552,N_3157,N_3183);
or U4553 (N_4553,N_3619,N_2756);
xnor U4554 (N_4554,N_3727,N_3055);
nor U4555 (N_4555,N_2692,N_3288);
and U4556 (N_4556,N_2613,N_2615);
nand U4557 (N_4557,N_3695,N_2532);
xnor U4558 (N_4558,N_2666,N_3664);
xnor U4559 (N_4559,N_2654,N_2537);
or U4560 (N_4560,N_2528,N_3034);
nor U4561 (N_4561,N_2782,N_2607);
xor U4562 (N_4562,N_3404,N_2524);
nand U4563 (N_4563,N_2523,N_3178);
nand U4564 (N_4564,N_3047,N_3275);
or U4565 (N_4565,N_2592,N_3642);
or U4566 (N_4566,N_3051,N_2636);
or U4567 (N_4567,N_3049,N_2533);
or U4568 (N_4568,N_3612,N_3726);
and U4569 (N_4569,N_3202,N_3013);
or U4570 (N_4570,N_3483,N_3054);
xnor U4571 (N_4571,N_3449,N_2511);
and U4572 (N_4572,N_2642,N_3297);
and U4573 (N_4573,N_3710,N_3315);
and U4574 (N_4574,N_3128,N_3525);
and U4575 (N_4575,N_3736,N_2512);
or U4576 (N_4576,N_3487,N_3645);
and U4577 (N_4577,N_3645,N_2926);
or U4578 (N_4578,N_3268,N_3397);
nand U4579 (N_4579,N_3166,N_3237);
nor U4580 (N_4580,N_3608,N_2642);
and U4581 (N_4581,N_3559,N_2544);
or U4582 (N_4582,N_2959,N_3743);
nand U4583 (N_4583,N_2724,N_3671);
nor U4584 (N_4584,N_3598,N_2773);
xor U4585 (N_4585,N_2991,N_3438);
nand U4586 (N_4586,N_2711,N_3239);
and U4587 (N_4587,N_3420,N_2919);
nand U4588 (N_4588,N_2654,N_3008);
and U4589 (N_4589,N_3188,N_2628);
nand U4590 (N_4590,N_3219,N_3350);
or U4591 (N_4591,N_3662,N_3635);
nor U4592 (N_4592,N_2999,N_3299);
and U4593 (N_4593,N_3544,N_2528);
nand U4594 (N_4594,N_3728,N_2639);
nor U4595 (N_4595,N_2634,N_2502);
nand U4596 (N_4596,N_2552,N_3354);
and U4597 (N_4597,N_2569,N_3364);
and U4598 (N_4598,N_3524,N_3562);
xor U4599 (N_4599,N_2979,N_3538);
and U4600 (N_4600,N_2745,N_3693);
and U4601 (N_4601,N_2586,N_3022);
xor U4602 (N_4602,N_3444,N_2792);
nand U4603 (N_4603,N_3013,N_2768);
xor U4604 (N_4604,N_3019,N_2786);
nor U4605 (N_4605,N_3583,N_3482);
nor U4606 (N_4606,N_3180,N_3474);
xnor U4607 (N_4607,N_3168,N_2719);
nand U4608 (N_4608,N_3398,N_3179);
and U4609 (N_4609,N_3211,N_2762);
and U4610 (N_4610,N_2923,N_3212);
nand U4611 (N_4611,N_2796,N_3244);
nand U4612 (N_4612,N_3534,N_2742);
and U4613 (N_4613,N_3331,N_2740);
and U4614 (N_4614,N_2665,N_2841);
nand U4615 (N_4615,N_2920,N_2619);
and U4616 (N_4616,N_2745,N_3553);
nor U4617 (N_4617,N_2622,N_2636);
and U4618 (N_4618,N_3345,N_2851);
or U4619 (N_4619,N_3349,N_3071);
nor U4620 (N_4620,N_2839,N_3639);
nor U4621 (N_4621,N_3592,N_2715);
xor U4622 (N_4622,N_3006,N_2594);
xnor U4623 (N_4623,N_2684,N_3543);
nor U4624 (N_4624,N_2587,N_3602);
xor U4625 (N_4625,N_3707,N_3463);
and U4626 (N_4626,N_3565,N_2867);
nand U4627 (N_4627,N_3491,N_3089);
xor U4628 (N_4628,N_3354,N_2751);
nand U4629 (N_4629,N_2873,N_3105);
or U4630 (N_4630,N_3194,N_3100);
nand U4631 (N_4631,N_2703,N_3319);
and U4632 (N_4632,N_3386,N_3286);
and U4633 (N_4633,N_3610,N_3229);
nor U4634 (N_4634,N_3473,N_3449);
nand U4635 (N_4635,N_2523,N_3112);
or U4636 (N_4636,N_3353,N_2574);
nand U4637 (N_4637,N_3050,N_2896);
xor U4638 (N_4638,N_3022,N_3591);
or U4639 (N_4639,N_3043,N_3194);
and U4640 (N_4640,N_2624,N_3434);
or U4641 (N_4641,N_2631,N_2754);
nand U4642 (N_4642,N_3488,N_3329);
and U4643 (N_4643,N_3252,N_3010);
and U4644 (N_4644,N_3097,N_3055);
nor U4645 (N_4645,N_2617,N_2629);
nand U4646 (N_4646,N_3622,N_2926);
nand U4647 (N_4647,N_2980,N_3179);
or U4648 (N_4648,N_2665,N_2722);
or U4649 (N_4649,N_3443,N_2715);
nand U4650 (N_4650,N_3267,N_3088);
nor U4651 (N_4651,N_2845,N_3674);
or U4652 (N_4652,N_2885,N_3257);
or U4653 (N_4653,N_2613,N_2544);
and U4654 (N_4654,N_3429,N_2518);
and U4655 (N_4655,N_2510,N_2541);
or U4656 (N_4656,N_3474,N_2655);
xnor U4657 (N_4657,N_2727,N_3129);
xor U4658 (N_4658,N_2595,N_3105);
nand U4659 (N_4659,N_3186,N_2942);
or U4660 (N_4660,N_3036,N_3663);
and U4661 (N_4661,N_3545,N_2907);
or U4662 (N_4662,N_2515,N_3719);
nor U4663 (N_4663,N_3265,N_3029);
xor U4664 (N_4664,N_3128,N_3184);
nor U4665 (N_4665,N_2527,N_2712);
nand U4666 (N_4666,N_3053,N_2870);
xnor U4667 (N_4667,N_2601,N_3073);
xnor U4668 (N_4668,N_3395,N_3423);
and U4669 (N_4669,N_3013,N_2877);
nor U4670 (N_4670,N_2728,N_2727);
xor U4671 (N_4671,N_2817,N_3442);
or U4672 (N_4672,N_2874,N_3651);
nand U4673 (N_4673,N_2797,N_3567);
xor U4674 (N_4674,N_3360,N_2911);
nor U4675 (N_4675,N_2519,N_2637);
or U4676 (N_4676,N_3019,N_2942);
and U4677 (N_4677,N_2901,N_2802);
nor U4678 (N_4678,N_3590,N_3108);
nor U4679 (N_4679,N_2617,N_2581);
or U4680 (N_4680,N_3383,N_3122);
xor U4681 (N_4681,N_2919,N_2592);
or U4682 (N_4682,N_2813,N_2814);
nor U4683 (N_4683,N_2938,N_2930);
xnor U4684 (N_4684,N_3498,N_3280);
nand U4685 (N_4685,N_2785,N_3295);
nor U4686 (N_4686,N_3409,N_2983);
and U4687 (N_4687,N_2679,N_3293);
and U4688 (N_4688,N_2885,N_2917);
and U4689 (N_4689,N_2702,N_3585);
xor U4690 (N_4690,N_3049,N_2601);
xor U4691 (N_4691,N_3159,N_3665);
and U4692 (N_4692,N_3466,N_2607);
nor U4693 (N_4693,N_2569,N_2604);
and U4694 (N_4694,N_3428,N_2759);
and U4695 (N_4695,N_3280,N_2631);
and U4696 (N_4696,N_3251,N_2674);
and U4697 (N_4697,N_2950,N_2538);
or U4698 (N_4698,N_2734,N_3215);
and U4699 (N_4699,N_2811,N_2524);
nand U4700 (N_4700,N_3117,N_3404);
or U4701 (N_4701,N_2703,N_2679);
xnor U4702 (N_4702,N_3296,N_3470);
xor U4703 (N_4703,N_3497,N_2997);
or U4704 (N_4704,N_2966,N_2569);
or U4705 (N_4705,N_3095,N_3628);
nor U4706 (N_4706,N_3641,N_2945);
and U4707 (N_4707,N_3050,N_3580);
nor U4708 (N_4708,N_3671,N_2745);
xnor U4709 (N_4709,N_3234,N_3506);
xnor U4710 (N_4710,N_3210,N_3696);
xnor U4711 (N_4711,N_2964,N_3112);
nor U4712 (N_4712,N_3346,N_3113);
xor U4713 (N_4713,N_3365,N_3376);
nand U4714 (N_4714,N_3320,N_3145);
nor U4715 (N_4715,N_3348,N_2549);
and U4716 (N_4716,N_3111,N_2793);
and U4717 (N_4717,N_3712,N_3171);
nand U4718 (N_4718,N_3694,N_2616);
nand U4719 (N_4719,N_3686,N_2951);
nor U4720 (N_4720,N_2942,N_3037);
xnor U4721 (N_4721,N_3428,N_2980);
xor U4722 (N_4722,N_2984,N_2530);
nor U4723 (N_4723,N_2690,N_2543);
xnor U4724 (N_4724,N_2537,N_3070);
nor U4725 (N_4725,N_2662,N_3109);
xnor U4726 (N_4726,N_3393,N_2934);
nand U4727 (N_4727,N_3009,N_3137);
xor U4728 (N_4728,N_2538,N_2741);
nor U4729 (N_4729,N_3565,N_2624);
or U4730 (N_4730,N_2667,N_2652);
nor U4731 (N_4731,N_3231,N_3463);
xnor U4732 (N_4732,N_3664,N_3694);
and U4733 (N_4733,N_3738,N_3242);
or U4734 (N_4734,N_3017,N_2670);
nor U4735 (N_4735,N_3736,N_2940);
xnor U4736 (N_4736,N_2501,N_2769);
and U4737 (N_4737,N_3227,N_3105);
xor U4738 (N_4738,N_3443,N_2547);
and U4739 (N_4739,N_3741,N_3082);
and U4740 (N_4740,N_3028,N_2517);
or U4741 (N_4741,N_3532,N_3582);
nand U4742 (N_4742,N_2857,N_3460);
xor U4743 (N_4743,N_2972,N_2548);
or U4744 (N_4744,N_3501,N_3565);
and U4745 (N_4745,N_3020,N_3536);
and U4746 (N_4746,N_3689,N_3306);
xnor U4747 (N_4747,N_3319,N_3682);
xor U4748 (N_4748,N_2665,N_3023);
nor U4749 (N_4749,N_3232,N_2787);
nand U4750 (N_4750,N_3741,N_2730);
nor U4751 (N_4751,N_3714,N_3181);
and U4752 (N_4752,N_2849,N_3303);
and U4753 (N_4753,N_3304,N_3180);
or U4754 (N_4754,N_3062,N_3454);
xnor U4755 (N_4755,N_3205,N_3437);
or U4756 (N_4756,N_3362,N_2889);
nand U4757 (N_4757,N_3005,N_2902);
or U4758 (N_4758,N_2805,N_3200);
nand U4759 (N_4759,N_2686,N_2524);
xnor U4760 (N_4760,N_2907,N_2592);
or U4761 (N_4761,N_3464,N_2938);
nor U4762 (N_4762,N_3561,N_3483);
and U4763 (N_4763,N_2690,N_2749);
or U4764 (N_4764,N_3441,N_3061);
or U4765 (N_4765,N_2767,N_2600);
nor U4766 (N_4766,N_2517,N_3313);
xor U4767 (N_4767,N_3008,N_3502);
or U4768 (N_4768,N_3462,N_2846);
nor U4769 (N_4769,N_2654,N_3119);
nor U4770 (N_4770,N_3298,N_2829);
or U4771 (N_4771,N_3723,N_2970);
or U4772 (N_4772,N_2976,N_2995);
nor U4773 (N_4773,N_2923,N_3074);
xnor U4774 (N_4774,N_2881,N_3440);
or U4775 (N_4775,N_3265,N_2820);
nor U4776 (N_4776,N_2853,N_3144);
and U4777 (N_4777,N_2862,N_2934);
nor U4778 (N_4778,N_2625,N_3007);
and U4779 (N_4779,N_3258,N_3097);
or U4780 (N_4780,N_2550,N_3008);
nand U4781 (N_4781,N_2843,N_2675);
nand U4782 (N_4782,N_2833,N_3061);
or U4783 (N_4783,N_2570,N_3075);
nor U4784 (N_4784,N_3205,N_3518);
xor U4785 (N_4785,N_3414,N_3352);
xnor U4786 (N_4786,N_3486,N_3004);
nand U4787 (N_4787,N_2505,N_3042);
and U4788 (N_4788,N_3090,N_3437);
xor U4789 (N_4789,N_3702,N_3115);
nor U4790 (N_4790,N_3683,N_2619);
nor U4791 (N_4791,N_2603,N_3101);
xnor U4792 (N_4792,N_2634,N_3401);
nand U4793 (N_4793,N_3479,N_3376);
nor U4794 (N_4794,N_2932,N_3527);
xor U4795 (N_4795,N_2570,N_2648);
or U4796 (N_4796,N_2787,N_2589);
or U4797 (N_4797,N_3513,N_2772);
xnor U4798 (N_4798,N_2809,N_3051);
and U4799 (N_4799,N_3437,N_2624);
and U4800 (N_4800,N_3728,N_2971);
nand U4801 (N_4801,N_2909,N_3354);
and U4802 (N_4802,N_3374,N_3716);
xor U4803 (N_4803,N_3607,N_2858);
and U4804 (N_4804,N_2764,N_2631);
or U4805 (N_4805,N_2628,N_3574);
or U4806 (N_4806,N_3165,N_2945);
nor U4807 (N_4807,N_2653,N_3568);
nand U4808 (N_4808,N_3052,N_3715);
or U4809 (N_4809,N_2685,N_2813);
and U4810 (N_4810,N_3152,N_2979);
xor U4811 (N_4811,N_3019,N_3491);
xnor U4812 (N_4812,N_2761,N_3694);
or U4813 (N_4813,N_3308,N_2693);
nand U4814 (N_4814,N_3156,N_2600);
nor U4815 (N_4815,N_3712,N_3100);
xnor U4816 (N_4816,N_3686,N_2832);
nand U4817 (N_4817,N_3744,N_2639);
or U4818 (N_4818,N_3564,N_3712);
nor U4819 (N_4819,N_2934,N_2760);
or U4820 (N_4820,N_3259,N_3024);
nor U4821 (N_4821,N_3544,N_3527);
nor U4822 (N_4822,N_2854,N_2837);
nand U4823 (N_4823,N_3214,N_3604);
or U4824 (N_4824,N_2733,N_2764);
or U4825 (N_4825,N_2518,N_2517);
or U4826 (N_4826,N_3255,N_3491);
nand U4827 (N_4827,N_2997,N_3262);
nor U4828 (N_4828,N_3316,N_2991);
nor U4829 (N_4829,N_3644,N_2528);
nor U4830 (N_4830,N_3053,N_2630);
xor U4831 (N_4831,N_3453,N_3496);
xnor U4832 (N_4832,N_3170,N_2904);
and U4833 (N_4833,N_3060,N_3149);
nand U4834 (N_4834,N_3457,N_2679);
nand U4835 (N_4835,N_3109,N_3514);
nor U4836 (N_4836,N_2583,N_3268);
xor U4837 (N_4837,N_2914,N_2858);
and U4838 (N_4838,N_3035,N_2944);
and U4839 (N_4839,N_3073,N_2582);
xnor U4840 (N_4840,N_3607,N_3066);
and U4841 (N_4841,N_2648,N_3123);
and U4842 (N_4842,N_2558,N_2586);
or U4843 (N_4843,N_2605,N_3134);
and U4844 (N_4844,N_3648,N_2940);
or U4845 (N_4845,N_3048,N_2561);
nor U4846 (N_4846,N_3325,N_2506);
nand U4847 (N_4847,N_3666,N_2566);
nand U4848 (N_4848,N_3112,N_3318);
xor U4849 (N_4849,N_2914,N_3090);
nand U4850 (N_4850,N_2709,N_2666);
and U4851 (N_4851,N_3485,N_3412);
nor U4852 (N_4852,N_3623,N_3178);
and U4853 (N_4853,N_2738,N_2605);
and U4854 (N_4854,N_2657,N_3063);
and U4855 (N_4855,N_3102,N_3694);
xnor U4856 (N_4856,N_2598,N_3043);
or U4857 (N_4857,N_2892,N_2954);
or U4858 (N_4858,N_2826,N_3086);
xnor U4859 (N_4859,N_2855,N_3334);
nand U4860 (N_4860,N_3514,N_2782);
xor U4861 (N_4861,N_3111,N_3021);
or U4862 (N_4862,N_2955,N_2751);
and U4863 (N_4863,N_2649,N_3192);
or U4864 (N_4864,N_3702,N_2578);
and U4865 (N_4865,N_3554,N_2667);
or U4866 (N_4866,N_3262,N_3424);
xnor U4867 (N_4867,N_3495,N_3267);
xor U4868 (N_4868,N_2910,N_3330);
or U4869 (N_4869,N_2695,N_2588);
xor U4870 (N_4870,N_2749,N_2698);
nor U4871 (N_4871,N_3285,N_3367);
or U4872 (N_4872,N_3009,N_3236);
and U4873 (N_4873,N_2583,N_3378);
nor U4874 (N_4874,N_3159,N_3673);
nand U4875 (N_4875,N_3606,N_2529);
nand U4876 (N_4876,N_3387,N_3298);
or U4877 (N_4877,N_2667,N_3352);
nand U4878 (N_4878,N_2504,N_3080);
nor U4879 (N_4879,N_3686,N_2563);
nand U4880 (N_4880,N_2551,N_3196);
xor U4881 (N_4881,N_3308,N_3481);
nor U4882 (N_4882,N_2802,N_2544);
nand U4883 (N_4883,N_2816,N_3385);
and U4884 (N_4884,N_2963,N_3363);
xor U4885 (N_4885,N_2551,N_3463);
xor U4886 (N_4886,N_3591,N_3414);
nand U4887 (N_4887,N_3012,N_3141);
and U4888 (N_4888,N_3133,N_2803);
xnor U4889 (N_4889,N_3322,N_2803);
nor U4890 (N_4890,N_2964,N_3099);
nor U4891 (N_4891,N_3237,N_3114);
or U4892 (N_4892,N_3453,N_2913);
and U4893 (N_4893,N_3116,N_3435);
and U4894 (N_4894,N_2569,N_2626);
and U4895 (N_4895,N_3434,N_3057);
xor U4896 (N_4896,N_3656,N_3696);
nand U4897 (N_4897,N_2900,N_3216);
xnor U4898 (N_4898,N_3372,N_3441);
nor U4899 (N_4899,N_3634,N_2537);
nor U4900 (N_4900,N_2890,N_3578);
xor U4901 (N_4901,N_3253,N_3118);
or U4902 (N_4902,N_3677,N_3329);
or U4903 (N_4903,N_2707,N_2608);
or U4904 (N_4904,N_3109,N_3486);
and U4905 (N_4905,N_3512,N_3748);
nand U4906 (N_4906,N_3734,N_3160);
and U4907 (N_4907,N_3736,N_3565);
or U4908 (N_4908,N_3094,N_3277);
xnor U4909 (N_4909,N_3138,N_3451);
nand U4910 (N_4910,N_3304,N_3271);
and U4911 (N_4911,N_3096,N_3651);
xnor U4912 (N_4912,N_3510,N_2855);
nor U4913 (N_4913,N_3231,N_2511);
and U4914 (N_4914,N_3052,N_3472);
and U4915 (N_4915,N_3746,N_3061);
and U4916 (N_4916,N_3303,N_2834);
and U4917 (N_4917,N_3722,N_2927);
nand U4918 (N_4918,N_2846,N_2864);
nand U4919 (N_4919,N_3070,N_3242);
nand U4920 (N_4920,N_3445,N_3287);
nor U4921 (N_4921,N_3239,N_3389);
xor U4922 (N_4922,N_2604,N_3563);
nor U4923 (N_4923,N_3747,N_3232);
xor U4924 (N_4924,N_2551,N_2697);
nor U4925 (N_4925,N_3033,N_3420);
nand U4926 (N_4926,N_3520,N_3527);
nand U4927 (N_4927,N_3537,N_3348);
or U4928 (N_4928,N_2614,N_3127);
nor U4929 (N_4929,N_2673,N_2706);
and U4930 (N_4930,N_2597,N_3393);
nor U4931 (N_4931,N_3415,N_3529);
and U4932 (N_4932,N_2870,N_2537);
xnor U4933 (N_4933,N_3140,N_3537);
xnor U4934 (N_4934,N_3513,N_3540);
nor U4935 (N_4935,N_2529,N_2592);
nor U4936 (N_4936,N_2601,N_2924);
or U4937 (N_4937,N_3673,N_3189);
nand U4938 (N_4938,N_3198,N_3326);
or U4939 (N_4939,N_3336,N_3215);
and U4940 (N_4940,N_3114,N_3406);
xor U4941 (N_4941,N_3335,N_3647);
or U4942 (N_4942,N_2975,N_3178);
xnor U4943 (N_4943,N_3085,N_3178);
xor U4944 (N_4944,N_2984,N_3267);
nand U4945 (N_4945,N_2706,N_3721);
or U4946 (N_4946,N_2679,N_3690);
or U4947 (N_4947,N_3665,N_3488);
and U4948 (N_4948,N_2604,N_3214);
nor U4949 (N_4949,N_3052,N_2775);
and U4950 (N_4950,N_2847,N_3481);
xnor U4951 (N_4951,N_2742,N_3156);
and U4952 (N_4952,N_2601,N_3601);
nand U4953 (N_4953,N_2832,N_2740);
nand U4954 (N_4954,N_3028,N_3009);
and U4955 (N_4955,N_3161,N_3297);
and U4956 (N_4956,N_3538,N_3158);
nor U4957 (N_4957,N_2696,N_2874);
nor U4958 (N_4958,N_2647,N_3695);
xnor U4959 (N_4959,N_3126,N_3485);
nor U4960 (N_4960,N_2986,N_2756);
xor U4961 (N_4961,N_2691,N_2899);
xnor U4962 (N_4962,N_3690,N_3270);
and U4963 (N_4963,N_3081,N_3171);
or U4964 (N_4964,N_2827,N_3180);
nand U4965 (N_4965,N_2988,N_3173);
nand U4966 (N_4966,N_2832,N_2700);
xnor U4967 (N_4967,N_2890,N_2941);
xnor U4968 (N_4968,N_3156,N_2835);
xor U4969 (N_4969,N_2997,N_3441);
or U4970 (N_4970,N_3644,N_3283);
xor U4971 (N_4971,N_3738,N_3723);
nand U4972 (N_4972,N_3638,N_3258);
nor U4973 (N_4973,N_2561,N_2563);
and U4974 (N_4974,N_2712,N_3089);
nand U4975 (N_4975,N_3602,N_2580);
xnor U4976 (N_4976,N_2788,N_2632);
nand U4977 (N_4977,N_3323,N_2889);
nor U4978 (N_4978,N_3523,N_2636);
and U4979 (N_4979,N_2715,N_3422);
and U4980 (N_4980,N_3658,N_3365);
and U4981 (N_4981,N_2876,N_3535);
xor U4982 (N_4982,N_2723,N_3042);
nor U4983 (N_4983,N_2885,N_3303);
nand U4984 (N_4984,N_2682,N_3663);
nor U4985 (N_4985,N_3095,N_3358);
xor U4986 (N_4986,N_3470,N_3139);
and U4987 (N_4987,N_2685,N_3010);
or U4988 (N_4988,N_3283,N_2841);
xnor U4989 (N_4989,N_2870,N_2676);
nand U4990 (N_4990,N_3210,N_3019);
or U4991 (N_4991,N_3635,N_3741);
and U4992 (N_4992,N_2777,N_3173);
xnor U4993 (N_4993,N_3551,N_3237);
nand U4994 (N_4994,N_2850,N_2742);
and U4995 (N_4995,N_2778,N_3007);
or U4996 (N_4996,N_2644,N_3296);
or U4997 (N_4997,N_2701,N_2976);
or U4998 (N_4998,N_2533,N_2626);
nor U4999 (N_4999,N_2944,N_3219);
nand U5000 (N_5000,N_4226,N_4499);
xor U5001 (N_5001,N_3958,N_4215);
nor U5002 (N_5002,N_3770,N_4726);
and U5003 (N_5003,N_4189,N_4936);
and U5004 (N_5004,N_4692,N_3843);
or U5005 (N_5005,N_4086,N_4573);
and U5006 (N_5006,N_3993,N_4797);
nor U5007 (N_5007,N_4221,N_3754);
and U5008 (N_5008,N_4230,N_4701);
xnor U5009 (N_5009,N_4591,N_4103);
or U5010 (N_5010,N_4392,N_4153);
nand U5011 (N_5011,N_4930,N_4382);
xnor U5012 (N_5012,N_4229,N_4580);
and U5013 (N_5013,N_4436,N_4245);
or U5014 (N_5014,N_4719,N_4916);
xor U5015 (N_5015,N_4061,N_4073);
and U5016 (N_5016,N_4234,N_4879);
or U5017 (N_5017,N_4020,N_4462);
nand U5018 (N_5018,N_4022,N_3886);
or U5019 (N_5019,N_4278,N_4492);
xnor U5020 (N_5020,N_4568,N_3762);
nand U5021 (N_5021,N_4708,N_3774);
nand U5022 (N_5022,N_4470,N_3920);
xor U5023 (N_5023,N_4270,N_4503);
nor U5024 (N_5024,N_4748,N_3827);
nor U5025 (N_5025,N_4199,N_3907);
or U5026 (N_5026,N_4364,N_3941);
and U5027 (N_5027,N_4794,N_4267);
nand U5028 (N_5028,N_4063,N_4722);
xnor U5029 (N_5029,N_4046,N_3985);
or U5030 (N_5030,N_4228,N_4256);
and U5031 (N_5031,N_3847,N_4030);
nand U5032 (N_5032,N_4912,N_4539);
nor U5033 (N_5033,N_4292,N_4995);
and U5034 (N_5034,N_4316,N_4097);
or U5035 (N_5035,N_3942,N_4579);
nor U5036 (N_5036,N_3905,N_4000);
nand U5037 (N_5037,N_4965,N_4446);
and U5038 (N_5038,N_4924,N_4831);
nor U5039 (N_5039,N_4166,N_4901);
nor U5040 (N_5040,N_4812,N_4322);
xor U5041 (N_5041,N_3791,N_4062);
or U5042 (N_5042,N_4069,N_3910);
nand U5043 (N_5043,N_4172,N_4272);
nor U5044 (N_5044,N_4639,N_4110);
nor U5045 (N_5045,N_4369,N_4979);
nor U5046 (N_5046,N_4567,N_3798);
xnor U5047 (N_5047,N_4452,N_4982);
and U5048 (N_5048,N_4635,N_4105);
or U5049 (N_5049,N_3950,N_4188);
or U5050 (N_5050,N_3819,N_3927);
or U5051 (N_5051,N_4331,N_4059);
nor U5052 (N_5052,N_4755,N_4949);
or U5053 (N_5053,N_3975,N_4140);
and U5054 (N_5054,N_4301,N_4420);
nand U5055 (N_5055,N_4574,N_4943);
nand U5056 (N_5056,N_4606,N_4888);
and U5057 (N_5057,N_4792,N_4804);
nor U5058 (N_5058,N_4422,N_4183);
and U5059 (N_5059,N_4225,N_4866);
nand U5060 (N_5060,N_4773,N_4564);
or U5061 (N_5061,N_4762,N_3872);
xor U5062 (N_5062,N_4808,N_4674);
or U5063 (N_5063,N_4088,N_4058);
xnor U5064 (N_5064,N_4175,N_3790);
nand U5065 (N_5065,N_4132,N_3814);
nand U5066 (N_5066,N_4513,N_4233);
xor U5067 (N_5067,N_3919,N_4501);
nor U5068 (N_5068,N_4625,N_4778);
nand U5069 (N_5069,N_4959,N_4883);
or U5070 (N_5070,N_4992,N_4456);
xnor U5071 (N_5071,N_4377,N_3932);
and U5072 (N_5072,N_4896,N_4727);
nand U5073 (N_5073,N_3994,N_4145);
xnor U5074 (N_5074,N_3881,N_4401);
and U5075 (N_5075,N_4307,N_4554);
or U5076 (N_5076,N_4205,N_4344);
xnor U5077 (N_5077,N_3971,N_3787);
xnor U5078 (N_5078,N_3831,N_4569);
nor U5079 (N_5079,N_3880,N_4351);
xor U5080 (N_5080,N_4889,N_4317);
and U5081 (N_5081,N_4908,N_4682);
and U5082 (N_5082,N_4438,N_4133);
and U5083 (N_5083,N_3828,N_4330);
or U5084 (N_5084,N_4024,N_4483);
and U5085 (N_5085,N_4581,N_3989);
and U5086 (N_5086,N_4620,N_4867);
nand U5087 (N_5087,N_4282,N_4614);
or U5088 (N_5088,N_4083,N_4884);
nor U5089 (N_5089,N_4303,N_4193);
xnor U5090 (N_5090,N_3865,N_3758);
and U5091 (N_5091,N_4666,N_4336);
nor U5092 (N_5092,N_4841,N_4589);
nand U5093 (N_5093,N_4440,N_4066);
xnor U5094 (N_5094,N_4514,N_4938);
or U5095 (N_5095,N_4681,N_4846);
xor U5096 (N_5096,N_4173,N_3873);
and U5097 (N_5097,N_3810,N_3833);
nand U5098 (N_5098,N_4285,N_4911);
nand U5099 (N_5099,N_3851,N_4329);
or U5100 (N_5100,N_3914,N_4551);
and U5101 (N_5101,N_3874,N_4207);
nand U5102 (N_5102,N_4665,N_4842);
xnor U5103 (N_5103,N_4134,N_4476);
or U5104 (N_5104,N_4856,N_4826);
nor U5105 (N_5105,N_4647,N_3879);
xor U5106 (N_5106,N_4092,N_4227);
nand U5107 (N_5107,N_4745,N_4389);
and U5108 (N_5108,N_4990,N_3906);
nor U5109 (N_5109,N_4008,N_4975);
nor U5110 (N_5110,N_4181,N_4239);
nor U5111 (N_5111,N_3784,N_4624);
xnor U5112 (N_5112,N_4286,N_4169);
and U5113 (N_5113,N_4853,N_3858);
and U5114 (N_5114,N_4506,N_3908);
nand U5115 (N_5115,N_4012,N_4774);
or U5116 (N_5116,N_4104,N_4191);
or U5117 (N_5117,N_4343,N_4333);
and U5118 (N_5118,N_4976,N_4816);
nand U5119 (N_5119,N_4155,N_3964);
xor U5120 (N_5120,N_4439,N_4464);
nor U5121 (N_5121,N_3806,N_4815);
nand U5122 (N_5122,N_4860,N_4018);
or U5123 (N_5123,N_4249,N_4386);
nor U5124 (N_5124,N_4209,N_4006);
or U5125 (N_5125,N_4787,N_4053);
and U5126 (N_5126,N_4964,N_4102);
nand U5127 (N_5127,N_4048,N_4490);
nor U5128 (N_5128,N_4031,N_4194);
and U5129 (N_5129,N_4472,N_4461);
or U5130 (N_5130,N_4766,N_4426);
or U5131 (N_5131,N_4118,N_4873);
xnor U5132 (N_5132,N_4327,N_4120);
and U5133 (N_5133,N_4325,N_4621);
or U5134 (N_5134,N_3924,N_4880);
xor U5135 (N_5135,N_4318,N_4547);
or U5136 (N_5136,N_4360,N_3753);
or U5137 (N_5137,N_4448,N_4541);
xnor U5138 (N_5138,N_4491,N_4383);
or U5139 (N_5139,N_3887,N_4280);
and U5140 (N_5140,N_4847,N_4302);
and U5141 (N_5141,N_3915,N_4743);
and U5142 (N_5142,N_3936,N_4044);
or U5143 (N_5143,N_4457,N_3997);
or U5144 (N_5144,N_3939,N_4148);
nor U5145 (N_5145,N_4437,N_4754);
or U5146 (N_5146,N_4002,N_4690);
or U5147 (N_5147,N_4339,N_4224);
and U5148 (N_5148,N_4277,N_4341);
nand U5149 (N_5149,N_4531,N_4546);
or U5150 (N_5150,N_3938,N_4763);
nand U5151 (N_5151,N_4131,N_4545);
nand U5152 (N_5152,N_4416,N_4347);
xnor U5153 (N_5153,N_4315,N_4459);
and U5154 (N_5154,N_4704,N_4984);
nor U5155 (N_5155,N_4297,N_4216);
nand U5156 (N_5156,N_4335,N_4289);
xor U5157 (N_5157,N_3891,N_4396);
nand U5158 (N_5158,N_4683,N_4074);
and U5159 (N_5159,N_4356,N_3781);
and U5160 (N_5160,N_4068,N_3957);
or U5161 (N_5161,N_4433,N_4390);
xnor U5162 (N_5162,N_4076,N_4370);
xor U5163 (N_5163,N_3978,N_4848);
nand U5164 (N_5164,N_3970,N_3959);
nand U5165 (N_5165,N_4179,N_4124);
nor U5166 (N_5166,N_4991,N_4451);
nand U5167 (N_5167,N_4299,N_4746);
nor U5168 (N_5168,N_4864,N_3948);
xnor U5169 (N_5169,N_4863,N_4675);
xnor U5170 (N_5170,N_3952,N_4662);
nand U5171 (N_5171,N_4178,N_4345);
or U5172 (N_5172,N_4144,N_4667);
or U5173 (N_5173,N_4791,N_4242);
or U5174 (N_5174,N_4247,N_4028);
or U5175 (N_5175,N_4740,N_3793);
nand U5176 (N_5176,N_4003,N_4139);
or U5177 (N_5177,N_4806,N_4693);
nand U5178 (N_5178,N_4572,N_4146);
nand U5179 (N_5179,N_4811,N_4837);
or U5180 (N_5180,N_4290,N_4999);
or U5181 (N_5181,N_4288,N_4604);
nand U5182 (N_5182,N_4544,N_4897);
nor U5183 (N_5183,N_4730,N_4449);
or U5184 (N_5184,N_4016,N_3982);
or U5185 (N_5185,N_4255,N_4180);
nor U5186 (N_5186,N_4537,N_4612);
nand U5187 (N_5187,N_3811,N_4308);
and U5188 (N_5188,N_4269,N_4010);
or U5189 (N_5189,N_4578,N_4885);
or U5190 (N_5190,N_4136,N_4468);
or U5191 (N_5191,N_4946,N_4477);
nand U5192 (N_5192,N_4907,N_4698);
and U5193 (N_5193,N_4737,N_4805);
nand U5194 (N_5194,N_4689,N_4958);
nand U5195 (N_5195,N_4858,N_4653);
nor U5196 (N_5196,N_4640,N_4757);
or U5197 (N_5197,N_4397,N_4919);
nand U5198 (N_5198,N_3943,N_4482);
or U5199 (N_5199,N_4521,N_4414);
nand U5200 (N_5200,N_4259,N_4529);
and U5201 (N_5201,N_4109,N_3889);
and U5202 (N_5202,N_3783,N_4123);
nand U5203 (N_5203,N_3911,N_4096);
nor U5204 (N_5204,N_4340,N_4713);
or U5205 (N_5205,N_3895,N_4953);
nor U5206 (N_5206,N_4300,N_4467);
and U5207 (N_5207,N_3866,N_4825);
xor U5208 (N_5208,N_4817,N_4781);
nor U5209 (N_5209,N_3849,N_4899);
or U5210 (N_5210,N_4429,N_4342);
nand U5211 (N_5211,N_4672,N_4354);
and U5212 (N_5212,N_4947,N_4363);
or U5213 (N_5213,N_4651,N_4232);
nand U5214 (N_5214,N_4152,N_4937);
and U5215 (N_5215,N_4955,N_4696);
nor U5216 (N_5216,N_4332,N_4184);
and U5217 (N_5217,N_3800,N_4425);
nor U5218 (N_5218,N_4534,N_4571);
and U5219 (N_5219,N_4660,N_3990);
or U5220 (N_5220,N_3893,N_4321);
or U5221 (N_5221,N_4934,N_4213);
xor U5222 (N_5222,N_4526,N_3750);
nand U5223 (N_5223,N_4887,N_3869);
or U5224 (N_5224,N_4619,N_4618);
nand U5225 (N_5225,N_4284,N_3995);
xnor U5226 (N_5226,N_4945,N_4485);
nor U5227 (N_5227,N_4789,N_4542);
xor U5228 (N_5228,N_4978,N_4081);
xor U5229 (N_5229,N_4409,N_4231);
nor U5230 (N_5230,N_3884,N_4500);
nand U5231 (N_5231,N_4196,N_4126);
xnor U5232 (N_5232,N_4441,N_4989);
nor U5233 (N_5233,N_4695,N_4268);
nand U5234 (N_5234,N_4981,N_4516);
nand U5235 (N_5235,N_4821,N_4128);
xor U5236 (N_5236,N_4957,N_4361);
nand U5237 (N_5237,N_4379,N_4328);
nand U5238 (N_5238,N_4687,N_4005);
nand U5239 (N_5239,N_4820,N_4963);
or U5240 (N_5240,N_4014,N_4434);
xor U5241 (N_5241,N_4750,N_4742);
nand U5242 (N_5242,N_3859,N_4865);
or U5243 (N_5243,N_4706,N_4548);
nor U5244 (N_5244,N_4786,N_3755);
or U5245 (N_5245,N_4636,N_4271);
nand U5246 (N_5246,N_3900,N_4273);
nand U5247 (N_5247,N_4839,N_4998);
nor U5248 (N_5248,N_4223,N_4428);
and U5249 (N_5249,N_4266,N_4725);
or U5250 (N_5250,N_4611,N_4644);
or U5251 (N_5251,N_4552,N_4495);
and U5252 (N_5252,N_4484,N_4956);
nand U5253 (N_5253,N_4163,N_4056);
and U5254 (N_5254,N_3923,N_4717);
and U5255 (N_5255,N_4854,N_4029);
or U5256 (N_5256,N_3760,N_4047);
or U5257 (N_5257,N_4966,N_4412);
and U5258 (N_5258,N_4079,N_4111);
nor U5259 (N_5259,N_3961,N_4025);
nand U5260 (N_5260,N_4993,N_4098);
or U5261 (N_5261,N_4089,N_3944);
or U5262 (N_5262,N_3871,N_4450);
and U5263 (N_5263,N_3969,N_4067);
or U5264 (N_5264,N_4900,N_4657);
nand U5265 (N_5265,N_4803,N_4380);
or U5266 (N_5266,N_4394,N_4844);
nand U5267 (N_5267,N_4862,N_3862);
nand U5268 (N_5268,N_3983,N_4894);
nor U5269 (N_5269,N_4494,N_4882);
or U5270 (N_5270,N_4275,N_4852);
xor U5271 (N_5271,N_4508,N_4685);
xor U5272 (N_5272,N_4313,N_4823);
and U5273 (N_5273,N_3826,N_4415);
and U5274 (N_5274,N_4217,N_4594);
nor U5275 (N_5275,N_4469,N_4645);
nor U5276 (N_5276,N_4940,N_3780);
nor U5277 (N_5277,N_4631,N_4941);
nand U5278 (N_5278,N_4809,N_3853);
nor U5279 (N_5279,N_3894,N_4013);
nor U5280 (N_5280,N_4793,N_4496);
and U5281 (N_5281,N_3976,N_4237);
nand U5282 (N_5282,N_4649,N_4822);
nand U5283 (N_5283,N_4115,N_4609);
xnor U5284 (N_5284,N_3965,N_3921);
nor U5285 (N_5285,N_3928,N_4749);
and U5286 (N_5286,N_4473,N_4466);
nor U5287 (N_5287,N_4444,N_4813);
or U5288 (N_5288,N_4855,N_3935);
nand U5289 (N_5289,N_4019,N_4637);
nor U5290 (N_5290,N_4423,N_4796);
or U5291 (N_5291,N_4920,N_4540);
or U5292 (N_5292,N_4027,N_4776);
nand U5293 (N_5293,N_4630,N_4753);
nand U5294 (N_5294,N_3788,N_4556);
xor U5295 (N_5295,N_4782,N_4658);
and U5296 (N_5296,N_3877,N_4186);
nor U5297 (N_5297,N_4119,N_3759);
nand U5298 (N_5298,N_4263,N_4460);
xor U5299 (N_5299,N_4203,N_3898);
or U5300 (N_5300,N_3803,N_4718);
nor U5301 (N_5301,N_4362,N_4393);
or U5302 (N_5302,N_4142,N_4723);
or U5303 (N_5303,N_4465,N_4075);
xnor U5304 (N_5304,N_4085,N_3918);
and U5305 (N_5305,N_4358,N_4033);
nor U5306 (N_5306,N_4678,N_3897);
nor U5307 (N_5307,N_4697,N_4036);
or U5308 (N_5308,N_4582,N_4158);
or U5309 (N_5309,N_4721,N_4929);
xor U5310 (N_5310,N_3808,N_4661);
nand U5311 (N_5311,N_4970,N_4599);
nor U5312 (N_5312,N_3912,N_3813);
nor U5313 (N_5313,N_4893,N_4087);
and U5314 (N_5314,N_4149,N_4543);
nand U5315 (N_5315,N_4932,N_4788);
nand U5316 (N_5316,N_4218,N_4488);
nand U5317 (N_5317,N_4810,N_4504);
nand U5318 (N_5318,N_4702,N_4387);
and U5319 (N_5319,N_4914,N_4590);
and U5320 (N_5320,N_3817,N_4095);
xnor U5321 (N_5321,N_3934,N_4629);
nand U5322 (N_5322,N_4261,N_4703);
or U5323 (N_5323,N_3776,N_4607);
and U5324 (N_5324,N_4442,N_4248);
xnor U5325 (N_5325,N_4253,N_4628);
or U5326 (N_5326,N_3967,N_4592);
and U5327 (N_5327,N_4034,N_4669);
nor U5328 (N_5328,N_4668,N_4765);
nand U5329 (N_5329,N_3821,N_3856);
nor U5330 (N_5330,N_4107,N_4600);
and U5331 (N_5331,N_4349,N_3863);
xor U5332 (N_5332,N_4807,N_4598);
and U5333 (N_5333,N_4405,N_4877);
nand U5334 (N_5334,N_4659,N_4587);
or U5335 (N_5335,N_3904,N_4670);
nand U5336 (N_5336,N_4694,N_4834);
or U5337 (N_5337,N_4747,N_3785);
xnor U5338 (N_5338,N_3868,N_4274);
nor U5339 (N_5339,N_4913,N_4518);
and U5340 (N_5340,N_4260,N_3789);
or U5341 (N_5341,N_4174,N_4479);
and U5342 (N_5342,N_4710,N_4072);
and U5343 (N_5343,N_4154,N_4641);
xnor U5344 (N_5344,N_4212,N_4064);
nor U5345 (N_5345,N_4655,N_4909);
and U5346 (N_5346,N_4617,N_3882);
or U5347 (N_5347,N_4264,N_3875);
xnor U5348 (N_5348,N_4368,N_4802);
xnor U5349 (N_5349,N_4244,N_4741);
nand U5350 (N_5350,N_3794,N_4601);
xnor U5351 (N_5351,N_4023,N_4711);
nor U5352 (N_5352,N_4375,N_4951);
xor U5353 (N_5353,N_4734,N_4391);
nand U5354 (N_5354,N_4395,N_4738);
nand U5355 (N_5355,N_4051,N_4241);
and U5356 (N_5356,N_4827,N_4801);
xor U5357 (N_5357,N_4654,N_3962);
nor U5358 (N_5358,N_3992,N_3852);
nand U5359 (N_5359,N_3963,N_4206);
or U5360 (N_5360,N_4593,N_4502);
nand U5361 (N_5361,N_4679,N_4575);
and U5362 (N_5362,N_3930,N_4171);
or U5363 (N_5363,N_4724,N_4832);
nor U5364 (N_5364,N_4764,N_4851);
or U5365 (N_5365,N_4293,N_4829);
and U5366 (N_5366,N_4314,N_4384);
nor U5367 (N_5367,N_4407,N_3955);
nor U5368 (N_5368,N_4366,N_4532);
or U5369 (N_5369,N_4530,N_4677);
or U5370 (N_5370,N_4200,N_4004);
or U5371 (N_5371,N_4836,N_3778);
and U5372 (N_5372,N_4652,N_4404);
nand U5373 (N_5373,N_4161,N_4985);
xnor U5374 (N_5374,N_4872,N_4091);
xor U5375 (N_5375,N_4254,N_4664);
nand U5376 (N_5376,N_4838,N_4962);
nand U5377 (N_5377,N_3807,N_3837);
nand U5378 (N_5378,N_4994,N_4114);
nor U5379 (N_5379,N_4728,N_4622);
nand U5380 (N_5380,N_4001,N_4559);
nor U5381 (N_5381,N_4850,N_3835);
nand U5382 (N_5382,N_3772,N_4870);
and U5383 (N_5383,N_4182,N_3903);
xor U5384 (N_5384,N_4135,N_3765);
nor U5385 (N_5385,N_4767,N_4973);
or U5386 (N_5386,N_4287,N_4463);
or U5387 (N_5387,N_3933,N_4310);
xnor U5388 (N_5388,N_4312,N_4967);
nand U5389 (N_5389,N_4157,N_3820);
xnor U5390 (N_5390,N_4480,N_3973);
xnor U5391 (N_5391,N_3966,N_4533);
xor U5392 (N_5392,N_4324,N_4319);
and U5393 (N_5393,N_4453,N_4814);
nor U5394 (N_5394,N_4235,N_4381);
nor U5395 (N_5395,N_4458,N_4486);
or U5396 (N_5396,N_4626,N_3854);
xnor U5397 (N_5397,N_4830,N_4777);
or U5398 (N_5398,N_4795,N_4077);
and U5399 (N_5399,N_4898,N_4122);
or U5400 (N_5400,N_4605,N_4202);
and U5401 (N_5401,N_4106,N_3981);
and U5402 (N_5402,N_3799,N_4137);
xor U5403 (N_5403,N_4961,N_4219);
nand U5404 (N_5404,N_4201,N_4510);
xnor U5405 (N_5405,N_4535,N_4770);
xor U5406 (N_5406,N_3842,N_4116);
or U5407 (N_5407,N_3857,N_4560);
xor U5408 (N_5408,N_3949,N_4565);
and U5409 (N_5409,N_4167,N_4859);
or U5410 (N_5410,N_4583,N_4987);
nand U5411 (N_5411,N_4265,N_4164);
nand U5412 (N_5412,N_4198,N_4052);
or U5413 (N_5413,N_4243,N_4041);
or U5414 (N_5414,N_4355,N_4121);
and U5415 (N_5415,N_4160,N_4819);
nand U5416 (N_5416,N_3945,N_4972);
xnor U5417 (N_5417,N_4861,N_3954);
or U5418 (N_5418,N_3860,N_4733);
or U5419 (N_5419,N_3757,N_4151);
or U5420 (N_5420,N_4262,N_3804);
and U5421 (N_5421,N_4402,N_3829);
xor U5422 (N_5422,N_4365,N_4931);
or U5423 (N_5423,N_3916,N_4113);
and U5424 (N_5424,N_4471,N_3864);
nor U5425 (N_5425,N_4969,N_4296);
and U5426 (N_5426,N_4835,N_4378);
xnor U5427 (N_5427,N_4739,N_4357);
nand U5428 (N_5428,N_4707,N_3896);
or U5429 (N_5429,N_4735,N_4939);
nor U5430 (N_5430,N_4915,N_4731);
nand U5431 (N_5431,N_4528,N_4258);
and U5432 (N_5432,N_3848,N_4876);
and U5433 (N_5433,N_4760,N_4603);
nand U5434 (N_5434,N_4177,N_4663);
nand U5435 (N_5435,N_3885,N_4099);
xor U5436 (N_5436,N_3913,N_4878);
xnor U5437 (N_5437,N_4623,N_4165);
xor U5438 (N_5438,N_3940,N_3892);
nor U5439 (N_5439,N_4306,N_4080);
or U5440 (N_5440,N_4926,N_4917);
and U5441 (N_5441,N_3796,N_4413);
nor U5442 (N_5442,N_3752,N_4236);
and U5443 (N_5443,N_3947,N_4895);
or U5444 (N_5444,N_4276,N_3922);
and U5445 (N_5445,N_4125,N_4138);
and U5446 (N_5446,N_4720,N_4891);
or U5447 (N_5447,N_4828,N_4779);
and U5448 (N_5448,N_4562,N_4352);
and U5449 (N_5449,N_4950,N_4638);
nand U5450 (N_5450,N_3956,N_3931);
nand U5451 (N_5451,N_4454,N_4032);
nor U5452 (N_5452,N_4840,N_4129);
or U5453 (N_5453,N_4211,N_4597);
and U5454 (N_5454,N_4039,N_4082);
nor U5455 (N_5455,N_3792,N_4561);
xnor U5456 (N_5456,N_4986,N_4060);
nor U5457 (N_5457,N_4676,N_4084);
or U5458 (N_5458,N_4769,N_3777);
nor U5459 (N_5459,N_3823,N_4869);
xor U5460 (N_5460,N_4517,N_3977);
xor U5461 (N_5461,N_4736,N_4557);
xnor U5462 (N_5462,N_4952,N_4055);
xnor U5463 (N_5463,N_4045,N_3917);
xor U5464 (N_5464,N_4699,N_4902);
nor U5465 (N_5465,N_4642,N_4643);
xnor U5466 (N_5466,N_4373,N_3960);
nor U5467 (N_5467,N_4147,N_4214);
nand U5468 (N_5468,N_4065,N_3839);
xor U5469 (N_5469,N_4057,N_4222);
xor U5470 (N_5470,N_4525,N_4511);
or U5471 (N_5471,N_4419,N_4112);
nor U5472 (N_5472,N_4455,N_3996);
and U5473 (N_5473,N_4935,N_4563);
xor U5474 (N_5474,N_4800,N_4944);
nand U5475 (N_5475,N_4187,N_4633);
nand U5476 (N_5476,N_3838,N_4481);
nand U5477 (N_5477,N_3855,N_4007);
and U5478 (N_5478,N_4026,N_4168);
nand U5479 (N_5479,N_3883,N_4520);
or U5480 (N_5480,N_3937,N_4427);
nor U5481 (N_5481,N_3825,N_4399);
or U5482 (N_5482,N_4596,N_4353);
or U5483 (N_5483,N_3998,N_4190);
xor U5484 (N_5484,N_4948,N_4549);
xnor U5485 (N_5485,N_3801,N_4634);
nand U5486 (N_5486,N_4371,N_4585);
and U5487 (N_5487,N_3979,N_3901);
nor U5488 (N_5488,N_3809,N_4432);
or U5489 (N_5489,N_3953,N_4326);
xnor U5490 (N_5490,N_3812,N_4613);
xor U5491 (N_5491,N_4505,N_4881);
nand U5492 (N_5492,N_4709,N_4376);
nor U5493 (N_5493,N_4691,N_4195);
nor U5494 (N_5494,N_4700,N_4705);
or U5495 (N_5495,N_4772,N_3767);
or U5496 (N_5496,N_4100,N_4550);
xor U5497 (N_5497,N_4751,N_4204);
nand U5498 (N_5498,N_4049,N_4996);
nor U5499 (N_5499,N_4348,N_4833);
xnor U5500 (N_5500,N_4988,N_4759);
nand U5501 (N_5501,N_4374,N_4192);
xor U5502 (N_5502,N_3974,N_3797);
and U5503 (N_5503,N_4197,N_3841);
and U5504 (N_5504,N_4576,N_4279);
or U5505 (N_5505,N_3786,N_3899);
nand U5506 (N_5506,N_4954,N_3929);
and U5507 (N_5507,N_4430,N_4780);
nand U5508 (N_5508,N_4616,N_4980);
xor U5509 (N_5509,N_4385,N_4977);
nor U5510 (N_5510,N_3795,N_4714);
nor U5511 (N_5511,N_4009,N_4523);
nor U5512 (N_5512,N_4435,N_4602);
nor U5513 (N_5513,N_3756,N_4928);
xnor U5514 (N_5514,N_4117,N_4043);
or U5515 (N_5515,N_4159,N_4338);
xnor U5516 (N_5516,N_4408,N_4684);
and U5517 (N_5517,N_3773,N_4410);
nor U5518 (N_5518,N_3909,N_4927);
or U5519 (N_5519,N_4431,N_4761);
xor U5520 (N_5520,N_4400,N_4558);
and U5521 (N_5521,N_4752,N_3822);
or U5522 (N_5522,N_4176,N_4968);
nand U5523 (N_5523,N_4493,N_3830);
and U5524 (N_5524,N_3840,N_4553);
xnor U5525 (N_5525,N_3986,N_4337);
or U5526 (N_5526,N_4101,N_4447);
xor U5527 (N_5527,N_3988,N_4475);
nand U5528 (N_5528,N_4997,N_4732);
nand U5529 (N_5529,N_4359,N_4252);
nand U5530 (N_5530,N_3751,N_3805);
nor U5531 (N_5531,N_4798,N_4487);
nand U5532 (N_5532,N_4824,N_3766);
or U5533 (N_5533,N_4871,N_4141);
xor U5534 (N_5534,N_4130,N_4648);
nor U5535 (N_5535,N_4411,N_4323);
or U5536 (N_5536,N_4350,N_4843);
nor U5537 (N_5537,N_4903,N_3987);
xnor U5538 (N_5538,N_3834,N_4078);
nor U5539 (N_5539,N_3763,N_4785);
nand U5540 (N_5540,N_4311,N_4890);
or U5541 (N_5541,N_3782,N_4892);
nor U5542 (N_5542,N_4035,N_4108);
or U5543 (N_5543,N_4783,N_4744);
nand U5544 (N_5544,N_4868,N_4588);
nor U5545 (N_5545,N_3861,N_4942);
and U5546 (N_5546,N_4921,N_4775);
and U5547 (N_5547,N_4509,N_4886);
or U5548 (N_5548,N_4017,N_4040);
and U5549 (N_5549,N_4346,N_4586);
nor U5550 (N_5550,N_4673,N_3761);
nor U5551 (N_5551,N_4686,N_3968);
xor U5552 (N_5552,N_3925,N_3816);
nand U5553 (N_5553,N_4555,N_3775);
and U5554 (N_5554,N_4650,N_4627);
nand U5555 (N_5555,N_3991,N_3779);
nor U5556 (N_5556,N_3836,N_3876);
nand U5557 (N_5557,N_3972,N_4646);
nand U5558 (N_5558,N_4688,N_4756);
and U5559 (N_5559,N_3878,N_4071);
nor U5560 (N_5560,N_4298,N_4610);
or U5561 (N_5561,N_4474,N_4875);
nand U5562 (N_5562,N_4251,N_3850);
or U5563 (N_5563,N_4294,N_4498);
or U5564 (N_5564,N_4818,N_4093);
nor U5565 (N_5565,N_4515,N_4021);
xnor U5566 (N_5566,N_4156,N_4406);
or U5567 (N_5567,N_4905,N_3844);
xor U5568 (N_5568,N_4933,N_4845);
nand U5569 (N_5569,N_3984,N_4632);
nor U5570 (N_5570,N_4372,N_3870);
xor U5571 (N_5571,N_4729,N_4922);
nand U5572 (N_5572,N_3946,N_4443);
nand U5573 (N_5573,N_4170,N_4584);
nor U5574 (N_5574,N_3824,N_4246);
or U5575 (N_5575,N_4304,N_4418);
xnor U5576 (N_5576,N_4445,N_4712);
xor U5577 (N_5577,N_4220,N_4185);
nand U5578 (N_5578,N_4038,N_4042);
or U5579 (N_5579,N_3845,N_4790);
nor U5580 (N_5580,N_4538,N_4536);
or U5581 (N_5581,N_4570,N_4758);
nor U5582 (N_5582,N_3768,N_4388);
nor U5583 (N_5583,N_3802,N_4291);
xnor U5584 (N_5584,N_4680,N_3846);
xor U5585 (N_5585,N_4768,N_4305);
xor U5586 (N_5586,N_4925,N_3999);
xor U5587 (N_5587,N_4011,N_4566);
and U5588 (N_5588,N_4367,N_4417);
nand U5589 (N_5589,N_4070,N_4527);
xor U5590 (N_5590,N_4238,N_4320);
and U5591 (N_5591,N_3771,N_3888);
nor U5592 (N_5592,N_3832,N_4210);
or U5593 (N_5593,N_4497,N_4595);
nand U5594 (N_5594,N_4334,N_4403);
nand U5595 (N_5595,N_4519,N_4522);
nor U5596 (N_5596,N_3764,N_4150);
or U5597 (N_5597,N_4162,N_4309);
nand U5598 (N_5598,N_3951,N_4478);
xnor U5599 (N_5599,N_4857,N_4424);
xnor U5600 (N_5600,N_3926,N_4923);
xnor U5601 (N_5601,N_4577,N_3818);
nand U5602 (N_5602,N_4507,N_4489);
nor U5603 (N_5603,N_4090,N_3815);
nor U5604 (N_5604,N_4799,N_4918);
and U5605 (N_5605,N_3890,N_4037);
xor U5606 (N_5606,N_4671,N_4874);
and U5607 (N_5607,N_4283,N_4524);
nand U5608 (N_5608,N_4971,N_4608);
nand U5609 (N_5609,N_4960,N_4257);
nand U5610 (N_5610,N_4398,N_3867);
or U5611 (N_5611,N_4904,N_4784);
xnor U5612 (N_5612,N_4281,N_4054);
nand U5613 (N_5613,N_4656,N_4974);
nand U5614 (N_5614,N_4849,N_4208);
or U5615 (N_5615,N_4910,N_4015);
nand U5616 (N_5616,N_4715,N_4421);
and U5617 (N_5617,N_3769,N_4295);
or U5618 (N_5618,N_4240,N_4050);
or U5619 (N_5619,N_4127,N_4512);
and U5620 (N_5620,N_4143,N_4771);
nor U5621 (N_5621,N_4615,N_4250);
or U5622 (N_5622,N_4716,N_4094);
nand U5623 (N_5623,N_3980,N_3902);
xnor U5624 (N_5624,N_4983,N_4906);
and U5625 (N_5625,N_3753,N_4276);
xnor U5626 (N_5626,N_3960,N_3875);
nor U5627 (N_5627,N_3760,N_4324);
nor U5628 (N_5628,N_3822,N_4535);
xor U5629 (N_5629,N_4671,N_4948);
nor U5630 (N_5630,N_3863,N_4300);
nand U5631 (N_5631,N_4753,N_4590);
nand U5632 (N_5632,N_4105,N_4364);
nand U5633 (N_5633,N_4640,N_4945);
or U5634 (N_5634,N_4401,N_3922);
or U5635 (N_5635,N_4899,N_4944);
xor U5636 (N_5636,N_4312,N_4303);
nor U5637 (N_5637,N_3966,N_4292);
nor U5638 (N_5638,N_4925,N_3794);
nand U5639 (N_5639,N_4762,N_3861);
or U5640 (N_5640,N_4108,N_4151);
and U5641 (N_5641,N_4824,N_4048);
or U5642 (N_5642,N_4050,N_4423);
nand U5643 (N_5643,N_4932,N_4460);
and U5644 (N_5644,N_4921,N_4154);
and U5645 (N_5645,N_4847,N_4823);
and U5646 (N_5646,N_4729,N_4816);
nand U5647 (N_5647,N_4872,N_4171);
nor U5648 (N_5648,N_4807,N_3875);
and U5649 (N_5649,N_4800,N_4471);
nor U5650 (N_5650,N_4133,N_4404);
nor U5651 (N_5651,N_3982,N_4556);
xor U5652 (N_5652,N_4293,N_4813);
and U5653 (N_5653,N_4405,N_4139);
and U5654 (N_5654,N_4267,N_4430);
and U5655 (N_5655,N_4679,N_3857);
or U5656 (N_5656,N_3762,N_4614);
nor U5657 (N_5657,N_4728,N_4120);
nand U5658 (N_5658,N_4481,N_3890);
nor U5659 (N_5659,N_4282,N_4539);
nand U5660 (N_5660,N_4762,N_3875);
and U5661 (N_5661,N_4366,N_4910);
nand U5662 (N_5662,N_4996,N_4346);
and U5663 (N_5663,N_4451,N_4239);
nand U5664 (N_5664,N_4404,N_4054);
xnor U5665 (N_5665,N_4372,N_4321);
nor U5666 (N_5666,N_4624,N_4695);
nand U5667 (N_5667,N_4607,N_3902);
xnor U5668 (N_5668,N_4959,N_3828);
xnor U5669 (N_5669,N_4348,N_4846);
and U5670 (N_5670,N_4370,N_3953);
and U5671 (N_5671,N_4462,N_4291);
nor U5672 (N_5672,N_4636,N_4982);
xnor U5673 (N_5673,N_4394,N_4929);
nand U5674 (N_5674,N_4209,N_3951);
nand U5675 (N_5675,N_4371,N_4572);
nand U5676 (N_5676,N_4663,N_4743);
nand U5677 (N_5677,N_4765,N_3931);
or U5678 (N_5678,N_4235,N_4999);
and U5679 (N_5679,N_4187,N_4568);
nand U5680 (N_5680,N_3987,N_3785);
nand U5681 (N_5681,N_4633,N_4161);
nand U5682 (N_5682,N_4874,N_4377);
and U5683 (N_5683,N_3822,N_4165);
or U5684 (N_5684,N_4003,N_4615);
nand U5685 (N_5685,N_4085,N_4515);
xor U5686 (N_5686,N_4981,N_3892);
nor U5687 (N_5687,N_3804,N_4323);
nor U5688 (N_5688,N_4681,N_4294);
and U5689 (N_5689,N_4845,N_4311);
nor U5690 (N_5690,N_3907,N_3995);
xor U5691 (N_5691,N_4588,N_4038);
and U5692 (N_5692,N_4293,N_4313);
and U5693 (N_5693,N_4614,N_4856);
and U5694 (N_5694,N_4795,N_4322);
or U5695 (N_5695,N_4445,N_4865);
nand U5696 (N_5696,N_4251,N_4499);
nor U5697 (N_5697,N_4974,N_4866);
nand U5698 (N_5698,N_4944,N_4239);
nand U5699 (N_5699,N_4724,N_4815);
or U5700 (N_5700,N_4203,N_4457);
or U5701 (N_5701,N_3863,N_4255);
nand U5702 (N_5702,N_3901,N_4165);
xnor U5703 (N_5703,N_4596,N_3785);
nand U5704 (N_5704,N_4007,N_3843);
and U5705 (N_5705,N_4148,N_4364);
nor U5706 (N_5706,N_4875,N_4342);
nand U5707 (N_5707,N_3989,N_4693);
or U5708 (N_5708,N_4707,N_4100);
nand U5709 (N_5709,N_4879,N_4804);
and U5710 (N_5710,N_4080,N_4139);
nand U5711 (N_5711,N_4074,N_3772);
nor U5712 (N_5712,N_4408,N_4945);
nand U5713 (N_5713,N_4352,N_4079);
and U5714 (N_5714,N_4072,N_4903);
nand U5715 (N_5715,N_4449,N_4275);
nor U5716 (N_5716,N_3841,N_3929);
xor U5717 (N_5717,N_4074,N_4274);
and U5718 (N_5718,N_3915,N_4051);
or U5719 (N_5719,N_4383,N_4975);
or U5720 (N_5720,N_3940,N_4231);
and U5721 (N_5721,N_4682,N_4077);
nand U5722 (N_5722,N_3788,N_4779);
xor U5723 (N_5723,N_4353,N_4100);
or U5724 (N_5724,N_4246,N_4421);
and U5725 (N_5725,N_4774,N_4177);
or U5726 (N_5726,N_4304,N_4943);
nor U5727 (N_5727,N_4500,N_3794);
xor U5728 (N_5728,N_4699,N_4426);
xor U5729 (N_5729,N_4272,N_4764);
nand U5730 (N_5730,N_4551,N_4891);
or U5731 (N_5731,N_4605,N_4459);
nand U5732 (N_5732,N_4917,N_4008);
nand U5733 (N_5733,N_4411,N_3916);
nor U5734 (N_5734,N_4825,N_3790);
nand U5735 (N_5735,N_4077,N_4459);
xor U5736 (N_5736,N_4659,N_4145);
and U5737 (N_5737,N_4556,N_4620);
nor U5738 (N_5738,N_3825,N_4577);
xor U5739 (N_5739,N_3783,N_4312);
nand U5740 (N_5740,N_3851,N_4567);
or U5741 (N_5741,N_3804,N_4991);
nand U5742 (N_5742,N_4315,N_4530);
nor U5743 (N_5743,N_3938,N_4130);
or U5744 (N_5744,N_4605,N_4194);
xnor U5745 (N_5745,N_4245,N_4088);
nor U5746 (N_5746,N_4717,N_4563);
xnor U5747 (N_5747,N_3933,N_3987);
or U5748 (N_5748,N_4730,N_4416);
xor U5749 (N_5749,N_4980,N_4609);
xor U5750 (N_5750,N_3768,N_4523);
nand U5751 (N_5751,N_4758,N_4347);
nor U5752 (N_5752,N_4186,N_4826);
or U5753 (N_5753,N_4975,N_3850);
or U5754 (N_5754,N_4586,N_3961);
nand U5755 (N_5755,N_3814,N_4309);
or U5756 (N_5756,N_3896,N_4332);
or U5757 (N_5757,N_4033,N_4079);
or U5758 (N_5758,N_4539,N_4897);
nor U5759 (N_5759,N_4227,N_4052);
xnor U5760 (N_5760,N_4536,N_4059);
nand U5761 (N_5761,N_3775,N_3859);
xnor U5762 (N_5762,N_3801,N_4591);
nand U5763 (N_5763,N_4631,N_3881);
nor U5764 (N_5764,N_4338,N_4925);
and U5765 (N_5765,N_4487,N_4314);
nor U5766 (N_5766,N_3911,N_4272);
or U5767 (N_5767,N_4377,N_4036);
and U5768 (N_5768,N_4888,N_4843);
and U5769 (N_5769,N_4169,N_4613);
or U5770 (N_5770,N_4615,N_3778);
xor U5771 (N_5771,N_4225,N_4914);
xor U5772 (N_5772,N_4827,N_4997);
xor U5773 (N_5773,N_4126,N_4545);
or U5774 (N_5774,N_4127,N_3983);
and U5775 (N_5775,N_4387,N_4000);
nor U5776 (N_5776,N_4705,N_4557);
nand U5777 (N_5777,N_4427,N_4842);
and U5778 (N_5778,N_4470,N_4998);
nor U5779 (N_5779,N_3980,N_4674);
nor U5780 (N_5780,N_4569,N_4596);
nand U5781 (N_5781,N_4564,N_4343);
and U5782 (N_5782,N_3879,N_3790);
or U5783 (N_5783,N_3877,N_4026);
and U5784 (N_5784,N_4664,N_4895);
nand U5785 (N_5785,N_4247,N_3964);
xnor U5786 (N_5786,N_4049,N_4225);
nor U5787 (N_5787,N_4267,N_4126);
nand U5788 (N_5788,N_4210,N_3921);
nor U5789 (N_5789,N_4854,N_4896);
nand U5790 (N_5790,N_4605,N_4825);
nor U5791 (N_5791,N_4826,N_3952);
nand U5792 (N_5792,N_4373,N_4236);
nor U5793 (N_5793,N_3793,N_4699);
and U5794 (N_5794,N_4889,N_4230);
nor U5795 (N_5795,N_4356,N_4224);
or U5796 (N_5796,N_4633,N_4103);
and U5797 (N_5797,N_3781,N_4139);
and U5798 (N_5798,N_4727,N_4733);
xnor U5799 (N_5799,N_4487,N_3920);
and U5800 (N_5800,N_4660,N_4153);
nor U5801 (N_5801,N_4477,N_4744);
nor U5802 (N_5802,N_4255,N_4931);
and U5803 (N_5803,N_4802,N_4976);
nor U5804 (N_5804,N_4205,N_4289);
and U5805 (N_5805,N_4053,N_4540);
xor U5806 (N_5806,N_3975,N_3967);
nand U5807 (N_5807,N_4352,N_4654);
nand U5808 (N_5808,N_4924,N_4692);
and U5809 (N_5809,N_4985,N_4481);
xor U5810 (N_5810,N_4099,N_4948);
or U5811 (N_5811,N_4961,N_4093);
nor U5812 (N_5812,N_4282,N_4910);
xor U5813 (N_5813,N_4771,N_3826);
nand U5814 (N_5814,N_4476,N_4198);
or U5815 (N_5815,N_4564,N_3864);
and U5816 (N_5816,N_4285,N_4150);
and U5817 (N_5817,N_4995,N_3866);
and U5818 (N_5818,N_4881,N_4095);
nor U5819 (N_5819,N_4777,N_4438);
or U5820 (N_5820,N_4769,N_3967);
nand U5821 (N_5821,N_3779,N_3876);
or U5822 (N_5822,N_3921,N_3813);
nand U5823 (N_5823,N_4554,N_3982);
and U5824 (N_5824,N_4561,N_4205);
xor U5825 (N_5825,N_4886,N_4284);
or U5826 (N_5826,N_4632,N_4046);
xor U5827 (N_5827,N_4234,N_4546);
nand U5828 (N_5828,N_3781,N_4326);
nor U5829 (N_5829,N_3763,N_4777);
and U5830 (N_5830,N_4605,N_4637);
or U5831 (N_5831,N_3945,N_3757);
xnor U5832 (N_5832,N_4125,N_3775);
nand U5833 (N_5833,N_4600,N_4704);
nor U5834 (N_5834,N_4507,N_4430);
or U5835 (N_5835,N_4236,N_4899);
or U5836 (N_5836,N_4588,N_4385);
and U5837 (N_5837,N_4047,N_4221);
or U5838 (N_5838,N_3858,N_3829);
and U5839 (N_5839,N_3817,N_4701);
or U5840 (N_5840,N_4717,N_4015);
xnor U5841 (N_5841,N_3867,N_4397);
and U5842 (N_5842,N_4750,N_3949);
or U5843 (N_5843,N_3946,N_4158);
nor U5844 (N_5844,N_3947,N_4853);
nor U5845 (N_5845,N_4675,N_4381);
nor U5846 (N_5846,N_4885,N_4689);
nand U5847 (N_5847,N_3902,N_4621);
nand U5848 (N_5848,N_4782,N_3837);
or U5849 (N_5849,N_4888,N_3895);
and U5850 (N_5850,N_4879,N_4341);
nor U5851 (N_5851,N_4761,N_4916);
and U5852 (N_5852,N_4575,N_3884);
and U5853 (N_5853,N_4400,N_3947);
and U5854 (N_5854,N_4705,N_4136);
nand U5855 (N_5855,N_4137,N_4643);
or U5856 (N_5856,N_4019,N_3836);
nor U5857 (N_5857,N_4139,N_4097);
and U5858 (N_5858,N_4180,N_4402);
or U5859 (N_5859,N_4711,N_3794);
or U5860 (N_5860,N_4339,N_4487);
nand U5861 (N_5861,N_3900,N_4840);
nand U5862 (N_5862,N_4456,N_4287);
and U5863 (N_5863,N_3995,N_4861);
xnor U5864 (N_5864,N_4245,N_4221);
nand U5865 (N_5865,N_3803,N_3837);
and U5866 (N_5866,N_3964,N_4878);
nor U5867 (N_5867,N_4332,N_4763);
xnor U5868 (N_5868,N_4549,N_4375);
nor U5869 (N_5869,N_4055,N_4274);
or U5870 (N_5870,N_4983,N_3848);
nor U5871 (N_5871,N_4266,N_3816);
or U5872 (N_5872,N_4753,N_4042);
xnor U5873 (N_5873,N_3810,N_4138);
nand U5874 (N_5874,N_4612,N_3767);
and U5875 (N_5875,N_4414,N_4506);
nand U5876 (N_5876,N_4905,N_3833);
nor U5877 (N_5877,N_4696,N_4872);
nand U5878 (N_5878,N_4103,N_3844);
and U5879 (N_5879,N_3969,N_4138);
and U5880 (N_5880,N_4905,N_4152);
nor U5881 (N_5881,N_4758,N_4447);
nand U5882 (N_5882,N_4486,N_3752);
nor U5883 (N_5883,N_4529,N_3825);
nand U5884 (N_5884,N_4694,N_4017);
and U5885 (N_5885,N_4597,N_4406);
nand U5886 (N_5886,N_4657,N_4434);
xor U5887 (N_5887,N_4441,N_4913);
and U5888 (N_5888,N_3780,N_3940);
nand U5889 (N_5889,N_4003,N_4961);
or U5890 (N_5890,N_4660,N_4502);
nand U5891 (N_5891,N_4245,N_4824);
and U5892 (N_5892,N_4464,N_4293);
or U5893 (N_5893,N_4124,N_4435);
and U5894 (N_5894,N_4357,N_4923);
or U5895 (N_5895,N_4859,N_4181);
nor U5896 (N_5896,N_3957,N_4758);
and U5897 (N_5897,N_4524,N_3794);
or U5898 (N_5898,N_4135,N_3992);
and U5899 (N_5899,N_4973,N_4134);
nor U5900 (N_5900,N_4858,N_4898);
nor U5901 (N_5901,N_4547,N_4163);
or U5902 (N_5902,N_4218,N_3866);
xor U5903 (N_5903,N_4647,N_4021);
xor U5904 (N_5904,N_4107,N_4208);
and U5905 (N_5905,N_3997,N_4433);
nor U5906 (N_5906,N_4414,N_4312);
nand U5907 (N_5907,N_4490,N_4343);
xnor U5908 (N_5908,N_4564,N_3845);
or U5909 (N_5909,N_4476,N_4307);
nand U5910 (N_5910,N_4092,N_4124);
nor U5911 (N_5911,N_4274,N_3871);
nor U5912 (N_5912,N_3974,N_4074);
nand U5913 (N_5913,N_4805,N_4040);
and U5914 (N_5914,N_4292,N_4388);
xnor U5915 (N_5915,N_4623,N_4944);
and U5916 (N_5916,N_4038,N_4856);
or U5917 (N_5917,N_4332,N_4645);
nand U5918 (N_5918,N_4309,N_3925);
nand U5919 (N_5919,N_3884,N_3902);
nand U5920 (N_5920,N_3754,N_4185);
and U5921 (N_5921,N_4774,N_4408);
or U5922 (N_5922,N_4996,N_4488);
and U5923 (N_5923,N_4082,N_4816);
nor U5924 (N_5924,N_3875,N_4147);
nand U5925 (N_5925,N_4601,N_4528);
and U5926 (N_5926,N_3798,N_3950);
nand U5927 (N_5927,N_4057,N_4132);
nand U5928 (N_5928,N_4701,N_4386);
and U5929 (N_5929,N_4610,N_4814);
nand U5930 (N_5930,N_4373,N_4163);
nand U5931 (N_5931,N_4867,N_4381);
nand U5932 (N_5932,N_4607,N_4139);
or U5933 (N_5933,N_3800,N_4288);
and U5934 (N_5934,N_4697,N_4825);
nand U5935 (N_5935,N_4210,N_4639);
nand U5936 (N_5936,N_4242,N_4124);
xor U5937 (N_5937,N_4319,N_3850);
or U5938 (N_5938,N_4026,N_4707);
xnor U5939 (N_5939,N_3902,N_4623);
xor U5940 (N_5940,N_3930,N_4322);
and U5941 (N_5941,N_4133,N_4039);
xor U5942 (N_5942,N_4642,N_4037);
xor U5943 (N_5943,N_4657,N_4841);
or U5944 (N_5944,N_4631,N_4553);
nand U5945 (N_5945,N_4983,N_4284);
xnor U5946 (N_5946,N_4513,N_4069);
and U5947 (N_5947,N_4914,N_4108);
xnor U5948 (N_5948,N_4422,N_4274);
nor U5949 (N_5949,N_4607,N_4432);
nand U5950 (N_5950,N_4503,N_4408);
and U5951 (N_5951,N_4762,N_4241);
or U5952 (N_5952,N_4338,N_4576);
nand U5953 (N_5953,N_4246,N_3759);
nand U5954 (N_5954,N_4721,N_4675);
and U5955 (N_5955,N_3806,N_4665);
nand U5956 (N_5956,N_4282,N_4635);
or U5957 (N_5957,N_4441,N_4607);
or U5958 (N_5958,N_4472,N_4085);
and U5959 (N_5959,N_4069,N_3767);
or U5960 (N_5960,N_3945,N_4935);
nor U5961 (N_5961,N_4894,N_3807);
and U5962 (N_5962,N_4714,N_4311);
nor U5963 (N_5963,N_4229,N_3887);
or U5964 (N_5964,N_4482,N_4191);
or U5965 (N_5965,N_4020,N_4114);
or U5966 (N_5966,N_4052,N_4830);
xor U5967 (N_5967,N_4225,N_4963);
or U5968 (N_5968,N_4158,N_4238);
or U5969 (N_5969,N_4328,N_4531);
nor U5970 (N_5970,N_4708,N_4817);
or U5971 (N_5971,N_4020,N_4359);
xnor U5972 (N_5972,N_3791,N_4740);
nand U5973 (N_5973,N_4034,N_4334);
or U5974 (N_5974,N_3897,N_3851);
nor U5975 (N_5975,N_4755,N_4641);
or U5976 (N_5976,N_4844,N_4843);
or U5977 (N_5977,N_3886,N_4342);
or U5978 (N_5978,N_4411,N_4554);
xor U5979 (N_5979,N_4882,N_4011);
or U5980 (N_5980,N_3988,N_4680);
nor U5981 (N_5981,N_4423,N_4073);
xor U5982 (N_5982,N_4814,N_4073);
and U5983 (N_5983,N_4557,N_4778);
nor U5984 (N_5984,N_3921,N_3989);
nor U5985 (N_5985,N_4612,N_4319);
or U5986 (N_5986,N_4164,N_3891);
nor U5987 (N_5987,N_4909,N_4085);
xnor U5988 (N_5988,N_3925,N_3986);
xnor U5989 (N_5989,N_4284,N_3795);
and U5990 (N_5990,N_4915,N_4391);
xnor U5991 (N_5991,N_4189,N_4542);
or U5992 (N_5992,N_4921,N_4423);
or U5993 (N_5993,N_4546,N_4385);
nor U5994 (N_5994,N_4100,N_4511);
nor U5995 (N_5995,N_4847,N_4764);
and U5996 (N_5996,N_3820,N_4267);
nor U5997 (N_5997,N_4513,N_4701);
or U5998 (N_5998,N_3972,N_4068);
or U5999 (N_5999,N_4706,N_4775);
nand U6000 (N_6000,N_4270,N_3779);
and U6001 (N_6001,N_4705,N_4454);
nor U6002 (N_6002,N_4140,N_4767);
or U6003 (N_6003,N_3888,N_4357);
and U6004 (N_6004,N_4174,N_4929);
nor U6005 (N_6005,N_3991,N_4674);
nand U6006 (N_6006,N_4072,N_4917);
and U6007 (N_6007,N_4674,N_3808);
and U6008 (N_6008,N_4404,N_4309);
xor U6009 (N_6009,N_4390,N_3760);
and U6010 (N_6010,N_4678,N_4563);
nand U6011 (N_6011,N_4690,N_4674);
nand U6012 (N_6012,N_4946,N_4274);
nand U6013 (N_6013,N_4576,N_4309);
nand U6014 (N_6014,N_4223,N_4646);
or U6015 (N_6015,N_4611,N_4027);
nand U6016 (N_6016,N_3851,N_4437);
or U6017 (N_6017,N_3929,N_4999);
and U6018 (N_6018,N_3921,N_4671);
or U6019 (N_6019,N_3966,N_4843);
or U6020 (N_6020,N_4007,N_4346);
nand U6021 (N_6021,N_4371,N_4332);
xnor U6022 (N_6022,N_4160,N_4861);
nand U6023 (N_6023,N_3945,N_4343);
xor U6024 (N_6024,N_4595,N_3826);
and U6025 (N_6025,N_4817,N_4551);
and U6026 (N_6026,N_4214,N_4473);
nand U6027 (N_6027,N_4987,N_4652);
xor U6028 (N_6028,N_4644,N_4414);
and U6029 (N_6029,N_4082,N_4298);
or U6030 (N_6030,N_4197,N_4585);
and U6031 (N_6031,N_4812,N_3913);
nand U6032 (N_6032,N_4709,N_4904);
xor U6033 (N_6033,N_4754,N_4902);
nand U6034 (N_6034,N_4406,N_4177);
or U6035 (N_6035,N_4115,N_3812);
and U6036 (N_6036,N_4617,N_3822);
nor U6037 (N_6037,N_4713,N_4202);
xnor U6038 (N_6038,N_4973,N_4459);
and U6039 (N_6039,N_4722,N_4927);
and U6040 (N_6040,N_4515,N_4637);
nand U6041 (N_6041,N_4850,N_4293);
and U6042 (N_6042,N_4710,N_4544);
nor U6043 (N_6043,N_4938,N_4846);
xnor U6044 (N_6044,N_4177,N_4271);
or U6045 (N_6045,N_4079,N_4861);
or U6046 (N_6046,N_4309,N_4231);
and U6047 (N_6047,N_4805,N_3830);
or U6048 (N_6048,N_4294,N_4295);
and U6049 (N_6049,N_4411,N_3895);
xnor U6050 (N_6050,N_4419,N_4357);
xnor U6051 (N_6051,N_3887,N_3858);
xnor U6052 (N_6052,N_3819,N_4066);
or U6053 (N_6053,N_4228,N_4466);
nand U6054 (N_6054,N_4582,N_3816);
xor U6055 (N_6055,N_4078,N_4181);
or U6056 (N_6056,N_4676,N_4079);
and U6057 (N_6057,N_4158,N_3991);
and U6058 (N_6058,N_3760,N_3781);
or U6059 (N_6059,N_4561,N_4926);
or U6060 (N_6060,N_4318,N_4099);
and U6061 (N_6061,N_4883,N_4412);
and U6062 (N_6062,N_4845,N_3785);
and U6063 (N_6063,N_4968,N_4239);
nor U6064 (N_6064,N_4207,N_4532);
nor U6065 (N_6065,N_3817,N_4223);
nand U6066 (N_6066,N_4650,N_3792);
and U6067 (N_6067,N_4819,N_4455);
xnor U6068 (N_6068,N_4981,N_3750);
nand U6069 (N_6069,N_4646,N_4265);
and U6070 (N_6070,N_4839,N_4900);
nor U6071 (N_6071,N_4712,N_4867);
or U6072 (N_6072,N_4095,N_4346);
xnor U6073 (N_6073,N_4321,N_4732);
and U6074 (N_6074,N_4756,N_4457);
nor U6075 (N_6075,N_4445,N_4340);
nand U6076 (N_6076,N_4278,N_4010);
xnor U6077 (N_6077,N_4476,N_4700);
nor U6078 (N_6078,N_4860,N_3786);
nand U6079 (N_6079,N_4459,N_4731);
nor U6080 (N_6080,N_4400,N_4902);
and U6081 (N_6081,N_4821,N_4084);
or U6082 (N_6082,N_4257,N_4619);
xnor U6083 (N_6083,N_3778,N_4067);
or U6084 (N_6084,N_4141,N_4936);
xnor U6085 (N_6085,N_4608,N_4874);
xor U6086 (N_6086,N_3822,N_4353);
nand U6087 (N_6087,N_4196,N_3801);
nor U6088 (N_6088,N_4238,N_4964);
and U6089 (N_6089,N_4213,N_4015);
nand U6090 (N_6090,N_4051,N_3796);
xnor U6091 (N_6091,N_4020,N_4757);
nand U6092 (N_6092,N_3840,N_4919);
or U6093 (N_6093,N_3791,N_4145);
xor U6094 (N_6094,N_4004,N_4334);
and U6095 (N_6095,N_4461,N_3955);
nand U6096 (N_6096,N_4431,N_3990);
xor U6097 (N_6097,N_4666,N_3959);
or U6098 (N_6098,N_3985,N_3853);
nor U6099 (N_6099,N_3805,N_4851);
xor U6100 (N_6100,N_4429,N_3858);
and U6101 (N_6101,N_3890,N_4605);
and U6102 (N_6102,N_4838,N_4041);
xnor U6103 (N_6103,N_4371,N_3871);
xor U6104 (N_6104,N_3907,N_4937);
nor U6105 (N_6105,N_3874,N_4153);
and U6106 (N_6106,N_4991,N_4877);
nor U6107 (N_6107,N_4893,N_3837);
xor U6108 (N_6108,N_4862,N_4778);
or U6109 (N_6109,N_4263,N_3984);
nand U6110 (N_6110,N_3888,N_4542);
xor U6111 (N_6111,N_3862,N_4333);
nand U6112 (N_6112,N_4531,N_4547);
nor U6113 (N_6113,N_4858,N_4797);
nand U6114 (N_6114,N_3815,N_4303);
or U6115 (N_6115,N_3925,N_4511);
nor U6116 (N_6116,N_4880,N_4373);
nand U6117 (N_6117,N_4060,N_4090);
nand U6118 (N_6118,N_4891,N_4920);
and U6119 (N_6119,N_3771,N_4349);
or U6120 (N_6120,N_4351,N_4732);
or U6121 (N_6121,N_4396,N_4729);
nor U6122 (N_6122,N_4611,N_4747);
xor U6123 (N_6123,N_4956,N_4980);
nor U6124 (N_6124,N_4715,N_4279);
nor U6125 (N_6125,N_4814,N_4304);
and U6126 (N_6126,N_3942,N_4406);
or U6127 (N_6127,N_3945,N_4697);
or U6128 (N_6128,N_4013,N_4416);
nor U6129 (N_6129,N_3987,N_4252);
nor U6130 (N_6130,N_4884,N_3889);
nor U6131 (N_6131,N_4954,N_4751);
and U6132 (N_6132,N_3778,N_3761);
nand U6133 (N_6133,N_4421,N_4090);
or U6134 (N_6134,N_3891,N_3764);
nand U6135 (N_6135,N_4999,N_4669);
or U6136 (N_6136,N_4808,N_4430);
nand U6137 (N_6137,N_4123,N_3751);
nand U6138 (N_6138,N_4913,N_3951);
nor U6139 (N_6139,N_3994,N_4762);
nor U6140 (N_6140,N_4717,N_3930);
or U6141 (N_6141,N_3955,N_4982);
nor U6142 (N_6142,N_3860,N_4323);
nor U6143 (N_6143,N_3996,N_4711);
xnor U6144 (N_6144,N_4975,N_4521);
nand U6145 (N_6145,N_4379,N_4897);
nor U6146 (N_6146,N_3869,N_3802);
xor U6147 (N_6147,N_4400,N_4638);
or U6148 (N_6148,N_3914,N_4329);
nor U6149 (N_6149,N_4817,N_4463);
xor U6150 (N_6150,N_3755,N_3982);
nand U6151 (N_6151,N_4970,N_4219);
nor U6152 (N_6152,N_4266,N_4277);
nand U6153 (N_6153,N_4370,N_4353);
nor U6154 (N_6154,N_4617,N_4499);
nand U6155 (N_6155,N_4413,N_4487);
nor U6156 (N_6156,N_4829,N_4718);
xor U6157 (N_6157,N_4889,N_4328);
nand U6158 (N_6158,N_3767,N_4295);
xnor U6159 (N_6159,N_4146,N_4229);
or U6160 (N_6160,N_4854,N_4843);
nand U6161 (N_6161,N_4357,N_4437);
nand U6162 (N_6162,N_4714,N_3931);
xnor U6163 (N_6163,N_4496,N_4572);
or U6164 (N_6164,N_3790,N_4834);
or U6165 (N_6165,N_4835,N_4014);
xnor U6166 (N_6166,N_3753,N_3830);
nor U6167 (N_6167,N_4264,N_4331);
and U6168 (N_6168,N_4901,N_4221);
nor U6169 (N_6169,N_3844,N_3933);
nand U6170 (N_6170,N_3839,N_4204);
nand U6171 (N_6171,N_4330,N_4136);
nor U6172 (N_6172,N_4872,N_4059);
and U6173 (N_6173,N_3884,N_3941);
xor U6174 (N_6174,N_3970,N_3879);
nand U6175 (N_6175,N_3903,N_4558);
nor U6176 (N_6176,N_4719,N_3864);
xor U6177 (N_6177,N_4491,N_4897);
and U6178 (N_6178,N_4135,N_3995);
and U6179 (N_6179,N_4934,N_4308);
xnor U6180 (N_6180,N_4998,N_4181);
xnor U6181 (N_6181,N_4960,N_4047);
and U6182 (N_6182,N_4046,N_3795);
nand U6183 (N_6183,N_4057,N_4500);
xor U6184 (N_6184,N_4554,N_4551);
xor U6185 (N_6185,N_4098,N_4410);
or U6186 (N_6186,N_4243,N_4698);
nand U6187 (N_6187,N_4121,N_4897);
and U6188 (N_6188,N_4998,N_4517);
nand U6189 (N_6189,N_4330,N_4998);
nor U6190 (N_6190,N_4409,N_3750);
nor U6191 (N_6191,N_4173,N_4589);
nand U6192 (N_6192,N_4280,N_4601);
xor U6193 (N_6193,N_4722,N_4228);
or U6194 (N_6194,N_4819,N_4791);
nor U6195 (N_6195,N_4318,N_4550);
xnor U6196 (N_6196,N_4592,N_4355);
or U6197 (N_6197,N_4860,N_4485);
xnor U6198 (N_6198,N_4386,N_4179);
and U6199 (N_6199,N_4036,N_4068);
nand U6200 (N_6200,N_4893,N_4263);
xnor U6201 (N_6201,N_3756,N_4211);
nand U6202 (N_6202,N_4843,N_4963);
nor U6203 (N_6203,N_4928,N_3860);
or U6204 (N_6204,N_4317,N_4165);
or U6205 (N_6205,N_4425,N_4515);
nand U6206 (N_6206,N_3918,N_4909);
or U6207 (N_6207,N_4044,N_4872);
xnor U6208 (N_6208,N_4724,N_4216);
or U6209 (N_6209,N_4863,N_3806);
or U6210 (N_6210,N_4191,N_3833);
nand U6211 (N_6211,N_4058,N_4176);
nand U6212 (N_6212,N_4974,N_4977);
xnor U6213 (N_6213,N_4780,N_4278);
nor U6214 (N_6214,N_4899,N_3864);
or U6215 (N_6215,N_4472,N_4855);
and U6216 (N_6216,N_4028,N_4320);
or U6217 (N_6217,N_4790,N_4473);
and U6218 (N_6218,N_4835,N_4012);
xor U6219 (N_6219,N_3803,N_4181);
and U6220 (N_6220,N_4697,N_4851);
nand U6221 (N_6221,N_4382,N_4269);
nor U6222 (N_6222,N_3853,N_4416);
nor U6223 (N_6223,N_4520,N_4717);
nor U6224 (N_6224,N_4836,N_3881);
nand U6225 (N_6225,N_4496,N_4332);
and U6226 (N_6226,N_4939,N_4482);
xnor U6227 (N_6227,N_3802,N_4655);
nand U6228 (N_6228,N_4401,N_4383);
xnor U6229 (N_6229,N_4454,N_3992);
and U6230 (N_6230,N_4972,N_4282);
and U6231 (N_6231,N_4854,N_4908);
and U6232 (N_6232,N_4503,N_4917);
nand U6233 (N_6233,N_4455,N_4991);
xor U6234 (N_6234,N_4393,N_4936);
or U6235 (N_6235,N_4287,N_3761);
or U6236 (N_6236,N_4250,N_3867);
nor U6237 (N_6237,N_4609,N_4335);
or U6238 (N_6238,N_3867,N_4192);
xor U6239 (N_6239,N_3845,N_4409);
or U6240 (N_6240,N_4698,N_4383);
and U6241 (N_6241,N_4348,N_3890);
and U6242 (N_6242,N_4224,N_4730);
or U6243 (N_6243,N_4673,N_4761);
nand U6244 (N_6244,N_3947,N_4855);
or U6245 (N_6245,N_4260,N_4098);
nor U6246 (N_6246,N_4490,N_4110);
nor U6247 (N_6247,N_4466,N_4691);
nor U6248 (N_6248,N_3867,N_4220);
and U6249 (N_6249,N_4452,N_4903);
and U6250 (N_6250,N_5113,N_6060);
nand U6251 (N_6251,N_5631,N_6048);
nor U6252 (N_6252,N_5796,N_5763);
or U6253 (N_6253,N_5454,N_5683);
xor U6254 (N_6254,N_6011,N_5692);
or U6255 (N_6255,N_6161,N_5883);
nor U6256 (N_6256,N_5753,N_5147);
nor U6257 (N_6257,N_5643,N_5702);
or U6258 (N_6258,N_5444,N_5350);
and U6259 (N_6259,N_5060,N_5042);
xor U6260 (N_6260,N_6067,N_5292);
nor U6261 (N_6261,N_5899,N_5625);
nand U6262 (N_6262,N_5035,N_5626);
xor U6263 (N_6263,N_6043,N_5485);
or U6264 (N_6264,N_6158,N_5175);
or U6265 (N_6265,N_5975,N_5548);
nand U6266 (N_6266,N_5623,N_6113);
or U6267 (N_6267,N_6170,N_5349);
and U6268 (N_6268,N_5114,N_5351);
or U6269 (N_6269,N_5602,N_5432);
xor U6270 (N_6270,N_5000,N_6036);
and U6271 (N_6271,N_6102,N_5262);
nand U6272 (N_6272,N_5857,N_5322);
xor U6273 (N_6273,N_5335,N_5368);
nor U6274 (N_6274,N_5747,N_6024);
nor U6275 (N_6275,N_5571,N_5270);
nand U6276 (N_6276,N_5544,N_5779);
and U6277 (N_6277,N_5961,N_5674);
or U6278 (N_6278,N_5831,N_5284);
xnor U6279 (N_6279,N_5734,N_5026);
nor U6280 (N_6280,N_5439,N_5204);
nand U6281 (N_6281,N_5810,N_5421);
nor U6282 (N_6282,N_5278,N_5545);
nand U6283 (N_6283,N_5696,N_5888);
and U6284 (N_6284,N_5480,N_5921);
nand U6285 (N_6285,N_5176,N_5312);
nor U6286 (N_6286,N_5789,N_5954);
nor U6287 (N_6287,N_5627,N_5046);
xor U6288 (N_6288,N_5797,N_5572);
or U6289 (N_6289,N_5400,N_5814);
nand U6290 (N_6290,N_5006,N_5091);
or U6291 (N_6291,N_5574,N_5622);
nor U6292 (N_6292,N_5196,N_5890);
nor U6293 (N_6293,N_6079,N_6109);
xnor U6294 (N_6294,N_6042,N_5277);
nand U6295 (N_6295,N_5785,N_5985);
xor U6296 (N_6296,N_5962,N_5952);
nor U6297 (N_6297,N_5908,N_5704);
and U6298 (N_6298,N_6236,N_5462);
and U6299 (N_6299,N_5745,N_5477);
nand U6300 (N_6300,N_5705,N_5461);
nor U6301 (N_6301,N_6146,N_5902);
or U6302 (N_6302,N_5144,N_5467);
and U6303 (N_6303,N_5105,N_5898);
nor U6304 (N_6304,N_5510,N_5654);
xor U6305 (N_6305,N_5458,N_5378);
nor U6306 (N_6306,N_5135,N_5912);
xnor U6307 (N_6307,N_5313,N_5877);
nand U6308 (N_6308,N_5079,N_5728);
xor U6309 (N_6309,N_5443,N_5101);
and U6310 (N_6310,N_5793,N_5275);
nand U6311 (N_6311,N_5129,N_5276);
or U6312 (N_6312,N_5839,N_6132);
nor U6313 (N_6313,N_5494,N_5208);
or U6314 (N_6314,N_5021,N_5542);
nor U6315 (N_6315,N_5562,N_5725);
and U6316 (N_6316,N_6037,N_5846);
and U6317 (N_6317,N_6019,N_6093);
or U6318 (N_6318,N_5509,N_5279);
nand U6319 (N_6319,N_5182,N_5832);
or U6320 (N_6320,N_5288,N_6123);
nand U6321 (N_6321,N_6081,N_5490);
xor U6322 (N_6322,N_5892,N_5629);
nor U6323 (N_6323,N_5223,N_5811);
or U6324 (N_6324,N_5809,N_5450);
and U6325 (N_6325,N_6172,N_5066);
nand U6326 (N_6326,N_5741,N_5382);
nand U6327 (N_6327,N_5404,N_5180);
or U6328 (N_6328,N_5185,N_5521);
and U6329 (N_6329,N_5740,N_6050);
nor U6330 (N_6330,N_6099,N_5259);
or U6331 (N_6331,N_5580,N_5146);
or U6332 (N_6332,N_6182,N_6001);
xnor U6333 (N_6333,N_6226,N_6160);
xnor U6334 (N_6334,N_5198,N_5007);
xnor U6335 (N_6335,N_5413,N_5529);
nand U6336 (N_6336,N_5969,N_5013);
nor U6337 (N_6337,N_5314,N_5511);
and U6338 (N_6338,N_5024,N_5932);
xnor U6339 (N_6339,N_5418,N_5102);
nand U6340 (N_6340,N_5972,N_5257);
nor U6341 (N_6341,N_5910,N_5344);
nand U6342 (N_6342,N_6041,N_5124);
nand U6343 (N_6343,N_5425,N_5286);
xnor U6344 (N_6344,N_5345,N_5547);
nor U6345 (N_6345,N_5800,N_5502);
and U6346 (N_6346,N_5863,N_5836);
or U6347 (N_6347,N_5723,N_6035);
and U6348 (N_6348,N_5229,N_5134);
xnor U6349 (N_6349,N_5078,N_5770);
nand U6350 (N_6350,N_5103,N_5441);
nand U6351 (N_6351,N_5127,N_5923);
or U6352 (N_6352,N_5249,N_6143);
or U6353 (N_6353,N_6125,N_5377);
or U6354 (N_6354,N_5434,N_5804);
or U6355 (N_6355,N_5915,N_5901);
nor U6356 (N_6356,N_5179,N_5009);
and U6357 (N_6357,N_5807,N_5130);
nor U6358 (N_6358,N_6204,N_6090);
and U6359 (N_6359,N_6219,N_6137);
nor U6360 (N_6360,N_5553,N_5104);
xor U6361 (N_6361,N_5436,N_5872);
and U6362 (N_6362,N_5506,N_6030);
or U6363 (N_6363,N_5841,N_6101);
or U6364 (N_6364,N_5080,N_5583);
xnor U6365 (N_6365,N_5946,N_5442);
and U6366 (N_6366,N_5301,N_5758);
xnor U6367 (N_6367,N_5760,N_5659);
xnor U6368 (N_6368,N_5524,N_5755);
nand U6369 (N_6369,N_5522,N_5520);
xor U6370 (N_6370,N_5816,N_5154);
nor U6371 (N_6371,N_5460,N_5268);
and U6372 (N_6372,N_5656,N_5099);
nor U6373 (N_6373,N_6120,N_6175);
xnor U6374 (N_6374,N_5749,N_6085);
or U6375 (N_6375,N_5153,N_5222);
and U6376 (N_6376,N_5483,N_5756);
and U6377 (N_6377,N_5493,N_5448);
nor U6378 (N_6378,N_5107,N_5855);
or U6379 (N_6379,N_5928,N_5210);
nor U6380 (N_6380,N_6179,N_5744);
and U6381 (N_6381,N_5012,N_6197);
or U6382 (N_6382,N_5087,N_5944);
or U6383 (N_6383,N_5355,N_5497);
xor U6384 (N_6384,N_6185,N_5022);
and U6385 (N_6385,N_6045,N_5976);
nand U6386 (N_6386,N_6054,N_5058);
nand U6387 (N_6387,N_5428,N_5539);
and U6388 (N_6388,N_5453,N_6095);
or U6389 (N_6389,N_5711,N_5380);
nor U6390 (N_6390,N_5289,N_6218);
or U6391 (N_6391,N_5295,N_5721);
xor U6392 (N_6392,N_6005,N_5171);
nand U6393 (N_6393,N_5470,N_6063);
xnor U6394 (N_6394,N_5389,N_5260);
nor U6395 (N_6395,N_6248,N_6205);
nand U6396 (N_6396,N_5181,N_5261);
nand U6397 (N_6397,N_6121,N_6243);
and U6398 (N_6398,N_5372,N_5516);
xnor U6399 (N_6399,N_5590,N_5820);
xnor U6400 (N_6400,N_6075,N_5251);
nor U6401 (N_6401,N_5407,N_6070);
or U6402 (N_6402,N_5291,N_5660);
xnor U6403 (N_6403,N_5406,N_5010);
xor U6404 (N_6404,N_5219,N_6114);
nor U6405 (N_6405,N_5423,N_5774);
nand U6406 (N_6406,N_6106,N_5451);
nand U6407 (N_6407,N_5968,N_5849);
and U6408 (N_6408,N_6016,N_5513);
nor U6409 (N_6409,N_5717,N_5430);
or U6410 (N_6410,N_5537,N_5614);
or U6411 (N_6411,N_5033,N_5570);
or U6412 (N_6412,N_5017,N_5854);
or U6413 (N_6413,N_5325,N_5881);
xnor U6414 (N_6414,N_6088,N_6006);
xnor U6415 (N_6415,N_5575,N_5618);
xnor U6416 (N_6416,N_6202,N_6003);
and U6417 (N_6417,N_5665,N_5040);
and U6418 (N_6418,N_5348,N_5212);
nor U6419 (N_6419,N_6163,N_5504);
nand U6420 (N_6420,N_5447,N_5694);
and U6421 (N_6421,N_5764,N_5896);
xor U6422 (N_6422,N_6141,N_5310);
nand U6423 (N_6423,N_5055,N_5194);
nand U6424 (N_6424,N_5853,N_5459);
nand U6425 (N_6425,N_5334,N_5369);
xnor U6426 (N_6426,N_5356,N_5482);
xnor U6427 (N_6427,N_5318,N_5588);
nor U6428 (N_6428,N_5018,N_5746);
or U6429 (N_6429,N_5847,N_5671);
or U6430 (N_6430,N_5907,N_6129);
nor U6431 (N_6431,N_6025,N_5165);
xnor U6432 (N_6432,N_5246,N_5503);
xor U6433 (N_6433,N_5851,N_5403);
xnor U6434 (N_6434,N_6139,N_5609);
xor U6435 (N_6435,N_5294,N_6018);
nand U6436 (N_6436,N_5038,N_5424);
nor U6437 (N_6437,N_5002,N_5422);
and U6438 (N_6438,N_5900,N_5818);
nand U6439 (N_6439,N_5339,N_5027);
or U6440 (N_6440,N_5267,N_5947);
and U6441 (N_6441,N_5940,N_5971);
nand U6442 (N_6442,N_5093,N_5655);
nand U6443 (N_6443,N_5071,N_5752);
and U6444 (N_6444,N_5148,N_6176);
nand U6445 (N_6445,N_6159,N_5801);
nand U6446 (N_6446,N_6191,N_5190);
nand U6447 (N_6447,N_5455,N_5004);
nand U6448 (N_6448,N_5750,N_6015);
nor U6449 (N_6449,N_6216,N_5393);
xor U6450 (N_6450,N_5221,N_6046);
nor U6451 (N_6451,N_5864,N_5668);
nand U6452 (N_6452,N_5767,N_5019);
nor U6453 (N_6453,N_6150,N_5894);
nor U6454 (N_6454,N_5648,N_5199);
nand U6455 (N_6455,N_5645,N_5069);
xor U6456 (N_6456,N_5142,N_5159);
nand U6457 (N_6457,N_5293,N_5925);
or U6458 (N_6458,N_5475,N_5230);
and U6459 (N_6459,N_5346,N_5156);
nand U6460 (N_6460,N_6242,N_5234);
xor U6461 (N_6461,N_5474,N_5476);
nor U6462 (N_6462,N_5433,N_5657);
nand U6463 (N_6463,N_6224,N_5637);
or U6464 (N_6464,N_5938,N_5773);
or U6465 (N_6465,N_5158,N_5535);
xnor U6466 (N_6466,N_5578,N_5446);
and U6467 (N_6467,N_5751,N_5929);
and U6468 (N_6468,N_5576,N_6117);
or U6469 (N_6469,N_5543,N_5712);
and U6470 (N_6470,N_6214,N_5644);
or U6471 (N_6471,N_5769,N_6165);
xor U6472 (N_6472,N_5964,N_5978);
nand U6473 (N_6473,N_5084,N_5560);
xnor U6474 (N_6474,N_5003,N_5664);
and U6475 (N_6475,N_5498,N_5799);
nand U6476 (N_6476,N_5738,N_5517);
or U6477 (N_6477,N_6154,N_5097);
or U6478 (N_6478,N_6166,N_5365);
nor U6479 (N_6479,N_6134,N_5620);
and U6480 (N_6480,N_5170,N_5209);
xor U6481 (N_6481,N_5612,N_5936);
xor U6482 (N_6482,N_5754,N_5466);
and U6483 (N_6483,N_5077,N_6076);
nand U6484 (N_6484,N_6103,N_5601);
nor U6485 (N_6485,N_5473,N_5160);
and U6486 (N_6486,N_5856,N_5265);
xor U6487 (N_6487,N_5036,N_5116);
nor U6488 (N_6488,N_6147,N_5384);
nor U6489 (N_6489,N_5174,N_5586);
nor U6490 (N_6490,N_5667,N_6157);
nand U6491 (N_6491,N_5837,N_5765);
nand U6492 (N_6492,N_6225,N_6174);
and U6493 (N_6493,N_5076,N_5616);
nand U6494 (N_6494,N_5020,N_5039);
xnor U6495 (N_6495,N_5669,N_5743);
or U6496 (N_6496,N_5239,N_6246);
nand U6497 (N_6497,N_5955,N_5970);
or U6498 (N_6498,N_5218,N_5806);
and U6499 (N_6499,N_5998,N_5685);
or U6500 (N_6500,N_6211,N_5280);
xor U6501 (N_6501,N_6116,N_5507);
xor U6502 (N_6502,N_5053,N_5876);
xor U6503 (N_6503,N_6014,N_5508);
and U6504 (N_6504,N_5647,N_5865);
nand U6505 (N_6505,N_5163,N_5942);
xor U6506 (N_6506,N_5487,N_5098);
nor U6507 (N_6507,N_5634,N_5759);
or U6508 (N_6508,N_6039,N_5317);
and U6509 (N_6509,N_5783,N_5850);
nor U6510 (N_6510,N_5787,N_5304);
and U6511 (N_6511,N_5577,N_5869);
nand U6512 (N_6512,N_5109,N_5074);
xor U6513 (N_6513,N_5440,N_5405);
or U6514 (N_6514,N_6020,N_5125);
or U6515 (N_6515,N_5882,N_5981);
xnor U6516 (N_6516,N_5719,N_5603);
and U6517 (N_6517,N_5662,N_5953);
and U6518 (N_6518,N_5893,N_5132);
nand U6519 (N_6519,N_6027,N_5197);
xor U6520 (N_6520,N_5703,N_5370);
or U6521 (N_6521,N_5164,N_5701);
nor U6522 (N_6522,N_5242,N_5757);
nor U6523 (N_6523,N_6002,N_5023);
xor U6524 (N_6524,N_5161,N_5786);
nor U6525 (N_6525,N_5691,N_5227);
or U6526 (N_6526,N_5409,N_5905);
or U6527 (N_6527,N_6056,N_5252);
nand U6528 (N_6528,N_6249,N_5327);
or U6529 (N_6529,N_5730,N_5862);
and U6530 (N_6530,N_5607,N_5306);
or U6531 (N_6531,N_5819,N_5519);
or U6532 (N_6532,N_5067,N_5469);
or U6533 (N_6533,N_6082,N_6124);
xnor U6534 (N_6534,N_5065,N_5488);
and U6535 (N_6535,N_5561,N_5859);
or U6536 (N_6536,N_5646,N_5826);
nor U6537 (N_6537,N_5047,N_6031);
or U6538 (N_6538,N_5481,N_5256);
nor U6539 (N_6539,N_5619,N_5167);
nand U6540 (N_6540,N_5988,N_5889);
xor U6541 (N_6541,N_5059,N_5394);
nor U6542 (N_6542,N_5068,N_5357);
xnor U6543 (N_6543,N_5914,N_5297);
xor U6544 (N_6544,N_5420,N_6119);
or U6545 (N_6545,N_5136,N_5056);
nand U6546 (N_6546,N_6091,N_5670);
nand U6547 (N_6547,N_5429,N_6013);
nor U6548 (N_6548,N_5328,N_5302);
xor U6549 (N_6549,N_5532,N_6084);
nand U6550 (N_6550,N_5780,N_5387);
nand U6551 (N_6551,N_6180,N_5214);
and U6552 (N_6552,N_5546,N_5825);
nand U6553 (N_6553,N_6138,N_5585);
and U6554 (N_6554,N_5299,N_5679);
or U6555 (N_6555,N_6233,N_6089);
xor U6556 (N_6556,N_5120,N_5373);
xnor U6557 (N_6557,N_5792,N_5917);
xor U6558 (N_6558,N_5762,N_5283);
nand U6559 (N_6559,N_6231,N_5188);
and U6560 (N_6560,N_5551,N_5803);
nor U6561 (N_6561,N_6028,N_5639);
nand U6562 (N_6562,N_5641,N_6112);
or U6563 (N_6563,N_5438,N_5965);
xor U6564 (N_6564,N_5282,N_6087);
and U6565 (N_6565,N_6100,N_6122);
nor U6566 (N_6566,N_5922,N_5566);
xnor U6567 (N_6567,N_6128,N_6047);
xnor U6568 (N_6568,N_5977,N_6073);
nor U6569 (N_6569,N_6086,N_6072);
nor U6570 (N_6570,N_5189,N_6133);
nand U6571 (N_6571,N_5139,N_5879);
xor U6572 (N_6572,N_5584,N_6033);
nand U6573 (N_6573,N_5699,N_5296);
and U6574 (N_6574,N_5709,N_6038);
xnor U6575 (N_6575,N_5361,N_6221);
or U6576 (N_6576,N_5737,N_5790);
nand U6577 (N_6577,N_6130,N_6104);
nor U6578 (N_6578,N_5569,N_5123);
and U6579 (N_6579,N_5152,N_5408);
nor U6580 (N_6580,N_6229,N_5943);
nand U6581 (N_6581,N_5332,N_5732);
or U6582 (N_6582,N_5827,N_5540);
nor U6583 (N_6583,N_5070,N_5911);
nand U6584 (N_6584,N_5724,N_5817);
nand U6585 (N_6585,N_5258,N_6156);
nand U6586 (N_6586,N_5595,N_5396);
xor U6587 (N_6587,N_6068,N_5650);
nand U6588 (N_6588,N_6107,N_5383);
nor U6589 (N_6589,N_5984,N_5062);
xnor U6590 (N_6590,N_5842,N_6162);
nand U6591 (N_6591,N_5579,N_5829);
and U6592 (N_6592,N_6186,N_5772);
and U6593 (N_6593,N_5359,N_6203);
nand U6594 (N_6594,N_5303,N_6212);
nor U6595 (N_6595,N_5515,N_5379);
or U6596 (N_6596,N_5815,N_6171);
xor U6597 (N_6597,N_5512,N_5966);
or U6598 (N_6598,N_5761,N_5824);
and U6599 (N_6599,N_5155,N_5329);
or U6600 (N_6600,N_6227,N_5564);
or U6601 (N_6601,N_5178,N_5032);
nor U6602 (N_6602,N_5630,N_5742);
or U6603 (N_6603,N_5948,N_5255);
xor U6604 (N_6604,N_5308,N_5581);
and U6605 (N_6605,N_5162,N_5090);
or U6606 (N_6606,N_5871,N_5845);
nand U6607 (N_6607,N_5933,N_6012);
nand U6608 (N_6608,N_6110,N_5216);
and U6609 (N_6609,N_5813,N_6238);
or U6610 (N_6610,N_5802,N_5464);
xor U6611 (N_6611,N_5395,N_6195);
and U6612 (N_6612,N_6000,N_6052);
xnor U6613 (N_6613,N_5909,N_5633);
xor U6614 (N_6614,N_5126,N_5663);
xnor U6615 (N_6615,N_5203,N_5235);
nor U6616 (N_6616,N_5687,N_5342);
nand U6617 (N_6617,N_5568,N_5926);
or U6618 (N_6618,N_5456,N_6168);
nand U6619 (N_6619,N_5658,N_5200);
xor U6620 (N_6620,N_5727,N_5778);
and U6621 (N_6621,N_5638,N_5768);
and U6622 (N_6622,N_5238,N_5886);
nand U6623 (N_6623,N_5140,N_5011);
nand U6624 (N_6624,N_5353,N_5589);
or U6625 (N_6625,N_5596,N_5360);
and U6626 (N_6626,N_5177,N_5300);
xor U6627 (N_6627,N_5245,N_5224);
xor U6628 (N_6628,N_5573,N_6007);
and U6629 (N_6629,N_5788,N_5064);
xor U6630 (N_6630,N_5552,N_5594);
nand U6631 (N_6631,N_6098,N_6223);
xor U6632 (N_6632,N_5587,N_5145);
nand U6633 (N_6633,N_5617,N_5254);
and U6634 (N_6634,N_5479,N_5731);
and U6635 (N_6635,N_5860,N_5632);
or U6636 (N_6636,N_5324,N_5202);
nor U6637 (N_6637,N_5782,N_5228);
nand U6638 (N_6638,N_5061,N_5514);
or U6639 (N_6639,N_5885,N_5499);
nand U6640 (N_6640,N_6198,N_5031);
xor U6641 (N_6641,N_5949,N_6008);
or U6642 (N_6642,N_5599,N_5613);
and U6643 (N_6643,N_5449,N_5014);
nor U6644 (N_6644,N_5600,N_5821);
nand U6645 (N_6645,N_6144,N_5138);
xnor U6646 (N_6646,N_5094,N_6062);
or U6647 (N_6647,N_5415,N_5822);
nor U6648 (N_6648,N_6239,N_5274);
nor U6649 (N_6649,N_5715,N_5385);
or U6650 (N_6650,N_5973,N_5343);
and U6651 (N_6651,N_5315,N_5285);
or U6652 (N_6652,N_5417,N_5191);
nand U6653 (N_6653,N_5848,N_5858);
or U6654 (N_6654,N_5089,N_5192);
nor U6655 (N_6655,N_5320,N_5615);
or U6656 (N_6656,N_5690,N_5528);
nand U6657 (N_6657,N_5555,N_5939);
or U6658 (N_6658,N_5414,N_5184);
or U6659 (N_6659,N_5592,N_6055);
or U6660 (N_6660,N_5426,N_5941);
nand U6661 (N_6661,N_6234,N_5833);
nor U6662 (N_6662,N_5688,N_5290);
and U6663 (N_6663,N_5452,N_5533);
nor U6664 (N_6664,N_5682,N_5686);
nand U6665 (N_6665,N_5776,N_5591);
xnor U6666 (N_6666,N_5748,N_6058);
xor U6667 (N_6667,N_5963,N_5495);
nand U6668 (N_6668,N_5131,N_5083);
xnor U6669 (N_6669,N_5037,N_5527);
nor U6670 (N_6670,N_6097,N_5427);
or U6671 (N_6671,N_5100,N_5025);
nor U6672 (N_6672,N_5034,N_5672);
and U6673 (N_6673,N_5710,N_6004);
nand U6674 (N_6674,N_5281,N_5726);
nor U6675 (N_6675,N_5677,N_5934);
nand U6676 (N_6676,N_6187,N_5713);
nor U6677 (N_6677,N_5232,N_5247);
nand U6678 (N_6678,N_5416,N_5960);
and U6679 (N_6679,N_5895,N_5500);
or U6680 (N_6680,N_5777,N_5676);
nor U6681 (N_6681,N_5990,N_5410);
and U6682 (N_6682,N_5205,N_5463);
nor U6683 (N_6683,N_5974,N_6145);
xor U6684 (N_6684,N_5844,N_5697);
nor U6685 (N_6685,N_5986,N_5904);
nor U6686 (N_6686,N_5997,N_5693);
or U6687 (N_6687,N_5689,N_6044);
nor U6688 (N_6688,N_5412,N_6164);
xnor U6689 (N_6689,N_5605,N_6064);
xor U6690 (N_6690,N_5891,N_5225);
xor U6691 (N_6691,N_6069,N_5918);
nand U6692 (N_6692,N_6240,N_5491);
xnor U6693 (N_6693,N_6235,N_5331);
nor U6694 (N_6694,N_5995,N_5729);
nor U6695 (N_6695,N_5298,N_5237);
xor U6696 (N_6696,N_5549,N_6148);
or U6697 (N_6697,N_6201,N_6053);
xnor U6698 (N_6698,N_5133,N_5112);
or U6699 (N_6699,N_5471,N_6149);
or U6700 (N_6700,N_5347,N_5606);
nor U6701 (N_6701,N_5501,N_5005);
nand U6702 (N_6702,N_5722,N_5989);
nand U6703 (N_6703,N_5538,N_6142);
nand U6704 (N_6704,N_5598,N_5110);
or U6705 (N_6705,N_5082,N_5927);
nand U6706 (N_6706,N_5051,N_5287);
nand U6707 (N_6707,N_5897,N_5050);
nand U6708 (N_6708,N_5808,N_5128);
and U6709 (N_6709,N_5137,N_6022);
or U6710 (N_6710,N_6220,N_5044);
and U6711 (N_6711,N_5445,N_5736);
nand U6712 (N_6712,N_5358,N_6151);
and U6713 (N_6713,N_5784,N_5830);
nand U6714 (N_6714,N_6111,N_5195);
xor U6715 (N_6715,N_6051,N_5095);
nand U6716 (N_6716,N_5707,N_5582);
xor U6717 (N_6717,N_6115,N_5675);
xor U6718 (N_6718,N_5550,N_5115);
nand U6719 (N_6719,N_6167,N_5075);
nand U6720 (N_6720,N_5367,N_5795);
and U6721 (N_6721,N_5880,N_5534);
and U6722 (N_6722,N_5402,N_5391);
and U6723 (N_6723,N_6094,N_5610);
nor U6724 (N_6724,N_5642,N_5903);
nor U6725 (N_6725,N_5781,N_5472);
and U6726 (N_6726,N_5307,N_5906);
nor U6727 (N_6727,N_5431,N_5653);
or U6728 (N_6728,N_5217,N_5798);
xnor U6729 (N_6729,N_5363,N_5264);
xor U6730 (N_6730,N_5651,N_5706);
nor U6731 (N_6731,N_6199,N_6178);
or U6732 (N_6732,N_5766,N_5266);
and U6733 (N_6733,N_5492,N_6017);
xor U6734 (N_6734,N_5233,N_5805);
and U6735 (N_6735,N_5994,N_5956);
or U6736 (N_6736,N_5340,N_6209);
nand U6737 (N_6737,N_5951,N_5272);
xnor U6738 (N_6738,N_5937,N_6222);
or U6739 (N_6739,N_5371,N_6105);
nor U6740 (N_6740,N_5041,N_5323);
nor U6741 (N_6741,N_5326,N_5484);
xnor U6742 (N_6742,N_5073,N_5118);
and U6743 (N_6743,N_5931,N_5168);
nor U6744 (N_6744,N_5874,N_5680);
and U6745 (N_6745,N_5835,N_5072);
and U6746 (N_6746,N_6206,N_5366);
or U6747 (N_6747,N_6010,N_5673);
or U6748 (N_6748,N_5186,N_5330);
nor U6749 (N_6749,N_5983,N_5193);
xnor U6750 (N_6750,N_5496,N_5187);
or U6751 (N_6751,N_5950,N_6215);
xnor U6752 (N_6752,N_5565,N_5628);
and U6753 (N_6753,N_5250,N_5913);
and U6754 (N_6754,N_5088,N_6177);
and U6755 (N_6755,N_5611,N_5733);
nor U6756 (N_6756,N_6021,N_5958);
nor U6757 (N_6757,N_6009,N_5794);
nand U6758 (N_6758,N_5057,N_6065);
nand U6759 (N_6759,N_5624,N_6181);
nor U6760 (N_6760,N_5838,N_5852);
and U6761 (N_6761,N_5309,N_5119);
or U6762 (N_6762,N_5563,N_6173);
nand U6763 (N_6763,N_5478,N_5341);
or U6764 (N_6764,N_5559,N_5604);
or U6765 (N_6765,N_5437,N_6066);
xnor U6766 (N_6766,N_5401,N_6127);
nor U6767 (N_6767,N_5649,N_5338);
and U6768 (N_6768,N_5244,N_5884);
nand U6769 (N_6769,N_6237,N_5567);
nor U6770 (N_6770,N_5008,N_5530);
or U6771 (N_6771,N_5987,N_5157);
xor U6772 (N_6772,N_5735,N_5999);
xor U6773 (N_6773,N_5086,N_5684);
or U6774 (N_6774,N_6080,N_5333);
nor U6775 (N_6775,N_5980,N_6188);
and U6776 (N_6776,N_5878,N_5957);
xnor U6777 (N_6777,N_6077,N_6241);
nand U6778 (N_6778,N_5718,N_5166);
or U6779 (N_6779,N_5541,N_6245);
and U6780 (N_6780,N_5241,N_5273);
and U6781 (N_6781,N_5708,N_5045);
nand U6782 (N_6782,N_5411,N_5823);
nor U6783 (N_6783,N_5049,N_5593);
nor U6784 (N_6784,N_5678,N_6183);
and U6785 (N_6785,N_5141,N_5812);
nor U6786 (N_6786,N_5868,N_5111);
xnor U6787 (N_6787,N_5263,N_5640);
and U6788 (N_6788,N_5143,N_6152);
or U6789 (N_6789,N_5840,N_5468);
nor U6790 (N_6790,N_5364,N_6213);
and U6791 (N_6791,N_5375,N_5399);
or U6792 (N_6792,N_5398,N_6083);
and U6793 (N_6793,N_5220,N_6118);
and U6794 (N_6794,N_5996,N_6135);
and U6795 (N_6795,N_6193,N_5362);
nand U6796 (N_6796,N_5681,N_5698);
and U6797 (N_6797,N_5390,N_5695);
xor U6798 (N_6798,N_5828,N_5714);
and U6799 (N_6799,N_5875,N_5489);
or U6800 (N_6800,N_5945,N_6126);
xor U6801 (N_6801,N_5661,N_5523);
or U6802 (N_6802,N_5226,N_5666);
nand U6803 (N_6803,N_6140,N_6194);
xnor U6804 (N_6804,N_5392,N_5001);
nand U6805 (N_6805,N_6153,N_5531);
or U6806 (N_6806,N_6217,N_6061);
xnor U6807 (N_6807,N_5397,N_5652);
xnor U6808 (N_6808,N_5621,N_6207);
nor U6809 (N_6809,N_6074,N_5211);
nand U6810 (N_6810,N_5183,N_5419);
xnor U6811 (N_6811,N_6029,N_6034);
xor U6812 (N_6812,N_6190,N_5775);
and U6813 (N_6813,N_5149,N_5096);
and U6814 (N_6814,N_5048,N_5213);
or U6815 (N_6815,N_5015,N_5982);
nand U6816 (N_6816,N_5526,N_5374);
nor U6817 (N_6817,N_5992,N_5321);
xnor U6818 (N_6818,N_5240,N_5376);
nor U6819 (N_6819,N_5556,N_5243);
nand U6820 (N_6820,N_6155,N_6136);
nor U6821 (N_6821,N_5959,N_5030);
or U6822 (N_6822,N_5486,N_6200);
nor U6823 (N_6823,N_5354,N_5108);
xor U6824 (N_6824,N_5597,N_6023);
nor U6825 (N_6825,N_5866,N_6078);
or U6826 (N_6826,N_5720,N_5867);
or U6827 (N_6827,N_5791,N_5554);
xor U6828 (N_6828,N_5993,N_6026);
nor U6829 (N_6829,N_5151,N_6230);
or U6830 (N_6830,N_5924,N_5248);
and U6831 (N_6831,N_5316,N_6131);
or U6832 (N_6832,N_5435,N_5979);
xnor U6833 (N_6833,N_5206,N_5092);
xor U6834 (N_6834,N_5236,N_5207);
xnor U6835 (N_6835,N_5319,N_5930);
and U6836 (N_6836,N_6247,N_5381);
nand U6837 (N_6837,N_6169,N_5231);
or U6838 (N_6838,N_6232,N_5043);
nor U6839 (N_6839,N_6210,N_5608);
nor U6840 (N_6840,N_5150,N_5700);
or U6841 (N_6841,N_5336,N_5536);
or U6842 (N_6842,N_5063,N_5271);
or U6843 (N_6843,N_5935,N_5465);
and U6844 (N_6844,N_5843,N_5305);
nand U6845 (N_6845,N_5919,N_5834);
xnor U6846 (N_6846,N_5081,N_5558);
or U6847 (N_6847,N_5635,N_6196);
xnor U6848 (N_6848,N_5557,N_6059);
and U6849 (N_6849,N_5201,N_5525);
and U6850 (N_6850,N_5636,N_5054);
nor U6851 (N_6851,N_6092,N_5173);
nor U6852 (N_6852,N_6228,N_5028);
nand U6853 (N_6853,N_5457,N_6184);
nor U6854 (N_6854,N_5337,N_5388);
xnor U6855 (N_6855,N_6071,N_5117);
or U6856 (N_6856,N_5920,N_6049);
nand U6857 (N_6857,N_5172,N_5861);
xnor U6858 (N_6858,N_5870,N_5269);
xor U6859 (N_6859,N_5716,N_5518);
xor U6860 (N_6860,N_5771,N_5386);
xnor U6861 (N_6861,N_5169,N_6189);
nand U6862 (N_6862,N_5052,N_5352);
nand U6863 (N_6863,N_6057,N_5215);
nand U6864 (N_6864,N_5991,N_5887);
nand U6865 (N_6865,N_6244,N_6108);
nor U6866 (N_6866,N_5016,N_5253);
xnor U6867 (N_6867,N_6096,N_5505);
or U6868 (N_6868,N_5085,N_5739);
nor U6869 (N_6869,N_5311,N_6208);
nor U6870 (N_6870,N_5106,N_5916);
nand U6871 (N_6871,N_5029,N_6192);
nor U6872 (N_6872,N_6032,N_5122);
or U6873 (N_6873,N_6040,N_5873);
nand U6874 (N_6874,N_5967,N_5121);
or U6875 (N_6875,N_6056,N_5524);
or U6876 (N_6876,N_5180,N_5639);
nor U6877 (N_6877,N_5541,N_5977);
xnor U6878 (N_6878,N_5034,N_5510);
and U6879 (N_6879,N_5891,N_6071);
xor U6880 (N_6880,N_5732,N_5133);
nor U6881 (N_6881,N_5891,N_5415);
or U6882 (N_6882,N_6239,N_5706);
nand U6883 (N_6883,N_5815,N_5216);
and U6884 (N_6884,N_5744,N_5101);
nand U6885 (N_6885,N_5563,N_5077);
nor U6886 (N_6886,N_5762,N_5099);
nor U6887 (N_6887,N_5232,N_6167);
and U6888 (N_6888,N_5062,N_5675);
or U6889 (N_6889,N_5661,N_6088);
nand U6890 (N_6890,N_5048,N_5284);
and U6891 (N_6891,N_6184,N_5583);
nand U6892 (N_6892,N_5042,N_6002);
or U6893 (N_6893,N_5780,N_5722);
or U6894 (N_6894,N_5679,N_5846);
and U6895 (N_6895,N_5957,N_5291);
or U6896 (N_6896,N_5678,N_5460);
nor U6897 (N_6897,N_5651,N_5467);
nand U6898 (N_6898,N_5632,N_5158);
and U6899 (N_6899,N_5441,N_6240);
xor U6900 (N_6900,N_5694,N_6158);
or U6901 (N_6901,N_5067,N_5511);
nand U6902 (N_6902,N_5368,N_5391);
nor U6903 (N_6903,N_5053,N_5995);
or U6904 (N_6904,N_5572,N_5765);
nand U6905 (N_6905,N_5107,N_5727);
nor U6906 (N_6906,N_5750,N_6004);
or U6907 (N_6907,N_5789,N_5810);
nand U6908 (N_6908,N_5068,N_6223);
or U6909 (N_6909,N_6054,N_5263);
nand U6910 (N_6910,N_6170,N_5405);
or U6911 (N_6911,N_5398,N_5224);
or U6912 (N_6912,N_5532,N_5652);
and U6913 (N_6913,N_5251,N_5326);
and U6914 (N_6914,N_5339,N_5710);
or U6915 (N_6915,N_5524,N_5448);
nand U6916 (N_6916,N_5246,N_5120);
nand U6917 (N_6917,N_5361,N_6029);
nor U6918 (N_6918,N_5935,N_5669);
xnor U6919 (N_6919,N_5400,N_5264);
and U6920 (N_6920,N_6076,N_6245);
and U6921 (N_6921,N_5111,N_6208);
nand U6922 (N_6922,N_5339,N_5305);
or U6923 (N_6923,N_5961,N_5920);
xor U6924 (N_6924,N_5328,N_5782);
nand U6925 (N_6925,N_5581,N_5813);
xor U6926 (N_6926,N_5711,N_5363);
nor U6927 (N_6927,N_5740,N_5515);
nand U6928 (N_6928,N_5756,N_5609);
or U6929 (N_6929,N_5909,N_5461);
nor U6930 (N_6930,N_5636,N_5159);
nor U6931 (N_6931,N_5420,N_5433);
and U6932 (N_6932,N_5825,N_5762);
nor U6933 (N_6933,N_5580,N_5327);
and U6934 (N_6934,N_5800,N_5150);
nor U6935 (N_6935,N_5219,N_5747);
and U6936 (N_6936,N_5153,N_5969);
or U6937 (N_6937,N_5344,N_5620);
or U6938 (N_6938,N_5627,N_6040);
and U6939 (N_6939,N_6188,N_5134);
nor U6940 (N_6940,N_5813,N_5668);
or U6941 (N_6941,N_5262,N_5542);
nor U6942 (N_6942,N_5476,N_6010);
nor U6943 (N_6943,N_6030,N_6084);
nand U6944 (N_6944,N_6205,N_5817);
nor U6945 (N_6945,N_5447,N_6149);
xor U6946 (N_6946,N_5746,N_5001);
xnor U6947 (N_6947,N_5507,N_5488);
or U6948 (N_6948,N_5316,N_6049);
nand U6949 (N_6949,N_6078,N_5960);
or U6950 (N_6950,N_5489,N_5814);
xor U6951 (N_6951,N_5812,N_5795);
nand U6952 (N_6952,N_5761,N_6057);
xnor U6953 (N_6953,N_6156,N_5458);
or U6954 (N_6954,N_5419,N_5630);
nand U6955 (N_6955,N_5705,N_5623);
nand U6956 (N_6956,N_5986,N_5730);
nor U6957 (N_6957,N_5986,N_5495);
or U6958 (N_6958,N_5619,N_6218);
or U6959 (N_6959,N_5016,N_5607);
and U6960 (N_6960,N_5385,N_5184);
or U6961 (N_6961,N_5164,N_5557);
nor U6962 (N_6962,N_5010,N_5613);
nor U6963 (N_6963,N_5636,N_6102);
xnor U6964 (N_6964,N_5479,N_6236);
and U6965 (N_6965,N_5569,N_5469);
or U6966 (N_6966,N_5711,N_5427);
and U6967 (N_6967,N_5173,N_5134);
xor U6968 (N_6968,N_5082,N_5197);
and U6969 (N_6969,N_5242,N_5878);
xnor U6970 (N_6970,N_5684,N_5190);
or U6971 (N_6971,N_5365,N_5566);
and U6972 (N_6972,N_6149,N_5883);
nand U6973 (N_6973,N_5024,N_5036);
nor U6974 (N_6974,N_5413,N_6190);
and U6975 (N_6975,N_5886,N_5680);
or U6976 (N_6976,N_5056,N_5656);
nand U6977 (N_6977,N_5602,N_6099);
or U6978 (N_6978,N_6068,N_6184);
or U6979 (N_6979,N_5601,N_5099);
nand U6980 (N_6980,N_5096,N_6217);
nand U6981 (N_6981,N_5547,N_5365);
nor U6982 (N_6982,N_6195,N_5058);
or U6983 (N_6983,N_5184,N_5127);
xnor U6984 (N_6984,N_5058,N_5337);
xor U6985 (N_6985,N_5061,N_5671);
or U6986 (N_6986,N_5141,N_5319);
nand U6987 (N_6987,N_5316,N_6164);
and U6988 (N_6988,N_6188,N_6015);
xnor U6989 (N_6989,N_5108,N_6047);
and U6990 (N_6990,N_5725,N_5090);
nor U6991 (N_6991,N_5751,N_5198);
nand U6992 (N_6992,N_5318,N_5077);
or U6993 (N_6993,N_5554,N_5649);
nor U6994 (N_6994,N_6217,N_5311);
nand U6995 (N_6995,N_5385,N_6221);
or U6996 (N_6996,N_5035,N_5392);
nand U6997 (N_6997,N_5824,N_5703);
nand U6998 (N_6998,N_5386,N_6085);
nor U6999 (N_6999,N_6233,N_5988);
and U7000 (N_7000,N_5251,N_5110);
and U7001 (N_7001,N_6222,N_5810);
nand U7002 (N_7002,N_5341,N_5550);
or U7003 (N_7003,N_5987,N_5552);
or U7004 (N_7004,N_5127,N_5677);
nand U7005 (N_7005,N_6039,N_5951);
or U7006 (N_7006,N_6018,N_5848);
and U7007 (N_7007,N_5233,N_5190);
nor U7008 (N_7008,N_5039,N_5785);
and U7009 (N_7009,N_5434,N_5985);
nand U7010 (N_7010,N_5487,N_6066);
and U7011 (N_7011,N_5753,N_5792);
xor U7012 (N_7012,N_5464,N_5189);
xor U7013 (N_7013,N_5681,N_5769);
xor U7014 (N_7014,N_6167,N_6231);
and U7015 (N_7015,N_6155,N_5068);
and U7016 (N_7016,N_5093,N_5836);
xnor U7017 (N_7017,N_5516,N_5487);
or U7018 (N_7018,N_5190,N_6081);
or U7019 (N_7019,N_5792,N_5500);
xnor U7020 (N_7020,N_5524,N_5039);
nand U7021 (N_7021,N_5764,N_6060);
xor U7022 (N_7022,N_5071,N_5282);
xor U7023 (N_7023,N_6183,N_5556);
xnor U7024 (N_7024,N_5266,N_5134);
nand U7025 (N_7025,N_6154,N_5274);
xor U7026 (N_7026,N_5771,N_6200);
nand U7027 (N_7027,N_5353,N_5189);
xor U7028 (N_7028,N_5573,N_6231);
and U7029 (N_7029,N_5042,N_5926);
and U7030 (N_7030,N_5796,N_5498);
nor U7031 (N_7031,N_5492,N_6065);
and U7032 (N_7032,N_5023,N_5118);
nor U7033 (N_7033,N_5943,N_5833);
or U7034 (N_7034,N_5751,N_5710);
nor U7035 (N_7035,N_5747,N_5788);
or U7036 (N_7036,N_5118,N_5212);
nor U7037 (N_7037,N_5180,N_5268);
or U7038 (N_7038,N_5772,N_5629);
xor U7039 (N_7039,N_5328,N_5122);
and U7040 (N_7040,N_5515,N_5105);
nand U7041 (N_7041,N_5972,N_5250);
and U7042 (N_7042,N_5880,N_5515);
and U7043 (N_7043,N_6191,N_5268);
or U7044 (N_7044,N_5370,N_6048);
xnor U7045 (N_7045,N_5265,N_5759);
nor U7046 (N_7046,N_5273,N_5829);
and U7047 (N_7047,N_5837,N_6206);
xor U7048 (N_7048,N_5331,N_5364);
nor U7049 (N_7049,N_5397,N_5733);
nand U7050 (N_7050,N_5153,N_5653);
or U7051 (N_7051,N_5391,N_5804);
or U7052 (N_7052,N_6159,N_5945);
nand U7053 (N_7053,N_5096,N_5125);
and U7054 (N_7054,N_5513,N_6146);
nor U7055 (N_7055,N_5550,N_5329);
and U7056 (N_7056,N_5475,N_5675);
xnor U7057 (N_7057,N_6034,N_5971);
nand U7058 (N_7058,N_6080,N_5374);
xor U7059 (N_7059,N_5088,N_5963);
nor U7060 (N_7060,N_5349,N_6135);
nand U7061 (N_7061,N_5453,N_5607);
nor U7062 (N_7062,N_5635,N_5922);
and U7063 (N_7063,N_6019,N_5716);
nand U7064 (N_7064,N_5821,N_5251);
nor U7065 (N_7065,N_5995,N_5919);
and U7066 (N_7066,N_5286,N_5188);
and U7067 (N_7067,N_5837,N_5990);
or U7068 (N_7068,N_5391,N_6080);
xnor U7069 (N_7069,N_6087,N_5966);
or U7070 (N_7070,N_5970,N_5046);
and U7071 (N_7071,N_5583,N_5994);
and U7072 (N_7072,N_5424,N_5040);
nand U7073 (N_7073,N_6075,N_6171);
xnor U7074 (N_7074,N_5459,N_6209);
or U7075 (N_7075,N_5969,N_5858);
nor U7076 (N_7076,N_5210,N_5539);
nand U7077 (N_7077,N_6159,N_5608);
xnor U7078 (N_7078,N_5592,N_5427);
and U7079 (N_7079,N_5476,N_5776);
and U7080 (N_7080,N_5356,N_5854);
nand U7081 (N_7081,N_5087,N_5219);
xnor U7082 (N_7082,N_5805,N_5909);
nand U7083 (N_7083,N_5399,N_5068);
nand U7084 (N_7084,N_5321,N_5312);
or U7085 (N_7085,N_5218,N_5713);
xnor U7086 (N_7086,N_5009,N_6115);
and U7087 (N_7087,N_5645,N_5164);
nor U7088 (N_7088,N_5012,N_5548);
or U7089 (N_7089,N_5955,N_5939);
xnor U7090 (N_7090,N_5160,N_6116);
or U7091 (N_7091,N_5697,N_6220);
nor U7092 (N_7092,N_5781,N_5524);
nor U7093 (N_7093,N_6052,N_6074);
nand U7094 (N_7094,N_5642,N_5704);
or U7095 (N_7095,N_6037,N_5588);
or U7096 (N_7096,N_5400,N_5394);
xor U7097 (N_7097,N_5664,N_6239);
or U7098 (N_7098,N_6110,N_5579);
xor U7099 (N_7099,N_5610,N_5857);
and U7100 (N_7100,N_5709,N_5107);
xnor U7101 (N_7101,N_6218,N_5048);
nor U7102 (N_7102,N_5437,N_5421);
and U7103 (N_7103,N_5747,N_5458);
and U7104 (N_7104,N_5545,N_5512);
xnor U7105 (N_7105,N_5886,N_5306);
or U7106 (N_7106,N_5738,N_5271);
xor U7107 (N_7107,N_5232,N_6040);
nor U7108 (N_7108,N_6205,N_5029);
and U7109 (N_7109,N_5815,N_5396);
nor U7110 (N_7110,N_6050,N_6108);
nor U7111 (N_7111,N_5309,N_5301);
nor U7112 (N_7112,N_6057,N_6245);
and U7113 (N_7113,N_5737,N_5677);
and U7114 (N_7114,N_5374,N_5890);
xnor U7115 (N_7115,N_5904,N_5683);
nor U7116 (N_7116,N_6020,N_6190);
or U7117 (N_7117,N_5506,N_5702);
or U7118 (N_7118,N_6150,N_6088);
or U7119 (N_7119,N_5977,N_5007);
and U7120 (N_7120,N_5254,N_5459);
nand U7121 (N_7121,N_5317,N_5505);
xnor U7122 (N_7122,N_5906,N_5441);
nor U7123 (N_7123,N_5259,N_6105);
xnor U7124 (N_7124,N_6244,N_5691);
or U7125 (N_7125,N_5645,N_5305);
and U7126 (N_7126,N_5468,N_6162);
xnor U7127 (N_7127,N_5549,N_5646);
or U7128 (N_7128,N_5176,N_5578);
nor U7129 (N_7129,N_5568,N_5428);
xnor U7130 (N_7130,N_6114,N_5403);
xnor U7131 (N_7131,N_5663,N_5232);
and U7132 (N_7132,N_5951,N_5931);
nand U7133 (N_7133,N_5094,N_5180);
and U7134 (N_7134,N_5216,N_5257);
and U7135 (N_7135,N_5884,N_6108);
or U7136 (N_7136,N_5835,N_5579);
xor U7137 (N_7137,N_5051,N_5358);
nor U7138 (N_7138,N_5059,N_5381);
nor U7139 (N_7139,N_5097,N_5508);
or U7140 (N_7140,N_5524,N_5897);
nand U7141 (N_7141,N_5882,N_5617);
and U7142 (N_7142,N_5281,N_5440);
or U7143 (N_7143,N_5633,N_5002);
nor U7144 (N_7144,N_5823,N_5875);
and U7145 (N_7145,N_5506,N_5061);
or U7146 (N_7146,N_5848,N_5759);
nand U7147 (N_7147,N_5149,N_5813);
and U7148 (N_7148,N_5536,N_6110);
and U7149 (N_7149,N_5626,N_5539);
or U7150 (N_7150,N_5789,N_5816);
or U7151 (N_7151,N_5299,N_5977);
or U7152 (N_7152,N_5387,N_6047);
nand U7153 (N_7153,N_5576,N_5670);
or U7154 (N_7154,N_5851,N_5146);
nor U7155 (N_7155,N_5201,N_5788);
nand U7156 (N_7156,N_5341,N_5304);
xor U7157 (N_7157,N_5097,N_5902);
nor U7158 (N_7158,N_5209,N_5537);
or U7159 (N_7159,N_5371,N_5365);
or U7160 (N_7160,N_6037,N_6078);
nor U7161 (N_7161,N_5826,N_5551);
and U7162 (N_7162,N_5725,N_5475);
nor U7163 (N_7163,N_6093,N_5151);
nor U7164 (N_7164,N_5489,N_5322);
nor U7165 (N_7165,N_5726,N_6175);
xnor U7166 (N_7166,N_5317,N_5452);
xor U7167 (N_7167,N_5714,N_6167);
nand U7168 (N_7168,N_6249,N_5481);
nor U7169 (N_7169,N_5368,N_5233);
or U7170 (N_7170,N_6141,N_5094);
xor U7171 (N_7171,N_5465,N_5779);
nand U7172 (N_7172,N_5864,N_5259);
xnor U7173 (N_7173,N_5785,N_5889);
or U7174 (N_7174,N_5049,N_5093);
or U7175 (N_7175,N_5107,N_5274);
nor U7176 (N_7176,N_5588,N_5552);
nand U7177 (N_7177,N_5636,N_5526);
and U7178 (N_7178,N_5183,N_5891);
xnor U7179 (N_7179,N_6063,N_5437);
or U7180 (N_7180,N_6229,N_5048);
nor U7181 (N_7181,N_5309,N_5224);
nand U7182 (N_7182,N_5514,N_5342);
or U7183 (N_7183,N_5979,N_5658);
or U7184 (N_7184,N_5568,N_6205);
xnor U7185 (N_7185,N_5554,N_5988);
xnor U7186 (N_7186,N_5833,N_6009);
nor U7187 (N_7187,N_5718,N_5335);
nand U7188 (N_7188,N_6138,N_6139);
xor U7189 (N_7189,N_5638,N_6083);
xor U7190 (N_7190,N_5234,N_5052);
xor U7191 (N_7191,N_5241,N_5366);
nand U7192 (N_7192,N_5954,N_5936);
nand U7193 (N_7193,N_5858,N_6011);
nor U7194 (N_7194,N_5610,N_5364);
nand U7195 (N_7195,N_5580,N_5621);
nand U7196 (N_7196,N_6140,N_5877);
nand U7197 (N_7197,N_5495,N_5520);
xnor U7198 (N_7198,N_5521,N_5156);
nand U7199 (N_7199,N_5096,N_5234);
nand U7200 (N_7200,N_5558,N_5697);
nand U7201 (N_7201,N_5847,N_5403);
and U7202 (N_7202,N_5746,N_5034);
and U7203 (N_7203,N_5538,N_5740);
or U7204 (N_7204,N_5989,N_5138);
or U7205 (N_7205,N_5823,N_5568);
and U7206 (N_7206,N_5621,N_5432);
nand U7207 (N_7207,N_6111,N_5012);
nor U7208 (N_7208,N_5673,N_5180);
nor U7209 (N_7209,N_5221,N_6174);
and U7210 (N_7210,N_6145,N_5060);
nand U7211 (N_7211,N_5353,N_5611);
and U7212 (N_7212,N_5663,N_5042);
xnor U7213 (N_7213,N_5634,N_5561);
xor U7214 (N_7214,N_5032,N_5499);
nand U7215 (N_7215,N_6209,N_5973);
or U7216 (N_7216,N_5013,N_5463);
xor U7217 (N_7217,N_5495,N_6050);
or U7218 (N_7218,N_5646,N_5719);
or U7219 (N_7219,N_5662,N_6222);
or U7220 (N_7220,N_5803,N_5647);
or U7221 (N_7221,N_5250,N_6057);
xor U7222 (N_7222,N_5415,N_5907);
or U7223 (N_7223,N_5938,N_6074);
nor U7224 (N_7224,N_5758,N_6041);
nand U7225 (N_7225,N_5213,N_5551);
nand U7226 (N_7226,N_5048,N_5339);
xor U7227 (N_7227,N_5697,N_5497);
nand U7228 (N_7228,N_5497,N_5763);
or U7229 (N_7229,N_6070,N_5227);
or U7230 (N_7230,N_6034,N_6060);
nor U7231 (N_7231,N_5744,N_5381);
or U7232 (N_7232,N_5587,N_5840);
and U7233 (N_7233,N_6151,N_5919);
xor U7234 (N_7234,N_6004,N_6074);
nor U7235 (N_7235,N_5325,N_6142);
nor U7236 (N_7236,N_5747,N_5420);
nor U7237 (N_7237,N_6220,N_5310);
or U7238 (N_7238,N_5095,N_5920);
xnor U7239 (N_7239,N_5983,N_6098);
nand U7240 (N_7240,N_5261,N_5768);
nor U7241 (N_7241,N_6066,N_5497);
xor U7242 (N_7242,N_5520,N_6196);
and U7243 (N_7243,N_5935,N_5365);
xor U7244 (N_7244,N_5069,N_5544);
nand U7245 (N_7245,N_5111,N_5973);
or U7246 (N_7246,N_5305,N_5992);
nor U7247 (N_7247,N_5693,N_6032);
and U7248 (N_7248,N_5534,N_6073);
nor U7249 (N_7249,N_5922,N_5061);
or U7250 (N_7250,N_6012,N_5649);
or U7251 (N_7251,N_5177,N_5955);
and U7252 (N_7252,N_5864,N_6219);
nor U7253 (N_7253,N_5458,N_5060);
xor U7254 (N_7254,N_5823,N_6060);
and U7255 (N_7255,N_5780,N_5333);
xor U7256 (N_7256,N_5717,N_6026);
nand U7257 (N_7257,N_5669,N_5588);
and U7258 (N_7258,N_5075,N_5277);
nand U7259 (N_7259,N_5498,N_5284);
nor U7260 (N_7260,N_5992,N_5452);
nand U7261 (N_7261,N_5903,N_5019);
or U7262 (N_7262,N_5480,N_5115);
or U7263 (N_7263,N_5546,N_5922);
or U7264 (N_7264,N_6204,N_5025);
xor U7265 (N_7265,N_5656,N_5577);
and U7266 (N_7266,N_5756,N_5021);
and U7267 (N_7267,N_5055,N_5789);
nand U7268 (N_7268,N_5996,N_6248);
and U7269 (N_7269,N_5881,N_6217);
nor U7270 (N_7270,N_5656,N_5971);
and U7271 (N_7271,N_5721,N_5168);
and U7272 (N_7272,N_6050,N_5634);
nor U7273 (N_7273,N_5925,N_5372);
nor U7274 (N_7274,N_5734,N_5520);
nor U7275 (N_7275,N_5670,N_6097);
nor U7276 (N_7276,N_5016,N_5936);
nand U7277 (N_7277,N_5912,N_5292);
xor U7278 (N_7278,N_5002,N_5909);
nor U7279 (N_7279,N_5484,N_6204);
nand U7280 (N_7280,N_5342,N_5915);
nand U7281 (N_7281,N_5328,N_5786);
xor U7282 (N_7282,N_5345,N_5665);
nor U7283 (N_7283,N_5561,N_5345);
or U7284 (N_7284,N_5500,N_5197);
and U7285 (N_7285,N_5175,N_5915);
nor U7286 (N_7286,N_5895,N_5387);
xnor U7287 (N_7287,N_5168,N_5405);
nor U7288 (N_7288,N_5877,N_6039);
or U7289 (N_7289,N_6238,N_5103);
and U7290 (N_7290,N_5784,N_5218);
nand U7291 (N_7291,N_6216,N_5107);
xnor U7292 (N_7292,N_5767,N_6030);
nor U7293 (N_7293,N_5198,N_5897);
nand U7294 (N_7294,N_5355,N_6000);
xnor U7295 (N_7295,N_5466,N_5762);
and U7296 (N_7296,N_6081,N_5164);
nor U7297 (N_7297,N_6136,N_5699);
nand U7298 (N_7298,N_5121,N_5640);
nor U7299 (N_7299,N_5881,N_5830);
xor U7300 (N_7300,N_5093,N_5701);
nor U7301 (N_7301,N_6044,N_5361);
nand U7302 (N_7302,N_5733,N_6057);
and U7303 (N_7303,N_5790,N_6153);
nor U7304 (N_7304,N_5391,N_5162);
nand U7305 (N_7305,N_5533,N_5325);
nor U7306 (N_7306,N_6156,N_5001);
nand U7307 (N_7307,N_6117,N_5639);
xor U7308 (N_7308,N_5635,N_5552);
and U7309 (N_7309,N_6126,N_6101);
xnor U7310 (N_7310,N_5917,N_5848);
nand U7311 (N_7311,N_6138,N_5308);
nor U7312 (N_7312,N_5546,N_5703);
xnor U7313 (N_7313,N_5449,N_6038);
xnor U7314 (N_7314,N_6076,N_5076);
xnor U7315 (N_7315,N_5662,N_6172);
xor U7316 (N_7316,N_6065,N_5263);
nand U7317 (N_7317,N_6115,N_6017);
nand U7318 (N_7318,N_5595,N_5269);
xor U7319 (N_7319,N_5294,N_6159);
and U7320 (N_7320,N_5561,N_5616);
nor U7321 (N_7321,N_5259,N_5109);
nand U7322 (N_7322,N_5772,N_6017);
and U7323 (N_7323,N_5832,N_5774);
nand U7324 (N_7324,N_5925,N_5864);
nor U7325 (N_7325,N_5125,N_5683);
and U7326 (N_7326,N_5888,N_5795);
or U7327 (N_7327,N_5194,N_5514);
nand U7328 (N_7328,N_5357,N_5621);
xor U7329 (N_7329,N_5685,N_5780);
or U7330 (N_7330,N_5745,N_5865);
xnor U7331 (N_7331,N_5533,N_5891);
nor U7332 (N_7332,N_5161,N_6009);
nor U7333 (N_7333,N_5282,N_5822);
nor U7334 (N_7334,N_6233,N_5351);
or U7335 (N_7335,N_5395,N_6085);
xor U7336 (N_7336,N_5728,N_5659);
nor U7337 (N_7337,N_5897,N_5680);
or U7338 (N_7338,N_5967,N_5998);
xnor U7339 (N_7339,N_5287,N_5313);
nor U7340 (N_7340,N_5527,N_5695);
nor U7341 (N_7341,N_5547,N_5954);
and U7342 (N_7342,N_5719,N_5648);
or U7343 (N_7343,N_5817,N_5226);
and U7344 (N_7344,N_5429,N_5904);
nand U7345 (N_7345,N_5911,N_6172);
and U7346 (N_7346,N_5548,N_5239);
and U7347 (N_7347,N_5866,N_5427);
or U7348 (N_7348,N_5727,N_6101);
xnor U7349 (N_7349,N_5723,N_5185);
xnor U7350 (N_7350,N_5102,N_6101);
nand U7351 (N_7351,N_5663,N_5535);
nand U7352 (N_7352,N_5361,N_5685);
xnor U7353 (N_7353,N_5756,N_5247);
and U7354 (N_7354,N_5276,N_5306);
or U7355 (N_7355,N_5845,N_5882);
nor U7356 (N_7356,N_6218,N_5033);
nand U7357 (N_7357,N_5629,N_6034);
xor U7358 (N_7358,N_6131,N_5011);
xnor U7359 (N_7359,N_5663,N_5960);
or U7360 (N_7360,N_5645,N_5374);
or U7361 (N_7361,N_6094,N_5773);
or U7362 (N_7362,N_5168,N_5068);
nand U7363 (N_7363,N_6062,N_5231);
or U7364 (N_7364,N_5410,N_5291);
and U7365 (N_7365,N_5800,N_5342);
nor U7366 (N_7366,N_6158,N_5608);
xor U7367 (N_7367,N_5123,N_6040);
nand U7368 (N_7368,N_5267,N_6134);
xnor U7369 (N_7369,N_6154,N_6121);
xor U7370 (N_7370,N_5623,N_5941);
or U7371 (N_7371,N_5109,N_5219);
xor U7372 (N_7372,N_5510,N_6041);
nor U7373 (N_7373,N_5105,N_5368);
nor U7374 (N_7374,N_6192,N_5892);
nor U7375 (N_7375,N_5527,N_5045);
or U7376 (N_7376,N_5127,N_6205);
xnor U7377 (N_7377,N_6164,N_6119);
and U7378 (N_7378,N_5402,N_6063);
nor U7379 (N_7379,N_5622,N_5609);
nor U7380 (N_7380,N_6226,N_5127);
or U7381 (N_7381,N_5109,N_6082);
nand U7382 (N_7382,N_6239,N_5707);
nand U7383 (N_7383,N_5671,N_6027);
and U7384 (N_7384,N_5121,N_6217);
or U7385 (N_7385,N_6233,N_5272);
nand U7386 (N_7386,N_6035,N_5625);
nor U7387 (N_7387,N_5955,N_5155);
nand U7388 (N_7388,N_6073,N_5757);
xnor U7389 (N_7389,N_6061,N_5255);
xnor U7390 (N_7390,N_5109,N_6078);
and U7391 (N_7391,N_5832,N_6156);
xor U7392 (N_7392,N_5481,N_5032);
nand U7393 (N_7393,N_5730,N_6243);
nor U7394 (N_7394,N_6157,N_5317);
and U7395 (N_7395,N_6139,N_5431);
nor U7396 (N_7396,N_5068,N_5446);
nor U7397 (N_7397,N_5579,N_5009);
nor U7398 (N_7398,N_5629,N_6191);
nor U7399 (N_7399,N_6041,N_5304);
xor U7400 (N_7400,N_6148,N_5048);
xor U7401 (N_7401,N_5259,N_5410);
nor U7402 (N_7402,N_6173,N_5800);
or U7403 (N_7403,N_5857,N_5972);
xor U7404 (N_7404,N_5074,N_5188);
nor U7405 (N_7405,N_5959,N_5904);
nor U7406 (N_7406,N_6188,N_6136);
nor U7407 (N_7407,N_5936,N_6126);
or U7408 (N_7408,N_6204,N_6092);
xnor U7409 (N_7409,N_6095,N_6183);
xnor U7410 (N_7410,N_5576,N_5940);
nor U7411 (N_7411,N_5937,N_5932);
or U7412 (N_7412,N_5007,N_6229);
xor U7413 (N_7413,N_5289,N_5501);
nor U7414 (N_7414,N_5881,N_5390);
nand U7415 (N_7415,N_5550,N_5978);
or U7416 (N_7416,N_6240,N_5932);
or U7417 (N_7417,N_5949,N_5110);
nand U7418 (N_7418,N_5811,N_5222);
nor U7419 (N_7419,N_5901,N_5110);
and U7420 (N_7420,N_6175,N_5495);
nand U7421 (N_7421,N_6146,N_5670);
nand U7422 (N_7422,N_6146,N_5380);
and U7423 (N_7423,N_5731,N_5976);
nand U7424 (N_7424,N_5845,N_5247);
nor U7425 (N_7425,N_5919,N_5898);
nor U7426 (N_7426,N_5437,N_6219);
nor U7427 (N_7427,N_5718,N_5269);
or U7428 (N_7428,N_5879,N_6095);
and U7429 (N_7429,N_6210,N_5028);
nand U7430 (N_7430,N_5642,N_6154);
nand U7431 (N_7431,N_5143,N_5967);
nand U7432 (N_7432,N_6116,N_5258);
xor U7433 (N_7433,N_6084,N_5372);
or U7434 (N_7434,N_5365,N_5807);
nor U7435 (N_7435,N_5554,N_5371);
or U7436 (N_7436,N_5446,N_5631);
or U7437 (N_7437,N_5525,N_5328);
nand U7438 (N_7438,N_5513,N_5691);
and U7439 (N_7439,N_5072,N_5290);
or U7440 (N_7440,N_5024,N_5153);
or U7441 (N_7441,N_6230,N_5464);
xor U7442 (N_7442,N_5835,N_5319);
nand U7443 (N_7443,N_5748,N_6035);
nand U7444 (N_7444,N_6142,N_5341);
nand U7445 (N_7445,N_6160,N_5482);
or U7446 (N_7446,N_5716,N_6171);
nand U7447 (N_7447,N_5541,N_5836);
nor U7448 (N_7448,N_5507,N_5694);
or U7449 (N_7449,N_6205,N_5558);
and U7450 (N_7450,N_5553,N_5528);
nand U7451 (N_7451,N_5804,N_5759);
or U7452 (N_7452,N_5906,N_6182);
nor U7453 (N_7453,N_5365,N_6176);
or U7454 (N_7454,N_6021,N_5585);
xnor U7455 (N_7455,N_5421,N_5427);
or U7456 (N_7456,N_5884,N_6227);
nand U7457 (N_7457,N_5707,N_5655);
nand U7458 (N_7458,N_5830,N_5381);
or U7459 (N_7459,N_5123,N_5574);
nor U7460 (N_7460,N_5581,N_5958);
xnor U7461 (N_7461,N_5396,N_5602);
nand U7462 (N_7462,N_5424,N_5549);
xnor U7463 (N_7463,N_5250,N_5066);
xor U7464 (N_7464,N_5454,N_6236);
and U7465 (N_7465,N_5771,N_6067);
or U7466 (N_7466,N_5991,N_5742);
and U7467 (N_7467,N_6223,N_5044);
nor U7468 (N_7468,N_5832,N_5149);
nand U7469 (N_7469,N_6075,N_5254);
and U7470 (N_7470,N_5007,N_5695);
nand U7471 (N_7471,N_5844,N_5543);
nor U7472 (N_7472,N_5232,N_5962);
nand U7473 (N_7473,N_5144,N_5367);
nor U7474 (N_7474,N_6024,N_5918);
or U7475 (N_7475,N_5136,N_5755);
xor U7476 (N_7476,N_6174,N_5829);
or U7477 (N_7477,N_5539,N_5219);
nor U7478 (N_7478,N_6122,N_5039);
nor U7479 (N_7479,N_5807,N_5329);
and U7480 (N_7480,N_6102,N_5208);
and U7481 (N_7481,N_5624,N_5035);
and U7482 (N_7482,N_5827,N_5136);
nand U7483 (N_7483,N_5563,N_5844);
nand U7484 (N_7484,N_6187,N_6075);
nor U7485 (N_7485,N_5790,N_6242);
and U7486 (N_7486,N_5260,N_5086);
nor U7487 (N_7487,N_5678,N_5005);
nor U7488 (N_7488,N_5716,N_5496);
and U7489 (N_7489,N_5655,N_5366);
nor U7490 (N_7490,N_5426,N_5967);
xor U7491 (N_7491,N_5919,N_5251);
nor U7492 (N_7492,N_5558,N_5465);
or U7493 (N_7493,N_5607,N_6131);
or U7494 (N_7494,N_5712,N_5610);
nor U7495 (N_7495,N_6094,N_5735);
and U7496 (N_7496,N_5412,N_5184);
nor U7497 (N_7497,N_5266,N_5442);
or U7498 (N_7498,N_5482,N_5652);
nor U7499 (N_7499,N_5914,N_5152);
or U7500 (N_7500,N_6383,N_6650);
nand U7501 (N_7501,N_6276,N_6559);
xnor U7502 (N_7502,N_6342,N_7208);
and U7503 (N_7503,N_7349,N_6845);
xnor U7504 (N_7504,N_7047,N_7133);
nand U7505 (N_7505,N_6995,N_6493);
or U7506 (N_7506,N_6347,N_6320);
and U7507 (N_7507,N_7335,N_6973);
and U7508 (N_7508,N_7112,N_7196);
xnor U7509 (N_7509,N_7444,N_6808);
xnor U7510 (N_7510,N_7392,N_6687);
nand U7511 (N_7511,N_7316,N_6552);
nand U7512 (N_7512,N_6628,N_7077);
or U7513 (N_7513,N_6551,N_7287);
nand U7514 (N_7514,N_7021,N_6891);
nand U7515 (N_7515,N_6426,N_6366);
and U7516 (N_7516,N_6728,N_7419);
nor U7517 (N_7517,N_6315,N_7081);
nor U7518 (N_7518,N_6895,N_7480);
nor U7519 (N_7519,N_6609,N_6312);
nor U7520 (N_7520,N_6877,N_6361);
nand U7521 (N_7521,N_6952,N_7439);
nor U7522 (N_7522,N_6372,N_7085);
nor U7523 (N_7523,N_6457,N_6657);
nor U7524 (N_7524,N_7058,N_6985);
and U7525 (N_7525,N_7324,N_6799);
xnor U7526 (N_7526,N_6896,N_6658);
and U7527 (N_7527,N_7402,N_6554);
nor U7528 (N_7528,N_7028,N_6475);
or U7529 (N_7529,N_7215,N_7445);
and U7530 (N_7530,N_7141,N_7224);
nand U7531 (N_7531,N_7000,N_7129);
or U7532 (N_7532,N_6313,N_6682);
or U7533 (N_7533,N_6672,N_6613);
xor U7534 (N_7534,N_6731,N_6763);
nor U7535 (N_7535,N_7246,N_7049);
xor U7536 (N_7536,N_6723,N_6592);
or U7537 (N_7537,N_6926,N_7321);
or U7538 (N_7538,N_7189,N_6499);
nor U7539 (N_7539,N_6748,N_7309);
or U7540 (N_7540,N_6638,N_6913);
nand U7541 (N_7541,N_7163,N_6863);
nand U7542 (N_7542,N_7297,N_7422);
xnor U7543 (N_7543,N_6860,N_6667);
xor U7544 (N_7544,N_7030,N_6683);
nand U7545 (N_7545,N_6864,N_7383);
xnor U7546 (N_7546,N_7488,N_7139);
xor U7547 (N_7547,N_6829,N_6612);
nand U7548 (N_7548,N_7203,N_6573);
or U7549 (N_7549,N_7024,N_6935);
and U7550 (N_7550,N_6304,N_7225);
and U7551 (N_7551,N_6452,N_6744);
nor U7552 (N_7552,N_6351,N_6840);
xnor U7553 (N_7553,N_6645,N_6423);
and U7554 (N_7554,N_6948,N_6293);
xor U7555 (N_7555,N_6778,N_7126);
xnor U7556 (N_7556,N_7186,N_6635);
and U7557 (N_7557,N_6779,N_7078);
or U7558 (N_7558,N_6933,N_6602);
xor U7559 (N_7559,N_6663,N_6736);
or U7560 (N_7560,N_7122,N_6471);
nand U7561 (N_7561,N_7076,N_6572);
or U7562 (N_7562,N_6804,N_6869);
nand U7563 (N_7563,N_6535,N_6481);
nor U7564 (N_7564,N_7258,N_6812);
or U7565 (N_7565,N_6828,N_6563);
or U7566 (N_7566,N_6844,N_6598);
or U7567 (N_7567,N_6668,N_7157);
nand U7568 (N_7568,N_7451,N_6587);
nor U7569 (N_7569,N_6754,N_6455);
and U7570 (N_7570,N_7387,N_7442);
nand U7571 (N_7571,N_6394,N_7311);
nor U7572 (N_7572,N_6866,N_6795);
xor U7573 (N_7573,N_7219,N_6655);
or U7574 (N_7574,N_6319,N_6307);
and U7575 (N_7575,N_6287,N_6586);
and U7576 (N_7576,N_6620,N_6698);
nand U7577 (N_7577,N_6339,N_7485);
xnor U7578 (N_7578,N_7052,N_6327);
xnor U7579 (N_7579,N_7216,N_6502);
xor U7580 (N_7580,N_6711,N_6943);
and U7581 (N_7581,N_7100,N_6934);
nor U7582 (N_7582,N_7332,N_7271);
or U7583 (N_7583,N_7367,N_6399);
xnor U7584 (N_7584,N_7391,N_6953);
and U7585 (N_7585,N_6797,N_6922);
xor U7586 (N_7586,N_7088,N_7238);
nor U7587 (N_7587,N_6492,N_7009);
nand U7588 (N_7588,N_7120,N_6541);
or U7589 (N_7589,N_6318,N_6413);
nand U7590 (N_7590,N_6837,N_7036);
nor U7591 (N_7591,N_7338,N_6969);
and U7592 (N_7592,N_6940,N_7276);
xnor U7593 (N_7593,N_6478,N_7191);
and U7594 (N_7594,N_6856,N_7353);
nand U7595 (N_7595,N_7371,N_6273);
and U7596 (N_7596,N_7042,N_7341);
and U7597 (N_7597,N_6727,N_6803);
nor U7598 (N_7598,N_6382,N_7093);
xnor U7599 (N_7599,N_7170,N_7034);
nor U7600 (N_7600,N_7427,N_6430);
xnor U7601 (N_7601,N_6912,N_6855);
and U7602 (N_7602,N_6400,N_6718);
nand U7603 (N_7603,N_6278,N_6849);
xnor U7604 (N_7604,N_6782,N_6809);
xnor U7605 (N_7605,N_7428,N_6775);
or U7606 (N_7606,N_7357,N_6352);
nor U7607 (N_7607,N_6890,N_7064);
nor U7608 (N_7608,N_6525,N_6462);
xor U7609 (N_7609,N_6376,N_7339);
nor U7610 (N_7610,N_7183,N_7306);
and U7611 (N_7611,N_6691,N_7408);
and U7612 (N_7612,N_6739,N_7474);
nor U7613 (N_7613,N_6356,N_6871);
xor U7614 (N_7614,N_7273,N_7117);
nand U7615 (N_7615,N_6365,N_7452);
nand U7616 (N_7616,N_7421,N_6927);
nor U7617 (N_7617,N_6557,N_7075);
and U7618 (N_7618,N_7360,N_6373);
xnor U7619 (N_7619,N_6725,N_6652);
xnor U7620 (N_7620,N_6265,N_6666);
nor U7621 (N_7621,N_6360,N_7006);
and U7622 (N_7622,N_6729,N_7498);
and U7623 (N_7623,N_7063,N_7154);
xor U7624 (N_7624,N_7086,N_6870);
nor U7625 (N_7625,N_6343,N_6421);
nor U7626 (N_7626,N_6879,N_7411);
xor U7627 (N_7627,N_7396,N_7368);
and U7628 (N_7628,N_7050,N_6429);
nor U7629 (N_7629,N_6721,N_7403);
and U7630 (N_7630,N_7275,N_6401);
or U7631 (N_7631,N_7337,N_6824);
xnor U7632 (N_7632,N_6531,N_7331);
and U7633 (N_7633,N_6619,N_6646);
nor U7634 (N_7634,N_6751,N_6617);
xnor U7635 (N_7635,N_6636,N_7248);
nand U7636 (N_7636,N_6522,N_7267);
and U7637 (N_7637,N_7202,N_6410);
nand U7638 (N_7638,N_7443,N_6905);
nand U7639 (N_7639,N_7406,N_6689);
xor U7640 (N_7640,N_6815,N_6461);
xnor U7641 (N_7641,N_7264,N_6707);
and U7642 (N_7642,N_6988,N_6280);
or U7643 (N_7643,N_7210,N_6949);
xnor U7644 (N_7644,N_6906,N_7431);
nand U7645 (N_7645,N_6616,N_7027);
nand U7646 (N_7646,N_7207,N_6536);
and U7647 (N_7647,N_7294,N_7486);
xor U7648 (N_7648,N_6850,N_6370);
nand U7649 (N_7649,N_6450,N_7255);
or U7650 (N_7650,N_7146,N_7145);
xor U7651 (N_7651,N_7148,N_7471);
nor U7652 (N_7652,N_6848,N_6348);
xor U7653 (N_7653,N_6875,N_7231);
or U7654 (N_7654,N_7254,N_6738);
xnor U7655 (N_7655,N_7090,N_6303);
xor U7656 (N_7656,N_6390,N_6381);
xor U7657 (N_7657,N_7319,N_6605);
and U7658 (N_7658,N_6545,N_6703);
or U7659 (N_7659,N_6630,N_6791);
nand U7660 (N_7660,N_6363,N_6574);
or U7661 (N_7661,N_6811,N_6254);
and U7662 (N_7662,N_7001,N_6769);
or U7663 (N_7663,N_6677,N_6454);
xnor U7664 (N_7664,N_7212,N_6561);
xor U7665 (N_7665,N_7138,N_6966);
or U7666 (N_7666,N_6653,N_6567);
or U7667 (N_7667,N_7010,N_7347);
or U7668 (N_7668,N_6409,N_6514);
xor U7669 (N_7669,N_6286,N_6301);
and U7670 (N_7670,N_6353,N_6438);
xor U7671 (N_7671,N_6651,N_6833);
nor U7672 (N_7672,N_6579,N_6575);
and U7673 (N_7673,N_6957,N_7134);
xnor U7674 (N_7674,N_6669,N_6555);
and U7675 (N_7675,N_6649,N_6272);
or U7676 (N_7676,N_6865,N_6368);
or U7677 (N_7677,N_6539,N_6469);
xnor U7678 (N_7678,N_6416,N_6379);
xnor U7679 (N_7679,N_7320,N_6914);
xnor U7680 (N_7680,N_6606,N_6904);
and U7681 (N_7681,N_6862,N_6627);
or U7682 (N_7682,N_6810,N_6964);
or U7683 (N_7683,N_7462,N_6767);
or U7684 (N_7684,N_6302,N_6533);
nand U7685 (N_7685,N_6960,N_6827);
and U7686 (N_7686,N_6456,N_6634);
xor U7687 (N_7687,N_6623,N_7286);
and U7688 (N_7688,N_7364,N_7362);
nand U7689 (N_7689,N_7178,N_6476);
and U7690 (N_7690,N_7187,N_7323);
nand U7691 (N_7691,N_7489,N_7062);
nor U7692 (N_7692,N_7269,N_7053);
xor U7693 (N_7693,N_6578,N_6509);
xnor U7694 (N_7694,N_7281,N_6760);
or U7695 (N_7695,N_7430,N_7179);
and U7696 (N_7696,N_6780,N_7327);
nand U7697 (N_7697,N_6724,N_7025);
nand U7698 (N_7698,N_7315,N_7113);
nand U7699 (N_7699,N_6479,N_7102);
or U7700 (N_7700,N_6377,N_7334);
nand U7701 (N_7701,N_7200,N_7404);
and U7702 (N_7702,N_6640,N_6747);
nand U7703 (N_7703,N_6437,N_7328);
or U7704 (N_7704,N_6992,N_7017);
xnor U7705 (N_7705,N_6337,N_6886);
or U7706 (N_7706,N_7348,N_7222);
or U7707 (N_7707,N_6694,N_7366);
or U7708 (N_7708,N_6917,N_7164);
or U7709 (N_7709,N_7124,N_7336);
or U7710 (N_7710,N_7115,N_7140);
nand U7711 (N_7711,N_7342,N_6424);
and U7712 (N_7712,N_7097,N_6942);
nor U7713 (N_7713,N_6432,N_6486);
and U7714 (N_7714,N_6730,N_7051);
nand U7715 (N_7715,N_6283,N_6719);
nand U7716 (N_7716,N_6820,N_7478);
xnor U7717 (N_7717,N_6564,N_6622);
and U7718 (N_7718,N_7071,N_6295);
nand U7719 (N_7719,N_7293,N_6817);
and U7720 (N_7720,N_6521,N_7350);
or U7721 (N_7721,N_6624,N_7172);
or U7722 (N_7722,N_6392,N_7214);
and U7723 (N_7723,N_6793,N_6508);
nor U7724 (N_7724,N_6517,N_6961);
nor U7725 (N_7725,N_6333,N_6965);
and U7726 (N_7726,N_6451,N_6633);
nor U7727 (N_7727,N_7132,N_7162);
and U7728 (N_7728,N_6322,N_7167);
or U7729 (N_7729,N_6512,N_7165);
nand U7730 (N_7730,N_7476,N_7344);
xnor U7731 (N_7731,N_6534,N_7035);
nor U7732 (N_7732,N_7110,N_6671);
xnor U7733 (N_7733,N_6790,N_6527);
nor U7734 (N_7734,N_6997,N_6532);
xor U7735 (N_7735,N_6680,N_6956);
xor U7736 (N_7736,N_6746,N_6264);
xor U7737 (N_7737,N_6709,N_6299);
nand U7738 (N_7738,N_6321,N_6749);
or U7739 (N_7739,N_6702,N_7377);
nor U7740 (N_7740,N_7182,N_6524);
xnor U7741 (N_7741,N_6501,N_7026);
nand U7742 (N_7742,N_6305,N_6310);
or U7743 (N_7743,N_6753,N_6773);
or U7744 (N_7744,N_6899,N_7180);
and U7745 (N_7745,N_6897,N_6297);
or U7746 (N_7746,N_6459,N_7103);
nor U7747 (N_7747,N_6553,N_6362);
or U7748 (N_7748,N_6786,N_7069);
xor U7749 (N_7749,N_7380,N_6994);
or U7750 (N_7750,N_6334,N_6783);
nor U7751 (N_7751,N_7376,N_6446);
nand U7752 (N_7752,N_7308,N_7418);
nand U7753 (N_7753,N_6675,N_7232);
nor U7754 (N_7754,N_6407,N_6496);
nand U7755 (N_7755,N_6581,N_7363);
xor U7756 (N_7756,N_6838,N_6277);
or U7757 (N_7757,N_7416,N_6656);
nor U7758 (N_7758,N_6474,N_6951);
nand U7759 (N_7759,N_6428,N_6484);
nand U7760 (N_7760,N_6258,N_6632);
or U7761 (N_7761,N_6962,N_6583);
nor U7762 (N_7762,N_6503,N_6546);
nand U7763 (N_7763,N_7382,N_7358);
xor U7764 (N_7764,N_7241,N_7450);
xor U7765 (N_7765,N_6742,N_7011);
nor U7766 (N_7766,N_7277,N_7066);
nand U7767 (N_7767,N_7242,N_6745);
nand U7768 (N_7768,N_6910,N_6989);
nand U7769 (N_7769,N_7251,N_7155);
xor U7770 (N_7770,N_6349,N_6944);
xnor U7771 (N_7771,N_7268,N_6859);
and U7772 (N_7772,N_7453,N_7108);
nand U7773 (N_7773,N_6806,N_7262);
nor U7774 (N_7774,N_6530,N_6673);
or U7775 (N_7775,N_6420,N_6275);
or U7776 (N_7776,N_7057,N_6684);
nand U7777 (N_7777,N_6991,N_6594);
nor U7778 (N_7778,N_6449,N_6591);
nor U7779 (N_7779,N_6388,N_6821);
xor U7780 (N_7780,N_6878,N_6713);
nand U7781 (N_7781,N_6872,N_6516);
and U7782 (N_7782,N_6374,N_6393);
and U7783 (N_7783,N_6894,N_6902);
nor U7784 (N_7784,N_7313,N_6662);
nor U7785 (N_7785,N_7409,N_6996);
and U7786 (N_7786,N_7265,N_6528);
or U7787 (N_7787,N_6285,N_7061);
and U7788 (N_7788,N_7410,N_6369);
xnor U7789 (N_7789,N_7067,N_7394);
or U7790 (N_7790,N_7177,N_6971);
xnor U7791 (N_7791,N_7378,N_7407);
and U7792 (N_7792,N_6759,N_6857);
or U7793 (N_7793,N_7370,N_6851);
or U7794 (N_7794,N_7413,N_6785);
nand U7795 (N_7795,N_7239,N_7259);
nor U7796 (N_7796,N_7169,N_7470);
nand U7797 (N_7797,N_6411,N_6344);
xor U7798 (N_7798,N_6290,N_6441);
nand U7799 (N_7799,N_6483,N_6435);
and U7800 (N_7800,N_7247,N_7429);
or U7801 (N_7801,N_6898,N_6537);
nand U7802 (N_7802,N_6916,N_7361);
or U7803 (N_7803,N_7160,N_6291);
nor U7804 (N_7804,N_6358,N_6761);
or U7805 (N_7805,N_6805,N_6289);
or U7806 (N_7806,N_6936,N_7283);
nor U7807 (N_7807,N_7257,N_6678);
xnor U7808 (N_7808,N_6911,N_6954);
xor U7809 (N_7809,N_6968,N_7272);
or U7810 (N_7810,N_7487,N_6548);
and U7811 (N_7811,N_7374,N_6800);
xnor U7812 (N_7812,N_6571,N_6955);
xnor U7813 (N_7813,N_6984,N_6589);
nor U7814 (N_7814,N_6830,N_7468);
xor U7815 (N_7815,N_6284,N_6704);
xor U7816 (N_7816,N_6519,N_6389);
or U7817 (N_7817,N_6601,N_7424);
and U7818 (N_7818,N_6733,N_6562);
xor U7819 (N_7819,N_6696,N_7135);
nor U7820 (N_7820,N_6422,N_7496);
nor U7821 (N_7821,N_7068,N_7389);
xnor U7822 (N_7822,N_6919,N_6371);
nand U7823 (N_7823,N_7423,N_7318);
and U7824 (N_7824,N_7465,N_6737);
nand U7825 (N_7825,N_7171,N_6405);
nor U7826 (N_7826,N_7420,N_6776);
xor U7827 (N_7827,N_7074,N_6439);
xnor U7828 (N_7828,N_6357,N_6999);
nand U7829 (N_7829,N_6323,N_7070);
and U7830 (N_7830,N_7434,N_6543);
and U7831 (N_7831,N_7226,N_6329);
or U7832 (N_7832,N_6447,N_7379);
nand U7833 (N_7833,N_7083,N_6281);
nor U7834 (N_7834,N_6907,N_7044);
and U7835 (N_7835,N_7401,N_7352);
or U7836 (N_7836,N_6772,N_6887);
xor U7837 (N_7837,N_6367,N_6983);
xor U7838 (N_7838,N_7256,N_6507);
xor U7839 (N_7839,N_7400,N_6568);
xor U7840 (N_7840,N_7296,N_6274);
xor U7841 (N_7841,N_7305,N_7099);
xnor U7842 (N_7842,N_7073,N_6585);
or U7843 (N_7843,N_6963,N_6764);
xor U7844 (N_7844,N_6706,N_6929);
nand U7845 (N_7845,N_6482,N_6314);
nor U7846 (N_7846,N_6903,N_7091);
and U7847 (N_7847,N_7022,N_6686);
and U7848 (N_7848,N_6726,N_7312);
xnor U7849 (N_7849,N_7038,N_7121);
nor U7850 (N_7850,N_7436,N_6705);
xor U7851 (N_7851,N_7274,N_6882);
xor U7852 (N_7852,N_7373,N_6336);
or U7853 (N_7853,N_7045,N_6607);
and U7854 (N_7854,N_7019,N_6477);
or U7855 (N_7855,N_7475,N_6588);
nor U7856 (N_7856,N_6330,N_7125);
or U7857 (N_7857,N_6813,N_7221);
or U7858 (N_7858,N_6676,N_7249);
nor U7859 (N_7859,N_6270,N_7185);
xor U7860 (N_7860,N_6661,N_6271);
nand U7861 (N_7861,N_6980,N_6440);
xor U7862 (N_7862,N_7016,N_6506);
nor U7863 (N_7863,N_6354,N_7301);
xor U7864 (N_7864,N_7481,N_6970);
and U7865 (N_7865,N_6937,N_7447);
xnor U7866 (N_7866,N_6404,N_7142);
xnor U7867 (N_7867,N_6720,N_7218);
and U7868 (N_7868,N_6644,N_6801);
nand U7869 (N_7869,N_6993,N_7356);
or U7870 (N_7870,N_6267,N_6885);
xor U7871 (N_7871,N_7194,N_6834);
nand U7872 (N_7872,N_7493,N_6695);
and U7873 (N_7873,N_6752,N_7329);
nand U7874 (N_7874,N_7184,N_6266);
nor U7875 (N_7875,N_7456,N_7477);
nand U7876 (N_7876,N_6542,N_7414);
nor U7877 (N_7877,N_6335,N_6853);
or U7878 (N_7878,N_6768,N_6338);
xor U7879 (N_7879,N_7087,N_6639);
nor U7880 (N_7880,N_7227,N_7317);
or U7881 (N_7881,N_6331,N_6294);
or U7882 (N_7882,N_6978,N_6690);
nand U7883 (N_7883,N_6986,N_6659);
nor U7884 (N_7884,N_7046,N_7039);
nor U7885 (N_7885,N_6883,N_6974);
and U7886 (N_7886,N_7107,N_7033);
and U7887 (N_7887,N_6755,N_7278);
nor U7888 (N_7888,N_7054,N_7188);
xnor U7889 (N_7889,N_6489,N_7333);
and U7890 (N_7890,N_6414,N_7386);
nor U7891 (N_7891,N_6433,N_6664);
nor U7892 (N_7892,N_7193,N_7290);
nand U7893 (N_7893,N_6732,N_7197);
nand U7894 (N_7894,N_6681,N_6253);
xor U7895 (N_7895,N_7351,N_6831);
nor U7896 (N_7896,N_7398,N_7284);
nor U7897 (N_7897,N_6892,N_6480);
or U7898 (N_7898,N_7005,N_6495);
and U7899 (N_7899,N_7340,N_6444);
nor U7900 (N_7900,N_7065,N_7244);
xnor U7901 (N_7901,N_6740,N_6346);
xor U7902 (N_7902,N_6397,N_6685);
nand U7903 (N_7903,N_6466,N_7455);
nor U7904 (N_7904,N_6631,N_6771);
xor U7905 (N_7905,N_6538,N_6873);
nand U7906 (N_7906,N_7243,N_6549);
and U7907 (N_7907,N_7079,N_6491);
nand U7908 (N_7908,N_6975,N_7459);
or U7909 (N_7909,N_6463,N_6311);
nand U7910 (N_7910,N_6816,N_6615);
nor U7911 (N_7911,N_7472,N_6893);
nor U7912 (N_7912,N_7289,N_7003);
nand U7913 (N_7913,N_7282,N_7446);
or U7914 (N_7914,N_6500,N_6712);
or U7915 (N_7915,N_6257,N_6977);
or U7916 (N_7916,N_7192,N_6987);
and U7917 (N_7917,N_7143,N_7384);
nor U7918 (N_7918,N_6939,N_6692);
xor U7919 (N_7919,N_6596,N_7041);
or U7920 (N_7920,N_7303,N_7131);
or U7921 (N_7921,N_6570,N_7448);
nor U7922 (N_7922,N_7048,N_7111);
xnor U7923 (N_7923,N_6597,N_7291);
nand U7924 (N_7924,N_6443,N_7147);
xnor U7925 (N_7925,N_6908,N_6547);
nand U7926 (N_7926,N_7279,N_6436);
nor U7927 (N_7927,N_6510,N_6839);
nor U7928 (N_7928,N_7144,N_6340);
nor U7929 (N_7929,N_7372,N_6577);
xnor U7930 (N_7930,N_6359,N_7345);
or U7931 (N_7931,N_6317,N_6867);
nor U7932 (N_7932,N_7314,N_7151);
and U7933 (N_7933,N_6262,N_6654);
nor U7934 (N_7934,N_7096,N_7397);
and U7935 (N_7935,N_6590,N_7130);
and U7936 (N_7936,N_7014,N_6298);
and U7937 (N_7937,N_6544,N_6556);
and U7938 (N_7938,N_6881,N_6998);
nand U7939 (N_7939,N_6693,N_6900);
and U7940 (N_7940,N_6453,N_6292);
or U7941 (N_7941,N_6757,N_6378);
xor U7942 (N_7942,N_7173,N_6497);
xnor U7943 (N_7943,N_6473,N_6427);
nand U7944 (N_7944,N_7159,N_6259);
nor U7945 (N_7945,N_6279,N_6626);
and U7946 (N_7946,N_6464,N_6741);
or U7947 (N_7947,N_7458,N_7235);
and U7948 (N_7948,N_7490,N_6715);
xor U7949 (N_7949,N_7161,N_7007);
xnor U7950 (N_7950,N_7206,N_6814);
nor U7951 (N_7951,N_6398,N_6558);
or U7952 (N_7952,N_6920,N_6750);
nor U7953 (N_7953,N_7149,N_6967);
xor U7954 (N_7954,N_6802,N_7176);
xnor U7955 (N_7955,N_7181,N_6593);
and U7956 (N_7956,N_6408,N_6822);
nand U7957 (N_7957,N_7236,N_6402);
and U7958 (N_7958,N_6498,N_6316);
or U7959 (N_7959,N_7432,N_6637);
and U7960 (N_7960,N_6688,N_6674);
xnor U7961 (N_7961,N_7261,N_6854);
xor U7962 (N_7962,N_6520,N_6918);
nor U7963 (N_7963,N_7127,N_7116);
nand U7964 (N_7964,N_6874,N_7150);
or U7965 (N_7965,N_6487,N_7029);
xnor U7966 (N_7966,N_7388,N_7467);
or U7967 (N_7967,N_6982,N_6901);
or U7968 (N_7968,N_6858,N_7004);
nand U7969 (N_7969,N_6364,N_6580);
or U7970 (N_7970,N_7156,N_6511);
or U7971 (N_7971,N_6396,N_6326);
nand U7972 (N_7972,N_7092,N_6701);
nor U7973 (N_7973,N_7211,N_7417);
nor U7974 (N_7974,N_6700,N_7084);
nand U7975 (N_7975,N_7466,N_7449);
nor U7976 (N_7976,N_7094,N_6250);
nand U7977 (N_7977,N_6251,N_7304);
and U7978 (N_7978,N_7365,N_6756);
nand U7979 (N_7979,N_6979,N_7326);
nand U7980 (N_7980,N_6576,N_7385);
nand U7981 (N_7981,N_7454,N_6261);
xor U7982 (N_7982,N_7473,N_6976);
nand U7983 (N_7983,N_7056,N_6641);
nand U7984 (N_7984,N_7174,N_7395);
nor U7985 (N_7985,N_6419,N_6847);
nand U7986 (N_7986,N_7152,N_7233);
nor U7987 (N_7987,N_6990,N_6766);
nand U7988 (N_7988,N_7492,N_7295);
and U7989 (N_7989,N_6415,N_6610);
or U7990 (N_7990,N_6921,N_7082);
or U7991 (N_7991,N_6458,N_6505);
xor U7992 (N_7992,N_6826,N_6513);
nor U7993 (N_7993,N_7441,N_7204);
xor U7994 (N_7994,N_6472,N_7457);
xor U7995 (N_7995,N_6406,N_7325);
xor U7996 (N_7996,N_6526,N_6841);
nand U7997 (N_7997,N_6876,N_6599);
nor U7998 (N_7998,N_7205,N_6328);
and U7999 (N_7999,N_6660,N_6582);
or U8000 (N_8000,N_7482,N_6350);
nand U8001 (N_8001,N_6924,N_6621);
xor U8002 (N_8002,N_6595,N_6618);
xor U8003 (N_8003,N_6467,N_7435);
or U8004 (N_8004,N_7158,N_6395);
xnor U8005 (N_8005,N_7104,N_6306);
and U8006 (N_8006,N_6932,N_6665);
xnor U8007 (N_8007,N_6784,N_6494);
xor U8008 (N_8008,N_6403,N_6925);
or U8009 (N_8009,N_7060,N_7415);
xnor U8010 (N_8010,N_6470,N_6787);
nor U8011 (N_8011,N_7015,N_6614);
xnor U8012 (N_8012,N_6947,N_6386);
or U8013 (N_8013,N_6647,N_6515);
and U8014 (N_8014,N_7250,N_6565);
xor U8015 (N_8015,N_7072,N_6468);
or U8016 (N_8016,N_7032,N_6603);
nor U8017 (N_8017,N_7230,N_6774);
xor U8018 (N_8018,N_7491,N_6252);
xnor U8019 (N_8019,N_7240,N_7425);
xor U8020 (N_8020,N_7285,N_6923);
or U8021 (N_8021,N_6861,N_7002);
nand U8022 (N_8022,N_7037,N_6832);
or U8023 (N_8023,N_6324,N_7499);
xor U8024 (N_8024,N_6670,N_7310);
xnor U8025 (N_8025,N_6758,N_6269);
xnor U8026 (N_8026,N_6256,N_7288);
and U8027 (N_8027,N_7426,N_6309);
and U8028 (N_8028,N_7012,N_7043);
nor U8029 (N_8029,N_7234,N_7260);
nor U8030 (N_8030,N_7008,N_6611);
xor U8031 (N_8031,N_6889,N_6341);
nand U8032 (N_8032,N_6448,N_7031);
xor U8033 (N_8033,N_7263,N_7245);
xor U8034 (N_8034,N_6345,N_6716);
or U8035 (N_8035,N_7128,N_7330);
or U8036 (N_8036,N_6375,N_6485);
nor U8037 (N_8037,N_7137,N_6325);
nor U8038 (N_8038,N_6735,N_6425);
or U8039 (N_8039,N_6465,N_6762);
nand U8040 (N_8040,N_6648,N_6836);
nand U8041 (N_8041,N_6888,N_6958);
nor U8042 (N_8042,N_6807,N_6842);
nor U8043 (N_8043,N_7223,N_7055);
nand U8044 (N_8044,N_7101,N_6880);
xor U8045 (N_8045,N_6523,N_7381);
and U8046 (N_8046,N_7175,N_7299);
xnor U8047 (N_8047,N_6981,N_7059);
xor U8048 (N_8048,N_7040,N_7484);
and U8049 (N_8049,N_6296,N_7266);
xor U8050 (N_8050,N_6825,N_7106);
and U8051 (N_8051,N_7463,N_6387);
and U8052 (N_8052,N_6734,N_7018);
and U8053 (N_8053,N_6938,N_6460);
nand U8054 (N_8054,N_7461,N_7109);
xnor U8055 (N_8055,N_6868,N_6604);
and U8056 (N_8056,N_7440,N_6391);
xnor U8057 (N_8057,N_6308,N_7114);
nor U8058 (N_8058,N_6288,N_7433);
xnor U8059 (N_8059,N_6625,N_7322);
and U8060 (N_8060,N_6835,N_6434);
and U8061 (N_8061,N_6417,N_6412);
or U8062 (N_8062,N_7375,N_6798);
xnor U8063 (N_8063,N_6931,N_7209);
xnor U8064 (N_8064,N_7464,N_7198);
nor U8065 (N_8065,N_6781,N_7497);
and U8066 (N_8066,N_6819,N_7201);
or U8067 (N_8067,N_6300,N_6488);
xor U8068 (N_8068,N_6722,N_7118);
nand U8069 (N_8069,N_7343,N_7013);
nor U8070 (N_8070,N_6789,N_6743);
nor U8071 (N_8071,N_7119,N_7199);
or U8072 (N_8072,N_7080,N_7190);
or U8073 (N_8073,N_6629,N_6550);
or U8074 (N_8074,N_6490,N_7483);
and U8075 (N_8075,N_7228,N_6282);
or U8076 (N_8076,N_6915,N_7098);
and U8077 (N_8077,N_6959,N_7229);
nand U8078 (N_8078,N_6946,N_6717);
nor U8079 (N_8079,N_6796,N_6928);
and U8080 (N_8080,N_6699,N_7346);
or U8081 (N_8081,N_7494,N_6710);
or U8082 (N_8082,N_6600,N_6263);
and U8083 (N_8083,N_7405,N_6504);
or U8084 (N_8084,N_6445,N_6518);
or U8085 (N_8085,N_6418,N_7369);
nor U8086 (N_8086,N_7237,N_6945);
or U8087 (N_8087,N_6852,N_6788);
xor U8088 (N_8088,N_6384,N_6355);
xnor U8089 (N_8089,N_7355,N_6540);
nor U8090 (N_8090,N_6431,N_6909);
nor U8091 (N_8091,N_6714,N_6679);
xor U8092 (N_8092,N_7302,N_7123);
or U8093 (N_8093,N_6529,N_7166);
nor U8094 (N_8094,N_6566,N_6777);
or U8095 (N_8095,N_7217,N_6697);
xnor U8096 (N_8096,N_7359,N_6380);
nand U8097 (N_8097,N_6765,N_6941);
nand U8098 (N_8098,N_6823,N_6569);
or U8099 (N_8099,N_6708,N_6818);
xor U8100 (N_8100,N_7437,N_7495);
or U8101 (N_8101,N_6385,N_6643);
or U8102 (N_8102,N_7412,N_7300);
or U8103 (N_8103,N_6930,N_6792);
xor U8104 (N_8104,N_6950,N_6255);
or U8105 (N_8105,N_6608,N_7168);
and U8106 (N_8106,N_7298,N_7089);
nand U8107 (N_8107,N_7195,N_7469);
and U8108 (N_8108,N_7399,N_7479);
nor U8109 (N_8109,N_7136,N_6268);
xnor U8110 (N_8110,N_6794,N_7280);
nand U8111 (N_8111,N_7023,N_7105);
xnor U8112 (N_8112,N_7307,N_6260);
xor U8113 (N_8113,N_7153,N_7253);
or U8114 (N_8114,N_6846,N_7252);
nor U8115 (N_8115,N_7020,N_7095);
xor U8116 (N_8116,N_7270,N_7438);
or U8117 (N_8117,N_6560,N_7292);
and U8118 (N_8118,N_6770,N_6843);
and U8119 (N_8119,N_6584,N_7393);
and U8120 (N_8120,N_6332,N_6972);
xnor U8121 (N_8121,N_7390,N_6442);
nand U8122 (N_8122,N_7460,N_7354);
nor U8123 (N_8123,N_7213,N_7220);
nand U8124 (N_8124,N_6884,N_6642);
xnor U8125 (N_8125,N_6717,N_7169);
nand U8126 (N_8126,N_6526,N_7209);
or U8127 (N_8127,N_6532,N_7016);
nand U8128 (N_8128,N_6806,N_6610);
xor U8129 (N_8129,N_6969,N_6802);
nor U8130 (N_8130,N_6393,N_6816);
and U8131 (N_8131,N_7135,N_7110);
xnor U8132 (N_8132,N_6593,N_7362);
nand U8133 (N_8133,N_6498,N_7313);
or U8134 (N_8134,N_6632,N_6420);
nand U8135 (N_8135,N_6940,N_6301);
or U8136 (N_8136,N_6403,N_7291);
or U8137 (N_8137,N_6908,N_7014);
xnor U8138 (N_8138,N_6818,N_7492);
xor U8139 (N_8139,N_6580,N_7464);
nor U8140 (N_8140,N_7035,N_6853);
or U8141 (N_8141,N_7093,N_6725);
and U8142 (N_8142,N_6874,N_6572);
and U8143 (N_8143,N_6602,N_6309);
or U8144 (N_8144,N_6386,N_6469);
xnor U8145 (N_8145,N_7092,N_6681);
nand U8146 (N_8146,N_7258,N_7052);
nand U8147 (N_8147,N_6836,N_6280);
or U8148 (N_8148,N_7393,N_6891);
or U8149 (N_8149,N_7103,N_6891);
and U8150 (N_8150,N_6721,N_7486);
nand U8151 (N_8151,N_6267,N_7320);
or U8152 (N_8152,N_6774,N_7309);
or U8153 (N_8153,N_6966,N_6453);
or U8154 (N_8154,N_7017,N_6851);
nand U8155 (N_8155,N_6961,N_6767);
and U8156 (N_8156,N_7141,N_7498);
xnor U8157 (N_8157,N_6285,N_7107);
or U8158 (N_8158,N_7201,N_6733);
xor U8159 (N_8159,N_6288,N_6375);
xnor U8160 (N_8160,N_7455,N_7072);
or U8161 (N_8161,N_6336,N_6433);
and U8162 (N_8162,N_7306,N_7128);
nand U8163 (N_8163,N_7468,N_7445);
and U8164 (N_8164,N_6695,N_6436);
nand U8165 (N_8165,N_6903,N_6555);
or U8166 (N_8166,N_6703,N_7226);
nor U8167 (N_8167,N_7062,N_6695);
nor U8168 (N_8168,N_7380,N_6375);
nand U8169 (N_8169,N_7437,N_7303);
nor U8170 (N_8170,N_6710,N_6540);
nor U8171 (N_8171,N_7395,N_6737);
xnor U8172 (N_8172,N_6375,N_6312);
and U8173 (N_8173,N_6849,N_6881);
nor U8174 (N_8174,N_6614,N_7268);
and U8175 (N_8175,N_6958,N_6342);
or U8176 (N_8176,N_6906,N_6302);
or U8177 (N_8177,N_6874,N_6878);
nor U8178 (N_8178,N_6846,N_6451);
nand U8179 (N_8179,N_7240,N_6843);
nand U8180 (N_8180,N_7177,N_7130);
xnor U8181 (N_8181,N_6339,N_6549);
and U8182 (N_8182,N_6924,N_6557);
nand U8183 (N_8183,N_7096,N_6398);
xnor U8184 (N_8184,N_7463,N_6533);
or U8185 (N_8185,N_6963,N_7075);
xor U8186 (N_8186,N_6389,N_7029);
nand U8187 (N_8187,N_7097,N_7052);
xnor U8188 (N_8188,N_7323,N_6796);
and U8189 (N_8189,N_6257,N_6297);
nand U8190 (N_8190,N_6762,N_7213);
xnor U8191 (N_8191,N_6870,N_7092);
or U8192 (N_8192,N_6365,N_7239);
or U8193 (N_8193,N_6692,N_6818);
xor U8194 (N_8194,N_7209,N_6457);
xnor U8195 (N_8195,N_7305,N_6792);
nand U8196 (N_8196,N_7461,N_6324);
nand U8197 (N_8197,N_7271,N_6928);
or U8198 (N_8198,N_6869,N_6755);
xnor U8199 (N_8199,N_6562,N_6648);
nor U8200 (N_8200,N_6737,N_6687);
nor U8201 (N_8201,N_7341,N_7093);
and U8202 (N_8202,N_7051,N_6449);
nand U8203 (N_8203,N_7469,N_7319);
and U8204 (N_8204,N_6897,N_7337);
nand U8205 (N_8205,N_7186,N_7258);
or U8206 (N_8206,N_7304,N_6858);
or U8207 (N_8207,N_7334,N_6492);
or U8208 (N_8208,N_6939,N_7038);
xnor U8209 (N_8209,N_7228,N_6483);
xnor U8210 (N_8210,N_7003,N_6818);
nor U8211 (N_8211,N_6401,N_6873);
nor U8212 (N_8212,N_7280,N_6522);
and U8213 (N_8213,N_6980,N_6803);
or U8214 (N_8214,N_6545,N_7244);
xor U8215 (N_8215,N_7490,N_6331);
nor U8216 (N_8216,N_6824,N_6447);
xor U8217 (N_8217,N_6497,N_6287);
nor U8218 (N_8218,N_6719,N_7052);
and U8219 (N_8219,N_6338,N_6499);
and U8220 (N_8220,N_6594,N_6416);
xor U8221 (N_8221,N_7282,N_7209);
and U8222 (N_8222,N_7413,N_7255);
nor U8223 (N_8223,N_7153,N_6263);
nand U8224 (N_8224,N_6888,N_6541);
or U8225 (N_8225,N_7048,N_6503);
xnor U8226 (N_8226,N_6844,N_6420);
nand U8227 (N_8227,N_7387,N_6642);
nand U8228 (N_8228,N_7228,N_7450);
or U8229 (N_8229,N_7009,N_7325);
or U8230 (N_8230,N_6679,N_6413);
nor U8231 (N_8231,N_7259,N_7167);
and U8232 (N_8232,N_7311,N_7000);
or U8233 (N_8233,N_7213,N_7297);
xor U8234 (N_8234,N_6881,N_6879);
nor U8235 (N_8235,N_6685,N_6852);
nor U8236 (N_8236,N_6402,N_6938);
xor U8237 (N_8237,N_6909,N_6974);
nor U8238 (N_8238,N_7150,N_7062);
nor U8239 (N_8239,N_7056,N_6868);
nor U8240 (N_8240,N_6337,N_6864);
nor U8241 (N_8241,N_7143,N_6917);
and U8242 (N_8242,N_6644,N_7499);
nor U8243 (N_8243,N_6903,N_7089);
nand U8244 (N_8244,N_7144,N_7342);
xor U8245 (N_8245,N_6830,N_6484);
and U8246 (N_8246,N_7489,N_6754);
nand U8247 (N_8247,N_6909,N_6495);
nand U8248 (N_8248,N_7006,N_6254);
nor U8249 (N_8249,N_6303,N_7352);
nand U8250 (N_8250,N_7014,N_6473);
or U8251 (N_8251,N_6479,N_6586);
nor U8252 (N_8252,N_7284,N_6549);
nor U8253 (N_8253,N_7360,N_6981);
xor U8254 (N_8254,N_7443,N_6288);
or U8255 (N_8255,N_6294,N_6763);
xor U8256 (N_8256,N_6592,N_6605);
and U8257 (N_8257,N_6256,N_6696);
and U8258 (N_8258,N_7166,N_6799);
and U8259 (N_8259,N_7010,N_6804);
nor U8260 (N_8260,N_7274,N_7096);
and U8261 (N_8261,N_6933,N_7201);
nor U8262 (N_8262,N_6272,N_6929);
or U8263 (N_8263,N_7076,N_6362);
xnor U8264 (N_8264,N_7295,N_6630);
and U8265 (N_8265,N_6917,N_6518);
xor U8266 (N_8266,N_6520,N_6412);
nor U8267 (N_8267,N_7497,N_6858);
xor U8268 (N_8268,N_6906,N_7126);
nor U8269 (N_8269,N_6951,N_6682);
xor U8270 (N_8270,N_7192,N_6660);
xor U8271 (N_8271,N_7264,N_7206);
and U8272 (N_8272,N_7171,N_7036);
or U8273 (N_8273,N_6746,N_7309);
nand U8274 (N_8274,N_7398,N_6254);
and U8275 (N_8275,N_6919,N_6543);
and U8276 (N_8276,N_7229,N_6410);
nor U8277 (N_8277,N_6569,N_6783);
nand U8278 (N_8278,N_6478,N_6947);
or U8279 (N_8279,N_7386,N_7173);
nor U8280 (N_8280,N_6792,N_7436);
nand U8281 (N_8281,N_6614,N_7338);
nand U8282 (N_8282,N_6688,N_7002);
nor U8283 (N_8283,N_7111,N_6647);
xnor U8284 (N_8284,N_6688,N_6397);
and U8285 (N_8285,N_7031,N_7200);
and U8286 (N_8286,N_6583,N_6543);
and U8287 (N_8287,N_6429,N_6582);
nor U8288 (N_8288,N_6327,N_7276);
xnor U8289 (N_8289,N_6544,N_6745);
nor U8290 (N_8290,N_6415,N_6378);
nand U8291 (N_8291,N_6401,N_6864);
nor U8292 (N_8292,N_6455,N_7205);
nand U8293 (N_8293,N_6394,N_6404);
or U8294 (N_8294,N_7247,N_7356);
and U8295 (N_8295,N_7214,N_7358);
and U8296 (N_8296,N_6821,N_6363);
nor U8297 (N_8297,N_6735,N_6750);
or U8298 (N_8298,N_7314,N_6710);
or U8299 (N_8299,N_7246,N_6883);
or U8300 (N_8300,N_6451,N_7480);
nor U8301 (N_8301,N_6942,N_6606);
nand U8302 (N_8302,N_7205,N_6883);
nor U8303 (N_8303,N_6726,N_6940);
nand U8304 (N_8304,N_6570,N_6722);
nand U8305 (N_8305,N_7372,N_7324);
or U8306 (N_8306,N_6793,N_6276);
nand U8307 (N_8307,N_6521,N_7210);
or U8308 (N_8308,N_6392,N_6280);
xor U8309 (N_8309,N_6534,N_7072);
nand U8310 (N_8310,N_6428,N_7336);
and U8311 (N_8311,N_7038,N_6961);
nor U8312 (N_8312,N_7277,N_6301);
xnor U8313 (N_8313,N_7476,N_7104);
nor U8314 (N_8314,N_6476,N_6358);
xnor U8315 (N_8315,N_6717,N_6954);
nand U8316 (N_8316,N_6748,N_7295);
nand U8317 (N_8317,N_7237,N_7476);
and U8318 (N_8318,N_7414,N_7321);
nand U8319 (N_8319,N_7377,N_7316);
or U8320 (N_8320,N_6641,N_6626);
nand U8321 (N_8321,N_7179,N_7201);
or U8322 (N_8322,N_7366,N_6536);
or U8323 (N_8323,N_7176,N_6498);
xor U8324 (N_8324,N_6787,N_6733);
nand U8325 (N_8325,N_6686,N_7183);
nand U8326 (N_8326,N_7068,N_7288);
nor U8327 (N_8327,N_6340,N_7207);
or U8328 (N_8328,N_6772,N_6736);
xnor U8329 (N_8329,N_7467,N_6855);
nor U8330 (N_8330,N_6526,N_6886);
or U8331 (N_8331,N_6603,N_6526);
nand U8332 (N_8332,N_6616,N_6417);
nor U8333 (N_8333,N_7285,N_6508);
nand U8334 (N_8334,N_6783,N_7308);
xnor U8335 (N_8335,N_7177,N_7481);
nand U8336 (N_8336,N_7491,N_7212);
nand U8337 (N_8337,N_6850,N_7109);
or U8338 (N_8338,N_6496,N_7046);
nor U8339 (N_8339,N_7464,N_6933);
nand U8340 (N_8340,N_6363,N_6637);
xnor U8341 (N_8341,N_6447,N_7285);
xnor U8342 (N_8342,N_6479,N_6829);
xnor U8343 (N_8343,N_7469,N_6944);
nand U8344 (N_8344,N_7179,N_6958);
nor U8345 (N_8345,N_6813,N_7432);
nand U8346 (N_8346,N_6692,N_7391);
nor U8347 (N_8347,N_6786,N_6832);
nand U8348 (N_8348,N_6491,N_6729);
nand U8349 (N_8349,N_6860,N_7282);
and U8350 (N_8350,N_6486,N_7347);
nand U8351 (N_8351,N_6521,N_6562);
nor U8352 (N_8352,N_6297,N_7382);
or U8353 (N_8353,N_6639,N_6899);
and U8354 (N_8354,N_6537,N_7482);
or U8355 (N_8355,N_6890,N_6405);
xor U8356 (N_8356,N_6346,N_7156);
or U8357 (N_8357,N_7282,N_6261);
or U8358 (N_8358,N_6809,N_7069);
and U8359 (N_8359,N_7126,N_6947);
nor U8360 (N_8360,N_7259,N_6905);
or U8361 (N_8361,N_7199,N_7125);
nor U8362 (N_8362,N_7011,N_6813);
nor U8363 (N_8363,N_6829,N_6801);
xnor U8364 (N_8364,N_6370,N_6257);
xor U8365 (N_8365,N_6822,N_6650);
nor U8366 (N_8366,N_7236,N_7433);
nand U8367 (N_8367,N_6783,N_7054);
nor U8368 (N_8368,N_6789,N_6740);
xnor U8369 (N_8369,N_7466,N_7205);
or U8370 (N_8370,N_6895,N_6494);
and U8371 (N_8371,N_6770,N_7405);
xor U8372 (N_8372,N_6706,N_7276);
xnor U8373 (N_8373,N_6311,N_6282);
and U8374 (N_8374,N_7419,N_6737);
and U8375 (N_8375,N_6646,N_6309);
xnor U8376 (N_8376,N_7283,N_6788);
nor U8377 (N_8377,N_6420,N_7225);
nand U8378 (N_8378,N_7136,N_6839);
nand U8379 (N_8379,N_6657,N_7485);
nand U8380 (N_8380,N_6284,N_6799);
or U8381 (N_8381,N_7418,N_6381);
nand U8382 (N_8382,N_6775,N_7391);
nor U8383 (N_8383,N_7033,N_6859);
xnor U8384 (N_8384,N_7406,N_6949);
nor U8385 (N_8385,N_7162,N_6446);
nor U8386 (N_8386,N_6311,N_7323);
xor U8387 (N_8387,N_6891,N_6353);
nand U8388 (N_8388,N_6364,N_6699);
or U8389 (N_8389,N_6955,N_6402);
nor U8390 (N_8390,N_6647,N_7296);
xor U8391 (N_8391,N_6994,N_7130);
nor U8392 (N_8392,N_6326,N_6289);
and U8393 (N_8393,N_6647,N_6970);
or U8394 (N_8394,N_6531,N_6999);
and U8395 (N_8395,N_6766,N_6376);
or U8396 (N_8396,N_6817,N_6282);
nand U8397 (N_8397,N_7406,N_7478);
nor U8398 (N_8398,N_6670,N_7319);
nand U8399 (N_8399,N_7241,N_6415);
and U8400 (N_8400,N_7071,N_6323);
nor U8401 (N_8401,N_6559,N_6795);
nor U8402 (N_8402,N_7224,N_6436);
nand U8403 (N_8403,N_7045,N_7463);
and U8404 (N_8404,N_7454,N_6549);
xor U8405 (N_8405,N_7064,N_7192);
xnor U8406 (N_8406,N_6369,N_6930);
or U8407 (N_8407,N_6984,N_6256);
nand U8408 (N_8408,N_6634,N_6639);
nor U8409 (N_8409,N_6261,N_7343);
xor U8410 (N_8410,N_7482,N_6279);
nor U8411 (N_8411,N_6578,N_7390);
or U8412 (N_8412,N_6252,N_6463);
or U8413 (N_8413,N_7072,N_6582);
or U8414 (N_8414,N_7487,N_6776);
nand U8415 (N_8415,N_6596,N_6923);
xnor U8416 (N_8416,N_6537,N_6626);
nor U8417 (N_8417,N_6376,N_6655);
or U8418 (N_8418,N_6619,N_7308);
nor U8419 (N_8419,N_7417,N_6376);
nor U8420 (N_8420,N_7249,N_7286);
or U8421 (N_8421,N_6905,N_7064);
nand U8422 (N_8422,N_7050,N_6536);
xnor U8423 (N_8423,N_7377,N_7099);
nor U8424 (N_8424,N_6528,N_6653);
and U8425 (N_8425,N_7169,N_6918);
nand U8426 (N_8426,N_6600,N_7434);
or U8427 (N_8427,N_6455,N_6491);
xnor U8428 (N_8428,N_6682,N_6717);
xor U8429 (N_8429,N_7039,N_6547);
and U8430 (N_8430,N_6320,N_6647);
or U8431 (N_8431,N_6607,N_6580);
or U8432 (N_8432,N_6919,N_6958);
or U8433 (N_8433,N_6398,N_7348);
nand U8434 (N_8434,N_6341,N_7166);
nand U8435 (N_8435,N_7180,N_6731);
nand U8436 (N_8436,N_7329,N_6562);
and U8437 (N_8437,N_7470,N_6499);
and U8438 (N_8438,N_7303,N_7094);
or U8439 (N_8439,N_7207,N_6798);
nand U8440 (N_8440,N_6565,N_6897);
and U8441 (N_8441,N_7348,N_6771);
nor U8442 (N_8442,N_6829,N_6453);
and U8443 (N_8443,N_6395,N_6838);
nor U8444 (N_8444,N_7404,N_6322);
nand U8445 (N_8445,N_6904,N_6472);
xnor U8446 (N_8446,N_6606,N_7091);
nor U8447 (N_8447,N_6560,N_7453);
xnor U8448 (N_8448,N_6598,N_7154);
nand U8449 (N_8449,N_6289,N_6679);
nor U8450 (N_8450,N_6521,N_7178);
and U8451 (N_8451,N_6902,N_6331);
xnor U8452 (N_8452,N_6370,N_6774);
nor U8453 (N_8453,N_6312,N_7231);
xor U8454 (N_8454,N_7311,N_6730);
xnor U8455 (N_8455,N_7352,N_7326);
and U8456 (N_8456,N_7289,N_6844);
nor U8457 (N_8457,N_6796,N_6630);
nor U8458 (N_8458,N_6558,N_7232);
xor U8459 (N_8459,N_6758,N_7057);
nor U8460 (N_8460,N_6649,N_7121);
or U8461 (N_8461,N_7122,N_6488);
nand U8462 (N_8462,N_6535,N_7309);
and U8463 (N_8463,N_7226,N_6986);
or U8464 (N_8464,N_7056,N_7231);
nand U8465 (N_8465,N_7413,N_6606);
and U8466 (N_8466,N_7093,N_7321);
nor U8467 (N_8467,N_7432,N_7253);
nand U8468 (N_8468,N_6507,N_6501);
or U8469 (N_8469,N_6536,N_6893);
nand U8470 (N_8470,N_6974,N_6408);
or U8471 (N_8471,N_7335,N_7219);
nand U8472 (N_8472,N_7198,N_7444);
and U8473 (N_8473,N_6312,N_6938);
nor U8474 (N_8474,N_6606,N_7209);
and U8475 (N_8475,N_7424,N_6426);
xor U8476 (N_8476,N_6925,N_7016);
nor U8477 (N_8477,N_7358,N_7061);
nor U8478 (N_8478,N_6783,N_6828);
nor U8479 (N_8479,N_6834,N_6345);
nor U8480 (N_8480,N_7454,N_6910);
nand U8481 (N_8481,N_6714,N_7020);
nor U8482 (N_8482,N_6564,N_7033);
nor U8483 (N_8483,N_6500,N_6358);
xnor U8484 (N_8484,N_6934,N_6753);
and U8485 (N_8485,N_7196,N_6292);
and U8486 (N_8486,N_6377,N_6904);
or U8487 (N_8487,N_6621,N_6446);
and U8488 (N_8488,N_6551,N_7461);
and U8489 (N_8489,N_6569,N_7338);
nand U8490 (N_8490,N_7128,N_7466);
nor U8491 (N_8491,N_7172,N_7015);
and U8492 (N_8492,N_7435,N_6535);
nand U8493 (N_8493,N_6472,N_6845);
or U8494 (N_8494,N_6592,N_6620);
nand U8495 (N_8495,N_6939,N_6961);
or U8496 (N_8496,N_6978,N_7041);
and U8497 (N_8497,N_7374,N_6798);
nor U8498 (N_8498,N_6660,N_7019);
or U8499 (N_8499,N_6279,N_7489);
and U8500 (N_8500,N_7101,N_6709);
or U8501 (N_8501,N_7218,N_6601);
nand U8502 (N_8502,N_6617,N_6785);
and U8503 (N_8503,N_6903,N_7192);
nand U8504 (N_8504,N_7332,N_6774);
and U8505 (N_8505,N_7481,N_6624);
or U8506 (N_8506,N_6898,N_6847);
nor U8507 (N_8507,N_6672,N_7175);
and U8508 (N_8508,N_6981,N_6975);
nand U8509 (N_8509,N_6877,N_6565);
and U8510 (N_8510,N_7346,N_7476);
nand U8511 (N_8511,N_6375,N_6955);
and U8512 (N_8512,N_6573,N_7088);
or U8513 (N_8513,N_6993,N_6302);
nand U8514 (N_8514,N_6396,N_7417);
nor U8515 (N_8515,N_7458,N_6457);
nor U8516 (N_8516,N_7146,N_6433);
nor U8517 (N_8517,N_6622,N_7205);
and U8518 (N_8518,N_7336,N_6951);
nand U8519 (N_8519,N_6734,N_6923);
nor U8520 (N_8520,N_7415,N_6776);
xor U8521 (N_8521,N_6591,N_6851);
nand U8522 (N_8522,N_7294,N_7126);
nand U8523 (N_8523,N_7090,N_7123);
xor U8524 (N_8524,N_6756,N_7212);
nor U8525 (N_8525,N_6951,N_6319);
and U8526 (N_8526,N_6367,N_6379);
xor U8527 (N_8527,N_7485,N_6698);
and U8528 (N_8528,N_6520,N_7446);
xor U8529 (N_8529,N_6928,N_7131);
or U8530 (N_8530,N_6825,N_7438);
nand U8531 (N_8531,N_6473,N_6545);
xor U8532 (N_8532,N_6810,N_7271);
and U8533 (N_8533,N_6528,N_6267);
nor U8534 (N_8534,N_7401,N_6567);
xnor U8535 (N_8535,N_6584,N_6492);
or U8536 (N_8536,N_6742,N_6965);
or U8537 (N_8537,N_7304,N_6705);
or U8538 (N_8538,N_7424,N_6268);
xor U8539 (N_8539,N_6876,N_7305);
nand U8540 (N_8540,N_7094,N_7417);
nor U8541 (N_8541,N_6811,N_6973);
and U8542 (N_8542,N_6480,N_6398);
nor U8543 (N_8543,N_6310,N_7272);
nand U8544 (N_8544,N_6265,N_6506);
nor U8545 (N_8545,N_7006,N_7257);
xor U8546 (N_8546,N_7254,N_6708);
and U8547 (N_8547,N_6759,N_6776);
xor U8548 (N_8548,N_6412,N_6938);
nand U8549 (N_8549,N_6872,N_6376);
and U8550 (N_8550,N_7126,N_7323);
xor U8551 (N_8551,N_7162,N_6586);
and U8552 (N_8552,N_6903,N_6620);
nand U8553 (N_8553,N_7175,N_6641);
nand U8554 (N_8554,N_6485,N_6947);
nor U8555 (N_8555,N_6410,N_7053);
and U8556 (N_8556,N_6573,N_7069);
nand U8557 (N_8557,N_6448,N_7251);
nor U8558 (N_8558,N_7215,N_7155);
or U8559 (N_8559,N_6421,N_6908);
nand U8560 (N_8560,N_7353,N_7262);
nor U8561 (N_8561,N_6658,N_6625);
nor U8562 (N_8562,N_6816,N_6395);
or U8563 (N_8563,N_7084,N_6680);
xnor U8564 (N_8564,N_7454,N_6923);
nor U8565 (N_8565,N_6901,N_6457);
and U8566 (N_8566,N_6539,N_6987);
xnor U8567 (N_8567,N_6820,N_7481);
and U8568 (N_8568,N_7267,N_6453);
nand U8569 (N_8569,N_7235,N_6615);
xnor U8570 (N_8570,N_6507,N_6576);
and U8571 (N_8571,N_6672,N_7147);
or U8572 (N_8572,N_7025,N_6825);
or U8573 (N_8573,N_6399,N_6421);
nor U8574 (N_8574,N_6541,N_6629);
or U8575 (N_8575,N_7436,N_6959);
and U8576 (N_8576,N_7024,N_6493);
nand U8577 (N_8577,N_7005,N_6573);
or U8578 (N_8578,N_7479,N_7063);
nor U8579 (N_8579,N_7428,N_7277);
and U8580 (N_8580,N_6805,N_7158);
xnor U8581 (N_8581,N_6302,N_6310);
nor U8582 (N_8582,N_6955,N_7134);
nor U8583 (N_8583,N_7378,N_7239);
nor U8584 (N_8584,N_6331,N_6302);
xor U8585 (N_8585,N_7157,N_6286);
and U8586 (N_8586,N_6909,N_7092);
and U8587 (N_8587,N_7016,N_7061);
xor U8588 (N_8588,N_6341,N_6388);
xor U8589 (N_8589,N_6430,N_7178);
xnor U8590 (N_8590,N_6899,N_6699);
nor U8591 (N_8591,N_6268,N_6435);
nand U8592 (N_8592,N_6757,N_6932);
xor U8593 (N_8593,N_6533,N_6769);
nor U8594 (N_8594,N_7073,N_6567);
nand U8595 (N_8595,N_6444,N_7457);
xor U8596 (N_8596,N_6321,N_7375);
xor U8597 (N_8597,N_7377,N_6683);
nor U8598 (N_8598,N_7098,N_7170);
and U8599 (N_8599,N_6733,N_6470);
nor U8600 (N_8600,N_7457,N_6460);
or U8601 (N_8601,N_6360,N_6953);
or U8602 (N_8602,N_7053,N_6937);
or U8603 (N_8603,N_6387,N_6780);
or U8604 (N_8604,N_6419,N_7408);
xnor U8605 (N_8605,N_6687,N_6554);
or U8606 (N_8606,N_6546,N_6971);
and U8607 (N_8607,N_6305,N_6787);
and U8608 (N_8608,N_6815,N_6869);
or U8609 (N_8609,N_7014,N_7327);
and U8610 (N_8610,N_6276,N_6523);
nor U8611 (N_8611,N_6850,N_6274);
nor U8612 (N_8612,N_6703,N_6698);
nor U8613 (N_8613,N_7048,N_7192);
nor U8614 (N_8614,N_7269,N_6750);
and U8615 (N_8615,N_7341,N_6780);
nand U8616 (N_8616,N_6342,N_7198);
nor U8617 (N_8617,N_6772,N_7148);
and U8618 (N_8618,N_6861,N_6462);
xor U8619 (N_8619,N_6954,N_7471);
nor U8620 (N_8620,N_7136,N_7263);
nand U8621 (N_8621,N_6262,N_6319);
nand U8622 (N_8622,N_7377,N_6834);
xor U8623 (N_8623,N_6737,N_6695);
or U8624 (N_8624,N_6833,N_6617);
and U8625 (N_8625,N_6355,N_6623);
nand U8626 (N_8626,N_7270,N_6851);
or U8627 (N_8627,N_7113,N_6283);
nor U8628 (N_8628,N_6750,N_6906);
nand U8629 (N_8629,N_6756,N_7265);
or U8630 (N_8630,N_6990,N_6356);
and U8631 (N_8631,N_7092,N_7104);
xnor U8632 (N_8632,N_6307,N_6721);
nand U8633 (N_8633,N_7172,N_6732);
and U8634 (N_8634,N_6687,N_6551);
and U8635 (N_8635,N_7236,N_6719);
nor U8636 (N_8636,N_6344,N_7029);
or U8637 (N_8637,N_7188,N_6596);
or U8638 (N_8638,N_6282,N_7478);
or U8639 (N_8639,N_6485,N_7404);
or U8640 (N_8640,N_7174,N_6811);
xor U8641 (N_8641,N_6444,N_6901);
nor U8642 (N_8642,N_7475,N_7085);
or U8643 (N_8643,N_6495,N_7412);
nand U8644 (N_8644,N_6753,N_6421);
or U8645 (N_8645,N_6824,N_6924);
nor U8646 (N_8646,N_7016,N_6936);
nor U8647 (N_8647,N_6767,N_7110);
xor U8648 (N_8648,N_6561,N_6978);
xor U8649 (N_8649,N_6569,N_6491);
nor U8650 (N_8650,N_7299,N_6848);
and U8651 (N_8651,N_6352,N_7049);
and U8652 (N_8652,N_6713,N_7493);
nand U8653 (N_8653,N_7187,N_7189);
nor U8654 (N_8654,N_6926,N_6846);
nor U8655 (N_8655,N_6558,N_6868);
xor U8656 (N_8656,N_7295,N_6618);
nand U8657 (N_8657,N_7165,N_6476);
or U8658 (N_8658,N_6376,N_6946);
nand U8659 (N_8659,N_6429,N_6891);
nand U8660 (N_8660,N_6587,N_6469);
nand U8661 (N_8661,N_6722,N_6374);
xnor U8662 (N_8662,N_6294,N_6316);
xor U8663 (N_8663,N_6291,N_6251);
or U8664 (N_8664,N_6793,N_6689);
xor U8665 (N_8665,N_6885,N_6828);
nand U8666 (N_8666,N_7138,N_7406);
or U8667 (N_8667,N_6645,N_7184);
and U8668 (N_8668,N_6975,N_6492);
nand U8669 (N_8669,N_7200,N_7322);
nor U8670 (N_8670,N_6689,N_6562);
or U8671 (N_8671,N_6660,N_6376);
and U8672 (N_8672,N_7130,N_6339);
nor U8673 (N_8673,N_6583,N_7042);
and U8674 (N_8674,N_6659,N_6386);
and U8675 (N_8675,N_6789,N_7137);
nand U8676 (N_8676,N_7455,N_7245);
nor U8677 (N_8677,N_6859,N_7233);
xor U8678 (N_8678,N_7455,N_6928);
xnor U8679 (N_8679,N_6633,N_6547);
and U8680 (N_8680,N_7260,N_6681);
nor U8681 (N_8681,N_7043,N_7240);
or U8682 (N_8682,N_6266,N_6542);
nand U8683 (N_8683,N_7092,N_6839);
and U8684 (N_8684,N_6913,N_6666);
nor U8685 (N_8685,N_6614,N_6517);
nand U8686 (N_8686,N_6605,N_6403);
xor U8687 (N_8687,N_6342,N_7277);
and U8688 (N_8688,N_6898,N_7020);
xnor U8689 (N_8689,N_7369,N_7185);
and U8690 (N_8690,N_6651,N_7143);
and U8691 (N_8691,N_6722,N_6849);
and U8692 (N_8692,N_6376,N_6328);
or U8693 (N_8693,N_6748,N_6261);
nand U8694 (N_8694,N_7151,N_6624);
nand U8695 (N_8695,N_7166,N_6822);
xor U8696 (N_8696,N_6265,N_7059);
and U8697 (N_8697,N_7188,N_7143);
and U8698 (N_8698,N_7166,N_7014);
and U8699 (N_8699,N_7076,N_7280);
xnor U8700 (N_8700,N_7026,N_7412);
xor U8701 (N_8701,N_6314,N_7384);
or U8702 (N_8702,N_6903,N_6283);
and U8703 (N_8703,N_6428,N_7018);
or U8704 (N_8704,N_7226,N_7422);
nand U8705 (N_8705,N_7020,N_6619);
xnor U8706 (N_8706,N_6781,N_7164);
nand U8707 (N_8707,N_6593,N_6463);
xor U8708 (N_8708,N_6460,N_7064);
xnor U8709 (N_8709,N_6934,N_7336);
and U8710 (N_8710,N_7174,N_6557);
nor U8711 (N_8711,N_6616,N_6717);
nor U8712 (N_8712,N_7118,N_6478);
and U8713 (N_8713,N_6463,N_6923);
nor U8714 (N_8714,N_7468,N_7422);
or U8715 (N_8715,N_6299,N_7065);
or U8716 (N_8716,N_7119,N_7360);
nand U8717 (N_8717,N_7446,N_7223);
nor U8718 (N_8718,N_7265,N_6295);
and U8719 (N_8719,N_7180,N_6410);
or U8720 (N_8720,N_6389,N_7210);
xnor U8721 (N_8721,N_6562,N_7182);
nand U8722 (N_8722,N_7439,N_6611);
xnor U8723 (N_8723,N_6767,N_7135);
xnor U8724 (N_8724,N_6772,N_6412);
nand U8725 (N_8725,N_6393,N_6508);
nand U8726 (N_8726,N_7494,N_6814);
nor U8727 (N_8727,N_6321,N_6990);
nor U8728 (N_8728,N_6435,N_7142);
and U8729 (N_8729,N_6515,N_7401);
and U8730 (N_8730,N_7341,N_7087);
xnor U8731 (N_8731,N_7347,N_6422);
and U8732 (N_8732,N_6982,N_6966);
nand U8733 (N_8733,N_6924,N_6833);
or U8734 (N_8734,N_6890,N_6963);
nand U8735 (N_8735,N_7182,N_6770);
nor U8736 (N_8736,N_6280,N_6330);
nand U8737 (N_8737,N_7379,N_7300);
or U8738 (N_8738,N_7039,N_6625);
xnor U8739 (N_8739,N_7153,N_6291);
xnor U8740 (N_8740,N_6674,N_6727);
or U8741 (N_8741,N_7249,N_6311);
and U8742 (N_8742,N_7127,N_7174);
nor U8743 (N_8743,N_6370,N_7159);
xnor U8744 (N_8744,N_6856,N_7337);
and U8745 (N_8745,N_6455,N_7261);
nor U8746 (N_8746,N_6452,N_6703);
nor U8747 (N_8747,N_7380,N_6364);
nand U8748 (N_8748,N_6380,N_7104);
or U8749 (N_8749,N_7164,N_7435);
or U8750 (N_8750,N_7552,N_7683);
and U8751 (N_8751,N_8022,N_8217);
nand U8752 (N_8752,N_8606,N_7528);
and U8753 (N_8753,N_7847,N_8548);
nand U8754 (N_8754,N_8107,N_8491);
xor U8755 (N_8755,N_8525,N_8631);
nand U8756 (N_8756,N_7563,N_8578);
or U8757 (N_8757,N_8241,N_7742);
and U8758 (N_8758,N_8378,N_8070);
nand U8759 (N_8759,N_7638,N_8636);
or U8760 (N_8760,N_7749,N_8713);
nand U8761 (N_8761,N_8718,N_8674);
or U8762 (N_8762,N_8212,N_8392);
nor U8763 (N_8763,N_7519,N_8287);
and U8764 (N_8764,N_8711,N_8239);
and U8765 (N_8765,N_8366,N_8387);
nand U8766 (N_8766,N_8295,N_7549);
or U8767 (N_8767,N_8439,N_8633);
or U8768 (N_8768,N_8495,N_8467);
xor U8769 (N_8769,N_7670,N_7934);
xnor U8770 (N_8770,N_7983,N_7659);
and U8771 (N_8771,N_8486,N_7871);
nor U8772 (N_8772,N_8357,N_7759);
or U8773 (N_8773,N_7789,N_8659);
nand U8774 (N_8774,N_8140,N_8654);
or U8775 (N_8775,N_7525,N_8410);
or U8776 (N_8776,N_7610,N_7617);
nor U8777 (N_8777,N_8585,N_8211);
or U8778 (N_8778,N_8247,N_8501);
xor U8779 (N_8779,N_8530,N_7974);
nand U8780 (N_8780,N_7795,N_8675);
or U8781 (N_8781,N_8651,N_8114);
nor U8782 (N_8782,N_7529,N_8167);
xor U8783 (N_8783,N_8448,N_8516);
xnor U8784 (N_8784,N_8279,N_7567);
nor U8785 (N_8785,N_7600,N_8417);
and U8786 (N_8786,N_7671,N_7856);
and U8787 (N_8787,N_7786,N_7596);
nor U8788 (N_8788,N_8632,N_8215);
xnor U8789 (N_8789,N_8331,N_7655);
or U8790 (N_8790,N_8595,N_8619);
and U8791 (N_8791,N_8584,N_7571);
nor U8792 (N_8792,N_8009,N_7961);
or U8793 (N_8793,N_8480,N_8351);
or U8794 (N_8794,N_7783,N_7740);
or U8795 (N_8795,N_7521,N_8560);
and U8796 (N_8796,N_8028,N_7711);
xnor U8797 (N_8797,N_8268,N_7686);
or U8798 (N_8798,N_8608,N_8278);
and U8799 (N_8799,N_8669,N_8552);
xor U8800 (N_8800,N_7630,N_8405);
or U8801 (N_8801,N_8151,N_8094);
nand U8802 (N_8802,N_8186,N_7952);
nor U8803 (N_8803,N_7864,N_7574);
or U8804 (N_8804,N_8628,N_7717);
nand U8805 (N_8805,N_8492,N_8103);
xnor U8806 (N_8806,N_8526,N_8709);
or U8807 (N_8807,N_8313,N_7819);
or U8808 (N_8808,N_8593,N_8171);
and U8809 (N_8809,N_8712,N_7774);
or U8810 (N_8810,N_8087,N_8590);
and U8811 (N_8811,N_7784,N_7718);
xor U8812 (N_8812,N_7545,N_7603);
and U8813 (N_8813,N_8235,N_7910);
xor U8814 (N_8814,N_8393,N_7908);
nor U8815 (N_8815,N_7980,N_8170);
xnor U8816 (N_8816,N_7672,N_8722);
and U8817 (N_8817,N_8677,N_8250);
or U8818 (N_8818,N_8589,N_8510);
xor U8819 (N_8819,N_8728,N_8281);
or U8820 (N_8820,N_8451,N_8591);
or U8821 (N_8821,N_7623,N_8284);
nand U8822 (N_8822,N_8273,N_8721);
nand U8823 (N_8823,N_7767,N_7699);
or U8824 (N_8824,N_7509,N_7870);
and U8825 (N_8825,N_8242,N_7769);
and U8826 (N_8826,N_8213,N_7531);
nand U8827 (N_8827,N_7828,N_8694);
nor U8828 (N_8828,N_8611,N_8574);
and U8829 (N_8829,N_7933,N_8206);
nand U8830 (N_8830,N_7932,N_7682);
and U8831 (N_8831,N_7534,N_7809);
or U8832 (N_8832,N_7734,N_8688);
nor U8833 (N_8833,N_7698,N_7821);
nor U8834 (N_8834,N_8592,N_8325);
nor U8835 (N_8835,N_8126,N_7736);
or U8836 (N_8836,N_8164,N_8524);
nor U8837 (N_8837,N_7752,N_7562);
and U8838 (N_8838,N_8081,N_8428);
xor U8839 (N_8839,N_7693,N_8068);
xnor U8840 (N_8840,N_8230,N_8749);
nand U8841 (N_8841,N_8576,N_7741);
or U8842 (N_8842,N_8475,N_8187);
and U8843 (N_8843,N_7595,N_8104);
nand U8844 (N_8844,N_8105,N_8457);
or U8845 (N_8845,N_8293,N_8607);
nor U8846 (N_8846,N_8263,N_8384);
xnor U8847 (N_8847,N_7660,N_8733);
nor U8848 (N_8848,N_8562,N_8108);
nand U8849 (N_8849,N_7855,N_8265);
and U8850 (N_8850,N_8182,N_8536);
or U8851 (N_8851,N_7522,N_7515);
nand U8852 (N_8852,N_7707,N_7937);
nor U8853 (N_8853,N_7581,N_8412);
and U8854 (N_8854,N_7559,N_8442);
nand U8855 (N_8855,N_7973,N_8046);
or U8856 (N_8856,N_8080,N_8414);
xnor U8857 (N_8857,N_7653,N_8155);
nor U8858 (N_8858,N_7520,N_8460);
nor U8859 (N_8859,N_8237,N_8122);
nand U8860 (N_8860,N_8647,N_8408);
and U8861 (N_8861,N_8161,N_7625);
and U8862 (N_8862,N_8653,N_8021);
nand U8863 (N_8863,N_7613,N_7508);
nor U8864 (N_8864,N_7620,N_8554);
xor U8865 (N_8865,N_7743,N_7650);
nand U8866 (N_8866,N_7994,N_7942);
nor U8867 (N_8867,N_8493,N_7920);
and U8868 (N_8868,N_8544,N_8031);
xor U8869 (N_8869,N_8558,N_8372);
nand U8870 (N_8870,N_8111,N_7662);
xnor U8871 (N_8871,N_7967,N_7502);
nand U8872 (N_8872,N_7641,N_8397);
xor U8873 (N_8873,N_7888,N_8737);
nor U8874 (N_8874,N_8563,N_7751);
or U8875 (N_8875,N_7690,N_8542);
or U8876 (N_8876,N_8341,N_8676);
and U8877 (N_8877,N_8515,N_7703);
nand U8878 (N_8878,N_7730,N_8478);
or U8879 (N_8879,N_7962,N_7543);
xor U8880 (N_8880,N_7532,N_7599);
nand U8881 (N_8881,N_8184,N_7516);
xor U8882 (N_8882,N_7550,N_7723);
nor U8883 (N_8883,N_8090,N_7573);
and U8884 (N_8884,N_7503,N_8280);
nor U8885 (N_8885,N_8534,N_7527);
xor U8886 (N_8886,N_8540,N_7756);
xor U8887 (N_8887,N_8277,N_8024);
or U8888 (N_8888,N_7913,N_7796);
or U8889 (N_8889,N_7824,N_8599);
and U8890 (N_8890,N_8233,N_8613);
xnor U8891 (N_8891,N_7647,N_7981);
nor U8892 (N_8892,N_8203,N_8565);
xor U8893 (N_8893,N_7719,N_7547);
nor U8894 (N_8894,N_8400,N_7646);
and U8895 (N_8895,N_7586,N_7624);
or U8896 (N_8896,N_8625,N_7712);
nor U8897 (N_8897,N_8052,N_7854);
xor U8898 (N_8898,N_7689,N_8257);
and U8899 (N_8899,N_7897,N_7793);
or U8900 (N_8900,N_7523,N_8708);
nor U8901 (N_8901,N_8059,N_7544);
nand U8902 (N_8902,N_8577,N_8401);
nor U8903 (N_8903,N_7926,N_8190);
and U8904 (N_8904,N_8152,N_7969);
xnor U8905 (N_8905,N_8143,N_8468);
nand U8906 (N_8906,N_8588,N_7936);
and U8907 (N_8907,N_8739,N_8719);
nor U8908 (N_8908,N_7801,N_7797);
nor U8909 (N_8909,N_7989,N_8264);
or U8910 (N_8910,N_7998,N_7679);
nor U8911 (N_8911,N_7958,N_8083);
nor U8912 (N_8912,N_8707,N_8173);
nor U8913 (N_8913,N_8394,N_8621);
nand U8914 (N_8914,N_8504,N_7884);
nand U8915 (N_8915,N_7565,N_7606);
nor U8916 (N_8916,N_7745,N_7914);
or U8917 (N_8917,N_8147,N_8160);
and U8918 (N_8918,N_8195,N_8244);
or U8919 (N_8919,N_7852,N_7735);
and U8920 (N_8920,N_8289,N_8375);
xor U8921 (N_8921,N_7947,N_7637);
nand U8922 (N_8922,N_8359,N_7964);
nor U8923 (N_8923,N_8395,N_8370);
or U8924 (N_8924,N_7568,N_7744);
nor U8925 (N_8925,N_8096,N_7510);
or U8926 (N_8926,N_7953,N_7696);
and U8927 (N_8927,N_7803,N_8121);
nor U8928 (N_8928,N_7949,N_7765);
xnor U8929 (N_8929,N_8652,N_7772);
and U8930 (N_8930,N_7911,N_8715);
and U8931 (N_8931,N_8150,N_7838);
xnor U8932 (N_8932,N_8000,N_8041);
xnor U8933 (N_8933,N_8288,N_8483);
or U8934 (N_8934,N_7817,N_8145);
or U8935 (N_8935,N_8730,N_7538);
nor U8936 (N_8936,N_8700,N_7564);
or U8937 (N_8937,N_8455,N_8696);
nor U8938 (N_8938,N_8533,N_8686);
nand U8939 (N_8939,N_7748,N_8435);
or U8940 (N_8940,N_7731,N_7669);
nor U8941 (N_8941,N_8343,N_8680);
nand U8942 (N_8942,N_8354,N_7915);
and U8943 (N_8943,N_7780,N_7808);
nand U8944 (N_8944,N_8380,N_7835);
xor U8945 (N_8945,N_8610,N_8522);
xnor U8946 (N_8946,N_8340,N_7588);
nor U8947 (N_8947,N_8477,N_8386);
and U8948 (N_8948,N_7592,N_8500);
and U8949 (N_8949,N_8060,N_8687);
nor U8950 (N_8950,N_8208,N_8376);
and U8951 (N_8951,N_8396,N_8693);
nor U8952 (N_8952,N_8673,N_7940);
xor U8953 (N_8953,N_7901,N_8579);
nand U8954 (N_8954,N_7651,N_8446);
nand U8955 (N_8955,N_8466,N_7541);
nand U8956 (N_8956,N_8598,N_8317);
xnor U8957 (N_8957,N_7733,N_8229);
or U8958 (N_8958,N_7939,N_8640);
nor U8959 (N_8959,N_8614,N_8678);
nor U8960 (N_8960,N_7955,N_8745);
nor U8961 (N_8961,N_8472,N_7771);
nand U8962 (N_8962,N_8481,N_8447);
nand U8963 (N_8963,N_8617,N_7916);
or U8964 (N_8964,N_8549,N_8049);
nand U8965 (N_8965,N_8639,N_8272);
nor U8966 (N_8966,N_8645,N_7566);
or U8967 (N_8967,N_8546,N_8535);
or U8968 (N_8968,N_8063,N_8095);
or U8969 (N_8969,N_7825,N_7688);
nor U8970 (N_8970,N_8314,N_8443);
xor U8971 (N_8971,N_8283,N_8260);
nor U8972 (N_8972,N_8261,N_8307);
or U8973 (N_8973,N_8561,N_7880);
xnor U8974 (N_8974,N_7601,N_7876);
xor U8975 (N_8975,N_7676,N_8110);
nor U8976 (N_8976,N_7526,N_8130);
xor U8977 (N_8977,N_7842,N_7879);
nand U8978 (N_8978,N_8113,N_8403);
nor U8979 (N_8979,N_8334,N_8418);
xor U8980 (N_8980,N_8106,N_8587);
xnor U8981 (N_8981,N_8519,N_8583);
nor U8982 (N_8982,N_7822,N_7826);
nor U8983 (N_8983,N_8603,N_8484);
or U8984 (N_8984,N_8499,N_8169);
and U8985 (N_8985,N_8748,N_8197);
nand U8986 (N_8986,N_8228,N_7995);
nand U8987 (N_8987,N_8421,N_7997);
xnor U8988 (N_8988,N_8138,N_8176);
xor U8989 (N_8989,N_8627,N_8541);
xnor U8990 (N_8990,N_8048,N_7965);
xor U8991 (N_8991,N_7839,N_8142);
nor U8992 (N_8992,N_8348,N_7645);
nand U8993 (N_8993,N_7881,N_8685);
or U8994 (N_8994,N_8487,N_7999);
and U8995 (N_8995,N_8310,N_7867);
nor U8996 (N_8996,N_8148,N_7984);
and U8997 (N_8997,N_7517,N_8267);
and U8998 (N_8998,N_7773,N_7619);
xnor U8999 (N_8999,N_8178,N_8648);
xnor U9000 (N_9000,N_8315,N_7814);
nor U9001 (N_9001,N_8699,N_8282);
and U9002 (N_9002,N_8181,N_8005);
xor U9003 (N_9003,N_8234,N_8726);
and U9004 (N_9004,N_7979,N_8010);
xor U9005 (N_9005,N_8727,N_8091);
and U9006 (N_9006,N_7874,N_8390);
nand U9007 (N_9007,N_8596,N_7790);
or U9008 (N_9008,N_8124,N_7891);
or U9009 (N_9009,N_7900,N_8259);
or U9010 (N_9010,N_7524,N_8136);
nand U9011 (N_9011,N_8537,N_8735);
nand U9012 (N_9012,N_7572,N_8505);
and U9013 (N_9013,N_8660,N_8638);
and U9014 (N_9014,N_8223,N_7892);
nand U9015 (N_9015,N_8092,N_8471);
or U9016 (N_9016,N_7869,N_8030);
and U9017 (N_9017,N_8053,N_8337);
nand U9018 (N_9018,N_8328,N_7831);
or U9019 (N_9019,N_7678,N_8238);
and U9020 (N_9020,N_7605,N_8255);
or U9021 (N_9021,N_8692,N_7758);
xnor U9022 (N_9022,N_7504,N_7943);
or U9023 (N_9023,N_8612,N_8088);
xor U9024 (N_9024,N_7966,N_8074);
and U9025 (N_9025,N_8129,N_7702);
xor U9026 (N_9026,N_8306,N_7972);
or U9027 (N_9027,N_8600,N_8356);
xor U9028 (N_9028,N_8742,N_7656);
nor U9029 (N_9029,N_8649,N_8637);
nand U9030 (N_9030,N_8523,N_8624);
nor U9031 (N_9031,N_8319,N_7768);
xnor U9032 (N_9032,N_8670,N_7863);
and U9033 (N_9033,N_7763,N_8200);
or U9034 (N_9034,N_8077,N_8123);
or U9035 (N_9035,N_8252,N_8724);
or U9036 (N_9036,N_7704,N_8057);
nor U9037 (N_9037,N_7811,N_8717);
nor U9038 (N_9038,N_8013,N_8346);
xor U9039 (N_9039,N_8427,N_8362);
and U9040 (N_9040,N_8214,N_8275);
and U9041 (N_9041,N_7951,N_8476);
and U9042 (N_9042,N_7557,N_7575);
and U9043 (N_9043,N_8320,N_8019);
or U9044 (N_9044,N_7708,N_7886);
xor U9045 (N_9045,N_8034,N_7957);
and U9046 (N_9046,N_8690,N_8470);
xor U9047 (N_9047,N_7582,N_8342);
or U9048 (N_9048,N_7654,N_7628);
xnor U9049 (N_9049,N_8714,N_8168);
nor U9050 (N_9050,N_7787,N_8665);
or U9051 (N_9051,N_7633,N_7866);
or U9052 (N_9052,N_8672,N_8666);
nor U9053 (N_9053,N_7753,N_8622);
xor U9054 (N_9054,N_7665,N_7629);
nand U9055 (N_9055,N_7830,N_8157);
xnor U9056 (N_9056,N_7976,N_7500);
nand U9057 (N_9057,N_8099,N_8294);
xnor U9058 (N_9058,N_7597,N_8149);
xnor U9059 (N_9059,N_7877,N_8736);
xor U9060 (N_9060,N_8509,N_7858);
nor U9061 (N_9061,N_7561,N_8192);
or U9062 (N_9062,N_8667,N_8365);
and U9063 (N_9063,N_8744,N_7800);
and U9064 (N_9064,N_7627,N_7810);
and U9065 (N_9065,N_8017,N_7697);
nor U9066 (N_9066,N_8299,N_8517);
nor U9067 (N_9067,N_8497,N_8706);
xor U9068 (N_9068,N_8202,N_7829);
and U9069 (N_9069,N_8416,N_8419);
or U9070 (N_9070,N_7899,N_8564);
xnor U9071 (N_9071,N_8508,N_8226);
and U9072 (N_9072,N_8597,N_7945);
nand U9073 (N_9073,N_7583,N_8131);
nand U9074 (N_9074,N_8311,N_8026);
nand U9075 (N_9075,N_8249,N_8389);
nand U9076 (N_9076,N_7542,N_8664);
and U9077 (N_9077,N_7948,N_8703);
nor U9078 (N_9078,N_7579,N_7956);
and U9079 (N_9079,N_8067,N_7590);
and U9080 (N_9080,N_8231,N_7950);
nor U9081 (N_9081,N_8679,N_8322);
or U9082 (N_9082,N_8381,N_8078);
and U9083 (N_9083,N_8605,N_8423);
nor U9084 (N_9084,N_7622,N_7883);
xor U9085 (N_9085,N_7982,N_8165);
or U9086 (N_9086,N_8377,N_7978);
nor U9087 (N_9087,N_8166,N_8082);
or U9088 (N_9088,N_8601,N_8117);
nor U9089 (N_9089,N_7775,N_8566);
nand U9090 (N_9090,N_8144,N_7992);
and U9091 (N_9091,N_8368,N_8286);
and U9092 (N_9092,N_7692,N_7584);
nand U9093 (N_9093,N_8489,N_7918);
nand U9094 (N_9094,N_7668,N_8253);
and U9095 (N_9095,N_8004,N_7889);
xnor U9096 (N_9096,N_8269,N_7875);
and U9097 (N_9097,N_8236,N_8440);
or U9098 (N_9098,N_8058,N_8568);
nand U9099 (N_9099,N_7694,N_7539);
or U9100 (N_9100,N_8518,N_8188);
nor U9101 (N_9101,N_8141,N_8120);
xor U9102 (N_9102,N_8032,N_7776);
nor U9103 (N_9103,N_8623,N_7987);
nor U9104 (N_9104,N_7677,N_7558);
or U9105 (N_9105,N_8037,N_8602);
xor U9106 (N_9106,N_7546,N_8023);
nor U9107 (N_9107,N_7798,N_7639);
nor U9108 (N_9108,N_7805,N_7709);
and U9109 (N_9109,N_7827,N_7700);
xnor U9110 (N_9110,N_7729,N_7804);
nand U9111 (N_9111,N_8040,N_7815);
and U9112 (N_9112,N_8634,N_7816);
or U9113 (N_9113,N_7882,N_7684);
xnor U9114 (N_9114,N_8207,N_8291);
and U9115 (N_9115,N_7673,N_8521);
nor U9116 (N_9116,N_8333,N_7921);
xor U9117 (N_9117,N_8452,N_8329);
or U9118 (N_9118,N_8115,N_8352);
xnor U9119 (N_9119,N_8547,N_7928);
xor U9120 (N_9120,N_8292,N_8704);
or U9121 (N_9121,N_8404,N_8001);
nor U9122 (N_9122,N_8066,N_8641);
and U9123 (N_9123,N_8459,N_7924);
nand U9124 (N_9124,N_7537,N_8445);
nor U9125 (N_9125,N_8135,N_8132);
xnor U9126 (N_9126,N_8569,N_8681);
nor U9127 (N_9127,N_8650,N_7925);
nand U9128 (N_9128,N_7577,N_8006);
nor U9129 (N_9129,N_8513,N_7548);
and U9130 (N_9130,N_7813,N_8020);
nor U9131 (N_9131,N_7991,N_7865);
nand U9132 (N_9132,N_8551,N_8671);
nor U9133 (N_9133,N_8646,N_8185);
or U9134 (N_9134,N_8553,N_8434);
xnor U9135 (N_9135,N_7674,N_7781);
nand U9136 (N_9136,N_8199,N_8301);
nand U9137 (N_9137,N_8520,N_7929);
and U9138 (N_9138,N_8227,N_7975);
xor U9139 (N_9139,N_8304,N_7501);
xnor U9140 (N_9140,N_8353,N_8454);
nand U9141 (N_9141,N_7860,N_8193);
or U9142 (N_9142,N_8201,N_7608);
nand U9143 (N_9143,N_8413,N_8327);
xnor U9144 (N_9144,N_7612,N_8490);
nand U9145 (N_9145,N_8084,N_7853);
or U9146 (N_9146,N_7885,N_8629);
xnor U9147 (N_9147,N_7507,N_7642);
xor U9148 (N_9148,N_8011,N_7512);
and U9149 (N_9149,N_8433,N_7553);
nand U9150 (N_9150,N_7661,N_8134);
nor U9151 (N_9151,N_8258,N_7836);
xor U9152 (N_9152,N_8321,N_8496);
nand U9153 (N_9153,N_8731,N_8016);
nor U9154 (N_9154,N_8620,N_8543);
nor U9155 (N_9155,N_8642,N_7941);
and U9156 (N_9156,N_8316,N_7841);
xor U9157 (N_9157,N_8430,N_8159);
and U9158 (N_9158,N_8248,N_8385);
nand U9159 (N_9159,N_8586,N_7954);
and U9160 (N_9160,N_8179,N_7833);
nand U9161 (N_9161,N_8725,N_7862);
xor U9162 (N_9162,N_7580,N_8374);
nor U9163 (N_9163,N_8338,N_8180);
or U9164 (N_9164,N_8545,N_7585);
nand U9165 (N_9165,N_7513,N_8514);
xnor U9166 (N_9166,N_8008,N_8172);
or U9167 (N_9167,N_8065,N_7878);
nand U9168 (N_9168,N_8133,N_8689);
nor U9169 (N_9169,N_8409,N_8100);
nor U9170 (N_9170,N_8204,N_8656);
nor U9171 (N_9171,N_8324,N_8256);
or U9172 (N_9172,N_7578,N_7777);
nor U9173 (N_9173,N_7907,N_8086);
nor U9174 (N_9174,N_7701,N_7663);
nand U9175 (N_9175,N_7850,N_7687);
xor U9176 (N_9176,N_8661,N_8163);
and U9177 (N_9177,N_7664,N_8146);
or U9178 (N_9178,N_8474,N_7766);
nor U9179 (N_9179,N_7857,N_7594);
and U9180 (N_9180,N_7963,N_8194);
nand U9181 (N_9181,N_7898,N_8003);
nand U9182 (N_9182,N_8093,N_8644);
nand U9183 (N_9183,N_8507,N_8018);
xnor U9184 (N_9184,N_8436,N_7667);
or U9185 (N_9185,N_7569,N_7923);
nor U9186 (N_9186,N_8720,N_8738);
and U9187 (N_9187,N_8684,N_8240);
and U9188 (N_9188,N_8266,N_8101);
xnor U9189 (N_9189,N_7611,N_7761);
or U9190 (N_9190,N_7903,N_8027);
nor U9191 (N_9191,N_8038,N_7778);
nor U9192 (N_9192,N_7779,N_8503);
nand U9193 (N_9193,N_7649,N_8399);
xor U9194 (N_9194,N_8482,N_8139);
nor U9195 (N_9195,N_8033,N_7802);
nor U9196 (N_9196,N_7986,N_7846);
or U9197 (N_9197,N_7710,N_8303);
or U9198 (N_9198,N_7993,N_8682);
and U9199 (N_9199,N_7727,N_8296);
nor U9200 (N_9200,N_8079,N_8363);
nand U9201 (N_9201,N_8581,N_8097);
nor U9202 (N_9202,N_8056,N_8407);
xnor U9203 (N_9203,N_7631,N_8662);
or U9204 (N_9204,N_8618,N_8189);
or U9205 (N_9205,N_7732,N_7887);
nor U9206 (N_9206,N_8532,N_8064);
and U9207 (N_9207,N_8109,N_7757);
nor U9208 (N_9208,N_8305,N_8461);
xor U9209 (N_9209,N_8388,N_7812);
nand U9210 (N_9210,N_8626,N_8691);
nand U9211 (N_9211,N_7632,N_8391);
xnor U9212 (N_9212,N_8210,N_8369);
xor U9213 (N_9213,N_7738,N_7604);
or U9214 (N_9214,N_7675,N_8274);
nand U9215 (N_9215,N_8444,N_7782);
or U9216 (N_9216,N_7968,N_7591);
or U9217 (N_9217,N_8209,N_8162);
and U9218 (N_9218,N_8007,N_7726);
xnor U9219 (N_9219,N_8479,N_7715);
nand U9220 (N_9220,N_8550,N_8458);
or U9221 (N_9221,N_8734,N_8071);
nand U9222 (N_9222,N_8360,N_8246);
or U9223 (N_9223,N_7754,N_8220);
nand U9224 (N_9224,N_8498,N_7530);
nor U9225 (N_9225,N_8582,N_8073);
xor U9226 (N_9226,N_8668,N_7706);
or U9227 (N_9227,N_8658,N_8422);
or U9228 (N_9228,N_8432,N_7728);
or U9229 (N_9229,N_7681,N_7609);
nand U9230 (N_9230,N_8635,N_7560);
or U9231 (N_9231,N_7598,N_8571);
and U9232 (N_9232,N_7576,N_8371);
or U9233 (N_9233,N_7635,N_8488);
and U9234 (N_9234,N_8382,N_8456);
nor U9235 (N_9235,N_8297,N_8312);
xnor U9236 (N_9236,N_8431,N_8085);
or U9237 (N_9237,N_8119,N_8116);
xnor U9238 (N_9238,N_7799,N_7554);
nor U9239 (N_9239,N_8221,N_8183);
and U9240 (N_9240,N_8125,N_8746);
nor U9241 (N_9241,N_7551,N_8702);
or U9242 (N_9242,N_8300,N_8506);
and U9243 (N_9243,N_8663,N_7511);
nor U9244 (N_9244,N_8575,N_7807);
and U9245 (N_9245,N_8339,N_7621);
xor U9246 (N_9246,N_8072,N_8528);
nand U9247 (N_9247,N_8559,N_8361);
nor U9248 (N_9248,N_8415,N_8723);
xor U9249 (N_9249,N_7643,N_7634);
nor U9250 (N_9250,N_8285,N_7788);
nor U9251 (N_9251,N_7518,N_8137);
or U9252 (N_9252,N_8098,N_8347);
nand U9253 (N_9253,N_8655,N_8406);
nor U9254 (N_9254,N_8069,N_8463);
xnor U9255 (N_9255,N_7944,N_8014);
and U9256 (N_9256,N_8323,N_7556);
nand U9257 (N_9257,N_8335,N_8043);
nand U9258 (N_9258,N_8747,N_8411);
nor U9259 (N_9259,N_8462,N_8511);
and U9260 (N_9260,N_7680,N_7555);
nor U9261 (N_9261,N_8254,N_8309);
xor U9262 (N_9262,N_8450,N_7905);
nand U9263 (N_9263,N_7832,N_8042);
nand U9264 (N_9264,N_7806,N_7644);
nand U9265 (N_9265,N_7917,N_8383);
or U9266 (N_9266,N_8449,N_8055);
and U9267 (N_9267,N_7927,N_7893);
and U9268 (N_9268,N_7614,N_7843);
nand U9269 (N_9269,N_8572,N_8029);
or U9270 (N_9270,N_7849,N_8531);
nand U9271 (N_9271,N_8494,N_8336);
and U9272 (N_9272,N_8424,N_7602);
and U9273 (N_9273,N_7946,N_7912);
and U9274 (N_9274,N_7844,N_7626);
and U9275 (N_9275,N_7540,N_8426);
nor U9276 (N_9276,N_7837,N_7720);
and U9277 (N_9277,N_8175,N_8594);
or U9278 (N_9278,N_7977,N_8539);
xnor U9279 (N_9279,N_8198,N_8429);
xnor U9280 (N_9280,N_8191,N_8364);
nand U9281 (N_9281,N_7840,N_8045);
xor U9282 (N_9282,N_8061,N_7705);
nand U9283 (N_9283,N_7909,N_8025);
and U9284 (N_9284,N_8437,N_7895);
and U9285 (N_9285,N_8076,N_8398);
xor U9286 (N_9286,N_8243,N_7652);
nor U9287 (N_9287,N_7859,N_7666);
nand U9288 (N_9288,N_8464,N_7535);
and U9289 (N_9289,N_8345,N_8512);
nor U9290 (N_9290,N_8420,N_8196);
nor U9291 (N_9291,N_8349,N_8555);
or U9292 (N_9292,N_8615,N_8225);
xnor U9293 (N_9293,N_7791,N_8716);
nand U9294 (N_9294,N_7760,N_8224);
nand U9295 (N_9295,N_8465,N_8262);
xnor U9296 (N_9296,N_8358,N_7636);
xnor U9297 (N_9297,N_8153,N_8044);
and U9298 (N_9298,N_8219,N_7971);
or U9299 (N_9299,N_8270,N_8695);
nand U9300 (N_9300,N_8012,N_8705);
and U9301 (N_9301,N_7820,N_8743);
or U9302 (N_9302,N_8156,N_7861);
and U9303 (N_9303,N_8216,N_8318);
nor U9304 (N_9304,N_8741,N_7770);
and U9305 (N_9305,N_8697,N_7990);
xnor U9306 (N_9306,N_7691,N_7762);
nor U9307 (N_9307,N_8683,N_7716);
and U9308 (N_9308,N_8538,N_8271);
or U9309 (N_9309,N_7872,N_8616);
and U9310 (N_9310,N_8177,N_7919);
nor U9311 (N_9311,N_8089,N_8469);
nor U9312 (N_9312,N_8222,N_8290);
or U9313 (N_9313,N_8298,N_7970);
nor U9314 (N_9314,N_8015,N_7935);
nand U9315 (N_9315,N_8308,N_7640);
nand U9316 (N_9316,N_7904,N_8036);
or U9317 (N_9317,N_8402,N_7851);
and U9318 (N_9318,N_8112,N_8701);
and U9319 (N_9319,N_7737,N_7587);
xnor U9320 (N_9320,N_8127,N_7648);
nand U9321 (N_9321,N_7755,N_7593);
nand U9322 (N_9322,N_7615,N_8302);
nor U9323 (N_9323,N_7818,N_7505);
xor U9324 (N_9324,N_7902,N_8373);
nor U9325 (N_9325,N_8567,N_8102);
nor U9326 (N_9326,N_7868,N_7834);
nand U9327 (N_9327,N_7764,N_8604);
nor U9328 (N_9328,N_7506,N_7922);
nand U9329 (N_9329,N_8050,N_8205);
nor U9330 (N_9330,N_7536,N_7739);
nand U9331 (N_9331,N_7792,N_8502);
nand U9332 (N_9332,N_7873,N_7985);
or U9333 (N_9333,N_7845,N_7607);
xnor U9334 (N_9334,N_8232,N_8573);
or U9335 (N_9335,N_8054,N_8158);
nand U9336 (N_9336,N_8732,N_7725);
or U9337 (N_9337,N_8557,N_7906);
nor U9338 (N_9338,N_8367,N_8251);
and U9339 (N_9339,N_7890,N_8643);
or U9340 (N_9340,N_7750,N_8154);
nor U9341 (N_9341,N_8039,N_8062);
nand U9342 (N_9342,N_8438,N_8118);
or U9343 (N_9343,N_7996,N_7616);
or U9344 (N_9344,N_8529,N_7785);
nor U9345 (N_9345,N_8556,N_8441);
nand U9346 (N_9346,N_8047,N_8218);
nand U9347 (N_9347,N_7823,N_7713);
nand U9348 (N_9348,N_7930,N_8326);
nand U9349 (N_9349,N_7722,N_7724);
nor U9350 (N_9350,N_7514,N_7988);
xor U9351 (N_9351,N_7938,N_8425);
nand U9352 (N_9352,N_7896,N_7589);
nand U9353 (N_9353,N_8350,N_8051);
or U9354 (N_9354,N_7570,N_8035);
xor U9355 (N_9355,N_7959,N_8453);
or U9356 (N_9356,N_8527,N_7931);
or U9357 (N_9357,N_8379,N_8330);
or U9358 (N_9358,N_8276,N_7618);
nand U9359 (N_9359,N_8002,N_8245);
xnor U9360 (N_9360,N_8729,N_7746);
and U9361 (N_9361,N_7721,N_7794);
xor U9362 (N_9362,N_8570,N_7533);
xnor U9363 (N_9363,N_8740,N_8485);
nand U9364 (N_9364,N_8473,N_8698);
nor U9365 (N_9365,N_8355,N_8075);
nor U9366 (N_9366,N_8332,N_7714);
nor U9367 (N_9367,N_8128,N_7894);
xnor U9368 (N_9368,N_8344,N_7747);
or U9369 (N_9369,N_8174,N_7695);
nor U9370 (N_9370,N_8580,N_7685);
and U9371 (N_9371,N_7960,N_7848);
nor U9372 (N_9372,N_8630,N_8609);
nand U9373 (N_9373,N_8710,N_7658);
nor U9374 (N_9374,N_8657,N_7657);
xnor U9375 (N_9375,N_8246,N_8172);
and U9376 (N_9376,N_8469,N_7543);
and U9377 (N_9377,N_8084,N_8380);
nor U9378 (N_9378,N_8708,N_7866);
and U9379 (N_9379,N_7657,N_7747);
or U9380 (N_9380,N_7610,N_8162);
and U9381 (N_9381,N_7939,N_8338);
or U9382 (N_9382,N_8278,N_7649);
or U9383 (N_9383,N_7789,N_8172);
and U9384 (N_9384,N_7915,N_8507);
nor U9385 (N_9385,N_7614,N_7949);
nand U9386 (N_9386,N_8119,N_7666);
or U9387 (N_9387,N_8413,N_7524);
xnor U9388 (N_9388,N_8172,N_8705);
xnor U9389 (N_9389,N_8638,N_7590);
nor U9390 (N_9390,N_8189,N_8140);
and U9391 (N_9391,N_8309,N_8011);
or U9392 (N_9392,N_8101,N_8371);
or U9393 (N_9393,N_7934,N_7859);
nor U9394 (N_9394,N_7522,N_8038);
xor U9395 (N_9395,N_7967,N_7975);
or U9396 (N_9396,N_7881,N_8703);
and U9397 (N_9397,N_8187,N_8461);
or U9398 (N_9398,N_7725,N_7767);
and U9399 (N_9399,N_8673,N_7709);
and U9400 (N_9400,N_8399,N_7683);
xnor U9401 (N_9401,N_8558,N_8143);
and U9402 (N_9402,N_8383,N_8342);
nor U9403 (N_9403,N_7897,N_7938);
and U9404 (N_9404,N_7588,N_8280);
nor U9405 (N_9405,N_8054,N_7774);
and U9406 (N_9406,N_8502,N_8609);
nor U9407 (N_9407,N_8694,N_7517);
xnor U9408 (N_9408,N_7624,N_8517);
nand U9409 (N_9409,N_7670,N_7882);
xnor U9410 (N_9410,N_8593,N_7558);
nor U9411 (N_9411,N_7746,N_8717);
or U9412 (N_9412,N_8468,N_8749);
xor U9413 (N_9413,N_7968,N_8408);
nand U9414 (N_9414,N_7774,N_7502);
or U9415 (N_9415,N_8395,N_8263);
nand U9416 (N_9416,N_7725,N_7613);
nor U9417 (N_9417,N_7975,N_8748);
and U9418 (N_9418,N_8423,N_8661);
nor U9419 (N_9419,N_8346,N_8575);
or U9420 (N_9420,N_8288,N_8615);
xnor U9421 (N_9421,N_7743,N_8719);
and U9422 (N_9422,N_8302,N_7638);
and U9423 (N_9423,N_7725,N_8502);
and U9424 (N_9424,N_8304,N_7638);
and U9425 (N_9425,N_8701,N_7565);
nor U9426 (N_9426,N_8375,N_8056);
nand U9427 (N_9427,N_8301,N_8128);
xnor U9428 (N_9428,N_8659,N_7548);
nor U9429 (N_9429,N_7799,N_8420);
xor U9430 (N_9430,N_8558,N_8553);
or U9431 (N_9431,N_7535,N_7622);
xnor U9432 (N_9432,N_8219,N_7642);
and U9433 (N_9433,N_7828,N_7838);
or U9434 (N_9434,N_8370,N_8649);
xnor U9435 (N_9435,N_7656,N_8503);
xor U9436 (N_9436,N_8564,N_8152);
nor U9437 (N_9437,N_7698,N_8091);
nand U9438 (N_9438,N_8685,N_7698);
and U9439 (N_9439,N_8624,N_8682);
nand U9440 (N_9440,N_8177,N_7544);
nor U9441 (N_9441,N_8083,N_7665);
xor U9442 (N_9442,N_7952,N_8085);
and U9443 (N_9443,N_8540,N_7952);
or U9444 (N_9444,N_8431,N_7615);
nand U9445 (N_9445,N_7665,N_8132);
or U9446 (N_9446,N_7736,N_8389);
or U9447 (N_9447,N_7522,N_8664);
or U9448 (N_9448,N_8471,N_7858);
xor U9449 (N_9449,N_7928,N_7839);
or U9450 (N_9450,N_8505,N_7971);
and U9451 (N_9451,N_7791,N_7549);
nand U9452 (N_9452,N_7996,N_7986);
nor U9453 (N_9453,N_8125,N_8132);
nor U9454 (N_9454,N_7887,N_8417);
and U9455 (N_9455,N_8125,N_7909);
nand U9456 (N_9456,N_8040,N_8551);
xnor U9457 (N_9457,N_7901,N_8322);
or U9458 (N_9458,N_8304,N_8070);
and U9459 (N_9459,N_7868,N_7968);
and U9460 (N_9460,N_8601,N_8311);
xor U9461 (N_9461,N_8620,N_7561);
nand U9462 (N_9462,N_7526,N_8175);
nor U9463 (N_9463,N_7805,N_8615);
nand U9464 (N_9464,N_8564,N_7656);
or U9465 (N_9465,N_8493,N_8572);
nand U9466 (N_9466,N_7615,N_8419);
nand U9467 (N_9467,N_8409,N_8645);
or U9468 (N_9468,N_8128,N_8690);
xor U9469 (N_9469,N_8083,N_8677);
xnor U9470 (N_9470,N_8428,N_8465);
and U9471 (N_9471,N_8609,N_7902);
nand U9472 (N_9472,N_8069,N_7795);
and U9473 (N_9473,N_8556,N_7629);
nor U9474 (N_9474,N_7976,N_7730);
and U9475 (N_9475,N_7692,N_8172);
and U9476 (N_9476,N_8214,N_8285);
or U9477 (N_9477,N_7824,N_7594);
or U9478 (N_9478,N_8219,N_7531);
or U9479 (N_9479,N_8383,N_8530);
nand U9480 (N_9480,N_7706,N_7593);
nand U9481 (N_9481,N_7618,N_8009);
and U9482 (N_9482,N_7761,N_7645);
nor U9483 (N_9483,N_8159,N_7758);
nand U9484 (N_9484,N_8605,N_7829);
xnor U9485 (N_9485,N_7677,N_8353);
and U9486 (N_9486,N_8217,N_7884);
or U9487 (N_9487,N_8615,N_8081);
nand U9488 (N_9488,N_8133,N_7832);
nor U9489 (N_9489,N_8436,N_8271);
and U9490 (N_9490,N_8275,N_8748);
nand U9491 (N_9491,N_8025,N_8077);
or U9492 (N_9492,N_8021,N_7942);
xor U9493 (N_9493,N_8223,N_7989);
xor U9494 (N_9494,N_8063,N_8164);
nor U9495 (N_9495,N_8567,N_8361);
or U9496 (N_9496,N_7579,N_8021);
nand U9497 (N_9497,N_7871,N_7897);
xor U9498 (N_9498,N_8059,N_7798);
nand U9499 (N_9499,N_8595,N_7934);
nand U9500 (N_9500,N_8041,N_7722);
and U9501 (N_9501,N_8426,N_7933);
xnor U9502 (N_9502,N_7839,N_7925);
nor U9503 (N_9503,N_8203,N_7619);
xor U9504 (N_9504,N_7973,N_8119);
or U9505 (N_9505,N_8456,N_8153);
xnor U9506 (N_9506,N_8347,N_8017);
nand U9507 (N_9507,N_7981,N_7847);
and U9508 (N_9508,N_7960,N_8513);
nand U9509 (N_9509,N_7795,N_7608);
xnor U9510 (N_9510,N_8169,N_8435);
xor U9511 (N_9511,N_8582,N_8141);
nand U9512 (N_9512,N_8375,N_7553);
nand U9513 (N_9513,N_7505,N_8195);
or U9514 (N_9514,N_8724,N_7717);
nor U9515 (N_9515,N_8382,N_8086);
or U9516 (N_9516,N_8467,N_8384);
or U9517 (N_9517,N_7955,N_8264);
nand U9518 (N_9518,N_8458,N_8484);
nand U9519 (N_9519,N_8373,N_8709);
xnor U9520 (N_9520,N_7673,N_7519);
nor U9521 (N_9521,N_8150,N_8126);
and U9522 (N_9522,N_8747,N_7748);
nor U9523 (N_9523,N_8493,N_8071);
or U9524 (N_9524,N_8738,N_8558);
and U9525 (N_9525,N_7929,N_8650);
nor U9526 (N_9526,N_8285,N_7515);
nor U9527 (N_9527,N_7657,N_8004);
xnor U9528 (N_9528,N_7748,N_8144);
xnor U9529 (N_9529,N_7831,N_8224);
or U9530 (N_9530,N_8477,N_8058);
or U9531 (N_9531,N_8056,N_8333);
xnor U9532 (N_9532,N_8679,N_8555);
or U9533 (N_9533,N_8224,N_7512);
xnor U9534 (N_9534,N_7507,N_7651);
nand U9535 (N_9535,N_8332,N_8397);
or U9536 (N_9536,N_8309,N_7711);
nand U9537 (N_9537,N_8082,N_7805);
or U9538 (N_9538,N_7656,N_8640);
nor U9539 (N_9539,N_7510,N_8461);
xnor U9540 (N_9540,N_7584,N_8735);
nor U9541 (N_9541,N_8745,N_7959);
and U9542 (N_9542,N_7758,N_8335);
or U9543 (N_9543,N_8015,N_7763);
nor U9544 (N_9544,N_7935,N_7538);
and U9545 (N_9545,N_7646,N_7901);
nor U9546 (N_9546,N_8039,N_8285);
or U9547 (N_9547,N_7546,N_7949);
xor U9548 (N_9548,N_7903,N_8534);
or U9549 (N_9549,N_7743,N_7686);
xnor U9550 (N_9550,N_8464,N_8202);
nor U9551 (N_9551,N_7751,N_8594);
xor U9552 (N_9552,N_8050,N_8207);
xnor U9553 (N_9553,N_7892,N_8150);
nor U9554 (N_9554,N_8442,N_8655);
nor U9555 (N_9555,N_7771,N_7863);
and U9556 (N_9556,N_8031,N_8192);
nand U9557 (N_9557,N_8109,N_8062);
nor U9558 (N_9558,N_8689,N_8742);
and U9559 (N_9559,N_7693,N_7975);
xor U9560 (N_9560,N_8412,N_7833);
nand U9561 (N_9561,N_7900,N_7918);
nand U9562 (N_9562,N_7689,N_8304);
and U9563 (N_9563,N_8377,N_7750);
xor U9564 (N_9564,N_7633,N_8312);
nor U9565 (N_9565,N_8035,N_8400);
and U9566 (N_9566,N_8254,N_8303);
nor U9567 (N_9567,N_8266,N_7869);
xnor U9568 (N_9568,N_8589,N_8338);
nor U9569 (N_9569,N_8241,N_8229);
or U9570 (N_9570,N_7839,N_8042);
and U9571 (N_9571,N_7632,N_8128);
nor U9572 (N_9572,N_8158,N_8431);
nor U9573 (N_9573,N_7650,N_8331);
nor U9574 (N_9574,N_8711,N_8216);
xor U9575 (N_9575,N_7704,N_7849);
nor U9576 (N_9576,N_8381,N_7668);
or U9577 (N_9577,N_8225,N_8115);
and U9578 (N_9578,N_8156,N_7621);
xor U9579 (N_9579,N_8547,N_8344);
nand U9580 (N_9580,N_7878,N_8433);
nand U9581 (N_9581,N_7864,N_7613);
xor U9582 (N_9582,N_8531,N_7813);
and U9583 (N_9583,N_8660,N_8738);
or U9584 (N_9584,N_8586,N_8125);
nand U9585 (N_9585,N_7583,N_8294);
nor U9586 (N_9586,N_7675,N_8713);
or U9587 (N_9587,N_7729,N_7925);
or U9588 (N_9588,N_8657,N_8656);
or U9589 (N_9589,N_7766,N_7883);
xnor U9590 (N_9590,N_7909,N_7713);
or U9591 (N_9591,N_8006,N_7905);
nor U9592 (N_9592,N_7728,N_8235);
nand U9593 (N_9593,N_8196,N_7726);
nand U9594 (N_9594,N_8254,N_8311);
or U9595 (N_9595,N_8716,N_7845);
xor U9596 (N_9596,N_7628,N_7972);
nand U9597 (N_9597,N_8560,N_7843);
nor U9598 (N_9598,N_8240,N_8350);
or U9599 (N_9599,N_7867,N_8208);
xor U9600 (N_9600,N_8203,N_7871);
xnor U9601 (N_9601,N_8689,N_7837);
or U9602 (N_9602,N_8200,N_7720);
nor U9603 (N_9603,N_8746,N_7605);
xnor U9604 (N_9604,N_8022,N_7715);
xnor U9605 (N_9605,N_7687,N_7971);
xor U9606 (N_9606,N_8469,N_8223);
xor U9607 (N_9607,N_8050,N_8024);
xnor U9608 (N_9608,N_8573,N_7509);
xor U9609 (N_9609,N_8111,N_8222);
nor U9610 (N_9610,N_7520,N_8625);
nor U9611 (N_9611,N_8529,N_7681);
nor U9612 (N_9612,N_8088,N_7557);
nor U9613 (N_9613,N_8479,N_8399);
nand U9614 (N_9614,N_8647,N_8145);
or U9615 (N_9615,N_8225,N_7514);
nor U9616 (N_9616,N_8707,N_8526);
nand U9617 (N_9617,N_7750,N_7715);
nand U9618 (N_9618,N_8052,N_7802);
nand U9619 (N_9619,N_8685,N_7661);
xor U9620 (N_9620,N_8276,N_7860);
nand U9621 (N_9621,N_7943,N_8556);
and U9622 (N_9622,N_8696,N_7970);
or U9623 (N_9623,N_7609,N_8337);
nand U9624 (N_9624,N_8726,N_7570);
or U9625 (N_9625,N_8410,N_8492);
xor U9626 (N_9626,N_7996,N_8608);
xnor U9627 (N_9627,N_8579,N_8097);
xnor U9628 (N_9628,N_7802,N_8612);
nor U9629 (N_9629,N_8054,N_7869);
or U9630 (N_9630,N_8239,N_8074);
xnor U9631 (N_9631,N_7899,N_8307);
and U9632 (N_9632,N_7572,N_7552);
nor U9633 (N_9633,N_8076,N_7545);
nor U9634 (N_9634,N_8731,N_7686);
or U9635 (N_9635,N_7813,N_7996);
nor U9636 (N_9636,N_7507,N_7872);
xor U9637 (N_9637,N_7624,N_7669);
or U9638 (N_9638,N_8051,N_7899);
xor U9639 (N_9639,N_8110,N_7900);
nand U9640 (N_9640,N_7938,N_7516);
or U9641 (N_9641,N_7839,N_7723);
nand U9642 (N_9642,N_8348,N_7957);
xnor U9643 (N_9643,N_8316,N_8310);
nor U9644 (N_9644,N_8057,N_7956);
and U9645 (N_9645,N_7685,N_8495);
and U9646 (N_9646,N_8639,N_7535);
nand U9647 (N_9647,N_8495,N_7846);
nor U9648 (N_9648,N_8415,N_7854);
nor U9649 (N_9649,N_8272,N_7545);
and U9650 (N_9650,N_8494,N_8419);
nor U9651 (N_9651,N_8299,N_8619);
or U9652 (N_9652,N_8638,N_8581);
nand U9653 (N_9653,N_8505,N_7646);
or U9654 (N_9654,N_7756,N_8297);
xor U9655 (N_9655,N_8558,N_8071);
nand U9656 (N_9656,N_7716,N_8275);
and U9657 (N_9657,N_8120,N_7732);
and U9658 (N_9658,N_8538,N_8190);
xor U9659 (N_9659,N_8299,N_8705);
nand U9660 (N_9660,N_7894,N_8183);
nor U9661 (N_9661,N_8090,N_8020);
or U9662 (N_9662,N_7672,N_8740);
nand U9663 (N_9663,N_7926,N_8503);
nand U9664 (N_9664,N_7604,N_7984);
or U9665 (N_9665,N_7926,N_7997);
and U9666 (N_9666,N_7637,N_7891);
xnor U9667 (N_9667,N_7992,N_8336);
and U9668 (N_9668,N_8523,N_8671);
or U9669 (N_9669,N_8062,N_8627);
nor U9670 (N_9670,N_8244,N_8097);
and U9671 (N_9671,N_7682,N_7544);
or U9672 (N_9672,N_7531,N_8040);
nor U9673 (N_9673,N_7962,N_8251);
nor U9674 (N_9674,N_7824,N_7721);
or U9675 (N_9675,N_8295,N_8358);
or U9676 (N_9676,N_7511,N_8180);
nand U9677 (N_9677,N_8395,N_7906);
or U9678 (N_9678,N_8076,N_8690);
and U9679 (N_9679,N_7949,N_8501);
nor U9680 (N_9680,N_8162,N_8537);
nor U9681 (N_9681,N_8325,N_8014);
or U9682 (N_9682,N_8040,N_7890);
or U9683 (N_9683,N_8234,N_8690);
or U9684 (N_9684,N_8228,N_8441);
or U9685 (N_9685,N_7521,N_8694);
and U9686 (N_9686,N_7666,N_8442);
and U9687 (N_9687,N_8606,N_7856);
and U9688 (N_9688,N_7674,N_8624);
or U9689 (N_9689,N_7751,N_8567);
nor U9690 (N_9690,N_7935,N_8225);
or U9691 (N_9691,N_8511,N_8206);
nor U9692 (N_9692,N_8560,N_7634);
or U9693 (N_9693,N_8349,N_8506);
nor U9694 (N_9694,N_8541,N_8335);
nor U9695 (N_9695,N_8262,N_7606);
nor U9696 (N_9696,N_8414,N_7954);
xor U9697 (N_9697,N_8136,N_8497);
nor U9698 (N_9698,N_7884,N_7745);
and U9699 (N_9699,N_8638,N_7692);
xnor U9700 (N_9700,N_8131,N_7848);
or U9701 (N_9701,N_8180,N_7875);
and U9702 (N_9702,N_8630,N_7824);
nand U9703 (N_9703,N_8271,N_8474);
xor U9704 (N_9704,N_7502,N_8369);
nor U9705 (N_9705,N_7687,N_8312);
xnor U9706 (N_9706,N_8236,N_8339);
nor U9707 (N_9707,N_7695,N_7933);
and U9708 (N_9708,N_8174,N_8271);
and U9709 (N_9709,N_7938,N_7553);
nor U9710 (N_9710,N_7789,N_8204);
and U9711 (N_9711,N_7664,N_7734);
or U9712 (N_9712,N_8285,N_7621);
nand U9713 (N_9713,N_8330,N_8416);
nor U9714 (N_9714,N_8152,N_8647);
nor U9715 (N_9715,N_8437,N_8565);
nor U9716 (N_9716,N_8658,N_8194);
and U9717 (N_9717,N_8176,N_8580);
nand U9718 (N_9718,N_7812,N_8451);
xor U9719 (N_9719,N_8727,N_8192);
nand U9720 (N_9720,N_8152,N_7636);
and U9721 (N_9721,N_8718,N_7898);
nor U9722 (N_9722,N_7836,N_8561);
xnor U9723 (N_9723,N_7925,N_7667);
xnor U9724 (N_9724,N_8137,N_8181);
and U9725 (N_9725,N_8680,N_7878);
and U9726 (N_9726,N_8612,N_7501);
and U9727 (N_9727,N_7999,N_8315);
nand U9728 (N_9728,N_7548,N_7814);
xor U9729 (N_9729,N_8288,N_7992);
nand U9730 (N_9730,N_8640,N_8558);
xnor U9731 (N_9731,N_7664,N_7865);
xor U9732 (N_9732,N_8705,N_8102);
xnor U9733 (N_9733,N_7776,N_8502);
and U9734 (N_9734,N_8402,N_8585);
nand U9735 (N_9735,N_8030,N_8721);
xor U9736 (N_9736,N_8700,N_8728);
or U9737 (N_9737,N_8367,N_8695);
or U9738 (N_9738,N_7997,N_7888);
nand U9739 (N_9739,N_8116,N_8205);
or U9740 (N_9740,N_8688,N_7877);
nand U9741 (N_9741,N_8172,N_8416);
or U9742 (N_9742,N_8632,N_7678);
or U9743 (N_9743,N_7526,N_7730);
nor U9744 (N_9744,N_7635,N_7539);
xnor U9745 (N_9745,N_8300,N_8711);
xor U9746 (N_9746,N_7602,N_8168);
or U9747 (N_9747,N_7883,N_7838);
or U9748 (N_9748,N_8028,N_8146);
xor U9749 (N_9749,N_7869,N_8220);
nor U9750 (N_9750,N_7501,N_7609);
xor U9751 (N_9751,N_7636,N_8627);
and U9752 (N_9752,N_7571,N_7712);
xnor U9753 (N_9753,N_8648,N_7924);
nor U9754 (N_9754,N_8523,N_8748);
and U9755 (N_9755,N_8332,N_7511);
or U9756 (N_9756,N_7631,N_8156);
xnor U9757 (N_9757,N_7518,N_7677);
and U9758 (N_9758,N_8453,N_8080);
or U9759 (N_9759,N_8474,N_8735);
nor U9760 (N_9760,N_7996,N_7550);
and U9761 (N_9761,N_8394,N_7961);
nand U9762 (N_9762,N_8333,N_8683);
nand U9763 (N_9763,N_7796,N_7685);
nor U9764 (N_9764,N_8093,N_8623);
nand U9765 (N_9765,N_8024,N_8186);
nand U9766 (N_9766,N_7694,N_7728);
nand U9767 (N_9767,N_7972,N_7606);
nor U9768 (N_9768,N_8547,N_7522);
or U9769 (N_9769,N_8066,N_8165);
and U9770 (N_9770,N_7805,N_7855);
and U9771 (N_9771,N_7672,N_8277);
xor U9772 (N_9772,N_8282,N_8518);
xor U9773 (N_9773,N_7951,N_7745);
or U9774 (N_9774,N_7622,N_8067);
or U9775 (N_9775,N_7625,N_8129);
and U9776 (N_9776,N_8587,N_7840);
nand U9777 (N_9777,N_7930,N_8366);
and U9778 (N_9778,N_8456,N_8408);
nand U9779 (N_9779,N_7780,N_8649);
nand U9780 (N_9780,N_8518,N_7981);
and U9781 (N_9781,N_7680,N_8147);
nand U9782 (N_9782,N_8492,N_7728);
nand U9783 (N_9783,N_7785,N_8070);
or U9784 (N_9784,N_8129,N_8185);
and U9785 (N_9785,N_7899,N_8608);
nand U9786 (N_9786,N_8278,N_8142);
nand U9787 (N_9787,N_8262,N_8491);
nor U9788 (N_9788,N_8573,N_7911);
xnor U9789 (N_9789,N_7944,N_7541);
xor U9790 (N_9790,N_8354,N_8641);
or U9791 (N_9791,N_7819,N_7550);
nand U9792 (N_9792,N_8198,N_8077);
or U9793 (N_9793,N_7998,N_8544);
or U9794 (N_9794,N_7647,N_7805);
or U9795 (N_9795,N_7622,N_8314);
and U9796 (N_9796,N_7740,N_7591);
or U9797 (N_9797,N_7525,N_8396);
or U9798 (N_9798,N_7993,N_8585);
or U9799 (N_9799,N_8294,N_8003);
xor U9800 (N_9800,N_8391,N_7532);
nor U9801 (N_9801,N_8363,N_7651);
nand U9802 (N_9802,N_8150,N_8717);
or U9803 (N_9803,N_8167,N_8411);
or U9804 (N_9804,N_7785,N_8270);
or U9805 (N_9805,N_8417,N_8102);
and U9806 (N_9806,N_7722,N_7931);
nand U9807 (N_9807,N_7873,N_7710);
or U9808 (N_9808,N_8405,N_8048);
nor U9809 (N_9809,N_8636,N_8095);
xnor U9810 (N_9810,N_8504,N_7787);
nand U9811 (N_9811,N_8438,N_8244);
xor U9812 (N_9812,N_7731,N_8129);
xor U9813 (N_9813,N_8261,N_8503);
xor U9814 (N_9814,N_7667,N_8543);
xnor U9815 (N_9815,N_7972,N_7863);
and U9816 (N_9816,N_8424,N_7660);
and U9817 (N_9817,N_8174,N_8594);
or U9818 (N_9818,N_7523,N_7997);
and U9819 (N_9819,N_8396,N_8243);
nor U9820 (N_9820,N_8414,N_7691);
nand U9821 (N_9821,N_8181,N_7817);
xnor U9822 (N_9822,N_8280,N_8321);
xor U9823 (N_9823,N_8140,N_7900);
nor U9824 (N_9824,N_7993,N_7661);
nor U9825 (N_9825,N_7567,N_7765);
nand U9826 (N_9826,N_8747,N_8569);
xor U9827 (N_9827,N_7845,N_7624);
xnor U9828 (N_9828,N_7776,N_7923);
and U9829 (N_9829,N_7532,N_7626);
xor U9830 (N_9830,N_7949,N_8631);
and U9831 (N_9831,N_8738,N_8543);
or U9832 (N_9832,N_8335,N_8645);
or U9833 (N_9833,N_7965,N_8131);
nor U9834 (N_9834,N_7619,N_7707);
xnor U9835 (N_9835,N_8048,N_7558);
and U9836 (N_9836,N_8644,N_8390);
nor U9837 (N_9837,N_8168,N_8136);
or U9838 (N_9838,N_8523,N_8490);
or U9839 (N_9839,N_8360,N_8068);
nor U9840 (N_9840,N_8251,N_8527);
xnor U9841 (N_9841,N_8655,N_7788);
and U9842 (N_9842,N_8628,N_8513);
nand U9843 (N_9843,N_8089,N_7573);
nand U9844 (N_9844,N_8493,N_8745);
and U9845 (N_9845,N_8687,N_8244);
nor U9846 (N_9846,N_8162,N_8643);
nor U9847 (N_9847,N_8047,N_8592);
nand U9848 (N_9848,N_7666,N_7832);
xor U9849 (N_9849,N_7611,N_8652);
nor U9850 (N_9850,N_8116,N_8167);
xnor U9851 (N_9851,N_8115,N_8427);
and U9852 (N_9852,N_8391,N_8271);
or U9853 (N_9853,N_8198,N_8011);
and U9854 (N_9854,N_8195,N_7866);
nor U9855 (N_9855,N_7782,N_8730);
xor U9856 (N_9856,N_8101,N_8108);
and U9857 (N_9857,N_8098,N_8405);
nand U9858 (N_9858,N_8566,N_7709);
xnor U9859 (N_9859,N_8644,N_8300);
nor U9860 (N_9860,N_8326,N_8088);
xor U9861 (N_9861,N_8077,N_8343);
or U9862 (N_9862,N_8457,N_8426);
and U9863 (N_9863,N_7755,N_8655);
and U9864 (N_9864,N_8304,N_7686);
nor U9865 (N_9865,N_8485,N_8402);
nor U9866 (N_9866,N_8134,N_8323);
and U9867 (N_9867,N_8545,N_8055);
nor U9868 (N_9868,N_8642,N_7634);
or U9869 (N_9869,N_8139,N_7635);
xnor U9870 (N_9870,N_8323,N_7985);
or U9871 (N_9871,N_8504,N_8666);
nor U9872 (N_9872,N_7560,N_8582);
and U9873 (N_9873,N_8363,N_7593);
nor U9874 (N_9874,N_7733,N_8467);
nor U9875 (N_9875,N_8654,N_8111);
nor U9876 (N_9876,N_8419,N_7959);
and U9877 (N_9877,N_8023,N_8349);
and U9878 (N_9878,N_7934,N_7834);
nand U9879 (N_9879,N_8481,N_7644);
xnor U9880 (N_9880,N_7538,N_7671);
and U9881 (N_9881,N_7949,N_7623);
or U9882 (N_9882,N_8432,N_8189);
nor U9883 (N_9883,N_8525,N_8240);
nor U9884 (N_9884,N_7750,N_7605);
xnor U9885 (N_9885,N_7767,N_8584);
nand U9886 (N_9886,N_7596,N_7864);
nand U9887 (N_9887,N_7764,N_7904);
and U9888 (N_9888,N_8392,N_7847);
and U9889 (N_9889,N_8649,N_7869);
xor U9890 (N_9890,N_7629,N_8093);
xnor U9891 (N_9891,N_8163,N_7728);
xnor U9892 (N_9892,N_8247,N_8235);
xnor U9893 (N_9893,N_8125,N_8145);
and U9894 (N_9894,N_8428,N_7758);
nand U9895 (N_9895,N_8382,N_7632);
and U9896 (N_9896,N_7873,N_8014);
nand U9897 (N_9897,N_7636,N_7597);
or U9898 (N_9898,N_7593,N_8427);
nor U9899 (N_9899,N_8160,N_8710);
or U9900 (N_9900,N_7831,N_8032);
nand U9901 (N_9901,N_8531,N_7560);
nor U9902 (N_9902,N_8172,N_7951);
xnor U9903 (N_9903,N_8363,N_8464);
nand U9904 (N_9904,N_8313,N_7805);
xor U9905 (N_9905,N_8485,N_8541);
nor U9906 (N_9906,N_8616,N_7578);
xnor U9907 (N_9907,N_8178,N_8129);
xor U9908 (N_9908,N_7746,N_7599);
or U9909 (N_9909,N_7524,N_8077);
xor U9910 (N_9910,N_8563,N_8159);
nor U9911 (N_9911,N_7947,N_7838);
or U9912 (N_9912,N_7832,N_7775);
or U9913 (N_9913,N_8417,N_7793);
nand U9914 (N_9914,N_8285,N_8646);
and U9915 (N_9915,N_8629,N_8519);
and U9916 (N_9916,N_8554,N_7582);
nand U9917 (N_9917,N_8056,N_8530);
nand U9918 (N_9918,N_7963,N_8529);
or U9919 (N_9919,N_7587,N_7660);
and U9920 (N_9920,N_8007,N_7666);
nor U9921 (N_9921,N_8611,N_7955);
xor U9922 (N_9922,N_8211,N_8735);
and U9923 (N_9923,N_8020,N_8697);
xnor U9924 (N_9924,N_8452,N_7991);
and U9925 (N_9925,N_7695,N_7651);
and U9926 (N_9926,N_8603,N_8098);
nand U9927 (N_9927,N_7886,N_7667);
or U9928 (N_9928,N_8086,N_7692);
and U9929 (N_9929,N_7769,N_7608);
or U9930 (N_9930,N_8701,N_8391);
and U9931 (N_9931,N_7658,N_8080);
xnor U9932 (N_9932,N_7501,N_8603);
nand U9933 (N_9933,N_8469,N_8715);
or U9934 (N_9934,N_7916,N_8520);
or U9935 (N_9935,N_8195,N_7633);
nand U9936 (N_9936,N_7809,N_7620);
and U9937 (N_9937,N_7966,N_8326);
nor U9938 (N_9938,N_7717,N_8024);
and U9939 (N_9939,N_8075,N_8273);
and U9940 (N_9940,N_8504,N_8126);
nor U9941 (N_9941,N_7940,N_8232);
xnor U9942 (N_9942,N_8407,N_7878);
nand U9943 (N_9943,N_7726,N_8171);
nor U9944 (N_9944,N_8648,N_8745);
and U9945 (N_9945,N_7721,N_8088);
nand U9946 (N_9946,N_8120,N_7708);
xor U9947 (N_9947,N_7714,N_7672);
xnor U9948 (N_9948,N_8248,N_8631);
nand U9949 (N_9949,N_8542,N_8302);
or U9950 (N_9950,N_8603,N_8120);
and U9951 (N_9951,N_8142,N_7580);
xor U9952 (N_9952,N_8182,N_7562);
nand U9953 (N_9953,N_7507,N_7772);
or U9954 (N_9954,N_7781,N_8674);
nor U9955 (N_9955,N_8144,N_8244);
or U9956 (N_9956,N_8442,N_8583);
or U9957 (N_9957,N_7565,N_8175);
nor U9958 (N_9958,N_8502,N_7659);
and U9959 (N_9959,N_8745,N_7819);
xor U9960 (N_9960,N_8097,N_7508);
or U9961 (N_9961,N_7752,N_8219);
and U9962 (N_9962,N_7918,N_8087);
and U9963 (N_9963,N_8547,N_7881);
nand U9964 (N_9964,N_7560,N_8435);
or U9965 (N_9965,N_8645,N_7525);
and U9966 (N_9966,N_8308,N_8642);
nand U9967 (N_9967,N_7914,N_7736);
nor U9968 (N_9968,N_8639,N_8154);
nor U9969 (N_9969,N_7876,N_7609);
nor U9970 (N_9970,N_8322,N_7572);
or U9971 (N_9971,N_7816,N_7878);
nand U9972 (N_9972,N_8111,N_8627);
xnor U9973 (N_9973,N_8471,N_7706);
nor U9974 (N_9974,N_8733,N_8688);
nor U9975 (N_9975,N_7556,N_8074);
or U9976 (N_9976,N_7801,N_8452);
and U9977 (N_9977,N_7634,N_8281);
and U9978 (N_9978,N_8737,N_8076);
or U9979 (N_9979,N_8114,N_8234);
xor U9980 (N_9980,N_8574,N_8525);
nand U9981 (N_9981,N_8433,N_7938);
or U9982 (N_9982,N_7852,N_7653);
or U9983 (N_9983,N_7982,N_7629);
or U9984 (N_9984,N_8267,N_8158);
nor U9985 (N_9985,N_8161,N_8425);
nor U9986 (N_9986,N_8178,N_8229);
xnor U9987 (N_9987,N_7633,N_7980);
or U9988 (N_9988,N_8436,N_7794);
nand U9989 (N_9989,N_8267,N_7656);
nand U9990 (N_9990,N_8365,N_7659);
and U9991 (N_9991,N_7903,N_7509);
nor U9992 (N_9992,N_8226,N_8021);
nand U9993 (N_9993,N_7517,N_8702);
or U9994 (N_9994,N_7621,N_7973);
and U9995 (N_9995,N_7796,N_8080);
and U9996 (N_9996,N_8732,N_7679);
nor U9997 (N_9997,N_7775,N_7783);
and U9998 (N_9998,N_8501,N_7636);
nor U9999 (N_9999,N_8543,N_7772);
or U10000 (N_10000,N_9755,N_9447);
nand U10001 (N_10001,N_9488,N_9881);
and U10002 (N_10002,N_9534,N_9609);
or U10003 (N_10003,N_9984,N_9915);
nor U10004 (N_10004,N_8777,N_9162);
xnor U10005 (N_10005,N_9853,N_9882);
xnor U10006 (N_10006,N_9077,N_9401);
nor U10007 (N_10007,N_9250,N_9178);
and U10008 (N_10008,N_8985,N_9639);
and U10009 (N_10009,N_9117,N_8858);
or U10010 (N_10010,N_9318,N_9390);
or U10011 (N_10011,N_9678,N_8942);
xor U10012 (N_10012,N_9416,N_8982);
xnor U10013 (N_10013,N_9163,N_8945);
nor U10014 (N_10014,N_9215,N_9223);
xor U10015 (N_10015,N_9619,N_9253);
xnor U10016 (N_10016,N_9079,N_9830);
nor U10017 (N_10017,N_9995,N_9975);
xnor U10018 (N_10018,N_9378,N_9402);
nand U10019 (N_10019,N_8826,N_9779);
or U10020 (N_10020,N_9459,N_8892);
and U10021 (N_10021,N_9651,N_9232);
or U10022 (N_10022,N_8809,N_9707);
nand U10023 (N_10023,N_9880,N_9093);
nor U10024 (N_10024,N_9928,N_8946);
nor U10025 (N_10025,N_8851,N_8980);
or U10026 (N_10026,N_9665,N_9538);
nor U10027 (N_10027,N_8827,N_8893);
or U10028 (N_10028,N_9905,N_9652);
xor U10029 (N_10029,N_9344,N_9108);
or U10030 (N_10030,N_9544,N_9576);
nor U10031 (N_10031,N_9969,N_9645);
or U10032 (N_10032,N_8878,N_9875);
or U10033 (N_10033,N_9785,N_9759);
nand U10034 (N_10034,N_9091,N_9356);
nand U10035 (N_10035,N_9897,N_8753);
and U10036 (N_10036,N_9919,N_9903);
and U10037 (N_10037,N_8975,N_8795);
xor U10038 (N_10038,N_9238,N_9690);
and U10039 (N_10039,N_9864,N_8845);
xor U10040 (N_10040,N_9986,N_8863);
xor U10041 (N_10041,N_9725,N_9071);
or U10042 (N_10042,N_9099,N_9925);
or U10043 (N_10043,N_9778,N_9649);
xor U10044 (N_10044,N_8833,N_8859);
nand U10045 (N_10045,N_9513,N_8774);
or U10046 (N_10046,N_9002,N_9047);
nand U10047 (N_10047,N_9822,N_9304);
nand U10048 (N_10048,N_9789,N_9902);
or U10049 (N_10049,N_9073,N_8829);
and U10050 (N_10050,N_8909,N_9536);
and U10051 (N_10051,N_9739,N_9227);
nor U10052 (N_10052,N_9279,N_9632);
and U10053 (N_10053,N_9243,N_9572);
nor U10054 (N_10054,N_8802,N_8947);
nand U10055 (N_10055,N_8908,N_8790);
or U10056 (N_10056,N_9202,N_8883);
or U10057 (N_10057,N_9765,N_9696);
xor U10058 (N_10058,N_9611,N_9630);
and U10059 (N_10059,N_9452,N_8761);
nand U10060 (N_10060,N_9418,N_9821);
and U10061 (N_10061,N_9848,N_9620);
nand U10062 (N_10062,N_8978,N_9657);
xnor U10063 (N_10063,N_9434,N_9626);
xnor U10064 (N_10064,N_9886,N_9122);
xnor U10065 (N_10065,N_9140,N_8819);
xnor U10066 (N_10066,N_9371,N_8903);
xor U10067 (N_10067,N_9066,N_9599);
xor U10068 (N_10068,N_9815,N_9319);
nand U10069 (N_10069,N_8806,N_9834);
xnor U10070 (N_10070,N_9503,N_8758);
or U10071 (N_10071,N_9644,N_9019);
xnor U10072 (N_10072,N_9266,N_8838);
nand U10073 (N_10073,N_9176,N_9365);
nand U10074 (N_10074,N_9024,N_9682);
xor U10075 (N_10075,N_9070,N_9633);
or U10076 (N_10076,N_9222,N_9018);
xor U10077 (N_10077,N_9661,N_9912);
nand U10078 (N_10078,N_9263,N_9820);
nor U10079 (N_10079,N_9526,N_9315);
nand U10080 (N_10080,N_9990,N_9480);
and U10081 (N_10081,N_9866,N_8900);
or U10082 (N_10082,N_9942,N_9210);
or U10083 (N_10083,N_9305,N_9982);
xnor U10084 (N_10084,N_9484,N_9092);
or U10085 (N_10085,N_8800,N_9107);
xnor U10086 (N_10086,N_9945,N_9306);
or U10087 (N_10087,N_9320,N_9081);
xnor U10088 (N_10088,N_9088,N_9411);
nor U10089 (N_10089,N_9336,N_9930);
or U10090 (N_10090,N_8990,N_9141);
nand U10091 (N_10091,N_9728,N_9148);
and U10092 (N_10092,N_8765,N_9258);
xnor U10093 (N_10093,N_9680,N_9623);
xor U10094 (N_10094,N_8867,N_8803);
and U10095 (N_10095,N_9338,N_9339);
nor U10096 (N_10096,N_9030,N_9464);
nor U10097 (N_10097,N_9221,N_8939);
xnor U10098 (N_10098,N_9958,N_9884);
and U10099 (N_10099,N_9589,N_9396);
xor U10100 (N_10100,N_9515,N_9486);
and U10101 (N_10101,N_9494,N_9563);
nand U10102 (N_10102,N_9564,N_9686);
or U10103 (N_10103,N_8979,N_8970);
or U10104 (N_10104,N_9348,N_9642);
or U10105 (N_10105,N_8805,N_9677);
xor U10106 (N_10106,N_8813,N_9133);
or U10107 (N_10107,N_9417,N_9581);
or U10108 (N_10108,N_8993,N_8756);
and U10109 (N_10109,N_9722,N_9800);
xnor U10110 (N_10110,N_8962,N_9802);
xor U10111 (N_10111,N_9493,N_9357);
nand U10112 (N_10112,N_9774,N_8861);
nor U10113 (N_10113,N_9907,N_9399);
nor U10114 (N_10114,N_9807,N_9264);
nor U10115 (N_10115,N_9110,N_9374);
or U10116 (N_10116,N_9870,N_8966);
or U10117 (N_10117,N_9072,N_9780);
xnor U10118 (N_10118,N_9615,N_8968);
xor U10119 (N_10119,N_8879,N_8987);
nor U10120 (N_10120,N_8793,N_8943);
xor U10121 (N_10121,N_9597,N_8926);
nor U10122 (N_10122,N_9783,N_8843);
or U10123 (N_10123,N_9941,N_9653);
nand U10124 (N_10124,N_8991,N_9198);
nand U10125 (N_10125,N_9695,N_8839);
nand U10126 (N_10126,N_9571,N_9316);
nand U10127 (N_10127,N_9156,N_9049);
and U10128 (N_10128,N_9004,N_9596);
nor U10129 (N_10129,N_9750,N_8910);
xor U10130 (N_10130,N_9764,N_9520);
xor U10131 (N_10131,N_9234,N_9766);
nand U10132 (N_10132,N_8814,N_8828);
or U10133 (N_10133,N_9429,N_9667);
or U10134 (N_10134,N_9660,N_9455);
nand U10135 (N_10135,N_9753,N_9101);
xnor U10136 (N_10136,N_8872,N_8894);
and U10137 (N_10137,N_9655,N_9640);
nand U10138 (N_10138,N_9453,N_8799);
and U10139 (N_10139,N_9681,N_9960);
xnor U10140 (N_10140,N_9900,N_9809);
and U10141 (N_10141,N_9281,N_9300);
or U10142 (N_10142,N_9956,N_9174);
xnor U10143 (N_10143,N_9270,N_9718);
xor U10144 (N_10144,N_9616,N_9331);
nor U10145 (N_10145,N_9663,N_9372);
nor U10146 (N_10146,N_9191,N_9435);
nor U10147 (N_10147,N_9702,N_8999);
nor U10148 (N_10148,N_9804,N_9468);
and U10149 (N_10149,N_9512,N_9008);
nand U10150 (N_10150,N_9014,N_9309);
and U10151 (N_10151,N_9353,N_9738);
nand U10152 (N_10152,N_9608,N_9631);
and U10153 (N_10153,N_8823,N_9237);
nand U10154 (N_10154,N_9368,N_8850);
and U10155 (N_10155,N_9481,N_9400);
or U10156 (N_10156,N_9289,N_9173);
xor U10157 (N_10157,N_9491,N_9217);
and U10158 (N_10158,N_9323,N_9694);
or U10159 (N_10159,N_9314,N_8954);
or U10160 (N_10160,N_9966,N_9303);
or U10161 (N_10161,N_8889,N_9857);
and U10162 (N_10162,N_9384,N_9543);
nand U10163 (N_10163,N_9909,N_9557);
xnor U10164 (N_10164,N_8837,N_8890);
and U10165 (N_10165,N_9825,N_9734);
nor U10166 (N_10166,N_9171,N_9426);
or U10167 (N_10167,N_9444,N_9770);
xor U10168 (N_10168,N_9393,N_9283);
or U10169 (N_10169,N_9273,N_9559);
xor U10170 (N_10170,N_9656,N_9022);
xor U10171 (N_10171,N_9190,N_9860);
or U10172 (N_10172,N_9132,N_9170);
nand U10173 (N_10173,N_9366,N_9768);
nor U10174 (N_10174,N_9038,N_9150);
nor U10175 (N_10175,N_8825,N_8928);
or U10176 (N_10176,N_9425,N_9805);
nand U10177 (N_10177,N_9751,N_8791);
xor U10178 (N_10178,N_9508,N_9240);
and U10179 (N_10179,N_9182,N_9554);
nand U10180 (N_10180,N_8992,N_8807);
or U10181 (N_10181,N_9333,N_9826);
nor U10182 (N_10182,N_9391,N_9206);
xor U10183 (N_10183,N_9871,N_8857);
or U10184 (N_10184,N_9181,N_9861);
nand U10185 (N_10185,N_9749,N_9890);
xnor U10186 (N_10186,N_9095,N_9010);
nor U10187 (N_10187,N_9062,N_9763);
or U10188 (N_10188,N_8997,N_9985);
nor U10189 (N_10189,N_9836,N_8834);
nand U10190 (N_10190,N_9595,N_8754);
and U10191 (N_10191,N_9478,N_9016);
and U10192 (N_10192,N_8797,N_9917);
and U10193 (N_10193,N_9529,N_9726);
nand U10194 (N_10194,N_9601,N_9911);
nand U10195 (N_10195,N_9793,N_8760);
or U10196 (N_10196,N_9052,N_9298);
xor U10197 (N_10197,N_9475,N_8976);
xor U10198 (N_10198,N_9724,N_9105);
and U10199 (N_10199,N_9743,N_9899);
and U10200 (N_10200,N_9509,N_9185);
nand U10201 (N_10201,N_8916,N_8844);
nor U10202 (N_10202,N_9450,N_9838);
nand U10203 (N_10203,N_8776,N_9214);
and U10204 (N_10204,N_9082,N_9719);
or U10205 (N_10205,N_9844,N_9668);
and U10206 (N_10206,N_9456,N_8852);
and U10207 (N_10207,N_9961,N_9683);
nor U10208 (N_10208,N_9812,N_8952);
and U10209 (N_10209,N_9457,N_8762);
nand U10210 (N_10210,N_8788,N_8959);
nand U10211 (N_10211,N_9327,N_9388);
nor U10212 (N_10212,N_9127,N_9037);
nor U10213 (N_10213,N_9271,N_9313);
nor U10214 (N_10214,N_9102,N_9256);
and U10215 (N_10215,N_9054,N_9579);
and U10216 (N_10216,N_9155,N_9203);
nand U10217 (N_10217,N_9562,N_9748);
nor U10218 (N_10218,N_9275,N_9407);
xor U10219 (N_10219,N_8881,N_9041);
nand U10220 (N_10220,N_9204,N_9220);
nor U10221 (N_10221,N_9514,N_9561);
xor U10222 (N_10222,N_9065,N_9614);
or U10223 (N_10223,N_8832,N_9498);
xor U10224 (N_10224,N_9585,N_9260);
nor U10225 (N_10225,N_8918,N_9261);
xnor U10226 (N_10226,N_9879,N_9709);
nor U10227 (N_10227,N_9693,N_9566);
or U10228 (N_10228,N_9228,N_9403);
nor U10229 (N_10229,N_9700,N_9923);
nand U10230 (N_10230,N_9458,N_9873);
xnor U10231 (N_10231,N_8911,N_9292);
and U10232 (N_10232,N_8927,N_9075);
nor U10233 (N_10233,N_9560,N_8960);
or U10234 (N_10234,N_9090,N_9799);
and U10235 (N_10235,N_8860,N_8923);
xor U10236 (N_10236,N_9532,N_9962);
nand U10237 (N_10237,N_9021,N_9193);
or U10238 (N_10238,N_8773,N_9013);
xor U10239 (N_10239,N_9672,N_9762);
nor U10240 (N_10240,N_9184,N_9046);
xor U10241 (N_10241,N_9638,N_9888);
or U10242 (N_10242,N_9867,N_9469);
or U10243 (N_10243,N_9612,N_9239);
nand U10244 (N_10244,N_8783,N_9111);
xnor U10245 (N_10245,N_9541,N_8816);
and U10246 (N_10246,N_9134,N_9151);
nand U10247 (N_10247,N_9685,N_9125);
nor U10248 (N_10248,N_9364,N_9126);
nor U10249 (N_10249,N_9546,N_9023);
and U10250 (N_10250,N_9510,N_9282);
nand U10251 (N_10251,N_9476,N_8986);
nor U10252 (N_10252,N_9235,N_9974);
nor U10253 (N_10253,N_9811,N_9533);
or U10254 (N_10254,N_9967,N_9332);
nor U10255 (N_10255,N_9575,N_9518);
xnor U10256 (N_10256,N_9664,N_8898);
and U10257 (N_10257,N_9029,N_9659);
xnor U10258 (N_10258,N_9744,N_9257);
or U10259 (N_10259,N_9592,N_8840);
nand U10260 (N_10260,N_8804,N_9994);
nand U10261 (N_10261,N_9496,N_9628);
nor U10262 (N_10262,N_9036,N_9965);
nor U10263 (N_10263,N_9908,N_9251);
nor U10264 (N_10264,N_8841,N_9600);
nand U10265 (N_10265,N_8831,N_9499);
and U10266 (N_10266,N_9130,N_9831);
and U10267 (N_10267,N_9621,N_9487);
nor U10268 (N_10268,N_9436,N_8836);
nor U10269 (N_10269,N_8874,N_8775);
nor U10270 (N_10270,N_9218,N_9445);
and U10271 (N_10271,N_9790,N_9076);
or U10272 (N_10272,N_9121,N_9729);
nor U10273 (N_10273,N_9955,N_9325);
and U10274 (N_10274,N_8853,N_9293);
nand U10275 (N_10275,N_8932,N_9442);
nor U10276 (N_10276,N_9858,N_9714);
xnor U10277 (N_10277,N_9688,N_9195);
or U10278 (N_10278,N_9482,N_9837);
or U10279 (N_10279,N_9009,N_9872);
nor U10280 (N_10280,N_8794,N_9540);
xor U10281 (N_10281,N_9236,N_9159);
xor U10282 (N_10282,N_9662,N_9776);
or U10283 (N_10283,N_9771,N_9058);
xor U10284 (N_10284,N_9926,N_9177);
nand U10285 (N_10285,N_9330,N_8862);
nand U10286 (N_10286,N_9634,N_9818);
or U10287 (N_10287,N_9689,N_8873);
xnor U10288 (N_10288,N_8875,N_8907);
xnor U10289 (N_10289,N_9551,N_9658);
and U10290 (N_10290,N_9500,N_9308);
nor U10291 (N_10291,N_9167,N_9832);
nor U10292 (N_10292,N_9797,N_8815);
or U10293 (N_10293,N_9794,N_8965);
and U10294 (N_10294,N_9792,N_9415);
and U10295 (N_10295,N_9717,N_9343);
nor U10296 (N_10296,N_9892,N_9676);
or U10297 (N_10297,N_9395,N_8796);
xor U10298 (N_10298,N_8757,N_8937);
nor U10299 (N_10299,N_9843,N_9430);
nor U10300 (N_10300,N_9129,N_9856);
nand U10301 (N_10301,N_9404,N_9865);
and U10302 (N_10302,N_8798,N_9641);
and U10303 (N_10303,N_9020,N_9959);
xor U10304 (N_10304,N_9613,N_8995);
and U10305 (N_10305,N_9354,N_9976);
xor U10306 (N_10306,N_9118,N_9582);
nor U10307 (N_10307,N_9135,N_9521);
or U10308 (N_10308,N_9466,N_9212);
nor U10309 (N_10309,N_9267,N_9211);
xor U10310 (N_10310,N_8905,N_9269);
nor U10311 (N_10311,N_9978,N_9893);
or U10312 (N_10312,N_9078,N_8808);
nand U10313 (N_10313,N_9904,N_9603);
or U10314 (N_10314,N_9742,N_9060);
and U10315 (N_10315,N_9326,N_9624);
xnor U10316 (N_10316,N_9322,N_9869);
and U10317 (N_10317,N_8885,N_8958);
or U10318 (N_10318,N_8887,N_9158);
nand U10319 (N_10319,N_9782,N_9252);
nand U10320 (N_10320,N_9069,N_8811);
nand U10321 (N_10321,N_9542,N_9376);
nand U10322 (N_10322,N_9987,N_9495);
nor U10323 (N_10323,N_9045,N_9650);
or U10324 (N_10324,N_9720,N_9003);
nand U10325 (N_10325,N_9501,N_9196);
or U10326 (N_10326,N_8769,N_9610);
and U10327 (N_10327,N_9979,N_9671);
or U10328 (N_10328,N_9361,N_9943);
nand U10329 (N_10329,N_9687,N_9625);
xor U10330 (N_10330,N_9337,N_9100);
nor U10331 (N_10331,N_9321,N_9511);
nand U10332 (N_10332,N_8974,N_9033);
and U10333 (N_10333,N_9341,N_8755);
xnor U10334 (N_10334,N_9083,N_9876);
xnor U10335 (N_10335,N_8830,N_9670);
nand U10336 (N_10336,N_9711,N_9017);
nand U10337 (N_10337,N_8801,N_9936);
xnor U10338 (N_10338,N_8854,N_8864);
nor U10339 (N_10339,N_9972,N_9397);
xor U10340 (N_10340,N_9147,N_9980);
xnor U10341 (N_10341,N_9983,N_8914);
nand U10342 (N_10342,N_9276,N_9934);
and U10343 (N_10343,N_9334,N_8820);
xnor U10344 (N_10344,N_8785,N_9461);
xor U10345 (N_10345,N_9565,N_9183);
or U10346 (N_10346,N_9723,N_9446);
or U10347 (N_10347,N_9152,N_8988);
and U10348 (N_10348,N_9992,N_9692);
nor U10349 (N_10349,N_9817,N_8877);
nand U10350 (N_10350,N_9863,N_8977);
nor U10351 (N_10351,N_9859,N_8882);
and U10352 (N_10352,N_9027,N_9438);
or U10353 (N_10353,N_9583,N_9827);
nor U10354 (N_10354,N_8984,N_9377);
or U10355 (N_10355,N_8835,N_9473);
xnor U10356 (N_10356,N_8780,N_9654);
or U10357 (N_10357,N_9086,N_9087);
xor U10358 (N_10358,N_9577,N_9422);
and U10359 (N_10359,N_9971,N_9142);
nand U10360 (N_10360,N_9507,N_9849);
nand U10361 (N_10361,N_9519,N_9379);
nand U10362 (N_10362,N_9754,N_9026);
and U10363 (N_10363,N_9089,N_9816);
xor U10364 (N_10364,N_9349,N_9015);
nor U10365 (N_10365,N_9001,N_9197);
or U10366 (N_10366,N_9244,N_9898);
nor U10367 (N_10367,N_8933,N_9067);
nor U10368 (N_10368,N_9405,N_8770);
nand U10369 (N_10369,N_9835,N_9727);
and U10370 (N_10370,N_9999,N_9342);
nor U10371 (N_10371,N_9381,N_9548);
nor U10372 (N_10372,N_9704,N_8963);
or U10373 (N_10373,N_9635,N_9440);
nor U10374 (N_10374,N_9057,N_9539);
and U10375 (N_10375,N_8886,N_9398);
or U10376 (N_10376,N_9957,N_9901);
or U10377 (N_10377,N_9767,N_8935);
or U10378 (N_10378,N_9741,N_9299);
xor U10379 (N_10379,N_9246,N_8767);
or U10380 (N_10380,N_9492,N_9179);
and U10381 (N_10381,N_8981,N_9225);
or U10382 (N_10382,N_9031,N_8964);
nor U10383 (N_10383,N_9460,N_9359);
nor U10384 (N_10384,N_9850,N_9553);
nor U10385 (N_10385,N_9347,N_9752);
xnor U10386 (N_10386,N_9721,N_9437);
xor U10387 (N_10387,N_9061,N_8789);
and U10388 (N_10388,N_9932,N_9549);
or U10389 (N_10389,N_9109,N_9906);
xor U10390 (N_10390,N_9697,N_9420);
nor U10391 (N_10391,N_9701,N_8822);
and U10392 (N_10392,N_9259,N_9977);
nand U10393 (N_10393,N_9814,N_8884);
xor U10394 (N_10394,N_8876,N_9032);
xnor U10395 (N_10395,N_8781,N_9998);
or U10396 (N_10396,N_9736,N_8759);
nand U10397 (N_10397,N_8866,N_9868);
xnor U10398 (N_10398,N_9255,N_8996);
xnor U10399 (N_10399,N_9042,N_9796);
nor U10400 (N_10400,N_9483,N_9028);
nor U10401 (N_10401,N_8944,N_9847);
nand U10402 (N_10402,N_9007,N_9209);
and U10403 (N_10403,N_8782,N_9242);
nand U10404 (N_10404,N_9991,N_8951);
nand U10405 (N_10405,N_9933,N_9840);
and U10406 (N_10406,N_9439,N_9997);
nand U10407 (N_10407,N_9527,N_9307);
xnor U10408 (N_10408,N_9213,N_9410);
nor U10409 (N_10409,N_9485,N_9737);
nand U10410 (N_10410,N_9747,N_8763);
nand U10411 (N_10411,N_9922,N_9039);
nand U10412 (N_10412,N_9443,N_9428);
xor U10413 (N_10413,N_9408,N_9187);
and U10414 (N_10414,N_9120,N_9708);
and U10415 (N_10415,N_9352,N_9556);
and U10416 (N_10416,N_9947,N_8949);
or U10417 (N_10417,N_8940,N_9363);
and U10418 (N_10418,N_9895,N_9346);
and U10419 (N_10419,N_9691,N_9643);
xnor U10420 (N_10420,N_9157,N_8768);
and U10421 (N_10421,N_8912,N_9387);
or U10422 (N_10422,N_8924,N_9114);
nand U10423 (N_10423,N_9192,N_9913);
xnor U10424 (N_10424,N_8934,N_9138);
or U10425 (N_10425,N_9231,N_9772);
nor U10426 (N_10426,N_9703,N_9383);
and U10427 (N_10427,N_9113,N_9716);
and U10428 (N_10428,N_9216,N_9679);
xor U10429 (N_10429,N_9940,N_9705);
and U10430 (N_10430,N_9851,N_9451);
xor U10431 (N_10431,N_9537,N_9784);
and U10432 (N_10432,N_9948,N_9698);
xor U10433 (N_10433,N_8901,N_9929);
xnor U10434 (N_10434,N_9732,N_9535);
and U10435 (N_10435,N_9277,N_9788);
and U10436 (N_10436,N_8817,N_8888);
nand U10437 (N_10437,N_9385,N_9116);
xor U10438 (N_10438,N_9874,N_9064);
or U10439 (N_10439,N_9637,N_9050);
or U10440 (N_10440,N_9489,N_8972);
nor U10441 (N_10441,N_9201,N_9011);
or U10442 (N_10442,N_9935,N_9761);
xnor U10443 (N_10443,N_8871,N_8750);
nor U10444 (N_10444,N_9301,N_9877);
nand U10445 (N_10445,N_9097,N_8810);
nor U10446 (N_10446,N_8771,N_9646);
nand U10447 (N_10447,N_8906,N_9944);
nand U10448 (N_10448,N_9074,N_9590);
and U10449 (N_10449,N_8921,N_9291);
nor U10450 (N_10450,N_9249,N_9845);
or U10451 (N_10451,N_9294,N_9351);
xnor U10452 (N_10452,N_9813,N_9593);
and U10453 (N_10453,N_9712,N_8897);
or U10454 (N_10454,N_9085,N_9477);
or U10455 (N_10455,N_9474,N_9574);
nor U10456 (N_10456,N_9648,N_9080);
or U10457 (N_10457,N_9842,N_9855);
or U10458 (N_10458,N_9427,N_9740);
nor U10459 (N_10459,N_8917,N_9528);
xor U10460 (N_10460,N_9505,N_9550);
xor U10461 (N_10461,N_9106,N_9810);
or U10462 (N_10462,N_9803,N_9618);
nor U10463 (N_10463,N_9569,N_9471);
nor U10464 (N_10464,N_9675,N_9161);
and U10465 (N_10465,N_9153,N_9841);
xor U10466 (N_10466,N_9931,N_8957);
nand U10467 (N_10467,N_9946,N_9523);
or U10468 (N_10468,N_9226,N_8904);
nand U10469 (N_10469,N_8953,N_8766);
or U10470 (N_10470,N_9448,N_9302);
nand U10471 (N_10471,N_9733,N_9139);
or U10472 (N_10472,N_9059,N_9605);
nor U10473 (N_10473,N_8821,N_9449);
nand U10474 (N_10474,N_9887,N_9604);
nor U10475 (N_10475,N_9517,N_8920);
and U10476 (N_10476,N_9801,N_9465);
nand U10477 (N_10477,N_9918,N_8869);
xor U10478 (N_10478,N_8848,N_9669);
or U10479 (N_10479,N_9823,N_9358);
xnor U10480 (N_10480,N_9262,N_9136);
nor U10481 (N_10481,N_9629,N_9852);
nor U10482 (N_10482,N_9380,N_9287);
nor U10483 (N_10483,N_9207,N_9573);
nor U10484 (N_10484,N_9188,N_9735);
xor U10485 (N_10485,N_9570,N_9144);
or U10486 (N_10486,N_8998,N_9854);
and U10487 (N_10487,N_9025,N_9128);
nor U10488 (N_10488,N_9787,N_9627);
or U10489 (N_10489,N_9413,N_8941);
nand U10490 (N_10490,N_8812,N_8913);
and U10491 (N_10491,N_9145,N_8956);
and U10492 (N_10492,N_8784,N_9149);
nand U10493 (N_10493,N_9914,N_9937);
and U10494 (N_10494,N_9164,N_9916);
or U10495 (N_10495,N_9272,N_9617);
nor U10496 (N_10496,N_8865,N_9254);
or U10497 (N_10497,N_9168,N_9103);
nand U10498 (N_10498,N_9175,N_9394);
xor U10499 (N_10499,N_9268,N_9808);
or U10500 (N_10500,N_9392,N_9715);
and U10501 (N_10501,N_9286,N_9345);
xor U10502 (N_10502,N_8969,N_9647);
or U10503 (N_10503,N_9927,N_9806);
nand U10504 (N_10504,N_9938,N_9317);
and U10505 (N_10505,N_9414,N_9964);
and U10506 (N_10506,N_9194,N_9584);
xor U10507 (N_10507,N_9910,N_8849);
nor U10508 (N_10508,N_9012,N_8919);
xnor U10509 (N_10509,N_9189,N_9939);
and U10510 (N_10510,N_9791,N_9829);
xnor U10511 (N_10511,N_9757,N_8915);
or U10512 (N_10512,N_9706,N_8994);
and U10513 (N_10513,N_9710,N_8930);
and U10514 (N_10514,N_9274,N_9516);
nand U10515 (N_10515,N_9123,N_9795);
or U10516 (N_10516,N_8787,N_9324);
nand U10517 (N_10517,N_9172,N_9921);
xnor U10518 (N_10518,N_8778,N_9530);
or U10519 (N_10519,N_8936,N_9781);
or U10520 (N_10520,N_9056,N_9247);
xnor U10521 (N_10521,N_9296,N_9051);
xor U10522 (N_10522,N_9522,N_9409);
nand U10523 (N_10523,N_9424,N_8772);
nand U10524 (N_10524,N_9048,N_9200);
xor U10525 (N_10525,N_9112,N_9362);
and U10526 (N_10526,N_9777,N_9894);
or U10527 (N_10527,N_9104,N_9745);
xor U10528 (N_10528,N_8880,N_9470);
xnor U10529 (N_10529,N_9288,N_9005);
nand U10530 (N_10530,N_9889,N_9479);
xnor U10531 (N_10531,N_9166,N_9040);
or U10532 (N_10532,N_9098,N_8855);
and U10533 (N_10533,N_9230,N_9970);
nand U10534 (N_10534,N_9578,N_9454);
nand U10535 (N_10535,N_9310,N_9472);
nand U10536 (N_10536,N_9160,N_9545);
nor U10537 (N_10537,N_9094,N_8818);
nor U10538 (N_10538,N_9839,N_9006);
nand U10539 (N_10539,N_9328,N_9245);
xnor U10540 (N_10540,N_8948,N_9423);
and U10541 (N_10541,N_9502,N_8971);
nand U10542 (N_10542,N_9035,N_9199);
xnor U10543 (N_10543,N_9055,N_9833);
nand U10544 (N_10544,N_9775,N_9205);
nand U10545 (N_10545,N_9208,N_8895);
xor U10546 (N_10546,N_9567,N_9878);
nor U10547 (N_10547,N_8922,N_9285);
xnor U10548 (N_10548,N_9146,N_9773);
xnor U10549 (N_10549,N_9996,N_8902);
and U10550 (N_10550,N_9137,N_8989);
or U10551 (N_10551,N_9756,N_9524);
nand U10552 (N_10552,N_9355,N_9369);
nand U10553 (N_10553,N_8967,N_9034);
nand U10554 (N_10554,N_9043,N_9607);
or U10555 (N_10555,N_9953,N_9386);
xnor U10556 (N_10556,N_9731,N_9636);
xnor U10557 (N_10557,N_9412,N_9993);
or U10558 (N_10558,N_8983,N_9504);
nor U10559 (N_10559,N_9713,N_9896);
and U10560 (N_10560,N_8856,N_9598);
xor U10561 (N_10561,N_9819,N_9862);
nand U10562 (N_10562,N_9673,N_8870);
nand U10563 (N_10563,N_9096,N_9143);
nor U10564 (N_10564,N_9406,N_9989);
xor U10565 (N_10565,N_9891,N_9265);
and U10566 (N_10566,N_9591,N_9963);
nor U10567 (N_10567,N_8847,N_9115);
xnor U10568 (N_10568,N_9952,N_9746);
nor U10569 (N_10569,N_8929,N_8896);
and U10570 (N_10570,N_8751,N_9463);
or U10571 (N_10571,N_9920,N_9131);
nor U10572 (N_10572,N_9084,N_8786);
xor U10573 (N_10573,N_9280,N_9382);
xor U10574 (N_10574,N_9846,N_9490);
and U10575 (N_10575,N_9506,N_8824);
nand U10576 (N_10576,N_9186,N_9547);
and U10577 (N_10577,N_8842,N_9433);
and U10578 (N_10578,N_9389,N_9360);
and U10579 (N_10579,N_9594,N_9241);
or U10580 (N_10580,N_9335,N_8961);
nor U10581 (N_10581,N_9431,N_9312);
and U10582 (N_10582,N_9284,N_9950);
xor U10583 (N_10583,N_9988,N_9370);
xor U10584 (N_10584,N_9531,N_8891);
and U10585 (N_10585,N_9419,N_9165);
or U10586 (N_10586,N_9568,N_8868);
nand U10587 (N_10587,N_9180,N_9730);
xnor U10588 (N_10588,N_9684,N_9053);
and U10589 (N_10589,N_9044,N_9350);
nand U10590 (N_10590,N_9068,N_9000);
and U10591 (N_10591,N_9219,N_9233);
nor U10592 (N_10592,N_9373,N_9311);
nand U10593 (N_10593,N_9555,N_9119);
and U10594 (N_10594,N_9375,N_9169);
and U10595 (N_10595,N_9552,N_9497);
nand U10596 (N_10596,N_9949,N_8792);
nand U10597 (N_10597,N_8779,N_9954);
nand U10598 (N_10598,N_9278,N_8973);
or U10599 (N_10599,N_9981,N_9828);
xor U10600 (N_10600,N_9329,N_9786);
or U10601 (N_10601,N_9666,N_9154);
nor U10602 (N_10602,N_9586,N_8931);
and U10603 (N_10603,N_9758,N_9699);
and U10604 (N_10604,N_9798,N_8846);
and U10605 (N_10605,N_9340,N_9606);
nand U10606 (N_10606,N_9588,N_9224);
nor U10607 (N_10607,N_9924,N_9622);
nor U10608 (N_10608,N_9968,N_9824);
nand U10609 (N_10609,N_9367,N_9290);
nand U10610 (N_10610,N_9124,N_9558);
or U10611 (N_10611,N_9462,N_9580);
and U10612 (N_10612,N_9602,N_9295);
and U10613 (N_10613,N_8938,N_9297);
or U10614 (N_10614,N_9063,N_9229);
nor U10615 (N_10615,N_9432,N_9951);
xnor U10616 (N_10616,N_9973,N_9467);
nand U10617 (N_10617,N_9883,N_9885);
nor U10618 (N_10618,N_9587,N_9769);
or U10619 (N_10619,N_8955,N_8752);
nor U10620 (N_10620,N_8925,N_8764);
and U10621 (N_10621,N_9421,N_9760);
or U10622 (N_10622,N_9441,N_9248);
and U10623 (N_10623,N_9525,N_8950);
xor U10624 (N_10624,N_9674,N_8899);
nor U10625 (N_10625,N_9708,N_9049);
and U10626 (N_10626,N_8755,N_9651);
nor U10627 (N_10627,N_9046,N_9048);
and U10628 (N_10628,N_9163,N_9856);
nand U10629 (N_10629,N_9788,N_9131);
nand U10630 (N_10630,N_9116,N_9746);
and U10631 (N_10631,N_9932,N_8976);
nor U10632 (N_10632,N_9770,N_9517);
nor U10633 (N_10633,N_8801,N_9753);
xor U10634 (N_10634,N_9243,N_9695);
xor U10635 (N_10635,N_8793,N_9615);
xor U10636 (N_10636,N_9152,N_9711);
xor U10637 (N_10637,N_9615,N_9435);
nor U10638 (N_10638,N_8838,N_9541);
and U10639 (N_10639,N_9468,N_9058);
and U10640 (N_10640,N_9639,N_9771);
nand U10641 (N_10641,N_9650,N_9206);
nand U10642 (N_10642,N_9958,N_9839);
and U10643 (N_10643,N_9709,N_9293);
nand U10644 (N_10644,N_9152,N_9367);
nor U10645 (N_10645,N_9880,N_9293);
xor U10646 (N_10646,N_9588,N_9294);
nor U10647 (N_10647,N_9507,N_8834);
and U10648 (N_10648,N_9816,N_9421);
nor U10649 (N_10649,N_9869,N_9591);
nand U10650 (N_10650,N_9092,N_8767);
nor U10651 (N_10651,N_9679,N_9800);
xnor U10652 (N_10652,N_9633,N_9799);
nand U10653 (N_10653,N_8841,N_9404);
and U10654 (N_10654,N_9236,N_9709);
xnor U10655 (N_10655,N_9999,N_9197);
xor U10656 (N_10656,N_9315,N_9480);
or U10657 (N_10657,N_9016,N_8784);
nand U10658 (N_10658,N_8950,N_9569);
nor U10659 (N_10659,N_9447,N_9381);
nand U10660 (N_10660,N_9635,N_9505);
nor U10661 (N_10661,N_9558,N_9634);
nand U10662 (N_10662,N_8875,N_8957);
or U10663 (N_10663,N_9498,N_8944);
xnor U10664 (N_10664,N_8869,N_9176);
xor U10665 (N_10665,N_8844,N_8910);
nor U10666 (N_10666,N_9502,N_9058);
xnor U10667 (N_10667,N_9832,N_9079);
nand U10668 (N_10668,N_9679,N_9289);
or U10669 (N_10669,N_9194,N_9550);
nand U10670 (N_10670,N_9063,N_9233);
or U10671 (N_10671,N_9212,N_9072);
xor U10672 (N_10672,N_9233,N_9499);
and U10673 (N_10673,N_9359,N_9458);
xnor U10674 (N_10674,N_9804,N_9486);
and U10675 (N_10675,N_9123,N_9277);
nand U10676 (N_10676,N_9068,N_9017);
xor U10677 (N_10677,N_8916,N_9341);
and U10678 (N_10678,N_8774,N_8798);
xor U10679 (N_10679,N_9887,N_9830);
and U10680 (N_10680,N_9119,N_9762);
or U10681 (N_10681,N_9276,N_8808);
nor U10682 (N_10682,N_9209,N_9445);
nor U10683 (N_10683,N_9893,N_9397);
nand U10684 (N_10684,N_9304,N_9587);
nor U10685 (N_10685,N_9000,N_9880);
xnor U10686 (N_10686,N_9235,N_9449);
nor U10687 (N_10687,N_9968,N_8931);
nor U10688 (N_10688,N_9989,N_8842);
nor U10689 (N_10689,N_9727,N_9029);
and U10690 (N_10690,N_9632,N_9147);
nor U10691 (N_10691,N_8836,N_9149);
nand U10692 (N_10692,N_9312,N_9726);
nor U10693 (N_10693,N_9239,N_9802);
and U10694 (N_10694,N_9640,N_9547);
and U10695 (N_10695,N_9261,N_8850);
and U10696 (N_10696,N_8928,N_9077);
xor U10697 (N_10697,N_9112,N_9768);
nand U10698 (N_10698,N_9390,N_9702);
nand U10699 (N_10699,N_9169,N_9581);
nand U10700 (N_10700,N_9140,N_8845);
nand U10701 (N_10701,N_9854,N_9185);
or U10702 (N_10702,N_8854,N_9415);
nor U10703 (N_10703,N_9299,N_9329);
nand U10704 (N_10704,N_8829,N_8820);
and U10705 (N_10705,N_9402,N_8791);
and U10706 (N_10706,N_8964,N_9463);
or U10707 (N_10707,N_9657,N_8990);
nand U10708 (N_10708,N_9661,N_9509);
and U10709 (N_10709,N_8765,N_9787);
or U10710 (N_10710,N_9801,N_9366);
xor U10711 (N_10711,N_9397,N_8927);
xor U10712 (N_10712,N_8815,N_8920);
or U10713 (N_10713,N_8858,N_9583);
and U10714 (N_10714,N_9643,N_9759);
nor U10715 (N_10715,N_9997,N_9390);
xnor U10716 (N_10716,N_9213,N_9379);
xor U10717 (N_10717,N_9941,N_8787);
nor U10718 (N_10718,N_9394,N_9598);
or U10719 (N_10719,N_9163,N_9331);
nor U10720 (N_10720,N_9356,N_8762);
xor U10721 (N_10721,N_9266,N_9680);
or U10722 (N_10722,N_9597,N_9805);
or U10723 (N_10723,N_9312,N_9870);
and U10724 (N_10724,N_8768,N_9455);
nand U10725 (N_10725,N_9558,N_8925);
nand U10726 (N_10726,N_9784,N_9618);
xnor U10727 (N_10727,N_9200,N_9613);
or U10728 (N_10728,N_9052,N_9656);
or U10729 (N_10729,N_9755,N_8945);
xor U10730 (N_10730,N_9711,N_9182);
nand U10731 (N_10731,N_8872,N_9621);
and U10732 (N_10732,N_9586,N_9992);
nand U10733 (N_10733,N_9295,N_8925);
and U10734 (N_10734,N_9169,N_8900);
and U10735 (N_10735,N_8805,N_9139);
or U10736 (N_10736,N_9153,N_9361);
and U10737 (N_10737,N_8943,N_9957);
nor U10738 (N_10738,N_8752,N_9557);
nand U10739 (N_10739,N_9452,N_9973);
nor U10740 (N_10740,N_9158,N_9224);
or U10741 (N_10741,N_8822,N_9690);
and U10742 (N_10742,N_9162,N_9547);
or U10743 (N_10743,N_9857,N_9017);
xor U10744 (N_10744,N_9852,N_9441);
nor U10745 (N_10745,N_9619,N_9167);
or U10746 (N_10746,N_9003,N_9766);
nor U10747 (N_10747,N_8969,N_9148);
nor U10748 (N_10748,N_9524,N_8922);
or U10749 (N_10749,N_9528,N_9937);
nand U10750 (N_10750,N_9595,N_9687);
or U10751 (N_10751,N_8788,N_9227);
xor U10752 (N_10752,N_9552,N_8950);
nand U10753 (N_10753,N_8927,N_9279);
xnor U10754 (N_10754,N_9240,N_8786);
nor U10755 (N_10755,N_8874,N_9901);
nand U10756 (N_10756,N_9700,N_9245);
and U10757 (N_10757,N_9306,N_9152);
nor U10758 (N_10758,N_9040,N_9436);
xor U10759 (N_10759,N_9310,N_8967);
nor U10760 (N_10760,N_8978,N_8831);
nand U10761 (N_10761,N_9764,N_9363);
xnor U10762 (N_10762,N_9388,N_9859);
nor U10763 (N_10763,N_9405,N_8786);
or U10764 (N_10764,N_9185,N_9060);
or U10765 (N_10765,N_9849,N_9590);
nor U10766 (N_10766,N_9653,N_9536);
or U10767 (N_10767,N_9925,N_9958);
xnor U10768 (N_10768,N_8919,N_9270);
nor U10769 (N_10769,N_9813,N_9316);
xor U10770 (N_10770,N_9586,N_9458);
or U10771 (N_10771,N_8793,N_9168);
and U10772 (N_10772,N_9096,N_9667);
and U10773 (N_10773,N_9152,N_9106);
xor U10774 (N_10774,N_9443,N_9346);
xor U10775 (N_10775,N_8864,N_9873);
nor U10776 (N_10776,N_8945,N_9636);
xor U10777 (N_10777,N_9158,N_9576);
or U10778 (N_10778,N_9069,N_9880);
nand U10779 (N_10779,N_9812,N_9623);
and U10780 (N_10780,N_9788,N_9031);
or U10781 (N_10781,N_9773,N_9296);
nor U10782 (N_10782,N_9040,N_9445);
xnor U10783 (N_10783,N_9771,N_9241);
and U10784 (N_10784,N_9508,N_9229);
or U10785 (N_10785,N_9112,N_9434);
nor U10786 (N_10786,N_9855,N_9501);
and U10787 (N_10787,N_9328,N_9337);
or U10788 (N_10788,N_8869,N_9600);
xnor U10789 (N_10789,N_9401,N_9298);
and U10790 (N_10790,N_8950,N_9958);
xor U10791 (N_10791,N_9785,N_9349);
and U10792 (N_10792,N_9481,N_9638);
or U10793 (N_10793,N_9266,N_9372);
nand U10794 (N_10794,N_8802,N_9277);
and U10795 (N_10795,N_8761,N_9426);
or U10796 (N_10796,N_8759,N_9372);
xnor U10797 (N_10797,N_9447,N_9201);
nand U10798 (N_10798,N_9763,N_8833);
nand U10799 (N_10799,N_9194,N_9635);
and U10800 (N_10800,N_9103,N_9327);
nor U10801 (N_10801,N_9977,N_9872);
and U10802 (N_10802,N_9004,N_9698);
and U10803 (N_10803,N_9535,N_9524);
nor U10804 (N_10804,N_8841,N_8755);
nand U10805 (N_10805,N_9465,N_8956);
xnor U10806 (N_10806,N_8948,N_8987);
nor U10807 (N_10807,N_9467,N_8918);
nand U10808 (N_10808,N_9070,N_8850);
and U10809 (N_10809,N_9523,N_9879);
nor U10810 (N_10810,N_9652,N_9908);
and U10811 (N_10811,N_9249,N_9564);
and U10812 (N_10812,N_9070,N_9181);
and U10813 (N_10813,N_9339,N_9581);
xnor U10814 (N_10814,N_9288,N_9714);
or U10815 (N_10815,N_9103,N_9188);
xnor U10816 (N_10816,N_9171,N_8959);
xnor U10817 (N_10817,N_9501,N_9036);
xor U10818 (N_10818,N_8813,N_9293);
or U10819 (N_10819,N_8819,N_9879);
nor U10820 (N_10820,N_9250,N_9879);
xnor U10821 (N_10821,N_8768,N_8956);
nand U10822 (N_10822,N_9890,N_9280);
nand U10823 (N_10823,N_9210,N_8925);
and U10824 (N_10824,N_9997,N_9127);
nand U10825 (N_10825,N_8783,N_8923);
or U10826 (N_10826,N_9235,N_9111);
nor U10827 (N_10827,N_9161,N_9358);
and U10828 (N_10828,N_9255,N_9834);
or U10829 (N_10829,N_9568,N_9933);
xor U10830 (N_10830,N_9355,N_9619);
nand U10831 (N_10831,N_9777,N_9825);
nor U10832 (N_10832,N_9641,N_9032);
xnor U10833 (N_10833,N_9007,N_9903);
nor U10834 (N_10834,N_8868,N_9996);
xor U10835 (N_10835,N_9019,N_9016);
or U10836 (N_10836,N_9474,N_8849);
xnor U10837 (N_10837,N_9431,N_8796);
and U10838 (N_10838,N_9405,N_9810);
nor U10839 (N_10839,N_9849,N_9900);
or U10840 (N_10840,N_8780,N_9169);
and U10841 (N_10841,N_9484,N_9628);
xor U10842 (N_10842,N_9474,N_9987);
nand U10843 (N_10843,N_8881,N_9154);
nor U10844 (N_10844,N_9480,N_8952);
and U10845 (N_10845,N_9408,N_9907);
xnor U10846 (N_10846,N_9948,N_9527);
and U10847 (N_10847,N_9713,N_8998);
nand U10848 (N_10848,N_9632,N_8904);
and U10849 (N_10849,N_8771,N_9593);
nand U10850 (N_10850,N_9210,N_9248);
nand U10851 (N_10851,N_9596,N_8988);
and U10852 (N_10852,N_9178,N_9069);
nor U10853 (N_10853,N_9637,N_9918);
or U10854 (N_10854,N_9530,N_9625);
nand U10855 (N_10855,N_9554,N_9584);
nand U10856 (N_10856,N_9266,N_9892);
nand U10857 (N_10857,N_9948,N_9004);
or U10858 (N_10858,N_9315,N_8805);
nand U10859 (N_10859,N_9891,N_9854);
nand U10860 (N_10860,N_8788,N_9259);
and U10861 (N_10861,N_9544,N_9365);
xor U10862 (N_10862,N_9795,N_9420);
xor U10863 (N_10863,N_8896,N_8980);
xnor U10864 (N_10864,N_9795,N_8991);
and U10865 (N_10865,N_9561,N_9413);
xor U10866 (N_10866,N_9165,N_9840);
or U10867 (N_10867,N_9404,N_9773);
nand U10868 (N_10868,N_9664,N_9992);
xor U10869 (N_10869,N_8974,N_9849);
nor U10870 (N_10870,N_9408,N_9221);
xor U10871 (N_10871,N_8890,N_9884);
nor U10872 (N_10872,N_9567,N_9441);
and U10873 (N_10873,N_9207,N_9436);
nor U10874 (N_10874,N_9851,N_9259);
nor U10875 (N_10875,N_9777,N_8890);
nand U10876 (N_10876,N_8989,N_9325);
xor U10877 (N_10877,N_9727,N_9228);
and U10878 (N_10878,N_9197,N_9897);
or U10879 (N_10879,N_9777,N_9942);
nor U10880 (N_10880,N_9489,N_9285);
nor U10881 (N_10881,N_8923,N_8827);
or U10882 (N_10882,N_9473,N_9832);
or U10883 (N_10883,N_9776,N_8792);
xor U10884 (N_10884,N_9712,N_9412);
nand U10885 (N_10885,N_9834,N_9299);
or U10886 (N_10886,N_9328,N_9665);
xor U10887 (N_10887,N_9540,N_9565);
or U10888 (N_10888,N_9216,N_9688);
nor U10889 (N_10889,N_8941,N_9083);
nand U10890 (N_10890,N_8925,N_9226);
or U10891 (N_10891,N_9481,N_9489);
and U10892 (N_10892,N_9150,N_9720);
or U10893 (N_10893,N_9070,N_9852);
xor U10894 (N_10894,N_8843,N_9369);
and U10895 (N_10895,N_9066,N_9663);
nand U10896 (N_10896,N_9958,N_9123);
xnor U10897 (N_10897,N_9036,N_9651);
nand U10898 (N_10898,N_9437,N_8879);
xor U10899 (N_10899,N_9580,N_8851);
or U10900 (N_10900,N_9649,N_9231);
nand U10901 (N_10901,N_9725,N_9426);
nor U10902 (N_10902,N_8889,N_9553);
xnor U10903 (N_10903,N_8915,N_9714);
nor U10904 (N_10904,N_9574,N_9033);
nand U10905 (N_10905,N_9639,N_9076);
nor U10906 (N_10906,N_9751,N_9352);
xnor U10907 (N_10907,N_9765,N_8842);
xor U10908 (N_10908,N_9486,N_9077);
nor U10909 (N_10909,N_9390,N_9066);
nor U10910 (N_10910,N_9353,N_9852);
nand U10911 (N_10911,N_9185,N_9317);
and U10912 (N_10912,N_8936,N_9777);
xnor U10913 (N_10913,N_9149,N_9362);
xnor U10914 (N_10914,N_9898,N_9488);
nor U10915 (N_10915,N_9485,N_9519);
nor U10916 (N_10916,N_9559,N_9993);
xor U10917 (N_10917,N_9086,N_9537);
or U10918 (N_10918,N_8983,N_9086);
nor U10919 (N_10919,N_8781,N_9306);
xor U10920 (N_10920,N_9212,N_9464);
and U10921 (N_10921,N_9320,N_8905);
or U10922 (N_10922,N_9315,N_9398);
xnor U10923 (N_10923,N_9025,N_9140);
or U10924 (N_10924,N_9430,N_9661);
or U10925 (N_10925,N_9902,N_9762);
or U10926 (N_10926,N_8808,N_9845);
nand U10927 (N_10927,N_9026,N_9367);
xor U10928 (N_10928,N_9520,N_9700);
xor U10929 (N_10929,N_9254,N_9374);
nor U10930 (N_10930,N_9008,N_9893);
nor U10931 (N_10931,N_8838,N_8785);
xnor U10932 (N_10932,N_8807,N_9159);
xor U10933 (N_10933,N_8924,N_9285);
nor U10934 (N_10934,N_9963,N_8802);
nand U10935 (N_10935,N_9276,N_9747);
nor U10936 (N_10936,N_9573,N_9040);
and U10937 (N_10937,N_9416,N_9461);
xnor U10938 (N_10938,N_9426,N_9493);
or U10939 (N_10939,N_9192,N_9033);
nand U10940 (N_10940,N_9855,N_9119);
nor U10941 (N_10941,N_9627,N_8908);
or U10942 (N_10942,N_8887,N_8894);
nand U10943 (N_10943,N_8804,N_9084);
nand U10944 (N_10944,N_9108,N_8950);
xnor U10945 (N_10945,N_9386,N_9660);
xnor U10946 (N_10946,N_9422,N_9938);
and U10947 (N_10947,N_9401,N_9868);
nor U10948 (N_10948,N_9527,N_9090);
nor U10949 (N_10949,N_9545,N_8766);
xor U10950 (N_10950,N_9092,N_8991);
or U10951 (N_10951,N_9902,N_8752);
and U10952 (N_10952,N_9095,N_9757);
xnor U10953 (N_10953,N_8777,N_9669);
and U10954 (N_10954,N_9763,N_9487);
nor U10955 (N_10955,N_9389,N_9407);
or U10956 (N_10956,N_9917,N_9024);
nand U10957 (N_10957,N_9262,N_9374);
xor U10958 (N_10958,N_9760,N_9630);
nor U10959 (N_10959,N_9349,N_9483);
nor U10960 (N_10960,N_9929,N_9434);
nor U10961 (N_10961,N_8852,N_8859);
and U10962 (N_10962,N_8926,N_9620);
xnor U10963 (N_10963,N_9047,N_9398);
nor U10964 (N_10964,N_9371,N_9648);
and U10965 (N_10965,N_9748,N_8947);
xnor U10966 (N_10966,N_9387,N_9092);
xnor U10967 (N_10967,N_9626,N_9590);
nand U10968 (N_10968,N_9154,N_9342);
nor U10969 (N_10969,N_9839,N_8815);
and U10970 (N_10970,N_8922,N_9457);
nor U10971 (N_10971,N_9116,N_9535);
and U10972 (N_10972,N_9689,N_9955);
xor U10973 (N_10973,N_9098,N_9799);
and U10974 (N_10974,N_9549,N_9129);
and U10975 (N_10975,N_9178,N_8833);
or U10976 (N_10976,N_9253,N_9744);
nor U10977 (N_10977,N_9256,N_9747);
nor U10978 (N_10978,N_9989,N_9379);
xnor U10979 (N_10979,N_9360,N_9771);
nand U10980 (N_10980,N_9912,N_9686);
nand U10981 (N_10981,N_9248,N_8781);
or U10982 (N_10982,N_8956,N_9478);
xor U10983 (N_10983,N_9117,N_8799);
xnor U10984 (N_10984,N_8811,N_9626);
or U10985 (N_10985,N_9196,N_9536);
nand U10986 (N_10986,N_8921,N_9114);
and U10987 (N_10987,N_9242,N_9040);
nor U10988 (N_10988,N_9716,N_8814);
nand U10989 (N_10989,N_9140,N_8872);
nand U10990 (N_10990,N_9271,N_8951);
or U10991 (N_10991,N_9029,N_9106);
nand U10992 (N_10992,N_9718,N_9040);
nand U10993 (N_10993,N_9622,N_9489);
nand U10994 (N_10994,N_8927,N_9293);
nor U10995 (N_10995,N_9052,N_9142);
or U10996 (N_10996,N_9755,N_9154);
and U10997 (N_10997,N_9450,N_9595);
nand U10998 (N_10998,N_9136,N_8981);
xor U10999 (N_10999,N_9450,N_9411);
nand U11000 (N_11000,N_9165,N_9952);
xor U11001 (N_11001,N_9773,N_9120);
and U11002 (N_11002,N_9079,N_9438);
nand U11003 (N_11003,N_9285,N_9907);
nand U11004 (N_11004,N_9431,N_9495);
nor U11005 (N_11005,N_9372,N_9364);
and U11006 (N_11006,N_9587,N_9948);
nor U11007 (N_11007,N_9047,N_9799);
and U11008 (N_11008,N_9889,N_8983);
xor U11009 (N_11009,N_9175,N_9471);
xnor U11010 (N_11010,N_9046,N_9252);
nand U11011 (N_11011,N_9270,N_9529);
xor U11012 (N_11012,N_9875,N_9222);
or U11013 (N_11013,N_9597,N_8986);
or U11014 (N_11014,N_9854,N_9380);
nand U11015 (N_11015,N_9080,N_8986);
and U11016 (N_11016,N_9224,N_9537);
xor U11017 (N_11017,N_8852,N_9837);
xor U11018 (N_11018,N_9185,N_8866);
nor U11019 (N_11019,N_9405,N_9125);
xor U11020 (N_11020,N_9542,N_9095);
nor U11021 (N_11021,N_9086,N_8857);
nor U11022 (N_11022,N_9828,N_9887);
or U11023 (N_11023,N_8879,N_9016);
nand U11024 (N_11024,N_8757,N_9308);
nor U11025 (N_11025,N_9242,N_9138);
nor U11026 (N_11026,N_8936,N_9719);
nand U11027 (N_11027,N_8751,N_9313);
nand U11028 (N_11028,N_9487,N_9425);
xor U11029 (N_11029,N_8896,N_9346);
nor U11030 (N_11030,N_9906,N_8880);
nor U11031 (N_11031,N_9787,N_9475);
and U11032 (N_11032,N_9541,N_8977);
xor U11033 (N_11033,N_9006,N_9618);
nand U11034 (N_11034,N_9978,N_9319);
xor U11035 (N_11035,N_9596,N_9428);
nor U11036 (N_11036,N_9231,N_9161);
xor U11037 (N_11037,N_9863,N_8883);
nand U11038 (N_11038,N_8973,N_9404);
and U11039 (N_11039,N_9984,N_8775);
nor U11040 (N_11040,N_9742,N_9767);
and U11041 (N_11041,N_9820,N_9660);
nand U11042 (N_11042,N_9705,N_8883);
nor U11043 (N_11043,N_9439,N_9581);
or U11044 (N_11044,N_9861,N_9653);
nor U11045 (N_11045,N_9056,N_9871);
nand U11046 (N_11046,N_9299,N_9473);
nand U11047 (N_11047,N_9049,N_8781);
nand U11048 (N_11048,N_9846,N_9655);
nor U11049 (N_11049,N_9951,N_9460);
xor U11050 (N_11050,N_9844,N_9655);
nor U11051 (N_11051,N_9559,N_8800);
nor U11052 (N_11052,N_9627,N_9915);
nand U11053 (N_11053,N_8764,N_9528);
nand U11054 (N_11054,N_9853,N_9789);
xnor U11055 (N_11055,N_9778,N_9854);
nand U11056 (N_11056,N_9401,N_9379);
and U11057 (N_11057,N_8858,N_9333);
nor U11058 (N_11058,N_8945,N_9200);
and U11059 (N_11059,N_9516,N_9913);
and U11060 (N_11060,N_8824,N_9343);
nor U11061 (N_11061,N_9208,N_9484);
or U11062 (N_11062,N_8990,N_9433);
xnor U11063 (N_11063,N_9277,N_8902);
xnor U11064 (N_11064,N_8832,N_8778);
nand U11065 (N_11065,N_9721,N_9539);
nor U11066 (N_11066,N_9527,N_9627);
and U11067 (N_11067,N_9246,N_9715);
or U11068 (N_11068,N_9167,N_9593);
xor U11069 (N_11069,N_8840,N_9053);
nand U11070 (N_11070,N_9929,N_9370);
xor U11071 (N_11071,N_9581,N_9777);
xnor U11072 (N_11072,N_8829,N_9589);
nand U11073 (N_11073,N_9870,N_9926);
and U11074 (N_11074,N_9679,N_9476);
xor U11075 (N_11075,N_8868,N_9080);
nand U11076 (N_11076,N_9116,N_9390);
and U11077 (N_11077,N_9507,N_9811);
and U11078 (N_11078,N_9273,N_9412);
and U11079 (N_11079,N_9216,N_9595);
nor U11080 (N_11080,N_9046,N_9826);
nand U11081 (N_11081,N_9332,N_9011);
xor U11082 (N_11082,N_9062,N_8905);
xnor U11083 (N_11083,N_9517,N_9455);
nor U11084 (N_11084,N_9559,N_9413);
and U11085 (N_11085,N_9080,N_9370);
and U11086 (N_11086,N_9989,N_9610);
nor U11087 (N_11087,N_8818,N_9146);
or U11088 (N_11088,N_8860,N_9675);
nor U11089 (N_11089,N_9412,N_9186);
nand U11090 (N_11090,N_8798,N_8784);
xor U11091 (N_11091,N_9398,N_9354);
and U11092 (N_11092,N_9528,N_9625);
or U11093 (N_11093,N_9585,N_9164);
or U11094 (N_11094,N_9879,N_9317);
nand U11095 (N_11095,N_9551,N_9803);
nand U11096 (N_11096,N_8786,N_8798);
or U11097 (N_11097,N_9143,N_9019);
xnor U11098 (N_11098,N_9361,N_9176);
nor U11099 (N_11099,N_9697,N_9028);
and U11100 (N_11100,N_9950,N_9893);
or U11101 (N_11101,N_9364,N_9385);
nor U11102 (N_11102,N_8833,N_8968);
nand U11103 (N_11103,N_9833,N_8762);
nor U11104 (N_11104,N_9547,N_9098);
or U11105 (N_11105,N_9988,N_9498);
or U11106 (N_11106,N_8811,N_9274);
nor U11107 (N_11107,N_9333,N_8783);
nor U11108 (N_11108,N_9257,N_9640);
nor U11109 (N_11109,N_9865,N_9241);
and U11110 (N_11110,N_9665,N_9563);
nor U11111 (N_11111,N_9701,N_9358);
and U11112 (N_11112,N_9682,N_9865);
xnor U11113 (N_11113,N_8999,N_9301);
and U11114 (N_11114,N_9517,N_9274);
xnor U11115 (N_11115,N_8926,N_9945);
nor U11116 (N_11116,N_9150,N_9993);
nor U11117 (N_11117,N_9643,N_9388);
xnor U11118 (N_11118,N_8973,N_9649);
or U11119 (N_11119,N_9452,N_8977);
xor U11120 (N_11120,N_9808,N_9257);
and U11121 (N_11121,N_9732,N_8808);
or U11122 (N_11122,N_9330,N_9933);
and U11123 (N_11123,N_9095,N_9416);
xor U11124 (N_11124,N_8898,N_9473);
nand U11125 (N_11125,N_9466,N_9323);
or U11126 (N_11126,N_9958,N_9174);
and U11127 (N_11127,N_9799,N_8784);
xnor U11128 (N_11128,N_9369,N_9139);
or U11129 (N_11129,N_8914,N_8810);
nor U11130 (N_11130,N_8912,N_9404);
nand U11131 (N_11131,N_9738,N_9146);
and U11132 (N_11132,N_8894,N_9304);
xnor U11133 (N_11133,N_9861,N_9303);
nand U11134 (N_11134,N_9718,N_9136);
nand U11135 (N_11135,N_8900,N_9581);
nor U11136 (N_11136,N_9187,N_9668);
and U11137 (N_11137,N_9594,N_9757);
and U11138 (N_11138,N_9921,N_9336);
xor U11139 (N_11139,N_9622,N_9741);
nor U11140 (N_11140,N_9896,N_9278);
or U11141 (N_11141,N_9939,N_8981);
xor U11142 (N_11142,N_9995,N_9771);
xnor U11143 (N_11143,N_9731,N_9092);
xnor U11144 (N_11144,N_9662,N_9616);
xnor U11145 (N_11145,N_9721,N_9923);
nor U11146 (N_11146,N_9526,N_8907);
nand U11147 (N_11147,N_8885,N_9522);
xor U11148 (N_11148,N_9039,N_9172);
nor U11149 (N_11149,N_9758,N_9662);
xnor U11150 (N_11150,N_9040,N_9901);
and U11151 (N_11151,N_9154,N_9168);
xnor U11152 (N_11152,N_8945,N_9241);
xor U11153 (N_11153,N_9611,N_9898);
xor U11154 (N_11154,N_9199,N_8878);
or U11155 (N_11155,N_9608,N_8820);
nor U11156 (N_11156,N_9793,N_9844);
and U11157 (N_11157,N_8924,N_9543);
nor U11158 (N_11158,N_8781,N_9574);
nand U11159 (N_11159,N_9930,N_9433);
or U11160 (N_11160,N_9916,N_9151);
or U11161 (N_11161,N_9432,N_9005);
nand U11162 (N_11162,N_8779,N_9556);
or U11163 (N_11163,N_9349,N_8760);
nor U11164 (N_11164,N_9394,N_9190);
or U11165 (N_11165,N_9561,N_9188);
xnor U11166 (N_11166,N_9272,N_9185);
nand U11167 (N_11167,N_9563,N_9480);
nor U11168 (N_11168,N_9867,N_9415);
and U11169 (N_11169,N_9270,N_9513);
and U11170 (N_11170,N_9324,N_9858);
nor U11171 (N_11171,N_9770,N_9947);
or U11172 (N_11172,N_9659,N_9786);
nand U11173 (N_11173,N_9664,N_9710);
and U11174 (N_11174,N_9228,N_9115);
nand U11175 (N_11175,N_9926,N_9660);
nand U11176 (N_11176,N_9513,N_9782);
nor U11177 (N_11177,N_9219,N_8875);
nor U11178 (N_11178,N_9689,N_9732);
and U11179 (N_11179,N_9028,N_9823);
or U11180 (N_11180,N_9732,N_9853);
nor U11181 (N_11181,N_8950,N_9903);
nand U11182 (N_11182,N_9809,N_8753);
nor U11183 (N_11183,N_9265,N_9010);
and U11184 (N_11184,N_9111,N_9451);
or U11185 (N_11185,N_8830,N_9266);
and U11186 (N_11186,N_9184,N_9250);
and U11187 (N_11187,N_8750,N_9054);
nand U11188 (N_11188,N_9040,N_9309);
and U11189 (N_11189,N_8880,N_9190);
nor U11190 (N_11190,N_8866,N_8930);
and U11191 (N_11191,N_8859,N_9204);
nor U11192 (N_11192,N_9845,N_9815);
nor U11193 (N_11193,N_9571,N_9988);
or U11194 (N_11194,N_9494,N_9522);
nor U11195 (N_11195,N_9531,N_8943);
xor U11196 (N_11196,N_9844,N_9001);
or U11197 (N_11197,N_9058,N_9175);
nand U11198 (N_11198,N_9667,N_8785);
nor U11199 (N_11199,N_9992,N_9624);
and U11200 (N_11200,N_9299,N_8824);
nand U11201 (N_11201,N_9919,N_9884);
nand U11202 (N_11202,N_9782,N_9687);
and U11203 (N_11203,N_9416,N_9805);
nor U11204 (N_11204,N_9278,N_9184);
and U11205 (N_11205,N_9095,N_9541);
or U11206 (N_11206,N_9567,N_9097);
nand U11207 (N_11207,N_8902,N_8839);
and U11208 (N_11208,N_8927,N_8836);
and U11209 (N_11209,N_9042,N_9872);
and U11210 (N_11210,N_8891,N_9137);
or U11211 (N_11211,N_9042,N_9702);
or U11212 (N_11212,N_8929,N_9596);
or U11213 (N_11213,N_9651,N_9421);
nor U11214 (N_11214,N_9222,N_8943);
nand U11215 (N_11215,N_9148,N_9707);
xnor U11216 (N_11216,N_9907,N_9013);
and U11217 (N_11217,N_8869,N_9133);
nand U11218 (N_11218,N_9316,N_9409);
and U11219 (N_11219,N_9191,N_9839);
nand U11220 (N_11220,N_9732,N_9671);
nor U11221 (N_11221,N_8939,N_9130);
and U11222 (N_11222,N_9486,N_9288);
xnor U11223 (N_11223,N_9533,N_8764);
and U11224 (N_11224,N_9050,N_9110);
or U11225 (N_11225,N_9169,N_9804);
or U11226 (N_11226,N_9691,N_8990);
nand U11227 (N_11227,N_8983,N_9683);
xor U11228 (N_11228,N_9385,N_9883);
xnor U11229 (N_11229,N_9931,N_9412);
nor U11230 (N_11230,N_8879,N_9312);
and U11231 (N_11231,N_9433,N_8902);
or U11232 (N_11232,N_8803,N_9461);
nand U11233 (N_11233,N_9898,N_9137);
or U11234 (N_11234,N_9028,N_9328);
or U11235 (N_11235,N_9206,N_9957);
nor U11236 (N_11236,N_8828,N_9948);
and U11237 (N_11237,N_9996,N_9271);
nor U11238 (N_11238,N_9313,N_9832);
nor U11239 (N_11239,N_9998,N_9118);
nor U11240 (N_11240,N_9647,N_8771);
and U11241 (N_11241,N_9544,N_9580);
or U11242 (N_11242,N_8857,N_9401);
and U11243 (N_11243,N_8767,N_9727);
xnor U11244 (N_11244,N_9302,N_9198);
and U11245 (N_11245,N_9809,N_9576);
or U11246 (N_11246,N_8996,N_9821);
or U11247 (N_11247,N_9649,N_8883);
or U11248 (N_11248,N_9216,N_9459);
nand U11249 (N_11249,N_9858,N_9332);
and U11250 (N_11250,N_11152,N_11081);
xnor U11251 (N_11251,N_10676,N_10851);
nor U11252 (N_11252,N_10808,N_10014);
and U11253 (N_11253,N_10771,N_10210);
nor U11254 (N_11254,N_11164,N_10393);
xnor U11255 (N_11255,N_11167,N_10553);
nand U11256 (N_11256,N_10708,N_10333);
and U11257 (N_11257,N_10248,N_10743);
nand U11258 (N_11258,N_10954,N_10143);
nand U11259 (N_11259,N_10192,N_11168);
nand U11260 (N_11260,N_11248,N_10421);
or U11261 (N_11261,N_10949,N_10088);
and U11262 (N_11262,N_10985,N_10779);
nand U11263 (N_11263,N_10660,N_10468);
nand U11264 (N_11264,N_11169,N_10629);
nor U11265 (N_11265,N_10993,N_10725);
nand U11266 (N_11266,N_10291,N_10238);
xor U11267 (N_11267,N_10580,N_10346);
or U11268 (N_11268,N_10140,N_10908);
and U11269 (N_11269,N_10811,N_10089);
and U11270 (N_11270,N_10073,N_10072);
xnor U11271 (N_11271,N_10788,N_10319);
nor U11272 (N_11272,N_10146,N_10994);
nand U11273 (N_11273,N_11021,N_10299);
and U11274 (N_11274,N_10723,N_10241);
nor U11275 (N_11275,N_11176,N_10847);
xnor U11276 (N_11276,N_10763,N_10338);
nand U11277 (N_11277,N_10481,N_10835);
and U11278 (N_11278,N_10643,N_10613);
nor U11279 (N_11279,N_10050,N_11231);
and U11280 (N_11280,N_10976,N_10106);
or U11281 (N_11281,N_10820,N_11118);
xor U11282 (N_11282,N_10011,N_10315);
xor U11283 (N_11283,N_10021,N_10699);
and U11284 (N_11284,N_10928,N_10173);
and U11285 (N_11285,N_10899,N_10194);
and U11286 (N_11286,N_10901,N_11063);
xor U11287 (N_11287,N_10437,N_10774);
nor U11288 (N_11288,N_10591,N_10681);
nor U11289 (N_11289,N_10412,N_10433);
or U11290 (N_11290,N_10170,N_10995);
nand U11291 (N_11291,N_10893,N_11001);
nand U11292 (N_11292,N_11095,N_11181);
nand U11293 (N_11293,N_10962,N_10652);
nand U11294 (N_11294,N_11247,N_10076);
xnor U11295 (N_11295,N_11124,N_10110);
and U11296 (N_11296,N_10565,N_10280);
nand U11297 (N_11297,N_10324,N_10450);
nand U11298 (N_11298,N_10493,N_10448);
and U11299 (N_11299,N_11173,N_11024);
nor U11300 (N_11300,N_10294,N_10748);
nand U11301 (N_11301,N_11237,N_11204);
or U11302 (N_11302,N_10312,N_10602);
or U11303 (N_11303,N_10509,N_10415);
nand U11304 (N_11304,N_10929,N_10256);
or U11305 (N_11305,N_10358,N_10517);
xor U11306 (N_11306,N_11080,N_10859);
nand U11307 (N_11307,N_11184,N_10869);
xnor U11308 (N_11308,N_11189,N_10527);
nand U11309 (N_11309,N_10706,N_10092);
xnor U11310 (N_11310,N_11244,N_10977);
or U11311 (N_11311,N_10815,N_10288);
or U11312 (N_11312,N_10220,N_10270);
or U11313 (N_11313,N_10939,N_11135);
xor U11314 (N_11314,N_10844,N_11030);
or U11315 (N_11315,N_11075,N_10673);
nor U11316 (N_11316,N_10239,N_10531);
xor U11317 (N_11317,N_10840,N_10176);
and U11318 (N_11318,N_10165,N_10009);
nand U11319 (N_11319,N_10938,N_10352);
nor U11320 (N_11320,N_10520,N_10368);
or U11321 (N_11321,N_10654,N_10547);
nor U11322 (N_11322,N_10378,N_10127);
xnor U11323 (N_11323,N_11051,N_10417);
nand U11324 (N_11324,N_11134,N_10419);
nand U11325 (N_11325,N_11241,N_10558);
xnor U11326 (N_11326,N_10218,N_10955);
or U11327 (N_11327,N_10258,N_10398);
nand U11328 (N_11328,N_10698,N_10310);
xnor U11329 (N_11329,N_10486,N_10455);
nor U11330 (N_11330,N_10060,N_10704);
and U11331 (N_11331,N_10484,N_10186);
xnor U11332 (N_11332,N_10584,N_10661);
and U11333 (N_11333,N_10967,N_10171);
nor U11334 (N_11334,N_10594,N_10752);
nor U11335 (N_11335,N_10714,N_11038);
nor U11336 (N_11336,N_10142,N_10878);
and U11337 (N_11337,N_11214,N_11066);
or U11338 (N_11338,N_10101,N_10790);
xnor U11339 (N_11339,N_10645,N_10814);
nor U11340 (N_11340,N_10330,N_10999);
nor U11341 (N_11341,N_11086,N_10151);
nand U11342 (N_11342,N_10983,N_10154);
and U11343 (N_11343,N_10927,N_11067);
xor U11344 (N_11344,N_10045,N_11005);
or U11345 (N_11345,N_10665,N_10215);
xor U11346 (N_11346,N_10858,N_10795);
nor U11347 (N_11347,N_11175,N_10839);
nand U11348 (N_11348,N_11212,N_10772);
nor U11349 (N_11349,N_10970,N_10617);
nor U11350 (N_11350,N_10742,N_10329);
and U11351 (N_11351,N_11076,N_10314);
or U11352 (N_11352,N_10592,N_10933);
nand U11353 (N_11353,N_10284,N_11070);
nor U11354 (N_11354,N_10129,N_10502);
nor U11355 (N_11355,N_10898,N_10668);
nor U11356 (N_11356,N_11120,N_11226);
and U11357 (N_11357,N_11018,N_10737);
and U11358 (N_11358,N_10349,N_11060);
xnor U11359 (N_11359,N_11009,N_11194);
nand U11360 (N_11360,N_10651,N_10888);
or U11361 (N_11361,N_11222,N_11172);
or U11362 (N_11362,N_10769,N_10169);
nand U11363 (N_11363,N_10867,N_10936);
or U11364 (N_11364,N_10785,N_10778);
and U11365 (N_11365,N_10264,N_10371);
nor U11366 (N_11366,N_10025,N_10286);
or U11367 (N_11367,N_10459,N_10124);
or U11368 (N_11368,N_10749,N_10897);
nand U11369 (N_11369,N_10189,N_10307);
xor U11370 (N_11370,N_10255,N_10724);
nor U11371 (N_11371,N_11129,N_10242);
xnor U11372 (N_11372,N_11242,N_10487);
nor U11373 (N_11373,N_11149,N_10671);
nor U11374 (N_11374,N_10640,N_11042);
or U11375 (N_11375,N_10287,N_10340);
nor U11376 (N_11376,N_10806,N_10235);
or U11377 (N_11377,N_10108,N_10951);
nand U11378 (N_11378,N_10079,N_10276);
nor U11379 (N_11379,N_10357,N_10107);
nand U11380 (N_11380,N_10544,N_10700);
nor U11381 (N_11381,N_10707,N_10818);
nor U11382 (N_11382,N_10712,N_10537);
and U11383 (N_11383,N_10722,N_10731);
nor U11384 (N_11384,N_10744,N_10870);
or U11385 (N_11385,N_10925,N_10168);
xnor U11386 (N_11386,N_10006,N_10667);
nor U11387 (N_11387,N_10332,N_11065);
or U11388 (N_11388,N_10426,N_10013);
and U11389 (N_11389,N_10262,N_10507);
nor U11390 (N_11390,N_10004,N_10562);
nand U11391 (N_11391,N_10805,N_10965);
nand U11392 (N_11392,N_10990,N_10822);
and U11393 (N_11393,N_10445,N_10508);
and U11394 (N_11394,N_11232,N_10285);
nand U11395 (N_11395,N_10497,N_10492);
nand U11396 (N_11396,N_10656,N_11137);
and U11397 (N_11397,N_10064,N_10826);
or U11398 (N_11398,N_10988,N_10595);
nor U11399 (N_11399,N_10540,N_10225);
nand U11400 (N_11400,N_10891,N_10546);
nor U11401 (N_11401,N_10259,N_10410);
nor U11402 (N_11402,N_10794,N_10126);
or U11403 (N_11403,N_10213,N_10669);
or U11404 (N_11404,N_11207,N_10601);
or U11405 (N_11405,N_10650,N_11049);
and U11406 (N_11406,N_10098,N_11087);
nand U11407 (N_11407,N_10701,N_10234);
nor U11408 (N_11408,N_10810,N_11015);
and U11409 (N_11409,N_10857,N_10968);
nand U11410 (N_11410,N_10401,N_10369);
nand U11411 (N_11411,N_10477,N_10399);
nand U11412 (N_11412,N_10561,N_10281);
and U11413 (N_11413,N_10906,N_10720);
nor U11414 (N_11414,N_11126,N_10780);
or U11415 (N_11415,N_10217,N_11190);
nand U11416 (N_11416,N_10001,N_10411);
and U11417 (N_11417,N_10155,N_11121);
nor U11418 (N_11418,N_11078,N_10766);
and U11419 (N_11419,N_11141,N_10265);
xor U11420 (N_11420,N_10512,N_11163);
xnor U11421 (N_11421,N_10717,N_10366);
xor U11422 (N_11422,N_10874,N_10231);
nand U11423 (N_11423,N_10078,N_10420);
xnor U11424 (N_11424,N_10776,N_10121);
nand U11425 (N_11425,N_10042,N_10000);
and U11426 (N_11426,N_10372,N_10488);
or U11427 (N_11427,N_10343,N_10458);
nand U11428 (N_11428,N_10958,N_10306);
nand U11429 (N_11429,N_10905,N_11031);
nor U11430 (N_11430,N_11174,N_10646);
or U11431 (N_11431,N_10666,N_10441);
nand U11432 (N_11432,N_10359,N_10439);
nor U11433 (N_11433,N_10379,N_10081);
and U11434 (N_11434,N_10581,N_10430);
nand U11435 (N_11435,N_11085,N_10289);
xor U11436 (N_11436,N_10798,N_10728);
xor U11437 (N_11437,N_10395,N_10047);
nand U11438 (N_11438,N_10103,N_10160);
nor U11439 (N_11439,N_11155,N_10523);
nand U11440 (N_11440,N_10606,N_10133);
xor U11441 (N_11441,N_10871,N_11227);
xnor U11442 (N_11442,N_10158,N_10387);
xnor U11443 (N_11443,N_11220,N_10917);
nand U11444 (N_11444,N_10185,N_11089);
nor U11445 (N_11445,N_10283,N_10515);
or U11446 (N_11446,N_10940,N_11161);
nor U11447 (N_11447,N_10896,N_10038);
nor U11448 (N_11448,N_10318,N_10052);
and U11449 (N_11449,N_10396,N_11157);
or U11450 (N_11450,N_10416,N_10273);
xnor U11451 (N_11451,N_10322,N_11041);
and U11452 (N_11452,N_10603,N_10061);
xnor U11453 (N_11453,N_11040,N_10691);
or U11454 (N_11454,N_10726,N_11111);
or U11455 (N_11455,N_10162,N_10791);
nand U11456 (N_11456,N_10068,N_10446);
nand U11457 (N_11457,N_10653,N_10271);
nor U11458 (N_11458,N_10695,N_11127);
xnor U11459 (N_11459,N_10243,N_10353);
or U11460 (N_11460,N_10658,N_10913);
and U11461 (N_11461,N_11073,N_10015);
nand U11462 (N_11462,N_11029,N_11002);
nand U11463 (N_11463,N_10555,N_10336);
nor U11464 (N_11464,N_10033,N_10586);
or U11465 (N_11465,N_10834,N_10112);
nand U11466 (N_11466,N_10381,N_11192);
xor U11467 (N_11467,N_10620,N_10755);
nor U11468 (N_11468,N_10926,N_10188);
nand U11469 (N_11469,N_10263,N_10086);
and U11470 (N_11470,N_10600,N_11069);
and U11471 (N_11471,N_10037,N_10556);
nor U11472 (N_11472,N_11160,N_11224);
and U11473 (N_11473,N_10282,N_10018);
nand U11474 (N_11474,N_10132,N_10644);
nand U11475 (N_11475,N_10915,N_10010);
nand U11476 (N_11476,N_10482,N_11228);
xor U11477 (N_11477,N_10510,N_11195);
or U11478 (N_11478,N_10466,N_10224);
xnor U11479 (N_11479,N_10662,N_11088);
and U11480 (N_11480,N_11000,N_10753);
or U11481 (N_11481,N_10607,N_10959);
nand U11482 (N_11482,N_10403,N_10104);
or U11483 (N_11483,N_11217,N_11147);
or U11484 (N_11484,N_10384,N_10309);
xnor U11485 (N_11485,N_10566,N_10963);
nand U11486 (N_11486,N_10885,N_10924);
nand U11487 (N_11487,N_10732,N_10229);
or U11488 (N_11488,N_11077,N_10094);
nand U11489 (N_11489,N_10449,N_10007);
nand U11490 (N_11490,N_10848,N_10118);
xor U11491 (N_11491,N_10111,N_10842);
nand U11492 (N_11492,N_10588,N_11183);
xnor U11493 (N_11493,N_10240,N_10342);
xnor U11494 (N_11494,N_10424,N_10552);
nand U11495 (N_11495,N_10300,N_11140);
or U11496 (N_11496,N_10219,N_10392);
xnor U11497 (N_11497,N_10051,N_11218);
or U11498 (N_11498,N_10303,N_10892);
nor U11499 (N_11499,N_10113,N_10305);
or U11500 (N_11500,N_10120,N_10746);
nor U11501 (N_11501,N_11008,N_10245);
nor U11502 (N_11502,N_10494,N_11110);
or U11503 (N_11503,N_10616,N_10721);
or U11504 (N_11504,N_10861,N_10438);
and U11505 (N_11505,N_10505,N_10180);
xor U11506 (N_11506,N_11210,N_10767);
or U11507 (N_11507,N_11216,N_10803);
nor U11508 (N_11508,N_10831,N_10406);
and U11509 (N_11509,N_10465,N_10096);
xnor U11510 (N_11510,N_10855,N_10944);
and U11511 (N_11511,N_10860,N_10907);
xor U11512 (N_11512,N_11205,N_10634);
xnor U11513 (N_11513,N_11145,N_10733);
and U11514 (N_11514,N_10498,N_11092);
nand U11515 (N_11515,N_10461,N_10930);
xnor U11516 (N_11516,N_10157,N_11128);
nand U11517 (N_11517,N_11072,N_10257);
nand U11518 (N_11518,N_11170,N_10541);
and U11519 (N_11519,N_10719,N_10872);
or U11520 (N_11520,N_10850,N_10134);
nor U11521 (N_11521,N_10941,N_10741);
nand U11522 (N_11522,N_10577,N_10102);
xnor U11523 (N_11523,N_11234,N_10682);
and U11524 (N_11524,N_11019,N_10711);
nor U11525 (N_11525,N_10277,N_11206);
nor U11526 (N_11526,N_10760,N_11125);
nor U11527 (N_11527,N_10130,N_10123);
and U11528 (N_11528,N_10386,N_10469);
xor U11529 (N_11529,N_10063,N_10216);
or U11530 (N_11530,N_11177,N_10054);
nor U11531 (N_11531,N_10783,N_10604);
xor U11532 (N_11532,N_10932,N_10879);
or U11533 (N_11533,N_10181,N_11054);
and U11534 (N_11534,N_10948,N_10796);
xnor U11535 (N_11535,N_10172,N_10389);
or U11536 (N_11536,N_10764,N_10442);
nor U11537 (N_11537,N_10316,N_10873);
or U11538 (N_11538,N_11166,N_10008);
nand U11539 (N_11539,N_10191,N_10039);
and U11540 (N_11540,N_10572,N_10308);
and U11541 (N_11541,N_10119,N_10302);
and U11542 (N_11542,N_10223,N_10297);
and U11543 (N_11543,N_11162,N_10201);
nor U11544 (N_11544,N_10718,N_10407);
and U11545 (N_11545,N_10383,N_10095);
nand U11546 (N_11546,N_10207,N_11182);
or U11547 (N_11547,N_10163,N_10524);
and U11548 (N_11548,N_10986,N_10511);
nor U11549 (N_11549,N_10193,N_11199);
nor U11550 (N_11550,N_11074,N_10237);
and U11551 (N_11551,N_11055,N_10589);
and U11552 (N_11552,N_10034,N_10647);
nor U11553 (N_11553,N_10997,N_10462);
and U11554 (N_11554,N_10829,N_10066);
and U11555 (N_11555,N_10451,N_11119);
xor U11556 (N_11556,N_11006,N_11208);
and U11557 (N_11557,N_10418,N_10131);
nor U11558 (N_11558,N_10206,N_10161);
nand U11559 (N_11559,N_10067,N_10841);
nor U11560 (N_11560,N_10910,N_10020);
or U11561 (N_11561,N_10423,N_10044);
and U11562 (N_11562,N_10882,N_11079);
or U11563 (N_11563,N_10320,N_11056);
nand U11564 (N_11564,N_10866,N_10895);
or U11565 (N_11565,N_10296,N_11003);
or U11566 (N_11566,N_10745,N_10619);
nor U11567 (N_11567,N_11053,N_11082);
nand U11568 (N_11568,N_10563,N_10812);
or U11569 (N_11569,N_10659,N_10799);
xor U11570 (N_11570,N_10894,N_11219);
nor U11571 (N_11571,N_10470,N_10272);
nor U11572 (N_11572,N_11059,N_10480);
nand U11573 (N_11573,N_10648,N_11093);
or U11574 (N_11574,N_10684,N_10250);
xnor U11575 (N_11575,N_10655,N_11123);
or U11576 (N_11576,N_10221,N_10705);
xor U11577 (N_11577,N_11198,N_10397);
xor U11578 (N_11578,N_10304,N_10813);
nor U11579 (N_11579,N_10491,N_10686);
nor U11580 (N_11580,N_11058,N_10058);
nor U11581 (N_11581,N_10890,N_10128);
or U11582 (N_11582,N_10618,N_10109);
or U11583 (N_11583,N_10327,N_11039);
and U11584 (N_11584,N_10090,N_10085);
and U11585 (N_11585,N_10902,N_10184);
and U11586 (N_11586,N_11035,N_10543);
nand U11587 (N_11587,N_10364,N_11114);
xor U11588 (N_11588,N_10382,N_10518);
nand U11589 (N_11589,N_10317,N_10784);
xor U11590 (N_11590,N_10614,N_10087);
nor U11591 (N_11591,N_10341,N_10542);
xor U11592 (N_11592,N_10175,N_11099);
nor U11593 (N_11593,N_10950,N_10361);
nor U11594 (N_11594,N_11165,N_10845);
nand U11595 (N_11595,N_10116,N_10135);
or U11596 (N_11596,N_10056,N_10198);
xor U11597 (N_11597,N_10226,N_10694);
nor U11598 (N_11598,N_10919,N_10961);
or U11599 (N_11599,N_10138,N_10496);
xnor U11600 (N_11600,N_11196,N_10624);
xnor U11601 (N_11601,N_10070,N_11235);
nand U11602 (N_11602,N_11185,N_10059);
or U11603 (N_11603,N_11156,N_10208);
and U11604 (N_11604,N_10570,N_10920);
and U11605 (N_11605,N_10447,N_10122);
nor U11606 (N_11606,N_11071,N_10884);
xor U11607 (N_11607,N_10865,N_10177);
xnor U11608 (N_11608,N_11037,N_10828);
nor U11609 (N_11609,N_10476,N_11193);
xnor U11610 (N_11610,N_11096,N_10922);
xnor U11611 (N_11611,N_11007,N_11201);
nor U11612 (N_11612,N_10337,N_10199);
nor U11613 (N_11613,N_10973,N_10539);
nor U11614 (N_11614,N_10754,N_10362);
nor U11615 (N_11615,N_10495,N_10639);
xor U11616 (N_11616,N_10472,N_10689);
nand U11617 (N_11617,N_10145,N_10679);
nor U11618 (N_11618,N_10290,N_10918);
and U11619 (N_11619,N_10750,N_10937);
and U11620 (N_11620,N_11109,N_10084);
xor U11621 (N_11621,N_10522,N_10598);
xor U11622 (N_11622,N_11188,N_10996);
or U11623 (N_11623,N_10267,N_10587);
and U11624 (N_11624,N_10335,N_10149);
or U11625 (N_11625,N_10621,N_10373);
nand U11626 (N_11626,N_10786,N_10880);
and U11627 (N_11627,N_11221,N_10457);
xor U11628 (N_11628,N_10503,N_11133);
or U11629 (N_11629,N_10852,N_10478);
or U11630 (N_11630,N_10675,N_10251);
nor U11631 (N_11631,N_10992,N_11249);
or U11632 (N_11632,N_10431,N_10887);
nor U11633 (N_11633,N_10574,N_10463);
and U11634 (N_11634,N_10610,N_10348);
and U11635 (N_11635,N_10022,N_10809);
xor U11636 (N_11636,N_10914,N_10713);
nand U11637 (N_11637,N_10232,N_10295);
xnor U11638 (N_11638,N_10971,N_10942);
nand U11639 (N_11639,N_10560,N_11211);
xor U11640 (N_11640,N_10388,N_10200);
nand U11641 (N_11641,N_10824,N_10615);
nand U11642 (N_11642,N_10853,N_11012);
and U11643 (N_11643,N_11105,N_10196);
and U11644 (N_11644,N_10576,N_11171);
or U11645 (N_11645,N_11014,N_10554);
and U11646 (N_11646,N_11179,N_11068);
nand U11647 (N_11647,N_10029,N_11036);
or U11648 (N_11648,N_10363,N_10693);
or U11649 (N_11649,N_10244,N_11143);
or U11650 (N_11650,N_10978,N_10298);
nand U11651 (N_11651,N_10460,N_11240);
nor U11652 (N_11652,N_10053,N_10247);
xor U11653 (N_11653,N_10947,N_10800);
and U11654 (N_11654,N_10156,N_10627);
nor U11655 (N_11655,N_10205,N_10773);
xnor U11656 (N_11656,N_10099,N_10252);
or U11657 (N_11657,N_10432,N_10819);
nand U11658 (N_11658,N_10150,N_10385);
and U11659 (N_11659,N_11028,N_10982);
nor U11660 (N_11660,N_10048,N_10670);
xor U11661 (N_11661,N_10514,N_11097);
and U11662 (N_11662,N_11187,N_11033);
xor U11663 (N_11663,N_10485,N_11104);
or U11664 (N_11664,N_10987,N_10139);
and U11665 (N_11665,N_10685,N_10641);
nor U11666 (N_11666,N_11025,N_11153);
nand U11667 (N_11667,N_10945,N_10233);
xnor U11668 (N_11668,N_10573,N_10253);
nand U11669 (N_11669,N_10854,N_10345);
and U11670 (N_11670,N_10881,N_10159);
nor U11671 (N_11671,N_10696,N_11102);
or U11672 (N_11672,N_10422,N_10757);
or U11673 (N_11673,N_10876,N_10952);
nand U11674 (N_11674,N_10026,N_10141);
and U11675 (N_11675,N_10115,N_10868);
nor U11676 (N_11676,N_10427,N_11113);
nand U11677 (N_11677,N_10916,N_10040);
and U11678 (N_11678,N_10579,N_10683);
and U11679 (N_11679,N_10152,N_10024);
and U11680 (N_11680,N_10727,N_10582);
and U11681 (N_11681,N_10091,N_10425);
nor U11682 (N_11682,N_11180,N_10016);
nand U11683 (N_11683,N_10956,N_11020);
nand U11684 (N_11684,N_10093,N_10729);
or U11685 (N_11685,N_10623,N_10414);
or U11686 (N_11686,N_10365,N_10549);
or U11687 (N_11687,N_10489,N_11103);
nor U11688 (N_11688,N_10227,N_11046);
and U11689 (N_11689,N_10404,N_10483);
nand U11690 (N_11690,N_10697,N_11047);
or U11691 (N_11691,N_10991,N_11061);
xnor U11692 (N_11692,N_10960,N_10912);
and U11693 (N_11693,N_10400,N_10946);
nand U11694 (N_11694,N_10585,N_10801);
nand U11695 (N_11695,N_10187,N_10921);
nor U11696 (N_11696,N_10453,N_10097);
and U11697 (N_11697,N_11215,N_10569);
xnor U11698 (N_11698,N_10370,N_10687);
nand U11699 (N_11699,N_10526,N_10551);
nor U11700 (N_11700,N_10246,N_10605);
xor U11701 (N_11701,N_10821,N_11050);
nand U11702 (N_11702,N_10049,N_10311);
nor U11703 (N_11703,N_10454,N_10532);
nor U11704 (N_11704,N_10355,N_11107);
xor U11705 (N_11705,N_10738,N_10534);
and U11706 (N_11706,N_10002,N_10292);
and U11707 (N_11707,N_10222,N_10394);
and U11708 (N_11708,N_10680,N_10428);
nor U11709 (N_11709,N_10409,N_10444);
xor U11710 (N_11710,N_10843,N_11200);
nor U11711 (N_11711,N_10323,N_10041);
nor U11712 (N_11712,N_10625,N_10083);
and U11713 (N_11713,N_10230,N_10777);
xnor U11714 (N_11714,N_10479,N_10817);
and U11715 (N_11715,N_10759,N_10536);
or U11716 (N_11716,N_11043,N_10190);
nand U11717 (N_11717,N_11225,N_10077);
nand U11718 (N_11718,N_10035,N_10443);
nor U11719 (N_11719,N_10023,N_10863);
nand U11720 (N_11720,N_11139,N_11203);
xor U11721 (N_11721,N_10195,N_10608);
nand U11722 (N_11722,N_10735,N_10166);
nand U11723 (N_11723,N_11026,N_10969);
and U11724 (N_11724,N_10374,N_10268);
and U11725 (N_11725,N_10762,N_10408);
or U11726 (N_11726,N_10183,N_10657);
or U11727 (N_11727,N_10182,N_11148);
nor U11728 (N_11728,N_11130,N_10269);
or U11729 (N_11729,N_10528,N_10931);
xnor U11730 (N_11730,N_11094,N_10301);
nor U11731 (N_11731,N_10350,N_10203);
nor U11732 (N_11732,N_10228,N_10214);
or U11733 (N_11733,N_10599,N_10525);
and U11734 (N_11734,N_11034,N_11083);
nor U11735 (N_11735,N_10197,N_11011);
and U11736 (N_11736,N_11243,N_11116);
or U11737 (N_11737,N_10593,N_10473);
or U11738 (N_11738,N_10003,N_10334);
and U11739 (N_11739,N_10031,N_10934);
and U11740 (N_11740,N_10635,N_10548);
and U11741 (N_11741,N_10575,N_10974);
nor U11742 (N_11742,N_10793,N_10328);
and U11743 (N_11743,N_11108,N_10792);
nor U11744 (N_11744,N_11004,N_10568);
or U11745 (N_11745,N_10027,N_11245);
nand U11746 (N_11746,N_10559,N_11136);
nor U11747 (N_11747,N_11186,N_10875);
or U11748 (N_11748,N_10849,N_10797);
and U11749 (N_11749,N_11223,N_11022);
nor U11750 (N_11750,N_10513,N_10664);
nor U11751 (N_11751,N_11131,N_10082);
nand U11752 (N_11752,N_10688,N_10434);
or U11753 (N_11753,N_10474,N_10405);
nand U11754 (N_11754,N_10475,N_10236);
nor U11755 (N_11755,N_10028,N_10730);
nor U11756 (N_11756,N_10979,N_10125);
and U11757 (N_11757,N_10578,N_10065);
nand U11758 (N_11758,N_10321,N_10981);
nor U11759 (N_11759,N_10464,N_10501);
xnor U11760 (N_11760,N_11013,N_10830);
xnor U11761 (N_11761,N_10611,N_10911);
or U11762 (N_11762,N_10703,N_10331);
nand U11763 (N_11763,N_10856,N_10943);
and U11764 (N_11764,N_10062,N_10765);
nor U11765 (N_11765,N_10758,N_10631);
or U11766 (N_11766,N_10538,N_10770);
nand U11767 (N_11767,N_10402,N_10690);
nand U11768 (N_11768,N_10375,N_10837);
and U11769 (N_11769,N_11010,N_10325);
nor U11770 (N_11770,N_10768,N_10204);
xor U11771 (N_11771,N_11158,N_10440);
and U11772 (N_11772,N_10521,N_10715);
or U11773 (N_11773,N_10360,N_11101);
and U11774 (N_11774,N_10756,N_10709);
nor U11775 (N_11775,N_10823,N_11146);
and U11776 (N_11776,N_10471,N_11213);
nand U11777 (N_11777,N_10339,N_10716);
or U11778 (N_11778,N_10075,N_10612);
nor U11779 (N_11779,N_10533,N_10490);
nand U11780 (N_11780,N_10909,N_10886);
nor U11781 (N_11781,N_10136,N_10266);
nor U11782 (N_11782,N_10274,N_10649);
nand U11783 (N_11783,N_10391,N_10692);
nor U11784 (N_11784,N_10825,N_10677);
and U11785 (N_11785,N_10043,N_10017);
or U11786 (N_11786,N_10144,N_10710);
nand U11787 (N_11787,N_11238,N_10260);
nor U11788 (N_11788,N_11144,N_11159);
and U11789 (N_11789,N_10903,N_10069);
nand U11790 (N_11790,N_10179,N_10816);
nand U11791 (N_11791,N_10019,N_10377);
or U11792 (N_11792,N_10499,N_10663);
nor U11793 (N_11793,N_10074,N_11191);
and U11794 (N_11794,N_10278,N_10998);
or U11795 (N_11795,N_10862,N_11044);
nor U11796 (N_11796,N_10628,N_10751);
xor U11797 (N_11797,N_10787,N_11016);
nor U11798 (N_11798,N_11122,N_10254);
and U11799 (N_11799,N_10500,N_10293);
xnor U11800 (N_11800,N_10080,N_10436);
and U11801 (N_11801,N_10836,N_10275);
nor U11802 (N_11802,N_11115,N_10636);
and U11803 (N_11803,N_10380,N_10279);
xnor U11804 (N_11804,N_11202,N_10005);
xor U11805 (N_11805,N_10564,N_10832);
and U11806 (N_11806,N_10736,N_10846);
xnor U11807 (N_11807,N_10597,N_10211);
and U11808 (N_11808,N_10529,N_10467);
xnor U11809 (N_11809,N_10590,N_11142);
nand U11810 (N_11810,N_11032,N_10775);
xor U11811 (N_11811,N_10148,N_10114);
nand U11812 (N_11812,N_10975,N_10747);
nor U11813 (N_11813,N_10889,N_10354);
nor U11814 (N_11814,N_10153,N_10036);
nand U11815 (N_11815,N_10838,N_10057);
and U11816 (N_11816,N_10071,N_11091);
nand U11817 (N_11817,N_10261,N_10557);
nand U11818 (N_11818,N_11084,N_10519);
xnor U11819 (N_11819,N_10782,N_10609);
xnor U11820 (N_11820,N_10164,N_10178);
nand U11821 (N_11821,N_10923,N_10100);
or U11822 (N_11822,N_11064,N_11154);
or U11823 (N_11823,N_10452,N_10877);
and U11824 (N_11824,N_10761,N_11239);
xor U11825 (N_11825,N_11017,N_10739);
or U11826 (N_11826,N_10633,N_10504);
xor U11827 (N_11827,N_10642,N_10953);
and U11828 (N_11828,N_10833,N_10734);
and U11829 (N_11829,N_10632,N_10802);
and U11830 (N_11830,N_11117,N_10137);
and U11831 (N_11831,N_10012,N_10347);
or U11832 (N_11832,N_10678,N_10030);
or U11833 (N_11833,N_10167,N_10957);
nor U11834 (N_11834,N_10550,N_10376);
or U11835 (N_11835,N_11106,N_11150);
and U11836 (N_11836,N_10638,N_10864);
and U11837 (N_11837,N_11057,N_10980);
nor U11838 (N_11838,N_10702,N_10571);
and U11839 (N_11839,N_10212,N_10596);
nand U11840 (N_11840,N_10105,N_10637);
nand U11841 (N_11841,N_10506,N_10966);
and U11842 (N_11842,N_11229,N_10516);
nand U11843 (N_11843,N_10390,N_10209);
nor U11844 (N_11844,N_10964,N_11098);
nor U11845 (N_11845,N_10989,N_11062);
nor U11846 (N_11846,N_11178,N_10984);
nand U11847 (N_11847,N_11197,N_10630);
nor U11848 (N_11848,N_10904,N_11233);
nor U11849 (N_11849,N_10147,N_10807);
xor U11850 (N_11850,N_10456,N_10530);
or U11851 (N_11851,N_10032,N_10055);
or U11852 (N_11852,N_10972,N_11045);
nand U11853 (N_11853,N_10202,N_10567);
and U11854 (N_11854,N_10827,N_11236);
xor U11855 (N_11855,N_10429,N_10356);
and U11856 (N_11856,N_10535,N_10883);
and U11857 (N_11857,N_11209,N_10435);
xnor U11858 (N_11858,N_10789,N_11230);
and U11859 (N_11859,N_10935,N_10351);
or U11860 (N_11860,N_11048,N_10672);
and U11861 (N_11861,N_10804,N_10545);
nor U11862 (N_11862,N_10249,N_10626);
xnor U11863 (N_11863,N_11100,N_10046);
nand U11864 (N_11864,N_10117,N_10326);
nand U11865 (N_11865,N_10367,N_11246);
xor U11866 (N_11866,N_11151,N_10674);
xnor U11867 (N_11867,N_11138,N_10344);
nor U11868 (N_11868,N_11112,N_10740);
and U11869 (N_11869,N_10174,N_10622);
or U11870 (N_11870,N_11027,N_11090);
nand U11871 (N_11871,N_10313,N_10583);
or U11872 (N_11872,N_11132,N_11052);
nand U11873 (N_11873,N_11023,N_10413);
xor U11874 (N_11874,N_10781,N_10900);
nand U11875 (N_11875,N_10267,N_10162);
or U11876 (N_11876,N_10558,N_11180);
or U11877 (N_11877,N_11202,N_10254);
and U11878 (N_11878,N_11007,N_10081);
or U11879 (N_11879,N_10870,N_10773);
nand U11880 (N_11880,N_10607,N_10237);
or U11881 (N_11881,N_10471,N_10801);
xor U11882 (N_11882,N_10809,N_10091);
xnor U11883 (N_11883,N_10286,N_10805);
nand U11884 (N_11884,N_11154,N_10457);
nand U11885 (N_11885,N_11069,N_10011);
xor U11886 (N_11886,N_10000,N_10933);
xnor U11887 (N_11887,N_10477,N_10694);
and U11888 (N_11888,N_10613,N_10212);
and U11889 (N_11889,N_10473,N_10154);
and U11890 (N_11890,N_10386,N_10810);
or U11891 (N_11891,N_10417,N_10997);
and U11892 (N_11892,N_11245,N_10985);
nand U11893 (N_11893,N_10660,N_10709);
or U11894 (N_11894,N_10904,N_10592);
and U11895 (N_11895,N_10586,N_10081);
or U11896 (N_11896,N_10558,N_10269);
xnor U11897 (N_11897,N_11163,N_11008);
and U11898 (N_11898,N_10504,N_11218);
nor U11899 (N_11899,N_10108,N_11005);
xor U11900 (N_11900,N_10485,N_10693);
nor U11901 (N_11901,N_10428,N_11080);
nor U11902 (N_11902,N_10097,N_10012);
nor U11903 (N_11903,N_10623,N_10320);
and U11904 (N_11904,N_10052,N_10272);
xor U11905 (N_11905,N_11063,N_10534);
and U11906 (N_11906,N_11029,N_10570);
or U11907 (N_11907,N_10055,N_11155);
and U11908 (N_11908,N_10343,N_10274);
nor U11909 (N_11909,N_11172,N_10895);
nand U11910 (N_11910,N_10335,N_11147);
nand U11911 (N_11911,N_10216,N_10986);
xor U11912 (N_11912,N_10193,N_10776);
nor U11913 (N_11913,N_10661,N_11135);
or U11914 (N_11914,N_10439,N_10832);
and U11915 (N_11915,N_10638,N_10271);
nor U11916 (N_11916,N_10846,N_10051);
or U11917 (N_11917,N_10428,N_11248);
or U11918 (N_11918,N_11171,N_11137);
and U11919 (N_11919,N_10880,N_10420);
nand U11920 (N_11920,N_10502,N_10700);
and U11921 (N_11921,N_10210,N_11116);
nand U11922 (N_11922,N_10646,N_10397);
nand U11923 (N_11923,N_10397,N_11082);
or U11924 (N_11924,N_10276,N_10450);
and U11925 (N_11925,N_10290,N_10301);
or U11926 (N_11926,N_10407,N_10364);
nand U11927 (N_11927,N_11137,N_11246);
nand U11928 (N_11928,N_10628,N_10796);
nor U11929 (N_11929,N_10298,N_11147);
nand U11930 (N_11930,N_10718,N_10781);
or U11931 (N_11931,N_10404,N_10907);
xor U11932 (N_11932,N_10925,N_11004);
nor U11933 (N_11933,N_10115,N_10616);
xnor U11934 (N_11934,N_10839,N_10778);
nor U11935 (N_11935,N_10357,N_11227);
nand U11936 (N_11936,N_10102,N_10492);
xor U11937 (N_11937,N_11003,N_10220);
xnor U11938 (N_11938,N_10806,N_10158);
and U11939 (N_11939,N_10515,N_10687);
xor U11940 (N_11940,N_11014,N_10214);
nor U11941 (N_11941,N_10105,N_10169);
and U11942 (N_11942,N_10272,N_11020);
xnor U11943 (N_11943,N_10722,N_10706);
and U11944 (N_11944,N_10430,N_11040);
nor U11945 (N_11945,N_10748,N_10516);
nand U11946 (N_11946,N_10954,N_10226);
or U11947 (N_11947,N_10163,N_10780);
nor U11948 (N_11948,N_10672,N_10891);
nand U11949 (N_11949,N_10685,N_10829);
nor U11950 (N_11950,N_10003,N_11083);
nand U11951 (N_11951,N_10059,N_10474);
xnor U11952 (N_11952,N_10011,N_10257);
and U11953 (N_11953,N_10023,N_10349);
nor U11954 (N_11954,N_10362,N_10435);
or U11955 (N_11955,N_11063,N_10909);
xnor U11956 (N_11956,N_10338,N_10534);
nand U11957 (N_11957,N_11125,N_10025);
xor U11958 (N_11958,N_10297,N_11007);
nand U11959 (N_11959,N_10207,N_10129);
xnor U11960 (N_11960,N_10666,N_11018);
and U11961 (N_11961,N_10386,N_10849);
and U11962 (N_11962,N_10902,N_10393);
xor U11963 (N_11963,N_10233,N_11111);
nor U11964 (N_11964,N_10462,N_11049);
and U11965 (N_11965,N_10205,N_10488);
or U11966 (N_11966,N_10809,N_10036);
and U11967 (N_11967,N_10530,N_11100);
and U11968 (N_11968,N_11188,N_10127);
or U11969 (N_11969,N_10247,N_10572);
or U11970 (N_11970,N_10408,N_10520);
or U11971 (N_11971,N_10439,N_10999);
or U11972 (N_11972,N_10523,N_10554);
xor U11973 (N_11973,N_10385,N_10303);
nand U11974 (N_11974,N_10482,N_10640);
and U11975 (N_11975,N_11119,N_10188);
nor U11976 (N_11976,N_10069,N_10354);
and U11977 (N_11977,N_10677,N_10420);
nand U11978 (N_11978,N_10432,N_10924);
nor U11979 (N_11979,N_10853,N_10079);
xor U11980 (N_11980,N_10768,N_10432);
xor U11981 (N_11981,N_10945,N_10356);
xnor U11982 (N_11982,N_11052,N_10501);
nor U11983 (N_11983,N_10351,N_11209);
xor U11984 (N_11984,N_10986,N_10388);
and U11985 (N_11985,N_10742,N_11067);
nand U11986 (N_11986,N_10009,N_10358);
nand U11987 (N_11987,N_10406,N_10593);
xnor U11988 (N_11988,N_11190,N_11054);
nand U11989 (N_11989,N_10721,N_10004);
and U11990 (N_11990,N_10991,N_10592);
xnor U11991 (N_11991,N_10591,N_10426);
nor U11992 (N_11992,N_11197,N_10329);
and U11993 (N_11993,N_10072,N_11168);
nand U11994 (N_11994,N_11198,N_10727);
or U11995 (N_11995,N_10969,N_10348);
and U11996 (N_11996,N_11118,N_10292);
xnor U11997 (N_11997,N_10857,N_10579);
or U11998 (N_11998,N_10410,N_10636);
xnor U11999 (N_11999,N_10902,N_10799);
or U12000 (N_12000,N_11081,N_10707);
and U12001 (N_12001,N_11199,N_10016);
xor U12002 (N_12002,N_10260,N_10716);
and U12003 (N_12003,N_11034,N_10843);
nor U12004 (N_12004,N_10756,N_10450);
or U12005 (N_12005,N_10464,N_10775);
or U12006 (N_12006,N_10221,N_10537);
nand U12007 (N_12007,N_10391,N_10159);
or U12008 (N_12008,N_10212,N_11227);
nor U12009 (N_12009,N_10832,N_10295);
xor U12010 (N_12010,N_10026,N_10551);
or U12011 (N_12011,N_10615,N_10488);
nor U12012 (N_12012,N_10732,N_10181);
nand U12013 (N_12013,N_11131,N_10043);
or U12014 (N_12014,N_10436,N_10072);
nand U12015 (N_12015,N_11086,N_10673);
xnor U12016 (N_12016,N_11122,N_10381);
nor U12017 (N_12017,N_10406,N_10357);
or U12018 (N_12018,N_11158,N_10415);
xor U12019 (N_12019,N_10440,N_10490);
or U12020 (N_12020,N_10763,N_11076);
and U12021 (N_12021,N_10579,N_11158);
nand U12022 (N_12022,N_10465,N_11066);
and U12023 (N_12023,N_10825,N_10663);
or U12024 (N_12024,N_10500,N_10691);
nor U12025 (N_12025,N_10656,N_10240);
or U12026 (N_12026,N_10736,N_10532);
or U12027 (N_12027,N_11034,N_10077);
nor U12028 (N_12028,N_10668,N_10494);
nand U12029 (N_12029,N_10914,N_10749);
or U12030 (N_12030,N_10398,N_10878);
nand U12031 (N_12031,N_10250,N_10673);
xor U12032 (N_12032,N_10653,N_10519);
and U12033 (N_12033,N_10502,N_10298);
xor U12034 (N_12034,N_10011,N_10673);
nand U12035 (N_12035,N_10251,N_11206);
xnor U12036 (N_12036,N_10286,N_10134);
xnor U12037 (N_12037,N_10304,N_10594);
xor U12038 (N_12038,N_11242,N_11212);
xnor U12039 (N_12039,N_10821,N_11230);
nor U12040 (N_12040,N_10466,N_11154);
xor U12041 (N_12041,N_11142,N_10883);
or U12042 (N_12042,N_10806,N_10837);
nor U12043 (N_12043,N_10698,N_10675);
nand U12044 (N_12044,N_11193,N_10406);
nand U12045 (N_12045,N_10589,N_10178);
or U12046 (N_12046,N_11247,N_10188);
or U12047 (N_12047,N_10267,N_10179);
nand U12048 (N_12048,N_11090,N_11244);
and U12049 (N_12049,N_10432,N_10842);
nand U12050 (N_12050,N_11144,N_10405);
and U12051 (N_12051,N_10999,N_11015);
and U12052 (N_12052,N_10861,N_10927);
nand U12053 (N_12053,N_10402,N_10043);
or U12054 (N_12054,N_10363,N_10423);
nand U12055 (N_12055,N_10096,N_10882);
nand U12056 (N_12056,N_11074,N_10550);
xnor U12057 (N_12057,N_10132,N_10716);
or U12058 (N_12058,N_10021,N_10101);
and U12059 (N_12059,N_10141,N_10273);
nor U12060 (N_12060,N_10987,N_10147);
nand U12061 (N_12061,N_10477,N_11248);
and U12062 (N_12062,N_10248,N_10502);
nor U12063 (N_12063,N_10456,N_10280);
nor U12064 (N_12064,N_10030,N_10967);
and U12065 (N_12065,N_11074,N_10823);
xor U12066 (N_12066,N_10698,N_10540);
nor U12067 (N_12067,N_11037,N_10716);
nor U12068 (N_12068,N_11249,N_10761);
or U12069 (N_12069,N_10838,N_10087);
nor U12070 (N_12070,N_10340,N_10261);
and U12071 (N_12071,N_11197,N_10974);
nand U12072 (N_12072,N_10154,N_10353);
xor U12073 (N_12073,N_11030,N_10958);
nor U12074 (N_12074,N_10413,N_11102);
and U12075 (N_12075,N_10807,N_10406);
and U12076 (N_12076,N_10167,N_10569);
xor U12077 (N_12077,N_10740,N_10737);
and U12078 (N_12078,N_10643,N_10558);
nor U12079 (N_12079,N_11165,N_10996);
xnor U12080 (N_12080,N_11054,N_10023);
xnor U12081 (N_12081,N_10663,N_10251);
and U12082 (N_12082,N_10083,N_10491);
nor U12083 (N_12083,N_10096,N_10707);
or U12084 (N_12084,N_10675,N_10076);
nand U12085 (N_12085,N_10467,N_10274);
xor U12086 (N_12086,N_10739,N_10980);
nand U12087 (N_12087,N_11024,N_10067);
or U12088 (N_12088,N_10613,N_10555);
nand U12089 (N_12089,N_10594,N_10436);
and U12090 (N_12090,N_10827,N_11159);
or U12091 (N_12091,N_10887,N_10422);
nor U12092 (N_12092,N_10541,N_10430);
nor U12093 (N_12093,N_11029,N_10043);
nand U12094 (N_12094,N_10458,N_10603);
xnor U12095 (N_12095,N_10620,N_11197);
or U12096 (N_12096,N_10388,N_10439);
xnor U12097 (N_12097,N_10048,N_11106);
xor U12098 (N_12098,N_10195,N_10321);
and U12099 (N_12099,N_10502,N_10360);
nor U12100 (N_12100,N_10562,N_10321);
or U12101 (N_12101,N_11166,N_10197);
xor U12102 (N_12102,N_10970,N_10140);
and U12103 (N_12103,N_10408,N_11040);
nand U12104 (N_12104,N_10837,N_11118);
nor U12105 (N_12105,N_10378,N_10628);
nor U12106 (N_12106,N_10221,N_10592);
and U12107 (N_12107,N_11152,N_11055);
nor U12108 (N_12108,N_10054,N_10586);
xnor U12109 (N_12109,N_10942,N_10840);
or U12110 (N_12110,N_10380,N_10116);
or U12111 (N_12111,N_10367,N_10021);
nand U12112 (N_12112,N_10270,N_10578);
nand U12113 (N_12113,N_11111,N_10043);
xnor U12114 (N_12114,N_10806,N_10600);
and U12115 (N_12115,N_10406,N_10136);
and U12116 (N_12116,N_11175,N_10119);
nor U12117 (N_12117,N_10188,N_10293);
nand U12118 (N_12118,N_10452,N_10907);
and U12119 (N_12119,N_10055,N_10469);
and U12120 (N_12120,N_10748,N_10806);
or U12121 (N_12121,N_10237,N_10017);
and U12122 (N_12122,N_10222,N_11225);
xor U12123 (N_12123,N_11085,N_10965);
xor U12124 (N_12124,N_10867,N_10397);
xor U12125 (N_12125,N_10932,N_10161);
and U12126 (N_12126,N_10302,N_10034);
nor U12127 (N_12127,N_10974,N_10243);
and U12128 (N_12128,N_10450,N_10113);
and U12129 (N_12129,N_10063,N_10441);
nand U12130 (N_12130,N_10635,N_10851);
xor U12131 (N_12131,N_10163,N_10107);
xnor U12132 (N_12132,N_11172,N_10991);
and U12133 (N_12133,N_10149,N_10627);
or U12134 (N_12134,N_10764,N_10488);
and U12135 (N_12135,N_10276,N_10638);
and U12136 (N_12136,N_10396,N_10270);
xnor U12137 (N_12137,N_10441,N_10090);
and U12138 (N_12138,N_10887,N_11180);
xnor U12139 (N_12139,N_10163,N_11187);
and U12140 (N_12140,N_10049,N_10303);
nand U12141 (N_12141,N_10255,N_10619);
nor U12142 (N_12142,N_11130,N_10126);
nor U12143 (N_12143,N_10457,N_10997);
or U12144 (N_12144,N_11208,N_10603);
xnor U12145 (N_12145,N_10637,N_11061);
and U12146 (N_12146,N_10636,N_10867);
and U12147 (N_12147,N_10388,N_11042);
and U12148 (N_12148,N_10266,N_11204);
nand U12149 (N_12149,N_10911,N_10191);
nor U12150 (N_12150,N_10717,N_10513);
nor U12151 (N_12151,N_10037,N_11143);
or U12152 (N_12152,N_10320,N_10280);
and U12153 (N_12153,N_10438,N_10436);
and U12154 (N_12154,N_10869,N_10240);
or U12155 (N_12155,N_10216,N_10660);
nand U12156 (N_12156,N_10092,N_10868);
and U12157 (N_12157,N_11158,N_10787);
or U12158 (N_12158,N_10712,N_10656);
nand U12159 (N_12159,N_11164,N_10056);
nand U12160 (N_12160,N_10623,N_10211);
nand U12161 (N_12161,N_10551,N_10982);
and U12162 (N_12162,N_10798,N_10642);
or U12163 (N_12163,N_10824,N_10712);
nand U12164 (N_12164,N_11175,N_10934);
nor U12165 (N_12165,N_10886,N_10913);
nand U12166 (N_12166,N_10793,N_11209);
nand U12167 (N_12167,N_10205,N_10639);
xnor U12168 (N_12168,N_10732,N_10204);
nor U12169 (N_12169,N_10800,N_10182);
xor U12170 (N_12170,N_10662,N_10515);
and U12171 (N_12171,N_10196,N_10345);
xor U12172 (N_12172,N_11123,N_10123);
xnor U12173 (N_12173,N_10510,N_10504);
and U12174 (N_12174,N_10883,N_10400);
xnor U12175 (N_12175,N_10543,N_10056);
or U12176 (N_12176,N_10649,N_11070);
and U12177 (N_12177,N_10360,N_10585);
xor U12178 (N_12178,N_10111,N_10673);
and U12179 (N_12179,N_10167,N_10102);
or U12180 (N_12180,N_10417,N_10223);
or U12181 (N_12181,N_10651,N_10873);
nand U12182 (N_12182,N_11049,N_10591);
nand U12183 (N_12183,N_10090,N_10741);
or U12184 (N_12184,N_10123,N_11194);
xor U12185 (N_12185,N_10981,N_10094);
and U12186 (N_12186,N_10766,N_11017);
or U12187 (N_12187,N_10020,N_10304);
and U12188 (N_12188,N_10425,N_11179);
and U12189 (N_12189,N_10739,N_11179);
and U12190 (N_12190,N_10475,N_10585);
nor U12191 (N_12191,N_11199,N_11216);
or U12192 (N_12192,N_11174,N_10975);
and U12193 (N_12193,N_10668,N_11205);
and U12194 (N_12194,N_10666,N_11144);
or U12195 (N_12195,N_10252,N_11199);
and U12196 (N_12196,N_10063,N_11071);
and U12197 (N_12197,N_10751,N_10792);
nor U12198 (N_12198,N_11138,N_10226);
or U12199 (N_12199,N_10996,N_10565);
xor U12200 (N_12200,N_11166,N_10013);
nand U12201 (N_12201,N_10123,N_11064);
and U12202 (N_12202,N_10351,N_10938);
or U12203 (N_12203,N_10189,N_10693);
nor U12204 (N_12204,N_10438,N_11139);
nor U12205 (N_12205,N_10651,N_10427);
or U12206 (N_12206,N_10325,N_10808);
and U12207 (N_12207,N_10551,N_10702);
and U12208 (N_12208,N_10479,N_10334);
nor U12209 (N_12209,N_11242,N_10387);
or U12210 (N_12210,N_10948,N_10871);
and U12211 (N_12211,N_10755,N_10839);
and U12212 (N_12212,N_10002,N_11219);
or U12213 (N_12213,N_10777,N_10630);
or U12214 (N_12214,N_10727,N_10624);
or U12215 (N_12215,N_10854,N_10478);
nor U12216 (N_12216,N_10964,N_10073);
nor U12217 (N_12217,N_10483,N_10649);
nand U12218 (N_12218,N_10104,N_11187);
and U12219 (N_12219,N_10483,N_11067);
xor U12220 (N_12220,N_10084,N_10456);
or U12221 (N_12221,N_10415,N_10527);
and U12222 (N_12222,N_10553,N_10018);
xnor U12223 (N_12223,N_11078,N_10969);
nor U12224 (N_12224,N_10159,N_10189);
or U12225 (N_12225,N_11146,N_10756);
nor U12226 (N_12226,N_10540,N_10946);
nand U12227 (N_12227,N_10174,N_11012);
nor U12228 (N_12228,N_10587,N_10032);
nor U12229 (N_12229,N_10878,N_10904);
nand U12230 (N_12230,N_10766,N_10681);
or U12231 (N_12231,N_10979,N_10328);
xnor U12232 (N_12232,N_10799,N_11191);
nor U12233 (N_12233,N_10337,N_10809);
nor U12234 (N_12234,N_10209,N_10087);
and U12235 (N_12235,N_11113,N_11177);
and U12236 (N_12236,N_10448,N_10554);
nand U12237 (N_12237,N_10733,N_10773);
and U12238 (N_12238,N_10948,N_10737);
nand U12239 (N_12239,N_10499,N_10823);
nand U12240 (N_12240,N_10631,N_10670);
xor U12241 (N_12241,N_10387,N_10856);
nand U12242 (N_12242,N_10181,N_10505);
xor U12243 (N_12243,N_10385,N_11247);
and U12244 (N_12244,N_10250,N_10408);
and U12245 (N_12245,N_10046,N_10132);
nand U12246 (N_12246,N_10435,N_11193);
nor U12247 (N_12247,N_10133,N_11018);
nand U12248 (N_12248,N_10375,N_10136);
xnor U12249 (N_12249,N_10999,N_11233);
xnor U12250 (N_12250,N_11205,N_11098);
or U12251 (N_12251,N_10623,N_11212);
xor U12252 (N_12252,N_10591,N_10447);
nor U12253 (N_12253,N_10358,N_10198);
nor U12254 (N_12254,N_10788,N_11138);
and U12255 (N_12255,N_10248,N_11132);
and U12256 (N_12256,N_10484,N_11044);
nand U12257 (N_12257,N_10936,N_11177);
nor U12258 (N_12258,N_11121,N_10394);
nor U12259 (N_12259,N_10508,N_10915);
nand U12260 (N_12260,N_11028,N_10201);
or U12261 (N_12261,N_10112,N_10101);
nand U12262 (N_12262,N_10420,N_10235);
nand U12263 (N_12263,N_10144,N_10763);
or U12264 (N_12264,N_10757,N_11039);
and U12265 (N_12265,N_10472,N_10376);
and U12266 (N_12266,N_10188,N_10526);
nand U12267 (N_12267,N_11155,N_11169);
and U12268 (N_12268,N_11229,N_11120);
and U12269 (N_12269,N_10443,N_10827);
or U12270 (N_12270,N_10915,N_10457);
and U12271 (N_12271,N_10047,N_10991);
nor U12272 (N_12272,N_10501,N_10766);
nor U12273 (N_12273,N_10473,N_11222);
or U12274 (N_12274,N_10773,N_11178);
and U12275 (N_12275,N_10607,N_10260);
or U12276 (N_12276,N_10752,N_10692);
or U12277 (N_12277,N_10512,N_11217);
nor U12278 (N_12278,N_10818,N_11244);
nand U12279 (N_12279,N_10203,N_10588);
nor U12280 (N_12280,N_10263,N_10131);
xor U12281 (N_12281,N_10023,N_10283);
nand U12282 (N_12282,N_10331,N_10589);
xnor U12283 (N_12283,N_10747,N_10594);
xor U12284 (N_12284,N_10635,N_10981);
or U12285 (N_12285,N_10064,N_10303);
xnor U12286 (N_12286,N_10652,N_10467);
nor U12287 (N_12287,N_11009,N_10385);
xnor U12288 (N_12288,N_10571,N_10921);
or U12289 (N_12289,N_11185,N_10669);
nor U12290 (N_12290,N_10730,N_10462);
or U12291 (N_12291,N_10945,N_10958);
xor U12292 (N_12292,N_10953,N_10835);
or U12293 (N_12293,N_10322,N_10391);
nor U12294 (N_12294,N_11062,N_11004);
or U12295 (N_12295,N_10175,N_11227);
or U12296 (N_12296,N_10911,N_10743);
xor U12297 (N_12297,N_10183,N_10269);
nand U12298 (N_12298,N_10932,N_10253);
and U12299 (N_12299,N_10493,N_10818);
or U12300 (N_12300,N_10498,N_10163);
nor U12301 (N_12301,N_11220,N_11015);
and U12302 (N_12302,N_10514,N_10268);
or U12303 (N_12303,N_10841,N_10371);
or U12304 (N_12304,N_10670,N_10507);
xor U12305 (N_12305,N_10916,N_10364);
or U12306 (N_12306,N_11046,N_10487);
xor U12307 (N_12307,N_10564,N_10619);
nand U12308 (N_12308,N_10945,N_11205);
nor U12309 (N_12309,N_10619,N_10094);
nor U12310 (N_12310,N_10600,N_10998);
and U12311 (N_12311,N_10783,N_10376);
or U12312 (N_12312,N_11012,N_10950);
nor U12313 (N_12313,N_10108,N_10635);
xor U12314 (N_12314,N_10045,N_10586);
xor U12315 (N_12315,N_10624,N_10869);
xor U12316 (N_12316,N_10384,N_10296);
and U12317 (N_12317,N_11218,N_10168);
xor U12318 (N_12318,N_10606,N_11236);
and U12319 (N_12319,N_10413,N_10636);
xnor U12320 (N_12320,N_10383,N_10821);
nor U12321 (N_12321,N_10199,N_10226);
nand U12322 (N_12322,N_11152,N_10769);
and U12323 (N_12323,N_11161,N_10577);
or U12324 (N_12324,N_11245,N_10602);
xnor U12325 (N_12325,N_11002,N_10673);
nand U12326 (N_12326,N_10841,N_10127);
nor U12327 (N_12327,N_10629,N_11127);
nand U12328 (N_12328,N_10550,N_10423);
xor U12329 (N_12329,N_10721,N_10639);
xnor U12330 (N_12330,N_10311,N_10228);
xnor U12331 (N_12331,N_10222,N_10689);
and U12332 (N_12332,N_10201,N_10668);
or U12333 (N_12333,N_10299,N_11230);
nor U12334 (N_12334,N_10676,N_11220);
xnor U12335 (N_12335,N_10358,N_10240);
nor U12336 (N_12336,N_10760,N_11104);
nor U12337 (N_12337,N_10488,N_10758);
xor U12338 (N_12338,N_10358,N_10762);
or U12339 (N_12339,N_10026,N_10336);
or U12340 (N_12340,N_10357,N_10455);
xor U12341 (N_12341,N_10389,N_10023);
nor U12342 (N_12342,N_10760,N_11058);
nor U12343 (N_12343,N_10922,N_11117);
xor U12344 (N_12344,N_10817,N_10393);
xor U12345 (N_12345,N_10834,N_10237);
or U12346 (N_12346,N_10762,N_10262);
nand U12347 (N_12347,N_10134,N_10583);
or U12348 (N_12348,N_10517,N_10575);
nor U12349 (N_12349,N_11105,N_10264);
nor U12350 (N_12350,N_10514,N_10339);
or U12351 (N_12351,N_10119,N_10673);
nand U12352 (N_12352,N_10522,N_10545);
xor U12353 (N_12353,N_10182,N_10985);
xnor U12354 (N_12354,N_10287,N_11234);
and U12355 (N_12355,N_10297,N_11172);
or U12356 (N_12356,N_10800,N_10913);
and U12357 (N_12357,N_10210,N_10890);
nor U12358 (N_12358,N_10422,N_11165);
or U12359 (N_12359,N_10053,N_10722);
or U12360 (N_12360,N_10230,N_11098);
or U12361 (N_12361,N_10634,N_10251);
and U12362 (N_12362,N_10061,N_10779);
xnor U12363 (N_12363,N_10048,N_10379);
and U12364 (N_12364,N_10454,N_10269);
nor U12365 (N_12365,N_11198,N_11013);
nor U12366 (N_12366,N_10175,N_10370);
nand U12367 (N_12367,N_10402,N_10512);
xnor U12368 (N_12368,N_10035,N_11160);
nand U12369 (N_12369,N_10152,N_11131);
nand U12370 (N_12370,N_10746,N_10185);
or U12371 (N_12371,N_10045,N_10351);
and U12372 (N_12372,N_10921,N_10634);
nor U12373 (N_12373,N_10318,N_10995);
and U12374 (N_12374,N_10743,N_10575);
and U12375 (N_12375,N_10693,N_11177);
nor U12376 (N_12376,N_10870,N_10763);
or U12377 (N_12377,N_10916,N_11065);
xor U12378 (N_12378,N_10310,N_10896);
and U12379 (N_12379,N_10202,N_10491);
nand U12380 (N_12380,N_10586,N_10264);
and U12381 (N_12381,N_10960,N_10518);
and U12382 (N_12382,N_10038,N_10305);
xnor U12383 (N_12383,N_10196,N_10565);
and U12384 (N_12384,N_10443,N_10233);
nand U12385 (N_12385,N_10009,N_11230);
nand U12386 (N_12386,N_10551,N_10412);
nor U12387 (N_12387,N_10969,N_10386);
nor U12388 (N_12388,N_10852,N_10723);
or U12389 (N_12389,N_10890,N_10238);
xor U12390 (N_12390,N_10035,N_10301);
nand U12391 (N_12391,N_10207,N_10249);
xor U12392 (N_12392,N_10148,N_10008);
or U12393 (N_12393,N_10495,N_10506);
and U12394 (N_12394,N_10148,N_10909);
or U12395 (N_12395,N_10994,N_10945);
or U12396 (N_12396,N_10602,N_10027);
xor U12397 (N_12397,N_10211,N_10744);
nor U12398 (N_12398,N_10860,N_10104);
nor U12399 (N_12399,N_10327,N_10342);
xor U12400 (N_12400,N_10188,N_10421);
nor U12401 (N_12401,N_10434,N_11018);
nand U12402 (N_12402,N_11114,N_11207);
and U12403 (N_12403,N_10567,N_10047);
and U12404 (N_12404,N_10072,N_11162);
nor U12405 (N_12405,N_10522,N_10159);
xor U12406 (N_12406,N_11089,N_11037);
or U12407 (N_12407,N_10711,N_10288);
or U12408 (N_12408,N_10884,N_11042);
and U12409 (N_12409,N_11103,N_11178);
and U12410 (N_12410,N_10808,N_11078);
xor U12411 (N_12411,N_11186,N_10452);
or U12412 (N_12412,N_10996,N_10109);
and U12413 (N_12413,N_10978,N_10625);
nor U12414 (N_12414,N_10374,N_10915);
or U12415 (N_12415,N_10567,N_10308);
or U12416 (N_12416,N_10861,N_10258);
or U12417 (N_12417,N_10170,N_10392);
and U12418 (N_12418,N_10527,N_10841);
xor U12419 (N_12419,N_10595,N_10306);
nand U12420 (N_12420,N_10602,N_11028);
and U12421 (N_12421,N_10221,N_10430);
nor U12422 (N_12422,N_10303,N_10813);
or U12423 (N_12423,N_10946,N_10986);
and U12424 (N_12424,N_11249,N_10913);
nor U12425 (N_12425,N_10903,N_10511);
and U12426 (N_12426,N_10582,N_10032);
nand U12427 (N_12427,N_10895,N_10106);
and U12428 (N_12428,N_10561,N_10366);
xor U12429 (N_12429,N_10431,N_10638);
nand U12430 (N_12430,N_10140,N_11039);
nand U12431 (N_12431,N_10980,N_10183);
xnor U12432 (N_12432,N_10246,N_10375);
and U12433 (N_12433,N_10217,N_11178);
and U12434 (N_12434,N_10339,N_10287);
xnor U12435 (N_12435,N_10804,N_10983);
nand U12436 (N_12436,N_10175,N_10309);
nand U12437 (N_12437,N_10624,N_10019);
nand U12438 (N_12438,N_10599,N_10695);
or U12439 (N_12439,N_11086,N_10834);
nand U12440 (N_12440,N_10398,N_11087);
nand U12441 (N_12441,N_10489,N_10950);
or U12442 (N_12442,N_11072,N_10259);
xor U12443 (N_12443,N_10615,N_11212);
nor U12444 (N_12444,N_10084,N_10965);
and U12445 (N_12445,N_10087,N_11038);
or U12446 (N_12446,N_11237,N_10847);
nor U12447 (N_12447,N_10737,N_10025);
nor U12448 (N_12448,N_11226,N_10971);
nor U12449 (N_12449,N_11107,N_10523);
nor U12450 (N_12450,N_11137,N_10150);
or U12451 (N_12451,N_10932,N_10672);
or U12452 (N_12452,N_10849,N_10677);
nand U12453 (N_12453,N_10595,N_11190);
nor U12454 (N_12454,N_10299,N_10368);
and U12455 (N_12455,N_11065,N_11139);
or U12456 (N_12456,N_10695,N_11198);
or U12457 (N_12457,N_10802,N_10247);
nand U12458 (N_12458,N_10857,N_10003);
or U12459 (N_12459,N_10595,N_10332);
and U12460 (N_12460,N_10489,N_10840);
nor U12461 (N_12461,N_10966,N_10495);
and U12462 (N_12462,N_10258,N_10440);
xnor U12463 (N_12463,N_10562,N_10285);
and U12464 (N_12464,N_10995,N_10841);
nor U12465 (N_12465,N_11098,N_10933);
nand U12466 (N_12466,N_10009,N_10922);
nor U12467 (N_12467,N_11212,N_10521);
xor U12468 (N_12468,N_10605,N_10839);
or U12469 (N_12469,N_11182,N_10047);
xnor U12470 (N_12470,N_10147,N_10104);
or U12471 (N_12471,N_10709,N_11074);
nor U12472 (N_12472,N_10397,N_10017);
xor U12473 (N_12473,N_10069,N_11020);
nor U12474 (N_12474,N_10648,N_10071);
and U12475 (N_12475,N_10465,N_11148);
nor U12476 (N_12476,N_10733,N_10530);
and U12477 (N_12477,N_10185,N_10061);
or U12478 (N_12478,N_10107,N_10164);
nor U12479 (N_12479,N_11021,N_11155);
and U12480 (N_12480,N_10717,N_10517);
nand U12481 (N_12481,N_11204,N_10103);
nand U12482 (N_12482,N_10922,N_10797);
nand U12483 (N_12483,N_11221,N_11234);
xnor U12484 (N_12484,N_10562,N_10904);
or U12485 (N_12485,N_10395,N_10246);
xnor U12486 (N_12486,N_10437,N_10304);
and U12487 (N_12487,N_10506,N_10691);
xnor U12488 (N_12488,N_10491,N_11157);
and U12489 (N_12489,N_10588,N_10125);
nand U12490 (N_12490,N_11122,N_10194);
nor U12491 (N_12491,N_10719,N_10070);
xnor U12492 (N_12492,N_10117,N_10768);
nand U12493 (N_12493,N_10701,N_10917);
xnor U12494 (N_12494,N_10130,N_10667);
or U12495 (N_12495,N_11187,N_10030);
or U12496 (N_12496,N_10632,N_10997);
nor U12497 (N_12497,N_10496,N_10494);
nor U12498 (N_12498,N_10363,N_10721);
nand U12499 (N_12499,N_10241,N_10396);
xor U12500 (N_12500,N_12181,N_11265);
or U12501 (N_12501,N_12256,N_11798);
xor U12502 (N_12502,N_12331,N_11693);
nor U12503 (N_12503,N_11803,N_11745);
nor U12504 (N_12504,N_12056,N_11593);
nand U12505 (N_12505,N_11450,N_12433);
nor U12506 (N_12506,N_12035,N_12067);
xor U12507 (N_12507,N_11274,N_12269);
and U12508 (N_12508,N_11864,N_11638);
xor U12509 (N_12509,N_11543,N_11284);
and U12510 (N_12510,N_11773,N_11464);
xor U12511 (N_12511,N_12032,N_11454);
nor U12512 (N_12512,N_11902,N_11588);
nor U12513 (N_12513,N_12237,N_12472);
nand U12514 (N_12514,N_11533,N_11566);
or U12515 (N_12515,N_11913,N_12248);
and U12516 (N_12516,N_11659,N_11525);
or U12517 (N_12517,N_12274,N_12159);
nand U12518 (N_12518,N_11760,N_12427);
or U12519 (N_12519,N_12136,N_12493);
xor U12520 (N_12520,N_12455,N_12088);
nor U12521 (N_12521,N_12359,N_12036);
or U12522 (N_12522,N_11639,N_12358);
nor U12523 (N_12523,N_11948,N_12339);
xor U12524 (N_12524,N_11433,N_11429);
nand U12525 (N_12525,N_12126,N_11757);
nand U12526 (N_12526,N_11635,N_12110);
or U12527 (N_12527,N_11865,N_12250);
nand U12528 (N_12528,N_11992,N_12327);
and U12529 (N_12529,N_11586,N_11342);
xnor U12530 (N_12530,N_12430,N_11895);
nor U12531 (N_12531,N_11774,N_11658);
or U12532 (N_12532,N_11893,N_12075);
xnor U12533 (N_12533,N_11997,N_11414);
nand U12534 (N_12534,N_12115,N_12309);
nand U12535 (N_12535,N_11351,N_12481);
nand U12536 (N_12536,N_12325,N_11544);
xnor U12537 (N_12537,N_11924,N_11797);
or U12538 (N_12538,N_11363,N_12361);
nand U12539 (N_12539,N_12293,N_11538);
and U12540 (N_12540,N_11617,N_12047);
and U12541 (N_12541,N_12192,N_12260);
or U12542 (N_12542,N_11619,N_11386);
and U12543 (N_12543,N_11636,N_12005);
or U12544 (N_12544,N_12442,N_11350);
nor U12545 (N_12545,N_11879,N_11633);
nor U12546 (N_12546,N_11297,N_11294);
xnor U12547 (N_12547,N_11648,N_11710);
nor U12548 (N_12548,N_11555,N_11828);
or U12549 (N_12549,N_11596,N_11308);
and U12550 (N_12550,N_11304,N_12412);
nand U12551 (N_12551,N_11730,N_11257);
nor U12552 (N_12552,N_11813,N_11576);
or U12553 (N_12553,N_11939,N_11394);
nand U12554 (N_12554,N_11335,N_12270);
or U12555 (N_12555,N_11569,N_11759);
xnor U12556 (N_12556,N_12188,N_12348);
or U12557 (N_12557,N_11741,N_11625);
and U12558 (N_12558,N_11604,N_11618);
and U12559 (N_12559,N_11768,N_11694);
and U12560 (N_12560,N_11653,N_11995);
or U12561 (N_12561,N_11951,N_11361);
and U12562 (N_12562,N_11330,N_11842);
xnor U12563 (N_12563,N_12151,N_12400);
and U12564 (N_12564,N_11396,N_11344);
xor U12565 (N_12565,N_12350,N_12410);
nor U12566 (N_12566,N_11354,N_11298);
and U12567 (N_12567,N_12020,N_11459);
nand U12568 (N_12568,N_12375,N_12132);
nor U12569 (N_12569,N_12085,N_11871);
nor U12570 (N_12570,N_11535,N_12284);
and U12571 (N_12571,N_12295,N_11852);
xor U12572 (N_12572,N_11824,N_12408);
nor U12573 (N_12573,N_11285,N_12103);
and U12574 (N_12574,N_11985,N_11993);
nor U12575 (N_12575,N_11419,N_11845);
or U12576 (N_12576,N_12378,N_12193);
xnor U12577 (N_12577,N_11607,N_12199);
nand U12578 (N_12578,N_11258,N_11744);
xor U12579 (N_12579,N_11502,N_11885);
xnor U12580 (N_12580,N_11458,N_12145);
nand U12581 (N_12581,N_12069,N_12211);
and U12582 (N_12582,N_11352,N_11889);
nor U12583 (N_12583,N_11950,N_12060);
xnor U12584 (N_12584,N_12104,N_11349);
xnor U12585 (N_12585,N_11435,N_11436);
nand U12586 (N_12586,N_12184,N_11686);
and U12587 (N_12587,N_12143,N_11290);
xnor U12588 (N_12588,N_12089,N_12386);
and U12589 (N_12589,N_11288,N_11630);
or U12590 (N_12590,N_12329,N_12464);
or U12591 (N_12591,N_11703,N_12081);
and U12592 (N_12592,N_11971,N_11496);
xnor U12593 (N_12593,N_11862,N_12167);
xor U12594 (N_12594,N_11603,N_11882);
or U12595 (N_12595,N_12160,N_12168);
xor U12596 (N_12596,N_11994,N_11927);
or U12597 (N_12597,N_11699,N_12275);
nand U12598 (N_12598,N_12368,N_11812);
or U12599 (N_12599,N_11403,N_12096);
nand U12600 (N_12600,N_11827,N_12303);
nor U12601 (N_12601,N_11987,N_12187);
nor U12602 (N_12602,N_11339,N_12180);
or U12603 (N_12603,N_11976,N_12068);
nor U12604 (N_12604,N_12156,N_12341);
or U12605 (N_12605,N_11484,N_11567);
and U12606 (N_12606,N_11552,N_11863);
xnor U12607 (N_12607,N_11704,N_11962);
and U12608 (N_12608,N_11687,N_11624);
xor U12609 (N_12609,N_11367,N_12117);
nand U12610 (N_12610,N_12478,N_11655);
nand U12611 (N_12611,N_12407,N_11790);
xnor U12612 (N_12612,N_11983,N_11613);
xor U12613 (N_12613,N_12317,N_11846);
or U12614 (N_12614,N_12241,N_11729);
nor U12615 (N_12615,N_12306,N_11837);
nand U12616 (N_12616,N_11343,N_12015);
or U12617 (N_12617,N_12182,N_11514);
nor U12618 (N_12618,N_12024,N_12240);
xnor U12619 (N_12619,N_11307,N_11558);
xnor U12620 (N_12620,N_11937,N_12245);
and U12621 (N_12621,N_12004,N_12223);
nor U12622 (N_12622,N_11584,N_11956);
and U12623 (N_12623,N_12229,N_12164);
nor U12624 (N_12624,N_12023,N_12191);
and U12625 (N_12625,N_11861,N_11945);
xnor U12626 (N_12626,N_11276,N_12029);
or U12627 (N_12627,N_11933,N_12337);
nand U12628 (N_12628,N_12179,N_11583);
and U12629 (N_12629,N_12129,N_11984);
or U12630 (N_12630,N_12402,N_11859);
nor U12631 (N_12631,N_11462,N_11407);
xor U12632 (N_12632,N_11366,N_11900);
and U12633 (N_12633,N_11542,N_11316);
nand U12634 (N_12634,N_11910,N_11707);
xor U12635 (N_12635,N_11391,N_11300);
or U12636 (N_12636,N_12013,N_12058);
or U12637 (N_12637,N_12468,N_12347);
and U12638 (N_12638,N_12153,N_12022);
xnor U12639 (N_12639,N_12246,N_12244);
and U12640 (N_12640,N_11884,N_11752);
or U12641 (N_12641,N_11899,N_11770);
xnor U12642 (N_12642,N_11410,N_11547);
or U12643 (N_12643,N_12321,N_11428);
and U12644 (N_12644,N_11749,N_11805);
xor U12645 (N_12645,N_12443,N_11277);
nor U12646 (N_12646,N_11578,N_12077);
and U12647 (N_12647,N_11627,N_12087);
and U12648 (N_12648,N_11826,N_11794);
and U12649 (N_12649,N_12310,N_11561);
and U12650 (N_12650,N_11631,N_12112);
nor U12651 (N_12651,N_11432,N_12285);
xor U12652 (N_12652,N_12173,N_11451);
nor U12653 (N_12653,N_12186,N_12473);
or U12654 (N_12654,N_12294,N_11712);
nand U12655 (N_12655,N_12054,N_12095);
nand U12656 (N_12656,N_11782,N_12009);
or U12657 (N_12657,N_11493,N_11515);
nand U12658 (N_12658,N_11814,N_11907);
or U12659 (N_12659,N_12076,N_11581);
nand U12660 (N_12660,N_11318,N_11917);
and U12661 (N_12661,N_11660,N_11684);
nor U12662 (N_12662,N_11427,N_11326);
nand U12663 (N_12663,N_12488,N_12485);
xnor U12664 (N_12664,N_11337,N_12271);
xnor U12665 (N_12665,N_11833,N_11676);
nand U12666 (N_12666,N_12286,N_12422);
and U12667 (N_12667,N_11611,N_11528);
and U12668 (N_12668,N_11751,N_12150);
xor U12669 (N_12669,N_11637,N_11320);
or U12670 (N_12670,N_12161,N_12099);
xor U12671 (N_12671,N_12233,N_12390);
xnor U12672 (N_12672,N_12268,N_12197);
or U12673 (N_12673,N_11775,N_11315);
xor U12674 (N_12674,N_11516,N_11867);
nor U12675 (N_12675,N_12259,N_11894);
xor U12676 (N_12676,N_12314,N_12203);
and U12677 (N_12677,N_12479,N_11973);
nand U12678 (N_12678,N_11357,N_12416);
or U12679 (N_12679,N_11989,N_11548);
nand U12680 (N_12680,N_11564,N_11299);
nand U12681 (N_12681,N_11416,N_12090);
nand U12682 (N_12682,N_12258,N_12195);
nor U12683 (N_12683,N_12239,N_11711);
and U12684 (N_12684,N_11271,N_11280);
xor U12685 (N_12685,N_12201,N_11551);
or U12686 (N_12686,N_11661,N_11720);
or U12687 (N_12687,N_11892,N_12082);
xor U12688 (N_12688,N_12225,N_12498);
and U12689 (N_12689,N_12196,N_11574);
xor U12690 (N_12690,N_11906,N_11847);
or U12691 (N_12691,N_12071,N_12097);
or U12692 (N_12692,N_12255,N_11856);
nand U12693 (N_12693,N_11415,N_11811);
and U12694 (N_12694,N_12387,N_11926);
and U12695 (N_12695,N_11761,N_12469);
and U12696 (N_12696,N_11261,N_11601);
and U12697 (N_12697,N_12038,N_11979);
nor U12698 (N_12698,N_11556,N_11356);
or U12699 (N_12699,N_12397,N_12226);
nand U12700 (N_12700,N_11830,N_11563);
and U12701 (N_12701,N_12190,N_11520);
or U12702 (N_12702,N_11292,N_12323);
nor U12703 (N_12703,N_11364,N_12492);
nand U12704 (N_12704,N_11788,N_11680);
or U12705 (N_12705,N_11918,N_11641);
xnor U12706 (N_12706,N_11473,N_11713);
or U12707 (N_12707,N_11968,N_11746);
xor U12708 (N_12708,N_12119,N_11944);
nand U12709 (N_12709,N_12102,N_12431);
or U12710 (N_12710,N_11263,N_11314);
nand U12711 (N_12711,N_11536,N_11501);
and U12712 (N_12712,N_11319,N_11401);
nand U12713 (N_12713,N_12266,N_12343);
xnor U12714 (N_12714,N_11640,N_11690);
nor U12715 (N_12715,N_11408,N_12041);
or U12716 (N_12716,N_11589,N_11998);
xnor U12717 (N_12717,N_12027,N_12449);
and U12718 (N_12718,N_12218,N_12124);
nand U12719 (N_12719,N_11286,N_12424);
or U12720 (N_12720,N_12432,N_11508);
xnor U12721 (N_12721,N_12326,N_11579);
xnor U12722 (N_12722,N_11598,N_11537);
or U12723 (N_12723,N_12253,N_11876);
or U12724 (N_12724,N_12006,N_12228);
or U12725 (N_12725,N_12073,N_11549);
xnor U12726 (N_12726,N_11850,N_12474);
nor U12727 (N_12727,N_11928,N_12122);
or U12728 (N_12728,N_11384,N_11999);
nor U12729 (N_12729,N_11853,N_11657);
or U12730 (N_12730,N_12360,N_12147);
and U12731 (N_12731,N_11438,N_12209);
nand U12732 (N_12732,N_12098,N_12030);
or U12733 (N_12733,N_11786,N_11465);
nand U12734 (N_12734,N_12373,N_11978);
or U12735 (N_12735,N_11735,N_12484);
nor U12736 (N_12736,N_11594,N_11480);
nand U12737 (N_12737,N_11634,N_12497);
nor U12738 (N_12738,N_11829,N_11969);
or U12739 (N_12739,N_11309,N_12388);
nor U12740 (N_12740,N_12437,N_11644);
nand U12741 (N_12741,N_11931,N_11888);
or U12742 (N_12742,N_11755,N_11503);
xnor U12743 (N_12743,N_12101,N_11460);
or U12744 (N_12744,N_11313,N_12208);
and U12745 (N_12745,N_11990,N_12419);
nand U12746 (N_12746,N_12206,N_12413);
and U12747 (N_12747,N_12205,N_12213);
nand U12748 (N_12748,N_11560,N_12055);
nor U12749 (N_12749,N_12062,N_11402);
or U12750 (N_12750,N_11818,N_12333);
or U12751 (N_12751,N_12012,N_11816);
or U12752 (N_12752,N_12018,N_11777);
nand U12753 (N_12753,N_11540,N_12300);
or U12754 (N_12754,N_11452,N_12251);
nor U12755 (N_12755,N_11397,N_12466);
or U12756 (N_12756,N_12026,N_11801);
xor U12757 (N_12757,N_12078,N_11447);
or U12758 (N_12758,N_11970,N_12417);
nor U12759 (N_12759,N_11375,N_12460);
nand U12760 (N_12760,N_11267,N_12086);
or U12761 (N_12761,N_11869,N_11650);
xor U12762 (N_12762,N_11259,N_11311);
and U12763 (N_12763,N_11936,N_11957);
and U12764 (N_12764,N_12344,N_11742);
nor U12765 (N_12765,N_12162,N_11943);
and U12766 (N_12766,N_11738,N_12169);
nor U12767 (N_12767,N_11651,N_11353);
nor U12768 (N_12768,N_11256,N_11389);
and U12769 (N_12769,N_11793,N_12396);
or U12770 (N_12770,N_12028,N_12007);
xnor U12771 (N_12771,N_12139,N_11466);
nand U12772 (N_12772,N_11521,N_11546);
or U12773 (N_12773,N_11963,N_11810);
xor U12774 (N_12774,N_11675,N_11721);
nor U12775 (N_12775,N_11443,N_11530);
xnor U12776 (N_12776,N_11570,N_12288);
and U12777 (N_12777,N_11492,N_12141);
xnor U12778 (N_12778,N_11779,N_11647);
nand U12779 (N_12779,N_11832,N_11495);
nor U12780 (N_12780,N_12401,N_11679);
nor U12781 (N_12781,N_11996,N_11310);
nor U12782 (N_12782,N_12157,N_11822);
xor U12783 (N_12783,N_11291,N_11670);
nor U12784 (N_12784,N_12003,N_11430);
and U12785 (N_12785,N_12052,N_11441);
and U12786 (N_12786,N_12272,N_12487);
nand U12787 (N_12787,N_11295,N_12283);
xor U12788 (N_12788,N_11714,N_11872);
nand U12789 (N_12789,N_11268,N_11500);
xor U12790 (N_12790,N_12355,N_12428);
and U12791 (N_12791,N_11609,N_12311);
xor U12792 (N_12792,N_11262,N_11572);
and U12793 (N_12793,N_12114,N_12074);
and U12794 (N_12794,N_11942,N_11289);
nand U12795 (N_12795,N_11792,N_11449);
or U12796 (N_12796,N_11270,N_12072);
nor U12797 (N_12797,N_12166,N_11483);
xnor U12798 (N_12798,N_11785,N_12261);
or U12799 (N_12799,N_12480,N_11623);
nor U12800 (N_12800,N_12334,N_11266);
or U12801 (N_12801,N_11370,N_12414);
or U12802 (N_12802,N_12016,N_12049);
and U12803 (N_12803,N_11602,N_11949);
nand U12804 (N_12804,N_12470,N_11632);
nor U12805 (N_12805,N_11748,N_12264);
and U12806 (N_12806,N_11666,N_12370);
and U12807 (N_12807,N_11565,N_11485);
xor U12808 (N_12808,N_12140,N_12454);
or U12809 (N_12809,N_11799,N_12371);
nand U12810 (N_12810,N_11743,N_12389);
and U12811 (N_12811,N_11740,N_11977);
nand U12812 (N_12812,N_11843,N_11629);
nand U12813 (N_12813,N_11595,N_12461);
xnor U12814 (N_12814,N_12491,N_11839);
nor U12815 (N_12815,N_12385,N_12249);
or U12816 (N_12816,N_11920,N_12037);
or U12817 (N_12817,N_11541,N_11840);
and U12818 (N_12818,N_12281,N_12262);
or U12819 (N_12819,N_12125,N_11504);
and U12820 (N_12820,N_12267,N_11374);
or U12821 (N_12821,N_11333,N_12083);
and U12822 (N_12822,N_11424,N_11420);
nor U12823 (N_12823,N_12031,N_11781);
or U12824 (N_12824,N_12420,N_11526);
and U12825 (N_12825,N_12489,N_12495);
and U12826 (N_12826,N_11269,N_12113);
nor U12827 (N_12827,N_11880,N_11417);
nor U12828 (N_12828,N_11802,N_11669);
nand U12829 (N_12829,N_11577,N_11406);
xor U12830 (N_12830,N_12135,N_11328);
and U12831 (N_12831,N_11513,N_11848);
and U12832 (N_12832,N_12265,N_12356);
and U12833 (N_12833,N_11692,N_11385);
nor U12834 (N_12834,N_11723,N_12123);
nand U12835 (N_12835,N_11695,N_11815);
nor U12836 (N_12836,N_11463,N_11327);
or U12837 (N_12837,N_12376,N_11964);
or U12838 (N_12838,N_11725,N_11605);
nor U12839 (N_12839,N_12425,N_11562);
nor U12840 (N_12840,N_12399,N_11487);
nor U12841 (N_12841,N_12155,N_11444);
xnor U12842 (N_12842,N_12450,N_12230);
and U12843 (N_12843,N_11708,N_12384);
nand U12844 (N_12844,N_11376,N_11534);
nand U12845 (N_12845,N_11702,N_11448);
nand U12846 (N_12846,N_11475,N_12138);
and U12847 (N_12847,N_12365,N_11897);
and U12848 (N_12848,N_12210,N_12377);
nor U12849 (N_12849,N_11445,N_12045);
nand U12850 (N_12850,N_12458,N_12064);
xnor U12851 (N_12851,N_11392,N_11947);
xor U12852 (N_12852,N_12404,N_11668);
or U12853 (N_12853,N_12475,N_12398);
nor U12854 (N_12854,N_11697,N_12330);
nor U12855 (N_12855,N_12263,N_12476);
nand U12856 (N_12856,N_11980,N_11851);
nand U12857 (N_12857,N_12335,N_11512);
nand U12858 (N_12858,N_11754,N_11698);
xor U12859 (N_12859,N_11717,N_11390);
nor U12860 (N_12860,N_11358,N_11592);
nor U12861 (N_12861,N_12456,N_12462);
nand U12862 (N_12862,N_11425,N_11360);
nor U12863 (N_12863,N_11296,N_11545);
nor U12864 (N_12864,N_11854,N_12381);
xor U12865 (N_12865,N_11345,N_11672);
and U12866 (N_12866,N_11935,N_11275);
nor U12867 (N_12867,N_11914,N_11791);
or U12868 (N_12868,N_12080,N_12448);
nand U12869 (N_12869,N_12308,N_11431);
nand U12870 (N_12870,N_12346,N_11388);
nand U12871 (N_12871,N_11610,N_11573);
and U12872 (N_12872,N_11426,N_11321);
nor U12873 (N_12873,N_11626,N_11709);
nor U12874 (N_12874,N_12447,N_12332);
nor U12875 (N_12875,N_11750,N_12152);
xnor U12876 (N_12876,N_11472,N_12217);
nand U12877 (N_12877,N_11446,N_12280);
xnor U12878 (N_12878,N_12391,N_12392);
nor U12879 (N_12879,N_11421,N_12301);
nand U12880 (N_12880,N_11857,N_11412);
xnor U12881 (N_12881,N_11568,N_11615);
nor U12882 (N_12882,N_11934,N_11762);
nand U12883 (N_12883,N_12178,N_11434);
xor U12884 (N_12884,N_12000,N_12395);
and U12885 (N_12885,N_12034,N_12234);
nor U12886 (N_12886,N_11681,N_11991);
xor U12887 (N_12887,N_11718,N_11336);
nand U12888 (N_12888,N_12440,N_12299);
or U12889 (N_12889,N_12127,N_11705);
nand U12890 (N_12890,N_11682,N_12278);
xnor U12891 (N_12891,N_11398,N_11477);
and U12892 (N_12892,N_11346,N_11628);
nor U12893 (N_12893,N_11727,N_11866);
xor U12894 (N_12894,N_12232,N_12222);
nor U12895 (N_12895,N_11952,N_11789);
nor U12896 (N_12896,N_12108,N_12379);
nor U12897 (N_12897,N_11481,N_11858);
and U12898 (N_12898,N_11453,N_11456);
or U12899 (N_12899,N_12434,N_11499);
nor U12900 (N_12900,N_11347,N_12421);
or U12901 (N_12901,N_11891,N_12297);
nand U12902 (N_12902,N_12242,N_12010);
nand U12903 (N_12903,N_12444,N_11597);
xor U12904 (N_12904,N_11612,N_12121);
nand U12905 (N_12905,N_12405,N_12482);
xnor U12906 (N_12906,N_11468,N_12224);
and U12907 (N_12907,N_11616,N_11645);
xnor U12908 (N_12908,N_11489,N_11808);
nor U12909 (N_12909,N_11518,N_11874);
nand U12910 (N_12910,N_12149,N_11890);
nand U12911 (N_12911,N_11758,N_11409);
or U12912 (N_12912,N_12289,N_12471);
nor U12913 (N_12913,N_12352,N_11395);
nor U12914 (N_12914,N_11505,N_11317);
or U12915 (N_12915,N_11780,N_11961);
nand U12916 (N_12916,N_11329,N_11509);
nor U12917 (N_12917,N_11469,N_12065);
or U12918 (N_12918,N_12276,N_11901);
and U12919 (N_12919,N_11958,N_11886);
xnor U12920 (N_12920,N_11733,N_11511);
and U12921 (N_12921,N_11557,N_11380);
nor U12922 (N_12922,N_11953,N_11362);
nand U12923 (N_12923,N_11959,N_12282);
or U12924 (N_12924,N_11706,N_12011);
and U12925 (N_12925,N_11835,N_12094);
and U12926 (N_12926,N_12048,N_12292);
nand U12927 (N_12927,N_12252,N_11301);
xnor U12928 (N_12928,N_12319,N_11938);
nor U12929 (N_12929,N_11372,N_11753);
or U12930 (N_12930,N_11807,N_12409);
nor U12931 (N_12931,N_12383,N_12134);
nand U12932 (N_12932,N_12367,N_12216);
and U12933 (N_12933,N_12100,N_11825);
nor U12934 (N_12934,N_11688,N_12436);
nor U12935 (N_12935,N_11278,N_11904);
nand U12936 (N_12936,N_12322,N_11369);
nor U12937 (N_12937,N_12320,N_12118);
nor U12938 (N_12938,N_11875,N_11771);
nand U12939 (N_12939,N_11622,N_11724);
or U12940 (N_12940,N_12185,N_12316);
nor U12941 (N_12941,N_11663,N_12445);
xor U12942 (N_12942,N_12084,N_12070);
and U12943 (N_12943,N_11471,N_11359);
nand U12944 (N_12944,N_11763,N_12486);
or U12945 (N_12945,N_11665,N_11716);
xor U12946 (N_12946,N_11728,N_12457);
nor U12947 (N_12947,N_11795,N_11981);
nor U12948 (N_12948,N_11689,N_11823);
and U12949 (N_12949,N_11834,N_12014);
nand U12950 (N_12950,N_11599,N_11849);
and U12951 (N_12951,N_12406,N_11523);
or U12952 (N_12952,N_12354,N_11671);
or U12953 (N_12953,N_12017,N_11772);
xnor U12954 (N_12954,N_11820,N_12351);
nor U12955 (N_12955,N_11870,N_11532);
xor U12956 (N_12956,N_12198,N_12109);
nand U12957 (N_12957,N_12357,N_12002);
nor U12958 (N_12958,N_11778,N_11476);
or U12959 (N_12959,N_12092,N_11965);
nor U12960 (N_12960,N_12312,N_11873);
nand U12961 (N_12961,N_11413,N_12133);
xnor U12962 (N_12962,N_11582,N_11696);
and U12963 (N_12963,N_11539,N_12340);
nand U12964 (N_12964,N_11273,N_11868);
or U12965 (N_12965,N_12175,N_12042);
nor U12966 (N_12966,N_11912,N_11507);
nand U12967 (N_12967,N_12043,N_11878);
nor U12968 (N_12968,N_11908,N_11348);
nand U12969 (N_12969,N_12353,N_11877);
xnor U12970 (N_12970,N_12363,N_12438);
nor U12971 (N_12971,N_11479,N_11381);
and U12972 (N_12972,N_12290,N_11306);
nand U12973 (N_12973,N_11331,N_11966);
xnor U12974 (N_12974,N_11510,N_11455);
nand U12975 (N_12975,N_11819,N_11932);
or U12976 (N_12976,N_11921,N_11281);
xor U12977 (N_12977,N_12345,N_11929);
and U12978 (N_12978,N_11355,N_11737);
xor U12979 (N_12979,N_11497,N_12061);
nand U12980 (N_12980,N_11734,N_11519);
nand U12981 (N_12981,N_11841,N_12494);
nor U12982 (N_12982,N_11379,N_11667);
or U12983 (N_12983,N_11272,N_11664);
nor U12984 (N_12984,N_12243,N_11662);
or U12985 (N_12985,N_12040,N_11796);
and U12986 (N_12986,N_12423,N_12142);
or U12987 (N_12987,N_11338,N_12362);
nor U12988 (N_12988,N_11855,N_11250);
xnor U12989 (N_12989,N_12051,N_12200);
or U12990 (N_12990,N_11252,N_12008);
or U12991 (N_12991,N_11422,N_12465);
nand U12992 (N_12992,N_12219,N_12291);
or U12993 (N_12993,N_12338,N_12374);
nand U12994 (N_12994,N_11804,N_12411);
nand U12995 (N_12995,N_12057,N_11643);
nor U12996 (N_12996,N_12053,N_11860);
and U12997 (N_12997,N_12496,N_12441);
nor U12998 (N_12998,N_12093,N_12439);
xor U12999 (N_12999,N_11371,N_12298);
or U13000 (N_13000,N_11283,N_11494);
xor U13001 (N_13001,N_12426,N_11303);
nor U13002 (N_13002,N_11930,N_11411);
and U13003 (N_13003,N_12220,N_11575);
and U13004 (N_13004,N_11305,N_11747);
nand U13005 (N_13005,N_11522,N_12336);
xor U13006 (N_13006,N_11490,N_11423);
nand U13007 (N_13007,N_11279,N_12307);
xor U13008 (N_13008,N_11498,N_11946);
nor U13009 (N_13009,N_11253,N_12116);
nor U13010 (N_13010,N_11550,N_11726);
nor U13011 (N_13011,N_11478,N_12063);
nand U13012 (N_13012,N_11368,N_11925);
or U13013 (N_13013,N_11817,N_11919);
nor U13014 (N_13014,N_12131,N_11382);
nor U13015 (N_13015,N_12296,N_11691);
nor U13016 (N_13016,N_11554,N_11756);
nor U13017 (N_13017,N_11736,N_11787);
xnor U13018 (N_13018,N_12477,N_12453);
xnor U13019 (N_13019,N_11764,N_12236);
xnor U13020 (N_13020,N_12170,N_11491);
or U13021 (N_13021,N_12158,N_12393);
and U13022 (N_13022,N_12091,N_12235);
xnor U13023 (N_13023,N_12025,N_12146);
or U13024 (N_13024,N_11767,N_11642);
nand U13025 (N_13025,N_12174,N_12154);
and U13026 (N_13026,N_12446,N_11683);
xnor U13027 (N_13027,N_11332,N_12499);
xor U13028 (N_13028,N_11646,N_11800);
xor U13029 (N_13029,N_11529,N_11685);
nand U13030 (N_13030,N_11608,N_11393);
or U13031 (N_13031,N_12418,N_11506);
xnor U13032 (N_13032,N_12369,N_12257);
or U13033 (N_13033,N_12305,N_11474);
nand U13034 (N_13034,N_11974,N_12247);
and U13035 (N_13035,N_12059,N_11766);
nor U13036 (N_13036,N_11399,N_12215);
and U13037 (N_13037,N_12451,N_12202);
or U13038 (N_13038,N_12349,N_12066);
xnor U13039 (N_13039,N_11282,N_12148);
nor U13040 (N_13040,N_11383,N_11722);
and U13041 (N_13041,N_12324,N_12366);
or U13042 (N_13042,N_12394,N_11905);
nor U13043 (N_13043,N_12120,N_11652);
xnor U13044 (N_13044,N_11260,N_11806);
nand U13045 (N_13045,N_12459,N_12050);
and U13046 (N_13046,N_12172,N_11986);
nand U13047 (N_13047,N_12463,N_11776);
nor U13048 (N_13048,N_11881,N_11769);
and U13049 (N_13049,N_11580,N_11915);
nor U13050 (N_13050,N_11302,N_11783);
and U13051 (N_13051,N_11255,N_11251);
or U13052 (N_13052,N_11517,N_11940);
nand U13053 (N_13053,N_12177,N_12452);
xor U13054 (N_13054,N_11656,N_12313);
xnor U13055 (N_13055,N_12273,N_12106);
nor U13056 (N_13056,N_11387,N_11553);
xor U13057 (N_13057,N_12315,N_12318);
nand U13058 (N_13058,N_11982,N_11587);
or U13059 (N_13059,N_11340,N_11440);
nand U13060 (N_13060,N_12183,N_12277);
nand U13061 (N_13061,N_11486,N_12221);
xor U13062 (N_13062,N_12165,N_11325);
xnor U13063 (N_13063,N_12171,N_11620);
nand U13064 (N_13064,N_12429,N_12033);
nor U13065 (N_13065,N_11527,N_12467);
nand U13066 (N_13066,N_11606,N_11591);
nand U13067 (N_13067,N_12214,N_12304);
nand U13068 (N_13068,N_11954,N_11467);
nor U13069 (N_13069,N_12194,N_11457);
nand U13070 (N_13070,N_11559,N_12001);
nor U13071 (N_13071,N_11418,N_12128);
nand U13072 (N_13072,N_11715,N_11341);
nor U13073 (N_13073,N_11975,N_12176);
xnor U13074 (N_13074,N_11400,N_12044);
and U13075 (N_13075,N_12483,N_11600);
xnor U13076 (N_13076,N_11461,N_11821);
nand U13077 (N_13077,N_11784,N_12021);
nand U13078 (N_13078,N_12105,N_11334);
or U13079 (N_13079,N_11442,N_11571);
and U13080 (N_13080,N_11887,N_12279);
and U13081 (N_13081,N_11439,N_12302);
or U13082 (N_13082,N_11405,N_11896);
nand U13083 (N_13083,N_11254,N_11923);
nand U13084 (N_13084,N_12107,N_11955);
nor U13085 (N_13085,N_11524,N_11323);
and U13086 (N_13086,N_12207,N_12144);
nand U13087 (N_13087,N_12287,N_11883);
xor U13088 (N_13088,N_12137,N_12079);
xor U13089 (N_13089,N_11836,N_11941);
and U13090 (N_13090,N_11911,N_12238);
or U13091 (N_13091,N_11488,N_11614);
or U13092 (N_13092,N_12382,N_11838);
and U13093 (N_13093,N_12415,N_12328);
nand U13094 (N_13094,N_12435,N_11972);
xnor U13095 (N_13095,N_12019,N_11739);
nor U13096 (N_13096,N_11673,N_11701);
and U13097 (N_13097,N_12227,N_11312);
and U13098 (N_13098,N_12364,N_11377);
xnor U13099 (N_13099,N_11470,N_11831);
nor U13100 (N_13100,N_11909,N_11765);
xor U13101 (N_13101,N_12254,N_12189);
and U13102 (N_13102,N_11404,N_12231);
xor U13103 (N_13103,N_11322,N_12490);
and U13104 (N_13104,N_11531,N_11365);
xor U13105 (N_13105,N_11988,N_11731);
xor U13106 (N_13106,N_11678,N_11373);
or U13107 (N_13107,N_11967,N_12039);
nand U13108 (N_13108,N_11844,N_12204);
xor U13109 (N_13109,N_11621,N_11585);
and U13110 (N_13110,N_11654,N_11378);
xnor U13111 (N_13111,N_12046,N_12372);
nand U13112 (N_13112,N_12111,N_11590);
xnor U13113 (N_13113,N_11482,N_11700);
or U13114 (N_13114,N_11293,N_11732);
and U13115 (N_13115,N_11677,N_11264);
and U13116 (N_13116,N_12212,N_12403);
xor U13117 (N_13117,N_12130,N_11287);
nand U13118 (N_13118,N_12380,N_11649);
and U13119 (N_13119,N_11324,N_11437);
or U13120 (N_13120,N_11674,N_11903);
and U13121 (N_13121,N_12342,N_11960);
or U13122 (N_13122,N_11809,N_11719);
nand U13123 (N_13123,N_11922,N_11898);
or U13124 (N_13124,N_12163,N_11916);
or U13125 (N_13125,N_12194,N_11437);
xnor U13126 (N_13126,N_11292,N_11635);
nand U13127 (N_13127,N_11356,N_11697);
nor U13128 (N_13128,N_12424,N_11347);
and U13129 (N_13129,N_11842,N_12317);
or U13130 (N_13130,N_11377,N_12419);
nor U13131 (N_13131,N_11534,N_11598);
and U13132 (N_13132,N_11581,N_11796);
or U13133 (N_13133,N_11767,N_11444);
and U13134 (N_13134,N_11399,N_11620);
and U13135 (N_13135,N_12074,N_11374);
and U13136 (N_13136,N_12175,N_11971);
nand U13137 (N_13137,N_12147,N_11835);
nor U13138 (N_13138,N_11375,N_12111);
or U13139 (N_13139,N_12249,N_12093);
xnor U13140 (N_13140,N_12235,N_11893);
and U13141 (N_13141,N_11970,N_11862);
xor U13142 (N_13142,N_11433,N_11291);
and U13143 (N_13143,N_11896,N_11479);
nand U13144 (N_13144,N_11530,N_12447);
or U13145 (N_13145,N_11310,N_11401);
or U13146 (N_13146,N_11557,N_11962);
nor U13147 (N_13147,N_11295,N_12478);
and U13148 (N_13148,N_12451,N_12161);
nand U13149 (N_13149,N_11775,N_11916);
and U13150 (N_13150,N_11940,N_12310);
nor U13151 (N_13151,N_11490,N_11655);
nor U13152 (N_13152,N_11522,N_12303);
nor U13153 (N_13153,N_11268,N_12291);
xor U13154 (N_13154,N_11265,N_12309);
xor U13155 (N_13155,N_11775,N_11824);
xor U13156 (N_13156,N_11396,N_12204);
or U13157 (N_13157,N_11470,N_12099);
and U13158 (N_13158,N_11858,N_11745);
or U13159 (N_13159,N_12499,N_11456);
or U13160 (N_13160,N_12472,N_12434);
nor U13161 (N_13161,N_11476,N_11582);
or U13162 (N_13162,N_11434,N_11538);
nand U13163 (N_13163,N_11838,N_11328);
nor U13164 (N_13164,N_12229,N_12185);
and U13165 (N_13165,N_11421,N_12374);
xnor U13166 (N_13166,N_11488,N_11976);
or U13167 (N_13167,N_11441,N_11580);
or U13168 (N_13168,N_12097,N_11755);
nand U13169 (N_13169,N_12024,N_11960);
nand U13170 (N_13170,N_12246,N_12174);
and U13171 (N_13171,N_12499,N_11809);
and U13172 (N_13172,N_11257,N_12224);
or U13173 (N_13173,N_12307,N_11606);
nand U13174 (N_13174,N_11836,N_12430);
and U13175 (N_13175,N_12009,N_12448);
or U13176 (N_13176,N_11996,N_11952);
nor U13177 (N_13177,N_11967,N_11999);
nor U13178 (N_13178,N_11542,N_12261);
nor U13179 (N_13179,N_12403,N_11997);
or U13180 (N_13180,N_12230,N_12082);
nor U13181 (N_13181,N_11762,N_11428);
or U13182 (N_13182,N_12311,N_11772);
nand U13183 (N_13183,N_12387,N_11835);
nor U13184 (N_13184,N_11661,N_12444);
xnor U13185 (N_13185,N_12182,N_11841);
and U13186 (N_13186,N_11408,N_11936);
nor U13187 (N_13187,N_12175,N_11779);
nor U13188 (N_13188,N_11422,N_11795);
nor U13189 (N_13189,N_11966,N_11392);
or U13190 (N_13190,N_12122,N_11489);
nand U13191 (N_13191,N_11977,N_11614);
or U13192 (N_13192,N_11742,N_11357);
or U13193 (N_13193,N_12418,N_12293);
nor U13194 (N_13194,N_11304,N_11349);
xor U13195 (N_13195,N_11963,N_11413);
nand U13196 (N_13196,N_11965,N_11331);
and U13197 (N_13197,N_11840,N_12462);
xnor U13198 (N_13198,N_12084,N_11527);
and U13199 (N_13199,N_11948,N_11477);
nor U13200 (N_13200,N_12155,N_11450);
or U13201 (N_13201,N_12142,N_12052);
and U13202 (N_13202,N_11503,N_11789);
and U13203 (N_13203,N_11412,N_12194);
nand U13204 (N_13204,N_11905,N_11702);
and U13205 (N_13205,N_11330,N_11692);
nor U13206 (N_13206,N_12421,N_12067);
or U13207 (N_13207,N_11998,N_12415);
xor U13208 (N_13208,N_11320,N_11706);
xor U13209 (N_13209,N_11788,N_11267);
and U13210 (N_13210,N_11699,N_11417);
xnor U13211 (N_13211,N_11607,N_11534);
or U13212 (N_13212,N_11302,N_11865);
nand U13213 (N_13213,N_11987,N_11667);
or U13214 (N_13214,N_11924,N_11441);
nor U13215 (N_13215,N_11926,N_12252);
or U13216 (N_13216,N_11301,N_12130);
or U13217 (N_13217,N_11692,N_12454);
nor U13218 (N_13218,N_11789,N_11274);
xor U13219 (N_13219,N_12432,N_11891);
and U13220 (N_13220,N_11682,N_11916);
or U13221 (N_13221,N_11483,N_11801);
or U13222 (N_13222,N_12023,N_11403);
nor U13223 (N_13223,N_11312,N_12456);
and U13224 (N_13224,N_12374,N_12434);
or U13225 (N_13225,N_12007,N_12452);
nor U13226 (N_13226,N_12405,N_12236);
and U13227 (N_13227,N_11610,N_11330);
and U13228 (N_13228,N_12164,N_12055);
and U13229 (N_13229,N_11761,N_12492);
xnor U13230 (N_13230,N_12009,N_12497);
nor U13231 (N_13231,N_12453,N_12387);
nand U13232 (N_13232,N_12486,N_11996);
nor U13233 (N_13233,N_11307,N_11327);
xnor U13234 (N_13234,N_11522,N_12086);
and U13235 (N_13235,N_11317,N_11694);
nand U13236 (N_13236,N_12377,N_12480);
and U13237 (N_13237,N_12314,N_11549);
or U13238 (N_13238,N_12062,N_11267);
and U13239 (N_13239,N_12331,N_12361);
nand U13240 (N_13240,N_11273,N_11282);
and U13241 (N_13241,N_11531,N_12251);
nor U13242 (N_13242,N_12157,N_12426);
nor U13243 (N_13243,N_11916,N_12369);
nand U13244 (N_13244,N_12255,N_12491);
nor U13245 (N_13245,N_12263,N_12410);
nand U13246 (N_13246,N_11597,N_11374);
or U13247 (N_13247,N_12264,N_12166);
xor U13248 (N_13248,N_12155,N_11884);
or U13249 (N_13249,N_12383,N_11808);
nor U13250 (N_13250,N_12136,N_12416);
xor U13251 (N_13251,N_12357,N_12025);
nand U13252 (N_13252,N_12293,N_11959);
xor U13253 (N_13253,N_11646,N_11913);
and U13254 (N_13254,N_11669,N_11942);
nor U13255 (N_13255,N_11428,N_11893);
and U13256 (N_13256,N_11534,N_11511);
xnor U13257 (N_13257,N_11724,N_11445);
and U13258 (N_13258,N_11629,N_11835);
and U13259 (N_13259,N_12351,N_12378);
nor U13260 (N_13260,N_12264,N_11439);
nand U13261 (N_13261,N_11645,N_11646);
nor U13262 (N_13262,N_11423,N_11700);
nor U13263 (N_13263,N_12043,N_11762);
and U13264 (N_13264,N_12370,N_11320);
nand U13265 (N_13265,N_11469,N_11468);
and U13266 (N_13266,N_12176,N_11318);
or U13267 (N_13267,N_11977,N_11929);
xor U13268 (N_13268,N_12241,N_12162);
nand U13269 (N_13269,N_12059,N_12425);
nand U13270 (N_13270,N_11576,N_11297);
nand U13271 (N_13271,N_12219,N_11628);
xnor U13272 (N_13272,N_11816,N_12160);
or U13273 (N_13273,N_11836,N_11805);
nand U13274 (N_13274,N_11682,N_11406);
xor U13275 (N_13275,N_11604,N_11529);
and U13276 (N_13276,N_12102,N_12436);
or U13277 (N_13277,N_11435,N_12290);
nand U13278 (N_13278,N_11447,N_12261);
nand U13279 (N_13279,N_11406,N_11929);
nor U13280 (N_13280,N_12146,N_11681);
and U13281 (N_13281,N_12342,N_12353);
or U13282 (N_13282,N_11287,N_11289);
nand U13283 (N_13283,N_11365,N_11778);
and U13284 (N_13284,N_11921,N_12241);
nand U13285 (N_13285,N_12055,N_11618);
nand U13286 (N_13286,N_12140,N_12436);
nor U13287 (N_13287,N_12027,N_11747);
nand U13288 (N_13288,N_11969,N_11414);
nor U13289 (N_13289,N_11296,N_12441);
or U13290 (N_13290,N_11294,N_11625);
xnor U13291 (N_13291,N_12184,N_11270);
or U13292 (N_13292,N_11519,N_12356);
nand U13293 (N_13293,N_11747,N_12227);
or U13294 (N_13294,N_12425,N_11636);
or U13295 (N_13295,N_12047,N_11341);
or U13296 (N_13296,N_11398,N_11993);
nand U13297 (N_13297,N_11971,N_11892);
nand U13298 (N_13298,N_12279,N_12203);
or U13299 (N_13299,N_11965,N_11773);
xnor U13300 (N_13300,N_11872,N_12212);
and U13301 (N_13301,N_11809,N_11397);
xor U13302 (N_13302,N_12212,N_11426);
nor U13303 (N_13303,N_11648,N_12024);
nor U13304 (N_13304,N_11286,N_12443);
xor U13305 (N_13305,N_12093,N_11741);
xnor U13306 (N_13306,N_12028,N_11758);
nor U13307 (N_13307,N_11355,N_11650);
xnor U13308 (N_13308,N_12085,N_11706);
or U13309 (N_13309,N_12033,N_11954);
or U13310 (N_13310,N_11775,N_11953);
nor U13311 (N_13311,N_11719,N_11412);
or U13312 (N_13312,N_11776,N_11981);
xnor U13313 (N_13313,N_11876,N_12332);
or U13314 (N_13314,N_11936,N_12276);
xnor U13315 (N_13315,N_11333,N_12037);
and U13316 (N_13316,N_12287,N_12164);
and U13317 (N_13317,N_11777,N_11346);
xor U13318 (N_13318,N_11332,N_12258);
nor U13319 (N_13319,N_12363,N_12264);
xnor U13320 (N_13320,N_11666,N_11567);
nand U13321 (N_13321,N_11635,N_11944);
or U13322 (N_13322,N_11457,N_11884);
nor U13323 (N_13323,N_11525,N_12044);
xnor U13324 (N_13324,N_11694,N_11853);
nor U13325 (N_13325,N_12218,N_11574);
nor U13326 (N_13326,N_12180,N_12261);
nand U13327 (N_13327,N_12133,N_12269);
or U13328 (N_13328,N_11655,N_11639);
nor U13329 (N_13329,N_12499,N_12311);
xnor U13330 (N_13330,N_12449,N_12428);
xnor U13331 (N_13331,N_12476,N_12169);
nor U13332 (N_13332,N_12431,N_11983);
and U13333 (N_13333,N_11651,N_12045);
nand U13334 (N_13334,N_11940,N_11319);
nand U13335 (N_13335,N_11450,N_11899);
nor U13336 (N_13336,N_11862,N_11994);
or U13337 (N_13337,N_11284,N_11530);
and U13338 (N_13338,N_11754,N_12170);
or U13339 (N_13339,N_11836,N_11445);
xnor U13340 (N_13340,N_11354,N_12248);
nand U13341 (N_13341,N_12462,N_11511);
or U13342 (N_13342,N_12223,N_11711);
and U13343 (N_13343,N_11794,N_12289);
and U13344 (N_13344,N_12493,N_12451);
nand U13345 (N_13345,N_12111,N_11736);
nor U13346 (N_13346,N_11753,N_11342);
or U13347 (N_13347,N_12091,N_12286);
nand U13348 (N_13348,N_11643,N_11849);
nand U13349 (N_13349,N_11751,N_11649);
nand U13350 (N_13350,N_11433,N_12475);
or U13351 (N_13351,N_11262,N_11475);
or U13352 (N_13352,N_12147,N_12362);
xor U13353 (N_13353,N_11528,N_11908);
nor U13354 (N_13354,N_11782,N_11704);
or U13355 (N_13355,N_12397,N_12037);
or U13356 (N_13356,N_11649,N_11484);
nand U13357 (N_13357,N_12282,N_12148);
and U13358 (N_13358,N_11445,N_11814);
and U13359 (N_13359,N_11922,N_11693);
or U13360 (N_13360,N_12008,N_12238);
xor U13361 (N_13361,N_12118,N_11800);
nand U13362 (N_13362,N_11901,N_12097);
nand U13363 (N_13363,N_11693,N_11753);
xnor U13364 (N_13364,N_12244,N_12032);
and U13365 (N_13365,N_12321,N_11849);
and U13366 (N_13366,N_11399,N_12329);
nor U13367 (N_13367,N_12491,N_12452);
and U13368 (N_13368,N_12141,N_11441);
nor U13369 (N_13369,N_12176,N_11783);
nand U13370 (N_13370,N_12323,N_12120);
and U13371 (N_13371,N_11455,N_11725);
and U13372 (N_13372,N_11436,N_11762);
nor U13373 (N_13373,N_11777,N_12225);
nand U13374 (N_13374,N_11762,N_11508);
nor U13375 (N_13375,N_11796,N_11888);
nand U13376 (N_13376,N_12149,N_12191);
nor U13377 (N_13377,N_11448,N_12067);
or U13378 (N_13378,N_12194,N_12117);
nor U13379 (N_13379,N_11798,N_11428);
or U13380 (N_13380,N_11700,N_12325);
nand U13381 (N_13381,N_12432,N_11832);
xnor U13382 (N_13382,N_12135,N_12298);
and U13383 (N_13383,N_12182,N_11935);
nor U13384 (N_13384,N_11974,N_12335);
xnor U13385 (N_13385,N_12216,N_12038);
or U13386 (N_13386,N_11790,N_11874);
nor U13387 (N_13387,N_12417,N_12080);
nor U13388 (N_13388,N_11711,N_11898);
nand U13389 (N_13389,N_11489,N_11900);
or U13390 (N_13390,N_12101,N_11773);
xnor U13391 (N_13391,N_11932,N_11275);
or U13392 (N_13392,N_11564,N_12367);
nand U13393 (N_13393,N_11281,N_12053);
nand U13394 (N_13394,N_11821,N_12427);
and U13395 (N_13395,N_12360,N_12436);
xnor U13396 (N_13396,N_11391,N_12167);
or U13397 (N_13397,N_12085,N_11335);
nor U13398 (N_13398,N_11545,N_11519);
nand U13399 (N_13399,N_12229,N_12476);
or U13400 (N_13400,N_11853,N_12395);
and U13401 (N_13401,N_11646,N_11515);
xnor U13402 (N_13402,N_12444,N_12150);
or U13403 (N_13403,N_11868,N_11774);
and U13404 (N_13404,N_11538,N_12350);
nor U13405 (N_13405,N_12268,N_11884);
xnor U13406 (N_13406,N_12468,N_11309);
and U13407 (N_13407,N_11359,N_11299);
or U13408 (N_13408,N_11707,N_11835);
xor U13409 (N_13409,N_11420,N_11288);
xnor U13410 (N_13410,N_12280,N_11499);
and U13411 (N_13411,N_11338,N_12369);
nor U13412 (N_13412,N_11982,N_12237);
nand U13413 (N_13413,N_12012,N_12313);
or U13414 (N_13414,N_11564,N_11940);
xnor U13415 (N_13415,N_11334,N_12323);
nor U13416 (N_13416,N_12336,N_11669);
nor U13417 (N_13417,N_12178,N_11457);
and U13418 (N_13418,N_12365,N_11657);
or U13419 (N_13419,N_11297,N_12179);
and U13420 (N_13420,N_12403,N_11270);
xnor U13421 (N_13421,N_11572,N_12054);
and U13422 (N_13422,N_11863,N_11530);
xor U13423 (N_13423,N_11792,N_11885);
xor U13424 (N_13424,N_11654,N_11738);
xor U13425 (N_13425,N_12257,N_12057);
xor U13426 (N_13426,N_11727,N_11495);
nand U13427 (N_13427,N_11719,N_11794);
nand U13428 (N_13428,N_12122,N_11990);
or U13429 (N_13429,N_12441,N_11401);
or U13430 (N_13430,N_11344,N_11637);
xnor U13431 (N_13431,N_11751,N_12102);
nand U13432 (N_13432,N_11612,N_12107);
nor U13433 (N_13433,N_11705,N_12466);
nor U13434 (N_13434,N_11669,N_12312);
nor U13435 (N_13435,N_11553,N_12145);
nor U13436 (N_13436,N_12294,N_12050);
xnor U13437 (N_13437,N_11405,N_11811);
or U13438 (N_13438,N_12406,N_12373);
or U13439 (N_13439,N_11976,N_11300);
and U13440 (N_13440,N_11752,N_12433);
nand U13441 (N_13441,N_11894,N_11621);
and U13442 (N_13442,N_11749,N_12067);
and U13443 (N_13443,N_12169,N_11759);
xor U13444 (N_13444,N_12196,N_11761);
nand U13445 (N_13445,N_12236,N_11869);
and U13446 (N_13446,N_11300,N_12372);
and U13447 (N_13447,N_11526,N_11893);
nand U13448 (N_13448,N_11977,N_11350);
nand U13449 (N_13449,N_11652,N_11839);
nor U13450 (N_13450,N_11497,N_12331);
xor U13451 (N_13451,N_12377,N_12217);
nand U13452 (N_13452,N_11252,N_11821);
nand U13453 (N_13453,N_12026,N_11264);
xnor U13454 (N_13454,N_11851,N_11664);
or U13455 (N_13455,N_11687,N_11638);
nor U13456 (N_13456,N_11775,N_11299);
xnor U13457 (N_13457,N_12478,N_12096);
nand U13458 (N_13458,N_11762,N_12387);
nor U13459 (N_13459,N_12483,N_11363);
nand U13460 (N_13460,N_11446,N_11950);
nand U13461 (N_13461,N_11524,N_12314);
nand U13462 (N_13462,N_12350,N_11698);
xnor U13463 (N_13463,N_11816,N_11796);
and U13464 (N_13464,N_11541,N_11858);
and U13465 (N_13465,N_12080,N_12045);
xnor U13466 (N_13466,N_11971,N_12448);
and U13467 (N_13467,N_12335,N_11272);
or U13468 (N_13468,N_12065,N_11354);
xnor U13469 (N_13469,N_11525,N_11425);
or U13470 (N_13470,N_12165,N_11960);
nor U13471 (N_13471,N_11317,N_11350);
and U13472 (N_13472,N_11954,N_12394);
xor U13473 (N_13473,N_12413,N_11487);
nor U13474 (N_13474,N_12082,N_12263);
xnor U13475 (N_13475,N_12199,N_11683);
nand U13476 (N_13476,N_11909,N_12436);
xnor U13477 (N_13477,N_11550,N_11791);
or U13478 (N_13478,N_11889,N_11291);
nand U13479 (N_13479,N_11320,N_12440);
xor U13480 (N_13480,N_11854,N_11451);
or U13481 (N_13481,N_12176,N_11439);
xnor U13482 (N_13482,N_11755,N_11901);
xnor U13483 (N_13483,N_11541,N_11614);
nand U13484 (N_13484,N_11968,N_12082);
and U13485 (N_13485,N_12327,N_11725);
and U13486 (N_13486,N_12125,N_11929);
xnor U13487 (N_13487,N_11998,N_11478);
and U13488 (N_13488,N_12388,N_11756);
and U13489 (N_13489,N_12344,N_11804);
xnor U13490 (N_13490,N_11802,N_12349);
or U13491 (N_13491,N_11664,N_11270);
nor U13492 (N_13492,N_11358,N_11340);
xor U13493 (N_13493,N_11703,N_11692);
and U13494 (N_13494,N_11678,N_11938);
nor U13495 (N_13495,N_11808,N_11801);
and U13496 (N_13496,N_12448,N_11649);
or U13497 (N_13497,N_12083,N_11251);
nand U13498 (N_13498,N_11329,N_11563);
xor U13499 (N_13499,N_12136,N_11899);
xor U13500 (N_13500,N_12121,N_12211);
nand U13501 (N_13501,N_12206,N_12289);
nand U13502 (N_13502,N_12014,N_12156);
nand U13503 (N_13503,N_12131,N_12398);
nor U13504 (N_13504,N_11714,N_11571);
nor U13505 (N_13505,N_12203,N_11736);
or U13506 (N_13506,N_11748,N_12042);
nand U13507 (N_13507,N_12182,N_11631);
xnor U13508 (N_13508,N_11409,N_12490);
xor U13509 (N_13509,N_11999,N_12349);
nor U13510 (N_13510,N_11783,N_11506);
and U13511 (N_13511,N_11861,N_11255);
xor U13512 (N_13512,N_12171,N_12115);
nor U13513 (N_13513,N_11782,N_11819);
nand U13514 (N_13514,N_12498,N_11816);
xnor U13515 (N_13515,N_12164,N_11713);
nand U13516 (N_13516,N_11974,N_11367);
xor U13517 (N_13517,N_11479,N_12034);
xor U13518 (N_13518,N_12272,N_11393);
and U13519 (N_13519,N_12012,N_11469);
xor U13520 (N_13520,N_12426,N_12383);
nand U13521 (N_13521,N_12023,N_11672);
xor U13522 (N_13522,N_11955,N_12438);
xnor U13523 (N_13523,N_11309,N_11888);
nor U13524 (N_13524,N_12185,N_11866);
and U13525 (N_13525,N_11872,N_12336);
xnor U13526 (N_13526,N_11253,N_12088);
and U13527 (N_13527,N_11511,N_12177);
xor U13528 (N_13528,N_11955,N_11671);
nand U13529 (N_13529,N_11763,N_12469);
or U13530 (N_13530,N_11585,N_11349);
or U13531 (N_13531,N_12495,N_12484);
xor U13532 (N_13532,N_12152,N_12025);
or U13533 (N_13533,N_11452,N_11375);
nand U13534 (N_13534,N_11441,N_11928);
xor U13535 (N_13535,N_11868,N_11659);
nand U13536 (N_13536,N_11508,N_11537);
and U13537 (N_13537,N_11897,N_11340);
nor U13538 (N_13538,N_11971,N_12000);
and U13539 (N_13539,N_11731,N_11632);
nand U13540 (N_13540,N_11503,N_12054);
nor U13541 (N_13541,N_11442,N_11593);
nand U13542 (N_13542,N_11701,N_12170);
nor U13543 (N_13543,N_11357,N_11913);
and U13544 (N_13544,N_11583,N_12157);
or U13545 (N_13545,N_11676,N_11925);
and U13546 (N_13546,N_11356,N_12161);
nor U13547 (N_13547,N_11536,N_11504);
nor U13548 (N_13548,N_11851,N_12386);
nand U13549 (N_13549,N_11406,N_11957);
and U13550 (N_13550,N_11678,N_11543);
xor U13551 (N_13551,N_12318,N_11964);
nand U13552 (N_13552,N_12205,N_12397);
or U13553 (N_13553,N_12413,N_11253);
or U13554 (N_13554,N_12328,N_12034);
or U13555 (N_13555,N_11818,N_11377);
nor U13556 (N_13556,N_11546,N_11259);
and U13557 (N_13557,N_12077,N_11838);
and U13558 (N_13558,N_11697,N_12208);
nor U13559 (N_13559,N_11736,N_11679);
or U13560 (N_13560,N_11384,N_12002);
nor U13561 (N_13561,N_11526,N_11811);
nor U13562 (N_13562,N_12172,N_11406);
and U13563 (N_13563,N_12059,N_12190);
xnor U13564 (N_13564,N_12377,N_11742);
and U13565 (N_13565,N_12045,N_12372);
or U13566 (N_13566,N_11836,N_12428);
xnor U13567 (N_13567,N_11919,N_12238);
or U13568 (N_13568,N_11440,N_11782);
nor U13569 (N_13569,N_12303,N_11954);
xnor U13570 (N_13570,N_11359,N_11418);
or U13571 (N_13571,N_12095,N_12284);
xor U13572 (N_13572,N_12162,N_12309);
nor U13573 (N_13573,N_11852,N_12316);
and U13574 (N_13574,N_11842,N_11827);
and U13575 (N_13575,N_11793,N_11462);
nor U13576 (N_13576,N_11572,N_12091);
nand U13577 (N_13577,N_12111,N_12265);
or U13578 (N_13578,N_11580,N_11644);
and U13579 (N_13579,N_12025,N_12486);
and U13580 (N_13580,N_12411,N_11549);
or U13581 (N_13581,N_11354,N_11570);
or U13582 (N_13582,N_11645,N_12388);
nand U13583 (N_13583,N_12479,N_12214);
xor U13584 (N_13584,N_11274,N_12109);
or U13585 (N_13585,N_11741,N_11815);
xor U13586 (N_13586,N_12198,N_12172);
and U13587 (N_13587,N_12434,N_12427);
xor U13588 (N_13588,N_11707,N_12101);
nor U13589 (N_13589,N_12413,N_12459);
xor U13590 (N_13590,N_11267,N_11936);
nor U13591 (N_13591,N_12132,N_12177);
nand U13592 (N_13592,N_11844,N_11674);
nand U13593 (N_13593,N_11504,N_11272);
xnor U13594 (N_13594,N_11975,N_11956);
or U13595 (N_13595,N_11839,N_12013);
xor U13596 (N_13596,N_12096,N_11856);
and U13597 (N_13597,N_11668,N_11868);
xnor U13598 (N_13598,N_12119,N_11675);
xor U13599 (N_13599,N_11541,N_11655);
and U13600 (N_13600,N_11338,N_11727);
nand U13601 (N_13601,N_12141,N_11514);
or U13602 (N_13602,N_11790,N_11567);
nand U13603 (N_13603,N_11835,N_11938);
or U13604 (N_13604,N_12365,N_11469);
xor U13605 (N_13605,N_11626,N_12247);
xnor U13606 (N_13606,N_12166,N_12102);
or U13607 (N_13607,N_12416,N_12364);
nor U13608 (N_13608,N_11296,N_12301);
nand U13609 (N_13609,N_12168,N_12379);
nor U13610 (N_13610,N_12129,N_11476);
nor U13611 (N_13611,N_11256,N_12438);
and U13612 (N_13612,N_11640,N_12318);
nor U13613 (N_13613,N_11877,N_11764);
and U13614 (N_13614,N_11952,N_11328);
xor U13615 (N_13615,N_12273,N_11676);
nor U13616 (N_13616,N_11765,N_11297);
nor U13617 (N_13617,N_12134,N_11950);
xnor U13618 (N_13618,N_12423,N_11329);
xnor U13619 (N_13619,N_11990,N_11598);
nand U13620 (N_13620,N_11782,N_11269);
and U13621 (N_13621,N_12067,N_12290);
or U13622 (N_13622,N_12465,N_12391);
xnor U13623 (N_13623,N_12494,N_11761);
xnor U13624 (N_13624,N_11919,N_12470);
or U13625 (N_13625,N_11367,N_11595);
xor U13626 (N_13626,N_11792,N_12220);
or U13627 (N_13627,N_12271,N_12498);
nand U13628 (N_13628,N_11586,N_12360);
and U13629 (N_13629,N_11678,N_12428);
and U13630 (N_13630,N_12453,N_12338);
nor U13631 (N_13631,N_12490,N_11275);
xor U13632 (N_13632,N_12008,N_11273);
and U13633 (N_13633,N_11734,N_11794);
and U13634 (N_13634,N_12170,N_12130);
xor U13635 (N_13635,N_12168,N_11461);
nor U13636 (N_13636,N_11804,N_12416);
nand U13637 (N_13637,N_11875,N_11680);
xor U13638 (N_13638,N_11617,N_11673);
nand U13639 (N_13639,N_12464,N_11952);
nor U13640 (N_13640,N_12079,N_11720);
and U13641 (N_13641,N_11614,N_11443);
or U13642 (N_13642,N_11313,N_11709);
nor U13643 (N_13643,N_11628,N_11287);
xnor U13644 (N_13644,N_11406,N_12454);
xor U13645 (N_13645,N_11473,N_11450);
xnor U13646 (N_13646,N_12423,N_11949);
or U13647 (N_13647,N_11471,N_11375);
and U13648 (N_13648,N_11784,N_12329);
and U13649 (N_13649,N_11641,N_11350);
nand U13650 (N_13650,N_11683,N_11714);
or U13651 (N_13651,N_11850,N_11426);
nor U13652 (N_13652,N_12374,N_11515);
and U13653 (N_13653,N_12014,N_11499);
and U13654 (N_13654,N_11541,N_12081);
xor U13655 (N_13655,N_12174,N_11768);
or U13656 (N_13656,N_12113,N_11964);
nor U13657 (N_13657,N_12221,N_11566);
nand U13658 (N_13658,N_12285,N_11602);
and U13659 (N_13659,N_12047,N_12140);
xnor U13660 (N_13660,N_12340,N_11884);
xor U13661 (N_13661,N_12446,N_12245);
xor U13662 (N_13662,N_12138,N_12031);
xnor U13663 (N_13663,N_11394,N_12271);
nor U13664 (N_13664,N_11703,N_11334);
xnor U13665 (N_13665,N_11292,N_11821);
nor U13666 (N_13666,N_11793,N_11742);
nor U13667 (N_13667,N_11762,N_12011);
nor U13668 (N_13668,N_12432,N_11534);
or U13669 (N_13669,N_11449,N_11741);
nand U13670 (N_13670,N_11966,N_12139);
xnor U13671 (N_13671,N_12269,N_11395);
xor U13672 (N_13672,N_12347,N_11400);
xor U13673 (N_13673,N_12280,N_12311);
or U13674 (N_13674,N_11767,N_12219);
nand U13675 (N_13675,N_12111,N_12256);
or U13676 (N_13676,N_11443,N_12257);
and U13677 (N_13677,N_12378,N_11728);
or U13678 (N_13678,N_12374,N_12011);
nand U13679 (N_13679,N_11263,N_11778);
and U13680 (N_13680,N_11532,N_11287);
and U13681 (N_13681,N_12010,N_11635);
or U13682 (N_13682,N_11566,N_12365);
nand U13683 (N_13683,N_11925,N_11937);
xnor U13684 (N_13684,N_12030,N_11514);
nor U13685 (N_13685,N_11910,N_11786);
nand U13686 (N_13686,N_12064,N_11610);
nor U13687 (N_13687,N_12214,N_11390);
and U13688 (N_13688,N_11880,N_11534);
xor U13689 (N_13689,N_12024,N_12274);
and U13690 (N_13690,N_11661,N_11479);
nor U13691 (N_13691,N_12328,N_11483);
nor U13692 (N_13692,N_12159,N_12452);
xnor U13693 (N_13693,N_11784,N_12411);
or U13694 (N_13694,N_11590,N_11421);
and U13695 (N_13695,N_11255,N_11694);
nor U13696 (N_13696,N_11732,N_11686);
and U13697 (N_13697,N_12240,N_11604);
or U13698 (N_13698,N_11621,N_12138);
nand U13699 (N_13699,N_12195,N_11779);
xnor U13700 (N_13700,N_12224,N_12002);
nor U13701 (N_13701,N_11444,N_12093);
nand U13702 (N_13702,N_12469,N_11765);
nand U13703 (N_13703,N_11645,N_12478);
or U13704 (N_13704,N_11741,N_12475);
nor U13705 (N_13705,N_11415,N_12215);
and U13706 (N_13706,N_12407,N_11557);
or U13707 (N_13707,N_12127,N_11682);
or U13708 (N_13708,N_12357,N_12218);
and U13709 (N_13709,N_12463,N_11643);
or U13710 (N_13710,N_12412,N_11682);
nand U13711 (N_13711,N_12452,N_11676);
or U13712 (N_13712,N_12177,N_12299);
nand U13713 (N_13713,N_11671,N_11977);
or U13714 (N_13714,N_12384,N_11659);
nor U13715 (N_13715,N_12154,N_12114);
and U13716 (N_13716,N_11662,N_12414);
nand U13717 (N_13717,N_12448,N_11742);
nand U13718 (N_13718,N_11255,N_12060);
xor U13719 (N_13719,N_11383,N_12283);
and U13720 (N_13720,N_11720,N_12240);
nand U13721 (N_13721,N_12213,N_11566);
nor U13722 (N_13722,N_11485,N_11338);
and U13723 (N_13723,N_11472,N_11987);
or U13724 (N_13724,N_11667,N_11578);
xor U13725 (N_13725,N_11878,N_11385);
nand U13726 (N_13726,N_12338,N_12358);
nand U13727 (N_13727,N_11693,N_12231);
xor U13728 (N_13728,N_12219,N_11424);
nor U13729 (N_13729,N_11578,N_12302);
or U13730 (N_13730,N_11667,N_12387);
nand U13731 (N_13731,N_11335,N_11489);
xor U13732 (N_13732,N_11680,N_11502);
nand U13733 (N_13733,N_12326,N_11333);
and U13734 (N_13734,N_11366,N_11469);
nor U13735 (N_13735,N_12144,N_12174);
xor U13736 (N_13736,N_12241,N_11614);
and U13737 (N_13737,N_11355,N_11859);
or U13738 (N_13738,N_11884,N_11923);
and U13739 (N_13739,N_11796,N_12158);
or U13740 (N_13740,N_11412,N_11764);
or U13741 (N_13741,N_11328,N_12033);
nor U13742 (N_13742,N_12077,N_11262);
xor U13743 (N_13743,N_12472,N_12423);
nor U13744 (N_13744,N_11442,N_12214);
nand U13745 (N_13745,N_11606,N_12135);
nor U13746 (N_13746,N_11690,N_11680);
nand U13747 (N_13747,N_12081,N_12489);
xor U13748 (N_13748,N_12332,N_11468);
and U13749 (N_13749,N_11990,N_11492);
or U13750 (N_13750,N_13269,N_12613);
nand U13751 (N_13751,N_12539,N_12866);
nand U13752 (N_13752,N_12808,N_13296);
xor U13753 (N_13753,N_13081,N_12833);
nor U13754 (N_13754,N_13365,N_12627);
and U13755 (N_13755,N_13682,N_12628);
xor U13756 (N_13756,N_13714,N_13724);
nand U13757 (N_13757,N_12590,N_12797);
nor U13758 (N_13758,N_12793,N_13194);
nand U13759 (N_13759,N_13693,N_13143);
xor U13760 (N_13760,N_13610,N_13174);
xor U13761 (N_13761,N_13014,N_13469);
xor U13762 (N_13762,N_13036,N_13543);
nand U13763 (N_13763,N_13115,N_12982);
xnor U13764 (N_13764,N_12665,N_12922);
or U13765 (N_13765,N_13352,N_13214);
nor U13766 (N_13766,N_12563,N_13116);
or U13767 (N_13767,N_13330,N_12557);
xor U13768 (N_13768,N_13519,N_13191);
or U13769 (N_13769,N_12689,N_13247);
and U13770 (N_13770,N_12946,N_13332);
and U13771 (N_13771,N_12556,N_13155);
nand U13772 (N_13772,N_13746,N_13413);
xnor U13773 (N_13773,N_12779,N_12679);
and U13774 (N_13774,N_13104,N_13311);
or U13775 (N_13775,N_13376,N_12515);
nor U13776 (N_13776,N_12669,N_12681);
and U13777 (N_13777,N_13454,N_13465);
xor U13778 (N_13778,N_12514,N_12545);
nor U13779 (N_13779,N_13007,N_12636);
nor U13780 (N_13780,N_13207,N_13414);
and U13781 (N_13781,N_13430,N_13442);
nor U13782 (N_13782,N_13696,N_12710);
and U13783 (N_13783,N_13704,N_13225);
nor U13784 (N_13784,N_12703,N_13466);
or U13785 (N_13785,N_12874,N_12610);
and U13786 (N_13786,N_13112,N_13148);
nor U13787 (N_13787,N_12961,N_13222);
and U13788 (N_13788,N_13158,N_12687);
xnor U13789 (N_13789,N_13183,N_13522);
nor U13790 (N_13790,N_13179,N_13651);
or U13791 (N_13791,N_13662,N_13310);
nor U13792 (N_13792,N_12912,N_13118);
xor U13793 (N_13793,N_12648,N_12646);
xor U13794 (N_13794,N_13653,N_13151);
nor U13795 (N_13795,N_12993,N_13540);
nand U13796 (N_13796,N_12644,N_13507);
xnor U13797 (N_13797,N_13274,N_12976);
xnor U13798 (N_13798,N_12879,N_12815);
and U13799 (N_13799,N_13588,N_13425);
nor U13800 (N_13800,N_13452,N_13495);
or U13801 (N_13801,N_13100,N_12668);
xor U13802 (N_13802,N_12920,N_13170);
nor U13803 (N_13803,N_13114,N_12738);
nand U13804 (N_13804,N_13068,N_12770);
or U13805 (N_13805,N_12864,N_13498);
nor U13806 (N_13806,N_12894,N_13153);
or U13807 (N_13807,N_13636,N_13339);
or U13808 (N_13808,N_13031,N_12881);
nand U13809 (N_13809,N_12754,N_12761);
nor U13810 (N_13810,N_13666,N_13131);
nand U13811 (N_13811,N_13694,N_13345);
nor U13812 (N_13812,N_13494,N_13475);
and U13813 (N_13813,N_13444,N_13085);
nor U13814 (N_13814,N_12573,N_13009);
xor U13815 (N_13815,N_12861,N_12649);
or U13816 (N_13816,N_13661,N_13152);
and U13817 (N_13817,N_13370,N_12849);
nor U13818 (N_13818,N_12705,N_13154);
xnor U13819 (N_13819,N_13595,N_13175);
and U13820 (N_13820,N_13450,N_12672);
and U13821 (N_13821,N_12870,N_13373);
nor U13822 (N_13822,N_12596,N_13099);
nand U13823 (N_13823,N_13052,N_13263);
xnor U13824 (N_13824,N_13398,N_13057);
or U13825 (N_13825,N_12571,N_13568);
or U13826 (N_13826,N_13573,N_12535);
nand U13827 (N_13827,N_12530,N_13002);
xnor U13828 (N_13828,N_12749,N_12823);
nand U13829 (N_13829,N_13602,N_13429);
nand U13830 (N_13830,N_13200,N_13576);
xor U13831 (N_13831,N_12900,N_12843);
nor U13832 (N_13832,N_13280,N_13501);
or U13833 (N_13833,N_13678,N_12811);
or U13834 (N_13834,N_13688,N_13043);
xnor U13835 (N_13835,N_13729,N_13403);
and U13836 (N_13836,N_13064,N_12734);
and U13837 (N_13837,N_12686,N_12730);
nor U13838 (N_13838,N_13410,N_13532);
nand U13839 (N_13839,N_13448,N_12683);
nor U13840 (N_13840,N_12847,N_13394);
xnor U13841 (N_13841,N_13087,N_13472);
nand U13842 (N_13842,N_13545,N_13333);
nor U13843 (N_13843,N_13667,N_13005);
and U13844 (N_13844,N_12972,N_13010);
nand U13845 (N_13845,N_12570,N_13203);
and U13846 (N_13846,N_13301,N_13416);
nor U13847 (N_13847,N_13074,N_12898);
xnor U13848 (N_13848,N_12549,N_13259);
xnor U13849 (N_13849,N_13205,N_13526);
nor U13850 (N_13850,N_13421,N_13531);
and U13851 (N_13851,N_13379,N_12918);
or U13852 (N_13852,N_13125,N_13627);
and U13853 (N_13853,N_13435,N_13169);
nor U13854 (N_13854,N_13298,N_13220);
or U13855 (N_13855,N_12618,N_13338);
nor U13856 (N_13856,N_13592,N_12924);
and U13857 (N_13857,N_13715,N_13309);
nand U13858 (N_13858,N_12830,N_12653);
xor U13859 (N_13859,N_12896,N_12954);
nand U13860 (N_13860,N_13490,N_12939);
nor U13861 (N_13861,N_13348,N_13385);
nand U13862 (N_13862,N_12914,N_12597);
and U13863 (N_13863,N_13483,N_13464);
xnor U13864 (N_13864,N_12625,N_13571);
and U13865 (N_13865,N_12521,N_13607);
and U13866 (N_13866,N_12842,N_12566);
nand U13867 (N_13867,N_13659,N_13184);
nand U13868 (N_13868,N_13146,N_13686);
nor U13869 (N_13869,N_13658,N_13008);
and U13870 (N_13870,N_13614,N_13334);
nand U13871 (N_13871,N_13648,N_13700);
nor U13872 (N_13872,N_12675,N_13198);
or U13873 (N_13873,N_13268,N_12587);
or U13874 (N_13874,N_13489,N_12561);
or U13875 (N_13875,N_13281,N_13147);
nor U13876 (N_13876,N_13423,N_13053);
or U13877 (N_13877,N_13605,N_13529);
xnor U13878 (N_13878,N_12763,N_12949);
nor U13879 (N_13879,N_13219,N_12887);
xor U13880 (N_13880,N_13020,N_13178);
and U13881 (N_13881,N_13077,N_12805);
xor U13882 (N_13882,N_12759,N_13091);
xnor U13883 (N_13883,N_13628,N_12747);
and U13884 (N_13884,N_13477,N_13652);
and U13885 (N_13885,N_13633,N_12764);
nor U13886 (N_13886,N_12586,N_13502);
xnor U13887 (N_13887,N_13242,N_12929);
nand U13888 (N_13888,N_13739,N_13346);
and U13889 (N_13889,N_13092,N_13608);
or U13890 (N_13890,N_12725,N_13341);
nand U13891 (N_13891,N_13082,N_13166);
xor U13892 (N_13892,N_13692,N_13024);
or U13893 (N_13893,N_12917,N_13030);
and U13894 (N_13894,N_12776,N_12777);
nand U13895 (N_13895,N_12877,N_13625);
xor U13896 (N_13896,N_13051,N_13336);
nand U13897 (N_13897,N_13725,N_13720);
nand U13898 (N_13898,N_12554,N_13418);
nand U13899 (N_13899,N_13749,N_12718);
nor U13900 (N_13900,N_13355,N_12869);
or U13901 (N_13901,N_13375,N_13619);
or U13902 (N_13902,N_12771,N_13037);
or U13903 (N_13903,N_12934,N_12603);
nand U13904 (N_13904,N_13378,N_13664);
and U13905 (N_13905,N_12731,N_12907);
and U13906 (N_13906,N_13655,N_13171);
or U13907 (N_13907,N_13478,N_13236);
nor U13908 (N_13908,N_12943,N_13457);
xnor U13909 (N_13909,N_13596,N_13270);
nand U13910 (N_13910,N_13362,N_13730);
xor U13911 (N_13911,N_13606,N_13387);
nand U13912 (N_13912,N_12757,N_12723);
nor U13913 (N_13913,N_12816,N_13539);
or U13914 (N_13914,N_13510,N_13535);
nand U13915 (N_13915,N_13572,N_13071);
or U13916 (N_13916,N_13109,N_13580);
nor U13917 (N_13917,N_13359,N_13491);
xnor U13918 (N_13918,N_12517,N_13073);
and U13919 (N_13919,N_13347,N_13331);
nor U13920 (N_13920,N_13745,N_12778);
nand U13921 (N_13921,N_12676,N_13621);
xor U13922 (N_13922,N_12591,N_12632);
and U13923 (N_13923,N_12606,N_12595);
xnor U13924 (N_13924,N_13230,N_13709);
nand U13925 (N_13925,N_13718,N_13547);
xor U13926 (N_13926,N_12553,N_13548);
and U13927 (N_13927,N_12602,N_12584);
xor U13928 (N_13928,N_12500,N_13395);
or U13929 (N_13929,N_13586,N_12645);
nand U13930 (N_13930,N_13319,N_13093);
xor U13931 (N_13931,N_13062,N_13396);
nand U13932 (N_13932,N_12975,N_13562);
or U13933 (N_13933,N_12701,N_13208);
xnor U13934 (N_13934,N_13328,N_12737);
or U13935 (N_13935,N_13463,N_13391);
xnor U13936 (N_13936,N_13368,N_13374);
nor U13937 (N_13937,N_13713,N_13106);
and U13938 (N_13938,N_13372,N_13699);
and U13939 (N_13939,N_13383,N_13716);
and U13940 (N_13940,N_13622,N_13011);
nor U13941 (N_13941,N_13340,N_13246);
nand U13942 (N_13942,N_12927,N_12550);
nand U13943 (N_13943,N_13524,N_12852);
nor U13944 (N_13944,N_13215,N_13672);
nand U13945 (N_13945,N_12992,N_12640);
and U13946 (N_13946,N_12501,N_12775);
nand U13947 (N_13947,N_13629,N_13432);
and U13948 (N_13948,N_12760,N_12791);
and U13949 (N_13949,N_13032,N_13351);
or U13950 (N_13950,N_13356,N_12643);
xnor U13951 (N_13951,N_13618,N_13380);
nor U13952 (N_13952,N_13590,N_12848);
and U13953 (N_13953,N_13569,N_13244);
nand U13954 (N_13954,N_13677,N_12519);
xor U13955 (N_13955,N_13128,N_13500);
nor U13956 (N_13956,N_12880,N_13212);
or U13957 (N_13957,N_13226,N_12674);
xnor U13958 (N_13958,N_12663,N_13079);
xor U13959 (N_13959,N_13058,N_12748);
and U13960 (N_13960,N_13742,N_12739);
or U13961 (N_13961,N_13275,N_12932);
or U13962 (N_13962,N_13412,N_13044);
or U13963 (N_13963,N_12647,N_12941);
nor U13964 (N_13964,N_13364,N_12820);
and U13965 (N_13965,N_13260,N_12913);
xnor U13966 (N_13966,N_13360,N_13180);
nor U13967 (N_13967,N_13527,N_13687);
xnor U13968 (N_13968,N_13623,N_13541);
or U13969 (N_13969,N_13204,N_13458);
or U13970 (N_13970,N_13353,N_13431);
nand U13971 (N_13971,N_13190,N_13451);
and U13972 (N_13972,N_12546,N_13690);
and U13973 (N_13973,N_13564,N_12987);
nor U13974 (N_13974,N_13015,N_12564);
nor U13975 (N_13975,N_13066,N_13211);
nor U13976 (N_13976,N_12846,N_12538);
nand U13977 (N_13977,N_13626,N_13486);
and U13978 (N_13978,N_12706,N_13684);
nor U13979 (N_13979,N_13257,N_13555);
or U13980 (N_13980,N_12736,N_12743);
nor U13981 (N_13981,N_12548,N_13028);
nor U13982 (N_13982,N_13556,N_13302);
or U13983 (N_13983,N_12988,N_13042);
and U13984 (N_13984,N_13025,N_13575);
xor U13985 (N_13985,N_13290,N_13119);
and U13986 (N_13986,N_13188,N_12873);
xor U13987 (N_13987,N_12933,N_13638);
and U13988 (N_13988,N_13101,N_12506);
nand U13989 (N_13989,N_13035,N_12901);
xor U13990 (N_13990,N_13449,N_13139);
nand U13991 (N_13991,N_12829,N_13343);
nand U13992 (N_13992,N_12867,N_12915);
or U13993 (N_13993,N_13000,N_12711);
or U13994 (N_13994,N_13135,N_13660);
nor U13995 (N_13995,N_12605,N_13297);
nor U13996 (N_13996,N_12804,N_12926);
and U13997 (N_13997,N_12615,N_12588);
xor U13998 (N_13998,N_13401,N_13689);
xnor U13999 (N_13999,N_13516,N_12970);
or U14000 (N_14000,N_13060,N_12965);
xor U14001 (N_14001,N_12762,N_12526);
nand U14002 (N_14002,N_12890,N_12774);
xnor U14003 (N_14003,N_13645,N_13133);
and U14004 (N_14004,N_12658,N_13278);
xor U14005 (N_14005,N_13499,N_13255);
xor U14006 (N_14006,N_13612,N_12825);
or U14007 (N_14007,N_13113,N_12742);
nand U14008 (N_14008,N_12630,N_13276);
nand U14009 (N_14009,N_12814,N_12678);
xnor U14010 (N_14010,N_12534,N_12611);
xnor U14011 (N_14011,N_13717,N_12655);
nand U14012 (N_14012,N_12772,N_13422);
or U14013 (N_14013,N_13668,N_12790);
nand U14014 (N_14014,N_12767,N_12902);
or U14015 (N_14015,N_12536,N_13040);
and U14016 (N_14016,N_13105,N_13703);
xor U14017 (N_14017,N_12968,N_13110);
and U14018 (N_14018,N_12802,N_13316);
nor U14019 (N_14019,N_13663,N_13615);
nand U14020 (N_14020,N_13251,N_13287);
and U14021 (N_14021,N_13434,N_13705);
xor U14022 (N_14022,N_13683,N_12612);
or U14023 (N_14023,N_13732,N_13631);
xnor U14024 (N_14024,N_13306,N_12953);
nand U14025 (N_14025,N_13632,N_13127);
xnor U14026 (N_14026,N_12923,N_13428);
and U14027 (N_14027,N_12872,N_12694);
nand U14028 (N_14028,N_13582,N_13181);
nor U14029 (N_14029,N_12634,N_13439);
or U14030 (N_14030,N_13460,N_12562);
xnor U14031 (N_14031,N_12555,N_12524);
and U14032 (N_14032,N_13329,N_12533);
nand U14033 (N_14033,N_13095,N_12891);
or U14034 (N_14034,N_12967,N_12529);
nor U14035 (N_14035,N_12592,N_12638);
nand U14036 (N_14036,N_13446,N_12544);
xnor U14037 (N_14037,N_13424,N_13307);
and U14038 (N_14038,N_13390,N_13574);
nand U14039 (N_14039,N_13484,N_13591);
nor U14040 (N_14040,N_12826,N_13673);
and U14041 (N_14041,N_12685,N_13377);
and U14042 (N_14042,N_13474,N_13293);
nor U14043 (N_14043,N_12765,N_13514);
nor U14044 (N_14044,N_13168,N_12997);
or U14045 (N_14045,N_13656,N_13240);
or U14046 (N_14046,N_13272,N_13137);
nand U14047 (N_14047,N_13141,N_12854);
nor U14048 (N_14048,N_12836,N_13049);
or U14049 (N_14049,N_13335,N_12641);
nand U14050 (N_14050,N_13577,N_12998);
and U14051 (N_14051,N_12691,N_12980);
xor U14052 (N_14052,N_13744,N_13406);
xnor U14053 (N_14053,N_13567,N_13604);
nor U14054 (N_14054,N_13741,N_12801);
nand U14055 (N_14055,N_13084,N_13589);
and U14056 (N_14056,N_12594,N_13680);
and U14057 (N_14057,N_12983,N_12863);
xnor U14058 (N_14058,N_13669,N_13234);
nand U14059 (N_14059,N_12696,N_12865);
xnor U14060 (N_14060,N_13089,N_12803);
nor U14061 (N_14061,N_12523,N_12857);
xor U14062 (N_14062,N_13273,N_12527);
nor U14063 (N_14063,N_12935,N_13399);
nand U14064 (N_14064,N_13560,N_12642);
xor U14065 (N_14065,N_13056,N_12569);
and U14066 (N_14066,N_12905,N_12837);
xnor U14067 (N_14067,N_13482,N_13402);
and U14068 (N_14068,N_12853,N_13509);
or U14069 (N_14069,N_13487,N_13312);
or U14070 (N_14070,N_12751,N_13706);
nand U14071 (N_14071,N_12728,N_13337);
or U14072 (N_14072,N_12719,N_12531);
nor U14073 (N_14073,N_12931,N_13261);
nor U14074 (N_14074,N_12977,N_13536);
nand U14075 (N_14075,N_12697,N_13162);
nand U14076 (N_14076,N_13707,N_12974);
nor U14077 (N_14077,N_12543,N_13445);
xor U14078 (N_14078,N_12821,N_13551);
nor U14079 (N_14079,N_13134,N_13069);
or U14080 (N_14080,N_12614,N_12741);
xnor U14081 (N_14081,N_13459,N_12709);
and U14082 (N_14082,N_13102,N_12945);
or U14083 (N_14083,N_13130,N_13038);
and U14084 (N_14084,N_13213,N_12732);
or U14085 (N_14085,N_13640,N_12824);
or U14086 (N_14086,N_13144,N_13644);
nor U14087 (N_14087,N_12773,N_13252);
xnor U14088 (N_14088,N_13600,N_13657);
xor U14089 (N_14089,N_13132,N_12575);
or U14090 (N_14090,N_13282,N_12944);
or U14091 (N_14091,N_12995,N_12813);
nand U14092 (N_14092,N_13238,N_12560);
and U14093 (N_14093,N_13476,N_12714);
or U14094 (N_14094,N_12585,N_13643);
or U14095 (N_14095,N_13517,N_13641);
nand U14096 (N_14096,N_13176,N_12657);
nand U14097 (N_14097,N_12850,N_13525);
and U14098 (N_14098,N_13308,N_13734);
or U14099 (N_14099,N_13492,N_12895);
nor U14100 (N_14100,N_13284,N_12583);
nand U14101 (N_14101,N_12572,N_12960);
or U14102 (N_14102,N_13521,N_13584);
and U14103 (N_14103,N_12661,N_13080);
xnor U14104 (N_14104,N_12860,N_12619);
and U14105 (N_14105,N_12921,N_12795);
or U14106 (N_14106,N_13047,N_13462);
or U14107 (N_14107,N_13542,N_12717);
xor U14108 (N_14108,N_12604,N_12715);
and U14109 (N_14109,N_13496,N_13515);
or U14110 (N_14110,N_13361,N_13473);
or U14111 (N_14111,N_12832,N_13254);
or U14112 (N_14112,N_13438,N_12551);
nand U14113 (N_14113,N_13075,N_12542);
nor U14114 (N_14114,N_12899,N_13721);
and U14115 (N_14115,N_12925,N_13096);
nor U14116 (N_14116,N_13003,N_12609);
nand U14117 (N_14117,N_12651,N_13570);
and U14118 (N_14118,N_12991,N_12722);
nor U14119 (N_14119,N_12904,N_13021);
nor U14120 (N_14120,N_12990,N_13033);
and U14121 (N_14121,N_12692,N_13493);
nor U14122 (N_14122,N_13506,N_12818);
or U14123 (N_14123,N_13579,N_12713);
or U14124 (N_14124,N_12938,N_12884);
xor U14125 (N_14125,N_12781,N_12859);
nand U14126 (N_14126,N_12707,N_13022);
or U14127 (N_14127,N_13453,N_12631);
or U14128 (N_14128,N_13553,N_12937);
xor U14129 (N_14129,N_13196,N_12673);
and U14130 (N_14130,N_13585,N_12916);
xnor U14131 (N_14131,N_13344,N_12897);
nor U14132 (N_14132,N_12744,N_13441);
xnor U14133 (N_14133,N_12875,N_12508);
and U14134 (N_14134,N_12840,N_12626);
xnor U14135 (N_14135,N_13248,N_12957);
nor U14136 (N_14136,N_13397,N_13065);
and U14137 (N_14137,N_13712,N_13323);
nand U14138 (N_14138,N_13286,N_13480);
or U14139 (N_14139,N_12580,N_12841);
and U14140 (N_14140,N_13722,N_13528);
nor U14141 (N_14141,N_13420,N_13723);
and U14142 (N_14142,N_12831,N_12834);
nor U14143 (N_14143,N_13691,N_12908);
and U14144 (N_14144,N_13538,N_13138);
xnor U14145 (N_14145,N_12888,N_12969);
nand U14146 (N_14146,N_13318,N_13149);
or U14147 (N_14147,N_12817,N_12822);
nor U14148 (N_14148,N_12948,N_12660);
nand U14149 (N_14149,N_13001,N_12502);
or U14150 (N_14150,N_13173,N_12704);
nand U14151 (N_14151,N_12806,N_12700);
nand U14152 (N_14152,N_13103,N_12903);
nor U14153 (N_14153,N_12783,N_13511);
and U14154 (N_14154,N_12788,N_12509);
nand U14155 (N_14155,N_12578,N_13006);
xnor U14156 (N_14156,N_13650,N_12733);
nand U14157 (N_14157,N_12537,N_12518);
nor U14158 (N_14158,N_13363,N_12633);
nor U14159 (N_14159,N_12567,N_12637);
nor U14160 (N_14160,N_13126,N_12950);
xnor U14161 (N_14161,N_12656,N_12919);
nor U14162 (N_14162,N_13736,N_12800);
nand U14163 (N_14163,N_13250,N_13665);
or U14164 (N_14164,N_13727,N_13740);
or U14165 (N_14165,N_13197,N_13670);
nor U14166 (N_14166,N_13367,N_13609);
xnor U14167 (N_14167,N_12652,N_12670);
nand U14168 (N_14168,N_13294,N_12989);
and U14169 (N_14169,N_13224,N_12973);
xor U14170 (N_14170,N_13735,N_13565);
xor U14171 (N_14171,N_13447,N_12671);
nor U14172 (N_14172,N_12650,N_13520);
nor U14173 (N_14173,N_12582,N_13737);
xnor U14174 (N_14174,N_12952,N_12750);
or U14175 (N_14175,N_13620,N_13358);
or U14176 (N_14176,N_13599,N_12942);
xnor U14177 (N_14177,N_12559,N_12827);
xnor U14178 (N_14178,N_13048,N_13411);
xor U14179 (N_14179,N_12593,N_13303);
and U14180 (N_14180,N_13566,N_13059);
and U14181 (N_14181,N_12624,N_12755);
nor U14182 (N_14182,N_12558,N_13468);
nor U14183 (N_14183,N_13209,N_12799);
or U14184 (N_14184,N_13505,N_12577);
nand U14185 (N_14185,N_13630,N_13613);
or U14186 (N_14186,N_13076,N_13485);
or U14187 (N_14187,N_13262,N_12871);
nand U14188 (N_14188,N_12684,N_13393);
and U14189 (N_14189,N_13313,N_12574);
or U14190 (N_14190,N_13233,N_13354);
or U14191 (N_14191,N_13315,N_13642);
or U14192 (N_14192,N_12726,N_12936);
xnor U14193 (N_14193,N_12766,N_13107);
nand U14194 (N_14194,N_13283,N_12708);
nor U14195 (N_14195,N_12856,N_13561);
nand U14196 (N_14196,N_13702,N_13697);
or U14197 (N_14197,N_13055,N_12893);
and U14198 (N_14198,N_13530,N_13544);
nor U14199 (N_14199,N_13601,N_13004);
xnor U14200 (N_14200,N_12807,N_13277);
and U14201 (N_14201,N_13503,N_13120);
or U14202 (N_14202,N_12810,N_12889);
nor U14203 (N_14203,N_13070,N_13288);
or U14204 (N_14204,N_13289,N_12855);
xor U14205 (N_14205,N_13083,N_12951);
or U14206 (N_14206,N_13150,N_13537);
nor U14207 (N_14207,N_13679,N_13164);
nand U14208 (N_14208,N_13369,N_13675);
nor U14209 (N_14209,N_13554,N_13549);
or U14210 (N_14210,N_13436,N_13583);
xnor U14211 (N_14211,N_13342,N_12680);
xor U14212 (N_14212,N_12712,N_13437);
xor U14213 (N_14213,N_13698,N_13140);
nor U14214 (N_14214,N_12654,N_13232);
and U14215 (N_14215,N_13227,N_13266);
and U14216 (N_14216,N_12909,N_12882);
nand U14217 (N_14217,N_12532,N_12516);
xnor U14218 (N_14218,N_12589,N_13546);
nor U14219 (N_14219,N_12693,N_13063);
or U14220 (N_14220,N_13228,N_12784);
xor U14221 (N_14221,N_13594,N_13639);
or U14222 (N_14222,N_12520,N_12878);
nand U14223 (N_14223,N_13518,N_12622);
nor U14224 (N_14224,N_13479,N_13265);
or U14225 (N_14225,N_13111,N_12984);
xnor U14226 (N_14226,N_12838,N_12796);
nand U14227 (N_14227,N_12851,N_12659);
xnor U14228 (N_14228,N_13067,N_13624);
xor U14229 (N_14229,N_12999,N_12503);
xnor U14230 (N_14230,N_13381,N_13533);
or U14231 (N_14231,N_13086,N_13534);
xnor U14232 (N_14232,N_13513,N_13674);
and U14233 (N_14233,N_13676,N_12964);
nand U14234 (N_14234,N_12522,N_13747);
nand U14235 (N_14235,N_12702,N_12729);
xnor U14236 (N_14236,N_12746,N_12758);
and U14237 (N_14237,N_13271,N_13165);
nand U14238 (N_14238,N_13285,N_12769);
or U14239 (N_14239,N_13467,N_13013);
xnor U14240 (N_14240,N_12621,N_13142);
nor U14241 (N_14241,N_12883,N_12930);
or U14242 (N_14242,N_13320,N_13404);
xnor U14243 (N_14243,N_12994,N_12565);
and U14244 (N_14244,N_13733,N_13189);
xor U14245 (N_14245,N_13384,N_12576);
xor U14246 (N_14246,N_12782,N_13045);
nand U14247 (N_14247,N_13634,N_13603);
nor U14248 (N_14248,N_13210,N_12735);
or U14249 (N_14249,N_13386,N_13160);
or U14250 (N_14250,N_13159,N_13264);
and U14251 (N_14251,N_13305,N_13321);
nand U14252 (N_14252,N_13719,N_13229);
nor U14253 (N_14253,N_13611,N_13578);
and U14254 (N_14254,N_13710,N_12699);
nor U14255 (N_14255,N_13292,N_12607);
nand U14256 (N_14256,N_13072,N_12780);
xnor U14257 (N_14257,N_12616,N_13192);
and U14258 (N_14258,N_13023,N_12885);
and U14259 (N_14259,N_13217,N_13046);
nand U14260 (N_14260,N_13185,N_13349);
and U14261 (N_14261,N_12690,N_13617);
or U14262 (N_14262,N_13206,N_13616);
nor U14263 (N_14263,N_13249,N_13090);
xor U14264 (N_14264,N_12608,N_13426);
nand U14265 (N_14265,N_12698,N_12981);
nand U14266 (N_14266,N_13427,N_13392);
nor U14267 (N_14267,N_12789,N_12629);
and U14268 (N_14268,N_12868,N_13433);
xnor U14269 (N_14269,N_12959,N_12507);
xor U14270 (N_14270,N_13193,N_12947);
nand U14271 (N_14271,N_13654,N_13117);
nand U14272 (N_14272,N_13098,N_13497);
xnor U14273 (N_14273,N_13400,N_13108);
nand U14274 (N_14274,N_13231,N_13597);
nor U14275 (N_14275,N_13748,N_12512);
xor U14276 (N_14276,N_12958,N_13408);
or U14277 (N_14277,N_13481,N_12978);
or U14278 (N_14278,N_13157,N_13026);
nand U14279 (N_14279,N_12695,N_13223);
and U14280 (N_14280,N_13471,N_13029);
nor U14281 (N_14281,N_13241,N_12962);
and U14282 (N_14282,N_13407,N_12568);
nand U14283 (N_14283,N_12756,N_13123);
or U14284 (N_14284,N_13388,N_12966);
nor U14285 (N_14285,N_13488,N_13054);
nand U14286 (N_14286,N_12688,N_13322);
xor U14287 (N_14287,N_13325,N_13455);
and U14288 (N_14288,N_13726,N_13243);
xnor U14289 (N_14289,N_12635,N_12812);
or U14290 (N_14290,N_13018,N_12745);
nand U14291 (N_14291,N_13314,N_13267);
or U14292 (N_14292,N_13324,N_13593);
and U14293 (N_14293,N_13129,N_13405);
or U14294 (N_14294,N_12862,N_13078);
nand U14295 (N_14295,N_13202,N_13258);
xnor U14296 (N_14296,N_13327,N_12911);
and U14297 (N_14297,N_12740,N_12956);
nor U14298 (N_14298,N_13237,N_13731);
nor U14299 (N_14299,N_13012,N_13235);
xor U14300 (N_14300,N_13245,N_12598);
or U14301 (N_14301,N_12720,N_13218);
and U14302 (N_14302,N_13136,N_12809);
nor U14303 (N_14303,N_13161,N_12785);
xor U14304 (N_14304,N_12892,N_13743);
and U14305 (N_14305,N_13163,N_13034);
or U14306 (N_14306,N_12906,N_13671);
nor U14307 (N_14307,N_12828,N_13409);
or U14308 (N_14308,N_13050,N_13017);
and U14309 (N_14309,N_13711,N_13097);
or U14310 (N_14310,N_12505,N_13317);
nor U14311 (N_14311,N_13121,N_13523);
nand U14312 (N_14312,N_13199,N_12928);
or U14313 (N_14313,N_12985,N_13216);
nand U14314 (N_14314,N_13559,N_13094);
nand U14315 (N_14315,N_13550,N_12682);
nand U14316 (N_14316,N_12786,N_13461);
or U14317 (N_14317,N_12617,N_13253);
nand U14318 (N_14318,N_12721,N_12623);
nor U14319 (N_14319,N_13470,N_12541);
xnor U14320 (N_14320,N_13186,N_13552);
or U14321 (N_14321,N_13016,N_13708);
nor U14322 (N_14322,N_13417,N_12839);
or U14323 (N_14323,N_13039,N_13512);
xor U14324 (N_14324,N_12601,N_13646);
xnor U14325 (N_14325,N_12798,N_13221);
nand U14326 (N_14326,N_13019,N_12963);
nand U14327 (N_14327,N_13635,N_13187);
nand U14328 (N_14328,N_13350,N_13728);
nor U14329 (N_14329,N_13061,N_13563);
nor U14330 (N_14330,N_13177,N_13124);
and U14331 (N_14331,N_12666,N_12858);
nor U14332 (N_14332,N_12768,N_13649);
nor U14333 (N_14333,N_13382,N_12724);
or U14334 (N_14334,N_12979,N_13195);
nand U14335 (N_14335,N_12677,N_13389);
nor U14336 (N_14336,N_13295,N_12552);
or U14337 (N_14337,N_13558,N_12940);
xor U14338 (N_14338,N_13172,N_13504);
nor U14339 (N_14339,N_13300,N_12794);
nor U14340 (N_14340,N_12579,N_12727);
and U14341 (N_14341,N_12639,N_13371);
xor U14342 (N_14342,N_12845,N_12620);
nand U14343 (N_14343,N_13695,N_12504);
and U14344 (N_14344,N_12910,N_12667);
or U14345 (N_14345,N_13256,N_13581);
or U14346 (N_14346,N_13156,N_12581);
or U14347 (N_14347,N_13027,N_13637);
or U14348 (N_14348,N_12716,N_13239);
or U14349 (N_14349,N_12600,N_12528);
or U14350 (N_14350,N_13443,N_12752);
xnor U14351 (N_14351,N_12513,N_13279);
xor U14352 (N_14352,N_13456,N_13122);
xor U14353 (N_14353,N_13304,N_13299);
or U14354 (N_14354,N_13415,N_12792);
nor U14355 (N_14355,N_13685,N_12819);
xnor U14356 (N_14356,N_13326,N_13701);
and U14357 (N_14357,N_13508,N_12662);
or U14358 (N_14358,N_12787,N_13182);
and U14359 (N_14359,N_13357,N_12996);
xnor U14360 (N_14360,N_12525,N_13041);
nor U14361 (N_14361,N_12540,N_12844);
or U14362 (N_14362,N_13291,N_12664);
nand U14363 (N_14363,N_12547,N_13440);
and U14364 (N_14364,N_13366,N_13681);
xnor U14365 (N_14365,N_12876,N_13738);
nor U14366 (N_14366,N_13598,N_12986);
xor U14367 (N_14367,N_13557,N_12511);
and U14368 (N_14368,N_13587,N_13647);
and U14369 (N_14369,N_12510,N_12753);
or U14370 (N_14370,N_13088,N_12599);
xor U14371 (N_14371,N_13145,N_12955);
xor U14372 (N_14372,N_12886,N_13419);
nand U14373 (N_14373,N_13167,N_12835);
xor U14374 (N_14374,N_12971,N_13201);
or U14375 (N_14375,N_13530,N_13488);
nand U14376 (N_14376,N_12657,N_13185);
and U14377 (N_14377,N_13692,N_13420);
or U14378 (N_14378,N_12785,N_12577);
nor U14379 (N_14379,N_12681,N_13139);
nand U14380 (N_14380,N_13688,N_13561);
and U14381 (N_14381,N_12881,N_13736);
xnor U14382 (N_14382,N_12788,N_12855);
and U14383 (N_14383,N_13529,N_12627);
or U14384 (N_14384,N_13281,N_12514);
xnor U14385 (N_14385,N_13131,N_13213);
nor U14386 (N_14386,N_12919,N_13356);
or U14387 (N_14387,N_12884,N_12751);
nand U14388 (N_14388,N_13056,N_13616);
or U14389 (N_14389,N_12652,N_13649);
or U14390 (N_14390,N_13357,N_13066);
nor U14391 (N_14391,N_13301,N_12720);
xor U14392 (N_14392,N_12720,N_13504);
xor U14393 (N_14393,N_13505,N_13682);
nand U14394 (N_14394,N_13180,N_13495);
nand U14395 (N_14395,N_12623,N_13183);
or U14396 (N_14396,N_12631,N_13666);
xnor U14397 (N_14397,N_12897,N_13498);
xnor U14398 (N_14398,N_13467,N_13551);
or U14399 (N_14399,N_13729,N_12564);
nand U14400 (N_14400,N_13304,N_13645);
xor U14401 (N_14401,N_13544,N_12706);
nor U14402 (N_14402,N_12986,N_13389);
nand U14403 (N_14403,N_12719,N_12862);
or U14404 (N_14404,N_12635,N_13412);
or U14405 (N_14405,N_13288,N_13223);
xnor U14406 (N_14406,N_13304,N_13558);
or U14407 (N_14407,N_12805,N_12988);
and U14408 (N_14408,N_13562,N_12655);
nand U14409 (N_14409,N_12596,N_13711);
nand U14410 (N_14410,N_13527,N_12607);
xor U14411 (N_14411,N_12691,N_12626);
and U14412 (N_14412,N_13262,N_13532);
and U14413 (N_14413,N_12555,N_12666);
or U14414 (N_14414,N_13745,N_13556);
nand U14415 (N_14415,N_13385,N_12590);
xnor U14416 (N_14416,N_12510,N_13503);
or U14417 (N_14417,N_13707,N_13727);
xnor U14418 (N_14418,N_13730,N_12786);
nor U14419 (N_14419,N_12720,N_13175);
xnor U14420 (N_14420,N_13025,N_13674);
nand U14421 (N_14421,N_12748,N_13489);
nor U14422 (N_14422,N_13543,N_12845);
and U14423 (N_14423,N_13651,N_13491);
xnor U14424 (N_14424,N_12973,N_13608);
or U14425 (N_14425,N_13669,N_12539);
nor U14426 (N_14426,N_12847,N_12820);
or U14427 (N_14427,N_13744,N_13557);
nand U14428 (N_14428,N_12875,N_13065);
and U14429 (N_14429,N_12516,N_13195);
nor U14430 (N_14430,N_13539,N_13285);
or U14431 (N_14431,N_13111,N_12577);
xor U14432 (N_14432,N_13010,N_12847);
and U14433 (N_14433,N_13221,N_13355);
nand U14434 (N_14434,N_13046,N_12863);
or U14435 (N_14435,N_13423,N_13371);
nor U14436 (N_14436,N_12969,N_13394);
nor U14437 (N_14437,N_13523,N_12632);
or U14438 (N_14438,N_12527,N_13390);
nor U14439 (N_14439,N_13730,N_13460);
nor U14440 (N_14440,N_13289,N_13541);
or U14441 (N_14441,N_13656,N_13191);
nand U14442 (N_14442,N_13007,N_12571);
xor U14443 (N_14443,N_13443,N_12535);
nand U14444 (N_14444,N_13422,N_12859);
nor U14445 (N_14445,N_12765,N_13174);
xor U14446 (N_14446,N_13248,N_12670);
and U14447 (N_14447,N_13500,N_13676);
nor U14448 (N_14448,N_13583,N_12895);
xor U14449 (N_14449,N_12884,N_12556);
nand U14450 (N_14450,N_13125,N_13255);
nor U14451 (N_14451,N_12944,N_12845);
nand U14452 (N_14452,N_12813,N_12966);
nor U14453 (N_14453,N_12890,N_13140);
or U14454 (N_14454,N_13334,N_13116);
or U14455 (N_14455,N_13517,N_13563);
nand U14456 (N_14456,N_12933,N_12983);
nand U14457 (N_14457,N_12945,N_12715);
nor U14458 (N_14458,N_13718,N_13379);
or U14459 (N_14459,N_12530,N_13494);
and U14460 (N_14460,N_12846,N_13040);
nor U14461 (N_14461,N_12513,N_13539);
or U14462 (N_14462,N_13224,N_13610);
nand U14463 (N_14463,N_12668,N_13158);
xor U14464 (N_14464,N_12605,N_13034);
or U14465 (N_14465,N_13310,N_12754);
and U14466 (N_14466,N_13680,N_13702);
and U14467 (N_14467,N_13477,N_12732);
xor U14468 (N_14468,N_13280,N_12737);
nand U14469 (N_14469,N_13402,N_13632);
and U14470 (N_14470,N_12882,N_12629);
nand U14471 (N_14471,N_13062,N_13313);
xnor U14472 (N_14472,N_12620,N_13725);
nand U14473 (N_14473,N_13641,N_13124);
xnor U14474 (N_14474,N_13381,N_13078);
nor U14475 (N_14475,N_13196,N_13613);
nor U14476 (N_14476,N_13330,N_13540);
or U14477 (N_14477,N_12699,N_13034);
nand U14478 (N_14478,N_13266,N_12940);
and U14479 (N_14479,N_13269,N_12579);
and U14480 (N_14480,N_12646,N_13736);
xnor U14481 (N_14481,N_12543,N_13555);
or U14482 (N_14482,N_13301,N_13739);
nand U14483 (N_14483,N_12535,N_12770);
and U14484 (N_14484,N_13007,N_13239);
and U14485 (N_14485,N_13426,N_13063);
or U14486 (N_14486,N_12744,N_13135);
or U14487 (N_14487,N_12697,N_13555);
nand U14488 (N_14488,N_12955,N_13747);
nor U14489 (N_14489,N_13171,N_13238);
nand U14490 (N_14490,N_12918,N_12999);
or U14491 (N_14491,N_12668,N_12926);
or U14492 (N_14492,N_12930,N_13480);
and U14493 (N_14493,N_13014,N_12767);
or U14494 (N_14494,N_13008,N_13225);
and U14495 (N_14495,N_13414,N_13437);
and U14496 (N_14496,N_12682,N_12640);
nor U14497 (N_14497,N_13355,N_12946);
or U14498 (N_14498,N_13034,N_13304);
or U14499 (N_14499,N_13352,N_12674);
or U14500 (N_14500,N_13187,N_13127);
nor U14501 (N_14501,N_12596,N_12815);
nand U14502 (N_14502,N_12867,N_12811);
and U14503 (N_14503,N_13021,N_13351);
nand U14504 (N_14504,N_13432,N_12544);
nor U14505 (N_14505,N_12731,N_13530);
or U14506 (N_14506,N_12988,N_12757);
or U14507 (N_14507,N_13169,N_13015);
nor U14508 (N_14508,N_13724,N_12859);
xnor U14509 (N_14509,N_12516,N_13075);
xor U14510 (N_14510,N_12888,N_12885);
xor U14511 (N_14511,N_12593,N_13424);
nand U14512 (N_14512,N_13689,N_12906);
or U14513 (N_14513,N_13365,N_13191);
or U14514 (N_14514,N_12599,N_12713);
or U14515 (N_14515,N_13422,N_13372);
or U14516 (N_14516,N_13163,N_13495);
nor U14517 (N_14517,N_13628,N_13498);
xor U14518 (N_14518,N_13200,N_13351);
and U14519 (N_14519,N_12501,N_13290);
nor U14520 (N_14520,N_12825,N_13625);
nor U14521 (N_14521,N_12930,N_13516);
and U14522 (N_14522,N_13714,N_12940);
nand U14523 (N_14523,N_13307,N_13200);
nand U14524 (N_14524,N_13364,N_13272);
nand U14525 (N_14525,N_13357,N_12981);
xnor U14526 (N_14526,N_12581,N_12761);
nor U14527 (N_14527,N_12766,N_13525);
nor U14528 (N_14528,N_13388,N_13662);
xor U14529 (N_14529,N_13214,N_12890);
nor U14530 (N_14530,N_12970,N_13706);
nor U14531 (N_14531,N_13140,N_12924);
or U14532 (N_14532,N_13471,N_13552);
and U14533 (N_14533,N_13348,N_13609);
or U14534 (N_14534,N_12871,N_12668);
nand U14535 (N_14535,N_12601,N_13290);
and U14536 (N_14536,N_12795,N_12869);
xnor U14537 (N_14537,N_12949,N_13716);
nor U14538 (N_14538,N_13178,N_12795);
or U14539 (N_14539,N_13714,N_12772);
xnor U14540 (N_14540,N_13687,N_12519);
xor U14541 (N_14541,N_13685,N_13018);
nor U14542 (N_14542,N_13684,N_13636);
xnor U14543 (N_14543,N_13352,N_13661);
or U14544 (N_14544,N_12666,N_12749);
and U14545 (N_14545,N_12827,N_12752);
or U14546 (N_14546,N_13559,N_12962);
or U14547 (N_14547,N_12687,N_12697);
nand U14548 (N_14548,N_12713,N_12936);
nand U14549 (N_14549,N_12876,N_12547);
nand U14550 (N_14550,N_12515,N_12808);
nand U14551 (N_14551,N_13250,N_12685);
nor U14552 (N_14552,N_13469,N_13661);
xor U14553 (N_14553,N_12903,N_12577);
nor U14554 (N_14554,N_13684,N_12630);
nand U14555 (N_14555,N_13179,N_13241);
or U14556 (N_14556,N_12691,N_13240);
nand U14557 (N_14557,N_13445,N_13439);
or U14558 (N_14558,N_12803,N_13327);
nor U14559 (N_14559,N_12799,N_13270);
nand U14560 (N_14560,N_12742,N_12533);
and U14561 (N_14561,N_12544,N_13248);
or U14562 (N_14562,N_13019,N_13192);
nand U14563 (N_14563,N_13015,N_13143);
nor U14564 (N_14564,N_13435,N_12924);
xor U14565 (N_14565,N_12549,N_12963);
nor U14566 (N_14566,N_13319,N_12954);
or U14567 (N_14567,N_12503,N_13085);
and U14568 (N_14568,N_13113,N_12506);
and U14569 (N_14569,N_12973,N_13132);
or U14570 (N_14570,N_13500,N_13388);
or U14571 (N_14571,N_13322,N_13095);
nand U14572 (N_14572,N_12540,N_13240);
nand U14573 (N_14573,N_12959,N_13135);
and U14574 (N_14574,N_12700,N_12976);
nand U14575 (N_14575,N_12939,N_13227);
and U14576 (N_14576,N_12725,N_12562);
nor U14577 (N_14577,N_13705,N_13035);
nand U14578 (N_14578,N_13025,N_12503);
and U14579 (N_14579,N_13276,N_13280);
xor U14580 (N_14580,N_13199,N_13095);
nor U14581 (N_14581,N_13566,N_12895);
or U14582 (N_14582,N_13201,N_13746);
xnor U14583 (N_14583,N_13644,N_12986);
or U14584 (N_14584,N_13503,N_13026);
nor U14585 (N_14585,N_12731,N_13664);
and U14586 (N_14586,N_12874,N_12786);
xnor U14587 (N_14587,N_12587,N_12699);
nand U14588 (N_14588,N_12930,N_12579);
and U14589 (N_14589,N_12689,N_12604);
or U14590 (N_14590,N_12502,N_12618);
xnor U14591 (N_14591,N_13282,N_12948);
or U14592 (N_14592,N_12951,N_12709);
xnor U14593 (N_14593,N_13404,N_12769);
xnor U14594 (N_14594,N_12516,N_12805);
xor U14595 (N_14595,N_13036,N_13700);
nor U14596 (N_14596,N_12645,N_13446);
xor U14597 (N_14597,N_13271,N_12954);
or U14598 (N_14598,N_13729,N_13282);
and U14599 (N_14599,N_12773,N_12627);
xnor U14600 (N_14600,N_12899,N_13715);
nand U14601 (N_14601,N_13334,N_13226);
or U14602 (N_14602,N_13702,N_12995);
or U14603 (N_14603,N_13322,N_13287);
nand U14604 (N_14604,N_13708,N_12562);
nand U14605 (N_14605,N_13160,N_13136);
xnor U14606 (N_14606,N_12551,N_12876);
nand U14607 (N_14607,N_13350,N_13467);
xnor U14608 (N_14608,N_12680,N_12878);
and U14609 (N_14609,N_13520,N_13280);
or U14610 (N_14610,N_13087,N_12553);
xor U14611 (N_14611,N_13001,N_13051);
and U14612 (N_14612,N_12628,N_13290);
nand U14613 (N_14613,N_13607,N_13444);
or U14614 (N_14614,N_13371,N_12501);
and U14615 (N_14615,N_12987,N_13059);
xnor U14616 (N_14616,N_12735,N_13507);
nor U14617 (N_14617,N_12767,N_12802);
nor U14618 (N_14618,N_13670,N_12502);
xnor U14619 (N_14619,N_12547,N_13628);
or U14620 (N_14620,N_13736,N_13379);
xor U14621 (N_14621,N_13263,N_13383);
xor U14622 (N_14622,N_12515,N_12693);
and U14623 (N_14623,N_13423,N_12596);
xnor U14624 (N_14624,N_12933,N_12888);
or U14625 (N_14625,N_13313,N_13361);
or U14626 (N_14626,N_12646,N_12967);
and U14627 (N_14627,N_13340,N_13013);
and U14628 (N_14628,N_12838,N_12695);
nor U14629 (N_14629,N_12894,N_12632);
nor U14630 (N_14630,N_12566,N_13724);
and U14631 (N_14631,N_12759,N_13430);
and U14632 (N_14632,N_13144,N_13633);
xor U14633 (N_14633,N_13503,N_12815);
nor U14634 (N_14634,N_12645,N_13411);
nand U14635 (N_14635,N_13065,N_13420);
xnor U14636 (N_14636,N_13274,N_12931);
nor U14637 (N_14637,N_12583,N_12625);
nand U14638 (N_14638,N_13659,N_13231);
and U14639 (N_14639,N_13191,N_13210);
xor U14640 (N_14640,N_13296,N_13081);
or U14641 (N_14641,N_13269,N_13029);
or U14642 (N_14642,N_13541,N_13048);
nand U14643 (N_14643,N_13164,N_12575);
xor U14644 (N_14644,N_12591,N_13250);
or U14645 (N_14645,N_13495,N_13276);
and U14646 (N_14646,N_12823,N_12877);
nor U14647 (N_14647,N_12697,N_12962);
xor U14648 (N_14648,N_13112,N_13056);
or U14649 (N_14649,N_13509,N_13289);
xnor U14650 (N_14650,N_12980,N_13086);
nor U14651 (N_14651,N_12569,N_12916);
nand U14652 (N_14652,N_13553,N_12631);
or U14653 (N_14653,N_13409,N_13425);
nor U14654 (N_14654,N_12834,N_12991);
or U14655 (N_14655,N_12670,N_12816);
nand U14656 (N_14656,N_13254,N_13624);
and U14657 (N_14657,N_12908,N_13579);
and U14658 (N_14658,N_13161,N_13468);
nor U14659 (N_14659,N_13596,N_12695);
xor U14660 (N_14660,N_12943,N_13244);
or U14661 (N_14661,N_12982,N_13391);
nand U14662 (N_14662,N_13134,N_12921);
or U14663 (N_14663,N_13356,N_12655);
nand U14664 (N_14664,N_13220,N_13300);
and U14665 (N_14665,N_12701,N_12936);
xor U14666 (N_14666,N_13229,N_12882);
and U14667 (N_14667,N_12932,N_13474);
or U14668 (N_14668,N_12986,N_13035);
nand U14669 (N_14669,N_12514,N_13067);
and U14670 (N_14670,N_13696,N_12586);
nor U14671 (N_14671,N_13316,N_13403);
xor U14672 (N_14672,N_12588,N_12822);
xor U14673 (N_14673,N_12872,N_13312);
and U14674 (N_14674,N_13251,N_12570);
and U14675 (N_14675,N_12557,N_12918);
nor U14676 (N_14676,N_13035,N_12868);
xnor U14677 (N_14677,N_13217,N_13009);
or U14678 (N_14678,N_13716,N_13490);
nor U14679 (N_14679,N_12561,N_13181);
nor U14680 (N_14680,N_13082,N_12748);
xnor U14681 (N_14681,N_12723,N_13024);
and U14682 (N_14682,N_13584,N_13631);
or U14683 (N_14683,N_13496,N_12614);
nand U14684 (N_14684,N_13028,N_12616);
xnor U14685 (N_14685,N_13601,N_13620);
or U14686 (N_14686,N_12788,N_13241);
nand U14687 (N_14687,N_13615,N_12825);
or U14688 (N_14688,N_12605,N_13577);
and U14689 (N_14689,N_13567,N_12767);
nor U14690 (N_14690,N_13010,N_13337);
nand U14691 (N_14691,N_12546,N_13631);
nand U14692 (N_14692,N_12929,N_13468);
and U14693 (N_14693,N_13345,N_13579);
xor U14694 (N_14694,N_12794,N_13363);
xor U14695 (N_14695,N_13389,N_12768);
and U14696 (N_14696,N_12777,N_12531);
and U14697 (N_14697,N_13497,N_13425);
nor U14698 (N_14698,N_12925,N_12802);
xnor U14699 (N_14699,N_12776,N_12947);
nand U14700 (N_14700,N_13349,N_13666);
and U14701 (N_14701,N_12853,N_12720);
nand U14702 (N_14702,N_12805,N_13686);
or U14703 (N_14703,N_13263,N_13256);
or U14704 (N_14704,N_12509,N_13598);
xnor U14705 (N_14705,N_12789,N_13710);
xor U14706 (N_14706,N_13413,N_13000);
nor U14707 (N_14707,N_13613,N_13486);
xor U14708 (N_14708,N_12807,N_13568);
nor U14709 (N_14709,N_13503,N_13634);
xor U14710 (N_14710,N_12723,N_13744);
nand U14711 (N_14711,N_13188,N_13207);
or U14712 (N_14712,N_12733,N_13661);
nor U14713 (N_14713,N_13555,N_12808);
nand U14714 (N_14714,N_13121,N_12702);
or U14715 (N_14715,N_12874,N_13604);
xor U14716 (N_14716,N_13042,N_13693);
or U14717 (N_14717,N_12689,N_12863);
nand U14718 (N_14718,N_12741,N_12545);
nor U14719 (N_14719,N_13440,N_12616);
or U14720 (N_14720,N_13612,N_13192);
nor U14721 (N_14721,N_12519,N_12958);
nor U14722 (N_14722,N_12809,N_13444);
and U14723 (N_14723,N_13464,N_13453);
and U14724 (N_14724,N_13270,N_13420);
nand U14725 (N_14725,N_13395,N_13497);
nand U14726 (N_14726,N_12581,N_12936);
nand U14727 (N_14727,N_13065,N_13542);
nand U14728 (N_14728,N_13489,N_12678);
nor U14729 (N_14729,N_13457,N_12976);
xnor U14730 (N_14730,N_13260,N_12654);
nand U14731 (N_14731,N_13158,N_13631);
xor U14732 (N_14732,N_12648,N_13283);
and U14733 (N_14733,N_13305,N_12714);
and U14734 (N_14734,N_12637,N_13549);
xor U14735 (N_14735,N_12734,N_12861);
xor U14736 (N_14736,N_13623,N_13259);
nand U14737 (N_14737,N_13642,N_12863);
nand U14738 (N_14738,N_13034,N_13169);
and U14739 (N_14739,N_13667,N_13179);
nand U14740 (N_14740,N_13092,N_12933);
nor U14741 (N_14741,N_12925,N_13469);
and U14742 (N_14742,N_12873,N_13531);
and U14743 (N_14743,N_13233,N_13186);
or U14744 (N_14744,N_13114,N_13496);
xnor U14745 (N_14745,N_12575,N_13223);
nand U14746 (N_14746,N_13547,N_13639);
nor U14747 (N_14747,N_13114,N_12559);
or U14748 (N_14748,N_13405,N_13675);
and U14749 (N_14749,N_13328,N_13400);
xor U14750 (N_14750,N_13696,N_12573);
xor U14751 (N_14751,N_13456,N_13154);
xor U14752 (N_14752,N_12615,N_13380);
nand U14753 (N_14753,N_12960,N_12939);
nor U14754 (N_14754,N_13161,N_13555);
xor U14755 (N_14755,N_13624,N_13389);
nand U14756 (N_14756,N_13416,N_13531);
xnor U14757 (N_14757,N_12733,N_13743);
xor U14758 (N_14758,N_12870,N_13430);
or U14759 (N_14759,N_13355,N_13482);
and U14760 (N_14760,N_12841,N_12768);
nor U14761 (N_14761,N_13042,N_13155);
nand U14762 (N_14762,N_13019,N_13395);
and U14763 (N_14763,N_13513,N_12621);
nor U14764 (N_14764,N_13518,N_13008);
and U14765 (N_14765,N_13578,N_13077);
and U14766 (N_14766,N_13025,N_12539);
xor U14767 (N_14767,N_13683,N_13103);
or U14768 (N_14768,N_13127,N_13051);
xor U14769 (N_14769,N_13606,N_13563);
and U14770 (N_14770,N_13588,N_13286);
nand U14771 (N_14771,N_12563,N_13560);
or U14772 (N_14772,N_12852,N_12944);
nand U14773 (N_14773,N_12934,N_13569);
nor U14774 (N_14774,N_12850,N_12515);
xor U14775 (N_14775,N_13066,N_12980);
and U14776 (N_14776,N_13449,N_13171);
or U14777 (N_14777,N_12702,N_12608);
nand U14778 (N_14778,N_12632,N_13259);
xor U14779 (N_14779,N_13498,N_13615);
nand U14780 (N_14780,N_12905,N_12658);
nand U14781 (N_14781,N_12758,N_13386);
and U14782 (N_14782,N_12684,N_13553);
nand U14783 (N_14783,N_13606,N_12974);
xor U14784 (N_14784,N_13346,N_12847);
nand U14785 (N_14785,N_13744,N_12759);
or U14786 (N_14786,N_12798,N_12617);
nor U14787 (N_14787,N_12541,N_12893);
nor U14788 (N_14788,N_12844,N_13693);
or U14789 (N_14789,N_13184,N_13409);
nand U14790 (N_14790,N_13114,N_13533);
xor U14791 (N_14791,N_12654,N_13119);
nand U14792 (N_14792,N_13721,N_12513);
nor U14793 (N_14793,N_13190,N_13401);
xor U14794 (N_14794,N_13049,N_13251);
nand U14795 (N_14795,N_12550,N_12794);
nor U14796 (N_14796,N_13254,N_13113);
nor U14797 (N_14797,N_12685,N_12604);
and U14798 (N_14798,N_13432,N_13074);
or U14799 (N_14799,N_13427,N_12912);
nor U14800 (N_14800,N_12802,N_13510);
nand U14801 (N_14801,N_13024,N_13695);
and U14802 (N_14802,N_13151,N_13707);
or U14803 (N_14803,N_13728,N_12649);
xnor U14804 (N_14804,N_12961,N_13047);
nand U14805 (N_14805,N_12599,N_13642);
nand U14806 (N_14806,N_12861,N_13665);
and U14807 (N_14807,N_12501,N_12802);
and U14808 (N_14808,N_13065,N_13282);
or U14809 (N_14809,N_13708,N_13361);
nand U14810 (N_14810,N_13727,N_13589);
and U14811 (N_14811,N_12566,N_12510);
nand U14812 (N_14812,N_13173,N_12851);
or U14813 (N_14813,N_13713,N_13526);
or U14814 (N_14814,N_13165,N_12503);
nor U14815 (N_14815,N_13348,N_13173);
and U14816 (N_14816,N_12836,N_13051);
nor U14817 (N_14817,N_12620,N_13115);
and U14818 (N_14818,N_13076,N_13505);
or U14819 (N_14819,N_13434,N_12921);
and U14820 (N_14820,N_12776,N_13320);
xnor U14821 (N_14821,N_13426,N_13407);
xnor U14822 (N_14822,N_12959,N_13189);
nor U14823 (N_14823,N_13487,N_13512);
nor U14824 (N_14824,N_12524,N_13564);
and U14825 (N_14825,N_13477,N_13657);
nor U14826 (N_14826,N_12898,N_13149);
xor U14827 (N_14827,N_13717,N_12714);
nor U14828 (N_14828,N_13426,N_12631);
nor U14829 (N_14829,N_13550,N_13342);
nor U14830 (N_14830,N_13717,N_13346);
and U14831 (N_14831,N_13121,N_12600);
or U14832 (N_14832,N_13167,N_12704);
and U14833 (N_14833,N_13165,N_12720);
and U14834 (N_14834,N_13107,N_13410);
nor U14835 (N_14835,N_12539,N_13424);
or U14836 (N_14836,N_12941,N_13740);
and U14837 (N_14837,N_12952,N_13446);
nor U14838 (N_14838,N_13058,N_12786);
nand U14839 (N_14839,N_13262,N_13207);
nand U14840 (N_14840,N_12657,N_12981);
or U14841 (N_14841,N_12544,N_12840);
or U14842 (N_14842,N_13087,N_12766);
and U14843 (N_14843,N_12530,N_13244);
nor U14844 (N_14844,N_13607,N_13336);
nand U14845 (N_14845,N_12874,N_13005);
xor U14846 (N_14846,N_12674,N_12609);
xnor U14847 (N_14847,N_13597,N_13451);
or U14848 (N_14848,N_13005,N_13348);
and U14849 (N_14849,N_12963,N_13692);
xor U14850 (N_14850,N_12671,N_13182);
xnor U14851 (N_14851,N_13316,N_12725);
nor U14852 (N_14852,N_13412,N_13268);
nor U14853 (N_14853,N_13100,N_13113);
and U14854 (N_14854,N_12845,N_13593);
xnor U14855 (N_14855,N_12706,N_12569);
nor U14856 (N_14856,N_12732,N_13185);
nor U14857 (N_14857,N_12818,N_13200);
and U14858 (N_14858,N_12747,N_12918);
nand U14859 (N_14859,N_13026,N_13057);
or U14860 (N_14860,N_12943,N_13312);
or U14861 (N_14861,N_12506,N_13519);
nor U14862 (N_14862,N_12778,N_12508);
and U14863 (N_14863,N_12864,N_12740);
xnor U14864 (N_14864,N_13028,N_12685);
nand U14865 (N_14865,N_13585,N_12746);
xnor U14866 (N_14866,N_12562,N_13262);
and U14867 (N_14867,N_13747,N_13101);
and U14868 (N_14868,N_13475,N_13228);
xnor U14869 (N_14869,N_12634,N_13610);
or U14870 (N_14870,N_13006,N_12696);
xnor U14871 (N_14871,N_13555,N_13226);
nand U14872 (N_14872,N_12637,N_12944);
nand U14873 (N_14873,N_13601,N_12928);
nor U14874 (N_14874,N_12519,N_13095);
nand U14875 (N_14875,N_12565,N_13040);
or U14876 (N_14876,N_13175,N_13305);
and U14877 (N_14877,N_13455,N_13335);
nor U14878 (N_14878,N_12515,N_13034);
and U14879 (N_14879,N_12835,N_13169);
xnor U14880 (N_14880,N_13119,N_13708);
nand U14881 (N_14881,N_13221,N_13193);
xnor U14882 (N_14882,N_13143,N_12577);
nand U14883 (N_14883,N_13619,N_12557);
nor U14884 (N_14884,N_13692,N_12542);
and U14885 (N_14885,N_13005,N_12857);
xor U14886 (N_14886,N_13735,N_13647);
nand U14887 (N_14887,N_13114,N_13643);
or U14888 (N_14888,N_12958,N_13182);
xnor U14889 (N_14889,N_13431,N_12738);
and U14890 (N_14890,N_12680,N_13165);
or U14891 (N_14891,N_13502,N_13748);
nand U14892 (N_14892,N_12531,N_13206);
nand U14893 (N_14893,N_12837,N_13273);
xnor U14894 (N_14894,N_12554,N_12931);
nand U14895 (N_14895,N_13097,N_13287);
or U14896 (N_14896,N_13232,N_12987);
nand U14897 (N_14897,N_12722,N_12734);
xnor U14898 (N_14898,N_12652,N_13107);
nor U14899 (N_14899,N_13229,N_13036);
or U14900 (N_14900,N_13037,N_12674);
xor U14901 (N_14901,N_13571,N_13164);
and U14902 (N_14902,N_13143,N_13492);
and U14903 (N_14903,N_13566,N_13025);
xor U14904 (N_14904,N_12995,N_12941);
nand U14905 (N_14905,N_13138,N_12562);
nand U14906 (N_14906,N_12867,N_12902);
nand U14907 (N_14907,N_13450,N_13590);
xor U14908 (N_14908,N_12883,N_13413);
or U14909 (N_14909,N_12500,N_12753);
or U14910 (N_14910,N_13140,N_13422);
nand U14911 (N_14911,N_13277,N_13354);
or U14912 (N_14912,N_13376,N_12558);
and U14913 (N_14913,N_13486,N_12829);
nor U14914 (N_14914,N_13525,N_13538);
nand U14915 (N_14915,N_13289,N_13248);
or U14916 (N_14916,N_13303,N_13288);
nor U14917 (N_14917,N_13453,N_12574);
nand U14918 (N_14918,N_13335,N_12558);
or U14919 (N_14919,N_13655,N_12856);
or U14920 (N_14920,N_12542,N_12948);
or U14921 (N_14921,N_13355,N_13376);
or U14922 (N_14922,N_12504,N_12986);
nor U14923 (N_14923,N_12749,N_12768);
nor U14924 (N_14924,N_13523,N_13306);
nand U14925 (N_14925,N_13691,N_12571);
or U14926 (N_14926,N_12891,N_12616);
and U14927 (N_14927,N_12899,N_12625);
and U14928 (N_14928,N_13240,N_12697);
or U14929 (N_14929,N_13511,N_12982);
nand U14930 (N_14930,N_12964,N_13089);
xor U14931 (N_14931,N_12809,N_12930);
or U14932 (N_14932,N_13724,N_13413);
xor U14933 (N_14933,N_12702,N_13407);
and U14934 (N_14934,N_13413,N_12953);
xnor U14935 (N_14935,N_13663,N_13320);
xor U14936 (N_14936,N_13056,N_13270);
and U14937 (N_14937,N_12582,N_13619);
nor U14938 (N_14938,N_13262,N_13611);
nor U14939 (N_14939,N_13245,N_13696);
xor U14940 (N_14940,N_13321,N_12937);
nand U14941 (N_14941,N_12780,N_13185);
nor U14942 (N_14942,N_12979,N_13481);
nand U14943 (N_14943,N_12609,N_13288);
and U14944 (N_14944,N_12583,N_13263);
nand U14945 (N_14945,N_12537,N_12875);
nand U14946 (N_14946,N_13732,N_12920);
nor U14947 (N_14947,N_13445,N_13135);
or U14948 (N_14948,N_13010,N_12521);
or U14949 (N_14949,N_13555,N_13174);
nor U14950 (N_14950,N_13168,N_12570);
nor U14951 (N_14951,N_13572,N_12786);
or U14952 (N_14952,N_13558,N_13259);
nand U14953 (N_14953,N_12895,N_12528);
and U14954 (N_14954,N_12749,N_13421);
nand U14955 (N_14955,N_13225,N_13643);
xnor U14956 (N_14956,N_13151,N_13748);
or U14957 (N_14957,N_12700,N_13004);
nand U14958 (N_14958,N_12788,N_13031);
nand U14959 (N_14959,N_13106,N_13493);
nor U14960 (N_14960,N_13178,N_12905);
nand U14961 (N_14961,N_12672,N_12583);
xor U14962 (N_14962,N_12907,N_13204);
xnor U14963 (N_14963,N_13673,N_13541);
and U14964 (N_14964,N_13614,N_12826);
or U14965 (N_14965,N_13439,N_13145);
or U14966 (N_14966,N_13589,N_13134);
nor U14967 (N_14967,N_12993,N_13454);
and U14968 (N_14968,N_12808,N_13693);
nor U14969 (N_14969,N_13718,N_12806);
xor U14970 (N_14970,N_12573,N_12977);
xnor U14971 (N_14971,N_13665,N_12559);
nand U14972 (N_14972,N_13645,N_12915);
nor U14973 (N_14973,N_12746,N_12705);
xor U14974 (N_14974,N_13672,N_13240);
and U14975 (N_14975,N_12543,N_13488);
nor U14976 (N_14976,N_12524,N_13202);
or U14977 (N_14977,N_13113,N_12931);
nor U14978 (N_14978,N_13221,N_13101);
nand U14979 (N_14979,N_12746,N_13443);
or U14980 (N_14980,N_12878,N_13590);
xnor U14981 (N_14981,N_13674,N_12690);
nor U14982 (N_14982,N_13596,N_13109);
nand U14983 (N_14983,N_12893,N_12664);
nand U14984 (N_14984,N_13174,N_13575);
and U14985 (N_14985,N_12561,N_12949);
nor U14986 (N_14986,N_12580,N_13230);
nand U14987 (N_14987,N_12752,N_12585);
and U14988 (N_14988,N_13667,N_12841);
nor U14989 (N_14989,N_12770,N_12965);
xor U14990 (N_14990,N_13520,N_12827);
nand U14991 (N_14991,N_12708,N_13416);
and U14992 (N_14992,N_13483,N_12643);
nor U14993 (N_14993,N_12730,N_12947);
or U14994 (N_14994,N_13587,N_13605);
nor U14995 (N_14995,N_12845,N_13275);
and U14996 (N_14996,N_13412,N_13038);
nand U14997 (N_14997,N_13199,N_12853);
or U14998 (N_14998,N_13280,N_12720);
or U14999 (N_14999,N_12891,N_12523);
nand U15000 (N_15000,N_14164,N_14122);
and U15001 (N_15001,N_14475,N_14366);
nand U15002 (N_15002,N_14446,N_13977);
or U15003 (N_15003,N_14489,N_14363);
nand U15004 (N_15004,N_14135,N_13768);
and U15005 (N_15005,N_14666,N_14712);
nor U15006 (N_15006,N_14685,N_14546);
xnor U15007 (N_15007,N_14837,N_14725);
nand U15008 (N_15008,N_14360,N_14701);
or U15009 (N_15009,N_14005,N_14927);
or U15010 (N_15010,N_14581,N_14250);
nand U15011 (N_15011,N_14645,N_13872);
nor U15012 (N_15012,N_14562,N_14430);
and U15013 (N_15013,N_14415,N_13946);
nand U15014 (N_15014,N_14442,N_14450);
and U15015 (N_15015,N_14378,N_14447);
or U15016 (N_15016,N_14848,N_14989);
nor U15017 (N_15017,N_13811,N_14826);
or U15018 (N_15018,N_13806,N_13925);
xor U15019 (N_15019,N_14106,N_14256);
or U15020 (N_15020,N_14000,N_14977);
or U15021 (N_15021,N_14802,N_14011);
and U15022 (N_15022,N_13966,N_14290);
nand U15023 (N_15023,N_14845,N_14313);
and U15024 (N_15024,N_13762,N_14786);
or U15025 (N_15025,N_13964,N_14714);
nor U15026 (N_15026,N_13788,N_14723);
or U15027 (N_15027,N_14515,N_14706);
xnor U15028 (N_15028,N_14914,N_14864);
or U15029 (N_15029,N_14206,N_14688);
or U15030 (N_15030,N_14642,N_14964);
and U15031 (N_15031,N_14060,N_13996);
nand U15032 (N_15032,N_13873,N_13834);
nor U15033 (N_15033,N_14233,N_13961);
nand U15034 (N_15034,N_14208,N_14851);
or U15035 (N_15035,N_13984,N_14920);
nor U15036 (N_15036,N_14896,N_14844);
nor U15037 (N_15037,N_14391,N_14659);
nor U15038 (N_15038,N_13971,N_13945);
and U15039 (N_15039,N_14228,N_14283);
and U15040 (N_15040,N_14982,N_14083);
or U15041 (N_15041,N_13929,N_14089);
nand U15042 (N_15042,N_14909,N_13855);
xor U15043 (N_15043,N_14556,N_13876);
xor U15044 (N_15044,N_14879,N_13874);
xnor U15045 (N_15045,N_14308,N_14270);
nor U15046 (N_15046,N_14793,N_13827);
nor U15047 (N_15047,N_14003,N_14499);
or U15048 (N_15048,N_14080,N_13794);
xor U15049 (N_15049,N_14690,N_14486);
nor U15050 (N_15050,N_14856,N_13767);
or U15051 (N_15051,N_14763,N_14470);
nor U15052 (N_15052,N_14658,N_14697);
xnor U15053 (N_15053,N_14467,N_14154);
or U15054 (N_15054,N_14610,N_14040);
xor U15055 (N_15055,N_14631,N_14477);
or U15056 (N_15056,N_14820,N_14482);
nor U15057 (N_15057,N_13800,N_13804);
nand U15058 (N_15058,N_13771,N_14750);
and U15059 (N_15059,N_14739,N_13969);
or U15060 (N_15060,N_14133,N_14893);
or U15061 (N_15061,N_14299,N_14112);
nor U15062 (N_15062,N_14632,N_14376);
and U15063 (N_15063,N_14777,N_14109);
and U15064 (N_15064,N_14464,N_13956);
or U15065 (N_15065,N_14967,N_13932);
nand U15066 (N_15066,N_14812,N_14630);
xor U15067 (N_15067,N_14662,N_14531);
xor U15068 (N_15068,N_13941,N_14222);
nand U15069 (N_15069,N_14755,N_14996);
nor U15070 (N_15070,N_14311,N_14787);
or U15071 (N_15071,N_14413,N_14510);
and U15072 (N_15072,N_13928,N_14634);
xnor U15073 (N_15073,N_14722,N_13757);
nor U15074 (N_15074,N_14111,N_14936);
or U15075 (N_15075,N_14340,N_14751);
nor U15076 (N_15076,N_14301,N_14361);
nand U15077 (N_15077,N_14560,N_13993);
xor U15078 (N_15078,N_14226,N_13813);
nor U15079 (N_15079,N_14321,N_14871);
nor U15080 (N_15080,N_14661,N_14764);
nand U15081 (N_15081,N_14997,N_14128);
nor U15082 (N_15082,N_14325,N_13818);
and U15083 (N_15083,N_13991,N_14389);
nand U15084 (N_15084,N_13791,N_14036);
and U15085 (N_15085,N_14142,N_14139);
nor U15086 (N_15086,N_14455,N_13882);
nand U15087 (N_15087,N_14552,N_14564);
xor U15088 (N_15088,N_13820,N_14059);
nand U15089 (N_15089,N_14922,N_14589);
or U15090 (N_15090,N_14950,N_14935);
nand U15091 (N_15091,N_13973,N_14863);
xor U15092 (N_15092,N_13761,N_14292);
nor U15093 (N_15093,N_14492,N_14377);
nand U15094 (N_15094,N_13952,N_13892);
nor U15095 (N_15095,N_14409,N_14002);
xor U15096 (N_15096,N_14969,N_14229);
nand U15097 (N_15097,N_14561,N_14892);
nand U15098 (N_15098,N_14015,N_14624);
or U15099 (N_15099,N_13891,N_14992);
nand U15100 (N_15100,N_14370,N_14007);
and U15101 (N_15101,N_13825,N_14807);
or U15102 (N_15102,N_14792,N_14495);
or U15103 (N_15103,N_14437,N_14537);
nand U15104 (N_15104,N_14307,N_14454);
and U15105 (N_15105,N_13954,N_14588);
and U15106 (N_15106,N_13845,N_13755);
xor U15107 (N_15107,N_14490,N_14754);
xnor U15108 (N_15108,N_14058,N_14114);
xor U15109 (N_15109,N_14933,N_14113);
or U15110 (N_15110,N_14895,N_14282);
nor U15111 (N_15111,N_14648,N_14646);
and U15112 (N_15112,N_14772,N_14986);
xor U15113 (N_15113,N_14065,N_14506);
or U15114 (N_15114,N_14407,N_13784);
nor U15115 (N_15115,N_14733,N_14381);
nor U15116 (N_15116,N_14101,N_14861);
nand U15117 (N_15117,N_13870,N_14253);
xnor U15118 (N_15118,N_13766,N_13840);
xor U15119 (N_15119,N_13819,N_13986);
xor U15120 (N_15120,N_14432,N_14239);
xor U15121 (N_15121,N_14857,N_14877);
or U15122 (N_15122,N_14183,N_14636);
or U15123 (N_15123,N_14756,N_13817);
nand U15124 (N_15124,N_14882,N_14371);
or U15125 (N_15125,N_13979,N_14334);
or U15126 (N_15126,N_14358,N_13764);
nand U15127 (N_15127,N_14052,N_14219);
nor U15128 (N_15128,N_13888,N_14356);
nor U15129 (N_15129,N_14663,N_14513);
nand U15130 (N_15130,N_14461,N_14126);
xor U15131 (N_15131,N_14074,N_14343);
and U15132 (N_15132,N_13894,N_14266);
xor U15133 (N_15133,N_14887,N_14988);
or U15134 (N_15134,N_14993,N_14459);
nand U15135 (N_15135,N_14070,N_14951);
and U15136 (N_15136,N_14500,N_14008);
nor U15137 (N_15137,N_14053,N_13812);
and U15138 (N_15138,N_14818,N_14766);
nor U15139 (N_15139,N_14593,N_13793);
nor U15140 (N_15140,N_14641,N_14584);
and U15141 (N_15141,N_14880,N_14251);
or U15142 (N_15142,N_14152,N_14130);
nor U15143 (N_15143,N_14110,N_14274);
or U15144 (N_15144,N_14453,N_14519);
or U15145 (N_15145,N_14627,N_14039);
nand U15146 (N_15146,N_14265,N_14141);
nor U15147 (N_15147,N_14921,N_14380);
or U15148 (N_15148,N_14606,N_14717);
xnor U15149 (N_15149,N_14966,N_13854);
nand U15150 (N_15150,N_14682,N_14819);
or U15151 (N_15151,N_14474,N_14840);
or U15152 (N_15152,N_13939,N_14201);
nor U15153 (N_15153,N_14276,N_14277);
xor U15154 (N_15154,N_14651,N_14230);
or U15155 (N_15155,N_14973,N_14735);
or U15156 (N_15156,N_14924,N_14899);
or U15157 (N_15157,N_13783,N_14720);
or U15158 (N_15158,N_13948,N_13871);
and U15159 (N_15159,N_14210,N_14695);
xor U15160 (N_15160,N_14497,N_14801);
nand U15161 (N_15161,N_14910,N_14445);
xor U15162 (N_15162,N_14509,N_14087);
and U15163 (N_15163,N_14945,N_14468);
and U15164 (N_15164,N_14255,N_14758);
nand U15165 (N_15165,N_13824,N_14412);
or U15166 (N_15166,N_14131,N_14719);
nand U15167 (N_15167,N_14403,N_14832);
or U15168 (N_15168,N_14320,N_14994);
nand U15169 (N_15169,N_14440,N_14779);
and U15170 (N_15170,N_13864,N_14709);
nand U15171 (N_15171,N_14852,N_14189);
and U15172 (N_15172,N_14638,N_14429);
and U15173 (N_15173,N_14349,N_14512);
or U15174 (N_15174,N_13885,N_14280);
and U15175 (N_15175,N_13769,N_14273);
or U15176 (N_15176,N_14516,N_14171);
nand U15177 (N_15177,N_14557,N_14215);
nor U15178 (N_15178,N_13786,N_14035);
and U15179 (N_15179,N_13797,N_14637);
xnor U15180 (N_15180,N_14975,N_14049);
and U15181 (N_15181,N_14175,N_14622);
nand U15182 (N_15182,N_14505,N_14703);
nand U15183 (N_15183,N_14140,N_14684);
nand U15184 (N_15184,N_14607,N_13918);
or U15185 (N_15185,N_14948,N_14245);
and U15186 (N_15186,N_14894,N_14125);
or U15187 (N_15187,N_14212,N_14158);
or U15188 (N_15188,N_14385,N_14835);
xor U15189 (N_15189,N_13987,N_14991);
xnor U15190 (N_15190,N_13897,N_14958);
or U15191 (N_15191,N_14476,N_14119);
and U15192 (N_15192,N_14773,N_14196);
and U15193 (N_15193,N_14174,N_14176);
nand U15194 (N_15194,N_14088,N_13799);
nor U15195 (N_15195,N_14309,N_14932);
and U15196 (N_15196,N_14872,N_14738);
xor U15197 (N_15197,N_14300,N_14514);
and U15198 (N_15198,N_13934,N_14466);
nand U15199 (N_15199,N_13865,N_14554);
or U15200 (N_15200,N_14165,N_14760);
xor U15201 (N_15201,N_14314,N_14145);
nor U15202 (N_15202,N_14286,N_13990);
nor U15203 (N_15203,N_13849,N_14368);
nand U15204 (N_15204,N_14567,N_14535);
or U15205 (N_15205,N_14783,N_14785);
or U15206 (N_15206,N_14649,N_14704);
or U15207 (N_15207,N_14328,N_13828);
nand U15208 (N_15208,N_14191,N_14677);
or U15209 (N_15209,N_14424,N_14116);
nor U15210 (N_15210,N_14383,N_14788);
xnor U15211 (N_15211,N_14103,N_14740);
xor U15212 (N_15212,N_13822,N_14451);
xnor U15213 (N_15213,N_14615,N_14798);
and U15214 (N_15214,N_13867,N_14107);
or U15215 (N_15215,N_14326,N_14898);
nand U15216 (N_15216,N_13949,N_14743);
or U15217 (N_15217,N_14906,N_14435);
nor U15218 (N_15218,N_13982,N_14578);
xnor U15219 (N_15219,N_13751,N_14582);
nand U15220 (N_15220,N_13866,N_14876);
and U15221 (N_15221,N_14179,N_14796);
nand U15222 (N_15222,N_14414,N_14518);
and U15223 (N_15223,N_13781,N_13816);
xor U15224 (N_15224,N_14938,N_14547);
nand U15225 (N_15225,N_14726,N_14124);
nand U15226 (N_15226,N_14504,N_14207);
or U15227 (N_15227,N_13779,N_14318);
or U15228 (N_15228,N_14134,N_14843);
and U15229 (N_15229,N_13838,N_14665);
nor U15230 (N_15230,N_13943,N_14972);
nand U15231 (N_15231,N_14285,N_14747);
and U15232 (N_15232,N_14260,N_14946);
nor U15233 (N_15233,N_14185,N_14616);
nor U15234 (N_15234,N_14243,N_14327);
or U15235 (N_15235,N_13841,N_13907);
xnor U15236 (N_15236,N_14617,N_14332);
or U15237 (N_15237,N_14971,N_14753);
xor U15238 (N_15238,N_14168,N_14350);
xor U15239 (N_15239,N_14604,N_13868);
or U15240 (N_15240,N_13980,N_14050);
nor U15241 (N_15241,N_14941,N_14485);
and U15242 (N_15242,N_14092,N_14017);
nor U15243 (N_15243,N_14242,N_14548);
or U15244 (N_15244,N_14231,N_14120);
and U15245 (N_15245,N_14064,N_14408);
xor U15246 (N_15246,N_14803,N_14540);
nor U15247 (N_15247,N_14528,N_14190);
and U15248 (N_15248,N_13947,N_14322);
xor U15249 (N_15249,N_14043,N_14744);
and U15250 (N_15250,N_14472,N_14655);
nor U15251 (N_15251,N_14082,N_14965);
or U15252 (N_15252,N_14503,N_14267);
or U15253 (N_15253,N_14691,N_14683);
nand U15254 (N_15254,N_14978,N_13860);
nor U15255 (N_15255,N_14170,N_14599);
and U15256 (N_15256,N_14609,N_13940);
nand U15257 (N_15257,N_14063,N_14729);
nor U15258 (N_15258,N_13837,N_14187);
xor U15259 (N_15259,N_14700,N_14962);
nor U15260 (N_15260,N_14078,N_14484);
nor U15261 (N_15261,N_13878,N_14374);
nor U15262 (N_15262,N_13758,N_13992);
nor U15263 (N_15263,N_14269,N_13808);
xor U15264 (N_15264,N_14223,N_13875);
nor U15265 (N_15265,N_14192,N_14865);
nand U15266 (N_15266,N_13750,N_14998);
xnor U15267 (N_15267,N_14066,N_14227);
nand U15268 (N_15268,N_14100,N_13859);
nor U15269 (N_15269,N_14335,N_14029);
nor U15270 (N_15270,N_14569,N_13908);
nand U15271 (N_15271,N_14724,N_14940);
or U15272 (N_15272,N_14883,N_14947);
nor U15273 (N_15273,N_14944,N_13778);
or U15274 (N_15274,N_14182,N_14317);
xnor U15275 (N_15275,N_14902,N_13848);
nand U15276 (N_15276,N_14960,N_13944);
and U15277 (N_15277,N_14153,N_14713);
xor U15278 (N_15278,N_14652,N_13974);
nand U15279 (N_15279,N_14316,N_14157);
or U15280 (N_15280,N_14853,N_14258);
nor U15281 (N_15281,N_13917,N_14224);
or U15282 (N_15282,N_13883,N_14937);
and U15283 (N_15283,N_14601,N_14791);
nor U15284 (N_15284,N_14384,N_14888);
nand U15285 (N_15285,N_14728,N_14983);
xnor U15286 (N_15286,N_14592,N_14585);
or U15287 (N_15287,N_14021,N_13965);
xor U15288 (N_15288,N_14167,N_13815);
nand U15289 (N_15289,N_14331,N_14248);
or U15290 (N_15290,N_14911,N_14889);
and U15291 (N_15291,N_13905,N_14395);
xnor U15292 (N_15292,N_14716,N_14054);
or U15293 (N_15293,N_14048,N_14108);
nand U15294 (N_15294,N_13893,N_14770);
nor U15295 (N_15295,N_13842,N_14970);
or U15296 (N_15296,N_14341,N_14929);
xor U15297 (N_15297,N_14344,N_14479);
xnor U15298 (N_15298,N_14875,N_14220);
and U15299 (N_15299,N_14668,N_14433);
nand U15300 (N_15300,N_14047,N_14918);
nor U15301 (N_15301,N_14338,N_14545);
nor U15302 (N_15302,N_14913,N_14759);
or U15303 (N_15303,N_14781,N_14102);
nand U15304 (N_15304,N_14062,N_13836);
nor U15305 (N_15305,N_14055,N_14057);
xor U15306 (N_15306,N_14908,N_14004);
or U15307 (N_15307,N_14247,N_14869);
or U15308 (N_15308,N_14069,N_14836);
nand U15309 (N_15309,N_14833,N_14394);
or U15310 (N_15310,N_14254,N_14073);
and U15311 (N_15311,N_14386,N_14841);
and U15312 (N_15312,N_14854,N_14001);
nor U15313 (N_15313,N_14521,N_13989);
nor U15314 (N_15314,N_14502,N_13881);
xor U15315 (N_15315,N_14912,N_13858);
nand U15316 (N_15316,N_14752,N_14161);
or U15317 (N_15317,N_14094,N_13765);
nor U15318 (N_15318,N_13937,N_14775);
and U15319 (N_15319,N_13752,N_14602);
and U15320 (N_15320,N_14917,N_14794);
or U15321 (N_15321,N_14498,N_14193);
and U15322 (N_15322,N_13920,N_14399);
nor U15323 (N_15323,N_14985,N_14959);
or U15324 (N_15324,N_14372,N_14225);
or U15325 (N_15325,N_14839,N_14046);
or U15326 (N_15326,N_14693,N_14232);
and U15327 (N_15327,N_14427,N_14473);
and U15328 (N_15328,N_13998,N_14890);
nand U15329 (N_15329,N_13904,N_13913);
or U15330 (N_15330,N_14213,N_14767);
xor U15331 (N_15331,N_14732,N_13844);
nor U15332 (N_15332,N_14354,N_14188);
and U15333 (N_15333,N_14692,N_14426);
or U15334 (N_15334,N_14822,N_14550);
nor U15335 (N_15335,N_14268,N_14626);
or U15336 (N_15336,N_14132,N_14897);
xor U15337 (N_15337,N_14653,N_14603);
and U15338 (N_15338,N_14949,N_13953);
xnor U15339 (N_15339,N_14681,N_14810);
nor U15340 (N_15340,N_14707,N_14180);
or U15341 (N_15341,N_14587,N_14401);
or U15342 (N_15342,N_14974,N_14397);
xnor U15343 (N_15343,N_13889,N_14469);
and U15344 (N_15344,N_14072,N_14579);
nor U15345 (N_15345,N_14298,N_14353);
and U15346 (N_15346,N_14037,N_13803);
or U15347 (N_15347,N_14352,N_14705);
nor U15348 (N_15348,N_13899,N_14980);
nand U15349 (N_15349,N_14644,N_14237);
nand U15350 (N_15350,N_14900,N_13775);
nand U15351 (N_15351,N_14137,N_14806);
and U15352 (N_15352,N_14821,N_13903);
nor U15353 (N_15353,N_14769,N_13985);
nand U15354 (N_15354,N_14202,N_14302);
nor U15355 (N_15355,N_13785,N_13770);
nor U15356 (N_15356,N_13886,N_14392);
or U15357 (N_15357,N_14388,N_14675);
and U15358 (N_15358,N_14571,N_13909);
xor U15359 (N_15359,N_14006,N_14151);
nor U15360 (N_15360,N_14942,N_14874);
nor U15361 (N_15361,N_13843,N_14214);
xnor U15362 (N_15362,N_13853,N_14923);
nor U15363 (N_15363,N_14359,N_14934);
and U15364 (N_15364,N_14041,N_14155);
or U15365 (N_15365,N_14099,N_14824);
nand U15366 (N_15366,N_14211,N_14337);
nor U15367 (N_15367,N_13995,N_14081);
nor U15368 (N_15368,N_14811,N_14995);
or U15369 (N_15369,N_14981,N_14591);
and U15370 (N_15370,N_14625,N_14291);
and U15371 (N_15371,N_14218,N_14526);
and U15372 (N_15372,N_14621,N_14529);
and U15373 (N_15373,N_14533,N_14357);
nor U15374 (N_15374,N_13839,N_14611);
nor U15375 (N_15375,N_14774,N_14575);
nand U15376 (N_15376,N_14375,N_14252);
or U15377 (N_15377,N_14804,N_13776);
nor U15378 (N_15378,N_13895,N_14742);
xnor U15379 (N_15379,N_14249,N_14650);
xnor U15380 (N_15380,N_14431,N_14441);
nand U15381 (N_15381,N_13798,N_14838);
or U15382 (N_15382,N_13959,N_14159);
nor U15383 (N_15383,N_14272,N_14295);
or U15384 (N_15384,N_14595,N_14471);
nor U15385 (N_15385,N_14095,N_14566);
xor U15386 (N_15386,N_14369,N_14680);
nand U15387 (N_15387,N_14708,N_14024);
and U15388 (N_15388,N_13830,N_14961);
nand U15389 (N_15389,N_14045,N_14768);
or U15390 (N_15390,N_14574,N_14448);
or U15391 (N_15391,N_13805,N_13774);
nand U15392 (N_15392,N_13950,N_13763);
and U15393 (N_15393,N_14289,N_14831);
nand U15394 (N_15394,N_14079,N_14163);
and U15395 (N_15395,N_13877,N_13922);
nor U15396 (N_15396,N_14138,N_14365);
nand U15397 (N_15397,N_13923,N_13862);
and U15398 (N_15398,N_14396,N_14460);
and U15399 (N_15399,N_13958,N_14678);
nand U15400 (N_15400,N_14629,N_14699);
xnor U15401 (N_15401,N_14957,N_14926);
nand U15402 (N_15402,N_14178,N_14979);
nand U15403 (N_15403,N_13898,N_13829);
nand U15404 (N_15404,N_13857,N_14643);
and U15405 (N_15405,N_14860,N_14782);
nand U15406 (N_15406,N_13810,N_14905);
xor U15407 (N_15407,N_14026,N_14023);
or U15408 (N_15408,N_14362,N_14881);
nor U15409 (N_15409,N_14034,N_13994);
xor U15410 (N_15410,N_14815,N_14056);
and U15411 (N_15411,N_14698,N_14315);
xnor U15412 (N_15412,N_14449,N_13890);
nand U15413 (N_15413,N_13955,N_14746);
and U15414 (N_15414,N_14736,N_14689);
xor U15415 (N_15415,N_14789,N_14999);
nor U15416 (N_15416,N_14907,N_13802);
xnor U15417 (N_15417,N_13963,N_13912);
nand U15418 (N_15418,N_14930,N_13821);
xnor U15419 (N_15419,N_14757,N_14613);
nor U15420 (N_15420,N_14954,N_14730);
or U15421 (N_15421,N_14238,N_13823);
nor U15422 (N_15422,N_13833,N_14493);
or U15423 (N_15423,N_14790,N_14085);
nand U15424 (N_15424,N_14419,N_14762);
nand U15425 (N_15425,N_14823,N_14136);
or U15426 (N_15426,N_14203,N_14955);
nand U15427 (N_15427,N_14197,N_14886);
or U15428 (N_15428,N_14576,N_13911);
nor U15429 (N_15429,N_13826,N_14373);
and U15430 (N_15430,N_14012,N_14071);
and U15431 (N_15431,N_14127,N_14205);
and U15432 (N_15432,N_14076,N_14259);
xor U15433 (N_15433,N_14425,N_14778);
xor U15434 (N_15434,N_14532,N_14633);
nor U15435 (N_15435,N_14329,N_14184);
or U15436 (N_15436,N_14244,N_14013);
nand U15437 (N_15437,N_14143,N_14097);
or U15438 (N_15438,N_13983,N_14016);
nand U15439 (N_15439,N_14508,N_14925);
xnor U15440 (N_15440,N_14568,N_14204);
nand U15441 (N_15441,N_14421,N_14828);
nand U15442 (N_15442,N_13852,N_14808);
xnor U15443 (N_15443,N_14916,N_14118);
nand U15444 (N_15444,N_14236,N_14261);
nor U15445 (N_15445,N_14452,N_14846);
or U15446 (N_15446,N_14483,N_14855);
or U15447 (N_15447,N_14813,N_14780);
or U15448 (N_15448,N_14620,N_14271);
and U15449 (N_15449,N_14339,N_14075);
nor U15450 (N_15450,N_14186,N_14600);
xnor U15451 (N_15451,N_14639,N_14849);
nor U15452 (N_15452,N_14160,N_13777);
xnor U15453 (N_15453,N_14827,N_13851);
nand U15454 (N_15454,N_13773,N_14195);
or U15455 (N_15455,N_14590,N_14166);
nor U15456 (N_15456,N_14393,N_14553);
xor U15457 (N_15457,N_13967,N_14799);
nor U15458 (N_15458,N_14891,N_13931);
and U15459 (N_15459,N_14549,N_14061);
nand U15460 (N_15460,N_14246,N_14303);
or U15461 (N_15461,N_14146,N_14367);
nand U15462 (N_15462,N_14858,N_14830);
nand U15463 (N_15463,N_14398,N_13902);
nor U15464 (N_15464,N_13962,N_14198);
and U15465 (N_15465,N_14987,N_14333);
nor U15466 (N_15466,N_14465,N_14517);
or U15467 (N_15467,N_14859,N_14458);
or U15468 (N_15468,N_14323,N_14169);
or U15469 (N_15469,N_14953,N_14669);
or U15470 (N_15470,N_14084,N_13756);
xnor U15471 (N_15471,N_14077,N_14541);
or U15472 (N_15472,N_14847,N_14814);
nor U15473 (N_15473,N_14117,N_14534);
nor U15474 (N_15474,N_14672,N_14288);
nand U15475 (N_15475,N_13936,N_14022);
and U15476 (N_15476,N_14121,N_14020);
and U15477 (N_15477,N_14287,N_13960);
xor U15478 (N_15478,N_14647,N_14150);
and U15479 (N_15479,N_14850,N_14028);
nand U15480 (N_15480,N_14216,N_13814);
nor U15481 (N_15481,N_13951,N_14051);
xnor U15482 (N_15482,N_14586,N_14542);
xor U15483 (N_15483,N_14727,N_14319);
nand U15484 (N_15484,N_14093,N_13919);
and U15485 (N_15485,N_14784,N_14086);
nand U15486 (N_15486,N_14748,N_13968);
nor U15487 (N_15487,N_14594,N_13792);
and U15488 (N_15488,N_14640,N_14217);
xnor U15489 (N_15489,N_14619,N_14355);
and U15490 (N_15490,N_14456,N_14968);
nor U15491 (N_15491,N_14067,N_14731);
nand U15492 (N_15492,N_14156,N_14664);
nor U15493 (N_15493,N_14771,N_14221);
xnor U15494 (N_15494,N_14524,N_14200);
and U15495 (N_15495,N_13915,N_14737);
nor U15496 (N_15496,N_14660,N_14346);
or U15497 (N_15497,N_13832,N_13831);
xor U15498 (N_15498,N_14539,N_14522);
or U15499 (N_15499,N_14281,N_14105);
nor U15500 (N_15500,N_14296,N_13921);
or U15501 (N_15501,N_14654,N_14928);
or U15502 (N_15502,N_14177,N_14009);
nor U15503 (N_15503,N_14596,N_14612);
nor U15504 (N_15504,N_14293,N_14817);
nor U15505 (N_15505,N_14149,N_14410);
or U15506 (N_15506,N_14657,N_14598);
or U15507 (N_15507,N_14573,N_13930);
nand U15508 (N_15508,N_14463,N_14129);
nand U15509 (N_15509,N_14104,N_14931);
and U15510 (N_15510,N_14749,N_14294);
nand U15511 (N_15511,N_14402,N_14147);
nand U15512 (N_15512,N_14297,N_14558);
nor U15513 (N_15513,N_14867,N_14873);
and U15514 (N_15514,N_14976,N_13935);
nor U15515 (N_15515,N_13807,N_13927);
nor U15516 (N_15516,N_14364,N_14525);
nand U15517 (N_15517,N_14347,N_14527);
or U15518 (N_15518,N_13988,N_13942);
and U15519 (N_15519,N_14496,N_14765);
xnor U15520 (N_15520,N_14702,N_14800);
xnor U15521 (N_15521,N_14656,N_14538);
nand U15522 (N_15522,N_14884,N_13900);
and U15523 (N_15523,N_13887,N_13809);
nand U15524 (N_15524,N_14241,N_14199);
and U15525 (N_15525,N_14304,N_13772);
nand U15526 (N_15526,N_14903,N_14842);
nand U15527 (N_15527,N_14551,N_14491);
nor U15528 (N_15528,N_13924,N_14511);
nor U15529 (N_15529,N_14032,N_14943);
nand U15530 (N_15530,N_14543,N_14257);
nor U15531 (N_15531,N_13976,N_14565);
xor U15532 (N_15532,N_14530,N_14330);
nor U15533 (N_15533,N_14834,N_14809);
nor U15534 (N_15534,N_13790,N_14608);
xor U15535 (N_15535,N_14278,N_14919);
xnor U15536 (N_15536,N_14577,N_13938);
nor U15537 (N_15537,N_14348,N_13753);
or U15538 (N_15538,N_14400,N_14027);
nor U15539 (N_15539,N_14878,N_14123);
nand U15540 (N_15540,N_14605,N_13869);
nand U15541 (N_15541,N_14444,N_14324);
or U15542 (N_15542,N_14162,N_14305);
nor U15543 (N_15543,N_14462,N_14181);
nand U15544 (N_15544,N_13787,N_14382);
or U15545 (N_15545,N_14715,N_13847);
xor U15546 (N_15546,N_13782,N_14336);
xor U15547 (N_15547,N_14711,N_14956);
nand U15548 (N_15548,N_14572,N_14696);
or U15549 (N_15549,N_14488,N_14096);
xor U15550 (N_15550,N_14901,N_14033);
or U15551 (N_15551,N_14673,N_14379);
and U15552 (N_15552,N_14406,N_14570);
or U15553 (N_15553,N_14115,N_14068);
nor U15554 (N_15554,N_14718,N_14523);
or U15555 (N_15555,N_14679,N_14721);
and U15556 (N_15556,N_13933,N_14172);
or U15557 (N_15557,N_14862,N_14583);
and U15558 (N_15558,N_14434,N_14443);
or U15559 (N_15559,N_14091,N_13796);
and U15560 (N_15560,N_14939,N_13901);
nand U15561 (N_15561,N_13926,N_13972);
xnor U15562 (N_15562,N_14417,N_14555);
nor U15563 (N_15563,N_14031,N_13795);
or U15564 (N_15564,N_14507,N_14984);
nand U15565 (N_15565,N_14480,N_14345);
nand U15566 (N_15566,N_14494,N_14310);
xnor U15567 (N_15567,N_14306,N_14671);
or U15568 (N_15568,N_13906,N_14025);
and U15569 (N_15569,N_14687,N_14262);
or U15570 (N_15570,N_14284,N_14423);
nor U15571 (N_15571,N_13879,N_13975);
xor U15572 (N_15572,N_13910,N_13884);
nor U15573 (N_15573,N_14618,N_13780);
and U15574 (N_15574,N_14428,N_14420);
xnor U15575 (N_15575,N_14580,N_14623);
or U15576 (N_15576,N_13999,N_14148);
xor U15577 (N_15577,N_14829,N_14904);
and U15578 (N_15578,N_14098,N_14915);
nor U15579 (N_15579,N_14816,N_14795);
nor U15580 (N_15580,N_14544,N_14275);
nand U15581 (N_15581,N_14390,N_14635);
or U15582 (N_15582,N_14825,N_14870);
nand U15583 (N_15583,N_14279,N_13861);
nor U15584 (N_15584,N_14209,N_14351);
or U15585 (N_15585,N_14481,N_14797);
and U15586 (N_15586,N_13880,N_14439);
nor U15587 (N_15587,N_14487,N_14411);
xnor U15588 (N_15588,N_14312,N_14990);
or U15589 (N_15589,N_14019,N_14240);
or U15590 (N_15590,N_14416,N_13846);
or U15591 (N_15591,N_13997,N_14090);
or U15592 (N_15592,N_14194,N_14776);
xor U15593 (N_15593,N_14342,N_13754);
and U15594 (N_15594,N_14734,N_14418);
nand U15595 (N_15595,N_14520,N_13760);
nand U15596 (N_15596,N_14044,N_14038);
nand U15597 (N_15597,N_13759,N_14710);
nand U15598 (N_15598,N_13801,N_13856);
nor U15599 (N_15599,N_14457,N_14422);
nand U15600 (N_15600,N_14670,N_13850);
nand U15601 (N_15601,N_14597,N_13863);
and U15602 (N_15602,N_14694,N_14866);
nand U15603 (N_15603,N_14404,N_14436);
nor U15604 (N_15604,N_14761,N_14676);
and U15605 (N_15605,N_14234,N_14478);
or U15606 (N_15606,N_14010,N_14042);
nand U15607 (N_15607,N_13789,N_13914);
and U15608 (N_15608,N_14667,N_13916);
and U15609 (N_15609,N_14674,N_13978);
or U15610 (N_15610,N_14885,N_14559);
or U15611 (N_15611,N_13970,N_14018);
or U15612 (N_15612,N_14387,N_14868);
and U15613 (N_15613,N_14741,N_14952);
and U15614 (N_15614,N_14628,N_13835);
xor U15615 (N_15615,N_14235,N_14144);
nor U15616 (N_15616,N_14501,N_14030);
and U15617 (N_15617,N_13957,N_13896);
nor U15618 (N_15618,N_14173,N_14745);
or U15619 (N_15619,N_14536,N_13981);
and U15620 (N_15620,N_14963,N_14405);
nor U15621 (N_15621,N_14563,N_14263);
xor U15622 (N_15622,N_14805,N_14014);
nand U15623 (N_15623,N_14686,N_14438);
or U15624 (N_15624,N_14264,N_14614);
xor U15625 (N_15625,N_14684,N_14074);
xnor U15626 (N_15626,N_13776,N_13813);
or U15627 (N_15627,N_14063,N_14613);
and U15628 (N_15628,N_14896,N_14519);
xnor U15629 (N_15629,N_14031,N_14275);
xor U15630 (N_15630,N_14885,N_14970);
or U15631 (N_15631,N_14344,N_14382);
nand U15632 (N_15632,N_13861,N_14435);
nor U15633 (N_15633,N_14822,N_14719);
and U15634 (N_15634,N_14389,N_14456);
or U15635 (N_15635,N_14537,N_14351);
nand U15636 (N_15636,N_14261,N_14699);
nor U15637 (N_15637,N_14162,N_14730);
or U15638 (N_15638,N_13995,N_14988);
and U15639 (N_15639,N_14652,N_14997);
or U15640 (N_15640,N_13764,N_14179);
xor U15641 (N_15641,N_14381,N_14770);
and U15642 (N_15642,N_14496,N_13969);
or U15643 (N_15643,N_14294,N_14335);
xnor U15644 (N_15644,N_14974,N_14759);
and U15645 (N_15645,N_14394,N_14131);
nand U15646 (N_15646,N_14776,N_14372);
nand U15647 (N_15647,N_13870,N_14593);
and U15648 (N_15648,N_14033,N_13761);
xor U15649 (N_15649,N_14989,N_14479);
and U15650 (N_15650,N_14052,N_14534);
or U15651 (N_15651,N_14099,N_13956);
and U15652 (N_15652,N_14258,N_14912);
or U15653 (N_15653,N_14943,N_14875);
xor U15654 (N_15654,N_14966,N_14346);
or U15655 (N_15655,N_14373,N_14008);
nor U15656 (N_15656,N_14609,N_14770);
nand U15657 (N_15657,N_14800,N_14299);
and U15658 (N_15658,N_14793,N_14974);
and U15659 (N_15659,N_14367,N_14553);
or U15660 (N_15660,N_14521,N_13824);
xnor U15661 (N_15661,N_14979,N_14770);
xnor U15662 (N_15662,N_13997,N_14014);
nand U15663 (N_15663,N_14001,N_14384);
xor U15664 (N_15664,N_14390,N_13813);
and U15665 (N_15665,N_14405,N_14227);
and U15666 (N_15666,N_14324,N_14877);
nand U15667 (N_15667,N_13778,N_14588);
nand U15668 (N_15668,N_13900,N_14300);
nand U15669 (N_15669,N_14223,N_13862);
or U15670 (N_15670,N_14602,N_14730);
xor U15671 (N_15671,N_14986,N_14818);
and U15672 (N_15672,N_13863,N_14577);
and U15673 (N_15673,N_14338,N_14259);
and U15674 (N_15674,N_14352,N_14554);
or U15675 (N_15675,N_14472,N_14157);
nand U15676 (N_15676,N_14157,N_13836);
nor U15677 (N_15677,N_14316,N_14539);
or U15678 (N_15678,N_14367,N_14686);
or U15679 (N_15679,N_14217,N_14598);
xnor U15680 (N_15680,N_13765,N_14021);
nand U15681 (N_15681,N_14459,N_14085);
nor U15682 (N_15682,N_14096,N_14730);
or U15683 (N_15683,N_13928,N_13976);
nand U15684 (N_15684,N_13859,N_14117);
or U15685 (N_15685,N_14722,N_14148);
or U15686 (N_15686,N_14062,N_13842);
nand U15687 (N_15687,N_14583,N_13825);
or U15688 (N_15688,N_14667,N_14627);
nand U15689 (N_15689,N_14367,N_14629);
and U15690 (N_15690,N_13759,N_14428);
nor U15691 (N_15691,N_13801,N_14902);
xnor U15692 (N_15692,N_14498,N_13940);
or U15693 (N_15693,N_14866,N_14821);
nand U15694 (N_15694,N_14566,N_14559);
and U15695 (N_15695,N_13973,N_13871);
or U15696 (N_15696,N_14198,N_14810);
xnor U15697 (N_15697,N_14165,N_14308);
nor U15698 (N_15698,N_14778,N_14871);
nand U15699 (N_15699,N_13785,N_14823);
nor U15700 (N_15700,N_13768,N_13904);
and U15701 (N_15701,N_14360,N_14594);
nor U15702 (N_15702,N_13996,N_14792);
or U15703 (N_15703,N_14821,N_14353);
xor U15704 (N_15704,N_14774,N_13987);
and U15705 (N_15705,N_14384,N_13833);
nor U15706 (N_15706,N_13834,N_14329);
and U15707 (N_15707,N_14620,N_13835);
or U15708 (N_15708,N_14450,N_13977);
nand U15709 (N_15709,N_14852,N_14599);
xnor U15710 (N_15710,N_14636,N_13813);
xor U15711 (N_15711,N_13912,N_14401);
nor U15712 (N_15712,N_14787,N_14036);
xor U15713 (N_15713,N_14987,N_13887);
xnor U15714 (N_15714,N_14514,N_13975);
and U15715 (N_15715,N_14908,N_13937);
xor U15716 (N_15716,N_14419,N_14617);
nand U15717 (N_15717,N_14007,N_14648);
nor U15718 (N_15718,N_13941,N_13761);
xor U15719 (N_15719,N_13882,N_14572);
nand U15720 (N_15720,N_14090,N_14713);
and U15721 (N_15721,N_14984,N_14192);
xor U15722 (N_15722,N_14040,N_14890);
nor U15723 (N_15723,N_14658,N_14455);
nand U15724 (N_15724,N_14657,N_14578);
nor U15725 (N_15725,N_13762,N_14189);
nor U15726 (N_15726,N_13912,N_14244);
nor U15727 (N_15727,N_14362,N_14399);
and U15728 (N_15728,N_14176,N_14608);
nor U15729 (N_15729,N_14021,N_14320);
nand U15730 (N_15730,N_14524,N_14017);
and U15731 (N_15731,N_13894,N_14236);
or U15732 (N_15732,N_14421,N_14519);
or U15733 (N_15733,N_14284,N_14760);
nor U15734 (N_15734,N_14882,N_14023);
nor U15735 (N_15735,N_14206,N_14112);
nand U15736 (N_15736,N_13896,N_13835);
nor U15737 (N_15737,N_14679,N_14086);
and U15738 (N_15738,N_13783,N_14987);
xor U15739 (N_15739,N_14531,N_14202);
and U15740 (N_15740,N_14289,N_14507);
nand U15741 (N_15741,N_14812,N_13798);
nand U15742 (N_15742,N_14153,N_14603);
or U15743 (N_15743,N_14711,N_14715);
nor U15744 (N_15744,N_14806,N_14331);
nor U15745 (N_15745,N_14223,N_14821);
nor U15746 (N_15746,N_14574,N_14600);
xor U15747 (N_15747,N_14991,N_14838);
nand U15748 (N_15748,N_13890,N_13937);
and U15749 (N_15749,N_14488,N_14776);
or U15750 (N_15750,N_14350,N_14577);
xor U15751 (N_15751,N_14809,N_14110);
and U15752 (N_15752,N_14011,N_14641);
or U15753 (N_15753,N_14940,N_14363);
xnor U15754 (N_15754,N_13878,N_14643);
xor U15755 (N_15755,N_14535,N_14674);
or U15756 (N_15756,N_14759,N_14643);
nor U15757 (N_15757,N_14005,N_13943);
xnor U15758 (N_15758,N_14177,N_14682);
or U15759 (N_15759,N_14276,N_14916);
and U15760 (N_15760,N_14067,N_14541);
or U15761 (N_15761,N_14274,N_14572);
nor U15762 (N_15762,N_14848,N_14030);
and U15763 (N_15763,N_14588,N_14253);
nor U15764 (N_15764,N_13933,N_14926);
nand U15765 (N_15765,N_14199,N_14417);
and U15766 (N_15766,N_14091,N_14685);
and U15767 (N_15767,N_14274,N_14579);
nand U15768 (N_15768,N_14929,N_14425);
and U15769 (N_15769,N_14834,N_14501);
nor U15770 (N_15770,N_14168,N_14689);
and U15771 (N_15771,N_14000,N_14333);
nor U15772 (N_15772,N_13850,N_14272);
and U15773 (N_15773,N_13836,N_14211);
and U15774 (N_15774,N_13785,N_14838);
or U15775 (N_15775,N_14575,N_14185);
nand U15776 (N_15776,N_14557,N_13886);
nor U15777 (N_15777,N_14366,N_13977);
xor U15778 (N_15778,N_14317,N_14127);
nor U15779 (N_15779,N_13808,N_14780);
or U15780 (N_15780,N_14513,N_14868);
nand U15781 (N_15781,N_14619,N_14756);
or U15782 (N_15782,N_14033,N_14216);
nor U15783 (N_15783,N_14627,N_14783);
nand U15784 (N_15784,N_14853,N_14199);
nor U15785 (N_15785,N_14804,N_14915);
nor U15786 (N_15786,N_14804,N_13938);
or U15787 (N_15787,N_14632,N_14085);
and U15788 (N_15788,N_13834,N_14246);
xnor U15789 (N_15789,N_13815,N_14335);
and U15790 (N_15790,N_13898,N_13872);
xnor U15791 (N_15791,N_14264,N_14082);
nor U15792 (N_15792,N_14671,N_14454);
nand U15793 (N_15793,N_14830,N_14556);
nand U15794 (N_15794,N_14342,N_14097);
or U15795 (N_15795,N_14642,N_14288);
nor U15796 (N_15796,N_14566,N_14190);
or U15797 (N_15797,N_14064,N_14947);
or U15798 (N_15798,N_14330,N_13880);
or U15799 (N_15799,N_14161,N_14197);
nand U15800 (N_15800,N_14879,N_14957);
nand U15801 (N_15801,N_14711,N_14020);
or U15802 (N_15802,N_14184,N_14475);
nor U15803 (N_15803,N_13999,N_14496);
xor U15804 (N_15804,N_14443,N_14317);
nor U15805 (N_15805,N_14756,N_13889);
nand U15806 (N_15806,N_14820,N_13948);
nand U15807 (N_15807,N_14044,N_14275);
and U15808 (N_15808,N_13890,N_14032);
nor U15809 (N_15809,N_14181,N_14202);
nor U15810 (N_15810,N_14217,N_14669);
and U15811 (N_15811,N_14421,N_14968);
nor U15812 (N_15812,N_14650,N_14874);
or U15813 (N_15813,N_14283,N_14385);
nand U15814 (N_15814,N_14075,N_13804);
or U15815 (N_15815,N_13810,N_14078);
nand U15816 (N_15816,N_13811,N_14123);
or U15817 (N_15817,N_13929,N_14011);
or U15818 (N_15818,N_14046,N_14509);
nand U15819 (N_15819,N_14589,N_14223);
and U15820 (N_15820,N_13890,N_14976);
nor U15821 (N_15821,N_14808,N_14873);
xnor U15822 (N_15822,N_14486,N_14290);
or U15823 (N_15823,N_14435,N_14695);
nor U15824 (N_15824,N_14835,N_14769);
nand U15825 (N_15825,N_14804,N_14875);
nor U15826 (N_15826,N_13913,N_14145);
nor U15827 (N_15827,N_14235,N_13800);
and U15828 (N_15828,N_14903,N_14957);
nand U15829 (N_15829,N_14335,N_13855);
xor U15830 (N_15830,N_14762,N_13804);
xor U15831 (N_15831,N_14383,N_14734);
nand U15832 (N_15832,N_14117,N_14503);
nor U15833 (N_15833,N_14829,N_13762);
nand U15834 (N_15834,N_14412,N_14204);
nor U15835 (N_15835,N_14936,N_14067);
nor U15836 (N_15836,N_14402,N_14325);
or U15837 (N_15837,N_14721,N_14345);
nor U15838 (N_15838,N_14378,N_13995);
and U15839 (N_15839,N_14532,N_13963);
xor U15840 (N_15840,N_14383,N_13947);
xnor U15841 (N_15841,N_14923,N_13988);
and U15842 (N_15842,N_14154,N_14577);
or U15843 (N_15843,N_14013,N_14346);
nor U15844 (N_15844,N_13919,N_14143);
xnor U15845 (N_15845,N_13930,N_14490);
nor U15846 (N_15846,N_14103,N_14362);
xnor U15847 (N_15847,N_14681,N_13758);
xor U15848 (N_15848,N_14589,N_13837);
or U15849 (N_15849,N_14010,N_14355);
or U15850 (N_15850,N_14732,N_14615);
or U15851 (N_15851,N_14152,N_14404);
or U15852 (N_15852,N_14845,N_14338);
nor U15853 (N_15853,N_14796,N_14400);
nand U15854 (N_15854,N_14337,N_14657);
or U15855 (N_15855,N_13929,N_14759);
or U15856 (N_15856,N_14667,N_14072);
and U15857 (N_15857,N_14494,N_14598);
xnor U15858 (N_15858,N_14197,N_14633);
or U15859 (N_15859,N_14195,N_14245);
or U15860 (N_15860,N_14687,N_13775);
or U15861 (N_15861,N_14285,N_14307);
or U15862 (N_15862,N_14310,N_14182);
and U15863 (N_15863,N_14655,N_13822);
xor U15864 (N_15864,N_14203,N_13990);
or U15865 (N_15865,N_14587,N_14172);
or U15866 (N_15866,N_13817,N_13754);
nand U15867 (N_15867,N_14578,N_14595);
or U15868 (N_15868,N_14408,N_14362);
nor U15869 (N_15869,N_14468,N_14152);
nand U15870 (N_15870,N_14040,N_14595);
or U15871 (N_15871,N_14302,N_14565);
or U15872 (N_15872,N_14190,N_14718);
nand U15873 (N_15873,N_14666,N_14047);
xor U15874 (N_15874,N_14295,N_14197);
xor U15875 (N_15875,N_14040,N_14232);
xnor U15876 (N_15876,N_14942,N_14723);
nor U15877 (N_15877,N_14182,N_13778);
xor U15878 (N_15878,N_14160,N_14954);
or U15879 (N_15879,N_14345,N_14860);
and U15880 (N_15880,N_14336,N_13941);
nor U15881 (N_15881,N_14291,N_14796);
nor U15882 (N_15882,N_13789,N_14300);
nand U15883 (N_15883,N_14251,N_13881);
xor U15884 (N_15884,N_14984,N_13979);
xor U15885 (N_15885,N_14780,N_14831);
and U15886 (N_15886,N_14130,N_14030);
or U15887 (N_15887,N_13906,N_14964);
nand U15888 (N_15888,N_13957,N_14572);
nand U15889 (N_15889,N_13813,N_13953);
xor U15890 (N_15890,N_14007,N_14334);
nand U15891 (N_15891,N_14022,N_14480);
nor U15892 (N_15892,N_14524,N_14331);
nor U15893 (N_15893,N_14451,N_14764);
or U15894 (N_15894,N_14742,N_13942);
or U15895 (N_15895,N_14975,N_14742);
nand U15896 (N_15896,N_14350,N_14732);
xor U15897 (N_15897,N_14499,N_14706);
and U15898 (N_15898,N_14383,N_14633);
nor U15899 (N_15899,N_14698,N_14304);
xor U15900 (N_15900,N_14617,N_14058);
nor U15901 (N_15901,N_14739,N_14866);
nor U15902 (N_15902,N_14746,N_14467);
and U15903 (N_15903,N_14154,N_13923);
or U15904 (N_15904,N_14728,N_14800);
and U15905 (N_15905,N_14864,N_13969);
nor U15906 (N_15906,N_14676,N_14700);
and U15907 (N_15907,N_14093,N_14786);
and U15908 (N_15908,N_13969,N_14761);
nand U15909 (N_15909,N_14437,N_13995);
or U15910 (N_15910,N_14767,N_13909);
nor U15911 (N_15911,N_14959,N_14467);
xnor U15912 (N_15912,N_13819,N_13846);
nor U15913 (N_15913,N_14669,N_14642);
or U15914 (N_15914,N_14998,N_14243);
and U15915 (N_15915,N_14010,N_14873);
or U15916 (N_15916,N_14108,N_13933);
or U15917 (N_15917,N_14788,N_14469);
nand U15918 (N_15918,N_13975,N_13922);
and U15919 (N_15919,N_14384,N_14569);
xor U15920 (N_15920,N_14852,N_14239);
nand U15921 (N_15921,N_14055,N_14612);
xnor U15922 (N_15922,N_14906,N_14946);
and U15923 (N_15923,N_13811,N_14289);
and U15924 (N_15924,N_14697,N_13856);
xnor U15925 (N_15925,N_14008,N_14566);
and U15926 (N_15926,N_14764,N_13973);
or U15927 (N_15927,N_14402,N_14734);
xor U15928 (N_15928,N_14856,N_14461);
or U15929 (N_15929,N_14179,N_13850);
xor U15930 (N_15930,N_13842,N_13914);
and U15931 (N_15931,N_14411,N_13950);
and U15932 (N_15932,N_14998,N_13885);
xnor U15933 (N_15933,N_14955,N_14536);
xor U15934 (N_15934,N_13983,N_14749);
xnor U15935 (N_15935,N_14050,N_14186);
nor U15936 (N_15936,N_14945,N_14141);
nand U15937 (N_15937,N_14009,N_14268);
nand U15938 (N_15938,N_14516,N_14016);
and U15939 (N_15939,N_14157,N_14950);
and U15940 (N_15940,N_14477,N_14652);
and U15941 (N_15941,N_14746,N_14405);
nand U15942 (N_15942,N_13925,N_14485);
xnor U15943 (N_15943,N_14178,N_14203);
or U15944 (N_15944,N_14033,N_14970);
nor U15945 (N_15945,N_14971,N_14388);
nand U15946 (N_15946,N_14917,N_14230);
xnor U15947 (N_15947,N_14964,N_14483);
nand U15948 (N_15948,N_14412,N_14239);
or U15949 (N_15949,N_14871,N_14354);
and U15950 (N_15950,N_14963,N_14368);
nor U15951 (N_15951,N_14650,N_14256);
and U15952 (N_15952,N_14553,N_14373);
xnor U15953 (N_15953,N_14322,N_14645);
nor U15954 (N_15954,N_14553,N_14579);
and U15955 (N_15955,N_13947,N_14043);
or U15956 (N_15956,N_14188,N_13872);
or U15957 (N_15957,N_14895,N_14818);
or U15958 (N_15958,N_14144,N_14719);
nand U15959 (N_15959,N_13992,N_14381);
xor U15960 (N_15960,N_14952,N_14673);
nand U15961 (N_15961,N_14426,N_14968);
nor U15962 (N_15962,N_14750,N_14882);
or U15963 (N_15963,N_13995,N_14761);
nand U15964 (N_15964,N_13769,N_14741);
xor U15965 (N_15965,N_13784,N_14962);
and U15966 (N_15966,N_13927,N_13829);
xor U15967 (N_15967,N_14907,N_14557);
nand U15968 (N_15968,N_13953,N_14389);
xor U15969 (N_15969,N_14369,N_14074);
nor U15970 (N_15970,N_13769,N_13914);
and U15971 (N_15971,N_14895,N_14351);
nand U15972 (N_15972,N_14486,N_14007);
nand U15973 (N_15973,N_14912,N_14116);
nor U15974 (N_15974,N_14577,N_14581);
nor U15975 (N_15975,N_14084,N_13857);
or U15976 (N_15976,N_14428,N_14505);
nor U15977 (N_15977,N_14261,N_14716);
nor U15978 (N_15978,N_14167,N_14103);
xnor U15979 (N_15979,N_13883,N_13867);
nand U15980 (N_15980,N_14477,N_13943);
and U15981 (N_15981,N_14855,N_13926);
and U15982 (N_15982,N_14921,N_14952);
xnor U15983 (N_15983,N_14303,N_14672);
nor U15984 (N_15984,N_14726,N_14192);
and U15985 (N_15985,N_14946,N_14032);
and U15986 (N_15986,N_13965,N_14749);
xnor U15987 (N_15987,N_14972,N_14463);
xor U15988 (N_15988,N_14130,N_14300);
xor U15989 (N_15989,N_13880,N_14746);
nor U15990 (N_15990,N_14175,N_14720);
and U15991 (N_15991,N_14838,N_14167);
and U15992 (N_15992,N_13937,N_14297);
and U15993 (N_15993,N_14215,N_14150);
and U15994 (N_15994,N_14274,N_14183);
nand U15995 (N_15995,N_13919,N_14665);
or U15996 (N_15996,N_14208,N_14821);
xor U15997 (N_15997,N_14228,N_14232);
xnor U15998 (N_15998,N_14418,N_14108);
and U15999 (N_15999,N_13843,N_14456);
xnor U16000 (N_16000,N_14999,N_14712);
nor U16001 (N_16001,N_14086,N_14203);
xor U16002 (N_16002,N_14663,N_14173);
and U16003 (N_16003,N_14154,N_13952);
xnor U16004 (N_16004,N_13897,N_14061);
and U16005 (N_16005,N_14823,N_14134);
or U16006 (N_16006,N_13977,N_14152);
or U16007 (N_16007,N_14548,N_14402);
and U16008 (N_16008,N_14730,N_14016);
and U16009 (N_16009,N_14871,N_14386);
xnor U16010 (N_16010,N_13984,N_14717);
or U16011 (N_16011,N_14015,N_14387);
xor U16012 (N_16012,N_14184,N_14103);
nor U16013 (N_16013,N_14065,N_14951);
or U16014 (N_16014,N_14249,N_14921);
and U16015 (N_16015,N_14972,N_14199);
nand U16016 (N_16016,N_13874,N_13982);
nand U16017 (N_16017,N_14382,N_14442);
xnor U16018 (N_16018,N_13754,N_14776);
nor U16019 (N_16019,N_14717,N_14008);
or U16020 (N_16020,N_14964,N_14566);
and U16021 (N_16021,N_14710,N_14361);
or U16022 (N_16022,N_13787,N_14237);
nor U16023 (N_16023,N_14292,N_14043);
nand U16024 (N_16024,N_13809,N_14849);
or U16025 (N_16025,N_14482,N_14475);
or U16026 (N_16026,N_14889,N_14617);
and U16027 (N_16027,N_14171,N_14490);
xnor U16028 (N_16028,N_14424,N_14145);
nand U16029 (N_16029,N_13874,N_14733);
nand U16030 (N_16030,N_14914,N_14890);
nand U16031 (N_16031,N_14584,N_14116);
xnor U16032 (N_16032,N_14453,N_14100);
nand U16033 (N_16033,N_14262,N_14795);
and U16034 (N_16034,N_14265,N_14070);
and U16035 (N_16035,N_14055,N_14508);
nor U16036 (N_16036,N_14408,N_13900);
nand U16037 (N_16037,N_14551,N_14415);
nand U16038 (N_16038,N_14598,N_14895);
or U16039 (N_16039,N_14756,N_14549);
and U16040 (N_16040,N_14957,N_14895);
and U16041 (N_16041,N_14563,N_14951);
and U16042 (N_16042,N_13781,N_14477);
xnor U16043 (N_16043,N_14591,N_14411);
nand U16044 (N_16044,N_14564,N_14788);
and U16045 (N_16045,N_14871,N_14857);
nor U16046 (N_16046,N_14337,N_13798);
and U16047 (N_16047,N_13991,N_14919);
xor U16048 (N_16048,N_14721,N_13937);
nand U16049 (N_16049,N_14650,N_14186);
nand U16050 (N_16050,N_14538,N_14242);
or U16051 (N_16051,N_14840,N_14383);
and U16052 (N_16052,N_14696,N_14898);
or U16053 (N_16053,N_14029,N_14605);
xnor U16054 (N_16054,N_14868,N_14017);
nand U16055 (N_16055,N_14566,N_14020);
nor U16056 (N_16056,N_14014,N_14870);
and U16057 (N_16057,N_14010,N_14490);
xor U16058 (N_16058,N_14305,N_14972);
or U16059 (N_16059,N_14039,N_14351);
nand U16060 (N_16060,N_14505,N_14427);
nor U16061 (N_16061,N_13997,N_14917);
or U16062 (N_16062,N_14766,N_14888);
xor U16063 (N_16063,N_14460,N_14641);
and U16064 (N_16064,N_14489,N_14081);
and U16065 (N_16065,N_14750,N_14260);
and U16066 (N_16066,N_13907,N_14412);
nand U16067 (N_16067,N_14947,N_14519);
nand U16068 (N_16068,N_14880,N_14102);
nand U16069 (N_16069,N_13942,N_14118);
nor U16070 (N_16070,N_14499,N_14048);
xnor U16071 (N_16071,N_14873,N_14697);
nand U16072 (N_16072,N_14824,N_14614);
nor U16073 (N_16073,N_14861,N_14851);
or U16074 (N_16074,N_14691,N_14899);
or U16075 (N_16075,N_14125,N_14717);
or U16076 (N_16076,N_14480,N_14544);
nor U16077 (N_16077,N_14340,N_14179);
nor U16078 (N_16078,N_14675,N_13891);
xor U16079 (N_16079,N_14256,N_14857);
or U16080 (N_16080,N_14652,N_14988);
and U16081 (N_16081,N_14853,N_14922);
nand U16082 (N_16082,N_14405,N_13992);
nand U16083 (N_16083,N_14903,N_14222);
or U16084 (N_16084,N_14596,N_14958);
and U16085 (N_16085,N_13941,N_14955);
and U16086 (N_16086,N_14861,N_14748);
nand U16087 (N_16087,N_13988,N_14961);
xor U16088 (N_16088,N_14818,N_14391);
xor U16089 (N_16089,N_14188,N_14861);
xor U16090 (N_16090,N_14895,N_14229);
nand U16091 (N_16091,N_14129,N_14621);
xor U16092 (N_16092,N_14194,N_14134);
nor U16093 (N_16093,N_13769,N_14486);
and U16094 (N_16094,N_14215,N_14345);
nand U16095 (N_16095,N_14073,N_14293);
nand U16096 (N_16096,N_14828,N_14578);
xor U16097 (N_16097,N_14882,N_14560);
or U16098 (N_16098,N_14274,N_14154);
nor U16099 (N_16099,N_14682,N_14783);
nor U16100 (N_16100,N_13843,N_13869);
nor U16101 (N_16101,N_14156,N_13812);
or U16102 (N_16102,N_14615,N_14571);
xor U16103 (N_16103,N_14523,N_13871);
or U16104 (N_16104,N_13866,N_14352);
xnor U16105 (N_16105,N_14734,N_14455);
nor U16106 (N_16106,N_14359,N_14144);
nor U16107 (N_16107,N_14587,N_14839);
xnor U16108 (N_16108,N_14548,N_14661);
nand U16109 (N_16109,N_14063,N_14520);
nor U16110 (N_16110,N_14298,N_13946);
xnor U16111 (N_16111,N_14929,N_13838);
nor U16112 (N_16112,N_14940,N_13985);
or U16113 (N_16113,N_14255,N_14477);
nor U16114 (N_16114,N_14204,N_14857);
or U16115 (N_16115,N_14409,N_14404);
or U16116 (N_16116,N_14552,N_14884);
nor U16117 (N_16117,N_14942,N_13988);
xor U16118 (N_16118,N_14632,N_14507);
and U16119 (N_16119,N_13933,N_13815);
and U16120 (N_16120,N_14157,N_14265);
or U16121 (N_16121,N_14404,N_14244);
and U16122 (N_16122,N_14341,N_14337);
nand U16123 (N_16123,N_14922,N_14331);
nor U16124 (N_16124,N_13773,N_13947);
xor U16125 (N_16125,N_14018,N_14427);
xor U16126 (N_16126,N_13882,N_14584);
nor U16127 (N_16127,N_14948,N_13839);
nand U16128 (N_16128,N_14432,N_13892);
nand U16129 (N_16129,N_14299,N_14623);
and U16130 (N_16130,N_13762,N_14888);
nor U16131 (N_16131,N_13903,N_14641);
xnor U16132 (N_16132,N_14372,N_14920);
nand U16133 (N_16133,N_14749,N_14805);
and U16134 (N_16134,N_13932,N_14229);
or U16135 (N_16135,N_14771,N_14789);
nor U16136 (N_16136,N_14464,N_14869);
and U16137 (N_16137,N_14857,N_14702);
or U16138 (N_16138,N_14984,N_14547);
xor U16139 (N_16139,N_14088,N_14269);
and U16140 (N_16140,N_14466,N_13819);
xor U16141 (N_16141,N_14842,N_13886);
nand U16142 (N_16142,N_14858,N_14020);
or U16143 (N_16143,N_14780,N_14413);
and U16144 (N_16144,N_13861,N_14606);
nand U16145 (N_16145,N_14730,N_14593);
nor U16146 (N_16146,N_14634,N_14156);
xnor U16147 (N_16147,N_14018,N_14045);
nor U16148 (N_16148,N_14295,N_14344);
xnor U16149 (N_16149,N_14677,N_14365);
nor U16150 (N_16150,N_14904,N_14053);
xnor U16151 (N_16151,N_14899,N_13831);
and U16152 (N_16152,N_14278,N_14117);
xnor U16153 (N_16153,N_14596,N_14905);
xor U16154 (N_16154,N_14927,N_14089);
and U16155 (N_16155,N_14565,N_14445);
and U16156 (N_16156,N_14380,N_14935);
nand U16157 (N_16157,N_14153,N_14027);
or U16158 (N_16158,N_14805,N_14747);
xnor U16159 (N_16159,N_14085,N_14860);
or U16160 (N_16160,N_14806,N_14903);
and U16161 (N_16161,N_13921,N_14191);
nand U16162 (N_16162,N_13956,N_13939);
or U16163 (N_16163,N_14724,N_14187);
or U16164 (N_16164,N_14579,N_14077);
nor U16165 (N_16165,N_14731,N_14054);
nand U16166 (N_16166,N_14406,N_14314);
and U16167 (N_16167,N_14475,N_14376);
xnor U16168 (N_16168,N_14952,N_14223);
xnor U16169 (N_16169,N_14660,N_13872);
xnor U16170 (N_16170,N_14430,N_13866);
and U16171 (N_16171,N_14268,N_14995);
and U16172 (N_16172,N_14916,N_13993);
xor U16173 (N_16173,N_14752,N_13819);
nand U16174 (N_16174,N_14651,N_14305);
nand U16175 (N_16175,N_14186,N_14762);
xnor U16176 (N_16176,N_13778,N_14558);
nor U16177 (N_16177,N_14205,N_14112);
xnor U16178 (N_16178,N_14049,N_14477);
nor U16179 (N_16179,N_14351,N_14914);
xnor U16180 (N_16180,N_14567,N_14453);
xnor U16181 (N_16181,N_14232,N_14364);
and U16182 (N_16182,N_14603,N_14147);
xnor U16183 (N_16183,N_14955,N_14605);
and U16184 (N_16184,N_14631,N_13932);
nand U16185 (N_16185,N_14434,N_14278);
or U16186 (N_16186,N_13997,N_14085);
nand U16187 (N_16187,N_14882,N_14526);
or U16188 (N_16188,N_13915,N_14168);
and U16189 (N_16189,N_14871,N_14745);
xnor U16190 (N_16190,N_14369,N_14118);
nand U16191 (N_16191,N_14658,N_14718);
nor U16192 (N_16192,N_14181,N_14985);
nor U16193 (N_16193,N_14661,N_14832);
nor U16194 (N_16194,N_14462,N_14183);
nor U16195 (N_16195,N_14105,N_14015);
xnor U16196 (N_16196,N_14144,N_13825);
xnor U16197 (N_16197,N_14485,N_13815);
and U16198 (N_16198,N_14276,N_14757);
or U16199 (N_16199,N_13961,N_13955);
nand U16200 (N_16200,N_13906,N_14507);
nor U16201 (N_16201,N_14342,N_14563);
and U16202 (N_16202,N_14872,N_14376);
nand U16203 (N_16203,N_14284,N_13824);
nor U16204 (N_16204,N_13919,N_14193);
nand U16205 (N_16205,N_13906,N_14135);
and U16206 (N_16206,N_14742,N_14659);
nand U16207 (N_16207,N_14152,N_14155);
xnor U16208 (N_16208,N_14642,N_13765);
and U16209 (N_16209,N_14833,N_14470);
and U16210 (N_16210,N_14849,N_14264);
and U16211 (N_16211,N_13790,N_13771);
or U16212 (N_16212,N_14762,N_14576);
nor U16213 (N_16213,N_14913,N_14771);
xnor U16214 (N_16214,N_14392,N_14880);
nor U16215 (N_16215,N_14858,N_14117);
and U16216 (N_16216,N_14708,N_14906);
and U16217 (N_16217,N_13871,N_14279);
xnor U16218 (N_16218,N_13993,N_14311);
nor U16219 (N_16219,N_14804,N_14995);
or U16220 (N_16220,N_14099,N_14358);
or U16221 (N_16221,N_13889,N_14819);
xnor U16222 (N_16222,N_14323,N_14607);
nor U16223 (N_16223,N_14642,N_13949);
xnor U16224 (N_16224,N_14569,N_14009);
nand U16225 (N_16225,N_13890,N_14764);
nor U16226 (N_16226,N_14460,N_14585);
nand U16227 (N_16227,N_13985,N_14256);
and U16228 (N_16228,N_14573,N_14756);
or U16229 (N_16229,N_14817,N_14495);
nor U16230 (N_16230,N_13756,N_14540);
xor U16231 (N_16231,N_14648,N_14368);
and U16232 (N_16232,N_14862,N_14864);
nor U16233 (N_16233,N_14119,N_14477);
xor U16234 (N_16234,N_14533,N_13805);
nand U16235 (N_16235,N_14378,N_14845);
xor U16236 (N_16236,N_14169,N_14149);
and U16237 (N_16237,N_14506,N_14046);
nor U16238 (N_16238,N_13870,N_13816);
and U16239 (N_16239,N_13853,N_14140);
or U16240 (N_16240,N_14248,N_14483);
nand U16241 (N_16241,N_14178,N_14657);
and U16242 (N_16242,N_14046,N_13810);
xor U16243 (N_16243,N_14868,N_14719);
xor U16244 (N_16244,N_14989,N_14739);
xor U16245 (N_16245,N_14839,N_14044);
nand U16246 (N_16246,N_13809,N_14891);
nor U16247 (N_16247,N_13798,N_14721);
nand U16248 (N_16248,N_14553,N_14802);
nand U16249 (N_16249,N_14082,N_14574);
xnor U16250 (N_16250,N_15775,N_15933);
nand U16251 (N_16251,N_16237,N_16115);
nand U16252 (N_16252,N_15592,N_15413);
and U16253 (N_16253,N_15444,N_15229);
nor U16254 (N_16254,N_15453,N_15499);
xor U16255 (N_16255,N_15323,N_15707);
and U16256 (N_16256,N_15184,N_15642);
nand U16257 (N_16257,N_16002,N_15722);
nor U16258 (N_16258,N_15944,N_16154);
nand U16259 (N_16259,N_15825,N_15056);
and U16260 (N_16260,N_15377,N_16119);
nor U16261 (N_16261,N_15454,N_16001);
nor U16262 (N_16262,N_15689,N_15862);
or U16263 (N_16263,N_15107,N_16139);
xnor U16264 (N_16264,N_15298,N_15653);
nand U16265 (N_16265,N_16005,N_16182);
and U16266 (N_16266,N_16113,N_16076);
nand U16267 (N_16267,N_15017,N_15828);
and U16268 (N_16268,N_16206,N_15824);
xor U16269 (N_16269,N_15437,N_16068);
nor U16270 (N_16270,N_15053,N_15030);
or U16271 (N_16271,N_15640,N_15218);
nand U16272 (N_16272,N_15540,N_15532);
nand U16273 (N_16273,N_15975,N_15335);
xnor U16274 (N_16274,N_15637,N_15925);
nand U16275 (N_16275,N_16046,N_15246);
or U16276 (N_16276,N_15957,N_15114);
nand U16277 (N_16277,N_16123,N_15522);
nand U16278 (N_16278,N_15514,N_15461);
and U16279 (N_16279,N_15368,N_15013);
or U16280 (N_16280,N_15567,N_15068);
nor U16281 (N_16281,N_15673,N_16210);
xor U16282 (N_16282,N_15595,N_15216);
nor U16283 (N_16283,N_15877,N_16169);
nor U16284 (N_16284,N_15575,N_15728);
and U16285 (N_16285,N_15544,N_15482);
nor U16286 (N_16286,N_15835,N_15027);
and U16287 (N_16287,N_15442,N_15733);
nor U16288 (N_16288,N_16231,N_15194);
nand U16289 (N_16289,N_16177,N_15886);
nand U16290 (N_16290,N_15913,N_15311);
or U16291 (N_16291,N_15993,N_15654);
nor U16292 (N_16292,N_15249,N_15100);
and U16293 (N_16293,N_16197,N_15672);
nor U16294 (N_16294,N_15005,N_15766);
or U16295 (N_16295,N_15716,N_15521);
xor U16296 (N_16296,N_15570,N_15702);
xnor U16297 (N_16297,N_15346,N_15996);
nand U16298 (N_16298,N_15945,N_15140);
and U16299 (N_16299,N_15968,N_15051);
xnor U16300 (N_16300,N_15032,N_15602);
nand U16301 (N_16301,N_15598,N_15739);
nand U16302 (N_16302,N_15034,N_15579);
nor U16303 (N_16303,N_15819,N_15020);
nand U16304 (N_16304,N_15538,N_16134);
or U16305 (N_16305,N_15650,N_15666);
nand U16306 (N_16306,N_15907,N_15258);
nor U16307 (N_16307,N_15900,N_15665);
xnor U16308 (N_16308,N_16081,N_15037);
or U16309 (N_16309,N_15080,N_15787);
and U16310 (N_16310,N_15755,N_15314);
xor U16311 (N_16311,N_15790,N_15822);
nor U16312 (N_16312,N_15199,N_15067);
xor U16313 (N_16313,N_15102,N_15447);
or U16314 (N_16314,N_15742,N_15711);
nor U16315 (N_16315,N_15542,N_16207);
and U16316 (N_16316,N_15125,N_15606);
or U16317 (N_16317,N_16017,N_15240);
xor U16318 (N_16318,N_15856,N_15322);
xor U16319 (N_16319,N_15338,N_15276);
or U16320 (N_16320,N_15266,N_15631);
xnor U16321 (N_16321,N_15554,N_16122);
nand U16322 (N_16322,N_15381,N_16215);
nand U16323 (N_16323,N_16128,N_15093);
nor U16324 (N_16324,N_15360,N_15457);
or U16325 (N_16325,N_15046,N_16241);
nand U16326 (N_16326,N_15195,N_15963);
xor U16327 (N_16327,N_15226,N_15717);
nor U16328 (N_16328,N_15632,N_15127);
nand U16329 (N_16329,N_15513,N_15006);
xor U16330 (N_16330,N_15679,N_15841);
nor U16331 (N_16331,N_15915,N_15677);
or U16332 (N_16332,N_16175,N_15830);
xnor U16333 (N_16333,N_15430,N_15799);
nor U16334 (N_16334,N_15315,N_16082);
and U16335 (N_16335,N_15112,N_16011);
xor U16336 (N_16336,N_15419,N_15057);
or U16337 (N_16337,N_15337,N_16194);
xor U16338 (N_16338,N_15780,N_15872);
or U16339 (N_16339,N_15487,N_16141);
nor U16340 (N_16340,N_15713,N_15424);
nand U16341 (N_16341,N_16042,N_15065);
nor U16342 (N_16342,N_15596,N_15254);
xor U16343 (N_16343,N_16060,N_15397);
nor U16344 (N_16344,N_15069,N_15452);
and U16345 (N_16345,N_15366,N_15611);
and U16346 (N_16346,N_15163,N_15206);
or U16347 (N_16347,N_15991,N_15591);
or U16348 (N_16348,N_15519,N_15279);
nor U16349 (N_16349,N_15155,N_16008);
nand U16350 (N_16350,N_15232,N_15467);
nand U16351 (N_16351,N_15643,N_16025);
or U16352 (N_16352,N_15543,N_16108);
and U16353 (N_16353,N_15325,N_15211);
or U16354 (N_16354,N_15283,N_15883);
nand U16355 (N_16355,N_15089,N_15864);
xnor U16356 (N_16356,N_15443,N_15831);
nand U16357 (N_16357,N_15001,N_15026);
or U16358 (N_16358,N_15261,N_15025);
xor U16359 (N_16359,N_16245,N_15850);
nor U16360 (N_16360,N_15160,N_15428);
nor U16361 (N_16361,N_15663,N_15729);
and U16362 (N_16362,N_15779,N_16171);
or U16363 (N_16363,N_16069,N_15772);
and U16364 (N_16364,N_15192,N_15369);
nand U16365 (N_16365,N_15358,N_16190);
nand U16366 (N_16366,N_16054,N_16013);
or U16367 (N_16367,N_15556,N_15892);
nand U16368 (N_16368,N_15130,N_15984);
and U16369 (N_16369,N_15152,N_15588);
nand U16370 (N_16370,N_15881,N_15549);
xnor U16371 (N_16371,N_15282,N_15297);
nand U16372 (N_16372,N_15584,N_15559);
nand U16373 (N_16373,N_15607,N_15148);
nand U16374 (N_16374,N_15463,N_16044);
nand U16375 (N_16375,N_15275,N_16118);
xnor U16376 (N_16376,N_15170,N_16070);
xnor U16377 (N_16377,N_15762,N_15939);
xor U16378 (N_16378,N_15081,N_15349);
nor U16379 (N_16379,N_15541,N_15614);
nor U16380 (N_16380,N_15660,N_15820);
nand U16381 (N_16381,N_15574,N_15210);
or U16382 (N_16382,N_15484,N_15867);
or U16383 (N_16383,N_15878,N_15274);
nand U16384 (N_16384,N_15052,N_15674);
nor U16385 (N_16385,N_15146,N_16238);
and U16386 (N_16386,N_16105,N_15106);
xor U16387 (N_16387,N_15931,N_15497);
xnor U16388 (N_16388,N_15569,N_15238);
xor U16389 (N_16389,N_16212,N_15151);
or U16390 (N_16390,N_15235,N_15562);
xor U16391 (N_16391,N_15885,N_15694);
nand U16392 (N_16392,N_15414,N_15408);
nor U16393 (N_16393,N_15789,N_16133);
or U16394 (N_16394,N_15998,N_15410);
nand U16395 (N_16395,N_16196,N_16145);
xnor U16396 (N_16396,N_15664,N_15609);
and U16397 (N_16397,N_15122,N_15060);
xor U16398 (N_16398,N_15743,N_15581);
xnor U16399 (N_16399,N_15669,N_15491);
or U16400 (N_16400,N_15839,N_15851);
or U16401 (N_16401,N_15383,N_15488);
and U16402 (N_16402,N_15055,N_15372);
xnor U16403 (N_16403,N_15919,N_15402);
nor U16404 (N_16404,N_15597,N_15623);
nand U16405 (N_16405,N_15604,N_15019);
or U16406 (N_16406,N_16028,N_15866);
and U16407 (N_16407,N_15794,N_15593);
nor U16408 (N_16408,N_16007,N_15128);
or U16409 (N_16409,N_16092,N_15200);
and U16410 (N_16410,N_15807,N_15000);
nand U16411 (N_16411,N_16151,N_15399);
and U16412 (N_16412,N_15712,N_15531);
nor U16413 (N_16413,N_16100,N_15373);
xnor U16414 (N_16414,N_15259,N_15244);
nor U16415 (N_16415,N_15063,N_15546);
and U16416 (N_16416,N_15667,N_15126);
and U16417 (N_16417,N_16243,N_15262);
xor U16418 (N_16418,N_15264,N_15662);
nand U16419 (N_16419,N_15979,N_16120);
nor U16420 (N_16420,N_15021,N_15117);
and U16421 (N_16421,N_16148,N_15064);
xnor U16422 (N_16422,N_15243,N_15684);
and U16423 (N_16423,N_16058,N_15459);
and U16424 (N_16424,N_16107,N_15857);
xor U16425 (N_16425,N_15012,N_15110);
nand U16426 (N_16426,N_15781,N_15028);
nor U16427 (N_16427,N_15409,N_15073);
nand U16428 (N_16428,N_15004,N_15858);
and U16429 (N_16429,N_16091,N_15967);
or U16430 (N_16430,N_15201,N_15247);
nor U16431 (N_16431,N_15964,N_15942);
xnor U16432 (N_16432,N_16063,N_15286);
xor U16433 (N_16433,N_16126,N_15087);
and U16434 (N_16434,N_15329,N_15500);
and U16435 (N_16435,N_15084,N_15086);
or U16436 (N_16436,N_15995,N_15096);
and U16437 (N_16437,N_15113,N_16136);
and U16438 (N_16438,N_15888,N_15882);
nand U16439 (N_16439,N_15633,N_15761);
xnor U16440 (N_16440,N_15507,N_15853);
and U16441 (N_16441,N_15134,N_15950);
and U16442 (N_16442,N_16235,N_15977);
or U16443 (N_16443,N_15193,N_15121);
nor U16444 (N_16444,N_15111,N_15432);
or U16445 (N_16445,N_15852,N_15250);
nand U16446 (N_16446,N_15328,N_15986);
or U16447 (N_16447,N_15267,N_15388);
xor U16448 (N_16448,N_16110,N_15989);
nor U16449 (N_16449,N_15608,N_16036);
or U16450 (N_16450,N_15357,N_15670);
or U16451 (N_16451,N_15908,N_16072);
nor U16452 (N_16452,N_15417,N_15924);
or U16453 (N_16453,N_15342,N_15198);
nand U16454 (N_16454,N_16249,N_16168);
or U16455 (N_16455,N_15777,N_15699);
nor U16456 (N_16456,N_16078,N_15203);
nand U16457 (N_16457,N_16211,N_15760);
nand U16458 (N_16458,N_15874,N_16247);
or U16459 (N_16459,N_15813,N_15626);
and U16460 (N_16460,N_15320,N_15331);
or U16461 (N_16461,N_15010,N_16203);
nor U16462 (N_16462,N_15651,N_16221);
and U16463 (N_16463,N_16234,N_15680);
or U16464 (N_16464,N_15186,N_16097);
nand U16465 (N_16465,N_15044,N_15480);
xor U16466 (N_16466,N_15691,N_15868);
nor U16467 (N_16467,N_15610,N_15798);
or U16468 (N_16468,N_16156,N_15404);
or U16469 (N_16469,N_16112,N_15510);
nand U16470 (N_16470,N_15758,N_15618);
or U16471 (N_16471,N_16102,N_15304);
or U16472 (N_16472,N_15759,N_15518);
xnor U16473 (N_16473,N_15854,N_15916);
nor U16474 (N_16474,N_15131,N_15038);
nor U16475 (N_16475,N_15587,N_15551);
and U16476 (N_16476,N_15740,N_15164);
and U16477 (N_16477,N_15054,N_16174);
and U16478 (N_16478,N_15829,N_16020);
nand U16479 (N_16479,N_15123,N_15720);
and U16480 (N_16480,N_16075,N_15230);
and U16481 (N_16481,N_16117,N_15464);
or U16482 (N_16482,N_15603,N_15774);
nand U16483 (N_16483,N_15710,N_15345);
or U16484 (N_16484,N_15517,N_15321);
or U16485 (N_16485,N_15451,N_15827);
nand U16486 (N_16486,N_15895,N_16019);
and U16487 (N_16487,N_16099,N_15108);
xnor U16488 (N_16488,N_15241,N_15936);
or U16489 (N_16489,N_15659,N_15171);
nor U16490 (N_16490,N_15031,N_15706);
xnor U16491 (N_16491,N_15990,N_15696);
or U16492 (N_16492,N_15429,N_16216);
or U16493 (N_16493,N_15217,N_15287);
nor U16494 (N_16494,N_16012,N_15771);
or U16495 (N_16495,N_15115,N_15622);
nand U16496 (N_16496,N_15179,N_16173);
nor U16497 (N_16497,N_16111,N_15586);
nor U16498 (N_16498,N_15747,N_15422);
nor U16499 (N_16499,N_15547,N_16181);
xor U16500 (N_16500,N_15745,N_16109);
or U16501 (N_16501,N_15700,N_15844);
nand U16502 (N_16502,N_15951,N_15132);
or U16503 (N_16503,N_15668,N_15492);
xnor U16504 (N_16504,N_15840,N_15553);
nor U16505 (N_16505,N_15135,N_15224);
nand U16506 (N_16506,N_16236,N_16202);
or U16507 (N_16507,N_15293,N_15292);
and U16508 (N_16508,N_16027,N_15571);
or U16509 (N_16509,N_15374,N_16233);
nand U16510 (N_16510,N_16204,N_15016);
or U16511 (N_16511,N_16057,N_15088);
nand U16512 (N_16512,N_15066,N_15784);
nand U16513 (N_16513,N_15426,N_15280);
or U16514 (N_16514,N_15578,N_16155);
and U16515 (N_16515,N_15601,N_15455);
and U16516 (N_16516,N_16159,N_15281);
nand U16517 (N_16517,N_15860,N_15434);
and U16518 (N_16518,N_15972,N_15450);
nand U16519 (N_16519,N_15528,N_15641);
and U16520 (N_16520,N_15182,N_15803);
nand U16521 (N_16521,N_15221,N_15589);
xor U16522 (N_16522,N_15736,N_15009);
or U16523 (N_16523,N_15548,N_15692);
or U16524 (N_16524,N_15277,N_15231);
or U16525 (N_16525,N_15726,N_15458);
or U16526 (N_16526,N_15786,N_15072);
xnor U16527 (N_16527,N_15384,N_15178);
nor U16528 (N_16528,N_15855,N_15278);
and U16529 (N_16529,N_15501,N_15912);
and U16530 (N_16530,N_15927,N_15634);
nand U16531 (N_16531,N_15048,N_16138);
or U16532 (N_16532,N_16003,N_15049);
nand U16533 (N_16533,N_15161,N_15062);
nor U16534 (N_16534,N_15169,N_15209);
xor U16535 (N_16535,N_15253,N_15156);
or U16536 (N_16536,N_15473,N_16022);
nand U16537 (N_16537,N_15564,N_15506);
or U16538 (N_16538,N_15023,N_16192);
nor U16539 (N_16539,N_15884,N_15658);
nor U16540 (N_16540,N_15339,N_16144);
xor U16541 (N_16541,N_15675,N_15953);
nand U16542 (N_16542,N_15425,N_16180);
nand U16543 (N_16543,N_16062,N_16176);
nor U16544 (N_16544,N_15616,N_15836);
xor U16545 (N_16545,N_15175,N_15185);
nor U16546 (N_16546,N_15272,N_15502);
xor U16547 (N_16547,N_16152,N_15050);
xnor U16548 (N_16548,N_16071,N_15316);
xnor U16549 (N_16549,N_15917,N_15365);
xor U16550 (N_16550,N_15572,N_15776);
and U16551 (N_16551,N_16161,N_15645);
nand U16552 (N_16552,N_15959,N_15291);
xor U16553 (N_16553,N_15600,N_15303);
nand U16554 (N_16554,N_15763,N_15937);
and U16555 (N_16555,N_15412,N_15225);
or U16556 (N_16556,N_16055,N_15002);
nor U16557 (N_16557,N_15811,N_15237);
or U16558 (N_16558,N_15465,N_15703);
and U16559 (N_16559,N_16074,N_16188);
and U16560 (N_16560,N_15719,N_16077);
nand U16561 (N_16561,N_15701,N_15697);
and U16562 (N_16562,N_16198,N_15804);
and U16563 (N_16563,N_15647,N_16096);
nor U16564 (N_16564,N_15767,N_15764);
xor U16565 (N_16565,N_15234,N_15566);
and U16566 (N_16566,N_15035,N_15753);
xnor U16567 (N_16567,N_15334,N_15678);
nand U16568 (N_16568,N_15797,N_15555);
nand U16569 (N_16569,N_15008,N_15635);
and U16570 (N_16570,N_16021,N_16140);
xnor U16571 (N_16571,N_15375,N_15406);
nor U16572 (N_16572,N_15573,N_15498);
and U16573 (N_16573,N_15838,N_15150);
and U16574 (N_16574,N_15439,N_15978);
nand U16575 (N_16575,N_15731,N_15071);
and U16576 (N_16576,N_15904,N_15153);
nor U16577 (N_16577,N_15735,N_15379);
nand U16578 (N_16578,N_16131,N_15214);
nand U16579 (N_16579,N_16164,N_15715);
nor U16580 (N_16580,N_15350,N_15393);
nor U16581 (N_16581,N_16093,N_15188);
xor U16582 (N_16582,N_16178,N_15421);
nor U16583 (N_16583,N_16172,N_15898);
nand U16584 (N_16584,N_15103,N_15343);
nor U16585 (N_16585,N_15585,N_15652);
or U16586 (N_16586,N_15557,N_15392);
nor U16587 (N_16587,N_15208,N_15920);
nand U16588 (N_16588,N_15983,N_15612);
or U16589 (N_16589,N_15795,N_15897);
xnor U16590 (N_16590,N_15928,N_15583);
xnor U16591 (N_16591,N_15173,N_15353);
or U16592 (N_16592,N_15997,N_15503);
nor U16593 (N_16593,N_15778,N_15594);
xor U16594 (N_16594,N_16226,N_15223);
nand U16595 (N_16595,N_16048,N_15638);
and U16596 (N_16596,N_16153,N_15400);
and U16597 (N_16597,N_15535,N_15961);
xnor U16598 (N_16598,N_16129,N_15903);
nor U16599 (N_16599,N_16040,N_15815);
and U16600 (N_16600,N_15168,N_15943);
xnor U16601 (N_16601,N_15284,N_15981);
nand U16602 (N_16602,N_15495,N_15523);
nor U16603 (N_16603,N_16009,N_15524);
nor U16604 (N_16604,N_15333,N_15980);
xnor U16605 (N_16605,N_15411,N_15215);
xnor U16606 (N_16606,N_15746,N_15085);
nor U16607 (N_16607,N_16085,N_15992);
xor U16608 (N_16608,N_15129,N_15976);
and U16609 (N_16609,N_16121,N_16000);
and U16610 (N_16610,N_15007,N_15141);
or U16611 (N_16611,N_15505,N_16183);
nand U16612 (N_16612,N_15630,N_15552);
nand U16613 (N_16613,N_15183,N_15773);
xnor U16614 (N_16614,N_15971,N_15751);
nor U16615 (N_16615,N_15625,N_15090);
nor U16616 (N_16616,N_15685,N_16014);
xor U16617 (N_16617,N_15441,N_15041);
and U16618 (N_16618,N_15833,N_16087);
nor U16619 (N_16619,N_15525,N_15661);
or U16620 (N_16620,N_16065,N_15639);
nand U16621 (N_16621,N_15157,N_15876);
and U16622 (N_16622,N_15987,N_15485);
nand U16623 (N_16623,N_15704,N_15288);
and U16624 (N_16624,N_15896,N_15880);
and U16625 (N_16625,N_15248,N_16049);
or U16626 (N_16626,N_15098,N_15905);
or U16627 (N_16627,N_15970,N_16061);
and U16628 (N_16628,N_15732,N_15255);
nor U16629 (N_16629,N_16227,N_15355);
nor U16630 (N_16630,N_15965,N_15265);
xor U16631 (N_16631,N_15627,N_15843);
xnor U16632 (N_16632,N_15520,N_15094);
and U16633 (N_16633,N_15871,N_16205);
and U16634 (N_16634,N_15910,N_15327);
nor U16635 (N_16635,N_15801,N_15344);
and U16636 (N_16636,N_16244,N_15015);
nand U16637 (N_16637,N_16162,N_15202);
xor U16638 (N_16638,N_15988,N_16127);
and U16639 (N_16639,N_15440,N_15516);
and U16640 (N_16640,N_16135,N_15101);
xor U16641 (N_16641,N_15370,N_15619);
xor U16642 (N_16642,N_15821,N_16130);
and U16643 (N_16643,N_15352,N_15033);
nand U16644 (N_16644,N_16089,N_16199);
nor U16645 (N_16645,N_15563,N_16064);
xnor U16646 (N_16646,N_16222,N_15723);
or U16647 (N_16647,N_15059,N_15083);
nor U16648 (N_16648,N_15361,N_15040);
or U16649 (N_16649,N_15312,N_15922);
nand U16650 (N_16650,N_16220,N_15909);
and U16651 (N_16651,N_16142,N_15222);
or U16652 (N_16652,N_15470,N_16189);
nand U16653 (N_16653,N_15351,N_15539);
nand U16654 (N_16654,N_15295,N_15362);
nand U16655 (N_16655,N_15166,N_15834);
nor U16656 (N_16656,N_15309,N_15962);
nor U16657 (N_16657,N_15236,N_15705);
nand U16658 (N_16658,N_16114,N_15865);
nor U16659 (N_16659,N_16137,N_15847);
nand U16660 (N_16660,N_15879,N_16094);
xor U16661 (N_16661,N_15737,N_15077);
nand U16662 (N_16662,N_15445,N_15239);
and U16663 (N_16663,N_15918,N_16026);
nand U16664 (N_16664,N_15769,N_15300);
and U16665 (N_16665,N_15873,N_16125);
or U16666 (N_16666,N_15802,N_15657);
nand U16667 (N_16667,N_15395,N_15471);
nor U16668 (N_16668,N_15104,N_15436);
xnor U16669 (N_16669,N_15788,N_15472);
nor U16670 (N_16670,N_15142,N_15527);
nor U16671 (N_16671,N_15940,N_15512);
and U16672 (N_16672,N_16149,N_15149);
nand U16673 (N_16673,N_15613,N_15816);
nor U16674 (N_16674,N_15263,N_15207);
and U16675 (N_16675,N_15205,N_15796);
nor U16676 (N_16676,N_15615,N_15386);
nor U16677 (N_16677,N_16179,N_16195);
xnor U16678 (N_16678,N_15730,N_15305);
or U16679 (N_16679,N_15427,N_16052);
or U16680 (N_16680,N_15823,N_15966);
or U16681 (N_16681,N_15415,N_15228);
nand U16682 (N_16682,N_16051,N_16147);
nand U16683 (N_16683,N_15143,N_15478);
xor U16684 (N_16684,N_15893,N_15158);
nor U16685 (N_16685,N_15911,N_15407);
and U16686 (N_16686,N_16059,N_15568);
and U16687 (N_16687,N_15646,N_15952);
xnor U16688 (N_16688,N_15744,N_15809);
xor U16689 (N_16689,N_15565,N_16223);
and U16690 (N_16690,N_15655,N_16037);
xor U16691 (N_16691,N_15105,N_15845);
or U16692 (N_16692,N_15245,N_15537);
nor U16693 (N_16693,N_15124,N_15621);
nand U16694 (N_16694,N_16230,N_16083);
nor U16695 (N_16695,N_15709,N_15926);
nor U16696 (N_16696,N_15174,N_15139);
xnor U16697 (N_16697,N_15268,N_15934);
or U16698 (N_16698,N_16080,N_16116);
or U16699 (N_16699,N_15133,N_15036);
and U16700 (N_16700,N_15466,N_15863);
nor U16701 (N_16701,N_15047,N_15545);
or U16702 (N_16702,N_15974,N_15826);
xor U16703 (N_16703,N_15354,N_16101);
and U16704 (N_16704,N_15011,N_15097);
xor U16705 (N_16705,N_15791,N_15190);
or U16706 (N_16706,N_15378,N_15681);
or U16707 (N_16707,N_15750,N_15800);
xor U16708 (N_16708,N_15902,N_15212);
xor U16709 (N_16709,N_16157,N_15116);
or U16710 (N_16710,N_15341,N_15561);
nor U16711 (N_16711,N_16219,N_16143);
or U16712 (N_16712,N_15376,N_16246);
or U16713 (N_16713,N_16186,N_15024);
nor U16714 (N_16714,N_15859,N_15782);
xnor U16715 (N_16715,N_16030,N_15754);
or U16716 (N_16716,N_15177,N_15363);
nand U16717 (N_16717,N_16038,N_16029);
nand U16718 (N_16718,N_15837,N_15748);
or U16719 (N_16719,N_15628,N_15162);
or U16720 (N_16720,N_15889,N_15165);
xor U16721 (N_16721,N_15418,N_15687);
or U16722 (N_16722,N_15960,N_15725);
or U16723 (N_16723,N_15887,N_16056);
or U16724 (N_16724,N_15332,N_16239);
nor U16725 (N_16725,N_16218,N_15810);
xnor U16726 (N_16726,N_15695,N_15636);
xor U16727 (N_16727,N_15849,N_15935);
and U16728 (N_16728,N_15446,N_16084);
nor U16729 (N_16729,N_15949,N_15973);
xnor U16730 (N_16730,N_15074,N_15929);
nand U16731 (N_16731,N_15435,N_16150);
xnor U16732 (N_16732,N_15219,N_16045);
nor U16733 (N_16733,N_15405,N_15508);
and U16734 (N_16734,N_15220,N_15812);
and U16735 (N_16735,N_15714,N_16217);
xnor U16736 (N_16736,N_15617,N_15738);
nand U16737 (N_16737,N_15227,N_15580);
or U16738 (N_16738,N_15317,N_15906);
nand U16739 (N_16739,N_16047,N_15805);
xor U16740 (N_16740,N_15137,N_15382);
or U16741 (N_16741,N_15948,N_15842);
nand U16742 (N_16742,N_15260,N_16015);
nand U16743 (N_16743,N_15191,N_16228);
nor U16744 (N_16744,N_15955,N_15061);
or U16745 (N_16745,N_15494,N_15197);
nand U16746 (N_16746,N_15167,N_16185);
and U16747 (N_16747,N_16043,N_16034);
nand U16748 (N_16748,N_16106,N_15682);
nand U16749 (N_16749,N_15749,N_15693);
nand U16750 (N_16750,N_16229,N_15741);
and U16751 (N_16751,N_15076,N_15832);
xor U16752 (N_16752,N_15792,N_15285);
nand U16753 (N_16753,N_16201,N_16248);
and U16754 (N_16754,N_16088,N_15371);
xnor U16755 (N_16755,N_15187,N_16016);
xor U16756 (N_16756,N_16103,N_15449);
nand U16757 (N_16757,N_15433,N_15476);
or U16758 (N_16758,N_15814,N_15489);
and U16759 (N_16759,N_16053,N_15785);
and U16760 (N_16760,N_15756,N_15994);
nor U16761 (N_16761,N_16209,N_15319);
xor U16762 (N_16762,N_15708,N_15923);
nor U16763 (N_16763,N_15095,N_15396);
xnor U16764 (N_16764,N_15330,N_16004);
or U16765 (N_16765,N_15385,N_15490);
or U16766 (N_16766,N_15536,N_16167);
xor U16767 (N_16767,N_15932,N_15560);
nand U16768 (N_16768,N_15196,N_15752);
xor U16769 (N_16769,N_16010,N_15213);
and U16770 (N_16770,N_15003,N_16193);
nand U16771 (N_16771,N_15770,N_15969);
and U16772 (N_16772,N_15154,N_15014);
xor U16773 (N_16773,N_15387,N_15954);
xnor U16774 (N_16774,N_15686,N_15999);
nor U16775 (N_16775,N_15515,N_15483);
nor U16776 (N_16776,N_15721,N_15313);
xor U16777 (N_16777,N_16200,N_15416);
or U16778 (N_16778,N_15347,N_15577);
nand U16779 (N_16779,N_16006,N_16208);
or U16780 (N_16780,N_15765,N_15550);
and U16781 (N_16781,N_15438,N_15138);
and U16782 (N_16782,N_15189,N_15119);
or U16783 (N_16783,N_15423,N_15043);
nor U16784 (N_16784,N_15846,N_15486);
nand U16785 (N_16785,N_15091,N_15683);
nand U16786 (N_16786,N_15270,N_16165);
nor U16787 (N_16787,N_15511,N_16041);
and U16788 (N_16788,N_15359,N_16090);
nor U16789 (N_16789,N_15899,N_15269);
or U16790 (N_16790,N_15914,N_15136);
and U16791 (N_16791,N_15172,N_15783);
nor U16792 (N_16792,N_15118,N_15394);
and U16793 (N_16793,N_15294,N_16079);
nor U16794 (N_16794,N_15982,N_16033);
and U16795 (N_16795,N_15958,N_15475);
xor U16796 (N_16796,N_16039,N_15947);
and U16797 (N_16797,N_15380,N_16214);
or U16798 (N_16798,N_15289,N_15290);
xor U16799 (N_16799,N_15318,N_15890);
or U16800 (N_16800,N_15869,N_15676);
nor U16801 (N_16801,N_15901,N_15147);
nand U16802 (N_16802,N_16213,N_16170);
nand U16803 (N_16803,N_15448,N_15310);
or U16804 (N_16804,N_15894,N_15252);
and U16805 (N_16805,N_15045,N_15534);
nor U16806 (N_16806,N_15364,N_15326);
nor U16807 (N_16807,N_15389,N_15757);
nand U16808 (N_16808,N_15891,N_15671);
or U16809 (N_16809,N_16073,N_15082);
nand U16810 (N_16810,N_16098,N_15509);
nand U16811 (N_16811,N_15956,N_16132);
nor U16812 (N_16812,N_15605,N_15398);
or U16813 (N_16813,N_15469,N_16067);
xnor U16814 (N_16814,N_15808,N_16023);
nor U16815 (N_16815,N_15092,N_16124);
xor U16816 (N_16816,N_15724,N_15529);
nand U16817 (N_16817,N_15058,N_15768);
nand U16818 (N_16818,N_15526,N_16146);
or U16819 (N_16819,N_15029,N_15861);
or U16820 (N_16820,N_15946,N_16225);
and U16821 (N_16821,N_15624,N_15301);
nor U16822 (N_16822,N_15109,N_15649);
and U16823 (N_16823,N_16050,N_15734);
or U16824 (N_16824,N_15985,N_15629);
nand U16825 (N_16825,N_15930,N_15299);
nand U16826 (N_16826,N_15180,N_15590);
nor U16827 (N_16827,N_16031,N_15599);
and U16828 (N_16828,N_15493,N_15075);
and U16829 (N_16829,N_15144,N_15582);
xnor U16830 (N_16830,N_15039,N_15941);
nor U16831 (N_16831,N_15533,N_15817);
or U16832 (N_16832,N_15302,N_15271);
nand U16833 (N_16833,N_15718,N_16035);
xor U16834 (N_16834,N_16191,N_15620);
and U16835 (N_16835,N_16018,N_15481);
nand U16836 (N_16836,N_16166,N_15460);
and U16837 (N_16837,N_15022,N_16104);
or U16838 (N_16838,N_15356,N_16066);
nor U16839 (N_16839,N_15018,N_16095);
nand U16840 (N_16840,N_15420,N_15181);
nand U16841 (N_16841,N_15648,N_15306);
nand U16842 (N_16842,N_15479,N_15296);
xnor U16843 (N_16843,N_15690,N_15159);
nor U16844 (N_16844,N_16224,N_15462);
or U16845 (N_16845,N_15938,N_15727);
xor U16846 (N_16846,N_15204,N_15698);
and U16847 (N_16847,N_16184,N_15070);
and U16848 (N_16848,N_16158,N_15806);
nand U16849 (N_16849,N_15504,N_15474);
nor U16850 (N_16850,N_15324,N_15308);
nand U16851 (N_16851,N_15233,N_15079);
nand U16852 (N_16852,N_15391,N_16242);
or U16853 (N_16853,N_15145,N_15257);
or U16854 (N_16854,N_15530,N_15818);
xnor U16855 (N_16855,N_16024,N_15431);
nor U16856 (N_16856,N_15848,N_15042);
or U16857 (N_16857,N_15688,N_15078);
nor U16858 (N_16858,N_15307,N_15251);
nor U16859 (N_16859,N_15793,N_16163);
nor U16860 (N_16860,N_15120,N_16240);
and U16861 (N_16861,N_15099,N_16032);
nor U16862 (N_16862,N_16086,N_15870);
or U16863 (N_16863,N_15367,N_15644);
or U16864 (N_16864,N_15875,N_16160);
nand U16865 (N_16865,N_15273,N_15576);
or U16866 (N_16866,N_16232,N_15340);
or U16867 (N_16867,N_15558,N_16187);
xor U16868 (N_16868,N_15468,N_15336);
and U16869 (N_16869,N_15242,N_15348);
nor U16870 (N_16870,N_15921,N_15256);
xnor U16871 (N_16871,N_15390,N_15176);
nand U16872 (N_16872,N_15656,N_15403);
or U16873 (N_16873,N_15477,N_15456);
xnor U16874 (N_16874,N_15401,N_15496);
or U16875 (N_16875,N_15568,N_15739);
or U16876 (N_16876,N_15079,N_15320);
xnor U16877 (N_16877,N_15682,N_15723);
and U16878 (N_16878,N_15119,N_15193);
and U16879 (N_16879,N_15965,N_15890);
nand U16880 (N_16880,N_15650,N_15013);
or U16881 (N_16881,N_15689,N_16036);
nand U16882 (N_16882,N_15296,N_15651);
nand U16883 (N_16883,N_15386,N_15635);
or U16884 (N_16884,N_15206,N_15568);
nor U16885 (N_16885,N_15532,N_15665);
and U16886 (N_16886,N_15951,N_15905);
and U16887 (N_16887,N_16166,N_15837);
nor U16888 (N_16888,N_15712,N_16177);
and U16889 (N_16889,N_15383,N_15019);
nand U16890 (N_16890,N_15382,N_15963);
nand U16891 (N_16891,N_15492,N_15644);
or U16892 (N_16892,N_15200,N_15084);
xor U16893 (N_16893,N_16024,N_16093);
nand U16894 (N_16894,N_15081,N_15126);
and U16895 (N_16895,N_15963,N_15153);
and U16896 (N_16896,N_16021,N_15808);
nand U16897 (N_16897,N_15484,N_15240);
nand U16898 (N_16898,N_16172,N_15603);
nor U16899 (N_16899,N_15417,N_15757);
nand U16900 (N_16900,N_15660,N_15932);
and U16901 (N_16901,N_15574,N_15852);
nor U16902 (N_16902,N_15801,N_15449);
and U16903 (N_16903,N_15740,N_15620);
nand U16904 (N_16904,N_15677,N_15089);
or U16905 (N_16905,N_16078,N_15364);
nor U16906 (N_16906,N_15717,N_15895);
and U16907 (N_16907,N_15586,N_16158);
xnor U16908 (N_16908,N_16012,N_15754);
nand U16909 (N_16909,N_15626,N_15632);
and U16910 (N_16910,N_15896,N_16007);
or U16911 (N_16911,N_15134,N_15362);
and U16912 (N_16912,N_15776,N_16099);
xnor U16913 (N_16913,N_15788,N_15513);
nor U16914 (N_16914,N_15153,N_15925);
or U16915 (N_16915,N_15457,N_15331);
xor U16916 (N_16916,N_16081,N_15466);
nand U16917 (N_16917,N_15462,N_15997);
or U16918 (N_16918,N_16144,N_16125);
and U16919 (N_16919,N_15841,N_15387);
and U16920 (N_16920,N_16188,N_15114);
xor U16921 (N_16921,N_15565,N_15628);
and U16922 (N_16922,N_15949,N_15706);
nor U16923 (N_16923,N_15145,N_15536);
xor U16924 (N_16924,N_15874,N_16246);
xnor U16925 (N_16925,N_15771,N_15727);
nor U16926 (N_16926,N_15090,N_15397);
and U16927 (N_16927,N_15245,N_15968);
nand U16928 (N_16928,N_16124,N_15934);
or U16929 (N_16929,N_15535,N_15311);
xnor U16930 (N_16930,N_15112,N_15168);
xnor U16931 (N_16931,N_16115,N_15757);
and U16932 (N_16932,N_15352,N_15368);
nand U16933 (N_16933,N_15080,N_15781);
or U16934 (N_16934,N_15459,N_16240);
and U16935 (N_16935,N_15357,N_15826);
or U16936 (N_16936,N_15879,N_15156);
nor U16937 (N_16937,N_15134,N_15676);
xor U16938 (N_16938,N_15369,N_15325);
or U16939 (N_16939,N_15885,N_15591);
nand U16940 (N_16940,N_15559,N_15948);
nand U16941 (N_16941,N_15582,N_15456);
or U16942 (N_16942,N_15269,N_15740);
xnor U16943 (N_16943,N_15508,N_15826);
xnor U16944 (N_16944,N_15525,N_15027);
xnor U16945 (N_16945,N_15174,N_15554);
or U16946 (N_16946,N_15014,N_15328);
nor U16947 (N_16947,N_15397,N_15913);
nand U16948 (N_16948,N_15952,N_15750);
and U16949 (N_16949,N_15795,N_15089);
nand U16950 (N_16950,N_16067,N_15155);
or U16951 (N_16951,N_15897,N_16023);
nand U16952 (N_16952,N_15618,N_16096);
xor U16953 (N_16953,N_15472,N_15104);
and U16954 (N_16954,N_15951,N_15486);
nor U16955 (N_16955,N_15438,N_15833);
xor U16956 (N_16956,N_16099,N_15539);
nand U16957 (N_16957,N_15015,N_15992);
or U16958 (N_16958,N_15657,N_15939);
and U16959 (N_16959,N_15870,N_15024);
or U16960 (N_16960,N_15796,N_15266);
and U16961 (N_16961,N_15273,N_15585);
nand U16962 (N_16962,N_15325,N_16151);
nor U16963 (N_16963,N_15343,N_16125);
nand U16964 (N_16964,N_15445,N_15608);
nor U16965 (N_16965,N_15528,N_15366);
nor U16966 (N_16966,N_15269,N_16050);
nor U16967 (N_16967,N_15736,N_15699);
or U16968 (N_16968,N_15820,N_15678);
xor U16969 (N_16969,N_15500,N_15760);
nand U16970 (N_16970,N_15332,N_16126);
nand U16971 (N_16971,N_16174,N_15066);
or U16972 (N_16972,N_16144,N_15126);
and U16973 (N_16973,N_15131,N_15622);
or U16974 (N_16974,N_15329,N_15187);
xor U16975 (N_16975,N_16149,N_15466);
xnor U16976 (N_16976,N_15307,N_15798);
nand U16977 (N_16977,N_15274,N_15704);
xnor U16978 (N_16978,N_15876,N_15740);
and U16979 (N_16979,N_15271,N_16186);
xor U16980 (N_16980,N_15827,N_16180);
xor U16981 (N_16981,N_15996,N_15737);
nor U16982 (N_16982,N_15098,N_15790);
and U16983 (N_16983,N_15127,N_15851);
or U16984 (N_16984,N_15107,N_15040);
or U16985 (N_16985,N_16022,N_15655);
nand U16986 (N_16986,N_15466,N_15457);
or U16987 (N_16987,N_15579,N_15469);
or U16988 (N_16988,N_15831,N_15237);
and U16989 (N_16989,N_15180,N_16094);
nand U16990 (N_16990,N_15224,N_15476);
xor U16991 (N_16991,N_16124,N_15226);
xor U16992 (N_16992,N_15273,N_15986);
xnor U16993 (N_16993,N_15950,N_15605);
nor U16994 (N_16994,N_16183,N_15691);
and U16995 (N_16995,N_15119,N_15240);
nor U16996 (N_16996,N_16029,N_15630);
xor U16997 (N_16997,N_15397,N_15112);
xnor U16998 (N_16998,N_15819,N_15471);
nand U16999 (N_16999,N_15788,N_15775);
xnor U17000 (N_17000,N_15561,N_15078);
and U17001 (N_17001,N_15328,N_16200);
or U17002 (N_17002,N_15635,N_15000);
or U17003 (N_17003,N_16223,N_15850);
xnor U17004 (N_17004,N_15556,N_16189);
or U17005 (N_17005,N_15651,N_15164);
nand U17006 (N_17006,N_15561,N_16091);
nor U17007 (N_17007,N_15480,N_15805);
xor U17008 (N_17008,N_16235,N_15423);
nand U17009 (N_17009,N_15538,N_15263);
xnor U17010 (N_17010,N_15002,N_15890);
nand U17011 (N_17011,N_15170,N_15923);
nor U17012 (N_17012,N_15195,N_15663);
nand U17013 (N_17013,N_15475,N_15536);
xor U17014 (N_17014,N_15538,N_15852);
xnor U17015 (N_17015,N_15254,N_16051);
nand U17016 (N_17016,N_15585,N_15281);
xor U17017 (N_17017,N_15321,N_15399);
nor U17018 (N_17018,N_15336,N_16041);
and U17019 (N_17019,N_15750,N_15308);
and U17020 (N_17020,N_15226,N_15786);
nand U17021 (N_17021,N_15254,N_15587);
nand U17022 (N_17022,N_15933,N_15325);
xnor U17023 (N_17023,N_15648,N_15071);
xnor U17024 (N_17024,N_16098,N_15317);
and U17025 (N_17025,N_15998,N_15758);
nand U17026 (N_17026,N_16217,N_15586);
nor U17027 (N_17027,N_15519,N_15306);
or U17028 (N_17028,N_15727,N_16091);
xnor U17029 (N_17029,N_15689,N_15052);
and U17030 (N_17030,N_15083,N_15903);
nand U17031 (N_17031,N_15409,N_16110);
nand U17032 (N_17032,N_15282,N_15813);
and U17033 (N_17033,N_15277,N_15259);
nand U17034 (N_17034,N_15632,N_15530);
or U17035 (N_17035,N_15009,N_15602);
xor U17036 (N_17036,N_15318,N_16028);
or U17037 (N_17037,N_15423,N_15902);
and U17038 (N_17038,N_15817,N_16164);
xor U17039 (N_17039,N_15100,N_15701);
nand U17040 (N_17040,N_15701,N_15833);
nand U17041 (N_17041,N_15627,N_15958);
or U17042 (N_17042,N_16187,N_15500);
or U17043 (N_17043,N_15518,N_15885);
nand U17044 (N_17044,N_15020,N_15062);
nand U17045 (N_17045,N_15527,N_16235);
and U17046 (N_17046,N_15565,N_16057);
xnor U17047 (N_17047,N_15360,N_15499);
and U17048 (N_17048,N_16165,N_15570);
xnor U17049 (N_17049,N_15663,N_15521);
nor U17050 (N_17050,N_15063,N_15790);
and U17051 (N_17051,N_15328,N_15972);
and U17052 (N_17052,N_15362,N_15973);
nand U17053 (N_17053,N_15708,N_16026);
xor U17054 (N_17054,N_15280,N_16108);
and U17055 (N_17055,N_16247,N_15357);
nor U17056 (N_17056,N_16207,N_15133);
xor U17057 (N_17057,N_15069,N_15273);
and U17058 (N_17058,N_15257,N_15685);
nor U17059 (N_17059,N_15211,N_15642);
and U17060 (N_17060,N_15709,N_15217);
nand U17061 (N_17061,N_15007,N_16227);
xor U17062 (N_17062,N_15078,N_15672);
xor U17063 (N_17063,N_15686,N_16109);
or U17064 (N_17064,N_15708,N_15614);
xnor U17065 (N_17065,N_15557,N_15390);
nor U17066 (N_17066,N_15844,N_16187);
xor U17067 (N_17067,N_15124,N_16227);
nor U17068 (N_17068,N_15096,N_15238);
xor U17069 (N_17069,N_15305,N_15557);
xor U17070 (N_17070,N_15648,N_16217);
nor U17071 (N_17071,N_15980,N_15607);
nand U17072 (N_17072,N_15595,N_15957);
or U17073 (N_17073,N_15498,N_15579);
or U17074 (N_17074,N_15256,N_15594);
nor U17075 (N_17075,N_15073,N_15801);
nor U17076 (N_17076,N_15750,N_15936);
or U17077 (N_17077,N_15582,N_15853);
or U17078 (N_17078,N_16181,N_15735);
or U17079 (N_17079,N_15441,N_15353);
or U17080 (N_17080,N_15636,N_15377);
or U17081 (N_17081,N_15332,N_15781);
or U17082 (N_17082,N_15458,N_15632);
nand U17083 (N_17083,N_15776,N_15837);
nor U17084 (N_17084,N_15559,N_15078);
xor U17085 (N_17085,N_15323,N_16033);
xnor U17086 (N_17086,N_15406,N_15968);
nand U17087 (N_17087,N_16020,N_15418);
nor U17088 (N_17088,N_15780,N_15959);
nand U17089 (N_17089,N_15574,N_15884);
nand U17090 (N_17090,N_15987,N_16102);
and U17091 (N_17091,N_15595,N_15846);
nor U17092 (N_17092,N_15078,N_16104);
xor U17093 (N_17093,N_15196,N_15540);
and U17094 (N_17094,N_16063,N_15197);
and U17095 (N_17095,N_15164,N_15855);
nand U17096 (N_17096,N_15861,N_15674);
nor U17097 (N_17097,N_15676,N_15963);
nand U17098 (N_17098,N_15001,N_15778);
nor U17099 (N_17099,N_15066,N_15917);
and U17100 (N_17100,N_16222,N_16035);
or U17101 (N_17101,N_15271,N_15053);
nor U17102 (N_17102,N_16133,N_16228);
xnor U17103 (N_17103,N_15744,N_16187);
or U17104 (N_17104,N_15100,N_16046);
xor U17105 (N_17105,N_15758,N_16150);
and U17106 (N_17106,N_15994,N_15981);
xor U17107 (N_17107,N_15001,N_15781);
xor U17108 (N_17108,N_15523,N_15673);
or U17109 (N_17109,N_15750,N_15272);
nor U17110 (N_17110,N_15683,N_15857);
xor U17111 (N_17111,N_15546,N_15330);
and U17112 (N_17112,N_16096,N_15266);
or U17113 (N_17113,N_15312,N_15459);
nand U17114 (N_17114,N_15278,N_15188);
xnor U17115 (N_17115,N_15739,N_16204);
or U17116 (N_17116,N_16095,N_15354);
and U17117 (N_17117,N_15577,N_15293);
xnor U17118 (N_17118,N_15473,N_15989);
or U17119 (N_17119,N_15478,N_15065);
nor U17120 (N_17120,N_16224,N_15703);
and U17121 (N_17121,N_15131,N_15801);
nand U17122 (N_17122,N_15825,N_15557);
nand U17123 (N_17123,N_16231,N_15743);
nand U17124 (N_17124,N_15632,N_15862);
nor U17125 (N_17125,N_16138,N_15760);
nor U17126 (N_17126,N_15947,N_16132);
nand U17127 (N_17127,N_15943,N_16091);
or U17128 (N_17128,N_15651,N_15167);
or U17129 (N_17129,N_15266,N_15118);
or U17130 (N_17130,N_15504,N_15147);
xnor U17131 (N_17131,N_15318,N_15103);
xor U17132 (N_17132,N_15217,N_15190);
and U17133 (N_17133,N_15735,N_15793);
nand U17134 (N_17134,N_15603,N_15384);
xnor U17135 (N_17135,N_16005,N_15682);
or U17136 (N_17136,N_15553,N_16049);
or U17137 (N_17137,N_15174,N_15544);
nand U17138 (N_17138,N_16209,N_15349);
nand U17139 (N_17139,N_16211,N_16156);
nor U17140 (N_17140,N_15463,N_15206);
nor U17141 (N_17141,N_15276,N_16244);
or U17142 (N_17142,N_16214,N_15203);
nand U17143 (N_17143,N_15626,N_16107);
or U17144 (N_17144,N_15715,N_15830);
nor U17145 (N_17145,N_15175,N_15064);
and U17146 (N_17146,N_16039,N_15395);
or U17147 (N_17147,N_15369,N_16158);
xnor U17148 (N_17148,N_15930,N_15102);
xnor U17149 (N_17149,N_15099,N_15265);
and U17150 (N_17150,N_15799,N_16015);
nor U17151 (N_17151,N_15382,N_15127);
nor U17152 (N_17152,N_15642,N_15785);
and U17153 (N_17153,N_16157,N_16128);
nand U17154 (N_17154,N_15077,N_15475);
or U17155 (N_17155,N_15147,N_15536);
and U17156 (N_17156,N_15925,N_15808);
or U17157 (N_17157,N_15714,N_15462);
or U17158 (N_17158,N_16152,N_16228);
and U17159 (N_17159,N_16173,N_15392);
nand U17160 (N_17160,N_15243,N_16061);
xnor U17161 (N_17161,N_15364,N_15021);
nand U17162 (N_17162,N_15187,N_15084);
nand U17163 (N_17163,N_15072,N_15893);
or U17164 (N_17164,N_16183,N_15542);
nor U17165 (N_17165,N_15135,N_15843);
nor U17166 (N_17166,N_15437,N_15425);
nand U17167 (N_17167,N_15134,N_15349);
xnor U17168 (N_17168,N_16165,N_16033);
or U17169 (N_17169,N_15063,N_16233);
and U17170 (N_17170,N_15404,N_15476);
and U17171 (N_17171,N_16092,N_15361);
nand U17172 (N_17172,N_15103,N_15295);
nor U17173 (N_17173,N_16029,N_15431);
xnor U17174 (N_17174,N_15737,N_15258);
and U17175 (N_17175,N_15790,N_15726);
xor U17176 (N_17176,N_15781,N_16094);
and U17177 (N_17177,N_15836,N_15721);
nor U17178 (N_17178,N_16017,N_16075);
or U17179 (N_17179,N_15014,N_15582);
and U17180 (N_17180,N_15539,N_16023);
nand U17181 (N_17181,N_15840,N_15804);
xnor U17182 (N_17182,N_16235,N_15333);
nand U17183 (N_17183,N_15031,N_15779);
xor U17184 (N_17184,N_15387,N_15969);
and U17185 (N_17185,N_15214,N_16210);
nor U17186 (N_17186,N_15997,N_16238);
nor U17187 (N_17187,N_15829,N_15013);
nor U17188 (N_17188,N_15723,N_16085);
xor U17189 (N_17189,N_15565,N_15700);
and U17190 (N_17190,N_15518,N_15209);
nor U17191 (N_17191,N_16019,N_15490);
xnor U17192 (N_17192,N_15821,N_16134);
or U17193 (N_17193,N_15116,N_15956);
nor U17194 (N_17194,N_15632,N_15506);
xnor U17195 (N_17195,N_15475,N_16225);
and U17196 (N_17196,N_16109,N_15459);
nor U17197 (N_17197,N_15439,N_15501);
or U17198 (N_17198,N_15979,N_15848);
and U17199 (N_17199,N_15389,N_16130);
nor U17200 (N_17200,N_15008,N_15312);
and U17201 (N_17201,N_16138,N_16199);
xor U17202 (N_17202,N_15819,N_15588);
nand U17203 (N_17203,N_15069,N_15045);
nand U17204 (N_17204,N_16011,N_15472);
nor U17205 (N_17205,N_15932,N_16104);
xnor U17206 (N_17206,N_15362,N_15024);
xor U17207 (N_17207,N_15193,N_15699);
xor U17208 (N_17208,N_15853,N_15982);
nor U17209 (N_17209,N_16245,N_15226);
xor U17210 (N_17210,N_15678,N_15003);
xnor U17211 (N_17211,N_16157,N_15287);
or U17212 (N_17212,N_15087,N_16172);
nand U17213 (N_17213,N_16183,N_15281);
or U17214 (N_17214,N_16076,N_15041);
nor U17215 (N_17215,N_15141,N_16072);
xnor U17216 (N_17216,N_15242,N_15041);
nor U17217 (N_17217,N_15947,N_15880);
and U17218 (N_17218,N_15639,N_16165);
nor U17219 (N_17219,N_16169,N_16194);
nand U17220 (N_17220,N_15395,N_15785);
nand U17221 (N_17221,N_16187,N_15743);
xnor U17222 (N_17222,N_16015,N_15237);
or U17223 (N_17223,N_15570,N_15148);
or U17224 (N_17224,N_15520,N_15091);
and U17225 (N_17225,N_16247,N_16231);
nand U17226 (N_17226,N_15930,N_15032);
xor U17227 (N_17227,N_15094,N_15532);
nand U17228 (N_17228,N_15046,N_15649);
nand U17229 (N_17229,N_15640,N_15143);
xnor U17230 (N_17230,N_15698,N_15945);
and U17231 (N_17231,N_15012,N_15544);
xnor U17232 (N_17232,N_15449,N_15874);
and U17233 (N_17233,N_15599,N_15794);
nand U17234 (N_17234,N_15534,N_15904);
nor U17235 (N_17235,N_15777,N_15479);
or U17236 (N_17236,N_15582,N_15974);
or U17237 (N_17237,N_16086,N_15043);
or U17238 (N_17238,N_15191,N_15933);
nor U17239 (N_17239,N_15005,N_15861);
and U17240 (N_17240,N_15236,N_16243);
xnor U17241 (N_17241,N_16248,N_15768);
nor U17242 (N_17242,N_15932,N_15971);
and U17243 (N_17243,N_15976,N_16132);
and U17244 (N_17244,N_15134,N_15876);
nand U17245 (N_17245,N_15434,N_15603);
or U17246 (N_17246,N_15821,N_15720);
xnor U17247 (N_17247,N_15100,N_15407);
nand U17248 (N_17248,N_15432,N_15830);
and U17249 (N_17249,N_15586,N_15467);
and U17250 (N_17250,N_15778,N_15532);
nor U17251 (N_17251,N_15358,N_15700);
and U17252 (N_17252,N_15816,N_15733);
nor U17253 (N_17253,N_15827,N_15696);
nand U17254 (N_17254,N_15009,N_15829);
xor U17255 (N_17255,N_15357,N_16034);
nand U17256 (N_17256,N_15962,N_15694);
xor U17257 (N_17257,N_15772,N_15953);
nor U17258 (N_17258,N_15906,N_15713);
nand U17259 (N_17259,N_16201,N_15977);
nor U17260 (N_17260,N_15811,N_15969);
or U17261 (N_17261,N_16181,N_15029);
and U17262 (N_17262,N_15272,N_16217);
nor U17263 (N_17263,N_16136,N_16049);
xor U17264 (N_17264,N_15766,N_15780);
and U17265 (N_17265,N_16150,N_15781);
or U17266 (N_17266,N_15794,N_15139);
nand U17267 (N_17267,N_16163,N_15696);
or U17268 (N_17268,N_16008,N_15915);
or U17269 (N_17269,N_15653,N_15988);
or U17270 (N_17270,N_16086,N_15136);
xnor U17271 (N_17271,N_15681,N_15422);
nand U17272 (N_17272,N_15654,N_15823);
xor U17273 (N_17273,N_15606,N_15545);
nand U17274 (N_17274,N_15170,N_15184);
nor U17275 (N_17275,N_15002,N_15866);
or U17276 (N_17276,N_15530,N_16223);
nor U17277 (N_17277,N_15008,N_15928);
or U17278 (N_17278,N_15686,N_15260);
nor U17279 (N_17279,N_15693,N_15457);
or U17280 (N_17280,N_15194,N_15170);
xor U17281 (N_17281,N_16011,N_15176);
nand U17282 (N_17282,N_16123,N_15250);
nand U17283 (N_17283,N_15271,N_15581);
nand U17284 (N_17284,N_15183,N_15643);
nand U17285 (N_17285,N_15016,N_16246);
xnor U17286 (N_17286,N_16248,N_15133);
xor U17287 (N_17287,N_15867,N_15640);
nor U17288 (N_17288,N_15359,N_16182);
or U17289 (N_17289,N_16000,N_15461);
or U17290 (N_17290,N_15386,N_15329);
nor U17291 (N_17291,N_15069,N_15378);
and U17292 (N_17292,N_15007,N_15409);
and U17293 (N_17293,N_15615,N_15861);
and U17294 (N_17294,N_15389,N_16028);
nor U17295 (N_17295,N_15577,N_15416);
xor U17296 (N_17296,N_15778,N_16114);
nand U17297 (N_17297,N_15742,N_15611);
or U17298 (N_17298,N_16229,N_15937);
or U17299 (N_17299,N_15153,N_15690);
and U17300 (N_17300,N_15481,N_16141);
and U17301 (N_17301,N_15265,N_16090);
nor U17302 (N_17302,N_15874,N_15296);
and U17303 (N_17303,N_16127,N_16105);
and U17304 (N_17304,N_15050,N_15720);
and U17305 (N_17305,N_15382,N_16135);
and U17306 (N_17306,N_15367,N_15438);
xor U17307 (N_17307,N_16059,N_15362);
nor U17308 (N_17308,N_15890,N_15716);
nand U17309 (N_17309,N_15271,N_16065);
nor U17310 (N_17310,N_15580,N_16017);
xor U17311 (N_17311,N_15227,N_15388);
xnor U17312 (N_17312,N_15998,N_15316);
nor U17313 (N_17313,N_15362,N_15649);
and U17314 (N_17314,N_15241,N_15007);
nand U17315 (N_17315,N_15477,N_16168);
or U17316 (N_17316,N_15798,N_15241);
or U17317 (N_17317,N_15518,N_15121);
nand U17318 (N_17318,N_16128,N_15571);
or U17319 (N_17319,N_16061,N_15161);
xnor U17320 (N_17320,N_15855,N_16091);
or U17321 (N_17321,N_15541,N_15233);
or U17322 (N_17322,N_15945,N_16230);
or U17323 (N_17323,N_15603,N_16219);
and U17324 (N_17324,N_15753,N_15499);
and U17325 (N_17325,N_16053,N_15118);
nand U17326 (N_17326,N_16080,N_15681);
xnor U17327 (N_17327,N_15739,N_15625);
xor U17328 (N_17328,N_15382,N_15996);
nand U17329 (N_17329,N_16104,N_15774);
nand U17330 (N_17330,N_16180,N_15738);
nand U17331 (N_17331,N_15346,N_16219);
xor U17332 (N_17332,N_15171,N_15805);
and U17333 (N_17333,N_15071,N_15814);
and U17334 (N_17334,N_16189,N_16243);
and U17335 (N_17335,N_15186,N_15488);
nand U17336 (N_17336,N_15100,N_15656);
and U17337 (N_17337,N_15127,N_16182);
nor U17338 (N_17338,N_15015,N_15495);
xnor U17339 (N_17339,N_16200,N_15152);
nand U17340 (N_17340,N_15854,N_15689);
and U17341 (N_17341,N_15844,N_15538);
and U17342 (N_17342,N_15555,N_15636);
or U17343 (N_17343,N_15075,N_15728);
nand U17344 (N_17344,N_16139,N_15603);
nand U17345 (N_17345,N_15598,N_15668);
or U17346 (N_17346,N_15552,N_15773);
nand U17347 (N_17347,N_15370,N_15364);
nor U17348 (N_17348,N_15523,N_16059);
nand U17349 (N_17349,N_15557,N_15217);
or U17350 (N_17350,N_15414,N_16111);
xnor U17351 (N_17351,N_15569,N_15171);
nor U17352 (N_17352,N_15103,N_16028);
xnor U17353 (N_17353,N_15680,N_15193);
and U17354 (N_17354,N_15313,N_16248);
nor U17355 (N_17355,N_15714,N_15361);
or U17356 (N_17356,N_15581,N_15751);
and U17357 (N_17357,N_15663,N_16081);
nand U17358 (N_17358,N_15982,N_15722);
and U17359 (N_17359,N_15019,N_15986);
xor U17360 (N_17360,N_15318,N_15364);
nand U17361 (N_17361,N_15105,N_15243);
and U17362 (N_17362,N_15169,N_16238);
xor U17363 (N_17363,N_16123,N_16166);
nand U17364 (N_17364,N_15450,N_15720);
xnor U17365 (N_17365,N_15813,N_15499);
or U17366 (N_17366,N_15970,N_16183);
xor U17367 (N_17367,N_15783,N_16032);
and U17368 (N_17368,N_15820,N_15091);
and U17369 (N_17369,N_16143,N_15650);
xnor U17370 (N_17370,N_15560,N_15581);
nor U17371 (N_17371,N_15410,N_15309);
xor U17372 (N_17372,N_16050,N_15316);
nand U17373 (N_17373,N_15485,N_15618);
nand U17374 (N_17374,N_15678,N_15766);
xnor U17375 (N_17375,N_15541,N_16031);
nor U17376 (N_17376,N_15581,N_15887);
nand U17377 (N_17377,N_15722,N_16092);
nand U17378 (N_17378,N_16187,N_15932);
nor U17379 (N_17379,N_15786,N_15766);
nand U17380 (N_17380,N_15135,N_15449);
nor U17381 (N_17381,N_15045,N_15477);
and U17382 (N_17382,N_15828,N_15276);
xor U17383 (N_17383,N_15624,N_15892);
nand U17384 (N_17384,N_15609,N_15672);
nor U17385 (N_17385,N_15233,N_15107);
nand U17386 (N_17386,N_15168,N_15915);
or U17387 (N_17387,N_15467,N_15260);
nor U17388 (N_17388,N_15821,N_15644);
xor U17389 (N_17389,N_15488,N_15414);
xor U17390 (N_17390,N_16230,N_15901);
or U17391 (N_17391,N_15168,N_15959);
and U17392 (N_17392,N_15391,N_15529);
and U17393 (N_17393,N_15757,N_15527);
or U17394 (N_17394,N_15352,N_15082);
nand U17395 (N_17395,N_15006,N_15926);
or U17396 (N_17396,N_16090,N_16191);
and U17397 (N_17397,N_15669,N_16081);
and U17398 (N_17398,N_15138,N_15041);
xor U17399 (N_17399,N_15841,N_15110);
nor U17400 (N_17400,N_16212,N_15444);
or U17401 (N_17401,N_15325,N_15020);
nor U17402 (N_17402,N_15686,N_15578);
nor U17403 (N_17403,N_15399,N_15262);
nand U17404 (N_17404,N_15610,N_15210);
or U17405 (N_17405,N_15136,N_16201);
xor U17406 (N_17406,N_15574,N_15309);
or U17407 (N_17407,N_15358,N_16127);
or U17408 (N_17408,N_16217,N_15619);
or U17409 (N_17409,N_15087,N_15972);
and U17410 (N_17410,N_15209,N_15330);
xnor U17411 (N_17411,N_15753,N_15420);
nand U17412 (N_17412,N_15623,N_15001);
and U17413 (N_17413,N_15611,N_16139);
and U17414 (N_17414,N_15591,N_15540);
and U17415 (N_17415,N_15514,N_15784);
or U17416 (N_17416,N_15831,N_15688);
or U17417 (N_17417,N_15116,N_15841);
nand U17418 (N_17418,N_16044,N_16022);
xnor U17419 (N_17419,N_15102,N_15438);
and U17420 (N_17420,N_16219,N_15170);
nor U17421 (N_17421,N_15913,N_15658);
nand U17422 (N_17422,N_16034,N_15795);
nand U17423 (N_17423,N_15925,N_15608);
xor U17424 (N_17424,N_15367,N_15369);
or U17425 (N_17425,N_15435,N_15762);
nand U17426 (N_17426,N_15476,N_15281);
nand U17427 (N_17427,N_15025,N_16249);
and U17428 (N_17428,N_15249,N_15792);
or U17429 (N_17429,N_15728,N_15494);
nand U17430 (N_17430,N_15170,N_15494);
nand U17431 (N_17431,N_15334,N_15402);
or U17432 (N_17432,N_16117,N_15322);
nor U17433 (N_17433,N_15983,N_15606);
xor U17434 (N_17434,N_15581,N_15629);
or U17435 (N_17435,N_15616,N_15910);
xnor U17436 (N_17436,N_15282,N_15683);
xor U17437 (N_17437,N_15799,N_15395);
and U17438 (N_17438,N_16037,N_15364);
and U17439 (N_17439,N_16166,N_15083);
nand U17440 (N_17440,N_15411,N_15764);
nand U17441 (N_17441,N_15777,N_15605);
or U17442 (N_17442,N_15859,N_15090);
nor U17443 (N_17443,N_15829,N_15206);
xor U17444 (N_17444,N_16245,N_15168);
and U17445 (N_17445,N_15516,N_15715);
or U17446 (N_17446,N_15863,N_16008);
and U17447 (N_17447,N_15276,N_15462);
or U17448 (N_17448,N_16005,N_16127);
xnor U17449 (N_17449,N_15189,N_15852);
nand U17450 (N_17450,N_15693,N_15159);
nand U17451 (N_17451,N_15709,N_15855);
or U17452 (N_17452,N_16020,N_15460);
nand U17453 (N_17453,N_15286,N_16096);
xor U17454 (N_17454,N_15466,N_16108);
nand U17455 (N_17455,N_15542,N_16115);
nand U17456 (N_17456,N_15477,N_15084);
nor U17457 (N_17457,N_15349,N_16117);
or U17458 (N_17458,N_15688,N_15808);
or U17459 (N_17459,N_15999,N_15980);
and U17460 (N_17460,N_16235,N_16134);
and U17461 (N_17461,N_15388,N_15170);
nor U17462 (N_17462,N_15000,N_15721);
nand U17463 (N_17463,N_16100,N_15705);
and U17464 (N_17464,N_16216,N_15136);
and U17465 (N_17465,N_15860,N_15420);
nand U17466 (N_17466,N_15147,N_15898);
xor U17467 (N_17467,N_15501,N_15025);
nand U17468 (N_17468,N_16132,N_15698);
and U17469 (N_17469,N_15771,N_15249);
and U17470 (N_17470,N_16070,N_16109);
xnor U17471 (N_17471,N_15453,N_15229);
nand U17472 (N_17472,N_15569,N_16230);
or U17473 (N_17473,N_15569,N_15726);
or U17474 (N_17474,N_15805,N_15826);
and U17475 (N_17475,N_15975,N_15715);
and U17476 (N_17476,N_15843,N_15118);
and U17477 (N_17477,N_15472,N_15587);
nor U17478 (N_17478,N_15450,N_16204);
nor U17479 (N_17479,N_15370,N_15893);
nor U17480 (N_17480,N_16047,N_15440);
and U17481 (N_17481,N_16235,N_15122);
nand U17482 (N_17482,N_15344,N_15259);
nor U17483 (N_17483,N_15208,N_16108);
nor U17484 (N_17484,N_16141,N_16064);
and U17485 (N_17485,N_15049,N_15377);
and U17486 (N_17486,N_15564,N_15968);
nor U17487 (N_17487,N_16225,N_15808);
nand U17488 (N_17488,N_15151,N_15514);
and U17489 (N_17489,N_16188,N_15262);
nor U17490 (N_17490,N_15200,N_15129);
or U17491 (N_17491,N_15617,N_15524);
or U17492 (N_17492,N_15648,N_15462);
xor U17493 (N_17493,N_15150,N_15876);
and U17494 (N_17494,N_15062,N_15881);
nand U17495 (N_17495,N_15054,N_15843);
nand U17496 (N_17496,N_15516,N_15428);
and U17497 (N_17497,N_15311,N_16054);
and U17498 (N_17498,N_15868,N_15087);
and U17499 (N_17499,N_15489,N_16047);
or U17500 (N_17500,N_16433,N_16637);
xor U17501 (N_17501,N_16408,N_17054);
nand U17502 (N_17502,N_17333,N_16532);
nor U17503 (N_17503,N_16299,N_16293);
or U17504 (N_17504,N_17415,N_16785);
or U17505 (N_17505,N_17194,N_16465);
or U17506 (N_17506,N_16554,N_17081);
or U17507 (N_17507,N_17278,N_16324);
or U17508 (N_17508,N_16929,N_16603);
or U17509 (N_17509,N_16930,N_16625);
and U17510 (N_17510,N_17236,N_17344);
or U17511 (N_17511,N_17384,N_17040);
nor U17512 (N_17512,N_17075,N_16672);
xor U17513 (N_17513,N_17338,N_17347);
or U17514 (N_17514,N_17055,N_16996);
nor U17515 (N_17515,N_16970,N_16624);
nand U17516 (N_17516,N_17290,N_17188);
nor U17517 (N_17517,N_17206,N_16897);
or U17518 (N_17518,N_16535,N_16830);
xor U17519 (N_17519,N_16456,N_16254);
xor U17520 (N_17520,N_16478,N_17400);
nand U17521 (N_17521,N_17355,N_17108);
nor U17522 (N_17522,N_17392,N_16597);
xor U17523 (N_17523,N_17218,N_17080);
nand U17524 (N_17524,N_17135,N_17057);
nand U17525 (N_17525,N_17285,N_17133);
or U17526 (N_17526,N_16960,N_16656);
or U17527 (N_17527,N_16702,N_16833);
nand U17528 (N_17528,N_16419,N_17026);
and U17529 (N_17529,N_16923,N_16865);
xnor U17530 (N_17530,N_17237,N_17484);
xor U17531 (N_17531,N_16545,N_16959);
or U17532 (N_17532,N_17000,N_16466);
xnor U17533 (N_17533,N_17198,N_16718);
or U17534 (N_17534,N_17024,N_17065);
or U17535 (N_17535,N_17430,N_17136);
xor U17536 (N_17536,N_16315,N_16491);
xor U17537 (N_17537,N_16292,N_16990);
nand U17538 (N_17538,N_17303,N_17174);
and U17539 (N_17539,N_17014,N_16398);
or U17540 (N_17540,N_17009,N_16796);
and U17541 (N_17541,N_17429,N_16751);
and U17542 (N_17542,N_17359,N_16296);
xnor U17543 (N_17543,N_16778,N_16924);
nand U17544 (N_17544,N_17106,N_17342);
nand U17545 (N_17545,N_16260,N_16594);
xor U17546 (N_17546,N_16732,N_17177);
nand U17547 (N_17547,N_17271,N_16684);
or U17548 (N_17548,N_16514,N_17127);
or U17549 (N_17549,N_16703,N_16898);
nand U17550 (N_17550,N_16396,N_16876);
xor U17551 (N_17551,N_17300,N_16372);
nor U17552 (N_17552,N_17310,N_16522);
and U17553 (N_17553,N_16968,N_16673);
nor U17554 (N_17554,N_16497,N_17109);
nand U17555 (N_17555,N_16568,N_16352);
or U17556 (N_17556,N_16682,N_17451);
xnor U17557 (N_17557,N_17130,N_17002);
and U17558 (N_17558,N_16979,N_17191);
xnor U17559 (N_17559,N_17425,N_16854);
xor U17560 (N_17560,N_17072,N_16531);
nand U17561 (N_17561,N_16748,N_17197);
or U17562 (N_17562,N_17403,N_16861);
and U17563 (N_17563,N_17287,N_17454);
nand U17564 (N_17564,N_17131,N_16837);
xnor U17565 (N_17565,N_17043,N_16920);
and U17566 (N_17566,N_17469,N_16917);
and U17567 (N_17567,N_16492,N_16255);
or U17568 (N_17568,N_16540,N_16809);
nor U17569 (N_17569,N_17424,N_17047);
xnor U17570 (N_17570,N_17418,N_16948);
nor U17571 (N_17571,N_17156,N_17113);
or U17572 (N_17572,N_17143,N_16676);
or U17573 (N_17573,N_16328,N_17440);
and U17574 (N_17574,N_16366,N_17394);
and U17575 (N_17575,N_17378,N_16584);
nand U17576 (N_17576,N_16781,N_17281);
nand U17577 (N_17577,N_17193,N_17018);
nor U17578 (N_17578,N_16422,N_17439);
and U17579 (N_17579,N_17452,N_16390);
nand U17580 (N_17580,N_16411,N_17293);
or U17581 (N_17581,N_17094,N_16269);
nand U17582 (N_17582,N_17460,N_17207);
nor U17583 (N_17583,N_16504,N_17169);
and U17584 (N_17584,N_16526,N_17467);
and U17585 (N_17585,N_17395,N_17251);
nand U17586 (N_17586,N_16563,N_16459);
or U17587 (N_17587,N_17426,N_16721);
and U17588 (N_17588,N_16962,N_16883);
nor U17589 (N_17589,N_16641,N_17324);
nand U17590 (N_17590,N_16694,N_17099);
xor U17591 (N_17591,N_16601,N_17470);
nor U17592 (N_17592,N_16519,N_17150);
nor U17593 (N_17593,N_16952,N_16753);
nor U17594 (N_17594,N_16734,N_17192);
nand U17595 (N_17595,N_16450,N_16683);
and U17596 (N_17596,N_17398,N_17462);
xnor U17597 (N_17597,N_16481,N_17337);
xor U17598 (N_17598,N_17435,N_16868);
or U17599 (N_17599,N_16974,N_17004);
xor U17600 (N_17600,N_17168,N_16725);
and U17601 (N_17601,N_16783,N_17480);
nand U17602 (N_17602,N_17098,N_16453);
xor U17603 (N_17603,N_17475,N_16512);
or U17604 (N_17604,N_17120,N_17297);
and U17605 (N_17605,N_16349,N_16815);
and U17606 (N_17606,N_16770,N_16558);
nor U17607 (N_17607,N_17468,N_16602);
and U17608 (N_17608,N_17496,N_17352);
nand U17609 (N_17609,N_17119,N_17114);
nand U17610 (N_17610,N_17204,N_17471);
or U17611 (N_17611,N_16280,N_16393);
nand U17612 (N_17612,N_17361,N_17404);
or U17613 (N_17613,N_17298,N_17301);
nor U17614 (N_17614,N_16319,N_16376);
or U17615 (N_17615,N_17226,N_16482);
nand U17616 (N_17616,N_16612,N_17128);
and U17617 (N_17617,N_16348,N_17005);
nor U17618 (N_17618,N_16832,N_16361);
and U17619 (N_17619,N_16967,N_16811);
or U17620 (N_17620,N_17124,N_16647);
nor U17621 (N_17621,N_16884,N_16759);
and U17622 (N_17622,N_17163,N_16981);
nand U17623 (N_17623,N_16617,N_16831);
nor U17624 (N_17624,N_17360,N_16928);
nor U17625 (N_17625,N_16304,N_16666);
and U17626 (N_17626,N_16891,N_17309);
or U17627 (N_17627,N_16580,N_17406);
and U17628 (N_17628,N_16992,N_16501);
xor U17629 (N_17629,N_16908,N_17195);
and U17630 (N_17630,N_17248,N_16600);
and U17631 (N_17631,N_16572,N_17368);
xnor U17632 (N_17632,N_17074,N_16305);
and U17633 (N_17633,N_17232,N_17134);
nand U17634 (N_17634,N_16590,N_16933);
nor U17635 (N_17635,N_17096,N_16303);
xnor U17636 (N_17636,N_16536,N_16417);
and U17637 (N_17637,N_16268,N_16586);
and U17638 (N_17638,N_16754,N_16511);
nand U17639 (N_17639,N_17048,N_16985);
nor U17640 (N_17640,N_16646,N_16388);
and U17641 (N_17641,N_16976,N_17147);
and U17642 (N_17642,N_16581,N_16705);
and U17643 (N_17643,N_17126,N_16921);
or U17644 (N_17644,N_16986,N_16687);
nor U17645 (N_17645,N_16316,N_17077);
nand U17646 (N_17646,N_16988,N_16307);
nand U17647 (N_17647,N_16740,N_17154);
xnor U17648 (N_17648,N_16932,N_16281);
nor U17649 (N_17649,N_16286,N_17386);
and U17650 (N_17650,N_16816,N_16351);
nand U17651 (N_17651,N_17388,N_16969);
nand U17652 (N_17652,N_17017,N_16670);
xnor U17653 (N_17653,N_16822,N_16464);
xnor U17654 (N_17654,N_16824,N_17222);
or U17655 (N_17655,N_17180,N_16791);
and U17656 (N_17656,N_16276,N_16378);
nand U17657 (N_17657,N_17046,N_16746);
nor U17658 (N_17658,N_17013,N_16297);
nand U17659 (N_17659,N_17068,N_16680);
nand U17660 (N_17660,N_17265,N_17350);
xnor U17661 (N_17661,N_16578,N_16631);
and U17662 (N_17662,N_17276,N_16652);
or U17663 (N_17663,N_16405,N_16318);
or U17664 (N_17664,N_16444,N_17159);
and U17665 (N_17665,N_16565,N_16437);
nand U17666 (N_17666,N_17042,N_17356);
and U17667 (N_17667,N_16452,N_17187);
nand U17668 (N_17668,N_17001,N_17443);
and U17669 (N_17669,N_16252,N_17292);
nand U17670 (N_17670,N_16493,N_16711);
or U17671 (N_17671,N_16915,N_16659);
nand U17672 (N_17672,N_16749,N_16851);
nand U17673 (N_17673,N_16345,N_17269);
nand U17674 (N_17674,N_16284,N_17267);
nor U17675 (N_17675,N_17070,N_17117);
nand U17676 (N_17676,N_17357,N_16760);
nand U17677 (N_17677,N_16724,N_17076);
nand U17678 (N_17678,N_17332,N_16454);
xnor U17679 (N_17679,N_17314,N_17489);
or U17680 (N_17680,N_17423,N_16779);
or U17681 (N_17681,N_16479,N_17030);
and U17682 (N_17682,N_17112,N_17259);
and U17683 (N_17683,N_16688,N_16424);
or U17684 (N_17684,N_17179,N_16742);
xnor U17685 (N_17685,N_17213,N_16495);
nand U17686 (N_17686,N_17358,N_16262);
nor U17687 (N_17687,N_16402,N_17302);
xor U17688 (N_17688,N_16954,N_16620);
nand U17689 (N_17689,N_16566,N_16812);
xor U17690 (N_17690,N_16692,N_16343);
and U17691 (N_17691,N_16731,N_16880);
nor U17692 (N_17692,N_16598,N_17479);
or U17693 (N_17693,N_17053,N_16889);
nand U17694 (N_17694,N_17405,N_17203);
xnor U17695 (N_17695,N_17160,N_16528);
xnor U17696 (N_17696,N_17478,N_16971);
and U17697 (N_17697,N_16485,N_17093);
xnor U17698 (N_17698,N_16523,N_17396);
xor U17699 (N_17699,N_17322,N_16775);
xor U17700 (N_17700,N_16313,N_16871);
nand U17701 (N_17701,N_17273,N_17086);
nand U17702 (N_17702,N_17421,N_16542);
nand U17703 (N_17703,N_17339,N_16342);
nand U17704 (N_17704,N_16642,N_16320);
nand U17705 (N_17705,N_16653,N_17158);
xor U17706 (N_17706,N_16685,N_16799);
or U17707 (N_17707,N_16657,N_16259);
xnor U17708 (N_17708,N_17308,N_16737);
and U17709 (N_17709,N_16729,N_17372);
xnor U17710 (N_17710,N_16606,N_16916);
xnor U17711 (N_17711,N_17370,N_17250);
xnor U17712 (N_17712,N_16382,N_16788);
nand U17713 (N_17713,N_17200,N_17363);
nor U17714 (N_17714,N_16829,N_17450);
nor U17715 (N_17715,N_16633,N_16364);
xor U17716 (N_17716,N_16604,N_16356);
nand U17717 (N_17717,N_16503,N_17381);
xnor U17718 (N_17718,N_16546,N_16384);
or U17719 (N_17719,N_16640,N_16322);
nand U17720 (N_17720,N_16622,N_17326);
and U17721 (N_17721,N_16525,N_16695);
xor U17722 (N_17722,N_17233,N_16573);
nor U17723 (N_17723,N_17211,N_16710);
nand U17724 (N_17724,N_16991,N_17049);
and U17725 (N_17725,N_16980,N_16906);
nand U17726 (N_17726,N_17167,N_16714);
xnor U17727 (N_17727,N_16644,N_17391);
or U17728 (N_17728,N_16965,N_16964);
nand U17729 (N_17729,N_17286,N_16850);
xor U17730 (N_17730,N_16945,N_17091);
nor U17731 (N_17731,N_16978,N_17428);
or U17732 (N_17732,N_17383,N_16505);
nor U17733 (N_17733,N_16432,N_17412);
or U17734 (N_17734,N_17064,N_16567);
nor U17735 (N_17735,N_16392,N_16807);
xor U17736 (N_17736,N_16870,N_16288);
xor U17737 (N_17737,N_16645,N_16490);
nor U17738 (N_17738,N_16669,N_16808);
xnor U17739 (N_17739,N_16311,N_17058);
or U17740 (N_17740,N_16671,N_16274);
nand U17741 (N_17741,N_16341,N_16258);
xnor U17742 (N_17742,N_16836,N_17264);
or U17743 (N_17743,N_17463,N_16613);
xor U17744 (N_17744,N_17183,N_17382);
nor U17745 (N_17745,N_17157,N_17092);
or U17746 (N_17746,N_17071,N_16776);
nand U17747 (N_17747,N_17051,N_16649);
or U17748 (N_17748,N_16368,N_16738);
or U17749 (N_17749,N_17353,N_16849);
nor U17750 (N_17750,N_17021,N_16661);
or U17751 (N_17751,N_16265,N_16943);
xnor U17752 (N_17752,N_16909,N_16530);
nand U17753 (N_17753,N_16263,N_16386);
or U17754 (N_17754,N_16484,N_17012);
or U17755 (N_17755,N_16471,N_16340);
nor U17756 (N_17756,N_16723,N_17448);
or U17757 (N_17757,N_16473,N_17015);
and U17758 (N_17758,N_16443,N_17182);
or U17759 (N_17759,N_17020,N_16543);
nor U17760 (N_17760,N_16267,N_16691);
and U17761 (N_17761,N_16527,N_17010);
nor U17762 (N_17762,N_17351,N_17441);
and U17763 (N_17763,N_16371,N_17417);
nand U17764 (N_17764,N_16939,N_16765);
nor U17765 (N_17765,N_17473,N_16560);
and U17766 (N_17766,N_16513,N_16735);
or U17767 (N_17767,N_17087,N_16662);
nand U17768 (N_17768,N_16406,N_16699);
nand U17769 (N_17769,N_16326,N_17413);
nand U17770 (N_17770,N_16475,N_16925);
or U17771 (N_17771,N_16539,N_16442);
nor U17772 (N_17772,N_16697,N_16935);
nand U17773 (N_17773,N_16903,N_17037);
or U17774 (N_17774,N_17335,N_16910);
nor U17775 (N_17775,N_17376,N_17490);
nor U17776 (N_17776,N_17317,N_16436);
xnor U17777 (N_17777,N_16461,N_16882);
nand U17778 (N_17778,N_17125,N_16818);
nand U17779 (N_17779,N_16713,N_16619);
nor U17780 (N_17780,N_16251,N_17432);
nand U17781 (N_17781,N_17216,N_17247);
xnor U17782 (N_17782,N_16877,N_16605);
or U17783 (N_17783,N_16472,N_16993);
xor U17784 (N_17784,N_16840,N_16582);
nand U17785 (N_17785,N_17186,N_17144);
nand U17786 (N_17786,N_17399,N_16847);
nand U17787 (N_17787,N_17066,N_16489);
and U17788 (N_17788,N_16843,N_16761);
nor U17789 (N_17789,N_16298,N_17107);
and U17790 (N_17790,N_16534,N_16961);
and U17791 (N_17791,N_16922,N_17377);
and U17792 (N_17792,N_16561,N_16814);
or U17793 (N_17793,N_17132,N_17465);
xnor U17794 (N_17794,N_17420,N_16404);
xor U17795 (N_17795,N_16810,N_16892);
xnor U17796 (N_17796,N_17458,N_17244);
or U17797 (N_17797,N_16559,N_16576);
nand U17798 (N_17798,N_16357,N_17022);
nand U17799 (N_17799,N_17366,N_16394);
xnor U17800 (N_17800,N_16629,N_16678);
xor U17801 (N_17801,N_16752,N_17275);
nor U17802 (N_17802,N_16755,N_17387);
nand U17803 (N_17803,N_16766,N_16813);
nor U17804 (N_17804,N_16693,N_16596);
nor U17805 (N_17805,N_16323,N_17482);
nor U17806 (N_17806,N_17393,N_17323);
or U17807 (N_17807,N_16719,N_16852);
nor U17808 (N_17808,N_16440,N_17348);
and U17809 (N_17809,N_16938,N_17312);
and U17810 (N_17810,N_16516,N_16574);
and U17811 (N_17811,N_16575,N_16998);
nor U17812 (N_17812,N_16480,N_16639);
nand U17813 (N_17813,N_17411,N_17060);
and U17814 (N_17814,N_16369,N_17477);
nand U17815 (N_17815,N_16679,N_16709);
or U17816 (N_17816,N_16664,N_16698);
nand U17817 (N_17817,N_16377,N_17164);
or U17818 (N_17818,N_16275,N_17414);
nor U17819 (N_17819,N_16337,N_16614);
nor U17820 (N_17820,N_17062,N_16899);
nor U17821 (N_17821,N_17217,N_17422);
nor U17822 (N_17822,N_16674,N_16977);
or U17823 (N_17823,N_16795,N_16399);
nand U17824 (N_17824,N_17041,N_16359);
or U17825 (N_17825,N_16885,N_17249);
nand U17826 (N_17826,N_17063,N_17330);
nand U17827 (N_17827,N_16367,N_17178);
nand U17828 (N_17828,N_17220,N_17436);
nor U17829 (N_17829,N_17472,N_16630);
nor U17830 (N_17830,N_17011,N_16677);
and U17831 (N_17831,N_16690,N_16462);
xnor U17832 (N_17832,N_17038,N_16828);
nand U17833 (N_17833,N_17279,N_16538);
or U17834 (N_17834,N_17036,N_16758);
nor U17835 (N_17835,N_16989,N_16730);
nand U17836 (N_17836,N_17209,N_16455);
and U17837 (N_17837,N_16446,N_16250);
or U17838 (N_17838,N_16768,N_16427);
nand U17839 (N_17839,N_16874,N_17008);
nand U17840 (N_17840,N_17385,N_17444);
and U17841 (N_17841,N_17045,N_16949);
xor U17842 (N_17842,N_16827,N_16468);
or U17843 (N_17843,N_16438,N_16354);
nand U17844 (N_17844,N_16449,N_17277);
xor U17845 (N_17845,N_16518,N_16434);
nand U17846 (N_17846,N_16762,N_16626);
xor U17847 (N_17847,N_16919,N_17044);
or U17848 (N_17848,N_17129,N_17409);
or U17849 (N_17849,N_17311,N_16277);
nor U17850 (N_17850,N_17274,N_16858);
nor U17851 (N_17851,N_16635,N_16936);
nand U17852 (N_17852,N_17345,N_16317);
and U17853 (N_17853,N_17390,N_16890);
or U17854 (N_17854,N_16675,N_16413);
and U17855 (N_17855,N_16310,N_17090);
nor U17856 (N_17856,N_16658,N_16994);
or U17857 (N_17857,N_17088,N_17397);
nand U17858 (N_17858,N_16409,N_17488);
or U17859 (N_17859,N_16834,N_16282);
nand U17860 (N_17860,N_17097,N_17139);
xor U17861 (N_17861,N_17142,N_16859);
xnor U17862 (N_17862,N_16700,N_16736);
or U17863 (N_17863,N_16391,N_17225);
and U17864 (N_17864,N_16912,N_17082);
nand U17865 (N_17865,N_16336,N_17419);
nor U17866 (N_17866,N_16798,N_16431);
nor U17867 (N_17867,N_17214,N_16494);
nand U17868 (N_17868,N_16537,N_16774);
nand U17869 (N_17869,N_17023,N_17219);
and U17870 (N_17870,N_16756,N_16733);
xor U17871 (N_17871,N_17485,N_17083);
nor U17872 (N_17872,N_17116,N_16529);
nor U17873 (N_17873,N_16823,N_16308);
xnor U17874 (N_17874,N_16804,N_16587);
xor U17875 (N_17875,N_16552,N_17016);
and U17876 (N_17876,N_17111,N_16447);
nand U17877 (N_17877,N_17145,N_17434);
xnor U17878 (N_17878,N_16893,N_17295);
or U17879 (N_17879,N_16982,N_17461);
and U17880 (N_17880,N_17028,N_16741);
nand U17881 (N_17881,N_16696,N_16797);
xnor U17882 (N_17882,N_17389,N_17095);
nand U17883 (N_17883,N_16663,N_16634);
or U17884 (N_17884,N_17263,N_16579);
and U17885 (N_17885,N_16660,N_16995);
and U17886 (N_17886,N_16956,N_17196);
and U17887 (N_17887,N_16717,N_16716);
xor U17888 (N_17888,N_17137,N_16701);
or U17889 (N_17889,N_16285,N_16887);
or U17890 (N_17890,N_16355,N_17228);
or U17891 (N_17891,N_16583,N_17170);
and U17892 (N_17892,N_17241,N_16826);
xor U17893 (N_17893,N_16708,N_17199);
and U17894 (N_17894,N_16681,N_16556);
and U17895 (N_17895,N_16306,N_16564);
nand U17896 (N_17896,N_16502,N_17085);
and U17897 (N_17897,N_17073,N_16562);
nor U17898 (N_17898,N_17364,N_16611);
nor U17899 (N_17899,N_16474,N_16913);
nor U17900 (N_17900,N_17123,N_17365);
nand U17901 (N_17901,N_16463,N_17464);
nor U17902 (N_17902,N_16667,N_16875);
nor U17903 (N_17903,N_16940,N_17343);
nand U17904 (N_17904,N_17175,N_17067);
xor U17905 (N_17905,N_16599,N_16458);
nor U17906 (N_17906,N_16900,N_17304);
xor U17907 (N_17907,N_16862,N_17079);
and U17908 (N_17908,N_16794,N_16524);
nand U17909 (N_17909,N_16855,N_17059);
or U17910 (N_17910,N_17056,N_17270);
and U17911 (N_17911,N_16872,N_17498);
nand U17912 (N_17912,N_16999,N_17238);
and U17913 (N_17913,N_17367,N_17299);
nand U17914 (N_17914,N_17283,N_16905);
or U17915 (N_17915,N_16358,N_16506);
and U17916 (N_17916,N_16955,N_16350);
nand U17917 (N_17917,N_17329,N_17401);
and U17918 (N_17918,N_17006,N_16773);
and U17919 (N_17919,N_16389,N_17374);
and U17920 (N_17920,N_17328,N_16334);
xnor U17921 (N_17921,N_16570,N_16435);
nor U17922 (N_17922,N_16975,N_17007);
nand U17923 (N_17923,N_17315,N_17492);
nor U17924 (N_17924,N_17223,N_16407);
nand U17925 (N_17925,N_17153,N_17155);
nand U17926 (N_17926,N_17486,N_16615);
xor U17927 (N_17927,N_17266,N_16873);
and U17928 (N_17928,N_16944,N_17165);
xnor U17929 (N_17929,N_16314,N_17115);
xor U17930 (N_17930,N_17491,N_16425);
nor U17931 (N_17931,N_16934,N_16423);
or U17932 (N_17932,N_16722,N_17340);
nand U17933 (N_17933,N_16441,N_16266);
or U17934 (N_17934,N_17313,N_17105);
xnor U17935 (N_17935,N_17371,N_17334);
or U17936 (N_17936,N_17327,N_17118);
nor U17937 (N_17937,N_17035,N_17138);
and U17938 (N_17938,N_16787,N_17446);
nor U17939 (N_17939,N_17284,N_17268);
and U17940 (N_17940,N_17438,N_17495);
nand U17941 (N_17941,N_17433,N_17257);
and U17942 (N_17942,N_17497,N_16360);
and U17943 (N_17943,N_16541,N_16846);
xor U17944 (N_17944,N_17140,N_16301);
xnor U17945 (N_17945,N_16483,N_16819);
or U17946 (N_17946,N_16375,N_16549);
xor U17947 (N_17947,N_16806,N_16747);
nand U17948 (N_17948,N_17272,N_17110);
nor U17949 (N_17949,N_17408,N_17296);
nand U17950 (N_17950,N_16784,N_16937);
nand U17951 (N_17951,N_16636,N_16972);
and U17952 (N_17952,N_17234,N_16628);
xnor U17953 (N_17953,N_17089,N_16312);
nand U17954 (N_17954,N_16720,N_16395);
and U17955 (N_17955,N_17061,N_16283);
xor U17956 (N_17956,N_17245,N_16668);
nor U17957 (N_17957,N_16764,N_17103);
nor U17958 (N_17958,N_16415,N_16383);
nor U17959 (N_17959,N_16866,N_16457);
xor U17960 (N_17960,N_16689,N_16557);
xnor U17961 (N_17961,N_17221,N_16618);
or U17962 (N_17962,N_16294,N_16591);
or U17963 (N_17963,N_16332,N_16295);
nor U17964 (N_17964,N_16835,N_17162);
or U17965 (N_17965,N_17261,N_16261);
xnor U17966 (N_17966,N_16253,N_16793);
nand U17967 (N_17967,N_16904,N_16926);
or U17968 (N_17968,N_16589,N_16374);
xnor U17969 (N_17969,N_17034,N_17341);
nand U17970 (N_17970,N_17325,N_16616);
xnor U17971 (N_17971,N_16895,N_16643);
nor U17972 (N_17972,N_16380,N_17039);
nor U17973 (N_17973,N_16953,N_16896);
and U17974 (N_17974,N_17294,N_16769);
and U17975 (N_17975,N_16888,N_16487);
nor U17976 (N_17976,N_17481,N_16894);
nor U17977 (N_17977,N_17362,N_17476);
and U17978 (N_17978,N_17050,N_17349);
nand U17979 (N_17979,N_16289,N_17084);
or U17980 (N_17980,N_16309,N_17246);
and U17981 (N_17981,N_16655,N_17242);
and U17982 (N_17982,N_16780,N_17459);
or U17983 (N_17983,N_16550,N_17210);
xor U17984 (N_17984,N_16420,N_17027);
xnor U17985 (N_17985,N_17141,N_16272);
or U17986 (N_17986,N_16428,N_17031);
nor U17987 (N_17987,N_17181,N_16863);
nor U17988 (N_17988,N_16712,N_17369);
xor U17989 (N_17989,N_16553,N_17487);
nor U17990 (N_17990,N_16844,N_17184);
nand U17991 (N_17991,N_17316,N_16987);
nand U17992 (N_17992,N_17019,N_16750);
or U17993 (N_17993,N_16686,N_17189);
xor U17994 (N_17994,N_16792,N_16418);
and U17995 (N_17995,N_16706,N_16802);
nand U17996 (N_17996,N_16745,N_16607);
nor U17997 (N_17997,N_16448,N_17202);
and U17998 (N_17998,N_16801,N_17201);
nor U17999 (N_17999,N_16400,N_17305);
or U18000 (N_18000,N_16918,N_16704);
xor U18001 (N_18001,N_16291,N_17255);
nand U18002 (N_18002,N_17240,N_16817);
nor U18003 (N_18003,N_17149,N_17208);
nor U18004 (N_18004,N_17483,N_16789);
and U18005 (N_18005,N_16445,N_16270);
nor U18006 (N_18006,N_16757,N_17104);
and U18007 (N_18007,N_16857,N_17466);
and U18008 (N_18008,N_17320,N_16477);
nand U18009 (N_18009,N_16498,N_16856);
nand U18010 (N_18010,N_17052,N_16520);
nand U18011 (N_18011,N_17025,N_16595);
or U18012 (N_18012,N_16256,N_17282);
nor U18013 (N_18013,N_16638,N_17121);
nor U18014 (N_18014,N_16416,N_16387);
nand U18015 (N_18015,N_17227,N_16344);
xnor U18016 (N_18016,N_16941,N_17258);
and U18017 (N_18017,N_16585,N_17171);
or U18018 (N_18018,N_16593,N_16327);
nand U18019 (N_18019,N_16451,N_16845);
xor U18020 (N_18020,N_16429,N_16782);
or U18021 (N_18021,N_16335,N_16632);
xnor U18022 (N_18022,N_16331,N_16726);
xor U18023 (N_18023,N_17205,N_17032);
nand U18024 (N_18024,N_16838,N_17449);
xor U18025 (N_18025,N_16821,N_16727);
and U18026 (N_18026,N_16610,N_16927);
nand U18027 (N_18027,N_16370,N_17161);
xnor U18028 (N_18028,N_16338,N_17442);
nand U18029 (N_18029,N_17319,N_16488);
and U18030 (N_18030,N_17447,N_17033);
nor U18031 (N_18031,N_16353,N_17260);
or U18032 (N_18032,N_16515,N_16278);
nor U18033 (N_18033,N_17291,N_16805);
xor U18034 (N_18034,N_17069,N_17453);
and U18035 (N_18035,N_16860,N_16300);
nand U18036 (N_18036,N_16555,N_16621);
and U18037 (N_18037,N_16914,N_16786);
nand U18038 (N_18038,N_16767,N_17375);
and U18039 (N_18039,N_16521,N_16651);
or U18040 (N_18040,N_16517,N_16623);
and U18041 (N_18041,N_17166,N_16544);
or U18042 (N_18042,N_17379,N_17289);
nor U18043 (N_18043,N_16800,N_16867);
nand U18044 (N_18044,N_16329,N_17151);
or U18045 (N_18045,N_16648,N_17306);
and U18046 (N_18046,N_16942,N_17173);
or U18047 (N_18047,N_17146,N_17457);
nand U18048 (N_18048,N_16469,N_17288);
nand U18049 (N_18049,N_16715,N_16825);
xnor U18050 (N_18050,N_16864,N_17410);
nand U18051 (N_18051,N_17102,N_17445);
xnor U18052 (N_18052,N_16931,N_17122);
nor U18053 (N_18053,N_17455,N_16412);
or U18054 (N_18054,N_16654,N_16901);
xor U18055 (N_18055,N_16507,N_16771);
nand U18056 (N_18056,N_16997,N_17321);
nand U18057 (N_18057,N_16510,N_16946);
nor U18058 (N_18058,N_16963,N_16869);
or U18059 (N_18059,N_17437,N_16362);
nor U18060 (N_18060,N_17318,N_16609);
nor U18061 (N_18061,N_17229,N_17456);
nand U18062 (N_18062,N_16346,N_16650);
nor U18063 (N_18063,N_16264,N_17152);
nor U18064 (N_18064,N_17101,N_17100);
nand U18065 (N_18065,N_16841,N_17431);
or U18066 (N_18066,N_16257,N_16973);
or U18067 (N_18067,N_16476,N_16947);
nand U18068 (N_18068,N_17243,N_16547);
and U18069 (N_18069,N_16739,N_17346);
nand U18070 (N_18070,N_16551,N_16777);
nand U18071 (N_18071,N_17493,N_16271);
or U18072 (N_18072,N_16772,N_16414);
xnor U18073 (N_18073,N_17254,N_17373);
nor U18074 (N_18074,N_17474,N_16878);
nor U18075 (N_18075,N_16373,N_17427);
and U18076 (N_18076,N_17336,N_17331);
xnor U18077 (N_18077,N_16744,N_16763);
nand U18078 (N_18078,N_16486,N_16881);
nor U18079 (N_18079,N_16842,N_16592);
xnor U18080 (N_18080,N_16509,N_17239);
nand U18081 (N_18081,N_17253,N_16902);
and U18082 (N_18082,N_17380,N_17307);
or U18083 (N_18083,N_16707,N_16325);
or U18084 (N_18084,N_16385,N_16470);
xor U18085 (N_18085,N_16627,N_17176);
or U18086 (N_18086,N_17499,N_16569);
or U18087 (N_18087,N_16983,N_17212);
xnor U18088 (N_18088,N_17185,N_16500);
nand U18089 (N_18089,N_17262,N_16379);
or U18090 (N_18090,N_16950,N_16403);
or U18091 (N_18091,N_16397,N_16911);
and U18092 (N_18092,N_16321,N_16460);
nor U18093 (N_18093,N_17256,N_16508);
xnor U18094 (N_18094,N_16588,N_16577);
nand U18095 (N_18095,N_16665,N_16839);
nand U18096 (N_18096,N_16879,N_16957);
and U18097 (N_18097,N_17190,N_17494);
or U18098 (N_18098,N_17354,N_17235);
nand U18099 (N_18099,N_16287,N_16290);
or U18100 (N_18100,N_16966,N_17231);
and U18101 (N_18101,N_16401,N_17230);
or U18102 (N_18102,N_16330,N_16439);
or U18103 (N_18103,N_16728,N_17416);
nor U18104 (N_18104,N_16365,N_16302);
and U18105 (N_18105,N_16467,N_16430);
xnor U18106 (N_18106,N_17252,N_17003);
and U18107 (N_18107,N_16421,N_17148);
xor U18108 (N_18108,N_16951,N_17029);
nor U18109 (N_18109,N_16548,N_17215);
nor U18110 (N_18110,N_16496,N_16347);
nand U18111 (N_18111,N_16907,N_17078);
or U18112 (N_18112,N_17280,N_16426);
and U18113 (N_18113,N_16273,N_16533);
or U18114 (N_18114,N_16743,N_17402);
nor U18115 (N_18115,N_17407,N_16790);
xnor U18116 (N_18116,N_16886,N_16803);
or U18117 (N_18117,N_16853,N_16381);
nor U18118 (N_18118,N_17172,N_16820);
or U18119 (N_18119,N_16339,N_16571);
nor U18120 (N_18120,N_16279,N_16608);
nor U18121 (N_18121,N_16499,N_16848);
nand U18122 (N_18122,N_16333,N_16363);
nand U18123 (N_18123,N_16410,N_16984);
and U18124 (N_18124,N_17224,N_16958);
nor U18125 (N_18125,N_16503,N_17227);
xor U18126 (N_18126,N_17116,N_17177);
nand U18127 (N_18127,N_16881,N_16271);
xnor U18128 (N_18128,N_17383,N_17004);
and U18129 (N_18129,N_17353,N_17457);
xnor U18130 (N_18130,N_16605,N_17405);
or U18131 (N_18131,N_17360,N_16966);
and U18132 (N_18132,N_16840,N_16576);
and U18133 (N_18133,N_17481,N_16779);
nor U18134 (N_18134,N_17118,N_17060);
and U18135 (N_18135,N_16788,N_17178);
and U18136 (N_18136,N_16500,N_17370);
xor U18137 (N_18137,N_16937,N_16585);
and U18138 (N_18138,N_16530,N_16933);
nor U18139 (N_18139,N_16850,N_16376);
xor U18140 (N_18140,N_16689,N_17079);
nand U18141 (N_18141,N_17378,N_16488);
xor U18142 (N_18142,N_16465,N_17421);
nand U18143 (N_18143,N_16544,N_16884);
nand U18144 (N_18144,N_16753,N_16724);
nand U18145 (N_18145,N_16877,N_16871);
xor U18146 (N_18146,N_16447,N_16636);
and U18147 (N_18147,N_17430,N_16683);
nand U18148 (N_18148,N_16566,N_16780);
nor U18149 (N_18149,N_17210,N_17143);
xor U18150 (N_18150,N_17209,N_17415);
and U18151 (N_18151,N_16571,N_16567);
xor U18152 (N_18152,N_17403,N_17498);
xnor U18153 (N_18153,N_17166,N_16341);
and U18154 (N_18154,N_17171,N_16920);
or U18155 (N_18155,N_17116,N_16537);
xor U18156 (N_18156,N_16949,N_16685);
xnor U18157 (N_18157,N_16984,N_16289);
or U18158 (N_18158,N_17302,N_16364);
nor U18159 (N_18159,N_16784,N_16360);
nand U18160 (N_18160,N_16482,N_17330);
or U18161 (N_18161,N_17344,N_17101);
and U18162 (N_18162,N_16817,N_17024);
and U18163 (N_18163,N_16371,N_17477);
nor U18164 (N_18164,N_16904,N_17329);
and U18165 (N_18165,N_16507,N_16996);
xor U18166 (N_18166,N_16541,N_16994);
or U18167 (N_18167,N_16658,N_16434);
nand U18168 (N_18168,N_16270,N_16719);
and U18169 (N_18169,N_16412,N_17292);
nor U18170 (N_18170,N_16695,N_16771);
xnor U18171 (N_18171,N_16900,N_17378);
nand U18172 (N_18172,N_17307,N_16485);
and U18173 (N_18173,N_17315,N_16288);
or U18174 (N_18174,N_17004,N_16335);
or U18175 (N_18175,N_16811,N_17383);
or U18176 (N_18176,N_17134,N_16570);
or U18177 (N_18177,N_16719,N_16444);
nand U18178 (N_18178,N_16659,N_16634);
nand U18179 (N_18179,N_16522,N_16691);
xnor U18180 (N_18180,N_17084,N_16966);
nor U18181 (N_18181,N_16785,N_16880);
nand U18182 (N_18182,N_17210,N_16882);
or U18183 (N_18183,N_16423,N_17030);
and U18184 (N_18184,N_16403,N_16417);
nor U18185 (N_18185,N_16350,N_16881);
nor U18186 (N_18186,N_16643,N_17346);
or U18187 (N_18187,N_16632,N_16550);
and U18188 (N_18188,N_17067,N_16921);
xor U18189 (N_18189,N_16264,N_16965);
nor U18190 (N_18190,N_17353,N_16789);
nor U18191 (N_18191,N_16612,N_16353);
nand U18192 (N_18192,N_17337,N_17103);
nand U18193 (N_18193,N_16328,N_16626);
nand U18194 (N_18194,N_16952,N_16726);
and U18195 (N_18195,N_16582,N_16304);
and U18196 (N_18196,N_16378,N_16602);
nor U18197 (N_18197,N_16441,N_17384);
nor U18198 (N_18198,N_16504,N_16985);
xnor U18199 (N_18199,N_16772,N_17498);
nand U18200 (N_18200,N_16328,N_16484);
xnor U18201 (N_18201,N_16303,N_17161);
xor U18202 (N_18202,N_17332,N_17394);
and U18203 (N_18203,N_16898,N_17300);
and U18204 (N_18204,N_16515,N_17280);
and U18205 (N_18205,N_16287,N_16789);
nand U18206 (N_18206,N_16475,N_16714);
xor U18207 (N_18207,N_17284,N_16326);
nand U18208 (N_18208,N_16966,N_17427);
or U18209 (N_18209,N_16600,N_17045);
or U18210 (N_18210,N_17118,N_17155);
or U18211 (N_18211,N_16598,N_17197);
and U18212 (N_18212,N_17333,N_16568);
xor U18213 (N_18213,N_17241,N_16518);
nand U18214 (N_18214,N_16358,N_17181);
xor U18215 (N_18215,N_17301,N_16626);
or U18216 (N_18216,N_16571,N_16570);
nor U18217 (N_18217,N_16352,N_17388);
nor U18218 (N_18218,N_17477,N_16411);
and U18219 (N_18219,N_17479,N_16567);
and U18220 (N_18220,N_16316,N_17007);
nor U18221 (N_18221,N_16543,N_16669);
and U18222 (N_18222,N_16510,N_16506);
nand U18223 (N_18223,N_16385,N_16821);
and U18224 (N_18224,N_16652,N_16675);
and U18225 (N_18225,N_17117,N_17456);
or U18226 (N_18226,N_16929,N_16383);
nor U18227 (N_18227,N_17414,N_17257);
xor U18228 (N_18228,N_16939,N_16397);
or U18229 (N_18229,N_17416,N_17309);
nand U18230 (N_18230,N_17194,N_17085);
or U18231 (N_18231,N_17366,N_17185);
or U18232 (N_18232,N_16949,N_16305);
nand U18233 (N_18233,N_16743,N_16836);
xnor U18234 (N_18234,N_16984,N_16383);
or U18235 (N_18235,N_16795,N_16869);
and U18236 (N_18236,N_16891,N_16271);
nand U18237 (N_18237,N_16400,N_17421);
nor U18238 (N_18238,N_17184,N_16358);
nor U18239 (N_18239,N_17341,N_16429);
or U18240 (N_18240,N_17284,N_17477);
or U18241 (N_18241,N_17006,N_17332);
nand U18242 (N_18242,N_17364,N_16524);
and U18243 (N_18243,N_16625,N_16512);
nor U18244 (N_18244,N_16681,N_17353);
and U18245 (N_18245,N_16445,N_16795);
and U18246 (N_18246,N_17066,N_17220);
nor U18247 (N_18247,N_17453,N_16502);
nand U18248 (N_18248,N_17139,N_16875);
or U18249 (N_18249,N_16523,N_16739);
xnor U18250 (N_18250,N_16301,N_17200);
and U18251 (N_18251,N_16735,N_17038);
and U18252 (N_18252,N_16605,N_17428);
nor U18253 (N_18253,N_17264,N_17273);
nor U18254 (N_18254,N_16745,N_17451);
nor U18255 (N_18255,N_17229,N_17007);
nor U18256 (N_18256,N_16667,N_16937);
nor U18257 (N_18257,N_17120,N_16899);
xnor U18258 (N_18258,N_16664,N_16952);
or U18259 (N_18259,N_17382,N_16683);
nor U18260 (N_18260,N_16382,N_16288);
nand U18261 (N_18261,N_16649,N_16366);
nand U18262 (N_18262,N_16416,N_16399);
nand U18263 (N_18263,N_16822,N_16480);
nor U18264 (N_18264,N_17180,N_17273);
nor U18265 (N_18265,N_16644,N_16532);
nor U18266 (N_18266,N_17017,N_17473);
and U18267 (N_18267,N_17345,N_16356);
or U18268 (N_18268,N_17489,N_16503);
nand U18269 (N_18269,N_17274,N_16285);
xor U18270 (N_18270,N_16620,N_17142);
nand U18271 (N_18271,N_16542,N_16727);
nor U18272 (N_18272,N_16883,N_17057);
nor U18273 (N_18273,N_16493,N_17484);
xnor U18274 (N_18274,N_16504,N_16718);
nor U18275 (N_18275,N_17339,N_16757);
nor U18276 (N_18276,N_16896,N_16434);
nor U18277 (N_18277,N_16831,N_16716);
or U18278 (N_18278,N_17265,N_16513);
xor U18279 (N_18279,N_17156,N_17461);
and U18280 (N_18280,N_16298,N_16734);
xor U18281 (N_18281,N_16859,N_16470);
and U18282 (N_18282,N_17367,N_16455);
xnor U18283 (N_18283,N_16410,N_17335);
nand U18284 (N_18284,N_16614,N_17467);
xnor U18285 (N_18285,N_16948,N_16491);
and U18286 (N_18286,N_16492,N_16878);
xnor U18287 (N_18287,N_17069,N_17468);
nand U18288 (N_18288,N_16255,N_16758);
nor U18289 (N_18289,N_16404,N_17075);
nor U18290 (N_18290,N_17445,N_16985);
and U18291 (N_18291,N_16901,N_17384);
xnor U18292 (N_18292,N_17160,N_16878);
nor U18293 (N_18293,N_16471,N_16456);
or U18294 (N_18294,N_16507,N_17407);
and U18295 (N_18295,N_17416,N_17458);
xor U18296 (N_18296,N_16891,N_17190);
and U18297 (N_18297,N_16715,N_16964);
nor U18298 (N_18298,N_17105,N_16880);
xnor U18299 (N_18299,N_17264,N_17023);
or U18300 (N_18300,N_16904,N_16968);
and U18301 (N_18301,N_17217,N_17499);
or U18302 (N_18302,N_16945,N_16582);
and U18303 (N_18303,N_16588,N_16391);
nor U18304 (N_18304,N_16571,N_16948);
xnor U18305 (N_18305,N_17046,N_16744);
and U18306 (N_18306,N_16608,N_17491);
nand U18307 (N_18307,N_16317,N_16733);
nor U18308 (N_18308,N_16968,N_17073);
xor U18309 (N_18309,N_16772,N_16300);
xnor U18310 (N_18310,N_16723,N_16386);
and U18311 (N_18311,N_16551,N_16553);
xnor U18312 (N_18312,N_16263,N_16850);
nor U18313 (N_18313,N_17420,N_16990);
nand U18314 (N_18314,N_16396,N_16981);
nor U18315 (N_18315,N_16588,N_16656);
nor U18316 (N_18316,N_16868,N_16587);
nand U18317 (N_18317,N_16318,N_17210);
nor U18318 (N_18318,N_17394,N_17287);
nand U18319 (N_18319,N_17318,N_16263);
and U18320 (N_18320,N_17082,N_16712);
nand U18321 (N_18321,N_16736,N_16277);
xor U18322 (N_18322,N_16725,N_16898);
nor U18323 (N_18323,N_16853,N_16750);
and U18324 (N_18324,N_16655,N_17368);
nand U18325 (N_18325,N_16661,N_16375);
nand U18326 (N_18326,N_16449,N_17316);
nor U18327 (N_18327,N_16364,N_16253);
nor U18328 (N_18328,N_16260,N_16858);
nand U18329 (N_18329,N_17190,N_16865);
xor U18330 (N_18330,N_17220,N_16920);
xnor U18331 (N_18331,N_17264,N_17050);
and U18332 (N_18332,N_17029,N_17239);
and U18333 (N_18333,N_16859,N_16707);
and U18334 (N_18334,N_17149,N_16973);
xor U18335 (N_18335,N_17191,N_16419);
or U18336 (N_18336,N_16680,N_16809);
nand U18337 (N_18337,N_16887,N_16566);
or U18338 (N_18338,N_17245,N_16955);
nand U18339 (N_18339,N_17471,N_16503);
and U18340 (N_18340,N_16875,N_16640);
and U18341 (N_18341,N_16700,N_16885);
or U18342 (N_18342,N_16760,N_17065);
or U18343 (N_18343,N_16689,N_17374);
nand U18344 (N_18344,N_16935,N_17245);
xor U18345 (N_18345,N_17176,N_17001);
nor U18346 (N_18346,N_17465,N_16423);
or U18347 (N_18347,N_16808,N_17012);
nor U18348 (N_18348,N_16951,N_16553);
nor U18349 (N_18349,N_16521,N_16696);
nand U18350 (N_18350,N_16811,N_17461);
or U18351 (N_18351,N_16282,N_17078);
or U18352 (N_18352,N_17253,N_17010);
xor U18353 (N_18353,N_16868,N_17277);
or U18354 (N_18354,N_16325,N_16653);
nor U18355 (N_18355,N_17092,N_16688);
nand U18356 (N_18356,N_16347,N_16552);
or U18357 (N_18357,N_16251,N_16844);
xnor U18358 (N_18358,N_17287,N_16318);
or U18359 (N_18359,N_16743,N_16768);
xnor U18360 (N_18360,N_16718,N_17234);
nor U18361 (N_18361,N_17260,N_16617);
xnor U18362 (N_18362,N_17489,N_16838);
or U18363 (N_18363,N_16980,N_16506);
nand U18364 (N_18364,N_16535,N_17278);
and U18365 (N_18365,N_16635,N_16269);
xor U18366 (N_18366,N_16250,N_16603);
xor U18367 (N_18367,N_17360,N_17375);
nand U18368 (N_18368,N_16602,N_17432);
nor U18369 (N_18369,N_16453,N_16876);
and U18370 (N_18370,N_16255,N_17495);
xnor U18371 (N_18371,N_17088,N_16848);
nor U18372 (N_18372,N_16821,N_16551);
or U18373 (N_18373,N_16612,N_17443);
xnor U18374 (N_18374,N_16735,N_16439);
nor U18375 (N_18375,N_16290,N_17080);
nor U18376 (N_18376,N_17118,N_16293);
xor U18377 (N_18377,N_17166,N_17245);
nor U18378 (N_18378,N_16935,N_17171);
or U18379 (N_18379,N_16921,N_16285);
nor U18380 (N_18380,N_16479,N_17444);
xor U18381 (N_18381,N_16892,N_16785);
nor U18382 (N_18382,N_17266,N_17420);
xor U18383 (N_18383,N_17223,N_17332);
or U18384 (N_18384,N_16706,N_16366);
or U18385 (N_18385,N_17122,N_16710);
and U18386 (N_18386,N_17066,N_17030);
nand U18387 (N_18387,N_16951,N_16887);
nand U18388 (N_18388,N_16328,N_16695);
nor U18389 (N_18389,N_16613,N_16262);
nor U18390 (N_18390,N_17497,N_16904);
xnor U18391 (N_18391,N_16619,N_16327);
nor U18392 (N_18392,N_17230,N_16702);
and U18393 (N_18393,N_17255,N_17115);
nor U18394 (N_18394,N_17357,N_16480);
xnor U18395 (N_18395,N_16470,N_16635);
and U18396 (N_18396,N_17364,N_16490);
nor U18397 (N_18397,N_16300,N_16380);
xor U18398 (N_18398,N_16823,N_16905);
and U18399 (N_18399,N_16286,N_16488);
nand U18400 (N_18400,N_16387,N_16852);
nand U18401 (N_18401,N_16987,N_17334);
and U18402 (N_18402,N_16355,N_16506);
nand U18403 (N_18403,N_16812,N_17192);
xor U18404 (N_18404,N_16502,N_16769);
and U18405 (N_18405,N_16959,N_16893);
nor U18406 (N_18406,N_17469,N_16550);
nor U18407 (N_18407,N_16625,N_17388);
and U18408 (N_18408,N_16891,N_16634);
nor U18409 (N_18409,N_17283,N_16699);
nor U18410 (N_18410,N_17067,N_16711);
or U18411 (N_18411,N_16636,N_17005);
xnor U18412 (N_18412,N_16306,N_16302);
nor U18413 (N_18413,N_17213,N_17485);
and U18414 (N_18414,N_16660,N_16436);
xnor U18415 (N_18415,N_17275,N_16988);
and U18416 (N_18416,N_16923,N_16950);
nor U18417 (N_18417,N_17415,N_17224);
or U18418 (N_18418,N_17492,N_16659);
and U18419 (N_18419,N_16676,N_17129);
nor U18420 (N_18420,N_16384,N_16649);
nand U18421 (N_18421,N_17102,N_16394);
xnor U18422 (N_18422,N_16601,N_17101);
nand U18423 (N_18423,N_17130,N_16863);
xor U18424 (N_18424,N_17088,N_16619);
xnor U18425 (N_18425,N_17278,N_17016);
and U18426 (N_18426,N_16388,N_17468);
nor U18427 (N_18427,N_16475,N_16486);
and U18428 (N_18428,N_17499,N_16693);
or U18429 (N_18429,N_17012,N_16827);
nand U18430 (N_18430,N_16891,N_16960);
nand U18431 (N_18431,N_17307,N_16846);
nor U18432 (N_18432,N_17228,N_17291);
xnor U18433 (N_18433,N_16878,N_16278);
and U18434 (N_18434,N_17066,N_17127);
nand U18435 (N_18435,N_16525,N_16955);
xor U18436 (N_18436,N_16354,N_16521);
nand U18437 (N_18437,N_16887,N_17384);
xor U18438 (N_18438,N_16797,N_16779);
nand U18439 (N_18439,N_16611,N_17315);
or U18440 (N_18440,N_16331,N_17216);
or U18441 (N_18441,N_16284,N_16380);
nor U18442 (N_18442,N_16954,N_17107);
nor U18443 (N_18443,N_16662,N_16677);
nor U18444 (N_18444,N_16767,N_16392);
or U18445 (N_18445,N_16610,N_17065);
nor U18446 (N_18446,N_16547,N_17140);
xor U18447 (N_18447,N_17241,N_16783);
nand U18448 (N_18448,N_16786,N_16984);
nor U18449 (N_18449,N_16588,N_16423);
or U18450 (N_18450,N_16981,N_17173);
or U18451 (N_18451,N_16442,N_17130);
xnor U18452 (N_18452,N_16938,N_16635);
or U18453 (N_18453,N_17499,N_17449);
and U18454 (N_18454,N_17310,N_17239);
nand U18455 (N_18455,N_17452,N_16326);
xnor U18456 (N_18456,N_17242,N_17448);
or U18457 (N_18457,N_16291,N_16305);
xor U18458 (N_18458,N_16304,N_16414);
nor U18459 (N_18459,N_16838,N_17477);
or U18460 (N_18460,N_17100,N_16756);
and U18461 (N_18461,N_16949,N_17143);
xor U18462 (N_18462,N_16747,N_17426);
or U18463 (N_18463,N_17465,N_16311);
nand U18464 (N_18464,N_17289,N_17250);
xnor U18465 (N_18465,N_16878,N_16426);
and U18466 (N_18466,N_16439,N_16564);
xnor U18467 (N_18467,N_17498,N_16722);
xor U18468 (N_18468,N_16368,N_16375);
nand U18469 (N_18469,N_16908,N_16337);
nor U18470 (N_18470,N_17104,N_16609);
xnor U18471 (N_18471,N_16429,N_17414);
nor U18472 (N_18472,N_16723,N_17221);
xor U18473 (N_18473,N_16908,N_17461);
xnor U18474 (N_18474,N_17125,N_16551);
nand U18475 (N_18475,N_16918,N_17397);
and U18476 (N_18476,N_16769,N_16908);
and U18477 (N_18477,N_16722,N_16287);
and U18478 (N_18478,N_16434,N_16344);
nand U18479 (N_18479,N_16584,N_16379);
or U18480 (N_18480,N_17069,N_17257);
and U18481 (N_18481,N_16848,N_16860);
nor U18482 (N_18482,N_16878,N_16664);
nor U18483 (N_18483,N_17003,N_17331);
or U18484 (N_18484,N_16329,N_16323);
xor U18485 (N_18485,N_16978,N_16790);
or U18486 (N_18486,N_16823,N_17442);
and U18487 (N_18487,N_16720,N_16542);
nand U18488 (N_18488,N_17000,N_16982);
xnor U18489 (N_18489,N_16965,N_16829);
or U18490 (N_18490,N_16782,N_16876);
xnor U18491 (N_18491,N_17278,N_16412);
xnor U18492 (N_18492,N_17214,N_17200);
or U18493 (N_18493,N_16508,N_16687);
and U18494 (N_18494,N_17230,N_16736);
or U18495 (N_18495,N_16261,N_16732);
nand U18496 (N_18496,N_16803,N_17239);
xnor U18497 (N_18497,N_17416,N_16837);
or U18498 (N_18498,N_16820,N_16920);
xor U18499 (N_18499,N_17375,N_16965);
nand U18500 (N_18500,N_17456,N_16312);
and U18501 (N_18501,N_16891,N_16997);
xnor U18502 (N_18502,N_17161,N_16628);
nand U18503 (N_18503,N_16906,N_17210);
nor U18504 (N_18504,N_17483,N_17046);
or U18505 (N_18505,N_17420,N_16626);
or U18506 (N_18506,N_17468,N_17253);
nor U18507 (N_18507,N_16887,N_16266);
nand U18508 (N_18508,N_17401,N_17246);
xnor U18509 (N_18509,N_17051,N_17312);
and U18510 (N_18510,N_16954,N_16648);
nor U18511 (N_18511,N_16808,N_17410);
and U18512 (N_18512,N_16730,N_16497);
and U18513 (N_18513,N_16825,N_17154);
nor U18514 (N_18514,N_16719,N_16836);
xor U18515 (N_18515,N_17378,N_17330);
xor U18516 (N_18516,N_17206,N_16822);
nand U18517 (N_18517,N_16322,N_17387);
nor U18518 (N_18518,N_16669,N_17412);
or U18519 (N_18519,N_16895,N_16347);
and U18520 (N_18520,N_17030,N_17475);
nand U18521 (N_18521,N_16898,N_16930);
or U18522 (N_18522,N_17333,N_17495);
nand U18523 (N_18523,N_17451,N_16800);
nor U18524 (N_18524,N_16998,N_16702);
nand U18525 (N_18525,N_17116,N_16521);
nor U18526 (N_18526,N_16460,N_16470);
and U18527 (N_18527,N_16408,N_17168);
nor U18528 (N_18528,N_16327,N_16847);
xor U18529 (N_18529,N_17303,N_17141);
or U18530 (N_18530,N_16354,N_16933);
and U18531 (N_18531,N_16969,N_16253);
or U18532 (N_18532,N_16913,N_17431);
nand U18533 (N_18533,N_16592,N_17487);
and U18534 (N_18534,N_16497,N_17424);
or U18535 (N_18535,N_16335,N_17092);
or U18536 (N_18536,N_16310,N_16570);
nor U18537 (N_18537,N_16277,N_16404);
nor U18538 (N_18538,N_16830,N_16514);
nand U18539 (N_18539,N_16291,N_16858);
or U18540 (N_18540,N_16281,N_17159);
xnor U18541 (N_18541,N_16487,N_17146);
nand U18542 (N_18542,N_17120,N_17269);
xnor U18543 (N_18543,N_17380,N_16497);
nand U18544 (N_18544,N_17122,N_16457);
and U18545 (N_18545,N_17442,N_16502);
nand U18546 (N_18546,N_16284,N_16630);
and U18547 (N_18547,N_16312,N_16395);
nor U18548 (N_18548,N_17340,N_17003);
xnor U18549 (N_18549,N_16574,N_17108);
nor U18550 (N_18550,N_16298,N_17408);
nor U18551 (N_18551,N_16650,N_17052);
xor U18552 (N_18552,N_16778,N_17159);
nand U18553 (N_18553,N_16544,N_17427);
xnor U18554 (N_18554,N_17433,N_17135);
or U18555 (N_18555,N_17399,N_17116);
nor U18556 (N_18556,N_16442,N_16627);
nand U18557 (N_18557,N_16469,N_16972);
or U18558 (N_18558,N_17400,N_17043);
or U18559 (N_18559,N_16369,N_16748);
or U18560 (N_18560,N_17051,N_16893);
nand U18561 (N_18561,N_16966,N_17155);
nand U18562 (N_18562,N_17200,N_16700);
or U18563 (N_18563,N_17438,N_17201);
xor U18564 (N_18564,N_16546,N_17224);
or U18565 (N_18565,N_16288,N_16265);
nor U18566 (N_18566,N_16921,N_16329);
or U18567 (N_18567,N_16615,N_16547);
nor U18568 (N_18568,N_16384,N_17198);
nand U18569 (N_18569,N_16808,N_17191);
and U18570 (N_18570,N_16595,N_16279);
nor U18571 (N_18571,N_17407,N_16730);
or U18572 (N_18572,N_16425,N_16976);
and U18573 (N_18573,N_16926,N_16534);
nor U18574 (N_18574,N_16951,N_17272);
or U18575 (N_18575,N_16300,N_16454);
or U18576 (N_18576,N_16336,N_16717);
xor U18577 (N_18577,N_16706,N_16939);
xnor U18578 (N_18578,N_16652,N_16950);
nor U18579 (N_18579,N_16997,N_16950);
nor U18580 (N_18580,N_16701,N_16743);
nor U18581 (N_18581,N_17389,N_16558);
nand U18582 (N_18582,N_17362,N_17211);
xnor U18583 (N_18583,N_16848,N_17462);
nor U18584 (N_18584,N_17092,N_16359);
xor U18585 (N_18585,N_17495,N_16377);
and U18586 (N_18586,N_16912,N_17409);
and U18587 (N_18587,N_17051,N_16952);
and U18588 (N_18588,N_16476,N_17091);
nand U18589 (N_18589,N_16319,N_16314);
nand U18590 (N_18590,N_17447,N_17110);
nand U18591 (N_18591,N_16354,N_16526);
nor U18592 (N_18592,N_16993,N_17420);
and U18593 (N_18593,N_16564,N_17085);
nor U18594 (N_18594,N_17446,N_16516);
nand U18595 (N_18595,N_16940,N_17292);
or U18596 (N_18596,N_16750,N_17459);
nor U18597 (N_18597,N_16570,N_17095);
nand U18598 (N_18598,N_16795,N_16461);
and U18599 (N_18599,N_17165,N_16824);
nor U18600 (N_18600,N_16696,N_16295);
or U18601 (N_18601,N_16758,N_17006);
or U18602 (N_18602,N_17376,N_17236);
nor U18603 (N_18603,N_16290,N_17152);
nand U18604 (N_18604,N_16725,N_16743);
nor U18605 (N_18605,N_16682,N_17304);
xor U18606 (N_18606,N_17412,N_16489);
or U18607 (N_18607,N_17420,N_16444);
and U18608 (N_18608,N_17270,N_17311);
xor U18609 (N_18609,N_16730,N_17486);
and U18610 (N_18610,N_17083,N_16852);
nor U18611 (N_18611,N_16539,N_16411);
or U18612 (N_18612,N_17139,N_16910);
nand U18613 (N_18613,N_16617,N_16640);
nor U18614 (N_18614,N_17496,N_16593);
nor U18615 (N_18615,N_16628,N_17346);
and U18616 (N_18616,N_16704,N_17284);
nor U18617 (N_18617,N_17259,N_16338);
nor U18618 (N_18618,N_16274,N_17123);
and U18619 (N_18619,N_17020,N_17175);
and U18620 (N_18620,N_17174,N_16544);
or U18621 (N_18621,N_16859,N_17363);
or U18622 (N_18622,N_16611,N_16273);
nor U18623 (N_18623,N_16411,N_16305);
and U18624 (N_18624,N_16889,N_16408);
xor U18625 (N_18625,N_17120,N_16603);
nor U18626 (N_18626,N_17375,N_17185);
and U18627 (N_18627,N_16781,N_16828);
nor U18628 (N_18628,N_16957,N_17431);
and U18629 (N_18629,N_16761,N_16937);
or U18630 (N_18630,N_17480,N_16348);
or U18631 (N_18631,N_17074,N_17383);
and U18632 (N_18632,N_16680,N_16312);
and U18633 (N_18633,N_16317,N_17112);
and U18634 (N_18634,N_16340,N_16503);
xnor U18635 (N_18635,N_16704,N_17030);
or U18636 (N_18636,N_16917,N_16357);
xor U18637 (N_18637,N_16438,N_17332);
or U18638 (N_18638,N_16639,N_16770);
xnor U18639 (N_18639,N_16402,N_16729);
nand U18640 (N_18640,N_17413,N_16572);
nor U18641 (N_18641,N_16585,N_16641);
or U18642 (N_18642,N_16967,N_17090);
nand U18643 (N_18643,N_16446,N_17160);
and U18644 (N_18644,N_16994,N_17132);
xnor U18645 (N_18645,N_16398,N_17249);
and U18646 (N_18646,N_16932,N_16470);
xor U18647 (N_18647,N_17162,N_16978);
or U18648 (N_18648,N_16668,N_17330);
nor U18649 (N_18649,N_17377,N_17126);
or U18650 (N_18650,N_16252,N_16462);
nand U18651 (N_18651,N_16909,N_17016);
or U18652 (N_18652,N_16737,N_17385);
nand U18653 (N_18653,N_17267,N_17359);
nand U18654 (N_18654,N_16495,N_16763);
or U18655 (N_18655,N_16282,N_17168);
or U18656 (N_18656,N_16968,N_16975);
nor U18657 (N_18657,N_17257,N_17223);
or U18658 (N_18658,N_16888,N_17158);
nand U18659 (N_18659,N_17188,N_16745);
nand U18660 (N_18660,N_17250,N_16648);
nand U18661 (N_18661,N_17133,N_17467);
xor U18662 (N_18662,N_17147,N_16653);
and U18663 (N_18663,N_17023,N_17155);
nand U18664 (N_18664,N_16664,N_16286);
nand U18665 (N_18665,N_16272,N_17274);
or U18666 (N_18666,N_16765,N_16893);
or U18667 (N_18667,N_17101,N_16295);
nor U18668 (N_18668,N_16257,N_17006);
and U18669 (N_18669,N_16753,N_16666);
or U18670 (N_18670,N_17326,N_16456);
nand U18671 (N_18671,N_16509,N_16865);
nand U18672 (N_18672,N_16426,N_17048);
nor U18673 (N_18673,N_16943,N_16702);
xnor U18674 (N_18674,N_17285,N_16825);
and U18675 (N_18675,N_16989,N_16654);
nand U18676 (N_18676,N_17344,N_16430);
and U18677 (N_18677,N_16939,N_16895);
and U18678 (N_18678,N_16697,N_16806);
xnor U18679 (N_18679,N_16984,N_17450);
or U18680 (N_18680,N_16505,N_17293);
nand U18681 (N_18681,N_16850,N_16434);
xnor U18682 (N_18682,N_17303,N_17206);
or U18683 (N_18683,N_16951,N_17382);
nor U18684 (N_18684,N_17110,N_16307);
nand U18685 (N_18685,N_17085,N_17498);
xnor U18686 (N_18686,N_17353,N_16856);
or U18687 (N_18687,N_17392,N_17445);
or U18688 (N_18688,N_16546,N_17034);
nor U18689 (N_18689,N_17144,N_16902);
and U18690 (N_18690,N_16580,N_17217);
xnor U18691 (N_18691,N_17246,N_17353);
xor U18692 (N_18692,N_17270,N_17447);
nand U18693 (N_18693,N_16457,N_17207);
or U18694 (N_18694,N_16311,N_16747);
xor U18695 (N_18695,N_16777,N_17327);
nand U18696 (N_18696,N_17093,N_16333);
xnor U18697 (N_18697,N_16933,N_17467);
nor U18698 (N_18698,N_16754,N_16803);
and U18699 (N_18699,N_16259,N_16674);
and U18700 (N_18700,N_16675,N_17118);
or U18701 (N_18701,N_17426,N_17031);
xor U18702 (N_18702,N_16886,N_17455);
and U18703 (N_18703,N_16543,N_17240);
nand U18704 (N_18704,N_17349,N_16672);
nor U18705 (N_18705,N_16840,N_16341);
nand U18706 (N_18706,N_16947,N_17270);
xor U18707 (N_18707,N_16802,N_16715);
nand U18708 (N_18708,N_16355,N_16298);
and U18709 (N_18709,N_17279,N_17379);
nand U18710 (N_18710,N_17114,N_16498);
xor U18711 (N_18711,N_16792,N_17194);
or U18712 (N_18712,N_16366,N_16661);
xor U18713 (N_18713,N_16976,N_16424);
nor U18714 (N_18714,N_16587,N_16490);
and U18715 (N_18715,N_16498,N_17182);
nand U18716 (N_18716,N_16669,N_16592);
nor U18717 (N_18717,N_16413,N_17161);
nand U18718 (N_18718,N_16800,N_17187);
nand U18719 (N_18719,N_16375,N_17109);
and U18720 (N_18720,N_16388,N_16328);
or U18721 (N_18721,N_17306,N_17390);
and U18722 (N_18722,N_17073,N_17183);
or U18723 (N_18723,N_17389,N_17034);
and U18724 (N_18724,N_17408,N_17456);
nand U18725 (N_18725,N_16760,N_16872);
nand U18726 (N_18726,N_16786,N_17033);
nor U18727 (N_18727,N_17482,N_17018);
or U18728 (N_18728,N_16756,N_16255);
and U18729 (N_18729,N_16663,N_16385);
and U18730 (N_18730,N_17258,N_16349);
xnor U18731 (N_18731,N_16755,N_16863);
nand U18732 (N_18732,N_16663,N_17249);
nor U18733 (N_18733,N_16531,N_17389);
nor U18734 (N_18734,N_16404,N_16961);
xnor U18735 (N_18735,N_17095,N_16339);
and U18736 (N_18736,N_17123,N_17196);
nand U18737 (N_18737,N_17274,N_17471);
and U18738 (N_18738,N_16960,N_17355);
nand U18739 (N_18739,N_16465,N_17307);
nand U18740 (N_18740,N_16809,N_17114);
or U18741 (N_18741,N_16750,N_16310);
or U18742 (N_18742,N_16687,N_17140);
or U18743 (N_18743,N_16947,N_16507);
nand U18744 (N_18744,N_17035,N_17358);
nand U18745 (N_18745,N_17149,N_16744);
nand U18746 (N_18746,N_16921,N_16512);
xnor U18747 (N_18747,N_16913,N_17242);
nand U18748 (N_18748,N_16854,N_16778);
xor U18749 (N_18749,N_17345,N_16312);
xor U18750 (N_18750,N_17915,N_17822);
or U18751 (N_18751,N_17987,N_18498);
nor U18752 (N_18752,N_18160,N_18549);
nand U18753 (N_18753,N_17639,N_18203);
nor U18754 (N_18754,N_17790,N_18178);
nor U18755 (N_18755,N_18249,N_17868);
and U18756 (N_18756,N_17894,N_18106);
and U18757 (N_18757,N_18024,N_18431);
or U18758 (N_18758,N_17953,N_18334);
nand U18759 (N_18759,N_18643,N_18046);
and U18760 (N_18760,N_17957,N_18580);
nor U18761 (N_18761,N_17964,N_17620);
xnor U18762 (N_18762,N_17540,N_18468);
nand U18763 (N_18763,N_18281,N_18522);
and U18764 (N_18764,N_17851,N_17580);
nand U18765 (N_18765,N_18328,N_18098);
and U18766 (N_18766,N_18224,N_17856);
nand U18767 (N_18767,N_18442,N_17763);
or U18768 (N_18768,N_18338,N_17810);
xor U18769 (N_18769,N_18245,N_18736);
or U18770 (N_18770,N_18672,N_17944);
nor U18771 (N_18771,N_18086,N_18258);
or U18772 (N_18772,N_18344,N_18256);
xor U18773 (N_18773,N_18227,N_18354);
xor U18774 (N_18774,N_17959,N_17507);
nand U18775 (N_18775,N_18676,N_18638);
xnor U18776 (N_18776,N_18564,N_17603);
or U18777 (N_18777,N_18018,N_18108);
xor U18778 (N_18778,N_18219,N_17629);
and U18779 (N_18779,N_17626,N_18659);
nand U18780 (N_18780,N_18165,N_17729);
xor U18781 (N_18781,N_18282,N_18154);
nor U18782 (N_18782,N_17656,N_17889);
and U18783 (N_18783,N_18409,N_18147);
and U18784 (N_18784,N_17897,N_18292);
and U18785 (N_18785,N_17947,N_17760);
nand U18786 (N_18786,N_18254,N_17885);
and U18787 (N_18787,N_18162,N_17689);
nor U18788 (N_18788,N_18398,N_17609);
and U18789 (N_18789,N_18402,N_18632);
nand U18790 (N_18790,N_17756,N_18126);
nand U18791 (N_18791,N_18304,N_18131);
or U18792 (N_18792,N_17844,N_18007);
and U18793 (N_18793,N_17651,N_17634);
and U18794 (N_18794,N_18566,N_18230);
nand U18795 (N_18795,N_18301,N_17981);
nand U18796 (N_18796,N_18235,N_18671);
or U18797 (N_18797,N_17666,N_18050);
nor U18798 (N_18798,N_17853,N_17882);
nor U18799 (N_18799,N_18691,N_18090);
nand U18800 (N_18800,N_17695,N_18618);
and U18801 (N_18801,N_18565,N_17751);
nor U18802 (N_18802,N_17727,N_18006);
and U18803 (N_18803,N_18319,N_18192);
or U18804 (N_18804,N_17646,N_18403);
nand U18805 (N_18805,N_18367,N_18146);
or U18806 (N_18806,N_18078,N_18323);
or U18807 (N_18807,N_17510,N_18217);
nor U18808 (N_18808,N_18137,N_17595);
and U18809 (N_18809,N_18302,N_17614);
nor U18810 (N_18810,N_17734,N_18547);
nor U18811 (N_18811,N_18183,N_18275);
and U18812 (N_18812,N_18239,N_17631);
xor U18813 (N_18813,N_17655,N_18128);
nand U18814 (N_18814,N_17584,N_17876);
xnor U18815 (N_18815,N_18746,N_18038);
and U18816 (N_18816,N_18163,N_17546);
or U18817 (N_18817,N_18170,N_18438);
xor U18818 (N_18818,N_18125,N_18175);
nand U18819 (N_18819,N_17926,N_17950);
or U18820 (N_18820,N_18336,N_18654);
or U18821 (N_18821,N_18148,N_18470);
nand U18822 (N_18822,N_18729,N_18238);
or U18823 (N_18823,N_18464,N_18532);
nand U18824 (N_18824,N_17969,N_17770);
or U18825 (N_18825,N_17526,N_17578);
or U18826 (N_18826,N_17663,N_18042);
or U18827 (N_18827,N_17705,N_18507);
nand U18828 (N_18828,N_18360,N_18544);
xor U18829 (N_18829,N_18020,N_18513);
nand U18830 (N_18830,N_17662,N_17766);
xnor U18831 (N_18831,N_17815,N_17949);
xor U18832 (N_18832,N_18538,N_18340);
and U18833 (N_18833,N_18359,N_18646);
and U18834 (N_18834,N_17768,N_18317);
nand U18835 (N_18835,N_18493,N_17874);
xor U18836 (N_18836,N_18491,N_18429);
nor U18837 (N_18837,N_17877,N_18705);
and U18838 (N_18838,N_18112,N_18697);
xnor U18839 (N_18839,N_18714,N_17862);
xnor U18840 (N_18840,N_18114,N_17759);
or U18841 (N_18841,N_18415,N_18517);
nand U18842 (N_18842,N_18229,N_18185);
xor U18843 (N_18843,N_17956,N_17861);
or U18844 (N_18844,N_17587,N_18719);
nor U18845 (N_18845,N_17625,N_17670);
nor U18846 (N_18846,N_17963,N_18121);
xor U18847 (N_18847,N_18297,N_17749);
and U18848 (N_18848,N_18370,N_18337);
nand U18849 (N_18849,N_17523,N_18169);
xor U18850 (N_18850,N_18315,N_17958);
nand U18851 (N_18851,N_17916,N_17652);
xor U18852 (N_18852,N_17781,N_18063);
nand U18853 (N_18853,N_18631,N_18070);
nand U18854 (N_18854,N_18716,N_17665);
nor U18855 (N_18855,N_17679,N_18629);
and U18856 (N_18856,N_18695,N_18324);
nor U18857 (N_18857,N_17518,N_18561);
nand U18858 (N_18858,N_18043,N_17994);
xor U18859 (N_18859,N_18193,N_18035);
or U18860 (N_18860,N_17521,N_17955);
nor U18861 (N_18861,N_18383,N_18504);
or U18862 (N_18862,N_18158,N_17951);
xor U18863 (N_18863,N_18142,N_18586);
xnor U18864 (N_18864,N_17736,N_17677);
or U18865 (N_18865,N_17921,N_17528);
and U18866 (N_18866,N_18543,N_18309);
or U18867 (N_18867,N_18333,N_18542);
or U18868 (N_18868,N_17989,N_18529);
xnor U18869 (N_18869,N_18712,N_17701);
nand U18870 (N_18870,N_18735,N_17813);
or U18871 (N_18871,N_17560,N_18311);
xor U18872 (N_18872,N_17683,N_18263);
or U18873 (N_18873,N_17806,N_17754);
nor U18874 (N_18874,N_17505,N_17924);
and U18875 (N_18875,N_18377,N_17986);
nand U18876 (N_18876,N_17574,N_17611);
nor U18877 (N_18877,N_17912,N_18553);
nand U18878 (N_18878,N_17918,N_18366);
or U18879 (N_18879,N_18450,N_18428);
nor U18880 (N_18880,N_18068,N_17500);
or U18881 (N_18881,N_18420,N_17616);
xor U18882 (N_18882,N_17588,N_18184);
nor U18883 (N_18883,N_17865,N_18584);
nand U18884 (N_18884,N_18573,N_17745);
and U18885 (N_18885,N_18049,N_18257);
nor U18886 (N_18886,N_18589,N_17961);
nor U18887 (N_18887,N_17910,N_18702);
nor U18888 (N_18888,N_18077,N_17901);
xor U18889 (N_18889,N_17791,N_18312);
xnor U18890 (N_18890,N_18482,N_18639);
xor U18891 (N_18891,N_18685,N_17577);
nand U18892 (N_18892,N_17693,N_17875);
nor U18893 (N_18893,N_18437,N_18467);
xnor U18894 (N_18894,N_18373,N_17906);
or U18895 (N_18895,N_18053,N_17890);
xnor U18896 (N_18896,N_17798,N_17575);
nor U18897 (N_18897,N_18644,N_18687);
nor U18898 (N_18898,N_18277,N_17511);
and U18899 (N_18899,N_17632,N_17896);
nand U18900 (N_18900,N_18455,N_18039);
nor U18901 (N_18901,N_18195,N_18447);
xnor U18902 (N_18902,N_17769,N_17873);
nor U18903 (N_18903,N_18255,N_18594);
nor U18904 (N_18904,N_18711,N_18481);
nor U18905 (N_18905,N_17681,N_18250);
nor U18906 (N_18906,N_18385,N_17606);
xnor U18907 (N_18907,N_18358,N_18454);
nand U18908 (N_18908,N_18088,N_17506);
nor U18909 (N_18909,N_17817,N_17517);
nand U18910 (N_18910,N_17613,N_18197);
and U18911 (N_18911,N_18571,N_18026);
nor U18912 (N_18912,N_17839,N_18591);
nor U18913 (N_18913,N_18032,N_18536);
or U18914 (N_18914,N_18044,N_18574);
nand U18915 (N_18915,N_18310,N_18089);
nand U18916 (N_18916,N_18130,N_18535);
and U18917 (N_18917,N_18436,N_17816);
and U18918 (N_18918,N_17501,N_18668);
nor U18919 (N_18919,N_18421,N_17602);
nor U18920 (N_18920,N_18500,N_17617);
nor U18921 (N_18921,N_18641,N_18202);
nor U18922 (N_18922,N_18099,N_18009);
xor U18923 (N_18923,N_17692,N_18365);
and U18924 (N_18924,N_18159,N_17836);
xnor U18925 (N_18925,N_18656,N_18484);
and U18926 (N_18926,N_18610,N_18602);
nor U18927 (N_18927,N_18033,N_18372);
or U18928 (N_18928,N_18588,N_17827);
xnor U18929 (N_18929,N_18023,N_17941);
nand U18930 (N_18930,N_18073,N_17649);
and U18931 (N_18931,N_17807,N_18546);
xor U18932 (N_18932,N_18269,N_17843);
xor U18933 (N_18933,N_18749,N_18397);
or U18934 (N_18934,N_17509,N_17700);
nand U18935 (N_18935,N_17732,N_18399);
and U18936 (N_18936,N_18011,N_18715);
and U18937 (N_18937,N_17852,N_18452);
xnor U18938 (N_18938,N_18512,N_18056);
and U18939 (N_18939,N_18012,N_18550);
or U18940 (N_18940,N_17668,N_18605);
and U18941 (N_18941,N_17908,N_18606);
or U18942 (N_18942,N_18223,N_18449);
and U18943 (N_18943,N_18597,N_18585);
and U18944 (N_18944,N_18666,N_18724);
xor U18945 (N_18945,N_18673,N_17669);
or U18946 (N_18946,N_17999,N_18489);
nand U18947 (N_18947,N_17858,N_18380);
nand U18948 (N_18948,N_18733,N_17582);
or U18949 (N_18949,N_17970,N_18052);
nor U18950 (N_18950,N_18448,N_18675);
and U18951 (N_18951,N_18630,N_17966);
and U18952 (N_18952,N_17787,N_18686);
or U18953 (N_18953,N_17537,N_18261);
xor U18954 (N_18954,N_17718,N_18303);
xnor U18955 (N_18955,N_17867,N_18293);
nand U18956 (N_18956,N_18700,N_18361);
nor U18957 (N_18957,N_17503,N_18527);
and U18958 (N_18958,N_18201,N_18037);
nor U18959 (N_18959,N_17686,N_17542);
nand U18960 (N_18960,N_18426,N_18047);
nand U18961 (N_18961,N_17674,N_17672);
xor U18962 (N_18962,N_17654,N_17715);
nand U18963 (N_18963,N_18087,N_18486);
nor U18964 (N_18964,N_17841,N_17737);
and U18965 (N_18965,N_18329,N_17741);
and U18966 (N_18966,N_18548,N_17911);
or U18967 (N_18967,N_17544,N_18608);
and U18968 (N_18968,N_18693,N_17747);
xor U18969 (N_18969,N_18575,N_17864);
and U18970 (N_18970,N_18458,N_17713);
nand U18971 (N_18971,N_18390,N_18339);
or U18972 (N_18972,N_18064,N_17800);
nor U18973 (N_18973,N_18296,N_18212);
nor U18974 (N_18974,N_18181,N_18701);
nand U18975 (N_18975,N_18036,N_18141);
nand U18976 (N_18976,N_18031,N_18093);
nor U18977 (N_18977,N_17982,N_18568);
or U18978 (N_18978,N_17569,N_17920);
nor U18979 (N_18979,N_18149,N_17673);
nand U18980 (N_18980,N_18534,N_18294);
nor U18981 (N_18981,N_18412,N_18097);
or U18982 (N_18982,N_18603,N_17840);
nand U18983 (N_18983,N_17962,N_17541);
and U18984 (N_18984,N_17678,N_17774);
xor U18985 (N_18985,N_17709,N_18213);
and U18986 (N_18986,N_18680,N_18220);
nand U18987 (N_18987,N_17746,N_18300);
or U18988 (N_18988,N_18071,N_17593);
xor U18989 (N_18989,N_18110,N_17567);
and U18990 (N_18990,N_18180,N_18207);
nor U18991 (N_18991,N_18003,N_18528);
nor U18992 (N_18992,N_18572,N_18472);
nand U18993 (N_18993,N_18253,N_18173);
nand U18994 (N_18994,N_18204,N_18080);
nor U18995 (N_18995,N_18353,N_18503);
or U18996 (N_18996,N_18351,N_17502);
and U18997 (N_18997,N_17828,N_18583);
or U18998 (N_18998,N_17870,N_17684);
nand U18999 (N_18999,N_17586,N_17863);
xnor U19000 (N_19000,N_17610,N_18494);
xnor U19001 (N_19001,N_17685,N_17550);
nor U19002 (N_19002,N_18153,N_17664);
nand U19003 (N_19003,N_18103,N_18587);
and U19004 (N_19004,N_17533,N_17619);
xor U19005 (N_19005,N_18595,N_17735);
or U19006 (N_19006,N_18352,N_18748);
xnor U19007 (N_19007,N_18663,N_18393);
or U19008 (N_19008,N_18647,N_18501);
nor U19009 (N_19009,N_18725,N_17762);
xor U19010 (N_19010,N_17902,N_18368);
nand U19011 (N_19011,N_18406,N_17777);
xnor U19012 (N_19012,N_17757,N_17690);
and U19013 (N_19013,N_17968,N_18322);
nand U19014 (N_19014,N_17566,N_18601);
and U19015 (N_19015,N_18267,N_17589);
nand U19016 (N_19016,N_18369,N_18382);
xor U19017 (N_19017,N_18410,N_17979);
or U19018 (N_19018,N_18286,N_17707);
and U19019 (N_19019,N_17596,N_18604);
or U19020 (N_19020,N_18161,N_18133);
and U19021 (N_19021,N_17764,N_18332);
or U19022 (N_19022,N_18030,N_18374);
nor U19023 (N_19023,N_18341,N_18091);
and U19024 (N_19024,N_17793,N_18578);
and U19025 (N_19025,N_18008,N_18205);
xor U19026 (N_19026,N_18119,N_17922);
or U19027 (N_19027,N_18623,N_17598);
nor U19028 (N_19028,N_18198,N_18665);
or U19029 (N_19029,N_17776,N_18567);
nor U19030 (N_19030,N_18191,N_18155);
nand U19031 (N_19031,N_18590,N_18433);
and U19032 (N_19032,N_18288,N_17708);
or U19033 (N_19033,N_17752,N_18556);
xnor U19034 (N_19034,N_17659,N_18726);
nand U19035 (N_19035,N_17733,N_18058);
nor U19036 (N_19036,N_17529,N_18034);
and U19037 (N_19037,N_17899,N_18682);
nand U19038 (N_19038,N_18274,N_18523);
nand U19039 (N_19039,N_18439,N_18408);
or U19040 (N_19040,N_17731,N_18704);
nand U19041 (N_19041,N_17880,N_18240);
nor U19042 (N_19042,N_18069,N_17772);
xnor U19043 (N_19043,N_17898,N_18389);
nor U19044 (N_19044,N_17641,N_18739);
xnor U19045 (N_19045,N_17795,N_17869);
and U19046 (N_19046,N_17967,N_17644);
or U19047 (N_19047,N_17702,N_18206);
or U19048 (N_19048,N_18327,N_17750);
nand U19049 (N_19049,N_18506,N_17536);
and U19050 (N_19050,N_17866,N_17719);
xnor U19051 (N_19051,N_18637,N_18626);
xor U19052 (N_19052,N_18537,N_18598);
or U19053 (N_19053,N_17960,N_18232);
nand U19054 (N_19054,N_17725,N_18717);
or U19055 (N_19055,N_18692,N_18622);
nor U19056 (N_19056,N_18435,N_17761);
and U19057 (N_19057,N_17627,N_17561);
or U19058 (N_19058,N_18264,N_18025);
or U19059 (N_19059,N_18194,N_17576);
nand U19060 (N_19060,N_18027,N_18718);
nor U19061 (N_19061,N_17721,N_18381);
xnor U19062 (N_19062,N_17753,N_17919);
xnor U19063 (N_19063,N_18525,N_17859);
xor U19064 (N_19064,N_18531,N_18345);
and U19065 (N_19065,N_17527,N_18016);
xnor U19066 (N_19066,N_17538,N_17653);
nor U19067 (N_19067,N_17618,N_17531);
nor U19068 (N_19068,N_17722,N_18115);
nand U19069 (N_19069,N_18396,N_17942);
nor U19070 (N_19070,N_17565,N_18388);
and U19071 (N_19071,N_18136,N_18278);
or U19072 (N_19072,N_17952,N_18335);
nand U19073 (N_19073,N_17796,N_17638);
nor U19074 (N_19074,N_18273,N_17743);
xor U19075 (N_19075,N_17543,N_18404);
and U19076 (N_19076,N_18135,N_17712);
nor U19077 (N_19077,N_18456,N_17564);
xnor U19078 (N_19078,N_18129,N_17993);
nand U19079 (N_19079,N_18346,N_17604);
nor U19080 (N_19080,N_18019,N_18331);
and U19081 (N_19081,N_18362,N_18391);
nand U19082 (N_19082,N_18650,N_17829);
or U19083 (N_19083,N_18246,N_17648);
or U19084 (N_19084,N_17711,N_17551);
and U19085 (N_19085,N_18225,N_18616);
or U19086 (N_19086,N_17514,N_17892);
or U19087 (N_19087,N_18539,N_18075);
and U19088 (N_19088,N_18416,N_18499);
and U19089 (N_19089,N_17730,N_17976);
xnor U19090 (N_19090,N_18411,N_17784);
nor U19091 (N_19091,N_17590,N_17972);
xnor U19092 (N_19092,N_17925,N_18295);
and U19093 (N_19093,N_18157,N_17913);
nor U19094 (N_19094,N_18242,N_17599);
and U19095 (N_19095,N_17535,N_18466);
nand U19096 (N_19096,N_18655,N_18620);
or U19097 (N_19097,N_18152,N_18330);
nor U19098 (N_19098,N_18740,N_17637);
nand U19099 (N_19099,N_17837,N_18526);
or U19100 (N_19100,N_18440,N_17824);
and U19101 (N_19101,N_17917,N_17739);
or U19102 (N_19102,N_18651,N_18265);
and U19103 (N_19103,N_18681,N_18459);
xor U19104 (N_19104,N_18617,N_18737);
xnor U19105 (N_19105,N_17568,N_17825);
or U19106 (N_19106,N_18515,N_18356);
nor U19107 (N_19107,N_18559,N_18579);
or U19108 (N_19108,N_18271,N_18200);
xnor U19109 (N_19109,N_17971,N_18101);
xor U19110 (N_19110,N_17927,N_17640);
xor U19111 (N_19111,N_17571,N_17887);
nor U19112 (N_19112,N_17519,N_18138);
and U19113 (N_19113,N_17516,N_18022);
nand U19114 (N_19114,N_17935,N_18395);
and U19115 (N_19115,N_18299,N_18083);
nand U19116 (N_19116,N_18187,N_18582);
and U19117 (N_19117,N_17939,N_17591);
nand U19118 (N_19118,N_17676,N_18678);
xor U19119 (N_19119,N_18095,N_18446);
xor U19120 (N_19120,N_17802,N_18017);
or U19121 (N_19121,N_18005,N_18285);
nor U19122 (N_19122,N_18371,N_18066);
nand U19123 (N_19123,N_18581,N_17767);
xor U19124 (N_19124,N_18713,N_17742);
nand U19125 (N_19125,N_18485,N_18518);
and U19126 (N_19126,N_18465,N_17539);
and U19127 (N_19127,N_17675,N_18479);
or U19128 (N_19128,N_18355,N_17884);
nor U19129 (N_19129,N_18703,N_18660);
nor U19130 (N_19130,N_18552,N_18541);
xnor U19131 (N_19131,N_17635,N_18478);
nor U19132 (N_19132,N_18427,N_18521);
and U19133 (N_19133,N_17650,N_18551);
nand U19134 (N_19134,N_18473,N_18308);
xor U19135 (N_19135,N_18054,N_18511);
nand U19136 (N_19136,N_17532,N_18600);
and U19137 (N_19137,N_18291,N_17835);
and U19138 (N_19138,N_17933,N_17623);
nand U19139 (N_19139,N_18540,N_17811);
nand U19140 (N_19140,N_17728,N_17534);
nand U19141 (N_19141,N_18607,N_18082);
or U19142 (N_19142,N_17988,N_18558);
and U19143 (N_19143,N_18744,N_18314);
or U19144 (N_19144,N_18621,N_18469);
nor U19145 (N_19145,N_17775,N_17907);
nand U19146 (N_19146,N_17965,N_17738);
nor U19147 (N_19147,N_17855,N_18145);
and U19148 (N_19148,N_18423,N_17846);
xor U19149 (N_19149,N_18055,N_18648);
xnor U19150 (N_19150,N_18096,N_18143);
or U19151 (N_19151,N_18196,N_18514);
nor U19152 (N_19152,N_18316,N_18488);
or U19153 (N_19153,N_17661,N_18658);
and U19154 (N_19154,N_18116,N_18653);
xor U19155 (N_19155,N_18021,N_17847);
or U19156 (N_19156,N_18674,N_17716);
nor U19157 (N_19157,N_18313,N_17928);
nand U19158 (N_19158,N_18599,N_18248);
xnor U19159 (N_19159,N_18533,N_17647);
or U19160 (N_19160,N_18731,N_18613);
nand U19161 (N_19161,N_17818,N_18460);
nor U19162 (N_19162,N_17779,N_18419);
xnor U19163 (N_19163,N_17682,N_18688);
nor U19164 (N_19164,N_18728,N_18306);
nand U19165 (N_19165,N_18576,N_18520);
xor U19166 (N_19166,N_18363,N_18502);
xor U19167 (N_19167,N_18350,N_17726);
or U19168 (N_19168,N_17985,N_18228);
nand U19169 (N_19169,N_18199,N_18280);
and U19170 (N_19170,N_18182,N_17934);
and U19171 (N_19171,N_18475,N_17996);
nor U19172 (N_19172,N_18505,N_18120);
or U19173 (N_19173,N_18188,N_17786);
nor U19174 (N_19174,N_17691,N_17891);
xor U19175 (N_19175,N_18722,N_18326);
nand U19176 (N_19176,N_17886,N_17983);
xnor U19177 (N_19177,N_17936,N_17687);
nor U19178 (N_19178,N_18732,N_18179);
or U19179 (N_19179,N_17724,N_17937);
nor U19180 (N_19180,N_18287,N_17973);
xnor U19181 (N_19181,N_18609,N_18134);
nor U19182 (N_19182,N_18487,N_18266);
or U19183 (N_19183,N_18172,N_18696);
and U19184 (N_19184,N_18625,N_18347);
or U19185 (N_19185,N_18298,N_18615);
nand U19186 (N_19186,N_18118,N_18243);
nor U19187 (N_19187,N_18276,N_18417);
nand U19188 (N_19188,N_18079,N_18124);
xnor U19189 (N_19189,N_17525,N_17694);
or U19190 (N_19190,N_18394,N_18122);
xor U19191 (N_19191,N_17990,N_18689);
xnor U19192 (N_19192,N_17717,N_17624);
xor U19193 (N_19193,N_17799,N_18186);
and U19194 (N_19194,N_18190,N_18318);
or U19195 (N_19195,N_17823,N_17878);
and U19196 (N_19196,N_17945,N_18413);
and U19197 (N_19197,N_18364,N_17923);
xnor U19198 (N_19198,N_18349,N_17833);
and U19199 (N_19199,N_18476,N_18209);
nor U19200 (N_19200,N_18259,N_18260);
nor U19201 (N_19201,N_18210,N_17758);
and U19202 (N_19202,N_18262,N_18062);
nand U19203 (N_19203,N_18222,N_18497);
nor U19204 (N_19204,N_18000,N_18721);
nand U19205 (N_19205,N_18268,N_17563);
xnor U19206 (N_19206,N_18176,N_17513);
xor U19207 (N_19207,N_18348,N_18102);
nand U19208 (N_19208,N_18694,N_18059);
and U19209 (N_19209,N_18628,N_18002);
nand U19210 (N_19210,N_18375,N_17946);
xnor U19211 (N_19211,N_17954,N_18156);
or U19212 (N_19212,N_18592,N_17792);
nand U19213 (N_19213,N_17992,N_17819);
nand U19214 (N_19214,N_17573,N_17932);
or U19215 (N_19215,N_18166,N_18414);
and U19216 (N_19216,N_17643,N_17904);
or U19217 (N_19217,N_17559,N_17831);
nand U19218 (N_19218,N_18177,N_18251);
xor U19219 (N_19219,N_18451,N_18117);
nand U19220 (N_19220,N_18509,N_17696);
or U19221 (N_19221,N_18569,N_17820);
xor U19222 (N_19222,N_18624,N_18508);
xnor U19223 (N_19223,N_18516,N_18457);
or U19224 (N_19224,N_18640,N_18560);
nor U19225 (N_19225,N_17879,N_18001);
nor U19226 (N_19226,N_17783,N_17771);
or U19227 (N_19227,N_18387,N_18252);
and U19228 (N_19228,N_17805,N_17515);
and U19229 (N_19229,N_17929,N_18664);
and U19230 (N_19230,N_18443,N_18144);
xnor U19231 (N_19231,N_17974,N_17710);
xor U19232 (N_19232,N_18679,N_18140);
xnor U19233 (N_19233,N_17621,N_18168);
or U19234 (N_19234,N_17740,N_18400);
and U19235 (N_19235,N_18418,N_17881);
nor U19236 (N_19236,N_17850,N_18441);
xor U19237 (N_19237,N_17572,N_17714);
and U19238 (N_19238,N_18554,N_18690);
xnor U19239 (N_19239,N_18305,N_18237);
and U19240 (N_19240,N_17612,N_17504);
nor U19241 (N_19241,N_17755,N_18378);
or U19242 (N_19242,N_17821,N_17801);
xor U19243 (N_19243,N_18284,N_17557);
nor U19244 (N_19244,N_18661,N_17583);
nor U19245 (N_19245,N_18065,N_17773);
xnor U19246 (N_19246,N_18215,N_17594);
xnor U19247 (N_19247,N_18430,N_18636);
nand U19248 (N_19248,N_18734,N_17699);
nor U19249 (N_19249,N_17748,N_18730);
and U19250 (N_19250,N_18463,N_17900);
and U19251 (N_19251,N_18004,N_18645);
xnor U19252 (N_19252,N_18105,N_18123);
and U19253 (N_19253,N_17797,N_18216);
nor U19254 (N_19254,N_17998,N_18727);
xor U19255 (N_19255,N_18167,N_18109);
xor U19256 (N_19256,N_17698,N_17903);
or U19257 (N_19257,N_18557,N_18614);
and U19258 (N_19258,N_18708,N_17788);
and U19259 (N_19259,N_18745,N_18434);
and U19260 (N_19260,N_18562,N_17553);
or U19261 (N_19261,N_17671,N_18226);
nand U19262 (N_19262,N_18270,N_17930);
nor U19263 (N_19263,N_17549,N_18627);
and U19264 (N_19264,N_17975,N_18113);
and U19265 (N_19265,N_18670,N_18524);
and U19266 (N_19266,N_18272,N_18074);
nand U19267 (N_19267,N_17636,N_18085);
nand U19268 (N_19268,N_17794,N_18593);
nor U19269 (N_19269,N_18057,N_18247);
and U19270 (N_19270,N_18342,N_18307);
xnor U19271 (N_19271,N_17622,N_17782);
nor U19272 (N_19272,N_17980,N_17812);
xnor U19273 (N_19273,N_17688,N_18425);
nand U19274 (N_19274,N_18379,N_18060);
nor U19275 (N_19275,N_17778,N_17615);
and U19276 (N_19276,N_18325,N_17842);
nand U19277 (N_19277,N_18401,N_18723);
nand U19278 (N_19278,N_17948,N_18040);
nand U19279 (N_19279,N_17592,N_17765);
xor U19280 (N_19280,N_17667,N_18657);
or U19281 (N_19281,N_17581,N_18111);
nand U19282 (N_19282,N_18432,N_18244);
nand U19283 (N_19283,N_18483,N_18015);
nand U19284 (N_19284,N_18480,N_18741);
and U19285 (N_19285,N_17660,N_18289);
nand U19286 (N_19286,N_18048,N_17789);
xor U19287 (N_19287,N_17940,N_18462);
nor U19288 (N_19288,N_18343,N_17545);
nand U19289 (N_19289,N_17914,N_18357);
or U19290 (N_19290,N_17991,N_18132);
xor U19291 (N_19291,N_18577,N_17871);
xor U19292 (N_19292,N_18014,N_17834);
nor U19293 (N_19293,N_17977,N_18422);
nand U19294 (N_19294,N_17838,N_18611);
and U19295 (N_19295,N_18510,N_17658);
or U19296 (N_19296,N_17814,N_17857);
nand U19297 (N_19297,N_18743,N_18445);
xnor U19298 (N_19298,N_17633,N_18231);
nor U19299 (N_19299,N_18471,N_18612);
xnor U19300 (N_19300,N_18208,N_18233);
nand U19301 (N_19301,N_17703,N_17888);
nand U19302 (N_19302,N_17893,N_18453);
nand U19303 (N_19303,N_17547,N_18649);
nor U19304 (N_19304,N_18684,N_18492);
nand U19305 (N_19305,N_18084,N_17605);
xor U19306 (N_19306,N_17720,N_17832);
nand U19307 (N_19307,N_18236,N_18706);
or U19308 (N_19308,N_17530,N_18710);
or U19309 (N_19309,N_17642,N_17931);
nand U19310 (N_19310,N_18189,N_17895);
or U19311 (N_19311,N_17809,N_17704);
or U19312 (N_19312,N_17597,N_18051);
nand U19313 (N_19313,N_17657,N_18634);
nor U19314 (N_19314,N_18010,N_18474);
nand U19315 (N_19315,N_18677,N_18596);
nand U19316 (N_19316,N_17803,N_18104);
and U19317 (N_19317,N_18642,N_17849);
or U19318 (N_19318,N_18392,N_17645);
and U19319 (N_19319,N_17845,N_18094);
xnor U19320 (N_19320,N_18635,N_18570);
xor U19321 (N_19321,N_18738,N_18013);
and U19322 (N_19322,N_17607,N_18709);
xor U19323 (N_19323,N_18683,N_18151);
xor U19324 (N_19324,N_18490,N_17520);
nand U19325 (N_19325,N_18386,N_17628);
or U19326 (N_19326,N_17570,N_17555);
nor U19327 (N_19327,N_17848,N_18290);
nor U19328 (N_19328,N_17608,N_18321);
and U19329 (N_19329,N_17984,N_18405);
xnor U19330 (N_19330,N_17905,N_18667);
and U19331 (N_19331,N_18241,N_18092);
xor U19332 (N_19332,N_18563,N_18041);
and U19333 (N_19333,N_17556,N_18633);
nand U19334 (N_19334,N_18067,N_18107);
and U19335 (N_19335,N_17680,N_18076);
nand U19336 (N_19336,N_18081,N_17854);
nand U19337 (N_19337,N_18028,N_17554);
nor U19338 (N_19338,N_18072,N_18619);
and U19339 (N_19339,N_17508,N_18234);
and U19340 (N_19340,N_17723,N_18720);
or U19341 (N_19341,N_17512,N_17548);
xor U19342 (N_19342,N_17585,N_17978);
xor U19343 (N_19343,N_18424,N_18742);
or U19344 (N_19344,N_17744,N_17522);
nand U19345 (N_19345,N_18519,N_18214);
xor U19346 (N_19346,N_18698,N_18127);
xor U19347 (N_19347,N_18747,N_18707);
and U19348 (N_19348,N_18461,N_17706);
nor U19349 (N_19349,N_18545,N_18384);
or U19350 (N_19350,N_17804,N_17872);
and U19351 (N_19351,N_17995,N_18211);
or U19352 (N_19352,N_18218,N_18652);
nor U19353 (N_19353,N_17943,N_18530);
xor U19354 (N_19354,N_18139,N_17830);
xnor U19355 (N_19355,N_18495,N_17860);
xor U19356 (N_19356,N_17780,N_18061);
xnor U19357 (N_19357,N_17558,N_17562);
xnor U19358 (N_19358,N_18174,N_18555);
or U19359 (N_19359,N_18100,N_17600);
nor U19360 (N_19360,N_18477,N_18496);
or U19361 (N_19361,N_18444,N_17579);
or U19362 (N_19362,N_18221,N_17997);
xor U19363 (N_19363,N_17808,N_17938);
nor U19364 (N_19364,N_17524,N_17883);
or U19365 (N_19365,N_18171,N_17909);
or U19366 (N_19366,N_17552,N_17785);
xor U19367 (N_19367,N_18150,N_18376);
nand U19368 (N_19368,N_18407,N_17630);
nor U19369 (N_19369,N_18669,N_18045);
nand U19370 (N_19370,N_18699,N_18320);
or U19371 (N_19371,N_18279,N_18283);
nor U19372 (N_19372,N_18164,N_17601);
nand U19373 (N_19373,N_18662,N_17697);
and U19374 (N_19374,N_17826,N_18029);
or U19375 (N_19375,N_17722,N_18310);
nand U19376 (N_19376,N_18263,N_17801);
nor U19377 (N_19377,N_18025,N_17957);
and U19378 (N_19378,N_17575,N_17986);
or U19379 (N_19379,N_17706,N_18682);
and U19380 (N_19380,N_17919,N_18235);
nand U19381 (N_19381,N_18718,N_18365);
xnor U19382 (N_19382,N_18355,N_17615);
nand U19383 (N_19383,N_17977,N_17936);
nand U19384 (N_19384,N_18295,N_17781);
xor U19385 (N_19385,N_17820,N_18668);
nor U19386 (N_19386,N_18574,N_18409);
xor U19387 (N_19387,N_18172,N_18267);
and U19388 (N_19388,N_18440,N_17675);
xor U19389 (N_19389,N_17804,N_17513);
xor U19390 (N_19390,N_17805,N_18053);
nand U19391 (N_19391,N_17941,N_17718);
nand U19392 (N_19392,N_17736,N_18505);
nand U19393 (N_19393,N_17954,N_18260);
and U19394 (N_19394,N_17936,N_17718);
nor U19395 (N_19395,N_18224,N_18609);
or U19396 (N_19396,N_18703,N_18237);
or U19397 (N_19397,N_18249,N_17955);
xnor U19398 (N_19398,N_17926,N_17794);
xor U19399 (N_19399,N_17838,N_18572);
nor U19400 (N_19400,N_17772,N_17635);
nand U19401 (N_19401,N_18087,N_18263);
or U19402 (N_19402,N_18159,N_18070);
or U19403 (N_19403,N_18566,N_18137);
and U19404 (N_19404,N_18188,N_18082);
nor U19405 (N_19405,N_17716,N_18159);
xor U19406 (N_19406,N_18698,N_17728);
nand U19407 (N_19407,N_18593,N_18449);
nor U19408 (N_19408,N_18144,N_17799);
nand U19409 (N_19409,N_17506,N_18235);
or U19410 (N_19410,N_17870,N_17827);
nor U19411 (N_19411,N_17771,N_18181);
or U19412 (N_19412,N_18033,N_18182);
and U19413 (N_19413,N_17931,N_17852);
nor U19414 (N_19414,N_17827,N_17508);
nand U19415 (N_19415,N_17560,N_18349);
or U19416 (N_19416,N_17917,N_18492);
nor U19417 (N_19417,N_18398,N_18162);
and U19418 (N_19418,N_17913,N_18144);
and U19419 (N_19419,N_17908,N_18721);
xor U19420 (N_19420,N_17646,N_17963);
or U19421 (N_19421,N_18746,N_17920);
and U19422 (N_19422,N_17933,N_18338);
nand U19423 (N_19423,N_18119,N_17563);
and U19424 (N_19424,N_18624,N_17897);
nor U19425 (N_19425,N_17530,N_17639);
nand U19426 (N_19426,N_17554,N_18126);
nor U19427 (N_19427,N_17741,N_18327);
nor U19428 (N_19428,N_17730,N_18499);
or U19429 (N_19429,N_17512,N_18627);
xnor U19430 (N_19430,N_18443,N_18598);
xnor U19431 (N_19431,N_17723,N_17735);
nand U19432 (N_19432,N_18219,N_18134);
and U19433 (N_19433,N_18001,N_18215);
or U19434 (N_19434,N_17694,N_18650);
nand U19435 (N_19435,N_18001,N_18604);
xor U19436 (N_19436,N_18321,N_17597);
xor U19437 (N_19437,N_18108,N_18599);
nand U19438 (N_19438,N_18001,N_17943);
nor U19439 (N_19439,N_18177,N_18174);
nor U19440 (N_19440,N_17997,N_18114);
and U19441 (N_19441,N_18001,N_18075);
and U19442 (N_19442,N_17655,N_18563);
nor U19443 (N_19443,N_18742,N_18049);
nand U19444 (N_19444,N_17704,N_17524);
nand U19445 (N_19445,N_18444,N_18315);
nand U19446 (N_19446,N_17837,N_18583);
xnor U19447 (N_19447,N_17799,N_18545);
and U19448 (N_19448,N_17952,N_18729);
or U19449 (N_19449,N_17508,N_17523);
xor U19450 (N_19450,N_17535,N_18703);
and U19451 (N_19451,N_18149,N_17629);
or U19452 (N_19452,N_17646,N_18414);
or U19453 (N_19453,N_18746,N_18706);
nand U19454 (N_19454,N_18470,N_18446);
xor U19455 (N_19455,N_17897,N_18555);
or U19456 (N_19456,N_17970,N_18047);
nor U19457 (N_19457,N_17602,N_17904);
and U19458 (N_19458,N_18087,N_18148);
xor U19459 (N_19459,N_18439,N_18183);
nand U19460 (N_19460,N_18122,N_17965);
nor U19461 (N_19461,N_18715,N_18691);
nor U19462 (N_19462,N_17953,N_17757);
nor U19463 (N_19463,N_18327,N_18347);
xnor U19464 (N_19464,N_18130,N_18035);
xor U19465 (N_19465,N_18309,N_18412);
nand U19466 (N_19466,N_17762,N_18458);
xor U19467 (N_19467,N_17853,N_18670);
nor U19468 (N_19468,N_18290,N_18627);
nor U19469 (N_19469,N_18126,N_17602);
nor U19470 (N_19470,N_18202,N_18203);
nand U19471 (N_19471,N_18493,N_17986);
xnor U19472 (N_19472,N_18528,N_18177);
or U19473 (N_19473,N_18183,N_18547);
nor U19474 (N_19474,N_17909,N_17787);
xnor U19475 (N_19475,N_18375,N_17530);
nand U19476 (N_19476,N_18302,N_17988);
nand U19477 (N_19477,N_17791,N_18160);
nor U19478 (N_19478,N_18309,N_18157);
nor U19479 (N_19479,N_18109,N_18625);
or U19480 (N_19480,N_17684,N_18022);
xnor U19481 (N_19481,N_18609,N_17952);
nand U19482 (N_19482,N_18273,N_18227);
or U19483 (N_19483,N_17651,N_18109);
and U19484 (N_19484,N_18658,N_17758);
nor U19485 (N_19485,N_17698,N_18470);
nand U19486 (N_19486,N_18054,N_18032);
nand U19487 (N_19487,N_18702,N_18149);
or U19488 (N_19488,N_17619,N_17674);
nor U19489 (N_19489,N_18092,N_17809);
or U19490 (N_19490,N_17945,N_17601);
or U19491 (N_19491,N_18636,N_18501);
nand U19492 (N_19492,N_18002,N_18036);
xnor U19493 (N_19493,N_17617,N_18676);
nand U19494 (N_19494,N_18548,N_17997);
nor U19495 (N_19495,N_18037,N_17880);
nor U19496 (N_19496,N_18463,N_18096);
nand U19497 (N_19497,N_17562,N_18303);
nand U19498 (N_19498,N_18252,N_17761);
xnor U19499 (N_19499,N_18497,N_17926);
and U19500 (N_19500,N_18470,N_18163);
nor U19501 (N_19501,N_17768,N_18423);
or U19502 (N_19502,N_18668,N_17809);
or U19503 (N_19503,N_17972,N_18034);
and U19504 (N_19504,N_18629,N_18247);
and U19505 (N_19505,N_18208,N_18422);
nand U19506 (N_19506,N_17593,N_18318);
xnor U19507 (N_19507,N_17911,N_18596);
nand U19508 (N_19508,N_18703,N_17554);
xor U19509 (N_19509,N_18120,N_17640);
nor U19510 (N_19510,N_17555,N_17594);
nor U19511 (N_19511,N_17819,N_18203);
nor U19512 (N_19512,N_18433,N_17944);
nor U19513 (N_19513,N_17816,N_18314);
or U19514 (N_19514,N_17938,N_18582);
and U19515 (N_19515,N_18156,N_18173);
xor U19516 (N_19516,N_17625,N_18186);
nor U19517 (N_19517,N_17917,N_17723);
xnor U19518 (N_19518,N_18348,N_18246);
nand U19519 (N_19519,N_18094,N_18220);
nand U19520 (N_19520,N_17506,N_18431);
and U19521 (N_19521,N_18269,N_18411);
xnor U19522 (N_19522,N_17766,N_18299);
xor U19523 (N_19523,N_18185,N_18364);
nor U19524 (N_19524,N_18153,N_17990);
and U19525 (N_19525,N_18326,N_18360);
or U19526 (N_19526,N_17949,N_18182);
nor U19527 (N_19527,N_18110,N_17551);
and U19528 (N_19528,N_18277,N_17524);
or U19529 (N_19529,N_17902,N_18185);
xor U19530 (N_19530,N_17901,N_17635);
nor U19531 (N_19531,N_18411,N_17752);
nor U19532 (N_19532,N_17883,N_17889);
and U19533 (N_19533,N_17625,N_17706);
nor U19534 (N_19534,N_18428,N_17979);
xor U19535 (N_19535,N_18160,N_18571);
nor U19536 (N_19536,N_18419,N_18146);
and U19537 (N_19537,N_17836,N_17581);
xor U19538 (N_19538,N_18128,N_17716);
or U19539 (N_19539,N_17851,N_18225);
xnor U19540 (N_19540,N_18702,N_18609);
nor U19541 (N_19541,N_18357,N_17969);
nor U19542 (N_19542,N_17659,N_18595);
and U19543 (N_19543,N_18212,N_17612);
and U19544 (N_19544,N_18514,N_17608);
and U19545 (N_19545,N_18232,N_17576);
or U19546 (N_19546,N_18324,N_18692);
xnor U19547 (N_19547,N_18261,N_17586);
or U19548 (N_19548,N_17707,N_18352);
and U19549 (N_19549,N_18180,N_17517);
nand U19550 (N_19550,N_18505,N_17700);
xnor U19551 (N_19551,N_18481,N_18629);
nand U19552 (N_19552,N_18464,N_17625);
xnor U19553 (N_19553,N_17992,N_18282);
and U19554 (N_19554,N_18194,N_17980);
or U19555 (N_19555,N_18703,N_18046);
xor U19556 (N_19556,N_18607,N_18439);
nand U19557 (N_19557,N_18743,N_17774);
nand U19558 (N_19558,N_18274,N_18449);
and U19559 (N_19559,N_18716,N_18258);
nand U19560 (N_19560,N_17651,N_18440);
or U19561 (N_19561,N_18681,N_18606);
xor U19562 (N_19562,N_17861,N_18624);
or U19563 (N_19563,N_17937,N_18240);
nand U19564 (N_19564,N_17654,N_18033);
and U19565 (N_19565,N_18659,N_18522);
nand U19566 (N_19566,N_18219,N_17693);
xor U19567 (N_19567,N_18326,N_17821);
and U19568 (N_19568,N_18246,N_18028);
nand U19569 (N_19569,N_17720,N_18632);
xor U19570 (N_19570,N_18259,N_18393);
xor U19571 (N_19571,N_18503,N_18104);
xor U19572 (N_19572,N_18518,N_18055);
and U19573 (N_19573,N_17909,N_18014);
nor U19574 (N_19574,N_18116,N_17829);
or U19575 (N_19575,N_17982,N_17997);
nor U19576 (N_19576,N_17977,N_17536);
nor U19577 (N_19577,N_18182,N_18447);
and U19578 (N_19578,N_17790,N_18508);
xor U19579 (N_19579,N_17539,N_18010);
or U19580 (N_19580,N_18065,N_18028);
xnor U19581 (N_19581,N_18024,N_18365);
and U19582 (N_19582,N_18560,N_18686);
nand U19583 (N_19583,N_18656,N_17770);
xnor U19584 (N_19584,N_18643,N_17757);
nand U19585 (N_19585,N_18530,N_18653);
xor U19586 (N_19586,N_17763,N_18057);
and U19587 (N_19587,N_17909,N_18442);
nor U19588 (N_19588,N_17686,N_18732);
nor U19589 (N_19589,N_18714,N_18491);
nor U19590 (N_19590,N_18162,N_17531);
nand U19591 (N_19591,N_18146,N_18262);
nand U19592 (N_19592,N_17686,N_18053);
xnor U19593 (N_19593,N_17943,N_18185);
xnor U19594 (N_19594,N_18657,N_17700);
nand U19595 (N_19595,N_17781,N_18058);
and U19596 (N_19596,N_18418,N_18229);
xnor U19597 (N_19597,N_18260,N_18436);
xnor U19598 (N_19598,N_17534,N_18065);
nand U19599 (N_19599,N_17864,N_17808);
or U19600 (N_19600,N_18608,N_17558);
xnor U19601 (N_19601,N_18585,N_18708);
nor U19602 (N_19602,N_18006,N_17641);
or U19603 (N_19603,N_17947,N_17832);
and U19604 (N_19604,N_18172,N_18447);
nor U19605 (N_19605,N_18441,N_18241);
nor U19606 (N_19606,N_17733,N_17892);
and U19607 (N_19607,N_18095,N_18484);
nand U19608 (N_19608,N_18298,N_18337);
xnor U19609 (N_19609,N_18487,N_17826);
nand U19610 (N_19610,N_17927,N_17816);
nand U19611 (N_19611,N_18439,N_17958);
or U19612 (N_19612,N_18582,N_18682);
nor U19613 (N_19613,N_18684,N_18734);
and U19614 (N_19614,N_18613,N_18733);
nand U19615 (N_19615,N_17901,N_18320);
nand U19616 (N_19616,N_18419,N_18283);
or U19617 (N_19617,N_18398,N_17870);
nor U19618 (N_19618,N_17810,N_17947);
nand U19619 (N_19619,N_17726,N_17846);
nand U19620 (N_19620,N_18709,N_17929);
nand U19621 (N_19621,N_17913,N_17661);
nor U19622 (N_19622,N_18527,N_18260);
nand U19623 (N_19623,N_18066,N_18257);
or U19624 (N_19624,N_18225,N_18345);
nand U19625 (N_19625,N_17880,N_18363);
xor U19626 (N_19626,N_17733,N_18593);
xnor U19627 (N_19627,N_18347,N_17665);
and U19628 (N_19628,N_17687,N_18487);
and U19629 (N_19629,N_18065,N_18049);
nand U19630 (N_19630,N_18486,N_17606);
and U19631 (N_19631,N_18554,N_17809);
xor U19632 (N_19632,N_17676,N_17593);
and U19633 (N_19633,N_18495,N_17888);
nand U19634 (N_19634,N_18165,N_18402);
nor U19635 (N_19635,N_18406,N_18505);
nand U19636 (N_19636,N_18435,N_17998);
xor U19637 (N_19637,N_18726,N_18553);
nor U19638 (N_19638,N_17541,N_18170);
nand U19639 (N_19639,N_17715,N_18726);
nand U19640 (N_19640,N_17708,N_17994);
or U19641 (N_19641,N_17885,N_17612);
nand U19642 (N_19642,N_17525,N_18144);
nand U19643 (N_19643,N_17672,N_18023);
nor U19644 (N_19644,N_18241,N_18192);
or U19645 (N_19645,N_17551,N_17965);
nor U19646 (N_19646,N_17689,N_18201);
or U19647 (N_19647,N_17833,N_17888);
xor U19648 (N_19648,N_18214,N_17511);
or U19649 (N_19649,N_18362,N_18747);
and U19650 (N_19650,N_17839,N_18747);
or U19651 (N_19651,N_18639,N_18613);
nor U19652 (N_19652,N_17577,N_17931);
xor U19653 (N_19653,N_17786,N_18740);
xor U19654 (N_19654,N_17645,N_18251);
nand U19655 (N_19655,N_18346,N_18284);
nor U19656 (N_19656,N_17660,N_18060);
nand U19657 (N_19657,N_18692,N_17678);
nor U19658 (N_19658,N_18028,N_18471);
or U19659 (N_19659,N_17805,N_18716);
xnor U19660 (N_19660,N_17710,N_17610);
or U19661 (N_19661,N_17652,N_18417);
xnor U19662 (N_19662,N_18113,N_18628);
xnor U19663 (N_19663,N_17943,N_18486);
or U19664 (N_19664,N_17771,N_17791);
or U19665 (N_19665,N_18566,N_18110);
and U19666 (N_19666,N_18459,N_17840);
nor U19667 (N_19667,N_17673,N_17631);
or U19668 (N_19668,N_17787,N_18172);
nand U19669 (N_19669,N_17747,N_18623);
nor U19670 (N_19670,N_17807,N_17533);
nor U19671 (N_19671,N_18121,N_17527);
xnor U19672 (N_19672,N_18198,N_17534);
nand U19673 (N_19673,N_18194,N_17749);
nor U19674 (N_19674,N_18606,N_17616);
or U19675 (N_19675,N_17882,N_17504);
or U19676 (N_19676,N_18644,N_18595);
nand U19677 (N_19677,N_18175,N_17899);
nor U19678 (N_19678,N_18429,N_18550);
nand U19679 (N_19679,N_18119,N_17808);
and U19680 (N_19680,N_17694,N_17903);
or U19681 (N_19681,N_18607,N_18130);
nand U19682 (N_19682,N_18681,N_18409);
xor U19683 (N_19683,N_17974,N_18126);
nor U19684 (N_19684,N_17721,N_17540);
and U19685 (N_19685,N_18188,N_18295);
nor U19686 (N_19686,N_18643,N_17706);
nand U19687 (N_19687,N_18185,N_17852);
nand U19688 (N_19688,N_18140,N_17699);
and U19689 (N_19689,N_17818,N_18341);
and U19690 (N_19690,N_18657,N_18551);
and U19691 (N_19691,N_18472,N_17904);
and U19692 (N_19692,N_17853,N_17798);
and U19693 (N_19693,N_17707,N_18655);
nand U19694 (N_19694,N_18692,N_18444);
or U19695 (N_19695,N_17788,N_17830);
xnor U19696 (N_19696,N_18393,N_18616);
and U19697 (N_19697,N_17679,N_18321);
nor U19698 (N_19698,N_17542,N_18110);
nor U19699 (N_19699,N_17753,N_18497);
xor U19700 (N_19700,N_17613,N_18052);
nand U19701 (N_19701,N_17938,N_18101);
and U19702 (N_19702,N_17723,N_17730);
xor U19703 (N_19703,N_17845,N_18103);
xor U19704 (N_19704,N_18051,N_18346);
nand U19705 (N_19705,N_17745,N_18323);
nor U19706 (N_19706,N_17924,N_17504);
nor U19707 (N_19707,N_18375,N_18525);
nor U19708 (N_19708,N_18548,N_17896);
or U19709 (N_19709,N_18720,N_18167);
or U19710 (N_19710,N_18583,N_18335);
nor U19711 (N_19711,N_18050,N_18324);
nand U19712 (N_19712,N_17547,N_17805);
nor U19713 (N_19713,N_18139,N_18205);
nor U19714 (N_19714,N_17759,N_17681);
nor U19715 (N_19715,N_18141,N_17977);
and U19716 (N_19716,N_18077,N_18666);
or U19717 (N_19717,N_17500,N_17534);
nor U19718 (N_19718,N_17753,N_18209);
and U19719 (N_19719,N_17820,N_18163);
or U19720 (N_19720,N_17735,N_17975);
or U19721 (N_19721,N_17931,N_17929);
and U19722 (N_19722,N_17774,N_17903);
nor U19723 (N_19723,N_17807,N_18019);
and U19724 (N_19724,N_17559,N_17799);
xnor U19725 (N_19725,N_18382,N_17739);
and U19726 (N_19726,N_18260,N_18067);
and U19727 (N_19727,N_18467,N_18500);
xor U19728 (N_19728,N_17977,N_17764);
and U19729 (N_19729,N_17704,N_18329);
xor U19730 (N_19730,N_18385,N_17809);
xor U19731 (N_19731,N_18015,N_17743);
nand U19732 (N_19732,N_17726,N_18610);
or U19733 (N_19733,N_18472,N_18703);
and U19734 (N_19734,N_17730,N_17578);
nor U19735 (N_19735,N_18612,N_17872);
and U19736 (N_19736,N_18567,N_18058);
and U19737 (N_19737,N_17596,N_17747);
and U19738 (N_19738,N_18454,N_17568);
nor U19739 (N_19739,N_18166,N_17916);
nor U19740 (N_19740,N_18273,N_18630);
nor U19741 (N_19741,N_17741,N_18305);
xor U19742 (N_19742,N_17549,N_18730);
xnor U19743 (N_19743,N_18015,N_18285);
nand U19744 (N_19744,N_17818,N_18233);
nor U19745 (N_19745,N_18391,N_18685);
and U19746 (N_19746,N_18145,N_17510);
xnor U19747 (N_19747,N_18645,N_18288);
nor U19748 (N_19748,N_18647,N_17937);
nand U19749 (N_19749,N_18492,N_18006);
nand U19750 (N_19750,N_18520,N_17617);
nand U19751 (N_19751,N_18468,N_18397);
nand U19752 (N_19752,N_18262,N_18025);
xnor U19753 (N_19753,N_17551,N_17862);
nand U19754 (N_19754,N_18400,N_18729);
and U19755 (N_19755,N_17885,N_18105);
nor U19756 (N_19756,N_18013,N_18529);
and U19757 (N_19757,N_17763,N_18526);
nand U19758 (N_19758,N_18098,N_17862);
nor U19759 (N_19759,N_18402,N_18046);
nand U19760 (N_19760,N_18661,N_18344);
nand U19761 (N_19761,N_17943,N_17724);
nand U19762 (N_19762,N_17930,N_18661);
xnor U19763 (N_19763,N_18661,N_17643);
nand U19764 (N_19764,N_17598,N_17591);
nor U19765 (N_19765,N_17993,N_17894);
or U19766 (N_19766,N_17895,N_17806);
or U19767 (N_19767,N_18078,N_17647);
and U19768 (N_19768,N_18161,N_18495);
xor U19769 (N_19769,N_18532,N_18231);
or U19770 (N_19770,N_18374,N_18068);
and U19771 (N_19771,N_18131,N_18421);
nor U19772 (N_19772,N_18575,N_18483);
or U19773 (N_19773,N_18524,N_18401);
nor U19774 (N_19774,N_17512,N_17790);
xnor U19775 (N_19775,N_17990,N_17833);
or U19776 (N_19776,N_17728,N_18064);
nand U19777 (N_19777,N_18218,N_18481);
nor U19778 (N_19778,N_18663,N_17593);
nand U19779 (N_19779,N_18252,N_18405);
and U19780 (N_19780,N_17599,N_18432);
nor U19781 (N_19781,N_17845,N_17807);
nand U19782 (N_19782,N_18271,N_17861);
or U19783 (N_19783,N_18126,N_17648);
and U19784 (N_19784,N_18443,N_17758);
and U19785 (N_19785,N_18185,N_18614);
and U19786 (N_19786,N_18124,N_17933);
and U19787 (N_19787,N_18484,N_18222);
xnor U19788 (N_19788,N_18610,N_17593);
nand U19789 (N_19789,N_18288,N_17814);
nand U19790 (N_19790,N_17745,N_17814);
nor U19791 (N_19791,N_18515,N_18412);
nand U19792 (N_19792,N_17558,N_17639);
or U19793 (N_19793,N_18466,N_18079);
and U19794 (N_19794,N_18221,N_17748);
nand U19795 (N_19795,N_17901,N_17845);
nand U19796 (N_19796,N_17747,N_18551);
nand U19797 (N_19797,N_18439,N_17790);
or U19798 (N_19798,N_17565,N_18383);
nand U19799 (N_19799,N_17610,N_17935);
or U19800 (N_19800,N_18699,N_18432);
or U19801 (N_19801,N_18724,N_17714);
xnor U19802 (N_19802,N_18011,N_17774);
nand U19803 (N_19803,N_18431,N_18590);
or U19804 (N_19804,N_18135,N_18157);
nand U19805 (N_19805,N_17985,N_18211);
or U19806 (N_19806,N_18382,N_17753);
or U19807 (N_19807,N_17936,N_18460);
nand U19808 (N_19808,N_17907,N_18381);
and U19809 (N_19809,N_18737,N_17558);
or U19810 (N_19810,N_18699,N_17612);
or U19811 (N_19811,N_18470,N_18269);
xor U19812 (N_19812,N_17994,N_17836);
nor U19813 (N_19813,N_18707,N_18129);
nand U19814 (N_19814,N_18439,N_18687);
and U19815 (N_19815,N_18235,N_17614);
or U19816 (N_19816,N_18222,N_18044);
xnor U19817 (N_19817,N_18316,N_17745);
or U19818 (N_19818,N_17526,N_18246);
nand U19819 (N_19819,N_17849,N_18190);
or U19820 (N_19820,N_18082,N_18268);
or U19821 (N_19821,N_17878,N_17868);
and U19822 (N_19822,N_18479,N_18651);
or U19823 (N_19823,N_18376,N_17696);
xnor U19824 (N_19824,N_17938,N_17867);
nor U19825 (N_19825,N_18384,N_17529);
xnor U19826 (N_19826,N_18344,N_18168);
nand U19827 (N_19827,N_18149,N_17970);
xor U19828 (N_19828,N_17753,N_17835);
and U19829 (N_19829,N_18430,N_18101);
or U19830 (N_19830,N_17824,N_18165);
and U19831 (N_19831,N_17770,N_17648);
nor U19832 (N_19832,N_17570,N_18661);
and U19833 (N_19833,N_18247,N_17991);
or U19834 (N_19834,N_18022,N_17728);
nand U19835 (N_19835,N_17627,N_18544);
xnor U19836 (N_19836,N_18243,N_17890);
and U19837 (N_19837,N_18196,N_18329);
nand U19838 (N_19838,N_17805,N_18705);
xor U19839 (N_19839,N_18686,N_18364);
nand U19840 (N_19840,N_18492,N_17973);
xor U19841 (N_19841,N_18532,N_18253);
or U19842 (N_19842,N_18526,N_18092);
nor U19843 (N_19843,N_17749,N_17939);
nand U19844 (N_19844,N_18709,N_18055);
xnor U19845 (N_19845,N_18467,N_18645);
xor U19846 (N_19846,N_17634,N_17654);
xor U19847 (N_19847,N_18267,N_18535);
or U19848 (N_19848,N_18285,N_18485);
or U19849 (N_19849,N_17850,N_17565);
xor U19850 (N_19850,N_17632,N_18115);
nand U19851 (N_19851,N_17944,N_18714);
or U19852 (N_19852,N_17635,N_17641);
xor U19853 (N_19853,N_18067,N_17872);
xnor U19854 (N_19854,N_17984,N_17951);
and U19855 (N_19855,N_18084,N_17869);
or U19856 (N_19856,N_17729,N_18358);
and U19857 (N_19857,N_17757,N_18288);
nand U19858 (N_19858,N_18348,N_18290);
and U19859 (N_19859,N_18171,N_17687);
or U19860 (N_19860,N_17851,N_18242);
xnor U19861 (N_19861,N_17707,N_18673);
and U19862 (N_19862,N_18339,N_17703);
nor U19863 (N_19863,N_17812,N_17637);
nand U19864 (N_19864,N_17709,N_18701);
or U19865 (N_19865,N_17528,N_17896);
and U19866 (N_19866,N_17940,N_18668);
nor U19867 (N_19867,N_17754,N_18381);
or U19868 (N_19868,N_17517,N_17819);
nor U19869 (N_19869,N_17590,N_18209);
or U19870 (N_19870,N_18462,N_17819);
xnor U19871 (N_19871,N_17632,N_18607);
nand U19872 (N_19872,N_18483,N_18262);
or U19873 (N_19873,N_17779,N_18612);
nand U19874 (N_19874,N_18316,N_17870);
nand U19875 (N_19875,N_18158,N_17836);
nor U19876 (N_19876,N_18100,N_18290);
xor U19877 (N_19877,N_17922,N_17826);
nor U19878 (N_19878,N_17585,N_17835);
and U19879 (N_19879,N_18018,N_18439);
or U19880 (N_19880,N_18513,N_17822);
nor U19881 (N_19881,N_17845,N_18575);
nor U19882 (N_19882,N_18174,N_17913);
and U19883 (N_19883,N_17663,N_17812);
xor U19884 (N_19884,N_18698,N_18660);
xnor U19885 (N_19885,N_17797,N_18335);
xor U19886 (N_19886,N_18454,N_18656);
and U19887 (N_19887,N_17739,N_18146);
nor U19888 (N_19888,N_17773,N_17956);
or U19889 (N_19889,N_18274,N_17609);
or U19890 (N_19890,N_18675,N_18727);
nor U19891 (N_19891,N_17909,N_17515);
nand U19892 (N_19892,N_17817,N_18604);
xnor U19893 (N_19893,N_18137,N_17964);
xor U19894 (N_19894,N_18286,N_17743);
xnor U19895 (N_19895,N_17835,N_17628);
xor U19896 (N_19896,N_18032,N_18500);
xnor U19897 (N_19897,N_18498,N_18277);
or U19898 (N_19898,N_18082,N_17799);
nor U19899 (N_19899,N_18455,N_18519);
or U19900 (N_19900,N_18126,N_18698);
and U19901 (N_19901,N_18410,N_17541);
nor U19902 (N_19902,N_18229,N_17531);
nand U19903 (N_19903,N_18445,N_18657);
nor U19904 (N_19904,N_18714,N_18254);
nor U19905 (N_19905,N_18277,N_17917);
or U19906 (N_19906,N_17661,N_18107);
or U19907 (N_19907,N_17602,N_18219);
nor U19908 (N_19908,N_17718,N_18611);
or U19909 (N_19909,N_18673,N_17858);
and U19910 (N_19910,N_18132,N_17981);
nand U19911 (N_19911,N_18278,N_18414);
and U19912 (N_19912,N_18264,N_17902);
or U19913 (N_19913,N_18316,N_18254);
xor U19914 (N_19914,N_17994,N_18576);
and U19915 (N_19915,N_18568,N_17609);
or U19916 (N_19916,N_18193,N_18605);
nor U19917 (N_19917,N_17835,N_17575);
and U19918 (N_19918,N_18749,N_17555);
nor U19919 (N_19919,N_17782,N_17922);
nor U19920 (N_19920,N_18686,N_18100);
xor U19921 (N_19921,N_17777,N_18586);
nand U19922 (N_19922,N_18348,N_18046);
xor U19923 (N_19923,N_18688,N_18309);
nand U19924 (N_19924,N_17593,N_18651);
and U19925 (N_19925,N_17801,N_17981);
or U19926 (N_19926,N_18635,N_17733);
and U19927 (N_19927,N_18171,N_18433);
nor U19928 (N_19928,N_18678,N_18399);
and U19929 (N_19929,N_18377,N_17784);
xnor U19930 (N_19930,N_17951,N_17802);
xnor U19931 (N_19931,N_17963,N_18239);
and U19932 (N_19932,N_17971,N_17819);
nand U19933 (N_19933,N_17638,N_18241);
or U19934 (N_19934,N_18183,N_18364);
or U19935 (N_19935,N_18438,N_17898);
nand U19936 (N_19936,N_18080,N_18596);
nand U19937 (N_19937,N_17599,N_17510);
xnor U19938 (N_19938,N_18709,N_18453);
nor U19939 (N_19939,N_17915,N_18700);
nor U19940 (N_19940,N_17575,N_18473);
xnor U19941 (N_19941,N_18549,N_17917);
xnor U19942 (N_19942,N_18037,N_17835);
nor U19943 (N_19943,N_17705,N_18704);
or U19944 (N_19944,N_17726,N_18265);
or U19945 (N_19945,N_17928,N_18485);
nand U19946 (N_19946,N_17914,N_18294);
xnor U19947 (N_19947,N_17664,N_17730);
or U19948 (N_19948,N_17748,N_18394);
and U19949 (N_19949,N_18589,N_17952);
or U19950 (N_19950,N_18053,N_17771);
and U19951 (N_19951,N_17637,N_18165);
or U19952 (N_19952,N_17897,N_18740);
nand U19953 (N_19953,N_18293,N_18608);
xor U19954 (N_19954,N_18485,N_17581);
and U19955 (N_19955,N_18599,N_18033);
and U19956 (N_19956,N_17811,N_17580);
nand U19957 (N_19957,N_18364,N_18414);
nor U19958 (N_19958,N_18358,N_18274);
xnor U19959 (N_19959,N_18693,N_18634);
nand U19960 (N_19960,N_17555,N_18003);
xnor U19961 (N_19961,N_17662,N_17729);
nor U19962 (N_19962,N_18534,N_18347);
xor U19963 (N_19963,N_18619,N_18452);
or U19964 (N_19964,N_18437,N_18278);
nor U19965 (N_19965,N_18367,N_17527);
nor U19966 (N_19966,N_18003,N_18329);
nand U19967 (N_19967,N_17656,N_18405);
and U19968 (N_19968,N_17872,N_17933);
xor U19969 (N_19969,N_17529,N_18242);
xor U19970 (N_19970,N_17562,N_17842);
nand U19971 (N_19971,N_17599,N_18365);
or U19972 (N_19972,N_17575,N_18073);
nor U19973 (N_19973,N_17622,N_18136);
and U19974 (N_19974,N_17996,N_18610);
or U19975 (N_19975,N_18294,N_18479);
nand U19976 (N_19976,N_18172,N_18630);
nor U19977 (N_19977,N_18646,N_18645);
nor U19978 (N_19978,N_17806,N_18076);
nand U19979 (N_19979,N_18372,N_18160);
nor U19980 (N_19980,N_18461,N_18434);
or U19981 (N_19981,N_17997,N_17607);
or U19982 (N_19982,N_17748,N_17994);
nor U19983 (N_19983,N_17871,N_17549);
or U19984 (N_19984,N_17550,N_18297);
xor U19985 (N_19985,N_18542,N_17957);
nor U19986 (N_19986,N_18348,N_17645);
xnor U19987 (N_19987,N_18072,N_18722);
nor U19988 (N_19988,N_17921,N_17942);
and U19989 (N_19989,N_17961,N_17938);
and U19990 (N_19990,N_17717,N_18679);
nand U19991 (N_19991,N_18472,N_17558);
and U19992 (N_19992,N_17554,N_17587);
and U19993 (N_19993,N_18493,N_17784);
nor U19994 (N_19994,N_18532,N_18088);
or U19995 (N_19995,N_17675,N_18504);
nand U19996 (N_19996,N_18561,N_18668);
and U19997 (N_19997,N_18687,N_17579);
nand U19998 (N_19998,N_18657,N_18404);
nor U19999 (N_19999,N_18155,N_17566);
or U20000 (N_20000,N_18853,N_19060);
and U20001 (N_20001,N_19829,N_18793);
xnor U20002 (N_20002,N_19814,N_19057);
nand U20003 (N_20003,N_19601,N_19744);
and U20004 (N_20004,N_19243,N_19447);
nor U20005 (N_20005,N_18760,N_19026);
nand U20006 (N_20006,N_19086,N_19401);
xnor U20007 (N_20007,N_18951,N_19083);
or U20008 (N_20008,N_19976,N_18885);
nand U20009 (N_20009,N_19492,N_19300);
xor U20010 (N_20010,N_19217,N_18815);
and U20011 (N_20011,N_19790,N_19600);
and U20012 (N_20012,N_19761,N_18971);
xor U20013 (N_20013,N_18854,N_19099);
or U20014 (N_20014,N_19091,N_19347);
xor U20015 (N_20015,N_19048,N_19452);
and U20016 (N_20016,N_19713,N_19552);
and U20017 (N_20017,N_18917,N_19621);
or U20018 (N_20018,N_19226,N_19515);
xnor U20019 (N_20019,N_18993,N_19111);
and U20020 (N_20020,N_19567,N_19671);
nor U20021 (N_20021,N_18758,N_19782);
and U20022 (N_20022,N_19274,N_19440);
or U20023 (N_20023,N_18829,N_19075);
nor U20024 (N_20024,N_19130,N_19542);
xnor U20025 (N_20025,N_19895,N_19908);
xor U20026 (N_20026,N_19649,N_19246);
or U20027 (N_20027,N_18870,N_18860);
nor U20028 (N_20028,N_19381,N_18952);
nor U20029 (N_20029,N_19741,N_19002);
or U20030 (N_20030,N_19162,N_18765);
and U20031 (N_20031,N_19667,N_19623);
xnor U20032 (N_20032,N_19509,N_19974);
nor U20033 (N_20033,N_19449,N_19993);
and U20034 (N_20034,N_19033,N_19052);
nand U20035 (N_20035,N_18929,N_19205);
xor U20036 (N_20036,N_19996,N_19535);
nor U20037 (N_20037,N_19998,N_19475);
xor U20038 (N_20038,N_19686,N_19405);
xor U20039 (N_20039,N_19166,N_19143);
and U20040 (N_20040,N_19982,N_19295);
or U20041 (N_20041,N_19896,N_19353);
nor U20042 (N_20042,N_19015,N_19851);
nor U20043 (N_20043,N_19954,N_19408);
or U20044 (N_20044,N_19210,N_19241);
or U20045 (N_20045,N_19602,N_19670);
and U20046 (N_20046,N_19138,N_19916);
or U20047 (N_20047,N_19659,N_18974);
nand U20048 (N_20048,N_19548,N_19283);
nor U20049 (N_20049,N_19731,N_19424);
nand U20050 (N_20050,N_19822,N_19160);
nand U20051 (N_20051,N_18784,N_18832);
or U20052 (N_20052,N_18944,N_18934);
and U20053 (N_20053,N_19796,N_19286);
or U20054 (N_20054,N_19047,N_18812);
and U20055 (N_20055,N_19745,N_19718);
nor U20056 (N_20056,N_19619,N_19069);
and U20057 (N_20057,N_19081,N_19827);
nor U20058 (N_20058,N_18798,N_19315);
xnor U20059 (N_20059,N_19904,N_19333);
xnor U20060 (N_20060,N_19643,N_19929);
xnor U20061 (N_20061,N_19931,N_18897);
and U20062 (N_20062,N_18777,N_19986);
and U20063 (N_20063,N_18789,N_18814);
xnor U20064 (N_20064,N_19197,N_19359);
xnor U20065 (N_20065,N_19953,N_19488);
or U20066 (N_20066,N_19324,N_19082);
nand U20067 (N_20067,N_19969,N_19934);
nor U20068 (N_20068,N_18809,N_19618);
or U20069 (N_20069,N_19590,N_19693);
nand U20070 (N_20070,N_19648,N_19748);
nand U20071 (N_20071,N_19787,N_19174);
and U20072 (N_20072,N_19821,N_19287);
xor U20073 (N_20073,N_19681,N_19470);
nand U20074 (N_20074,N_19736,N_19971);
xor U20075 (N_20075,N_19041,N_19946);
xnor U20076 (N_20076,N_19311,N_19863);
xnor U20077 (N_20077,N_18799,N_19094);
or U20078 (N_20078,N_18880,N_18878);
nand U20079 (N_20079,N_19914,N_19249);
xor U20080 (N_20080,N_19282,N_19533);
nor U20081 (N_20081,N_19239,N_19750);
nor U20082 (N_20082,N_19545,N_19296);
nand U20083 (N_20083,N_19753,N_19493);
xnor U20084 (N_20084,N_19635,N_19624);
or U20085 (N_20085,N_19029,N_19421);
and U20086 (N_20086,N_18973,N_19156);
nor U20087 (N_20087,N_19317,N_19939);
or U20088 (N_20088,N_19800,N_19293);
or U20089 (N_20089,N_18816,N_19222);
nand U20090 (N_20090,N_18902,N_19572);
and U20091 (N_20091,N_18856,N_19525);
and U20092 (N_20092,N_19819,N_18879);
xnor U20093 (N_20093,N_18997,N_19778);
nor U20094 (N_20094,N_19633,N_19377);
nor U20095 (N_20095,N_19740,N_19306);
nand U20096 (N_20096,N_18752,N_19154);
or U20097 (N_20097,N_19593,N_19661);
nor U20098 (N_20098,N_19785,N_18800);
and U20099 (N_20099,N_19224,N_19251);
xnor U20100 (N_20100,N_18811,N_19588);
nor U20101 (N_20101,N_19812,N_19944);
or U20102 (N_20102,N_19716,N_18764);
nor U20103 (N_20103,N_18767,N_19540);
nand U20104 (N_20104,N_19173,N_19897);
nor U20105 (N_20105,N_19276,N_19764);
nand U20106 (N_20106,N_19644,N_19958);
or U20107 (N_20107,N_19067,N_19385);
and U20108 (N_20108,N_19983,N_19115);
nand U20109 (N_20109,N_19049,N_19290);
or U20110 (N_20110,N_19503,N_19878);
nand U20111 (N_20111,N_19597,N_18762);
or U20112 (N_20112,N_19232,N_19402);
and U20113 (N_20113,N_18754,N_19445);
xnor U20114 (N_20114,N_19909,N_19096);
xor U20115 (N_20115,N_19411,N_18808);
nand U20116 (N_20116,N_19071,N_19990);
nor U20117 (N_20117,N_18850,N_19495);
xor U20118 (N_20118,N_19614,N_18913);
nand U20119 (N_20119,N_19936,N_18957);
and U20120 (N_20120,N_19114,N_19415);
nand U20121 (N_20121,N_19769,N_19746);
and U20122 (N_20122,N_19992,N_19979);
xnor U20123 (N_20123,N_19959,N_19265);
nand U20124 (N_20124,N_19781,N_19184);
or U20125 (N_20125,N_19834,N_19964);
nand U20126 (N_20126,N_19512,N_19948);
and U20127 (N_20127,N_19794,N_18955);
nand U20128 (N_20128,N_18969,N_19702);
nor U20129 (N_20129,N_19279,N_19087);
or U20130 (N_20130,N_19857,N_18932);
and U20131 (N_20131,N_19608,N_18940);
or U20132 (N_20132,N_19361,N_18939);
and U20133 (N_20133,N_18999,N_18865);
or U20134 (N_20134,N_19541,N_19483);
xnor U20135 (N_20135,N_19104,N_18889);
nand U20136 (N_20136,N_18887,N_19108);
and U20137 (N_20137,N_19373,N_19346);
nor U20138 (N_20138,N_19676,N_19984);
or U20139 (N_20139,N_18986,N_19978);
xor U20140 (N_20140,N_19610,N_18837);
nor U20141 (N_20141,N_19795,N_19259);
and U20142 (N_20142,N_19714,N_19862);
nor U20143 (N_20143,N_19097,N_19388);
nor U20144 (N_20144,N_19288,N_19137);
xnor U20145 (N_20145,N_19549,N_19009);
or U20146 (N_20146,N_19132,N_19013);
and U20147 (N_20147,N_19507,N_19064);
nand U20148 (N_20148,N_19870,N_19309);
or U20149 (N_20149,N_19650,N_19529);
and U20150 (N_20150,N_19640,N_19923);
xor U20151 (N_20151,N_19678,N_18864);
and U20152 (N_20152,N_19005,N_19054);
nor U20153 (N_20153,N_19085,N_18948);
xnor U20154 (N_20154,N_19941,N_19392);
and U20155 (N_20155,N_18991,N_19077);
and U20156 (N_20156,N_19574,N_19236);
and U20157 (N_20157,N_19023,N_19190);
or U20158 (N_20158,N_18847,N_19144);
nor U20159 (N_20159,N_19065,N_19281);
or U20160 (N_20160,N_18761,N_19647);
or U20161 (N_20161,N_19471,N_19182);
xor U20162 (N_20162,N_19758,N_19596);
and U20163 (N_20163,N_19364,N_19806);
nand U20164 (N_20164,N_19124,N_19587);
nor U20165 (N_20165,N_18757,N_18906);
and U20166 (N_20166,N_19799,N_18968);
xnor U20167 (N_20167,N_19839,N_19318);
nor U20168 (N_20168,N_18891,N_19489);
and U20169 (N_20169,N_19943,N_19269);
xor U20170 (N_20170,N_19968,N_19845);
nor U20171 (N_20171,N_19792,N_19204);
xnor U20172 (N_20172,N_19700,N_19701);
nor U20173 (N_20173,N_19774,N_18768);
nor U20174 (N_20174,N_19188,N_19739);
nor U20175 (N_20175,N_19335,N_18892);
or U20176 (N_20176,N_19890,N_19776);
or U20177 (N_20177,N_19207,N_19429);
nand U20178 (N_20178,N_19807,N_19975);
nand U20179 (N_20179,N_19842,N_18791);
or U20180 (N_20180,N_19285,N_18920);
and U20181 (N_20181,N_19294,N_19977);
nor U20182 (N_20182,N_19938,N_19654);
nand U20183 (N_20183,N_19187,N_19876);
and U20184 (N_20184,N_18872,N_18774);
nand U20185 (N_20185,N_19757,N_19692);
or U20186 (N_20186,N_19734,N_19727);
and U20187 (N_20187,N_19422,N_18964);
xor U20188 (N_20188,N_19487,N_19828);
nand U20189 (N_20189,N_19391,N_19902);
and U20190 (N_20190,N_19109,N_19398);
or U20191 (N_20191,N_19846,N_19140);
xor U20192 (N_20192,N_19418,N_18942);
and U20193 (N_20193,N_19245,N_19950);
xnor U20194 (N_20194,N_19028,N_19666);
nor U20195 (N_20195,N_19672,N_19456);
or U20196 (N_20196,N_19024,N_19328);
nand U20197 (N_20197,N_19711,N_19849);
nand U20198 (N_20198,N_19254,N_18867);
and U20199 (N_20199,N_19079,N_19380);
or U20200 (N_20200,N_19835,N_18950);
nand U20201 (N_20201,N_18894,N_19859);
and U20202 (N_20202,N_19133,N_18831);
xor U20203 (N_20203,N_19646,N_19510);
xnor U20204 (N_20204,N_19406,N_19523);
or U20205 (N_20205,N_19004,N_19036);
and U20206 (N_20206,N_19712,N_19342);
nand U20207 (N_20207,N_18898,N_19688);
and U20208 (N_20208,N_18849,N_19988);
nor U20209 (N_20209,N_19728,N_19848);
xnor U20210 (N_20210,N_19877,N_19486);
xnor U20211 (N_20211,N_19159,N_19961);
or U20212 (N_20212,N_19611,N_19334);
nand U20213 (N_20213,N_19165,N_18810);
nand U20214 (N_20214,N_19001,N_19066);
nor U20215 (N_20215,N_19524,N_19343);
or U20216 (N_20216,N_19536,N_18937);
nor U20217 (N_20217,N_19505,N_19061);
nor U20218 (N_20218,N_19354,N_19003);
nand U20219 (N_20219,N_19201,N_19497);
xnor U20220 (N_20220,N_19658,N_19312);
or U20221 (N_20221,N_19366,N_18817);
xor U20222 (N_20222,N_19725,N_19823);
nand U20223 (N_20223,N_19501,N_18928);
nor U20224 (N_20224,N_19238,N_19802);
nand U20225 (N_20225,N_19885,N_19291);
xor U20226 (N_20226,N_18982,N_19617);
nand U20227 (N_20227,N_19779,N_19092);
xor U20228 (N_20228,N_19363,N_19526);
nand U20229 (N_20229,N_19256,N_19737);
xnor U20230 (N_20230,N_19894,N_19039);
xor U20231 (N_20231,N_19338,N_19609);
nand U20232 (N_20232,N_19442,N_19050);
nand U20233 (N_20233,N_19168,N_18844);
nor U20234 (N_20234,N_19074,N_19818);
or U20235 (N_20235,N_19213,N_19194);
or U20236 (N_20236,N_19632,N_18763);
or U20237 (N_20237,N_19231,N_19784);
nor U20238 (N_20238,N_19559,N_19462);
nand U20239 (N_20239,N_19485,N_19551);
xor U20240 (N_20240,N_18954,N_18876);
and U20241 (N_20241,N_19668,N_19298);
and U20242 (N_20242,N_19738,N_19577);
and U20243 (N_20243,N_19682,N_19255);
or U20244 (N_20244,N_19917,N_19258);
xnor U20245 (N_20245,N_19145,N_19120);
nand U20246 (N_20246,N_18984,N_19762);
and U20247 (N_20247,N_19856,N_18908);
and U20248 (N_20248,N_19339,N_19119);
nand U20249 (N_20249,N_19479,N_19062);
and U20250 (N_20250,N_19833,N_19579);
nor U20251 (N_20251,N_19584,N_19230);
xnor U20252 (N_20252,N_19791,N_19933);
nand U20253 (N_20253,N_19652,N_19694);
nand U20254 (N_20254,N_18794,N_18750);
or U20255 (N_20255,N_19777,N_19451);
or U20256 (N_20256,N_19473,N_19019);
and U20257 (N_20257,N_18755,N_19244);
xor U20258 (N_20258,N_19257,N_19152);
or U20259 (N_20259,N_19208,N_19356);
xnor U20260 (N_20260,N_19301,N_19307);
and U20261 (N_20261,N_19164,N_19220);
nor U20262 (N_20262,N_19123,N_19808);
nand U20263 (N_20263,N_19726,N_18900);
xnor U20264 (N_20264,N_19893,N_19271);
nor U20265 (N_20265,N_19357,N_19742);
xnor U20266 (N_20266,N_19696,N_19056);
nand U20267 (N_20267,N_19825,N_19305);
and U20268 (N_20268,N_18949,N_19468);
or U20269 (N_20269,N_19582,N_18873);
or U20270 (N_20270,N_19922,N_19997);
nor U20271 (N_20271,N_19967,N_19443);
or U20272 (N_20272,N_19527,N_19185);
or U20273 (N_20273,N_18820,N_19289);
xnor U20274 (N_20274,N_19637,N_18890);
and U20275 (N_20275,N_19815,N_19889);
xnor U20276 (N_20276,N_18852,N_19566);
and U20277 (N_20277,N_19481,N_19556);
xor U20278 (N_20278,N_19474,N_19035);
nand U20279 (N_20279,N_19561,N_19397);
nand U20280 (N_20280,N_19565,N_18781);
nand U20281 (N_20281,N_19490,N_18838);
xnor U20282 (N_20282,N_18888,N_19040);
and U20283 (N_20283,N_19107,N_19102);
nand U20284 (N_20284,N_19053,N_19240);
or U20285 (N_20285,N_19826,N_19698);
nand U20286 (N_20286,N_19801,N_19368);
nand U20287 (N_20287,N_19464,N_19158);
and U20288 (N_20288,N_18845,N_18963);
or U20289 (N_20289,N_19273,N_18782);
xnor U20290 (N_20290,N_19011,N_19196);
xnor U20291 (N_20291,N_19463,N_19832);
nor U20292 (N_20292,N_19662,N_19389);
nor U20293 (N_20293,N_19117,N_18893);
or U20294 (N_20294,N_19598,N_19554);
nor U20295 (N_20295,N_19962,N_19683);
or U20296 (N_20296,N_19200,N_18786);
nor U20297 (N_20297,N_19433,N_19674);
or U20298 (N_20298,N_19118,N_19370);
nor U20299 (N_20299,N_19730,N_19543);
and U20300 (N_20300,N_19817,N_19297);
nand U20301 (N_20301,N_19687,N_18967);
nand U20302 (N_20302,N_19735,N_18881);
nand U20303 (N_20303,N_18927,N_19076);
nor U20304 (N_20304,N_18821,N_19477);
or U20305 (N_20305,N_18877,N_19871);
nor U20306 (N_20306,N_19417,N_19592);
nand U20307 (N_20307,N_19573,N_19260);
nand U20308 (N_20308,N_18995,N_19454);
or U20309 (N_20309,N_19715,N_19058);
and U20310 (N_20310,N_19136,N_19629);
and U20311 (N_20311,N_19034,N_18805);
xor U20312 (N_20312,N_19613,N_19199);
xor U20313 (N_20313,N_19498,N_19410);
or U20314 (N_20314,N_19907,N_19126);
and U20315 (N_20315,N_18988,N_19660);
and U20316 (N_20316,N_18976,N_19177);
xor U20317 (N_20317,N_19759,N_19743);
or U20318 (N_20318,N_19645,N_19995);
or U20319 (N_20319,N_19263,N_18922);
xnor U20320 (N_20320,N_19547,N_19513);
xnor U20321 (N_20321,N_19765,N_19396);
xor U20322 (N_20322,N_19824,N_18787);
nand U20323 (N_20323,N_19134,N_19191);
nor U20324 (N_20324,N_19991,N_18992);
xnor U20325 (N_20325,N_19973,N_19499);
and U20326 (N_20326,N_19706,N_19223);
or U20327 (N_20327,N_19027,N_19811);
nand U20328 (N_20328,N_19775,N_19721);
nand U20329 (N_20329,N_19112,N_19310);
and U20330 (N_20330,N_19416,N_19070);
or U20331 (N_20331,N_19772,N_19837);
nor U20332 (N_20332,N_19038,N_19369);
nand U20333 (N_20333,N_19450,N_19516);
or U20334 (N_20334,N_19980,N_19903);
and U20335 (N_20335,N_19684,N_18980);
or U20336 (N_20336,N_18771,N_18945);
xor U20337 (N_20337,N_19864,N_19446);
nor U20338 (N_20338,N_19733,N_19435);
or U20339 (N_20339,N_19448,N_19494);
and U20340 (N_20340,N_19330,N_19163);
nand U20341 (N_20341,N_18911,N_19006);
nor U20342 (N_20342,N_19403,N_19749);
xor U20343 (N_20343,N_19578,N_19927);
nand U20344 (N_20344,N_19280,N_19030);
or U20345 (N_20345,N_18835,N_19724);
xor U20346 (N_20346,N_18874,N_19703);
or U20347 (N_20347,N_19237,N_19816);
nand U20348 (N_20348,N_18827,N_18983);
or U20349 (N_20349,N_19267,N_19155);
or U20350 (N_20350,N_19341,N_19560);
xnor U20351 (N_20351,N_18904,N_19098);
or U20352 (N_20352,N_18778,N_19920);
nor U20353 (N_20353,N_19399,N_18943);
nor U20354 (N_20354,N_19690,N_19277);
nor U20355 (N_20355,N_19482,N_19371);
and U20356 (N_20356,N_18966,N_19689);
nor U20357 (N_20357,N_19860,N_18851);
nor U20358 (N_20358,N_19899,N_19639);
and U20359 (N_20359,N_19045,N_19657);
and U20360 (N_20360,N_19921,N_18962);
and U20361 (N_20361,N_18825,N_19010);
and U20362 (N_20362,N_18961,N_19225);
nor U20363 (N_20363,N_19461,N_19453);
and U20364 (N_20364,N_19100,N_19212);
xnor U20365 (N_20365,N_18915,N_19221);
nor U20366 (N_20366,N_19880,N_19534);
or U20367 (N_20367,N_19576,N_18753);
nand U20368 (N_20368,N_19502,N_19374);
and U20369 (N_20369,N_19585,N_19467);
nor U20370 (N_20370,N_18818,N_19372);
or U20371 (N_20371,N_19760,N_19375);
xor U20372 (N_20372,N_19874,N_19626);
xor U20373 (N_20373,N_19379,N_18916);
xor U20374 (N_20374,N_19472,N_19868);
or U20375 (N_20375,N_19439,N_18795);
nand U20376 (N_20376,N_19882,N_19570);
or U20377 (N_20377,N_19321,N_18965);
xor U20378 (N_20378,N_19088,N_19272);
xnor U20379 (N_20379,N_19981,N_19250);
xnor U20380 (N_20380,N_19836,N_18766);
nand U20381 (N_20381,N_19031,N_19970);
nor U20382 (N_20382,N_19669,N_18822);
or U20383 (N_20383,N_19723,N_19193);
or U20384 (N_20384,N_19999,N_19506);
or U20385 (N_20385,N_19072,N_18947);
and U20386 (N_20386,N_19571,N_18823);
or U20387 (N_20387,N_19393,N_19768);
or U20388 (N_20388,N_19940,N_19419);
and U20389 (N_20389,N_19875,N_18776);
or U20390 (N_20390,N_19089,N_19586);
xnor U20391 (N_20391,N_18836,N_18978);
nor U20392 (N_20392,N_19051,N_19518);
nand U20393 (N_20393,N_19809,N_19478);
nor U20394 (N_20394,N_19150,N_18796);
nand U20395 (N_20395,N_18979,N_18770);
nand U20396 (N_20396,N_19007,N_19705);
nand U20397 (N_20397,N_19055,N_19046);
and U20398 (N_20398,N_18803,N_19407);
nor U20399 (N_20399,N_18910,N_18855);
nor U20400 (N_20400,N_18959,N_19021);
nor U20401 (N_20401,N_19323,N_19020);
xor U20402 (N_20402,N_18958,N_19084);
nand U20403 (N_20403,N_19355,N_19722);
xnor U20404 (N_20404,N_19211,N_19583);
nand U20405 (N_20405,N_19638,N_19131);
or U20406 (N_20406,N_19413,N_19459);
nor U20407 (N_20407,N_19500,N_19951);
nor U20408 (N_20408,N_19891,N_19017);
nand U20409 (N_20409,N_19496,N_19351);
nor U20410 (N_20410,N_19717,N_19063);
nor U20411 (N_20411,N_19767,N_18804);
xnor U20412 (N_20412,N_19925,N_19195);
xor U20413 (N_20413,N_18819,N_18790);
nor U20414 (N_20414,N_19409,N_19830);
nor U20415 (N_20415,N_18918,N_19563);
and U20416 (N_20416,N_19892,N_18862);
xor U20417 (N_20417,N_18909,N_19386);
or U20418 (N_20418,N_19169,N_19581);
or U20419 (N_20419,N_19989,N_19180);
and U20420 (N_20420,N_19532,N_19268);
nor U20421 (N_20421,N_18833,N_19665);
or U20422 (N_20422,N_19455,N_19345);
nor U20423 (N_20423,N_19956,N_19378);
and U20424 (N_20424,N_19438,N_19437);
and U20425 (N_20425,N_19008,N_19865);
and U20426 (N_20426,N_19810,N_19151);
nand U20427 (N_20427,N_19022,N_19412);
and U20428 (N_20428,N_19589,N_18884);
nor U20429 (N_20429,N_19362,N_19831);
nor U20430 (N_20430,N_19171,N_19766);
nand U20431 (N_20431,N_19642,N_18806);
or U20432 (N_20432,N_19235,N_19469);
xor U20433 (N_20433,N_18807,N_19068);
nor U20434 (N_20434,N_19302,N_19604);
or U20435 (N_20435,N_19930,N_19358);
or U20436 (N_20436,N_18858,N_19558);
or U20437 (N_20437,N_19519,N_19770);
nor U20438 (N_20438,N_19480,N_19270);
nor U20439 (N_20439,N_19014,N_19325);
nor U20440 (N_20440,N_18756,N_19414);
nand U20441 (N_20441,N_19059,N_19663);
or U20442 (N_20442,N_18769,N_19018);
and U20443 (N_20443,N_19420,N_19395);
xor U20444 (N_20444,N_19919,N_19966);
or U20445 (N_20445,N_19476,N_19209);
and U20446 (N_20446,N_19400,N_19116);
nand U20447 (N_20447,N_19139,N_19595);
and U20448 (N_20448,N_19841,N_19928);
nor U20449 (N_20449,N_19153,N_19755);
and U20450 (N_20450,N_19322,N_19044);
or U20451 (N_20451,N_19537,N_19569);
nor U20452 (N_20452,N_19508,N_18924);
nand U20453 (N_20453,N_18826,N_19539);
or U20454 (N_20454,N_19331,N_18780);
or U20455 (N_20455,N_19128,N_19955);
nor U20456 (N_20456,N_19853,N_19350);
nor U20457 (N_20457,N_19677,N_19248);
or U20458 (N_20458,N_19348,N_18960);
nor U20459 (N_20459,N_19465,N_19599);
and U20460 (N_20460,N_19910,N_19219);
nand U20461 (N_20461,N_19215,N_18751);
xor U20462 (N_20462,N_19387,N_19016);
nor U20463 (N_20463,N_19316,N_19763);
and U20464 (N_20464,N_19491,N_19078);
nand U20465 (N_20465,N_19945,N_18759);
xnor U20466 (N_20466,N_19292,N_18846);
nand U20467 (N_20467,N_18834,N_19175);
nor U20468 (N_20468,N_19425,N_19783);
and U20469 (N_20469,N_18921,N_19216);
and U20470 (N_20470,N_19866,N_19773);
xnor U20471 (N_20471,N_19679,N_19844);
xor U20472 (N_20472,N_19729,N_19798);
nand U20473 (N_20473,N_19025,N_19101);
nor U20474 (N_20474,N_19987,N_19607);
nor U20475 (N_20475,N_19704,N_18866);
and U20476 (N_20476,N_19651,N_19858);
xnor U20477 (N_20477,N_19653,N_18895);
xnor U20478 (N_20478,N_19924,N_19697);
or U20479 (N_20479,N_19308,N_18785);
nand U20480 (N_20480,N_19553,N_19206);
and U20481 (N_20481,N_19756,N_19575);
or U20482 (N_20482,N_19262,N_19555);
nor U20483 (N_20483,N_19879,N_18886);
and U20484 (N_20484,N_19105,N_18848);
and U20485 (N_20485,N_18926,N_19546);
nand U20486 (N_20486,N_19229,N_18863);
nor U20487 (N_20487,N_19843,N_19458);
nor U20488 (N_20488,N_19847,N_19432);
xnor U20489 (N_20489,N_18996,N_18987);
nand U20490 (N_20490,N_19428,N_19630);
or U20491 (N_20491,N_19771,N_18938);
and U20492 (N_20492,N_19404,N_19867);
nor U20493 (N_20493,N_19352,N_19441);
nor U20494 (N_20494,N_19932,N_19313);
and U20495 (N_20495,N_18936,N_19531);
or U20496 (N_20496,N_19580,N_19113);
nor U20497 (N_20497,N_19228,N_18871);
nand U20498 (N_20498,N_19183,N_19935);
nor U20499 (N_20499,N_19142,N_19234);
nor U20500 (N_20500,N_19304,N_19179);
nand U20501 (N_20501,N_18931,N_19710);
nor U20502 (N_20502,N_18868,N_18901);
or U20503 (N_20503,N_18998,N_19685);
and U20504 (N_20504,N_19484,N_19320);
nand U20505 (N_20505,N_18946,N_19786);
xor U20506 (N_20506,N_19382,N_19591);
and U20507 (N_20507,N_19135,N_19360);
or U20508 (N_20508,N_19985,N_19616);
nor U20509 (N_20509,N_19247,N_19170);
or U20510 (N_20510,N_19838,N_19383);
xor U20511 (N_20511,N_19918,N_19275);
or U20512 (N_20512,N_19699,N_19965);
xor U20513 (N_20513,N_19957,N_19627);
nand U20514 (N_20514,N_19708,N_19073);
or U20515 (N_20515,N_19852,N_18923);
xor U20516 (N_20516,N_19314,N_19218);
or U20517 (N_20517,N_19625,N_18933);
and U20518 (N_20518,N_18907,N_18775);
nor U20519 (N_20519,N_18985,N_18783);
xnor U20520 (N_20520,N_18839,N_19511);
and U20521 (N_20521,N_19430,N_19202);
nor U20522 (N_20522,N_19544,N_19720);
nor U20523 (N_20523,N_19000,N_19037);
xnor U20524 (N_20524,N_19884,N_19615);
or U20525 (N_20525,N_19913,N_19203);
nor U20526 (N_20526,N_19517,N_19905);
or U20527 (N_20527,N_19106,N_19192);
xor U20528 (N_20528,N_19337,N_18841);
xnor U20529 (N_20529,N_18912,N_19901);
xnor U20530 (N_20530,N_19594,N_19628);
or U20531 (N_20531,N_18972,N_19780);
and U20532 (N_20532,N_18843,N_19797);
and U20533 (N_20533,N_18925,N_18981);
xnor U20534 (N_20534,N_19125,N_19198);
nand U20535 (N_20535,N_19804,N_19947);
and U20536 (N_20536,N_19167,N_19504);
xnor U20537 (N_20537,N_19095,N_19656);
nor U20538 (N_20538,N_19127,N_19227);
and U20539 (N_20539,N_18990,N_19568);
nor U20540 (N_20540,N_19675,N_19803);
nor U20541 (N_20541,N_19641,N_18773);
and U20542 (N_20542,N_18861,N_19178);
or U20543 (N_20543,N_19390,N_19336);
or U20544 (N_20544,N_19898,N_19911);
xor U20545 (N_20545,N_19789,N_19906);
nor U20546 (N_20546,N_19854,N_19186);
and U20547 (N_20547,N_19915,N_19326);
xor U20548 (N_20548,N_18919,N_19883);
and U20549 (N_20549,N_18956,N_19299);
nand U20550 (N_20550,N_19319,N_19960);
xor U20551 (N_20551,N_19886,N_19603);
xor U20552 (N_20552,N_18830,N_19752);
and U20553 (N_20553,N_18989,N_19521);
xor U20554 (N_20554,N_19994,N_19861);
nand U20555 (N_20555,N_19528,N_19181);
xnor U20556 (N_20556,N_19457,N_19655);
nand U20557 (N_20557,N_19278,N_19103);
nand U20558 (N_20558,N_19252,N_19367);
and U20559 (N_20559,N_19426,N_19444);
and U20560 (N_20560,N_19538,N_19754);
xor U20561 (N_20561,N_19942,N_19284);
nand U20562 (N_20562,N_19840,N_19242);
or U20563 (N_20563,N_19751,N_18797);
and U20564 (N_20564,N_18813,N_19673);
nand U20565 (N_20565,N_19732,N_19562);
and U20566 (N_20566,N_18772,N_19466);
nand U20567 (N_20567,N_19952,N_18896);
nand U20568 (N_20568,N_18914,N_19620);
xnor U20569 (N_20569,N_19172,N_19926);
nand U20570 (N_20570,N_19520,N_18905);
or U20571 (N_20571,N_19080,N_18970);
nor U20572 (N_20572,N_18788,N_19937);
or U20573 (N_20573,N_19664,N_19376);
nor U20574 (N_20574,N_19122,N_19365);
xnor U20575 (N_20575,N_19680,N_19963);
or U20576 (N_20576,N_18859,N_19329);
nand U20577 (N_20577,N_19149,N_19161);
or U20578 (N_20578,N_19394,N_19636);
nand U20579 (N_20579,N_18801,N_18828);
xnor U20580 (N_20580,N_19850,N_19522);
or U20581 (N_20581,N_18883,N_19912);
nand U20582 (N_20582,N_18977,N_19189);
and U20583 (N_20583,N_18953,N_19261);
and U20584 (N_20584,N_19253,N_19820);
nor U20585 (N_20585,N_19550,N_19514);
xor U20586 (N_20586,N_19093,N_18903);
xnor U20587 (N_20587,N_18824,N_19032);
and U20588 (N_20588,N_19427,N_19042);
nor U20589 (N_20589,N_19631,N_19233);
and U20590 (N_20590,N_19043,N_19605);
or U20591 (N_20591,N_19530,N_19327);
nand U20592 (N_20592,N_19121,N_19012);
nor U20593 (N_20593,N_19813,N_18975);
nand U20594 (N_20594,N_19634,N_18869);
and U20595 (N_20595,N_19129,N_19090);
nor U20596 (N_20596,N_19264,N_19881);
nand U20597 (N_20597,N_19423,N_19460);
nor U20598 (N_20598,N_19146,N_19972);
nand U20599 (N_20599,N_19793,N_18994);
xor U20600 (N_20600,N_18930,N_19707);
and U20601 (N_20601,N_18779,N_19873);
xnor U20602 (N_20602,N_18802,N_19434);
or U20603 (N_20603,N_19332,N_19157);
or U20604 (N_20604,N_19805,N_19266);
nor U20605 (N_20605,N_19872,N_19888);
and U20606 (N_20606,N_18935,N_19436);
and U20607 (N_20607,N_19695,N_18882);
or U20608 (N_20608,N_19340,N_19612);
nor U20609 (N_20609,N_19691,N_19349);
nor U20610 (N_20610,N_19176,N_19557);
and U20611 (N_20611,N_18899,N_19384);
or U20612 (N_20612,N_19214,N_19431);
nand U20613 (N_20613,N_19788,N_19110);
nand U20614 (N_20614,N_19564,N_18792);
or U20615 (N_20615,N_19719,N_19344);
xor U20616 (N_20616,N_19148,N_19141);
or U20617 (N_20617,N_18857,N_19303);
xor U20618 (N_20618,N_19949,N_19606);
nor U20619 (N_20619,N_19900,N_19747);
or U20620 (N_20620,N_19855,N_18875);
xor U20621 (N_20621,N_19709,N_19869);
nand U20622 (N_20622,N_19622,N_19887);
or U20623 (N_20623,N_18840,N_18842);
and U20624 (N_20624,N_18941,N_19147);
nor U20625 (N_20625,N_19399,N_19650);
nand U20626 (N_20626,N_19985,N_19583);
nand U20627 (N_20627,N_19065,N_19522);
nor U20628 (N_20628,N_19252,N_19398);
nor U20629 (N_20629,N_19894,N_19836);
and U20630 (N_20630,N_19645,N_19304);
and U20631 (N_20631,N_19694,N_19365);
nor U20632 (N_20632,N_18847,N_19978);
and U20633 (N_20633,N_19917,N_19315);
or U20634 (N_20634,N_19180,N_19695);
and U20635 (N_20635,N_19853,N_19585);
xnor U20636 (N_20636,N_19641,N_19467);
xnor U20637 (N_20637,N_18862,N_19133);
nor U20638 (N_20638,N_19099,N_19410);
nand U20639 (N_20639,N_18917,N_18934);
nor U20640 (N_20640,N_19436,N_18819);
and U20641 (N_20641,N_18814,N_19364);
xnor U20642 (N_20642,N_18985,N_19481);
xor U20643 (N_20643,N_18812,N_19188);
xor U20644 (N_20644,N_19880,N_18986);
or U20645 (N_20645,N_19214,N_19859);
nand U20646 (N_20646,N_19362,N_19570);
nand U20647 (N_20647,N_19959,N_19586);
nand U20648 (N_20648,N_19596,N_19034);
xnor U20649 (N_20649,N_19228,N_18940);
nand U20650 (N_20650,N_19894,N_19383);
or U20651 (N_20651,N_19206,N_19266);
and U20652 (N_20652,N_19270,N_18893);
nand U20653 (N_20653,N_19393,N_19325);
and U20654 (N_20654,N_19245,N_19125);
nand U20655 (N_20655,N_18760,N_19715);
or U20656 (N_20656,N_19394,N_18863);
xor U20657 (N_20657,N_18968,N_19755);
or U20658 (N_20658,N_19508,N_19681);
nand U20659 (N_20659,N_19159,N_19699);
or U20660 (N_20660,N_19315,N_19284);
and U20661 (N_20661,N_19674,N_19396);
and U20662 (N_20662,N_18923,N_19785);
nand U20663 (N_20663,N_18819,N_19751);
nor U20664 (N_20664,N_18889,N_19335);
and U20665 (N_20665,N_19429,N_19329);
nor U20666 (N_20666,N_19636,N_19670);
xnor U20667 (N_20667,N_19819,N_19113);
and U20668 (N_20668,N_19871,N_19437);
or U20669 (N_20669,N_18950,N_19207);
nand U20670 (N_20670,N_19466,N_19533);
nor U20671 (N_20671,N_19170,N_19149);
nand U20672 (N_20672,N_19012,N_18817);
nand U20673 (N_20673,N_19818,N_19506);
xor U20674 (N_20674,N_19784,N_19813);
xor U20675 (N_20675,N_18899,N_19615);
nor U20676 (N_20676,N_19977,N_18827);
nand U20677 (N_20677,N_19985,N_19493);
nor U20678 (N_20678,N_19377,N_19863);
or U20679 (N_20679,N_19518,N_19261);
and U20680 (N_20680,N_19353,N_19149);
nand U20681 (N_20681,N_19196,N_19837);
xor U20682 (N_20682,N_19414,N_18943);
xnor U20683 (N_20683,N_19033,N_19570);
xnor U20684 (N_20684,N_19737,N_19022);
and U20685 (N_20685,N_19072,N_19616);
and U20686 (N_20686,N_18780,N_19987);
xor U20687 (N_20687,N_19585,N_19774);
nand U20688 (N_20688,N_19675,N_19470);
or U20689 (N_20689,N_19473,N_19454);
or U20690 (N_20690,N_19535,N_19471);
and U20691 (N_20691,N_19762,N_19991);
and U20692 (N_20692,N_19956,N_19301);
or U20693 (N_20693,N_19291,N_18803);
and U20694 (N_20694,N_19745,N_19376);
nor U20695 (N_20695,N_19995,N_19979);
nand U20696 (N_20696,N_19518,N_19876);
xnor U20697 (N_20697,N_19126,N_18999);
xnor U20698 (N_20698,N_19775,N_19900);
nand U20699 (N_20699,N_18867,N_19891);
xor U20700 (N_20700,N_19099,N_19336);
xor U20701 (N_20701,N_19783,N_19084);
nand U20702 (N_20702,N_19313,N_19961);
nor U20703 (N_20703,N_19189,N_18916);
nor U20704 (N_20704,N_19043,N_18787);
xnor U20705 (N_20705,N_19329,N_19146);
or U20706 (N_20706,N_19261,N_19982);
and U20707 (N_20707,N_19460,N_19854);
xor U20708 (N_20708,N_18826,N_19392);
nor U20709 (N_20709,N_19357,N_19882);
xnor U20710 (N_20710,N_19388,N_19009);
xor U20711 (N_20711,N_19737,N_19887);
nor U20712 (N_20712,N_19459,N_18948);
xnor U20713 (N_20713,N_19311,N_19235);
nand U20714 (N_20714,N_19662,N_19490);
and U20715 (N_20715,N_19398,N_18791);
nor U20716 (N_20716,N_19374,N_18891);
or U20717 (N_20717,N_19715,N_19991);
xnor U20718 (N_20718,N_18779,N_19361);
and U20719 (N_20719,N_19426,N_19929);
nor U20720 (N_20720,N_19527,N_18768);
nor U20721 (N_20721,N_19421,N_19153);
and U20722 (N_20722,N_19732,N_18787);
nand U20723 (N_20723,N_18813,N_19007);
and U20724 (N_20724,N_19638,N_18996);
or U20725 (N_20725,N_18771,N_18860);
nor U20726 (N_20726,N_19314,N_19588);
xnor U20727 (N_20727,N_19358,N_19301);
nor U20728 (N_20728,N_18926,N_19938);
or U20729 (N_20729,N_19912,N_19387);
and U20730 (N_20730,N_18752,N_19036);
xor U20731 (N_20731,N_18847,N_19359);
nand U20732 (N_20732,N_18984,N_19722);
nor U20733 (N_20733,N_19186,N_19897);
nand U20734 (N_20734,N_19368,N_18772);
nand U20735 (N_20735,N_19353,N_19840);
xnor U20736 (N_20736,N_19581,N_19925);
nor U20737 (N_20737,N_19097,N_19384);
or U20738 (N_20738,N_19259,N_19452);
xnor U20739 (N_20739,N_19613,N_18922);
nor U20740 (N_20740,N_19757,N_19608);
and U20741 (N_20741,N_19393,N_19279);
nor U20742 (N_20742,N_19186,N_19357);
nor U20743 (N_20743,N_19956,N_19697);
or U20744 (N_20744,N_19493,N_19214);
nor U20745 (N_20745,N_19187,N_19473);
nor U20746 (N_20746,N_19089,N_19978);
and U20747 (N_20747,N_19828,N_18957);
and U20748 (N_20748,N_19445,N_19101);
and U20749 (N_20749,N_18761,N_19615);
nor U20750 (N_20750,N_19134,N_19951);
xnor U20751 (N_20751,N_19988,N_18938);
and U20752 (N_20752,N_19484,N_19268);
xnor U20753 (N_20753,N_18937,N_18877);
and U20754 (N_20754,N_19175,N_19888);
nor U20755 (N_20755,N_18920,N_19242);
and U20756 (N_20756,N_19373,N_19050);
xor U20757 (N_20757,N_19524,N_18770);
xnor U20758 (N_20758,N_19452,N_19611);
or U20759 (N_20759,N_19669,N_19921);
and U20760 (N_20760,N_19264,N_19183);
and U20761 (N_20761,N_19703,N_19632);
nand U20762 (N_20762,N_19154,N_19936);
or U20763 (N_20763,N_19432,N_19104);
nor U20764 (N_20764,N_19138,N_19986);
nand U20765 (N_20765,N_19524,N_19455);
or U20766 (N_20766,N_19984,N_19841);
xnor U20767 (N_20767,N_19678,N_19754);
xor U20768 (N_20768,N_18933,N_19424);
or U20769 (N_20769,N_19950,N_18970);
nand U20770 (N_20770,N_18765,N_19259);
nor U20771 (N_20771,N_18764,N_18871);
xor U20772 (N_20772,N_19062,N_19129);
xnor U20773 (N_20773,N_19559,N_19252);
or U20774 (N_20774,N_19081,N_19205);
or U20775 (N_20775,N_18764,N_19786);
or U20776 (N_20776,N_19519,N_19344);
nand U20777 (N_20777,N_19541,N_19010);
nor U20778 (N_20778,N_19121,N_19872);
or U20779 (N_20779,N_19547,N_19957);
nand U20780 (N_20780,N_18886,N_19560);
or U20781 (N_20781,N_18909,N_19609);
nor U20782 (N_20782,N_19216,N_19980);
nand U20783 (N_20783,N_19673,N_19388);
or U20784 (N_20784,N_19423,N_18798);
nand U20785 (N_20785,N_19070,N_18831);
nand U20786 (N_20786,N_19682,N_18973);
or U20787 (N_20787,N_19118,N_18764);
nor U20788 (N_20788,N_19154,N_19573);
and U20789 (N_20789,N_19346,N_19989);
nand U20790 (N_20790,N_19737,N_19847);
and U20791 (N_20791,N_19584,N_19231);
and U20792 (N_20792,N_19211,N_19132);
and U20793 (N_20793,N_19022,N_19952);
and U20794 (N_20794,N_18787,N_19625);
or U20795 (N_20795,N_19770,N_18839);
nand U20796 (N_20796,N_19326,N_18964);
or U20797 (N_20797,N_19828,N_19105);
xor U20798 (N_20798,N_19000,N_19771);
nor U20799 (N_20799,N_18782,N_19591);
nand U20800 (N_20800,N_19732,N_19051);
xnor U20801 (N_20801,N_19545,N_19179);
or U20802 (N_20802,N_19920,N_19831);
nand U20803 (N_20803,N_18930,N_18815);
nand U20804 (N_20804,N_19236,N_19017);
or U20805 (N_20805,N_19466,N_19985);
or U20806 (N_20806,N_19025,N_19548);
and U20807 (N_20807,N_19925,N_19617);
or U20808 (N_20808,N_19877,N_19370);
xor U20809 (N_20809,N_19559,N_19193);
nor U20810 (N_20810,N_19030,N_19078);
or U20811 (N_20811,N_18977,N_19362);
or U20812 (N_20812,N_19847,N_19219);
or U20813 (N_20813,N_18975,N_18941);
xor U20814 (N_20814,N_19128,N_19703);
nand U20815 (N_20815,N_19219,N_19263);
or U20816 (N_20816,N_18999,N_19395);
nor U20817 (N_20817,N_19085,N_19917);
xnor U20818 (N_20818,N_19419,N_19216);
xor U20819 (N_20819,N_18852,N_19976);
or U20820 (N_20820,N_19443,N_18953);
nor U20821 (N_20821,N_19178,N_19172);
xor U20822 (N_20822,N_19835,N_19280);
or U20823 (N_20823,N_19731,N_19794);
nor U20824 (N_20824,N_18868,N_19232);
nor U20825 (N_20825,N_19860,N_19066);
and U20826 (N_20826,N_19561,N_19120);
and U20827 (N_20827,N_19898,N_19092);
nand U20828 (N_20828,N_19451,N_19093);
or U20829 (N_20829,N_19779,N_19901);
nor U20830 (N_20830,N_19731,N_19802);
and U20831 (N_20831,N_19902,N_18842);
nand U20832 (N_20832,N_19965,N_19739);
nand U20833 (N_20833,N_19454,N_19267);
nor U20834 (N_20834,N_19000,N_19428);
xor U20835 (N_20835,N_18967,N_18870);
xnor U20836 (N_20836,N_19576,N_19008);
or U20837 (N_20837,N_19180,N_18779);
and U20838 (N_20838,N_19243,N_19649);
or U20839 (N_20839,N_19544,N_19976);
nor U20840 (N_20840,N_19544,N_19254);
nor U20841 (N_20841,N_19837,N_19080);
or U20842 (N_20842,N_19014,N_19247);
and U20843 (N_20843,N_18750,N_19757);
nor U20844 (N_20844,N_18764,N_19508);
xnor U20845 (N_20845,N_19059,N_19725);
nand U20846 (N_20846,N_19423,N_19802);
nand U20847 (N_20847,N_19419,N_19271);
nand U20848 (N_20848,N_19357,N_18935);
or U20849 (N_20849,N_19673,N_19423);
xnor U20850 (N_20850,N_19573,N_19982);
and U20851 (N_20851,N_19623,N_18794);
nor U20852 (N_20852,N_19067,N_19471);
and U20853 (N_20853,N_19881,N_19871);
xnor U20854 (N_20854,N_19498,N_19013);
xor U20855 (N_20855,N_19319,N_19188);
xnor U20856 (N_20856,N_18854,N_18926);
nand U20857 (N_20857,N_19530,N_19613);
or U20858 (N_20858,N_18889,N_19448);
nand U20859 (N_20859,N_19416,N_19305);
nor U20860 (N_20860,N_18993,N_19915);
nand U20861 (N_20861,N_18784,N_19712);
or U20862 (N_20862,N_19022,N_19215);
and U20863 (N_20863,N_19284,N_18947);
xnor U20864 (N_20864,N_19882,N_19602);
and U20865 (N_20865,N_19519,N_19250);
or U20866 (N_20866,N_18805,N_19808);
xnor U20867 (N_20867,N_19538,N_19957);
nand U20868 (N_20868,N_19925,N_19202);
and U20869 (N_20869,N_19075,N_19964);
nor U20870 (N_20870,N_19058,N_19203);
and U20871 (N_20871,N_19276,N_18974);
xnor U20872 (N_20872,N_19625,N_18951);
nor U20873 (N_20873,N_19869,N_19716);
nand U20874 (N_20874,N_18989,N_19047);
or U20875 (N_20875,N_19871,N_18891);
nor U20876 (N_20876,N_19040,N_19506);
or U20877 (N_20877,N_19118,N_18927);
nand U20878 (N_20878,N_19502,N_18980);
nand U20879 (N_20879,N_18794,N_19215);
nor U20880 (N_20880,N_18997,N_19005);
xnor U20881 (N_20881,N_19177,N_18864);
and U20882 (N_20882,N_18786,N_19971);
and U20883 (N_20883,N_19526,N_19655);
nor U20884 (N_20884,N_19412,N_19360);
nor U20885 (N_20885,N_18816,N_18861);
nand U20886 (N_20886,N_18894,N_19689);
nor U20887 (N_20887,N_19768,N_18760);
xor U20888 (N_20888,N_19195,N_18754);
xnor U20889 (N_20889,N_19013,N_19202);
or U20890 (N_20890,N_19951,N_19446);
and U20891 (N_20891,N_19787,N_19557);
and U20892 (N_20892,N_19209,N_18959);
and U20893 (N_20893,N_19422,N_18884);
xnor U20894 (N_20894,N_19364,N_18906);
or U20895 (N_20895,N_19573,N_19478);
or U20896 (N_20896,N_19879,N_19826);
and U20897 (N_20897,N_19029,N_19964);
nor U20898 (N_20898,N_19386,N_19557);
nor U20899 (N_20899,N_19836,N_19302);
xnor U20900 (N_20900,N_19903,N_19887);
nand U20901 (N_20901,N_19923,N_19497);
xnor U20902 (N_20902,N_19024,N_18893);
or U20903 (N_20903,N_19052,N_19100);
or U20904 (N_20904,N_18905,N_19929);
xnor U20905 (N_20905,N_19223,N_18941);
or U20906 (N_20906,N_18871,N_19365);
or U20907 (N_20907,N_19931,N_18851);
and U20908 (N_20908,N_18815,N_19034);
nand U20909 (N_20909,N_19230,N_19478);
nand U20910 (N_20910,N_18774,N_19658);
nand U20911 (N_20911,N_18998,N_19274);
or U20912 (N_20912,N_18767,N_18907);
nor U20913 (N_20913,N_19440,N_19385);
xor U20914 (N_20914,N_18986,N_19663);
xor U20915 (N_20915,N_19493,N_19684);
or U20916 (N_20916,N_19202,N_19836);
and U20917 (N_20917,N_19698,N_18963);
and U20918 (N_20918,N_18899,N_18949);
xnor U20919 (N_20919,N_18761,N_19965);
xnor U20920 (N_20920,N_19834,N_18855);
xnor U20921 (N_20921,N_19156,N_19429);
nand U20922 (N_20922,N_18962,N_19124);
xor U20923 (N_20923,N_19074,N_18986);
xor U20924 (N_20924,N_19902,N_19313);
or U20925 (N_20925,N_19089,N_19750);
xor U20926 (N_20926,N_19590,N_19917);
nor U20927 (N_20927,N_19327,N_19435);
xor U20928 (N_20928,N_19373,N_19527);
or U20929 (N_20929,N_18961,N_19241);
xor U20930 (N_20930,N_19405,N_19770);
and U20931 (N_20931,N_19189,N_18883);
nand U20932 (N_20932,N_19771,N_19361);
and U20933 (N_20933,N_19019,N_19751);
or U20934 (N_20934,N_19243,N_19434);
nor U20935 (N_20935,N_19879,N_18844);
nor U20936 (N_20936,N_19254,N_18917);
nor U20937 (N_20937,N_19408,N_19016);
nor U20938 (N_20938,N_19924,N_19180);
nand U20939 (N_20939,N_19349,N_18934);
nand U20940 (N_20940,N_19594,N_19060);
nand U20941 (N_20941,N_19423,N_19785);
nor U20942 (N_20942,N_19923,N_19025);
xor U20943 (N_20943,N_19853,N_19439);
nor U20944 (N_20944,N_18819,N_19620);
xor U20945 (N_20945,N_19270,N_18763);
and U20946 (N_20946,N_19649,N_19357);
and U20947 (N_20947,N_19329,N_19988);
nor U20948 (N_20948,N_19355,N_19740);
nand U20949 (N_20949,N_19764,N_19062);
xor U20950 (N_20950,N_19332,N_19134);
or U20951 (N_20951,N_18793,N_19912);
nand U20952 (N_20952,N_19444,N_19449);
or U20953 (N_20953,N_19206,N_18948);
and U20954 (N_20954,N_19075,N_19181);
and U20955 (N_20955,N_19077,N_19892);
nor U20956 (N_20956,N_19828,N_19091);
nor U20957 (N_20957,N_19307,N_19129);
nand U20958 (N_20958,N_19791,N_19952);
nand U20959 (N_20959,N_19783,N_19795);
nor U20960 (N_20960,N_19215,N_18819);
and U20961 (N_20961,N_19049,N_19941);
and U20962 (N_20962,N_18821,N_19557);
nor U20963 (N_20963,N_19559,N_19522);
xor U20964 (N_20964,N_19423,N_19983);
xor U20965 (N_20965,N_19799,N_19758);
or U20966 (N_20966,N_18976,N_19872);
nor U20967 (N_20967,N_19049,N_19786);
or U20968 (N_20968,N_19297,N_19366);
xor U20969 (N_20969,N_18773,N_19456);
nor U20970 (N_20970,N_18837,N_19650);
or U20971 (N_20971,N_19554,N_19203);
nand U20972 (N_20972,N_18842,N_18791);
and U20973 (N_20973,N_19079,N_19754);
or U20974 (N_20974,N_18858,N_19734);
or U20975 (N_20975,N_19752,N_19154);
and U20976 (N_20976,N_19662,N_19624);
or U20977 (N_20977,N_19067,N_19975);
xor U20978 (N_20978,N_18929,N_19920);
xor U20979 (N_20979,N_19447,N_19550);
xor U20980 (N_20980,N_19107,N_19626);
nor U20981 (N_20981,N_18801,N_19129);
or U20982 (N_20982,N_19352,N_19816);
xnor U20983 (N_20983,N_19846,N_19198);
nor U20984 (N_20984,N_19338,N_19190);
or U20985 (N_20985,N_19530,N_19685);
or U20986 (N_20986,N_19054,N_19886);
nand U20987 (N_20987,N_19523,N_19747);
and U20988 (N_20988,N_19083,N_18802);
xnor U20989 (N_20989,N_18867,N_19117);
xor U20990 (N_20990,N_19701,N_19760);
xnor U20991 (N_20991,N_19152,N_18902);
or U20992 (N_20992,N_18914,N_19277);
xnor U20993 (N_20993,N_19354,N_19981);
xor U20994 (N_20994,N_19874,N_19657);
or U20995 (N_20995,N_19319,N_19779);
xnor U20996 (N_20996,N_18810,N_18907);
nand U20997 (N_20997,N_19392,N_19144);
and U20998 (N_20998,N_19000,N_19466);
xnor U20999 (N_20999,N_18781,N_19663);
or U21000 (N_21000,N_19686,N_19321);
nand U21001 (N_21001,N_19436,N_19716);
or U21002 (N_21002,N_19213,N_19323);
and U21003 (N_21003,N_19103,N_18882);
nand U21004 (N_21004,N_19648,N_19995);
nand U21005 (N_21005,N_19446,N_19230);
nand U21006 (N_21006,N_19748,N_19737);
nor U21007 (N_21007,N_19115,N_19180);
and U21008 (N_21008,N_19709,N_19363);
or U21009 (N_21009,N_19610,N_19519);
nor U21010 (N_21010,N_19536,N_18861);
nand U21011 (N_21011,N_19852,N_19440);
xnor U21012 (N_21012,N_19039,N_19653);
nor U21013 (N_21013,N_19839,N_19532);
xnor U21014 (N_21014,N_19805,N_18884);
or U21015 (N_21015,N_19786,N_19841);
xor U21016 (N_21016,N_18898,N_18824);
and U21017 (N_21017,N_19638,N_19907);
xnor U21018 (N_21018,N_19702,N_18853);
nand U21019 (N_21019,N_19653,N_19778);
nand U21020 (N_21020,N_19997,N_18886);
xor U21021 (N_21021,N_19486,N_19470);
xnor U21022 (N_21022,N_19583,N_18996);
and U21023 (N_21023,N_19634,N_19244);
and U21024 (N_21024,N_19911,N_18773);
or U21025 (N_21025,N_19865,N_18992);
or U21026 (N_21026,N_19531,N_19189);
nand U21027 (N_21027,N_19102,N_19920);
or U21028 (N_21028,N_18829,N_19215);
or U21029 (N_21029,N_19029,N_19513);
or U21030 (N_21030,N_18848,N_19991);
nor U21031 (N_21031,N_19460,N_19640);
nand U21032 (N_21032,N_18921,N_18981);
xnor U21033 (N_21033,N_19171,N_19319);
xor U21034 (N_21034,N_18942,N_18831);
nand U21035 (N_21035,N_19150,N_19135);
nor U21036 (N_21036,N_19138,N_19429);
or U21037 (N_21037,N_18832,N_19186);
xnor U21038 (N_21038,N_19704,N_18795);
xnor U21039 (N_21039,N_19959,N_18945);
nor U21040 (N_21040,N_18781,N_19476);
nand U21041 (N_21041,N_19924,N_19696);
xnor U21042 (N_21042,N_19364,N_19356);
and U21043 (N_21043,N_19846,N_19809);
or U21044 (N_21044,N_19492,N_18992);
nor U21045 (N_21045,N_19326,N_19487);
or U21046 (N_21046,N_19901,N_19591);
nand U21047 (N_21047,N_19423,N_19194);
nor U21048 (N_21048,N_19446,N_18914);
nand U21049 (N_21049,N_19110,N_19808);
nand U21050 (N_21050,N_19281,N_19422);
and U21051 (N_21051,N_19281,N_19315);
or U21052 (N_21052,N_19370,N_19849);
xor U21053 (N_21053,N_18973,N_19050);
and U21054 (N_21054,N_18938,N_19155);
nor U21055 (N_21055,N_19346,N_18945);
or U21056 (N_21056,N_19401,N_18980);
nand U21057 (N_21057,N_19905,N_19077);
and U21058 (N_21058,N_18907,N_19529);
and U21059 (N_21059,N_19130,N_19800);
and U21060 (N_21060,N_19545,N_18997);
xor U21061 (N_21061,N_19748,N_19943);
nor U21062 (N_21062,N_19974,N_19832);
and U21063 (N_21063,N_19239,N_19788);
and U21064 (N_21064,N_19850,N_19816);
or U21065 (N_21065,N_19630,N_19138);
and U21066 (N_21066,N_18945,N_19518);
and U21067 (N_21067,N_19988,N_18928);
nor U21068 (N_21068,N_19430,N_19606);
xnor U21069 (N_21069,N_19039,N_19108);
and U21070 (N_21070,N_18815,N_19852);
nand U21071 (N_21071,N_18786,N_18976);
nor U21072 (N_21072,N_19992,N_19002);
xor U21073 (N_21073,N_19555,N_19588);
xor U21074 (N_21074,N_18812,N_19354);
or U21075 (N_21075,N_19238,N_19913);
nand U21076 (N_21076,N_19426,N_19977);
or U21077 (N_21077,N_19135,N_19967);
nor U21078 (N_21078,N_19675,N_18930);
nand U21079 (N_21079,N_19960,N_19044);
xor U21080 (N_21080,N_19065,N_19717);
and U21081 (N_21081,N_19726,N_19607);
nor U21082 (N_21082,N_19035,N_19284);
nor U21083 (N_21083,N_19181,N_19369);
xnor U21084 (N_21084,N_19588,N_19462);
and U21085 (N_21085,N_18795,N_19145);
or U21086 (N_21086,N_19338,N_18817);
nand U21087 (N_21087,N_19130,N_19633);
and U21088 (N_21088,N_19828,N_19585);
or U21089 (N_21089,N_19988,N_19916);
nand U21090 (N_21090,N_19049,N_19587);
nand U21091 (N_21091,N_19314,N_19897);
and U21092 (N_21092,N_19883,N_19202);
and U21093 (N_21093,N_18966,N_19283);
nor U21094 (N_21094,N_19089,N_19925);
and U21095 (N_21095,N_19575,N_19814);
nor U21096 (N_21096,N_19249,N_19655);
nand U21097 (N_21097,N_19747,N_19067);
and U21098 (N_21098,N_19616,N_19872);
nor U21099 (N_21099,N_19475,N_18896);
nand U21100 (N_21100,N_19708,N_19869);
xnor U21101 (N_21101,N_19691,N_19281);
and U21102 (N_21102,N_18980,N_19144);
and U21103 (N_21103,N_18855,N_19652);
nor U21104 (N_21104,N_19150,N_19848);
xnor U21105 (N_21105,N_19909,N_19031);
or U21106 (N_21106,N_19024,N_19817);
nand U21107 (N_21107,N_19481,N_18867);
xor U21108 (N_21108,N_19554,N_19223);
and U21109 (N_21109,N_19659,N_18760);
and U21110 (N_21110,N_19330,N_18763);
nor U21111 (N_21111,N_19261,N_18788);
and U21112 (N_21112,N_19883,N_19463);
nand U21113 (N_21113,N_19196,N_19637);
xor U21114 (N_21114,N_18998,N_19312);
or U21115 (N_21115,N_18813,N_19860);
or U21116 (N_21116,N_18882,N_19559);
nand U21117 (N_21117,N_19364,N_19292);
nand U21118 (N_21118,N_19790,N_18977);
nand U21119 (N_21119,N_19024,N_18838);
nor U21120 (N_21120,N_19685,N_19042);
or U21121 (N_21121,N_18977,N_19927);
nand U21122 (N_21122,N_19012,N_19308);
nand U21123 (N_21123,N_19222,N_19611);
xnor U21124 (N_21124,N_19700,N_19204);
xor U21125 (N_21125,N_19508,N_18939);
nand U21126 (N_21126,N_19943,N_19595);
or U21127 (N_21127,N_19504,N_19419);
nor U21128 (N_21128,N_19424,N_18801);
or U21129 (N_21129,N_19527,N_19844);
nor U21130 (N_21130,N_19726,N_19107);
nor U21131 (N_21131,N_19231,N_19398);
or U21132 (N_21132,N_19792,N_18890);
or U21133 (N_21133,N_18842,N_19609);
nor U21134 (N_21134,N_19374,N_19712);
nor U21135 (N_21135,N_19559,N_18811);
nand U21136 (N_21136,N_19129,N_19768);
xor U21137 (N_21137,N_19363,N_19547);
nand U21138 (N_21138,N_19907,N_19708);
or U21139 (N_21139,N_18791,N_19441);
or U21140 (N_21140,N_18780,N_19319);
nand U21141 (N_21141,N_19193,N_19733);
xnor U21142 (N_21142,N_19371,N_19501);
nor U21143 (N_21143,N_19925,N_19454);
or U21144 (N_21144,N_19238,N_18754);
xor U21145 (N_21145,N_18888,N_19248);
nor U21146 (N_21146,N_19466,N_19875);
nor U21147 (N_21147,N_19645,N_19852);
nor U21148 (N_21148,N_19504,N_19083);
nor U21149 (N_21149,N_18892,N_19715);
xnor U21150 (N_21150,N_18863,N_19488);
and U21151 (N_21151,N_18996,N_19260);
or U21152 (N_21152,N_18973,N_19201);
and U21153 (N_21153,N_18949,N_18800);
xor U21154 (N_21154,N_19963,N_19044);
nand U21155 (N_21155,N_19859,N_19375);
or U21156 (N_21156,N_19562,N_19412);
xor U21157 (N_21157,N_18901,N_19638);
nor U21158 (N_21158,N_19110,N_19009);
xnor U21159 (N_21159,N_19938,N_19364);
nand U21160 (N_21160,N_19459,N_19641);
xnor U21161 (N_21161,N_19854,N_19414);
and U21162 (N_21162,N_19980,N_19153);
and U21163 (N_21163,N_19698,N_19034);
xor U21164 (N_21164,N_19442,N_19294);
and U21165 (N_21165,N_19579,N_19087);
or U21166 (N_21166,N_19894,N_18955);
and U21167 (N_21167,N_19622,N_19618);
nor U21168 (N_21168,N_19189,N_19676);
and U21169 (N_21169,N_18784,N_19329);
and U21170 (N_21170,N_18896,N_18888);
xnor U21171 (N_21171,N_19935,N_18781);
or U21172 (N_21172,N_19431,N_18896);
xnor U21173 (N_21173,N_19588,N_18970);
nor U21174 (N_21174,N_19231,N_19498);
xor U21175 (N_21175,N_19623,N_18776);
nor U21176 (N_21176,N_19852,N_19746);
nand U21177 (N_21177,N_18801,N_19363);
xor U21178 (N_21178,N_19988,N_19560);
and U21179 (N_21179,N_19904,N_19358);
nand U21180 (N_21180,N_19178,N_19840);
or U21181 (N_21181,N_18940,N_19508);
or U21182 (N_21182,N_19700,N_19865);
xnor U21183 (N_21183,N_19023,N_19762);
xnor U21184 (N_21184,N_19686,N_19491);
or U21185 (N_21185,N_19739,N_19800);
or U21186 (N_21186,N_19629,N_19531);
xnor U21187 (N_21187,N_19118,N_19476);
nand U21188 (N_21188,N_18980,N_18986);
and U21189 (N_21189,N_19110,N_19572);
nand U21190 (N_21190,N_19952,N_19465);
xnor U21191 (N_21191,N_19353,N_19718);
nor U21192 (N_21192,N_19382,N_18894);
or U21193 (N_21193,N_19722,N_18850);
xnor U21194 (N_21194,N_19118,N_19904);
and U21195 (N_21195,N_18900,N_19171);
nor U21196 (N_21196,N_19752,N_18991);
and U21197 (N_21197,N_19438,N_19169);
nor U21198 (N_21198,N_19528,N_19268);
nand U21199 (N_21199,N_19943,N_19768);
nand U21200 (N_21200,N_18940,N_19539);
and U21201 (N_21201,N_19053,N_19792);
or U21202 (N_21202,N_19609,N_18901);
and U21203 (N_21203,N_19414,N_19346);
xor U21204 (N_21204,N_19517,N_19987);
nand U21205 (N_21205,N_19873,N_19635);
xor U21206 (N_21206,N_18998,N_19977);
or U21207 (N_21207,N_19780,N_19999);
and U21208 (N_21208,N_18760,N_19458);
nor U21209 (N_21209,N_19409,N_19368);
nor U21210 (N_21210,N_19123,N_19615);
xor U21211 (N_21211,N_19651,N_18778);
nor U21212 (N_21212,N_19200,N_19844);
nand U21213 (N_21213,N_19784,N_18782);
nand U21214 (N_21214,N_18791,N_19971);
or U21215 (N_21215,N_19070,N_19652);
nor U21216 (N_21216,N_18888,N_19141);
or U21217 (N_21217,N_19624,N_19387);
nand U21218 (N_21218,N_19975,N_19575);
and U21219 (N_21219,N_19752,N_19601);
xnor U21220 (N_21220,N_19455,N_19825);
nand U21221 (N_21221,N_19839,N_19952);
nand U21222 (N_21222,N_19968,N_19993);
nor U21223 (N_21223,N_19056,N_19048);
nor U21224 (N_21224,N_19439,N_19755);
and U21225 (N_21225,N_19322,N_18757);
or U21226 (N_21226,N_19889,N_19677);
nor U21227 (N_21227,N_19716,N_19010);
nand U21228 (N_21228,N_18866,N_19516);
or U21229 (N_21229,N_19816,N_18910);
nor U21230 (N_21230,N_18994,N_18972);
nand U21231 (N_21231,N_18945,N_19573);
or U21232 (N_21232,N_18822,N_19008);
and U21233 (N_21233,N_19379,N_19691);
nand U21234 (N_21234,N_19691,N_19117);
or U21235 (N_21235,N_19760,N_19705);
and U21236 (N_21236,N_19211,N_19732);
or U21237 (N_21237,N_19083,N_19721);
and U21238 (N_21238,N_19639,N_18933);
nand U21239 (N_21239,N_19524,N_18760);
nand U21240 (N_21240,N_19987,N_18868);
nand U21241 (N_21241,N_19760,N_18754);
xnor U21242 (N_21242,N_19893,N_19544);
nand U21243 (N_21243,N_18809,N_19783);
or U21244 (N_21244,N_19347,N_19393);
and U21245 (N_21245,N_19344,N_19947);
xor U21246 (N_21246,N_19041,N_19460);
xnor U21247 (N_21247,N_19229,N_19880);
xnor U21248 (N_21248,N_18918,N_18932);
nand U21249 (N_21249,N_19762,N_19659);
nand U21250 (N_21250,N_21164,N_20863);
or U21251 (N_21251,N_20247,N_20624);
and U21252 (N_21252,N_21145,N_20742);
xnor U21253 (N_21253,N_20349,N_21073);
xnor U21254 (N_21254,N_20836,N_20396);
or U21255 (N_21255,N_20948,N_20980);
and U21256 (N_21256,N_20075,N_20004);
nand U21257 (N_21257,N_21028,N_20890);
nand U21258 (N_21258,N_20780,N_20194);
xor U21259 (N_21259,N_20280,N_20486);
or U21260 (N_21260,N_20515,N_20435);
xor U21261 (N_21261,N_20124,N_20957);
nand U21262 (N_21262,N_20110,N_20489);
xnor U21263 (N_21263,N_20611,N_20900);
or U21264 (N_21264,N_20111,N_20255);
nand U21265 (N_21265,N_20456,N_20764);
nand U21266 (N_21266,N_21107,N_20552);
xnor U21267 (N_21267,N_20123,N_21103);
or U21268 (N_21268,N_20202,N_20471);
xnor U21269 (N_21269,N_21142,N_20267);
nand U21270 (N_21270,N_21171,N_20620);
and U21271 (N_21271,N_20967,N_21088);
xnor U21272 (N_21272,N_21032,N_20031);
xnor U21273 (N_21273,N_20180,N_20477);
or U21274 (N_21274,N_20057,N_21169);
xor U21275 (N_21275,N_21187,N_20120);
nand U21276 (N_21276,N_20532,N_20335);
and U21277 (N_21277,N_21000,N_20952);
nand U21278 (N_21278,N_20705,N_20023);
and U21279 (N_21279,N_20970,N_21012);
nand U21280 (N_21280,N_20511,N_20706);
nor U21281 (N_21281,N_20412,N_20974);
or U21282 (N_21282,N_20938,N_21120);
nand U21283 (N_21283,N_20039,N_21234);
and U21284 (N_21284,N_20136,N_20521);
and U21285 (N_21285,N_20723,N_20361);
and U21286 (N_21286,N_20106,N_20466);
and U21287 (N_21287,N_20577,N_20140);
xor U21288 (N_21288,N_20181,N_20072);
nand U21289 (N_21289,N_20698,N_20083);
or U21290 (N_21290,N_20289,N_21183);
nor U21291 (N_21291,N_20287,N_20442);
or U21292 (N_21292,N_20513,N_20953);
or U21293 (N_21293,N_20818,N_20768);
nand U21294 (N_21294,N_20531,N_21218);
nor U21295 (N_21295,N_20784,N_20528);
nand U21296 (N_21296,N_20363,N_20209);
nor U21297 (N_21297,N_20210,N_20258);
xnor U21298 (N_21298,N_20915,N_20218);
and U21299 (N_21299,N_20104,N_21002);
nor U21300 (N_21300,N_21152,N_20036);
nor U21301 (N_21301,N_20771,N_20386);
and U21302 (N_21302,N_20137,N_20714);
nor U21303 (N_21303,N_20642,N_20332);
and U21304 (N_21304,N_20944,N_20141);
or U21305 (N_21305,N_21087,N_20109);
nand U21306 (N_21306,N_20983,N_20382);
or U21307 (N_21307,N_20849,N_20082);
nor U21308 (N_21308,N_20084,N_20126);
xnor U21309 (N_21309,N_21024,N_20352);
xnor U21310 (N_21310,N_21137,N_21228);
or U21311 (N_21311,N_20519,N_20167);
or U21312 (N_21312,N_20282,N_21094);
nand U21313 (N_21313,N_20174,N_20512);
or U21314 (N_21314,N_20424,N_20516);
or U21315 (N_21315,N_20445,N_21082);
and U21316 (N_21316,N_20748,N_20778);
nor U21317 (N_21317,N_20872,N_20256);
nor U21318 (N_21318,N_21102,N_20024);
or U21319 (N_21319,N_21134,N_20753);
nor U21320 (N_21320,N_20372,N_20875);
and U21321 (N_21321,N_20285,N_21014);
nor U21322 (N_21322,N_20648,N_20862);
xnor U21323 (N_21323,N_20783,N_20584);
or U21324 (N_21324,N_20767,N_20251);
nand U21325 (N_21325,N_21104,N_20250);
xnor U21326 (N_21326,N_21056,N_20319);
or U21327 (N_21327,N_20030,N_20945);
and U21328 (N_21328,N_20409,N_20188);
xnor U21329 (N_21329,N_20143,N_20708);
xor U21330 (N_21330,N_21116,N_20990);
and U21331 (N_21331,N_21242,N_20431);
and U21332 (N_21332,N_20831,N_20520);
and U21333 (N_21333,N_20840,N_20861);
or U21334 (N_21334,N_20786,N_21226);
xnor U21335 (N_21335,N_20704,N_21208);
nor U21336 (N_21336,N_20594,N_21215);
and U21337 (N_21337,N_20310,N_20096);
xor U21338 (N_21338,N_20189,N_21007);
nand U21339 (N_21339,N_20581,N_21176);
nand U21340 (N_21340,N_20149,N_20749);
or U21341 (N_21341,N_20173,N_21243);
and U21342 (N_21342,N_20437,N_20331);
xor U21343 (N_21343,N_20606,N_20851);
xnor U21344 (N_21344,N_20514,N_20438);
xor U21345 (N_21345,N_21105,N_21182);
nor U21346 (N_21346,N_20654,N_20949);
nand U21347 (N_21347,N_21217,N_20660);
nand U21348 (N_21348,N_20160,N_20558);
and U21349 (N_21349,N_20345,N_20542);
nor U21350 (N_21350,N_20619,N_21184);
xnor U21351 (N_21351,N_20774,N_20572);
xnor U21352 (N_21352,N_20905,N_20709);
nor U21353 (N_21353,N_20668,N_21197);
nor U21354 (N_21354,N_20187,N_21106);
and U21355 (N_21355,N_20797,N_20587);
nand U21356 (N_21356,N_20919,N_20899);
xor U21357 (N_21357,N_20557,N_20377);
xor U21358 (N_21358,N_21231,N_21232);
xnor U21359 (N_21359,N_20071,N_20399);
and U21360 (N_21360,N_21009,N_20673);
nand U21361 (N_21361,N_20266,N_20378);
or U21362 (N_21362,N_20205,N_20088);
xor U21363 (N_21363,N_20789,N_20802);
nor U21364 (N_21364,N_20406,N_21011);
xnor U21365 (N_21365,N_21119,N_20598);
or U21366 (N_21366,N_20394,N_20597);
or U21367 (N_21367,N_20035,N_20834);
or U21368 (N_21368,N_20718,N_20400);
xnor U21369 (N_21369,N_20657,N_21241);
or U21370 (N_21370,N_20274,N_20573);
or U21371 (N_21371,N_20571,N_20485);
nand U21372 (N_21372,N_21008,N_21213);
nor U21373 (N_21373,N_20259,N_21147);
xnor U21374 (N_21374,N_20252,N_20719);
or U21375 (N_21375,N_20279,N_20956);
nor U21376 (N_21376,N_20042,N_21224);
xnor U21377 (N_21377,N_20468,N_20765);
nor U21378 (N_21378,N_20344,N_20968);
nand U21379 (N_21379,N_20248,N_20398);
or U21380 (N_21380,N_20551,N_20601);
nor U21381 (N_21381,N_20225,N_20314);
nand U21382 (N_21382,N_21239,N_20483);
nand U21383 (N_21383,N_20070,N_20965);
xnor U21384 (N_21384,N_21118,N_20014);
nor U21385 (N_21385,N_20249,N_20046);
nand U21386 (N_21386,N_21076,N_20716);
nand U21387 (N_21387,N_20121,N_21079);
and U21388 (N_21388,N_20053,N_20838);
xnor U21389 (N_21389,N_20565,N_21085);
nand U21390 (N_21390,N_20067,N_20493);
nand U21391 (N_21391,N_20393,N_20627);
or U21392 (N_21392,N_20777,N_20074);
or U21393 (N_21393,N_20504,N_20475);
xor U21394 (N_21394,N_20800,N_21175);
nor U21395 (N_21395,N_20446,N_21053);
nand U21396 (N_21396,N_20045,N_20626);
nand U21397 (N_21397,N_20755,N_21138);
xnor U21398 (N_21398,N_20901,N_20044);
nor U21399 (N_21399,N_20479,N_21036);
and U21400 (N_21400,N_20145,N_20237);
and U21401 (N_21401,N_20118,N_20293);
xor U21402 (N_21402,N_21127,N_20553);
nor U21403 (N_21403,N_21043,N_20159);
xor U21404 (N_21404,N_20478,N_20745);
or U21405 (N_21405,N_20644,N_21146);
nor U21406 (N_21406,N_20871,N_20633);
nand U21407 (N_21407,N_20991,N_20824);
xnor U21408 (N_21408,N_21030,N_20081);
nand U21409 (N_21409,N_20147,N_20452);
nand U21410 (N_21410,N_20895,N_20199);
or U21411 (N_21411,N_20533,N_20954);
nand U21412 (N_21412,N_20404,N_20391);
or U21413 (N_21413,N_20904,N_20823);
nor U21414 (N_21414,N_20505,N_20848);
or U21415 (N_21415,N_21021,N_20085);
or U21416 (N_21416,N_20821,N_20175);
xnor U21417 (N_21417,N_21029,N_21225);
nor U21418 (N_21418,N_21206,N_21204);
and U21419 (N_21419,N_21126,N_21202);
or U21420 (N_21420,N_21001,N_20882);
or U21421 (N_21421,N_20675,N_20560);
nor U21422 (N_21422,N_20865,N_20960);
and U21423 (N_21423,N_20304,N_20729);
xor U21424 (N_21424,N_21189,N_20739);
xor U21425 (N_21425,N_21086,N_20273);
nand U21426 (N_21426,N_20315,N_21018);
and U21427 (N_21427,N_20924,N_20766);
or U21428 (N_21428,N_21039,N_20530);
nor U21429 (N_21429,N_20506,N_20001);
and U21430 (N_21430,N_20610,N_20793);
and U21431 (N_21431,N_20829,N_20317);
nor U21432 (N_21432,N_20822,N_20782);
or U21433 (N_21433,N_20077,N_20029);
or U21434 (N_21434,N_20451,N_20996);
and U21435 (N_21435,N_21070,N_21060);
or U21436 (N_21436,N_20561,N_20734);
nor U21437 (N_21437,N_20699,N_21219);
or U21438 (N_21438,N_20725,N_20984);
nand U21439 (N_21439,N_20667,N_20387);
nand U21440 (N_21440,N_20320,N_20231);
nor U21441 (N_21441,N_20679,N_20607);
xor U21442 (N_21442,N_20423,N_20683);
xnor U21443 (N_21443,N_21214,N_20918);
nand U21444 (N_21444,N_20791,N_20737);
xnor U21445 (N_21445,N_20876,N_20336);
and U21446 (N_21446,N_20065,N_21095);
xnor U21447 (N_21447,N_21003,N_21025);
and U21448 (N_21448,N_20550,N_20888);
and U21449 (N_21449,N_20941,N_20186);
or U21450 (N_21450,N_20695,N_20977);
or U21451 (N_21451,N_21249,N_20214);
xnor U21452 (N_21452,N_20384,N_20041);
or U21453 (N_21453,N_20226,N_20321);
or U21454 (N_21454,N_21222,N_20054);
nor U21455 (N_21455,N_20963,N_20129);
nand U21456 (N_21456,N_21123,N_20694);
or U21457 (N_21457,N_20715,N_20578);
and U21458 (N_21458,N_20864,N_20211);
nand U21459 (N_21459,N_20652,N_20373);
nor U21460 (N_21460,N_20987,N_20613);
and U21461 (N_21461,N_20710,N_20858);
or U21462 (N_21462,N_21181,N_20116);
or U21463 (N_21463,N_20690,N_20665);
nor U21464 (N_21464,N_20548,N_20870);
or U21465 (N_21465,N_20212,N_20672);
and U21466 (N_21466,N_20405,N_20856);
and U21467 (N_21467,N_20702,N_21108);
and U21468 (N_21468,N_20019,N_20027);
xnor U21469 (N_21469,N_20228,N_20150);
and U21470 (N_21470,N_20501,N_20855);
or U21471 (N_21471,N_20312,N_21015);
nor U21472 (N_21472,N_20877,N_21122);
and U21473 (N_21473,N_20306,N_20687);
nor U21474 (N_21474,N_20241,N_20380);
or U21475 (N_21475,N_20508,N_20554);
xor U21476 (N_21476,N_20507,N_20425);
and U21477 (N_21477,N_20158,N_20916);
nand U21478 (N_21478,N_20402,N_20224);
nor U21479 (N_21479,N_21034,N_20495);
nor U21480 (N_21480,N_20682,N_20239);
or U21481 (N_21481,N_20850,N_21203);
nor U21482 (N_21482,N_21031,N_20462);
and U21483 (N_21483,N_21240,N_21020);
and U21484 (N_21484,N_21046,N_21083);
nand U21485 (N_21485,N_20102,N_20685);
and U21486 (N_21486,N_20887,N_20852);
nor U21487 (N_21487,N_20902,N_20647);
or U21488 (N_21488,N_21044,N_20847);
nand U21489 (N_21489,N_20482,N_21019);
nand U21490 (N_21490,N_20388,N_20222);
nand U21491 (N_21491,N_20217,N_20351);
or U21492 (N_21492,N_21063,N_20414);
and U21493 (N_21493,N_21190,N_20892);
xor U21494 (N_21494,N_21037,N_21067);
xor U21495 (N_21495,N_20153,N_20885);
and U21496 (N_21496,N_20333,N_20236);
xnor U21497 (N_21497,N_20411,N_20474);
nand U21498 (N_21498,N_20490,N_20113);
and U21499 (N_21499,N_21097,N_20208);
and U21500 (N_21500,N_20305,N_20366);
xnor U21501 (N_21501,N_21174,N_20549);
and U21502 (N_21502,N_20441,N_20804);
xor U21503 (N_21503,N_20176,N_20012);
xnor U21504 (N_21504,N_20357,N_20052);
and U21505 (N_21505,N_21080,N_20947);
or U21506 (N_21506,N_20229,N_20839);
nand U21507 (N_21507,N_20827,N_20166);
nand U21508 (N_21508,N_20711,N_20599);
or U21509 (N_21509,N_20061,N_20139);
or U21510 (N_21510,N_21022,N_20098);
xnor U21511 (N_21511,N_20650,N_20720);
and U21512 (N_21512,N_20105,N_20903);
nor U21513 (N_21513,N_20461,N_20368);
or U21514 (N_21514,N_21244,N_20112);
and U21515 (N_21515,N_21178,N_21074);
or U21516 (N_21516,N_20353,N_20346);
and U21517 (N_21517,N_20868,N_21235);
nand U21518 (N_21518,N_20591,N_20283);
nand U21519 (N_21519,N_20743,N_21196);
xnor U21520 (N_21520,N_20093,N_20763);
or U21521 (N_21521,N_20942,N_20590);
or U21522 (N_21522,N_20585,N_20544);
and U21523 (N_21523,N_20064,N_20617);
xor U21524 (N_21524,N_20204,N_21210);
and U21525 (N_21525,N_20732,N_20303);
and U21526 (N_21526,N_20575,N_20994);
and U21527 (N_21527,N_20663,N_20546);
and U21528 (N_21528,N_20661,N_20750);
or U21529 (N_21529,N_20263,N_20108);
or U21530 (N_21530,N_20889,N_21061);
nand U21531 (N_21531,N_20896,N_20701);
nand U21532 (N_21532,N_20801,N_20670);
and U21533 (N_21533,N_21033,N_20148);
or U21534 (N_21534,N_20284,N_20286);
nand U21535 (N_21535,N_21006,N_21200);
or U21536 (N_21536,N_20040,N_20612);
xnor U21537 (N_21537,N_20161,N_20527);
or U21538 (N_21538,N_20609,N_20751);
and U21539 (N_21539,N_20447,N_20658);
or U21540 (N_21540,N_21163,N_20815);
and U21541 (N_21541,N_20066,N_21059);
xnor U21542 (N_21542,N_20413,N_21177);
or U21543 (N_21543,N_20350,N_21193);
or U21544 (N_21544,N_20966,N_20635);
nand U21545 (N_21545,N_20260,N_20500);
nor U21546 (N_21546,N_20419,N_20828);
xnor U21547 (N_21547,N_20367,N_20130);
and U21548 (N_21548,N_20969,N_21151);
nor U21549 (N_21549,N_20195,N_20343);
and U21550 (N_21550,N_20232,N_20458);
nor U21551 (N_21551,N_20999,N_20676);
nand U21552 (N_21552,N_20817,N_20625);
nor U21553 (N_21553,N_20634,N_20922);
nor U21554 (N_21554,N_21180,N_21161);
and U21555 (N_21555,N_20997,N_20271);
nor U21556 (N_21556,N_20292,N_20989);
xor U21557 (N_21557,N_20788,N_20152);
nand U21558 (N_21558,N_20201,N_20296);
or U21559 (N_21559,N_20596,N_21040);
and U21560 (N_21560,N_20569,N_20993);
xor U21561 (N_21561,N_20666,N_21112);
and U21562 (N_21562,N_20092,N_20976);
and U21563 (N_21563,N_20826,N_20459);
or U21564 (N_21564,N_20308,N_20220);
nand U21565 (N_21565,N_20940,N_20009);
or U21566 (N_21566,N_20497,N_21153);
and U21567 (N_21567,N_20299,N_21064);
and U21568 (N_21568,N_20480,N_21078);
and U21569 (N_21569,N_20154,N_20428);
nor U21570 (N_21570,N_20741,N_20354);
and U21571 (N_21571,N_21004,N_20342);
xor U21572 (N_21572,N_20931,N_20509);
xor U21573 (N_21573,N_20262,N_20177);
or U21574 (N_21574,N_20873,N_20168);
and U21575 (N_21575,N_20146,N_20684);
nor U21576 (N_21576,N_20358,N_20586);
and U21577 (N_21577,N_20323,N_20355);
and U21578 (N_21578,N_20874,N_21090);
and U21579 (N_21579,N_20646,N_20752);
or U21580 (N_21580,N_20614,N_21160);
xor U21581 (N_21581,N_20713,N_20089);
or U21582 (N_21582,N_20866,N_20196);
xor U21583 (N_21583,N_20920,N_21065);
nor U21584 (N_21584,N_21212,N_20117);
or U21585 (N_21585,N_20328,N_20122);
or U21586 (N_21586,N_20978,N_20526);
and U21587 (N_21587,N_21130,N_20604);
nor U21588 (N_21588,N_20006,N_20488);
or U21589 (N_21589,N_21050,N_21049);
and U21590 (N_21590,N_21198,N_21055);
xor U21591 (N_21591,N_20772,N_20568);
or U21592 (N_21592,N_20639,N_20812);
nor U21593 (N_21593,N_20681,N_20392);
nor U21594 (N_21594,N_20295,N_20770);
or U21595 (N_21595,N_20570,N_20397);
nor U21596 (N_21596,N_20884,N_21109);
nor U21597 (N_21597,N_20165,N_20806);
nor U21598 (N_21598,N_20216,N_20517);
and U21599 (N_21599,N_20691,N_20653);
or U21600 (N_21600,N_21185,N_20465);
nor U21601 (N_21601,N_20207,N_21081);
nor U21602 (N_21602,N_20334,N_20934);
xnor U21603 (N_21603,N_20003,N_21236);
nand U21604 (N_21604,N_20359,N_20325);
nand U21605 (N_21605,N_20007,N_20757);
nor U21606 (N_21606,N_20680,N_20717);
and U21607 (N_21607,N_20339,N_20433);
nor U21608 (N_21608,N_21139,N_20923);
or U21609 (N_21609,N_20401,N_20936);
xnor U21610 (N_21610,N_20503,N_20499);
or U21611 (N_21611,N_20453,N_20986);
nor U21612 (N_21612,N_21237,N_21027);
xnor U21613 (N_21613,N_21069,N_20629);
or U21614 (N_21614,N_20525,N_21023);
and U21615 (N_21615,N_20820,N_20157);
and U21616 (N_21616,N_20979,N_20932);
xor U21617 (N_21617,N_20638,N_20700);
and U21618 (N_21618,N_20807,N_20277);
xnor U21619 (N_21619,N_21209,N_20728);
nor U21620 (N_21620,N_20671,N_21159);
or U21621 (N_21621,N_20559,N_20127);
nor U21622 (N_21622,N_20379,N_20927);
xnor U21623 (N_21623,N_20107,N_20811);
nand U21624 (N_21624,N_20078,N_20630);
nor U21625 (N_21625,N_21092,N_20011);
xor U21626 (N_21626,N_20600,N_20434);
nor U21627 (N_21627,N_20860,N_21052);
xnor U21628 (N_21628,N_20794,N_20950);
nor U21629 (N_21629,N_20664,N_20484);
or U21630 (N_21630,N_20450,N_20535);
nor U21631 (N_21631,N_20841,N_20191);
and U21632 (N_21632,N_20926,N_20050);
or U21633 (N_21633,N_20929,N_20537);
and U21634 (N_21634,N_21101,N_20254);
and U21635 (N_21635,N_20426,N_20440);
or U21636 (N_21636,N_20883,N_21140);
nor U21637 (N_21637,N_20301,N_20238);
nand U21638 (N_21638,N_20193,N_20076);
nor U21639 (N_21639,N_21038,N_21246);
nand U21640 (N_21640,N_20015,N_21093);
nand U21641 (N_21641,N_20534,N_20094);
or U21642 (N_21642,N_20416,N_20637);
xor U21643 (N_21643,N_20138,N_20142);
nor U21644 (N_21644,N_20917,N_20491);
and U21645 (N_21645,N_20724,N_20588);
or U21646 (N_21646,N_21229,N_20013);
and U21647 (N_21647,N_20132,N_20721);
nor U21648 (N_21648,N_20068,N_20798);
nand U21649 (N_21649,N_20540,N_20151);
and U21650 (N_21650,N_20879,N_20307);
nor U21651 (N_21651,N_20156,N_20463);
and U21652 (N_21652,N_20830,N_20454);
or U21653 (N_21653,N_20727,N_20432);
nand U21654 (N_21654,N_20813,N_20179);
and U21655 (N_21655,N_20645,N_20958);
nand U21656 (N_21656,N_20628,N_20869);
xnor U21657 (N_21657,N_20370,N_20444);
and U21658 (N_21658,N_20374,N_20880);
nor U21659 (N_21659,N_20790,N_21099);
and U21660 (N_21660,N_21141,N_20010);
xor U21661 (N_21661,N_21148,N_20261);
and U21662 (N_21662,N_21113,N_20291);
xor U21663 (N_21663,N_20131,N_20472);
or U21664 (N_21664,N_20857,N_20095);
xor U21665 (N_21665,N_20758,N_21111);
or U21666 (N_21666,N_20659,N_20881);
nor U21667 (N_21667,N_20785,N_20037);
nand U21668 (N_21668,N_20051,N_20300);
or U21669 (N_21669,N_20962,N_20893);
or U21670 (N_21670,N_20242,N_20618);
or U21671 (N_21671,N_20021,N_20135);
xnor U21672 (N_21672,N_20602,N_20169);
nand U21673 (N_21673,N_20853,N_21054);
and U21674 (N_21674,N_20819,N_20418);
and U21675 (N_21675,N_20086,N_21016);
and U21676 (N_21676,N_20443,N_20805);
xnor U21677 (N_21677,N_20476,N_20356);
nand U21678 (N_21678,N_21062,N_20898);
xnor U21679 (N_21679,N_20338,N_20097);
nand U21680 (N_21680,N_21121,N_20264);
xnor U21681 (N_21681,N_20290,N_20933);
and U21682 (N_21682,N_20100,N_20125);
or U21683 (N_21683,N_21077,N_20574);
nor U21684 (N_21684,N_21207,N_20810);
xnor U21685 (N_21685,N_20178,N_21071);
and U21686 (N_21686,N_20975,N_20746);
xor U21687 (N_21687,N_20925,N_20564);
and U21688 (N_21688,N_20422,N_21191);
xor U21689 (N_21689,N_20908,N_20047);
and U21690 (N_21690,N_20731,N_20198);
nor U21691 (N_21691,N_21168,N_21188);
and U21692 (N_21692,N_21117,N_20912);
or U21693 (N_21693,N_20469,N_20547);
nor U21694 (N_21694,N_20756,N_21047);
or U21695 (N_21695,N_20787,N_21084);
xnor U21696 (N_21696,N_20275,N_20326);
nand U21697 (N_21697,N_20803,N_20203);
or U21698 (N_21698,N_21201,N_20246);
nor U21699 (N_21699,N_20369,N_20430);
nor U21700 (N_21700,N_20971,N_20215);
or U21701 (N_21701,N_20556,N_20843);
and U21702 (N_21702,N_20641,N_21247);
nor U21703 (N_21703,N_20886,N_21173);
xnor U21704 (N_21704,N_20536,N_21133);
and U21705 (N_21705,N_21045,N_20808);
or U21706 (N_21706,N_20240,N_20740);
nand U21707 (N_21707,N_20025,N_20632);
nand U21708 (N_21708,N_20792,N_20562);
xor U21709 (N_21709,N_20910,N_21066);
or U21710 (N_21710,N_20921,N_20762);
xor U21711 (N_21711,N_20545,N_21096);
nand U21712 (N_21712,N_20055,N_20164);
nand U21713 (N_21713,N_20696,N_20381);
nand U21714 (N_21714,N_20090,N_20427);
nand U21715 (N_21715,N_20421,N_21010);
nor U21716 (N_21716,N_20779,N_20318);
and U21717 (N_21717,N_20867,N_20028);
or U21718 (N_21718,N_20605,N_20563);
or U21719 (N_21719,N_20733,N_20832);
nor U21720 (N_21720,N_20056,N_20649);
nor U21721 (N_21721,N_21230,N_20502);
nor U21722 (N_21722,N_20579,N_20846);
nor U21723 (N_21723,N_20906,N_20436);
nor U21724 (N_21724,N_20580,N_20878);
or U21725 (N_21725,N_20943,N_20735);
nand U21726 (N_21726,N_21026,N_20744);
or U21727 (N_21727,N_20079,N_20298);
nor U21728 (N_21728,N_20998,N_20073);
and U21729 (N_21729,N_20809,N_20230);
xnor U21730 (N_21730,N_21132,N_20730);
xor U21731 (N_21731,N_20567,N_20020);
or U21732 (N_21732,N_20457,N_20390);
xnor U21733 (N_21733,N_20995,N_20316);
and U21734 (N_21734,N_20134,N_20448);
nand U21735 (N_21735,N_20510,N_21098);
or U21736 (N_21736,N_20008,N_20223);
nand U21737 (N_21737,N_20183,N_21091);
xor U21738 (N_21738,N_20623,N_20651);
nor U21739 (N_21739,N_20738,N_20615);
or U21740 (N_21740,N_21089,N_20278);
xor U21741 (N_21741,N_20347,N_21248);
nand U21742 (N_21742,N_21042,N_20955);
or U21743 (N_21743,N_20747,N_20288);
xnor U21744 (N_21744,N_20907,N_20935);
nor U21745 (N_21745,N_21233,N_20403);
nand U21746 (N_21746,N_20498,N_20913);
xor U21747 (N_21747,N_20245,N_20760);
nor U21748 (N_21748,N_20928,N_20688);
nand U21749 (N_21749,N_20964,N_20281);
nand U21750 (N_21750,N_20854,N_20018);
nor U21751 (N_21751,N_20213,N_20487);
or U21752 (N_21752,N_20655,N_21166);
nor U21753 (N_21753,N_20985,N_20144);
and U21754 (N_21754,N_20060,N_21149);
and U21755 (N_21755,N_20313,N_20722);
nand U21756 (N_21756,N_20371,N_20219);
nand U21757 (N_21757,N_20257,N_20894);
nor U21758 (N_21758,N_20048,N_20043);
or U21759 (N_21759,N_21179,N_20033);
nor U21760 (N_21760,N_20101,N_21144);
or U21761 (N_21761,N_20128,N_20227);
and U21762 (N_21762,N_21135,N_20383);
xor U21763 (N_21763,N_20842,N_20621);
nor U21764 (N_21764,N_20939,N_20192);
xnor U21765 (N_21765,N_20270,N_20460);
or U21766 (N_21766,N_21154,N_21165);
nand U21767 (N_21767,N_20022,N_20197);
nor U21768 (N_21768,N_20759,N_21051);
or U21769 (N_21769,N_20470,N_20337);
nand U21770 (N_21770,N_20119,N_20837);
xnor U21771 (N_21771,N_20362,N_21220);
or U21772 (N_21772,N_20656,N_20322);
nor U21773 (N_21773,N_21172,N_20643);
xor U21774 (N_21774,N_21124,N_20375);
or U21775 (N_21775,N_21058,N_20686);
or U21776 (N_21776,N_21057,N_20327);
or U21777 (N_21777,N_20276,N_20162);
nand U21778 (N_21778,N_20297,N_20133);
nor U21779 (N_21779,N_20190,N_21136);
xnor U21780 (N_21780,N_20467,N_20539);
xor U21781 (N_21781,N_20496,N_20114);
or U21782 (N_21782,N_21170,N_20415);
nand U21783 (N_21783,N_21114,N_20034);
xor U21784 (N_21784,N_21199,N_20538);
xnor U21785 (N_21785,N_20522,N_21155);
xor U21786 (N_21786,N_20799,N_21223);
or U21787 (N_21787,N_21195,N_21156);
and U21788 (N_21788,N_20631,N_20844);
nor U21789 (N_21789,N_20449,N_20674);
and U21790 (N_21790,N_21048,N_20059);
and U21791 (N_21791,N_21150,N_21186);
and U21792 (N_21792,N_20340,N_21216);
nor U21793 (N_21793,N_20329,N_20017);
xnor U21794 (N_21794,N_20833,N_20341);
xnor U21795 (N_21795,N_20795,N_20524);
or U21796 (N_21796,N_20796,N_20172);
nand U21797 (N_21797,N_20330,N_20049);
nor U21798 (N_21798,N_20973,N_20395);
xnor U21799 (N_21799,N_20816,N_20677);
or U21800 (N_21800,N_21041,N_20376);
xor U21801 (N_21801,N_20541,N_20992);
or U21802 (N_21802,N_20669,N_20069);
nand U21803 (N_21803,N_20268,N_20603);
xor U21804 (N_21804,N_20776,N_20243);
and U21805 (N_21805,N_20184,N_20410);
and U21806 (N_21806,N_20171,N_20689);
xor U21807 (N_21807,N_20754,N_21194);
and U21808 (N_21808,N_20185,N_21005);
xnor U21809 (N_21809,N_20736,N_20062);
nand U21810 (N_21810,N_20555,N_20703);
or U21811 (N_21811,N_20407,N_20455);
nor U21812 (N_21812,N_20909,N_20937);
nor U21813 (N_21813,N_20099,N_20080);
or U21814 (N_21814,N_20163,N_21162);
xnor U21815 (N_21815,N_20032,N_21013);
and U21816 (N_21816,N_20726,N_21017);
or U21817 (N_21817,N_21227,N_20302);
xnor U21818 (N_21818,N_20439,N_20692);
nand U21819 (N_21819,N_20473,N_20385);
or U21820 (N_21820,N_21158,N_21068);
or U21821 (N_21821,N_20005,N_20182);
nand U21822 (N_21822,N_20103,N_21100);
or U21823 (N_21823,N_20417,N_21211);
nor U21824 (N_21824,N_20712,N_20707);
xor U21825 (N_21825,N_21128,N_20982);
nor U21826 (N_21826,N_20115,N_21143);
nand U21827 (N_21827,N_20859,N_20891);
nor U21828 (N_21828,N_20170,N_20972);
xnor U21829 (N_21829,N_20234,N_20200);
xor U21830 (N_21830,N_20492,N_20389);
nand U21831 (N_21831,N_20697,N_20761);
nor U21832 (N_21832,N_20640,N_20678);
nor U21833 (N_21833,N_20481,N_20616);
and U21834 (N_21834,N_20269,N_20294);
xnor U21835 (N_21835,N_20272,N_20155);
nand U21836 (N_21836,N_20592,N_20835);
nand U21837 (N_21837,N_20897,N_20063);
and U21838 (N_21838,N_20233,N_20000);
and U21839 (N_21839,N_20324,N_20576);
nor U21840 (N_21840,N_21157,N_20543);
nand U21841 (N_21841,N_20309,N_20773);
nor U21842 (N_21842,N_20529,N_20582);
and U21843 (N_21843,N_20566,N_20769);
nand U21844 (N_21844,N_20002,N_20583);
or U21845 (N_21845,N_20825,N_20693);
and U21846 (N_21846,N_20253,N_21072);
nand U21847 (N_21847,N_20981,N_21167);
or U21848 (N_21848,N_20589,N_21192);
nand U21849 (N_21849,N_20348,N_20593);
nor U21850 (N_21850,N_20016,N_20961);
or U21851 (N_21851,N_20429,N_21245);
or U21852 (N_21852,N_20523,N_20775);
nor U21853 (N_21853,N_21129,N_21075);
nand U21854 (N_21854,N_20518,N_20911);
nor U21855 (N_21855,N_20244,N_21115);
or U21856 (N_21856,N_20622,N_20365);
nand U21857 (N_21857,N_20091,N_21035);
and U21858 (N_21858,N_20058,N_20845);
nand U21859 (N_21859,N_20494,N_21221);
and U21860 (N_21860,N_21125,N_21238);
or U21861 (N_21861,N_20464,N_20026);
and U21862 (N_21862,N_20206,N_20087);
nand U21863 (N_21863,N_20420,N_20595);
or U21864 (N_21864,N_20988,N_20959);
and U21865 (N_21865,N_20265,N_20946);
nand U21866 (N_21866,N_20662,N_20781);
nor U21867 (N_21867,N_20408,N_20636);
and U21868 (N_21868,N_20930,N_20914);
and U21869 (N_21869,N_21205,N_20235);
xnor U21870 (N_21870,N_20038,N_20608);
nand U21871 (N_21871,N_20364,N_21110);
and U21872 (N_21872,N_20951,N_20311);
xnor U21873 (N_21873,N_21131,N_20814);
xor U21874 (N_21874,N_20221,N_20360);
xor U21875 (N_21875,N_20251,N_20475);
nor U21876 (N_21876,N_21201,N_20294);
nand U21877 (N_21877,N_20774,N_20525);
nand U21878 (N_21878,N_20008,N_20558);
and U21879 (N_21879,N_20159,N_20634);
nor U21880 (N_21880,N_20870,N_20959);
or U21881 (N_21881,N_20523,N_20597);
nand U21882 (N_21882,N_20845,N_20760);
xnor U21883 (N_21883,N_20829,N_20717);
nand U21884 (N_21884,N_21092,N_20954);
nor U21885 (N_21885,N_20769,N_20435);
xnor U21886 (N_21886,N_21113,N_20940);
xor U21887 (N_21887,N_20556,N_21094);
xor U21888 (N_21888,N_20923,N_21222);
and U21889 (N_21889,N_20216,N_20040);
xor U21890 (N_21890,N_20106,N_20955);
xnor U21891 (N_21891,N_20010,N_20188);
nand U21892 (N_21892,N_20043,N_20335);
or U21893 (N_21893,N_20600,N_20561);
xnor U21894 (N_21894,N_20528,N_20066);
or U21895 (N_21895,N_20689,N_20486);
nor U21896 (N_21896,N_20983,N_20005);
nor U21897 (N_21897,N_20109,N_20187);
nand U21898 (N_21898,N_20071,N_20769);
nand U21899 (N_21899,N_20450,N_20309);
nand U21900 (N_21900,N_20120,N_20069);
nand U21901 (N_21901,N_21218,N_21230);
and U21902 (N_21902,N_20363,N_20511);
nand U21903 (N_21903,N_20533,N_20266);
nand U21904 (N_21904,N_21115,N_20405);
nor U21905 (N_21905,N_20873,N_20288);
xnor U21906 (N_21906,N_21201,N_21042);
or U21907 (N_21907,N_20496,N_20808);
or U21908 (N_21908,N_20683,N_20692);
and U21909 (N_21909,N_20847,N_20927);
or U21910 (N_21910,N_21183,N_20251);
or U21911 (N_21911,N_20980,N_20626);
xnor U21912 (N_21912,N_21065,N_20290);
nand U21913 (N_21913,N_21115,N_20159);
nor U21914 (N_21914,N_21089,N_20560);
nor U21915 (N_21915,N_20299,N_20621);
or U21916 (N_21916,N_20906,N_21060);
and U21917 (N_21917,N_21107,N_20113);
or U21918 (N_21918,N_20707,N_20766);
nand U21919 (N_21919,N_20283,N_20180);
or U21920 (N_21920,N_20905,N_21155);
or U21921 (N_21921,N_21029,N_20969);
xor U21922 (N_21922,N_20608,N_20463);
xor U21923 (N_21923,N_21047,N_20353);
nand U21924 (N_21924,N_20054,N_20273);
nor U21925 (N_21925,N_20837,N_20568);
or U21926 (N_21926,N_20717,N_21223);
xor U21927 (N_21927,N_20802,N_21085);
xnor U21928 (N_21928,N_20163,N_20195);
and U21929 (N_21929,N_20681,N_20809);
xnor U21930 (N_21930,N_20381,N_20910);
nor U21931 (N_21931,N_20445,N_20328);
and U21932 (N_21932,N_21239,N_20521);
nand U21933 (N_21933,N_20000,N_20630);
xnor U21934 (N_21934,N_21187,N_20242);
xnor U21935 (N_21935,N_20785,N_20169);
xnor U21936 (N_21936,N_20849,N_20474);
nor U21937 (N_21937,N_20050,N_21047);
nand U21938 (N_21938,N_21054,N_20397);
and U21939 (N_21939,N_20972,N_20125);
nor U21940 (N_21940,N_21102,N_20426);
and U21941 (N_21941,N_20295,N_20124);
or U21942 (N_21942,N_20332,N_20418);
and U21943 (N_21943,N_20145,N_20747);
and U21944 (N_21944,N_21081,N_21052);
or U21945 (N_21945,N_21185,N_20865);
nor U21946 (N_21946,N_20321,N_20233);
or U21947 (N_21947,N_20748,N_21196);
nor U21948 (N_21948,N_21118,N_20251);
and U21949 (N_21949,N_20642,N_20752);
and U21950 (N_21950,N_20168,N_20603);
and U21951 (N_21951,N_20917,N_20379);
or U21952 (N_21952,N_21026,N_20387);
or U21953 (N_21953,N_20481,N_20036);
nand U21954 (N_21954,N_20422,N_20302);
nand U21955 (N_21955,N_20513,N_20112);
xnor U21956 (N_21956,N_20968,N_20158);
nand U21957 (N_21957,N_20648,N_21064);
xnor U21958 (N_21958,N_20107,N_20661);
or U21959 (N_21959,N_20112,N_21223);
nor U21960 (N_21960,N_21120,N_20742);
or U21961 (N_21961,N_20821,N_20861);
nand U21962 (N_21962,N_20944,N_20652);
and U21963 (N_21963,N_20887,N_20827);
nor U21964 (N_21964,N_20104,N_20613);
xor U21965 (N_21965,N_20092,N_20907);
or U21966 (N_21966,N_20608,N_20383);
xnor U21967 (N_21967,N_20388,N_20037);
xor U21968 (N_21968,N_20775,N_20045);
and U21969 (N_21969,N_20803,N_21011);
and U21970 (N_21970,N_20715,N_20844);
or U21971 (N_21971,N_20099,N_20943);
xor U21972 (N_21972,N_20332,N_20270);
nor U21973 (N_21973,N_20808,N_20351);
nand U21974 (N_21974,N_21007,N_21014);
nor U21975 (N_21975,N_20155,N_21076);
nand U21976 (N_21976,N_20831,N_20391);
and U21977 (N_21977,N_21011,N_20388);
nand U21978 (N_21978,N_20697,N_20152);
or U21979 (N_21979,N_20928,N_20618);
and U21980 (N_21980,N_20242,N_20773);
or U21981 (N_21981,N_20493,N_20761);
nand U21982 (N_21982,N_20249,N_20209);
and U21983 (N_21983,N_20222,N_20711);
and U21984 (N_21984,N_20329,N_20384);
and U21985 (N_21985,N_21118,N_20599);
and U21986 (N_21986,N_20842,N_20193);
or U21987 (N_21987,N_20339,N_20490);
nor U21988 (N_21988,N_20963,N_20160);
and U21989 (N_21989,N_20943,N_20728);
nor U21990 (N_21990,N_21173,N_20202);
nor U21991 (N_21991,N_20287,N_20587);
nand U21992 (N_21992,N_21249,N_20850);
nor U21993 (N_21993,N_20579,N_20435);
and U21994 (N_21994,N_20684,N_20676);
or U21995 (N_21995,N_20645,N_20271);
and U21996 (N_21996,N_20640,N_21093);
nor U21997 (N_21997,N_21133,N_20932);
nand U21998 (N_21998,N_20670,N_20434);
nor U21999 (N_21999,N_20729,N_20229);
nor U22000 (N_22000,N_20878,N_20833);
nand U22001 (N_22001,N_20339,N_20728);
xnor U22002 (N_22002,N_20342,N_20545);
nand U22003 (N_22003,N_20011,N_20348);
nor U22004 (N_22004,N_20457,N_20755);
nand U22005 (N_22005,N_20024,N_20961);
nand U22006 (N_22006,N_20933,N_20265);
nand U22007 (N_22007,N_20105,N_21228);
xor U22008 (N_22008,N_21170,N_20735);
nand U22009 (N_22009,N_20440,N_20291);
and U22010 (N_22010,N_21131,N_20846);
xnor U22011 (N_22011,N_20560,N_20128);
and U22012 (N_22012,N_20396,N_20175);
nand U22013 (N_22013,N_21011,N_20847);
and U22014 (N_22014,N_20527,N_20366);
or U22015 (N_22015,N_20597,N_20065);
nand U22016 (N_22016,N_20159,N_20319);
xor U22017 (N_22017,N_20109,N_20942);
nor U22018 (N_22018,N_20135,N_21179);
xnor U22019 (N_22019,N_21101,N_21084);
xnor U22020 (N_22020,N_20565,N_20583);
nor U22021 (N_22021,N_20484,N_20679);
nand U22022 (N_22022,N_20144,N_21105);
nor U22023 (N_22023,N_20169,N_20376);
nand U22024 (N_22024,N_21071,N_20946);
nand U22025 (N_22025,N_20339,N_20885);
or U22026 (N_22026,N_21060,N_20707);
nor U22027 (N_22027,N_20597,N_20339);
and U22028 (N_22028,N_20247,N_20793);
nor U22029 (N_22029,N_20685,N_20653);
or U22030 (N_22030,N_20529,N_20393);
and U22031 (N_22031,N_20167,N_20769);
xor U22032 (N_22032,N_21084,N_20051);
nor U22033 (N_22033,N_20191,N_20432);
nand U22034 (N_22034,N_20554,N_20961);
xor U22035 (N_22035,N_21141,N_20409);
nand U22036 (N_22036,N_20315,N_20308);
xor U22037 (N_22037,N_20271,N_20138);
xor U22038 (N_22038,N_20328,N_20415);
xnor U22039 (N_22039,N_20086,N_20985);
nor U22040 (N_22040,N_20941,N_21025);
or U22041 (N_22041,N_20341,N_20202);
and U22042 (N_22042,N_20759,N_20053);
and U22043 (N_22043,N_20193,N_21005);
and U22044 (N_22044,N_20985,N_20290);
or U22045 (N_22045,N_20704,N_21235);
nor U22046 (N_22046,N_20717,N_21018);
or U22047 (N_22047,N_20229,N_20014);
nor U22048 (N_22048,N_21190,N_20259);
xnor U22049 (N_22049,N_20460,N_21075);
or U22050 (N_22050,N_20405,N_20794);
nand U22051 (N_22051,N_20052,N_20131);
nand U22052 (N_22052,N_21072,N_20422);
xor U22053 (N_22053,N_20751,N_20951);
and U22054 (N_22054,N_21174,N_20543);
nor U22055 (N_22055,N_20893,N_20205);
and U22056 (N_22056,N_20559,N_20349);
nor U22057 (N_22057,N_20806,N_20671);
nand U22058 (N_22058,N_20174,N_20537);
xor U22059 (N_22059,N_20045,N_20162);
xor U22060 (N_22060,N_20552,N_21197);
nor U22061 (N_22061,N_20401,N_21167);
nand U22062 (N_22062,N_20597,N_21194);
xnor U22063 (N_22063,N_20616,N_20770);
and U22064 (N_22064,N_21249,N_20817);
and U22065 (N_22065,N_20977,N_20377);
nand U22066 (N_22066,N_21198,N_20753);
and U22067 (N_22067,N_20413,N_20877);
xor U22068 (N_22068,N_20816,N_20683);
nand U22069 (N_22069,N_20222,N_20698);
and U22070 (N_22070,N_20309,N_20136);
and U22071 (N_22071,N_20178,N_20115);
nand U22072 (N_22072,N_20670,N_20361);
xnor U22073 (N_22073,N_20305,N_20333);
xnor U22074 (N_22074,N_20784,N_20127);
nor U22075 (N_22075,N_20752,N_20454);
and U22076 (N_22076,N_20313,N_20302);
and U22077 (N_22077,N_20633,N_20277);
or U22078 (N_22078,N_20877,N_20108);
or U22079 (N_22079,N_20509,N_20127);
and U22080 (N_22080,N_20586,N_20438);
nor U22081 (N_22081,N_20478,N_20886);
nor U22082 (N_22082,N_20308,N_20187);
xnor U22083 (N_22083,N_20832,N_20270);
nand U22084 (N_22084,N_21084,N_21153);
nand U22085 (N_22085,N_21126,N_20333);
xnor U22086 (N_22086,N_20872,N_20509);
xor U22087 (N_22087,N_20867,N_21201);
nor U22088 (N_22088,N_20370,N_20854);
and U22089 (N_22089,N_21023,N_20250);
and U22090 (N_22090,N_20287,N_20282);
nor U22091 (N_22091,N_20875,N_20575);
xnor U22092 (N_22092,N_21054,N_20780);
nor U22093 (N_22093,N_20270,N_20645);
nor U22094 (N_22094,N_20867,N_20751);
nand U22095 (N_22095,N_20696,N_20151);
and U22096 (N_22096,N_20920,N_20867);
xnor U22097 (N_22097,N_20902,N_21242);
nor U22098 (N_22098,N_20154,N_20915);
or U22099 (N_22099,N_21104,N_20499);
or U22100 (N_22100,N_20089,N_21229);
xnor U22101 (N_22101,N_21149,N_20103);
or U22102 (N_22102,N_20894,N_20650);
nor U22103 (N_22103,N_20577,N_20050);
and U22104 (N_22104,N_20760,N_21111);
nor U22105 (N_22105,N_21068,N_20188);
nor U22106 (N_22106,N_20938,N_20692);
nor U22107 (N_22107,N_21024,N_21080);
xnor U22108 (N_22108,N_20542,N_20538);
and U22109 (N_22109,N_21004,N_20192);
nor U22110 (N_22110,N_20331,N_20299);
xor U22111 (N_22111,N_20126,N_20279);
nor U22112 (N_22112,N_21242,N_20386);
nor U22113 (N_22113,N_20393,N_20508);
and U22114 (N_22114,N_20630,N_20976);
nor U22115 (N_22115,N_20919,N_20653);
nand U22116 (N_22116,N_20857,N_21211);
and U22117 (N_22117,N_20473,N_21168);
nor U22118 (N_22118,N_20734,N_20449);
nand U22119 (N_22119,N_20774,N_20768);
nand U22120 (N_22120,N_21034,N_21171);
or U22121 (N_22121,N_20011,N_20270);
or U22122 (N_22122,N_20617,N_20548);
xor U22123 (N_22123,N_20108,N_20334);
and U22124 (N_22124,N_20471,N_20840);
or U22125 (N_22125,N_20472,N_21023);
nand U22126 (N_22126,N_20215,N_20995);
nor U22127 (N_22127,N_20341,N_20038);
and U22128 (N_22128,N_21189,N_20470);
nand U22129 (N_22129,N_20353,N_20622);
or U22130 (N_22130,N_20306,N_20313);
xnor U22131 (N_22131,N_20419,N_20461);
nand U22132 (N_22132,N_20009,N_20356);
or U22133 (N_22133,N_20980,N_20631);
and U22134 (N_22134,N_21163,N_21029);
nand U22135 (N_22135,N_20815,N_20877);
xor U22136 (N_22136,N_20164,N_20596);
and U22137 (N_22137,N_20042,N_20597);
nor U22138 (N_22138,N_20743,N_20132);
nor U22139 (N_22139,N_20502,N_20110);
nor U22140 (N_22140,N_21107,N_21175);
nor U22141 (N_22141,N_20767,N_20343);
nor U22142 (N_22142,N_20235,N_20424);
or U22143 (N_22143,N_20075,N_20389);
nor U22144 (N_22144,N_20759,N_20954);
or U22145 (N_22145,N_20736,N_20010);
or U22146 (N_22146,N_20861,N_20074);
or U22147 (N_22147,N_20979,N_20156);
nor U22148 (N_22148,N_20668,N_20186);
nor U22149 (N_22149,N_20714,N_20158);
nor U22150 (N_22150,N_20797,N_21014);
xnor U22151 (N_22151,N_21208,N_20752);
and U22152 (N_22152,N_20693,N_20428);
nand U22153 (N_22153,N_20170,N_20544);
xnor U22154 (N_22154,N_20447,N_20303);
nor U22155 (N_22155,N_20751,N_21227);
or U22156 (N_22156,N_20081,N_20662);
xor U22157 (N_22157,N_20295,N_20438);
nand U22158 (N_22158,N_20357,N_20379);
or U22159 (N_22159,N_20905,N_20361);
xor U22160 (N_22160,N_20913,N_20757);
xor U22161 (N_22161,N_20964,N_20030);
nor U22162 (N_22162,N_20801,N_20713);
or U22163 (N_22163,N_20083,N_20987);
nor U22164 (N_22164,N_20409,N_21049);
and U22165 (N_22165,N_21239,N_20627);
or U22166 (N_22166,N_20176,N_21005);
or U22167 (N_22167,N_20177,N_20516);
nor U22168 (N_22168,N_21100,N_20121);
nand U22169 (N_22169,N_21014,N_21097);
xor U22170 (N_22170,N_20284,N_20685);
or U22171 (N_22171,N_21060,N_20252);
and U22172 (N_22172,N_20129,N_20622);
nor U22173 (N_22173,N_21167,N_20824);
xor U22174 (N_22174,N_20914,N_20452);
nand U22175 (N_22175,N_20472,N_20649);
or U22176 (N_22176,N_20020,N_20622);
nor U22177 (N_22177,N_21221,N_20273);
or U22178 (N_22178,N_20283,N_21058);
or U22179 (N_22179,N_20545,N_20247);
nand U22180 (N_22180,N_21133,N_20733);
and U22181 (N_22181,N_20747,N_20873);
nand U22182 (N_22182,N_20644,N_20633);
and U22183 (N_22183,N_20616,N_20933);
and U22184 (N_22184,N_21184,N_20377);
or U22185 (N_22185,N_20352,N_20419);
xor U22186 (N_22186,N_21048,N_20144);
xor U22187 (N_22187,N_20165,N_20794);
xor U22188 (N_22188,N_20801,N_20307);
and U22189 (N_22189,N_20045,N_21013);
nand U22190 (N_22190,N_20144,N_20532);
xnor U22191 (N_22191,N_21039,N_21249);
nand U22192 (N_22192,N_20252,N_21046);
nand U22193 (N_22193,N_20433,N_20267);
nand U22194 (N_22194,N_20088,N_20418);
and U22195 (N_22195,N_20770,N_21218);
xor U22196 (N_22196,N_20002,N_20139);
nor U22197 (N_22197,N_20966,N_20998);
and U22198 (N_22198,N_20634,N_20419);
xor U22199 (N_22199,N_21217,N_20777);
nand U22200 (N_22200,N_20172,N_20903);
and U22201 (N_22201,N_20372,N_21078);
and U22202 (N_22202,N_20254,N_20803);
or U22203 (N_22203,N_20911,N_20504);
xnor U22204 (N_22204,N_20353,N_21216);
nor U22205 (N_22205,N_20660,N_20144);
xnor U22206 (N_22206,N_20005,N_20938);
or U22207 (N_22207,N_20408,N_20090);
and U22208 (N_22208,N_21127,N_20277);
nor U22209 (N_22209,N_20313,N_21161);
nor U22210 (N_22210,N_20166,N_21071);
nand U22211 (N_22211,N_20341,N_20194);
and U22212 (N_22212,N_20846,N_20158);
nor U22213 (N_22213,N_20653,N_20621);
nand U22214 (N_22214,N_20510,N_20812);
or U22215 (N_22215,N_20428,N_20544);
xor U22216 (N_22216,N_20680,N_20720);
or U22217 (N_22217,N_20640,N_20370);
or U22218 (N_22218,N_20645,N_20022);
and U22219 (N_22219,N_20125,N_20305);
and U22220 (N_22220,N_20723,N_20467);
or U22221 (N_22221,N_20613,N_21133);
or U22222 (N_22222,N_20565,N_21048);
and U22223 (N_22223,N_21142,N_21028);
xor U22224 (N_22224,N_20690,N_20097);
nor U22225 (N_22225,N_20340,N_20997);
nor U22226 (N_22226,N_20585,N_20754);
or U22227 (N_22227,N_20335,N_20173);
or U22228 (N_22228,N_20599,N_21163);
nand U22229 (N_22229,N_20638,N_20424);
or U22230 (N_22230,N_20136,N_20611);
nor U22231 (N_22231,N_20037,N_20390);
or U22232 (N_22232,N_20260,N_20371);
nor U22233 (N_22233,N_20174,N_20731);
or U22234 (N_22234,N_20624,N_21016);
nor U22235 (N_22235,N_20645,N_20178);
xnor U22236 (N_22236,N_21053,N_20515);
or U22237 (N_22237,N_20091,N_20850);
xor U22238 (N_22238,N_20774,N_20536);
nand U22239 (N_22239,N_20238,N_21242);
xor U22240 (N_22240,N_20801,N_20508);
and U22241 (N_22241,N_20816,N_20152);
nor U22242 (N_22242,N_20116,N_20554);
and U22243 (N_22243,N_20411,N_20610);
xnor U22244 (N_22244,N_20929,N_21093);
xor U22245 (N_22245,N_20365,N_20364);
nand U22246 (N_22246,N_20203,N_21151);
or U22247 (N_22247,N_20678,N_20938);
nor U22248 (N_22248,N_20417,N_20285);
nand U22249 (N_22249,N_20374,N_20086);
xor U22250 (N_22250,N_21127,N_21113);
nand U22251 (N_22251,N_20412,N_20505);
and U22252 (N_22252,N_20490,N_20614);
nor U22253 (N_22253,N_20520,N_20727);
nand U22254 (N_22254,N_20239,N_21130);
nand U22255 (N_22255,N_20508,N_20031);
and U22256 (N_22256,N_20148,N_20390);
and U22257 (N_22257,N_20518,N_20584);
nor U22258 (N_22258,N_20781,N_20407);
nor U22259 (N_22259,N_21137,N_21002);
xor U22260 (N_22260,N_20628,N_20023);
nand U22261 (N_22261,N_21019,N_20411);
and U22262 (N_22262,N_21145,N_20589);
nand U22263 (N_22263,N_21208,N_20202);
nand U22264 (N_22264,N_20725,N_20308);
nor U22265 (N_22265,N_20480,N_20795);
and U22266 (N_22266,N_20166,N_20458);
and U22267 (N_22267,N_21154,N_20128);
or U22268 (N_22268,N_20527,N_20511);
or U22269 (N_22269,N_20323,N_20658);
or U22270 (N_22270,N_20217,N_21173);
or U22271 (N_22271,N_20183,N_21123);
xnor U22272 (N_22272,N_20585,N_20893);
or U22273 (N_22273,N_20098,N_20734);
nand U22274 (N_22274,N_20335,N_20876);
xor U22275 (N_22275,N_20395,N_21014);
xnor U22276 (N_22276,N_20305,N_20286);
nand U22277 (N_22277,N_20824,N_20914);
xnor U22278 (N_22278,N_20379,N_20102);
nor U22279 (N_22279,N_20598,N_20692);
nand U22280 (N_22280,N_20320,N_20507);
or U22281 (N_22281,N_21077,N_20578);
nand U22282 (N_22282,N_20847,N_21034);
and U22283 (N_22283,N_20668,N_20637);
and U22284 (N_22284,N_20575,N_20060);
nor U22285 (N_22285,N_21113,N_20836);
and U22286 (N_22286,N_20044,N_20043);
or U22287 (N_22287,N_20448,N_20325);
nand U22288 (N_22288,N_20232,N_21077);
and U22289 (N_22289,N_20190,N_21131);
or U22290 (N_22290,N_20356,N_21192);
or U22291 (N_22291,N_21233,N_20558);
and U22292 (N_22292,N_20101,N_20484);
or U22293 (N_22293,N_20667,N_21243);
xor U22294 (N_22294,N_20393,N_21057);
and U22295 (N_22295,N_21196,N_20700);
nor U22296 (N_22296,N_21223,N_20394);
or U22297 (N_22297,N_21156,N_20218);
nor U22298 (N_22298,N_20542,N_20203);
and U22299 (N_22299,N_20888,N_20128);
nor U22300 (N_22300,N_20103,N_20528);
nor U22301 (N_22301,N_20493,N_20952);
xor U22302 (N_22302,N_20312,N_21073);
nand U22303 (N_22303,N_20189,N_20336);
or U22304 (N_22304,N_20552,N_20179);
or U22305 (N_22305,N_20321,N_20969);
nand U22306 (N_22306,N_20226,N_20463);
nand U22307 (N_22307,N_20908,N_20721);
nand U22308 (N_22308,N_20159,N_20200);
nor U22309 (N_22309,N_20558,N_20279);
xor U22310 (N_22310,N_20055,N_20420);
nand U22311 (N_22311,N_20557,N_20628);
xor U22312 (N_22312,N_20475,N_20392);
nor U22313 (N_22313,N_21045,N_20155);
or U22314 (N_22314,N_21137,N_21036);
and U22315 (N_22315,N_20661,N_20655);
and U22316 (N_22316,N_20254,N_20523);
nor U22317 (N_22317,N_20074,N_20533);
nand U22318 (N_22318,N_20444,N_20204);
nand U22319 (N_22319,N_21057,N_20571);
and U22320 (N_22320,N_21231,N_20336);
or U22321 (N_22321,N_21168,N_20053);
and U22322 (N_22322,N_20029,N_20637);
or U22323 (N_22323,N_21004,N_20875);
and U22324 (N_22324,N_20984,N_20642);
xor U22325 (N_22325,N_20297,N_20117);
and U22326 (N_22326,N_20624,N_20056);
nor U22327 (N_22327,N_20177,N_20017);
xor U22328 (N_22328,N_20959,N_20191);
nor U22329 (N_22329,N_21137,N_20168);
and U22330 (N_22330,N_21041,N_20174);
and U22331 (N_22331,N_20631,N_20439);
xor U22332 (N_22332,N_20596,N_20655);
and U22333 (N_22333,N_21130,N_20916);
and U22334 (N_22334,N_20517,N_20244);
xor U22335 (N_22335,N_21063,N_21110);
nor U22336 (N_22336,N_20493,N_20578);
xor U22337 (N_22337,N_20044,N_20128);
nand U22338 (N_22338,N_20618,N_20749);
xor U22339 (N_22339,N_20885,N_21088);
nor U22340 (N_22340,N_20695,N_20968);
nor U22341 (N_22341,N_20922,N_20783);
nand U22342 (N_22342,N_20071,N_20525);
and U22343 (N_22343,N_20055,N_21241);
nand U22344 (N_22344,N_20436,N_20057);
nand U22345 (N_22345,N_20606,N_20895);
or U22346 (N_22346,N_21184,N_20211);
and U22347 (N_22347,N_20412,N_21032);
xnor U22348 (N_22348,N_20290,N_20650);
nor U22349 (N_22349,N_20363,N_20099);
nand U22350 (N_22350,N_20147,N_20566);
nor U22351 (N_22351,N_20230,N_20854);
and U22352 (N_22352,N_21023,N_20779);
and U22353 (N_22353,N_20458,N_20409);
and U22354 (N_22354,N_20174,N_20733);
and U22355 (N_22355,N_21160,N_21180);
or U22356 (N_22356,N_20230,N_20176);
and U22357 (N_22357,N_20934,N_21079);
nor U22358 (N_22358,N_20454,N_20563);
or U22359 (N_22359,N_20853,N_20940);
and U22360 (N_22360,N_20118,N_20318);
xor U22361 (N_22361,N_21013,N_20599);
and U22362 (N_22362,N_20349,N_20873);
xor U22363 (N_22363,N_20225,N_20034);
nand U22364 (N_22364,N_20195,N_20251);
nor U22365 (N_22365,N_20583,N_21081);
xnor U22366 (N_22366,N_20595,N_20815);
nor U22367 (N_22367,N_20338,N_20291);
or U22368 (N_22368,N_20306,N_20207);
xnor U22369 (N_22369,N_20674,N_20453);
or U22370 (N_22370,N_20367,N_20625);
xor U22371 (N_22371,N_20501,N_20375);
nand U22372 (N_22372,N_20344,N_20629);
nor U22373 (N_22373,N_20654,N_20354);
nand U22374 (N_22374,N_21099,N_20309);
or U22375 (N_22375,N_20345,N_20252);
and U22376 (N_22376,N_20490,N_21116);
nor U22377 (N_22377,N_20330,N_20655);
and U22378 (N_22378,N_21013,N_20842);
or U22379 (N_22379,N_20611,N_20390);
or U22380 (N_22380,N_20220,N_20934);
xnor U22381 (N_22381,N_20512,N_20876);
nor U22382 (N_22382,N_20052,N_20215);
or U22383 (N_22383,N_20862,N_20650);
nand U22384 (N_22384,N_20507,N_20317);
and U22385 (N_22385,N_21009,N_21139);
nand U22386 (N_22386,N_20281,N_20767);
xnor U22387 (N_22387,N_20244,N_20922);
xor U22388 (N_22388,N_21190,N_20142);
nor U22389 (N_22389,N_20913,N_20486);
and U22390 (N_22390,N_20631,N_20646);
nand U22391 (N_22391,N_20152,N_21212);
xor U22392 (N_22392,N_21006,N_20190);
nor U22393 (N_22393,N_20980,N_20043);
or U22394 (N_22394,N_20366,N_21087);
and U22395 (N_22395,N_20317,N_20240);
and U22396 (N_22396,N_20743,N_20226);
nor U22397 (N_22397,N_20291,N_20143);
xnor U22398 (N_22398,N_20967,N_20834);
nor U22399 (N_22399,N_20270,N_20813);
and U22400 (N_22400,N_20205,N_20720);
or U22401 (N_22401,N_21165,N_20775);
xor U22402 (N_22402,N_20117,N_20390);
and U22403 (N_22403,N_20540,N_21195);
nand U22404 (N_22404,N_21181,N_20957);
nor U22405 (N_22405,N_20618,N_20036);
nand U22406 (N_22406,N_21080,N_20936);
xor U22407 (N_22407,N_20115,N_21076);
nor U22408 (N_22408,N_20876,N_21042);
or U22409 (N_22409,N_20903,N_21091);
nor U22410 (N_22410,N_20273,N_21160);
and U22411 (N_22411,N_21205,N_20651);
nor U22412 (N_22412,N_21123,N_21097);
nand U22413 (N_22413,N_20296,N_20758);
and U22414 (N_22414,N_20601,N_20967);
nand U22415 (N_22415,N_20032,N_21190);
nor U22416 (N_22416,N_20465,N_20580);
and U22417 (N_22417,N_20842,N_20111);
or U22418 (N_22418,N_20707,N_20595);
nor U22419 (N_22419,N_20161,N_21099);
or U22420 (N_22420,N_20442,N_21129);
nor U22421 (N_22421,N_20526,N_20134);
and U22422 (N_22422,N_20092,N_20086);
or U22423 (N_22423,N_20291,N_20589);
nor U22424 (N_22424,N_20761,N_20439);
or U22425 (N_22425,N_21170,N_20476);
xor U22426 (N_22426,N_20761,N_21095);
and U22427 (N_22427,N_21064,N_20158);
nor U22428 (N_22428,N_21001,N_20024);
or U22429 (N_22429,N_20831,N_20560);
and U22430 (N_22430,N_21217,N_20548);
nand U22431 (N_22431,N_20984,N_20518);
nand U22432 (N_22432,N_20214,N_20029);
nor U22433 (N_22433,N_20896,N_20025);
or U22434 (N_22434,N_20089,N_20783);
nand U22435 (N_22435,N_21089,N_20949);
nand U22436 (N_22436,N_20754,N_20105);
nand U22437 (N_22437,N_21200,N_20913);
or U22438 (N_22438,N_20745,N_20655);
or U22439 (N_22439,N_20316,N_20339);
xnor U22440 (N_22440,N_20008,N_20526);
or U22441 (N_22441,N_20986,N_20208);
or U22442 (N_22442,N_20497,N_20988);
and U22443 (N_22443,N_20212,N_20486);
and U22444 (N_22444,N_20333,N_20537);
nand U22445 (N_22445,N_20965,N_20301);
nor U22446 (N_22446,N_20736,N_20995);
nand U22447 (N_22447,N_21006,N_20976);
nand U22448 (N_22448,N_21106,N_20734);
xnor U22449 (N_22449,N_20337,N_20692);
and U22450 (N_22450,N_20184,N_20611);
nor U22451 (N_22451,N_21065,N_20422);
xnor U22452 (N_22452,N_20321,N_20362);
and U22453 (N_22453,N_21133,N_21164);
or U22454 (N_22454,N_21127,N_20430);
nor U22455 (N_22455,N_20509,N_21144);
nor U22456 (N_22456,N_20191,N_20093);
nor U22457 (N_22457,N_20545,N_20738);
and U22458 (N_22458,N_20364,N_20481);
nand U22459 (N_22459,N_21155,N_21003);
nand U22460 (N_22460,N_21021,N_21228);
nor U22461 (N_22461,N_20677,N_20167);
and U22462 (N_22462,N_20723,N_20288);
and U22463 (N_22463,N_20788,N_21171);
xnor U22464 (N_22464,N_20951,N_20091);
nand U22465 (N_22465,N_20826,N_20102);
xnor U22466 (N_22466,N_20355,N_20698);
nand U22467 (N_22467,N_20576,N_20685);
and U22468 (N_22468,N_20266,N_20724);
and U22469 (N_22469,N_20830,N_20420);
nor U22470 (N_22470,N_20139,N_20615);
or U22471 (N_22471,N_21085,N_20347);
nand U22472 (N_22472,N_20421,N_20621);
nand U22473 (N_22473,N_21169,N_20621);
nand U22474 (N_22474,N_20981,N_20806);
and U22475 (N_22475,N_20084,N_20633);
xnor U22476 (N_22476,N_21232,N_20132);
nor U22477 (N_22477,N_21238,N_20491);
or U22478 (N_22478,N_20995,N_20710);
nand U22479 (N_22479,N_20488,N_20620);
nand U22480 (N_22480,N_21187,N_21049);
nor U22481 (N_22481,N_20747,N_20312);
and U22482 (N_22482,N_20353,N_20839);
nand U22483 (N_22483,N_20075,N_20448);
nor U22484 (N_22484,N_20470,N_20676);
and U22485 (N_22485,N_21225,N_20893);
or U22486 (N_22486,N_20372,N_20703);
nor U22487 (N_22487,N_20068,N_20670);
xor U22488 (N_22488,N_20843,N_20866);
and U22489 (N_22489,N_20675,N_20187);
nor U22490 (N_22490,N_21128,N_20455);
and U22491 (N_22491,N_20129,N_20111);
xor U22492 (N_22492,N_20855,N_20966);
xnor U22493 (N_22493,N_20838,N_20071);
xnor U22494 (N_22494,N_21023,N_20570);
xor U22495 (N_22495,N_20332,N_21040);
nor U22496 (N_22496,N_20222,N_20719);
xor U22497 (N_22497,N_20735,N_20471);
nand U22498 (N_22498,N_21201,N_21009);
and U22499 (N_22499,N_21218,N_20891);
or U22500 (N_22500,N_22305,N_22024);
and U22501 (N_22501,N_21784,N_21370);
nor U22502 (N_22502,N_22037,N_21651);
or U22503 (N_22503,N_21641,N_21530);
nor U22504 (N_22504,N_21599,N_22252);
nand U22505 (N_22505,N_21267,N_22470);
xnor U22506 (N_22506,N_21503,N_22136);
and U22507 (N_22507,N_22028,N_22464);
nand U22508 (N_22508,N_21494,N_22277);
nor U22509 (N_22509,N_21319,N_21381);
and U22510 (N_22510,N_22055,N_21739);
and U22511 (N_22511,N_21302,N_21282);
nand U22512 (N_22512,N_21378,N_21970);
xor U22513 (N_22513,N_22357,N_22203);
or U22514 (N_22514,N_22057,N_22469);
and U22515 (N_22515,N_21300,N_22406);
or U22516 (N_22516,N_21422,N_22467);
or U22517 (N_22517,N_21813,N_21477);
nand U22518 (N_22518,N_21586,N_22325);
nor U22519 (N_22519,N_21421,N_21407);
or U22520 (N_22520,N_21674,N_21999);
xnor U22521 (N_22521,N_21353,N_22423);
nand U22522 (N_22522,N_22457,N_22010);
and U22523 (N_22523,N_21726,N_22463);
and U22524 (N_22524,N_21350,N_21301);
and U22525 (N_22525,N_21707,N_21334);
or U22526 (N_22526,N_21863,N_22150);
or U22527 (N_22527,N_22283,N_21786);
nor U22528 (N_22528,N_21688,N_21976);
or U22529 (N_22529,N_22090,N_21405);
and U22530 (N_22530,N_21352,N_21317);
xor U22531 (N_22531,N_21522,N_22061);
nor U22532 (N_22532,N_22263,N_22160);
or U22533 (N_22533,N_21584,N_22000);
nand U22534 (N_22534,N_22399,N_21454);
nand U22535 (N_22535,N_21942,N_21995);
xor U22536 (N_22536,N_21724,N_21457);
and U22537 (N_22537,N_22185,N_22494);
xnor U22538 (N_22538,N_21348,N_22431);
or U22539 (N_22539,N_22349,N_21746);
nor U22540 (N_22540,N_22339,N_22419);
nor U22541 (N_22541,N_21515,N_21977);
nand U22542 (N_22542,N_22293,N_21634);
nand U22543 (N_22543,N_22490,N_21495);
nor U22544 (N_22544,N_22096,N_22447);
nor U22545 (N_22545,N_21465,N_21807);
and U22546 (N_22546,N_21329,N_21581);
and U22547 (N_22547,N_22282,N_21671);
or U22548 (N_22548,N_22327,N_22178);
or U22549 (N_22549,N_21616,N_21921);
or U22550 (N_22550,N_22046,N_22340);
or U22551 (N_22551,N_22003,N_21516);
or U22552 (N_22552,N_21573,N_22221);
nand U22553 (N_22553,N_21935,N_21452);
xnor U22554 (N_22554,N_22155,N_21252);
nor U22555 (N_22555,N_22304,N_21964);
nand U22556 (N_22556,N_21768,N_21542);
nand U22557 (N_22557,N_21467,N_21589);
nor U22558 (N_22558,N_22446,N_21489);
nor U22559 (N_22559,N_22246,N_22384);
nand U22560 (N_22560,N_21536,N_22382);
and U22561 (N_22561,N_21974,N_22317);
nor U22562 (N_22562,N_22128,N_22303);
or U22563 (N_22563,N_22402,N_21949);
or U22564 (N_22564,N_22157,N_21758);
xnor U22565 (N_22565,N_21826,N_21720);
and U22566 (N_22566,N_21360,N_21502);
and U22567 (N_22567,N_21272,N_21862);
nand U22568 (N_22568,N_21954,N_21548);
nor U22569 (N_22569,N_22015,N_21366);
nand U22570 (N_22570,N_21534,N_22168);
nand U22571 (N_22571,N_22245,N_21956);
and U22572 (N_22572,N_22443,N_22329);
nand U22573 (N_22573,N_21346,N_22043);
or U22574 (N_22574,N_22104,N_21718);
nand U22575 (N_22575,N_21265,N_21521);
or U22576 (N_22576,N_22313,N_22348);
nand U22577 (N_22577,N_21873,N_22079);
xor U22578 (N_22578,N_21780,N_22275);
or U22579 (N_22579,N_22247,N_21770);
and U22580 (N_22580,N_21982,N_22224);
nor U22581 (N_22581,N_21484,N_21874);
xnor U22582 (N_22582,N_21753,N_22499);
nand U22583 (N_22583,N_21860,N_21670);
nand U22584 (N_22584,N_21391,N_21799);
nor U22585 (N_22585,N_21476,N_21968);
and U22586 (N_22586,N_21590,N_21751);
xnor U22587 (N_22587,N_21686,N_21473);
xor U22588 (N_22588,N_21915,N_21463);
nor U22589 (N_22589,N_21410,N_21565);
and U22590 (N_22590,N_21896,N_22364);
or U22591 (N_22591,N_21506,N_22218);
nor U22592 (N_22592,N_21870,N_21349);
xnor U22593 (N_22593,N_21654,N_22097);
or U22594 (N_22594,N_22065,N_21284);
xnor U22595 (N_22595,N_22425,N_21285);
or U22596 (N_22596,N_21369,N_21700);
and U22597 (N_22597,N_21273,N_22461);
nor U22598 (N_22598,N_22316,N_22021);
nand U22599 (N_22599,N_22146,N_21308);
xor U22600 (N_22600,N_21897,N_21355);
or U22601 (N_22601,N_22139,N_21636);
nand U22602 (N_22602,N_21450,N_22279);
and U22603 (N_22603,N_22385,N_21650);
nor U22604 (N_22604,N_22126,N_22331);
nor U22605 (N_22605,N_21895,N_21655);
or U22606 (N_22606,N_21932,N_21387);
nor U22607 (N_22607,N_22088,N_21434);
and U22608 (N_22608,N_21309,N_22292);
nor U22609 (N_22609,N_21509,N_21673);
xor U22610 (N_22610,N_22174,N_21492);
and U22611 (N_22611,N_21364,N_22239);
or U22612 (N_22612,N_21771,N_22318);
and U22613 (N_22613,N_22177,N_22394);
xnor U22614 (N_22614,N_22085,N_22369);
nor U22615 (N_22615,N_22243,N_21315);
xor U22616 (N_22616,N_21814,N_22397);
nor U22617 (N_22617,N_22105,N_22421);
nor U22618 (N_22618,N_22322,N_22320);
and U22619 (N_22619,N_21851,N_21729);
or U22620 (N_22620,N_22119,N_21250);
and U22621 (N_22621,N_21313,N_21431);
nand U22622 (N_22622,N_21879,N_21512);
or U22623 (N_22623,N_21606,N_21980);
xnor U22624 (N_22624,N_22452,N_21828);
and U22625 (N_22625,N_21871,N_22124);
nand U22626 (N_22626,N_21490,N_21464);
or U22627 (N_22627,N_22092,N_21392);
xnor U22628 (N_22628,N_21850,N_21886);
or U22629 (N_22629,N_22199,N_21772);
nor U22630 (N_22630,N_22188,N_22439);
or U22631 (N_22631,N_22276,N_22413);
or U22632 (N_22632,N_22069,N_21406);
and U22633 (N_22633,N_22241,N_21736);
or U22634 (N_22634,N_21263,N_21526);
or U22635 (N_22635,N_22392,N_22342);
and U22636 (N_22636,N_21507,N_21446);
and U22637 (N_22637,N_21774,N_21842);
nor U22638 (N_22638,N_21816,N_21335);
and U22639 (N_22639,N_22255,N_22307);
nand U22640 (N_22640,N_21764,N_22014);
nor U22641 (N_22641,N_22393,N_22374);
and U22642 (N_22642,N_21679,N_21733);
or U22643 (N_22643,N_21436,N_21281);
nand U22644 (N_22644,N_22491,N_21928);
and U22645 (N_22645,N_21337,N_22290);
nor U22646 (N_22646,N_21695,N_22038);
nor U22647 (N_22647,N_21268,N_21499);
or U22648 (N_22648,N_22341,N_22332);
xnor U22649 (N_22649,N_21640,N_21804);
nand U22650 (N_22650,N_22025,N_21571);
xnor U22651 (N_22651,N_21883,N_21510);
or U22652 (N_22652,N_21680,N_21439);
or U22653 (N_22653,N_21497,N_22023);
xnor U22654 (N_22654,N_21532,N_22445);
or U22655 (N_22655,N_21496,N_21880);
xnor U22656 (N_22656,N_22091,N_22171);
xor U22657 (N_22657,N_22089,N_21778);
or U22658 (N_22658,N_21822,N_21339);
nor U22659 (N_22659,N_22260,N_22344);
or U22660 (N_22660,N_21801,N_21931);
nor U22661 (N_22661,N_21953,N_21630);
or U22662 (N_22662,N_21667,N_22035);
nor U22663 (N_22663,N_21274,N_21519);
xor U22664 (N_22664,N_22248,N_21981);
nor U22665 (N_22665,N_21876,N_21320);
xnor U22666 (N_22666,N_22163,N_22066);
nand U22667 (N_22667,N_21504,N_22179);
or U22668 (N_22668,N_22067,N_22366);
and U22669 (N_22669,N_21330,N_22147);
nand U22670 (N_22670,N_21633,N_21270);
nand U22671 (N_22671,N_21607,N_22296);
nor U22672 (N_22672,N_21908,N_22280);
xor U22673 (N_22673,N_21404,N_21354);
xnor U22674 (N_22674,N_21619,N_21848);
xor U22675 (N_22675,N_21322,N_21692);
xor U22676 (N_22676,N_22440,N_22426);
nand U22677 (N_22677,N_21760,N_22027);
and U22678 (N_22678,N_22080,N_21613);
or U22679 (N_22679,N_21637,N_22272);
and U22680 (N_22680,N_22217,N_22372);
or U22681 (N_22681,N_21371,N_21750);
nand U22682 (N_22682,N_22359,N_22050);
and U22683 (N_22683,N_22148,N_22326);
nand U22684 (N_22684,N_21442,N_21798);
or U22685 (N_22685,N_21419,N_21991);
nor U22686 (N_22686,N_22367,N_22210);
and U22687 (N_22687,N_21259,N_22455);
nor U22688 (N_22688,N_22229,N_21539);
nor U22689 (N_22689,N_21311,N_21545);
nor U22690 (N_22690,N_21417,N_22291);
or U22691 (N_22691,N_21544,N_22338);
and U22692 (N_22692,N_22466,N_22140);
and U22693 (N_22693,N_21893,N_21951);
or U22694 (N_22694,N_22442,N_21668);
and U22695 (N_22695,N_22109,N_21549);
or U22696 (N_22696,N_22295,N_22278);
or U22697 (N_22697,N_21279,N_21971);
nand U22698 (N_22698,N_21540,N_22285);
nor U22699 (N_22699,N_22480,N_22074);
nand U22700 (N_22700,N_21552,N_22053);
and U22701 (N_22701,N_22266,N_21854);
or U22702 (N_22702,N_21911,N_21737);
nor U22703 (N_22703,N_22190,N_21594);
nand U22704 (N_22704,N_21817,N_22030);
or U22705 (N_22705,N_21938,N_21560);
nand U22706 (N_22706,N_21617,N_21550);
or U22707 (N_22707,N_21830,N_21420);
nor U22708 (N_22708,N_21435,N_22125);
xnor U22709 (N_22709,N_21837,N_22093);
xnor U22710 (N_22710,N_21656,N_21967);
nor U22711 (N_22711,N_21691,N_21525);
or U22712 (N_22712,N_21998,N_21644);
xnor U22713 (N_22713,N_21769,N_21832);
or U22714 (N_22714,N_22123,N_21277);
nand U22715 (N_22715,N_21403,N_21925);
and U22716 (N_22716,N_22132,N_22412);
and U22717 (N_22717,N_22441,N_21347);
and U22718 (N_22718,N_21635,N_21757);
or U22719 (N_22719,N_21393,N_21975);
or U22720 (N_22720,N_21759,N_21470);
and U22721 (N_22721,N_21821,N_21430);
nand U22722 (N_22722,N_22206,N_21443);
nor U22723 (N_22723,N_22383,N_21524);
nor U22724 (N_22724,N_21398,N_22100);
nand U22725 (N_22725,N_21914,N_21643);
or U22726 (N_22726,N_22355,N_21962);
and U22727 (N_22727,N_22152,N_21298);
nand U22728 (N_22728,N_21359,N_22267);
nor U22729 (N_22729,N_21264,N_22298);
xnor U22730 (N_22730,N_21557,N_21491);
or U22731 (N_22731,N_22352,N_21683);
nand U22732 (N_22732,N_22401,N_22254);
nand U22733 (N_22733,N_22219,N_21882);
xor U22734 (N_22734,N_22009,N_22005);
nor U22735 (N_22735,N_22118,N_21620);
xnor U22736 (N_22736,N_21262,N_21867);
nand U22737 (N_22737,N_22141,N_21459);
nand U22738 (N_22738,N_21944,N_21388);
xor U22739 (N_22739,N_21779,N_22204);
nor U22740 (N_22740,N_22052,N_21794);
nor U22741 (N_22741,N_21627,N_21414);
xnor U22742 (N_22742,N_22428,N_22004);
nor U22743 (N_22743,N_21919,N_21266);
nand U22744 (N_22744,N_21958,N_21845);
nor U22745 (N_22745,N_22324,N_22134);
nand U22746 (N_22746,N_22236,N_21400);
and U22747 (N_22747,N_21722,N_21864);
xor U22748 (N_22748,N_22368,N_21952);
xor U22749 (N_22749,N_21614,N_21593);
or U22750 (N_22750,N_22182,N_21732);
nand U22751 (N_22751,N_21833,N_21927);
or U22752 (N_22752,N_21642,N_21559);
nand U22753 (N_22753,N_22424,N_21567);
or U22754 (N_22754,N_21752,N_21781);
or U22755 (N_22755,N_21257,N_22437);
nor U22756 (N_22756,N_22197,N_21859);
and U22757 (N_22757,N_21676,N_21909);
xnor U22758 (N_22758,N_21986,N_21961);
or U22759 (N_22759,N_21500,N_21763);
xnor U22760 (N_22760,N_21699,N_21913);
xor U22761 (N_22761,N_22059,N_22208);
nand U22762 (N_22762,N_21289,N_21917);
nor U22763 (N_22763,N_21992,N_22498);
or U22764 (N_22764,N_22175,N_21611);
nor U22765 (N_22765,N_21356,N_21922);
nand U22766 (N_22766,N_21255,N_21415);
nand U22767 (N_22767,N_21802,N_21596);
nand U22768 (N_22768,N_22214,N_21994);
nor U22769 (N_22769,N_21479,N_22319);
nor U22770 (N_22770,N_22205,N_22220);
nand U22771 (N_22771,N_21527,N_22194);
or U22772 (N_22772,N_21844,N_21413);
xnor U22773 (N_22773,N_22429,N_21427);
and U22774 (N_22774,N_21747,N_22172);
nand U22775 (N_22775,N_21456,N_21462);
nor U22776 (N_22776,N_21741,N_22170);
or U22777 (N_22777,N_21541,N_22462);
and U22778 (N_22778,N_22351,N_21743);
or U22779 (N_22779,N_22230,N_22186);
and U22780 (N_22780,N_21866,N_21292);
or U22781 (N_22781,N_22371,N_21943);
and U22782 (N_22782,N_21725,N_21803);
or U22783 (N_22783,N_21978,N_21576);
or U22784 (N_22784,N_21451,N_21610);
nor U22785 (N_22785,N_22063,N_21409);
and U22786 (N_22786,N_22381,N_22191);
nor U22787 (N_22787,N_21299,N_22212);
or U22788 (N_22788,N_21648,N_21959);
nor U22789 (N_22789,N_21835,N_21626);
xor U22790 (N_22790,N_21773,N_21304);
nor U22791 (N_22791,N_22101,N_22213);
nand U22792 (N_22792,N_21416,N_21945);
xor U22793 (N_22793,N_21425,N_21818);
nor U22794 (N_22794,N_22169,N_21973);
and U22795 (N_22795,N_21411,N_21966);
nor U22796 (N_22796,N_21681,N_21710);
nor U22797 (N_22797,N_22225,N_22019);
nor U22798 (N_22798,N_22389,N_22299);
nand U22799 (N_22799,N_21295,N_22207);
xnor U22800 (N_22800,N_22216,N_22485);
nor U22801 (N_22801,N_22151,N_22112);
or U22802 (N_22802,N_22211,N_22311);
and U22803 (N_22803,N_21877,N_22453);
xor U22804 (N_22804,N_22144,N_21251);
nor U22805 (N_22805,N_21703,N_22472);
or U22806 (N_22806,N_21856,N_21554);
nor U22807 (N_22807,N_22111,N_22131);
nand U22808 (N_22808,N_21849,N_21878);
xnor U22809 (N_22809,N_21460,N_21809);
xnor U22810 (N_22810,N_22095,N_21969);
and U22811 (N_22811,N_21468,N_21592);
nand U22812 (N_22812,N_22117,N_22471);
nand U22813 (N_22813,N_22330,N_21579);
nand U22814 (N_22814,N_21664,N_21556);
nand U22815 (N_22815,N_21412,N_22378);
and U22816 (N_22816,N_22084,N_21852);
xnor U22817 (N_22817,N_22071,N_21776);
nand U22818 (N_22818,N_21984,N_21885);
nand U22819 (N_22819,N_21340,N_21918);
xnor U22820 (N_22820,N_21294,N_22232);
and U22821 (N_22821,N_21785,N_22200);
nand U22822 (N_22822,N_22240,N_22082);
and U22823 (N_22823,N_21615,N_22354);
or U22824 (N_22824,N_21881,N_21829);
xnor U22825 (N_22825,N_21365,N_21869);
xor U22826 (N_22826,N_22335,N_22281);
or U22827 (N_22827,N_21312,N_22237);
xor U22828 (N_22828,N_21493,N_21458);
and U22829 (N_22829,N_21820,N_21793);
or U22830 (N_22830,N_21399,N_21649);
nand U22831 (N_22831,N_21326,N_21694);
or U22832 (N_22832,N_22433,N_21865);
or U22833 (N_22833,N_22346,N_21537);
nand U22834 (N_22834,N_21638,N_21936);
and U22835 (N_22835,N_21291,N_21598);
nand U22836 (N_22836,N_22265,N_22184);
xnor U22837 (N_22837,N_21906,N_21677);
nor U22838 (N_22838,N_22400,N_22404);
nor U22839 (N_22839,N_21861,N_22432);
and U22840 (N_22840,N_22395,N_21841);
nand U22841 (N_22841,N_21890,N_21444);
or U22842 (N_22842,N_22031,N_22309);
or U22843 (N_22843,N_22410,N_21333);
nand U22844 (N_22844,N_21629,N_22365);
xnor U22845 (N_22845,N_21904,N_21745);
nand U22846 (N_22846,N_22013,N_22159);
nand U22847 (N_22847,N_22417,N_22405);
or U22848 (N_22848,N_21595,N_21343);
and U22849 (N_22849,N_21395,N_21332);
or U22850 (N_22850,N_22483,N_21934);
nand U22851 (N_22851,N_22409,N_21687);
nor U22852 (N_22852,N_22054,N_21327);
and U22853 (N_22853,N_21811,N_21646);
nand U22854 (N_22854,N_21543,N_22122);
and U22855 (N_22855,N_21709,N_22196);
nor U22856 (N_22856,N_22070,N_21380);
or U22857 (N_22857,N_22235,N_21384);
xnor U22858 (N_22858,N_21305,N_21997);
nand U22859 (N_22859,N_21603,N_21428);
nor U22860 (N_22860,N_21382,N_21386);
nor U22861 (N_22861,N_21993,N_21905);
nor U22862 (N_22862,N_21721,N_22176);
and U22863 (N_22863,N_21675,N_21318);
xnor U22864 (N_22864,N_22193,N_21987);
nand U22865 (N_22865,N_21754,N_22161);
or U22866 (N_22866,N_21253,N_22388);
nor U22867 (N_22867,N_22314,N_21738);
or U22868 (N_22868,N_21310,N_22045);
nor U22869 (N_22869,N_21572,N_22049);
or U22870 (N_22870,N_21702,N_21858);
and U22871 (N_22871,N_21437,N_21765);
nor U22872 (N_22872,N_21455,N_21461);
xor U22873 (N_22873,N_21812,N_22098);
xor U22874 (N_22874,N_22482,N_21666);
or U22875 (N_22875,N_22121,N_22192);
nor U22876 (N_22876,N_22120,N_21609);
xor U22877 (N_22877,N_21792,N_22073);
xor U22878 (N_22878,N_22058,N_21985);
xnor U22879 (N_22879,N_22026,N_22044);
nand U22880 (N_22880,N_21561,N_21625);
nand U22881 (N_22881,N_21892,N_22209);
and U22882 (N_22882,N_21796,N_22142);
and U22883 (N_22883,N_22257,N_22087);
nor U22884 (N_22884,N_21321,N_21508);
nand U22885 (N_22885,N_21296,N_21575);
or U22886 (N_22886,N_22181,N_21704);
nand U22887 (N_22887,N_21390,N_21955);
nand U22888 (N_22888,N_21547,N_21624);
nor U22889 (N_22889,N_21374,N_21731);
or U22890 (N_22890,N_22493,N_21868);
and U22891 (N_22891,N_22183,N_22343);
xor U22892 (N_22892,N_22274,N_21487);
xor U22893 (N_22893,N_22468,N_21853);
nand U22894 (N_22894,N_22001,N_21336);
nand U22895 (N_22895,N_22042,N_21834);
nand U22896 (N_22896,N_21728,N_21480);
and U22897 (N_22897,N_21665,N_22460);
xor U22898 (N_22898,N_21902,N_22064);
xor U22899 (N_22899,N_21795,N_22451);
nor U22900 (N_22900,N_21513,N_22201);
nand U22901 (N_22901,N_21341,N_22475);
xnor U22902 (N_22902,N_22422,N_21564);
nand U22903 (N_22903,N_21363,N_22488);
nand U22904 (N_22904,N_21286,N_21684);
or U22905 (N_22905,N_21505,N_22076);
nor U22906 (N_22906,N_21693,N_21511);
and U22907 (N_22907,N_21888,N_21488);
nand U22908 (N_22908,N_21855,N_21831);
nand U22909 (N_22909,N_21705,N_21587);
and U22910 (N_22910,N_21280,N_21481);
xnor U22911 (N_22911,N_22018,N_21303);
xor U22912 (N_22912,N_21408,N_21325);
or U22913 (N_22913,N_21440,N_22258);
or U22914 (N_22914,N_22473,N_21551);
and U22915 (N_22915,N_22376,N_22353);
nor U22916 (N_22916,N_22062,N_21520);
nor U22917 (N_22917,N_21808,N_22416);
nor U22918 (N_22918,N_21562,N_22008);
and U22919 (N_22919,N_22262,N_21258);
nand U22920 (N_22920,N_21269,N_22379);
or U22921 (N_22921,N_21278,N_21714);
and U22922 (N_22922,N_22036,N_21847);
nand U22923 (N_22923,N_21762,N_21884);
xnor U22924 (N_22924,N_21445,N_21501);
or U22925 (N_22925,N_21658,N_21585);
nor U22926 (N_22926,N_21689,N_21990);
xnor U22927 (N_22927,N_21815,N_21271);
and U22928 (N_22928,N_22006,N_21836);
xnor U22929 (N_22929,N_22138,N_21622);
nor U22930 (N_22930,N_22495,N_21910);
or U22931 (N_22931,N_21518,N_21946);
xnor U22932 (N_22932,N_21730,N_22114);
nand U22933 (N_22933,N_21988,N_21478);
nand U22934 (N_22934,N_22487,N_22328);
or U22935 (N_22935,N_22231,N_21800);
nand U22936 (N_22936,N_22300,N_22187);
nor U22937 (N_22937,N_21657,N_22474);
xor U22938 (N_22938,N_22115,N_21394);
and U22939 (N_22939,N_22040,N_21697);
nand U22940 (N_22940,N_22195,N_21357);
nand U22941 (N_22941,N_21385,N_21602);
or U22942 (N_22942,N_22129,N_21447);
xnor U22943 (N_22943,N_22306,N_21621);
xnor U22944 (N_22944,N_21889,N_21574);
and U22945 (N_22945,N_22337,N_22496);
and U22946 (N_22946,N_22312,N_21466);
nand U22947 (N_22947,N_21623,N_22476);
xor U22948 (N_22948,N_22390,N_22271);
and U22949 (N_22949,N_21577,N_22116);
xnor U22950 (N_22950,N_22198,N_22438);
or U22951 (N_22951,N_21612,N_21756);
xnor U22952 (N_22952,N_22167,N_22249);
or U22953 (N_22953,N_21483,N_22215);
xor U22954 (N_22954,N_22149,N_21361);
xor U22955 (N_22955,N_21344,N_22002);
nand U22956 (N_22956,N_22465,N_21482);
or U22957 (N_22957,N_22007,N_21901);
nand U22958 (N_22958,N_21474,N_22068);
nor U22959 (N_22959,N_22180,N_21486);
nor U22960 (N_22960,N_21661,N_21979);
xor U22961 (N_22961,N_21472,N_21805);
nand U22962 (N_22962,N_21569,N_21723);
or U22963 (N_22963,N_21523,N_22479);
or U22964 (N_22964,N_21789,N_22032);
nor U22965 (N_22965,N_21929,N_22350);
nand U22966 (N_22966,N_22396,N_22398);
xnor U22967 (N_22967,N_21872,N_21947);
nor U22968 (N_22968,N_22427,N_21555);
nand U22969 (N_22969,N_21583,N_21749);
or U22970 (N_22970,N_22264,N_22189);
nor U22971 (N_22971,N_21660,N_22321);
nor U22972 (N_22972,N_21631,N_21735);
and U22973 (N_22973,N_22108,N_22377);
xnor U22974 (N_22974,N_22286,N_22251);
nand U22975 (N_22975,N_21438,N_21256);
and U22976 (N_22976,N_21469,N_21535);
xor U22977 (N_22977,N_21367,N_22336);
nor U22978 (N_22978,N_22259,N_21517);
or U22979 (N_22979,N_21790,N_22238);
or U22980 (N_22980,N_21827,N_21734);
nor U22981 (N_22981,N_21568,N_21608);
and U22982 (N_22982,N_21783,N_22386);
nand U22983 (N_22983,N_21580,N_21429);
nand U22984 (N_22984,N_21426,N_22361);
and U22985 (N_22985,N_22288,N_22156);
nor U22986 (N_22986,N_21690,N_22310);
xor U22987 (N_22987,N_21293,N_22315);
nand U22988 (N_22988,N_21345,N_21423);
nor U22989 (N_22989,N_21432,N_22489);
nand U22990 (N_22990,N_22135,N_22477);
or U22991 (N_22991,N_22086,N_21601);
nand U22992 (N_22992,N_21538,N_21711);
xor U22993 (N_22993,N_21449,N_21351);
and U22994 (N_22994,N_21824,N_21948);
and U22995 (N_22995,N_22020,N_21715);
or U22996 (N_22996,N_21533,N_22102);
nand U22997 (N_22997,N_22387,N_21839);
or U22998 (N_22998,N_21396,N_21713);
or U22999 (N_22999,N_21698,N_22345);
and U23000 (N_23000,N_21900,N_21323);
xor U23001 (N_23001,N_22459,N_21838);
xor U23002 (N_23002,N_21563,N_22273);
or U23003 (N_23003,N_22017,N_22363);
nand U23004 (N_23004,N_21338,N_22164);
nand U23005 (N_23005,N_21960,N_21744);
and U23006 (N_23006,N_22347,N_21659);
nand U23007 (N_23007,N_22408,N_22268);
nor U23008 (N_23008,N_21401,N_21290);
xnor U23009 (N_23009,N_21843,N_21755);
nor U23010 (N_23010,N_21531,N_22244);
nand U23011 (N_23011,N_22041,N_21287);
and U23012 (N_23012,N_22486,N_22078);
or U23013 (N_23013,N_22481,N_21275);
nor U23014 (N_23014,N_21989,N_22250);
nand U23015 (N_23015,N_21939,N_22047);
and U23016 (N_23016,N_22033,N_21618);
or U23017 (N_23017,N_22039,N_22077);
xnor U23018 (N_23018,N_22162,N_22051);
or U23019 (N_23019,N_21924,N_21514);
xnor U23020 (N_23020,N_22403,N_21712);
nand U23021 (N_23021,N_21996,N_21448);
and U23022 (N_23022,N_21254,N_21553);
and U23023 (N_23023,N_22449,N_22233);
and U23024 (N_23024,N_21782,N_21941);
nand U23025 (N_23025,N_22407,N_21887);
or U23026 (N_23026,N_22289,N_22056);
nor U23027 (N_23027,N_22302,N_22034);
or U23028 (N_23028,N_22016,N_21761);
nand U23029 (N_23029,N_21328,N_21306);
nand U23030 (N_23030,N_22458,N_21528);
or U23031 (N_23031,N_21823,N_21940);
nand U23032 (N_23032,N_21600,N_22287);
xor U23033 (N_23033,N_22415,N_21717);
and U23034 (N_23034,N_21260,N_21375);
nand U23035 (N_23035,N_22360,N_21383);
xor U23036 (N_23036,N_22358,N_21570);
or U23037 (N_23037,N_21972,N_21604);
xnor U23038 (N_23038,N_22484,N_21652);
or U23039 (N_23039,N_21840,N_22256);
or U23040 (N_23040,N_22153,N_22418);
nor U23041 (N_23041,N_22110,N_22478);
nor U23042 (N_23042,N_22448,N_21857);
nand U23043 (N_23043,N_22094,N_22492);
nor U23044 (N_23044,N_22420,N_21907);
xor U23045 (N_23045,N_21740,N_22143);
xnor U23046 (N_23046,N_21376,N_22228);
xor U23047 (N_23047,N_21276,N_21358);
nor U23048 (N_23048,N_22436,N_21912);
xor U23049 (N_23049,N_22022,N_21748);
xor U23050 (N_23050,N_22430,N_21708);
xor U23051 (N_23051,N_22012,N_22411);
xor U23052 (N_23052,N_22414,N_21324);
nand U23053 (N_23053,N_21582,N_21632);
nor U23054 (N_23054,N_22301,N_21930);
xor U23055 (N_23055,N_21498,N_21806);
nor U23056 (N_23056,N_21588,N_21727);
xnor U23057 (N_23057,N_22270,N_21788);
and U23058 (N_23058,N_22269,N_21316);
xnor U23059 (N_23059,N_22380,N_21471);
or U23060 (N_23060,N_21402,N_21653);
and U23061 (N_23061,N_21957,N_22099);
nand U23062 (N_23062,N_22356,N_22434);
nand U23063 (N_23063,N_21742,N_21797);
nor U23064 (N_23064,N_21529,N_21372);
nand U23065 (N_23065,N_22107,N_21591);
and U23066 (N_23066,N_21983,N_21342);
nand U23067 (N_23067,N_21926,N_22165);
xor U23068 (N_23068,N_22106,N_21682);
and U23069 (N_23069,N_22154,N_21706);
nand U23070 (N_23070,N_22297,N_21418);
or U23071 (N_23071,N_21362,N_21307);
or U23072 (N_23072,N_21894,N_22294);
nor U23073 (N_23073,N_22234,N_21639);
nand U23074 (N_23074,N_22202,N_21923);
nor U23075 (N_23075,N_21331,N_22333);
or U23076 (N_23076,N_21368,N_22173);
xor U23077 (N_23077,N_21903,N_22456);
or U23078 (N_23078,N_21441,N_21696);
xor U23079 (N_23079,N_21433,N_21558);
nand U23080 (N_23080,N_21891,N_22133);
xnor U23081 (N_23081,N_21678,N_21819);
and U23082 (N_23082,N_21628,N_21647);
nor U23083 (N_23083,N_21933,N_22373);
nand U23084 (N_23084,N_21605,N_21578);
nor U23085 (N_23085,N_21283,N_21701);
and U23086 (N_23086,N_21389,N_22223);
nand U23087 (N_23087,N_21453,N_22454);
xnor U23088 (N_23088,N_22226,N_21672);
nand U23089 (N_23089,N_21373,N_21662);
xor U23090 (N_23090,N_21846,N_21791);
and U23091 (N_23091,N_22060,N_22113);
nor U23092 (N_23092,N_21810,N_21377);
xor U23093 (N_23093,N_22362,N_21898);
xnor U23094 (N_23094,N_21775,N_21963);
xnor U23095 (N_23095,N_21767,N_22137);
and U23096 (N_23096,N_21716,N_22261);
or U23097 (N_23097,N_21669,N_21766);
and U23098 (N_23098,N_22130,N_21379);
or U23099 (N_23099,N_22375,N_22158);
nor U23100 (N_23100,N_21920,N_22323);
xnor U23101 (N_23101,N_21663,N_22072);
nor U23102 (N_23102,N_22127,N_21777);
xor U23103 (N_23103,N_21645,N_21546);
or U23104 (N_23104,N_22029,N_21288);
nor U23105 (N_23105,N_22253,N_21937);
and U23106 (N_23106,N_22242,N_22166);
and U23107 (N_23107,N_21875,N_21787);
or U23108 (N_23108,N_21899,N_21719);
nand U23109 (N_23109,N_22075,N_22391);
xor U23110 (N_23110,N_21424,N_22145);
nand U23111 (N_23111,N_21685,N_22103);
or U23112 (N_23112,N_21297,N_22048);
nand U23113 (N_23113,N_22435,N_22227);
and U23114 (N_23114,N_22497,N_21475);
nand U23115 (N_23115,N_21597,N_22370);
or U23116 (N_23116,N_22222,N_21965);
and U23117 (N_23117,N_21566,N_22011);
nor U23118 (N_23118,N_21916,N_21261);
and U23119 (N_23119,N_21950,N_21397);
or U23120 (N_23120,N_22083,N_22444);
or U23121 (N_23121,N_21485,N_21825);
nor U23122 (N_23122,N_22308,N_21314);
nand U23123 (N_23123,N_22284,N_22081);
or U23124 (N_23124,N_22450,N_22334);
nand U23125 (N_23125,N_22041,N_22223);
nand U23126 (N_23126,N_21555,N_21716);
or U23127 (N_23127,N_22388,N_21376);
nand U23128 (N_23128,N_22044,N_21384);
xnor U23129 (N_23129,N_21829,N_22110);
nor U23130 (N_23130,N_21840,N_21449);
nand U23131 (N_23131,N_21635,N_21493);
and U23132 (N_23132,N_22407,N_22338);
nor U23133 (N_23133,N_21521,N_21786);
xor U23134 (N_23134,N_21634,N_22054);
xor U23135 (N_23135,N_21368,N_21485);
xor U23136 (N_23136,N_21265,N_21655);
nor U23137 (N_23137,N_22397,N_22359);
nor U23138 (N_23138,N_22154,N_22358);
nand U23139 (N_23139,N_21572,N_21357);
nor U23140 (N_23140,N_22359,N_22106);
nand U23141 (N_23141,N_22191,N_22120);
xnor U23142 (N_23142,N_21949,N_21840);
or U23143 (N_23143,N_22395,N_21531);
nor U23144 (N_23144,N_21940,N_21551);
nor U23145 (N_23145,N_21574,N_22491);
nor U23146 (N_23146,N_22444,N_21277);
nor U23147 (N_23147,N_22082,N_22381);
xnor U23148 (N_23148,N_22181,N_21807);
and U23149 (N_23149,N_21654,N_21640);
and U23150 (N_23150,N_21396,N_22084);
nor U23151 (N_23151,N_22448,N_22254);
xor U23152 (N_23152,N_22481,N_21882);
nand U23153 (N_23153,N_22134,N_22401);
or U23154 (N_23154,N_22354,N_21413);
xnor U23155 (N_23155,N_21378,N_21342);
and U23156 (N_23156,N_21677,N_22009);
xnor U23157 (N_23157,N_22423,N_22176);
nand U23158 (N_23158,N_21532,N_21910);
xor U23159 (N_23159,N_21401,N_21810);
and U23160 (N_23160,N_22056,N_21622);
xor U23161 (N_23161,N_21961,N_21701);
and U23162 (N_23162,N_21291,N_21797);
and U23163 (N_23163,N_21827,N_22301);
nor U23164 (N_23164,N_22037,N_22445);
nand U23165 (N_23165,N_21681,N_22494);
and U23166 (N_23166,N_22089,N_22025);
or U23167 (N_23167,N_21830,N_21509);
nand U23168 (N_23168,N_21496,N_21328);
nand U23169 (N_23169,N_21812,N_22017);
nor U23170 (N_23170,N_21872,N_22367);
nor U23171 (N_23171,N_21466,N_21855);
nand U23172 (N_23172,N_21634,N_22030);
xor U23173 (N_23173,N_21573,N_22227);
or U23174 (N_23174,N_22089,N_21626);
xor U23175 (N_23175,N_21578,N_22248);
xor U23176 (N_23176,N_21253,N_22145);
nand U23177 (N_23177,N_21365,N_21412);
or U23178 (N_23178,N_22121,N_22341);
xnor U23179 (N_23179,N_21323,N_22359);
or U23180 (N_23180,N_21649,N_21747);
or U23181 (N_23181,N_22054,N_21603);
xor U23182 (N_23182,N_22310,N_22028);
or U23183 (N_23183,N_21499,N_22242);
nor U23184 (N_23184,N_22190,N_22067);
nor U23185 (N_23185,N_21998,N_22199);
xnor U23186 (N_23186,N_22480,N_21430);
xnor U23187 (N_23187,N_22141,N_22160);
nand U23188 (N_23188,N_22335,N_21802);
and U23189 (N_23189,N_21290,N_22048);
nor U23190 (N_23190,N_22147,N_21490);
or U23191 (N_23191,N_22065,N_22367);
and U23192 (N_23192,N_22394,N_22031);
xor U23193 (N_23193,N_21503,N_22132);
and U23194 (N_23194,N_21743,N_21917);
or U23195 (N_23195,N_21879,N_22095);
nand U23196 (N_23196,N_21317,N_21890);
nor U23197 (N_23197,N_21991,N_22192);
nand U23198 (N_23198,N_22063,N_22103);
nand U23199 (N_23199,N_21550,N_22172);
or U23200 (N_23200,N_22020,N_22238);
nand U23201 (N_23201,N_22205,N_22182);
and U23202 (N_23202,N_21273,N_22105);
or U23203 (N_23203,N_21531,N_21642);
and U23204 (N_23204,N_21885,N_21322);
and U23205 (N_23205,N_21273,N_22406);
and U23206 (N_23206,N_21863,N_22201);
nand U23207 (N_23207,N_21955,N_21602);
or U23208 (N_23208,N_22300,N_21506);
nor U23209 (N_23209,N_22057,N_22430);
nand U23210 (N_23210,N_21276,N_21458);
and U23211 (N_23211,N_21699,N_22314);
nand U23212 (N_23212,N_22305,N_21793);
xor U23213 (N_23213,N_21778,N_21615);
or U23214 (N_23214,N_22092,N_22396);
xnor U23215 (N_23215,N_21281,N_21546);
nand U23216 (N_23216,N_21676,N_21973);
and U23217 (N_23217,N_22158,N_22168);
or U23218 (N_23218,N_22121,N_21951);
nor U23219 (N_23219,N_22463,N_21825);
or U23220 (N_23220,N_22425,N_22309);
or U23221 (N_23221,N_22142,N_21774);
and U23222 (N_23222,N_21256,N_21859);
xnor U23223 (N_23223,N_21381,N_22473);
and U23224 (N_23224,N_21912,N_21713);
nor U23225 (N_23225,N_21381,N_21833);
nand U23226 (N_23226,N_21530,N_21445);
xnor U23227 (N_23227,N_21867,N_21704);
nor U23228 (N_23228,N_22369,N_21714);
and U23229 (N_23229,N_22178,N_22111);
or U23230 (N_23230,N_21254,N_21278);
nor U23231 (N_23231,N_21597,N_22069);
or U23232 (N_23232,N_21729,N_22117);
or U23233 (N_23233,N_21688,N_22396);
or U23234 (N_23234,N_22436,N_21937);
and U23235 (N_23235,N_21819,N_22094);
or U23236 (N_23236,N_21460,N_21770);
and U23237 (N_23237,N_21864,N_22403);
and U23238 (N_23238,N_21597,N_21671);
nor U23239 (N_23239,N_21750,N_22153);
or U23240 (N_23240,N_21874,N_21888);
and U23241 (N_23241,N_21643,N_21771);
nor U23242 (N_23242,N_21648,N_21511);
or U23243 (N_23243,N_21918,N_21656);
nor U23244 (N_23244,N_21902,N_22246);
nor U23245 (N_23245,N_21961,N_21966);
xnor U23246 (N_23246,N_21536,N_21457);
or U23247 (N_23247,N_21832,N_21652);
xnor U23248 (N_23248,N_22174,N_22108);
or U23249 (N_23249,N_22492,N_21254);
or U23250 (N_23250,N_22062,N_22384);
xor U23251 (N_23251,N_21464,N_21527);
xnor U23252 (N_23252,N_21919,N_22096);
xor U23253 (N_23253,N_21755,N_22405);
xnor U23254 (N_23254,N_22010,N_22023);
nor U23255 (N_23255,N_21967,N_21807);
or U23256 (N_23256,N_21825,N_21713);
and U23257 (N_23257,N_21812,N_21384);
nor U23258 (N_23258,N_21421,N_22130);
nor U23259 (N_23259,N_21808,N_21875);
and U23260 (N_23260,N_22370,N_22187);
xor U23261 (N_23261,N_21418,N_21470);
nor U23262 (N_23262,N_22319,N_21372);
nor U23263 (N_23263,N_21368,N_22415);
or U23264 (N_23264,N_21479,N_22233);
nor U23265 (N_23265,N_22122,N_21595);
nand U23266 (N_23266,N_21803,N_21688);
nand U23267 (N_23267,N_22126,N_22122);
nor U23268 (N_23268,N_21478,N_21782);
nand U23269 (N_23269,N_22486,N_22179);
and U23270 (N_23270,N_21415,N_22279);
or U23271 (N_23271,N_21350,N_21730);
nor U23272 (N_23272,N_22408,N_21744);
nand U23273 (N_23273,N_21586,N_22039);
nor U23274 (N_23274,N_21800,N_22057);
and U23275 (N_23275,N_21309,N_22205);
nand U23276 (N_23276,N_22313,N_21299);
nand U23277 (N_23277,N_21775,N_21543);
nor U23278 (N_23278,N_22221,N_21377);
xnor U23279 (N_23279,N_21330,N_21337);
xor U23280 (N_23280,N_21798,N_22496);
and U23281 (N_23281,N_21295,N_22242);
or U23282 (N_23282,N_21681,N_21933);
xor U23283 (N_23283,N_22013,N_21883);
nand U23284 (N_23284,N_21800,N_22411);
nor U23285 (N_23285,N_21649,N_22368);
and U23286 (N_23286,N_21552,N_21486);
xor U23287 (N_23287,N_22018,N_22237);
or U23288 (N_23288,N_21662,N_22214);
or U23289 (N_23289,N_22080,N_22146);
nor U23290 (N_23290,N_21840,N_22083);
nand U23291 (N_23291,N_22233,N_21916);
and U23292 (N_23292,N_21342,N_21548);
xor U23293 (N_23293,N_22209,N_21866);
xnor U23294 (N_23294,N_22492,N_21655);
and U23295 (N_23295,N_21575,N_21562);
and U23296 (N_23296,N_21729,N_21831);
or U23297 (N_23297,N_21495,N_22232);
nor U23298 (N_23298,N_21602,N_21316);
and U23299 (N_23299,N_22168,N_22259);
nor U23300 (N_23300,N_21537,N_21803);
and U23301 (N_23301,N_21296,N_22051);
xor U23302 (N_23302,N_22434,N_22227);
and U23303 (N_23303,N_22212,N_22043);
nor U23304 (N_23304,N_21746,N_21462);
nor U23305 (N_23305,N_21929,N_22044);
or U23306 (N_23306,N_21261,N_21568);
or U23307 (N_23307,N_22075,N_22122);
xor U23308 (N_23308,N_21393,N_21261);
or U23309 (N_23309,N_21537,N_22354);
nand U23310 (N_23310,N_21982,N_21455);
or U23311 (N_23311,N_22067,N_21807);
and U23312 (N_23312,N_21265,N_22226);
nor U23313 (N_23313,N_21453,N_22248);
nor U23314 (N_23314,N_22035,N_21781);
nand U23315 (N_23315,N_21530,N_22194);
nand U23316 (N_23316,N_22339,N_22142);
nand U23317 (N_23317,N_21789,N_22069);
nand U23318 (N_23318,N_21902,N_21885);
or U23319 (N_23319,N_22332,N_21954);
nor U23320 (N_23320,N_21860,N_21768);
or U23321 (N_23321,N_21978,N_22486);
nand U23322 (N_23322,N_21678,N_21728);
nor U23323 (N_23323,N_22147,N_22180);
or U23324 (N_23324,N_22371,N_21453);
nand U23325 (N_23325,N_21638,N_21889);
nor U23326 (N_23326,N_21450,N_22276);
and U23327 (N_23327,N_22140,N_22188);
nor U23328 (N_23328,N_21342,N_21897);
or U23329 (N_23329,N_21492,N_21820);
nand U23330 (N_23330,N_22093,N_21623);
or U23331 (N_23331,N_21272,N_21585);
and U23332 (N_23332,N_22284,N_22302);
and U23333 (N_23333,N_21444,N_22206);
nor U23334 (N_23334,N_22285,N_21432);
nor U23335 (N_23335,N_22153,N_22357);
or U23336 (N_23336,N_21266,N_21431);
xnor U23337 (N_23337,N_21785,N_22427);
nor U23338 (N_23338,N_22292,N_21365);
nand U23339 (N_23339,N_22377,N_22260);
xor U23340 (N_23340,N_22443,N_21319);
or U23341 (N_23341,N_21653,N_21503);
xor U23342 (N_23342,N_22321,N_22158);
nand U23343 (N_23343,N_22061,N_21325);
and U23344 (N_23344,N_21449,N_22020);
xor U23345 (N_23345,N_22228,N_21523);
nand U23346 (N_23346,N_22430,N_21454);
xor U23347 (N_23347,N_21469,N_22078);
and U23348 (N_23348,N_21427,N_21413);
or U23349 (N_23349,N_22182,N_21444);
nor U23350 (N_23350,N_21780,N_21568);
xor U23351 (N_23351,N_21308,N_22344);
xor U23352 (N_23352,N_21447,N_22429);
nor U23353 (N_23353,N_21863,N_21828);
and U23354 (N_23354,N_21712,N_21939);
xor U23355 (N_23355,N_22386,N_22352);
or U23356 (N_23356,N_21741,N_22392);
or U23357 (N_23357,N_21933,N_21461);
nand U23358 (N_23358,N_22145,N_22235);
and U23359 (N_23359,N_22407,N_21458);
and U23360 (N_23360,N_21707,N_22446);
or U23361 (N_23361,N_22304,N_21730);
nand U23362 (N_23362,N_22315,N_22453);
xor U23363 (N_23363,N_21377,N_22400);
or U23364 (N_23364,N_22089,N_21598);
nand U23365 (N_23365,N_22069,N_22374);
nand U23366 (N_23366,N_22246,N_22285);
xor U23367 (N_23367,N_22495,N_21640);
nor U23368 (N_23368,N_21592,N_21595);
xor U23369 (N_23369,N_22462,N_22304);
nand U23370 (N_23370,N_21931,N_21563);
xnor U23371 (N_23371,N_21940,N_22280);
or U23372 (N_23372,N_21683,N_22165);
xnor U23373 (N_23373,N_21408,N_21380);
and U23374 (N_23374,N_21507,N_21869);
nor U23375 (N_23375,N_21385,N_22292);
or U23376 (N_23376,N_21659,N_21687);
and U23377 (N_23377,N_21285,N_21552);
nand U23378 (N_23378,N_22040,N_21771);
xor U23379 (N_23379,N_22274,N_22000);
nor U23380 (N_23380,N_22255,N_21754);
xnor U23381 (N_23381,N_21640,N_21322);
and U23382 (N_23382,N_21548,N_21814);
or U23383 (N_23383,N_21563,N_22423);
or U23384 (N_23384,N_21782,N_21329);
or U23385 (N_23385,N_22287,N_21771);
xor U23386 (N_23386,N_21745,N_21534);
xor U23387 (N_23387,N_21717,N_21513);
nor U23388 (N_23388,N_21405,N_21799);
and U23389 (N_23389,N_21851,N_22168);
and U23390 (N_23390,N_21287,N_21368);
or U23391 (N_23391,N_22028,N_22043);
or U23392 (N_23392,N_21525,N_21716);
xor U23393 (N_23393,N_21754,N_22280);
xor U23394 (N_23394,N_22142,N_22121);
or U23395 (N_23395,N_21778,N_22100);
or U23396 (N_23396,N_22228,N_22391);
or U23397 (N_23397,N_22352,N_21688);
nor U23398 (N_23398,N_21624,N_21302);
and U23399 (N_23399,N_21407,N_21561);
and U23400 (N_23400,N_22233,N_22034);
xor U23401 (N_23401,N_21847,N_21351);
and U23402 (N_23402,N_21840,N_21285);
and U23403 (N_23403,N_22399,N_22364);
xor U23404 (N_23404,N_21714,N_22186);
or U23405 (N_23405,N_22153,N_21660);
nand U23406 (N_23406,N_21299,N_21816);
nor U23407 (N_23407,N_21676,N_21746);
and U23408 (N_23408,N_21626,N_22420);
or U23409 (N_23409,N_22127,N_21910);
xor U23410 (N_23410,N_21871,N_21485);
or U23411 (N_23411,N_22490,N_21340);
or U23412 (N_23412,N_21778,N_21679);
and U23413 (N_23413,N_22278,N_21507);
xnor U23414 (N_23414,N_21429,N_21977);
xnor U23415 (N_23415,N_21885,N_21793);
and U23416 (N_23416,N_21519,N_22439);
nor U23417 (N_23417,N_21447,N_21885);
xnor U23418 (N_23418,N_21477,N_21520);
nor U23419 (N_23419,N_22372,N_21897);
xor U23420 (N_23420,N_22093,N_21988);
xor U23421 (N_23421,N_21355,N_22267);
and U23422 (N_23422,N_22067,N_21872);
nand U23423 (N_23423,N_22029,N_21389);
nor U23424 (N_23424,N_22028,N_22246);
nand U23425 (N_23425,N_21653,N_22023);
and U23426 (N_23426,N_21540,N_21867);
nand U23427 (N_23427,N_21814,N_22145);
xor U23428 (N_23428,N_22353,N_22400);
and U23429 (N_23429,N_22008,N_21554);
xor U23430 (N_23430,N_21850,N_21949);
xor U23431 (N_23431,N_21275,N_21705);
or U23432 (N_23432,N_22036,N_21791);
nor U23433 (N_23433,N_22225,N_22462);
xor U23434 (N_23434,N_21711,N_22271);
and U23435 (N_23435,N_22027,N_22359);
xnor U23436 (N_23436,N_21395,N_21664);
and U23437 (N_23437,N_22360,N_21453);
and U23438 (N_23438,N_22326,N_21307);
and U23439 (N_23439,N_21632,N_22237);
nand U23440 (N_23440,N_22153,N_21521);
or U23441 (N_23441,N_22267,N_21697);
nor U23442 (N_23442,N_22221,N_21919);
xor U23443 (N_23443,N_22385,N_22088);
nor U23444 (N_23444,N_22249,N_21651);
nor U23445 (N_23445,N_21744,N_21432);
xor U23446 (N_23446,N_22298,N_21435);
or U23447 (N_23447,N_21264,N_21872);
or U23448 (N_23448,N_21573,N_21252);
nor U23449 (N_23449,N_21806,N_21550);
nor U23450 (N_23450,N_22180,N_21536);
and U23451 (N_23451,N_21783,N_22276);
or U23452 (N_23452,N_22437,N_21445);
or U23453 (N_23453,N_21434,N_22364);
and U23454 (N_23454,N_22161,N_21441);
nand U23455 (N_23455,N_22150,N_21608);
nand U23456 (N_23456,N_21502,N_21763);
nand U23457 (N_23457,N_21447,N_21802);
nor U23458 (N_23458,N_22226,N_22370);
xnor U23459 (N_23459,N_22403,N_21926);
nand U23460 (N_23460,N_21696,N_22080);
or U23461 (N_23461,N_22011,N_22164);
and U23462 (N_23462,N_22279,N_21469);
nor U23463 (N_23463,N_21796,N_21332);
or U23464 (N_23464,N_21665,N_21267);
nor U23465 (N_23465,N_21283,N_22250);
nor U23466 (N_23466,N_21920,N_22392);
nand U23467 (N_23467,N_22211,N_22125);
or U23468 (N_23468,N_21824,N_21655);
xnor U23469 (N_23469,N_22233,N_22305);
and U23470 (N_23470,N_21703,N_21699);
nor U23471 (N_23471,N_21816,N_21898);
and U23472 (N_23472,N_22117,N_21958);
nor U23473 (N_23473,N_22201,N_21519);
xor U23474 (N_23474,N_22092,N_21717);
nor U23475 (N_23475,N_21824,N_21826);
or U23476 (N_23476,N_21979,N_21328);
and U23477 (N_23477,N_21903,N_22213);
or U23478 (N_23478,N_22043,N_22332);
nand U23479 (N_23479,N_21591,N_22222);
nor U23480 (N_23480,N_22334,N_21859);
xnor U23481 (N_23481,N_21716,N_21493);
and U23482 (N_23482,N_21902,N_21300);
nor U23483 (N_23483,N_21657,N_22095);
nand U23484 (N_23484,N_21726,N_21632);
and U23485 (N_23485,N_22122,N_21531);
or U23486 (N_23486,N_21632,N_21647);
and U23487 (N_23487,N_21920,N_22458);
xor U23488 (N_23488,N_21644,N_21548);
xor U23489 (N_23489,N_21939,N_21912);
nor U23490 (N_23490,N_21337,N_21386);
or U23491 (N_23491,N_21402,N_21472);
nor U23492 (N_23492,N_22380,N_22483);
or U23493 (N_23493,N_21971,N_21659);
nand U23494 (N_23494,N_21293,N_22000);
nand U23495 (N_23495,N_22313,N_21374);
xor U23496 (N_23496,N_22014,N_21842);
nand U23497 (N_23497,N_21593,N_22071);
and U23498 (N_23498,N_21682,N_21379);
xnor U23499 (N_23499,N_21963,N_22206);
nand U23500 (N_23500,N_22309,N_22449);
or U23501 (N_23501,N_22153,N_21456);
xor U23502 (N_23502,N_21711,N_22347);
nand U23503 (N_23503,N_22196,N_22088);
xnor U23504 (N_23504,N_21826,N_22086);
nor U23505 (N_23505,N_21710,N_21348);
nand U23506 (N_23506,N_22184,N_22079);
and U23507 (N_23507,N_21754,N_22102);
and U23508 (N_23508,N_21431,N_21353);
nand U23509 (N_23509,N_21504,N_21761);
and U23510 (N_23510,N_22063,N_21418);
or U23511 (N_23511,N_22052,N_21293);
and U23512 (N_23512,N_21985,N_22372);
nand U23513 (N_23513,N_22133,N_21471);
nand U23514 (N_23514,N_21624,N_22193);
and U23515 (N_23515,N_22290,N_21342);
nand U23516 (N_23516,N_22322,N_22372);
nor U23517 (N_23517,N_21579,N_22369);
nand U23518 (N_23518,N_21396,N_21903);
and U23519 (N_23519,N_22044,N_22017);
nand U23520 (N_23520,N_22129,N_22278);
xnor U23521 (N_23521,N_21464,N_21799);
or U23522 (N_23522,N_22059,N_21796);
xnor U23523 (N_23523,N_21508,N_22375);
and U23524 (N_23524,N_21636,N_22283);
xnor U23525 (N_23525,N_22295,N_22105);
nor U23526 (N_23526,N_22115,N_22047);
nor U23527 (N_23527,N_21880,N_22488);
and U23528 (N_23528,N_21759,N_21780);
and U23529 (N_23529,N_21358,N_21600);
nand U23530 (N_23530,N_21665,N_22262);
xor U23531 (N_23531,N_21479,N_21614);
xor U23532 (N_23532,N_21751,N_21536);
nand U23533 (N_23533,N_21810,N_21494);
nand U23534 (N_23534,N_22337,N_21784);
xnor U23535 (N_23535,N_21644,N_21699);
and U23536 (N_23536,N_21498,N_21516);
xnor U23537 (N_23537,N_21317,N_21301);
nor U23538 (N_23538,N_21445,N_22288);
xnor U23539 (N_23539,N_22021,N_22420);
xor U23540 (N_23540,N_21561,N_21653);
nand U23541 (N_23541,N_21254,N_22367);
nand U23542 (N_23542,N_22438,N_21585);
nand U23543 (N_23543,N_22205,N_21364);
or U23544 (N_23544,N_21526,N_22063);
or U23545 (N_23545,N_22449,N_21620);
and U23546 (N_23546,N_21442,N_22310);
xnor U23547 (N_23547,N_21664,N_21749);
nor U23548 (N_23548,N_21535,N_21259);
and U23549 (N_23549,N_21309,N_22406);
or U23550 (N_23550,N_21622,N_21697);
and U23551 (N_23551,N_21369,N_22374);
nor U23552 (N_23552,N_22230,N_22348);
xor U23553 (N_23553,N_21290,N_21996);
and U23554 (N_23554,N_21589,N_22420);
or U23555 (N_23555,N_21843,N_22477);
nand U23556 (N_23556,N_22208,N_22056);
and U23557 (N_23557,N_22079,N_22366);
or U23558 (N_23558,N_21610,N_22116);
or U23559 (N_23559,N_21718,N_22377);
and U23560 (N_23560,N_21391,N_21888);
nor U23561 (N_23561,N_22205,N_22498);
or U23562 (N_23562,N_21952,N_21502);
nand U23563 (N_23563,N_22055,N_21334);
nand U23564 (N_23564,N_21752,N_22180);
nor U23565 (N_23565,N_22382,N_21824);
or U23566 (N_23566,N_21684,N_22081);
nor U23567 (N_23567,N_21333,N_21534);
xnor U23568 (N_23568,N_21825,N_22414);
xnor U23569 (N_23569,N_22321,N_21682);
nor U23570 (N_23570,N_22126,N_22446);
nor U23571 (N_23571,N_21346,N_21945);
or U23572 (N_23572,N_21388,N_21949);
or U23573 (N_23573,N_22114,N_21363);
xnor U23574 (N_23574,N_22385,N_21315);
or U23575 (N_23575,N_21778,N_21400);
nand U23576 (N_23576,N_21441,N_21517);
nand U23577 (N_23577,N_21764,N_22058);
or U23578 (N_23578,N_22342,N_21492);
nand U23579 (N_23579,N_22421,N_21532);
nand U23580 (N_23580,N_21417,N_21596);
nand U23581 (N_23581,N_21791,N_21932);
nand U23582 (N_23582,N_22382,N_21925);
or U23583 (N_23583,N_22113,N_21597);
nor U23584 (N_23584,N_21774,N_21795);
nor U23585 (N_23585,N_22234,N_22166);
nor U23586 (N_23586,N_21943,N_22298);
and U23587 (N_23587,N_21947,N_21756);
and U23588 (N_23588,N_21808,N_21921);
xor U23589 (N_23589,N_22438,N_22040);
xor U23590 (N_23590,N_21529,N_22263);
nand U23591 (N_23591,N_21390,N_21500);
and U23592 (N_23592,N_22208,N_21669);
or U23593 (N_23593,N_22435,N_21744);
or U23594 (N_23594,N_22200,N_22251);
nor U23595 (N_23595,N_22067,N_21405);
and U23596 (N_23596,N_22313,N_22460);
xnor U23597 (N_23597,N_21493,N_21695);
nand U23598 (N_23598,N_21475,N_21765);
nand U23599 (N_23599,N_22076,N_21932);
and U23600 (N_23600,N_21515,N_22378);
or U23601 (N_23601,N_21316,N_21703);
nand U23602 (N_23602,N_21998,N_21351);
or U23603 (N_23603,N_22372,N_22392);
xnor U23604 (N_23604,N_21925,N_22046);
and U23605 (N_23605,N_21914,N_22408);
and U23606 (N_23606,N_21901,N_21933);
or U23607 (N_23607,N_22257,N_22024);
xnor U23608 (N_23608,N_22050,N_21564);
and U23609 (N_23609,N_21982,N_21643);
nor U23610 (N_23610,N_21773,N_21684);
or U23611 (N_23611,N_21460,N_22412);
nand U23612 (N_23612,N_21352,N_21796);
nor U23613 (N_23613,N_21760,N_21860);
and U23614 (N_23614,N_21608,N_22303);
nor U23615 (N_23615,N_21577,N_22298);
nand U23616 (N_23616,N_21606,N_21361);
nor U23617 (N_23617,N_21333,N_21490);
and U23618 (N_23618,N_21988,N_21875);
nand U23619 (N_23619,N_22005,N_21476);
xor U23620 (N_23620,N_21728,N_21717);
or U23621 (N_23621,N_22240,N_21572);
or U23622 (N_23622,N_21677,N_21897);
nand U23623 (N_23623,N_22024,N_22384);
nor U23624 (N_23624,N_21290,N_21428);
nand U23625 (N_23625,N_21691,N_21831);
nand U23626 (N_23626,N_21374,N_22045);
or U23627 (N_23627,N_21347,N_22001);
nor U23628 (N_23628,N_22133,N_22344);
xnor U23629 (N_23629,N_21744,N_22282);
or U23630 (N_23630,N_21766,N_22184);
nor U23631 (N_23631,N_22344,N_21752);
nand U23632 (N_23632,N_21888,N_21922);
nand U23633 (N_23633,N_21361,N_21390);
nor U23634 (N_23634,N_22481,N_21302);
or U23635 (N_23635,N_21362,N_21779);
nor U23636 (N_23636,N_22277,N_21381);
or U23637 (N_23637,N_21515,N_22093);
or U23638 (N_23638,N_21710,N_21530);
xor U23639 (N_23639,N_21251,N_21439);
and U23640 (N_23640,N_21294,N_22217);
or U23641 (N_23641,N_21281,N_22364);
nand U23642 (N_23642,N_22047,N_21293);
xnor U23643 (N_23643,N_21848,N_21940);
nand U23644 (N_23644,N_21379,N_21483);
nand U23645 (N_23645,N_21722,N_21501);
xnor U23646 (N_23646,N_22114,N_21309);
xor U23647 (N_23647,N_21882,N_21805);
nor U23648 (N_23648,N_21313,N_21657);
and U23649 (N_23649,N_22077,N_21460);
nor U23650 (N_23650,N_22026,N_21428);
xor U23651 (N_23651,N_21695,N_22233);
xor U23652 (N_23652,N_21894,N_21816);
or U23653 (N_23653,N_22278,N_21289);
nand U23654 (N_23654,N_22485,N_22409);
xor U23655 (N_23655,N_21395,N_22250);
nor U23656 (N_23656,N_21349,N_22270);
xor U23657 (N_23657,N_21931,N_22380);
nor U23658 (N_23658,N_21291,N_21603);
and U23659 (N_23659,N_22384,N_22032);
nor U23660 (N_23660,N_21858,N_21491);
or U23661 (N_23661,N_21366,N_22429);
or U23662 (N_23662,N_21869,N_22115);
and U23663 (N_23663,N_21308,N_22437);
and U23664 (N_23664,N_21431,N_22143);
nor U23665 (N_23665,N_21587,N_21633);
nand U23666 (N_23666,N_21696,N_21373);
and U23667 (N_23667,N_22152,N_21873);
or U23668 (N_23668,N_21961,N_21319);
or U23669 (N_23669,N_21984,N_21733);
xor U23670 (N_23670,N_21936,N_21434);
nor U23671 (N_23671,N_22478,N_21251);
and U23672 (N_23672,N_21265,N_22334);
nand U23673 (N_23673,N_21258,N_22011);
or U23674 (N_23674,N_22494,N_21908);
or U23675 (N_23675,N_21773,N_22132);
and U23676 (N_23676,N_21339,N_22486);
nor U23677 (N_23677,N_22151,N_21712);
xor U23678 (N_23678,N_22416,N_21576);
or U23679 (N_23679,N_21925,N_21521);
or U23680 (N_23680,N_22218,N_21376);
nand U23681 (N_23681,N_21969,N_22336);
nor U23682 (N_23682,N_21760,N_22037);
and U23683 (N_23683,N_22300,N_22038);
nor U23684 (N_23684,N_22393,N_21941);
xor U23685 (N_23685,N_22146,N_21523);
nor U23686 (N_23686,N_21305,N_22327);
or U23687 (N_23687,N_21839,N_21440);
and U23688 (N_23688,N_21413,N_22044);
nor U23689 (N_23689,N_22157,N_21426);
and U23690 (N_23690,N_22020,N_21837);
xor U23691 (N_23691,N_22311,N_22385);
or U23692 (N_23692,N_22198,N_21525);
nor U23693 (N_23693,N_22342,N_21776);
or U23694 (N_23694,N_22245,N_21922);
nand U23695 (N_23695,N_22473,N_21419);
or U23696 (N_23696,N_22303,N_22215);
nand U23697 (N_23697,N_21544,N_21653);
xor U23698 (N_23698,N_21429,N_22414);
xor U23699 (N_23699,N_22131,N_21566);
xor U23700 (N_23700,N_21794,N_21341);
and U23701 (N_23701,N_22318,N_21421);
xnor U23702 (N_23702,N_22047,N_21775);
nand U23703 (N_23703,N_21833,N_21604);
or U23704 (N_23704,N_21735,N_21437);
or U23705 (N_23705,N_21372,N_21986);
nor U23706 (N_23706,N_21834,N_21870);
xor U23707 (N_23707,N_22025,N_22382);
nand U23708 (N_23708,N_22129,N_22093);
nor U23709 (N_23709,N_21822,N_22120);
nor U23710 (N_23710,N_21290,N_22364);
nand U23711 (N_23711,N_21853,N_21359);
nor U23712 (N_23712,N_22067,N_21789);
and U23713 (N_23713,N_21744,N_21940);
or U23714 (N_23714,N_21486,N_21960);
nand U23715 (N_23715,N_21681,N_22407);
and U23716 (N_23716,N_21790,N_21784);
or U23717 (N_23717,N_21969,N_21789);
and U23718 (N_23718,N_21386,N_21668);
xor U23719 (N_23719,N_21450,N_22498);
nand U23720 (N_23720,N_21497,N_22065);
and U23721 (N_23721,N_21323,N_21563);
and U23722 (N_23722,N_22145,N_21872);
nand U23723 (N_23723,N_22102,N_22388);
nand U23724 (N_23724,N_21804,N_21612);
and U23725 (N_23725,N_21637,N_22184);
or U23726 (N_23726,N_21622,N_21359);
nand U23727 (N_23727,N_22469,N_21426);
or U23728 (N_23728,N_22385,N_21728);
or U23729 (N_23729,N_22381,N_21885);
and U23730 (N_23730,N_22086,N_22291);
nor U23731 (N_23731,N_21287,N_22476);
and U23732 (N_23732,N_22017,N_21631);
or U23733 (N_23733,N_21527,N_21542);
nor U23734 (N_23734,N_21658,N_21905);
or U23735 (N_23735,N_22361,N_21970);
or U23736 (N_23736,N_21812,N_21569);
xor U23737 (N_23737,N_21731,N_22013);
and U23738 (N_23738,N_21646,N_21483);
xnor U23739 (N_23739,N_22250,N_22470);
xnor U23740 (N_23740,N_21311,N_21643);
and U23741 (N_23741,N_21760,N_21641);
and U23742 (N_23742,N_21557,N_21621);
or U23743 (N_23743,N_21371,N_21262);
nor U23744 (N_23744,N_21713,N_21950);
nor U23745 (N_23745,N_21368,N_21488);
or U23746 (N_23746,N_21339,N_22493);
nor U23747 (N_23747,N_22429,N_22306);
nand U23748 (N_23748,N_22019,N_21351);
nor U23749 (N_23749,N_22363,N_21290);
nor U23750 (N_23750,N_23250,N_22617);
xnor U23751 (N_23751,N_22511,N_23583);
xnor U23752 (N_23752,N_23343,N_22592);
or U23753 (N_23753,N_22979,N_23216);
or U23754 (N_23754,N_23595,N_22889);
or U23755 (N_23755,N_22637,N_23081);
or U23756 (N_23756,N_23499,N_22639);
or U23757 (N_23757,N_22794,N_23197);
or U23758 (N_23758,N_23233,N_22585);
nand U23759 (N_23759,N_22700,N_23154);
or U23760 (N_23760,N_23692,N_23373);
or U23761 (N_23761,N_22580,N_23385);
nand U23762 (N_23762,N_23516,N_22613);
and U23763 (N_23763,N_23333,N_22551);
nand U23764 (N_23764,N_22542,N_23243);
or U23765 (N_23765,N_23533,N_22923);
or U23766 (N_23766,N_22936,N_23132);
and U23767 (N_23767,N_23658,N_23178);
nor U23768 (N_23768,N_23422,N_22833);
nor U23769 (N_23769,N_23183,N_23646);
nor U23770 (N_23770,N_22736,N_22912);
and U23771 (N_23771,N_22694,N_23127);
and U23772 (N_23772,N_23540,N_22876);
xnor U23773 (N_23773,N_23337,N_23372);
and U23774 (N_23774,N_23040,N_22775);
nand U23775 (N_23775,N_23245,N_23518);
nor U23776 (N_23776,N_22944,N_23689);
xnor U23777 (N_23777,N_23306,N_23211);
and U23778 (N_23778,N_22754,N_23588);
and U23779 (N_23779,N_23220,N_22558);
nor U23780 (N_23780,N_23443,N_23574);
or U23781 (N_23781,N_23485,N_23078);
xor U23782 (N_23782,N_23342,N_23427);
or U23783 (N_23783,N_23545,N_22610);
or U23784 (N_23784,N_22763,N_23137);
and U23785 (N_23785,N_22947,N_22892);
and U23786 (N_23786,N_22727,N_23575);
nand U23787 (N_23787,N_22945,N_23339);
nor U23788 (N_23788,N_22665,N_23676);
or U23789 (N_23789,N_23476,N_23323);
or U23790 (N_23790,N_23152,N_23394);
nor U23791 (N_23791,N_23696,N_23455);
or U23792 (N_23792,N_23087,N_22813);
nor U23793 (N_23793,N_23021,N_23043);
and U23794 (N_23794,N_23269,N_23527);
or U23795 (N_23795,N_22631,N_22744);
and U23796 (N_23796,N_23679,N_22709);
xnor U23797 (N_23797,N_23366,N_23254);
and U23798 (N_23798,N_22955,N_22629);
and U23799 (N_23799,N_23730,N_23016);
nand U23800 (N_23800,N_23426,N_23346);
and U23801 (N_23801,N_23633,N_22952);
nand U23802 (N_23802,N_23252,N_22850);
or U23803 (N_23803,N_22903,N_23118);
xor U23804 (N_23804,N_22735,N_23209);
nor U23805 (N_23805,N_22984,N_23739);
nor U23806 (N_23806,N_23454,N_23713);
xor U23807 (N_23807,N_23514,N_22674);
and U23808 (N_23808,N_23393,N_23542);
xnor U23809 (N_23809,N_23093,N_23044);
nand U23810 (N_23810,N_22960,N_23004);
or U23811 (N_23811,N_22968,N_23601);
xor U23812 (N_23812,N_22662,N_22910);
xnor U23813 (N_23813,N_22759,N_23557);
xnor U23814 (N_23814,N_22915,N_23684);
nand U23815 (N_23815,N_23203,N_22670);
xor U23816 (N_23816,N_22962,N_22913);
xor U23817 (N_23817,N_23065,N_22824);
nor U23818 (N_23818,N_23624,N_22619);
nor U23819 (N_23819,N_22855,N_22501);
and U23820 (N_23820,N_22796,N_23423);
nand U23821 (N_23821,N_22921,N_23212);
nor U23822 (N_23822,N_22967,N_23412);
and U23823 (N_23823,N_23215,N_23456);
or U23824 (N_23824,N_22929,N_23651);
nor U23825 (N_23825,N_22842,N_23086);
and U23826 (N_23826,N_23039,N_23429);
nand U23827 (N_23827,N_23502,N_23331);
nor U23828 (N_23828,N_22917,N_23058);
or U23829 (N_23829,N_22684,N_23210);
xnor U23830 (N_23830,N_23523,N_22618);
nand U23831 (N_23831,N_23280,N_22728);
nand U23832 (N_23832,N_22982,N_23508);
nor U23833 (N_23833,N_23510,N_22788);
and U23834 (N_23834,N_22989,N_23461);
xnor U23835 (N_23835,N_23128,N_22816);
or U23836 (N_23836,N_23293,N_22653);
or U23837 (N_23837,N_22598,N_23555);
or U23838 (N_23838,N_23386,N_22739);
nor U23839 (N_23839,N_23726,N_23591);
xor U23840 (N_23840,N_23258,N_23031);
nor U23841 (N_23841,N_23396,N_23490);
nand U23842 (N_23842,N_22671,N_23176);
or U23843 (N_23843,N_23101,N_22589);
or U23844 (N_23844,N_23489,N_22885);
or U23845 (N_23845,N_22612,N_23434);
and U23846 (N_23846,N_22931,N_23678);
nor U23847 (N_23847,N_23486,N_22904);
nor U23848 (N_23848,N_22607,N_23578);
or U23849 (N_23849,N_23656,N_23749);
nand U23850 (N_23850,N_22958,N_22741);
xnor U23851 (N_23851,N_23003,N_22840);
or U23852 (N_23852,N_23570,N_22822);
nand U23853 (N_23853,N_22819,N_23246);
xor U23854 (N_23854,N_23232,N_23159);
nor U23855 (N_23855,N_22680,N_23134);
nand U23856 (N_23856,N_22748,N_22811);
nor U23857 (N_23857,N_23096,N_23147);
or U23858 (N_23858,N_23686,N_22622);
nand U23859 (N_23859,N_22557,N_22559);
nand U23860 (N_23860,N_22996,N_23654);
or U23861 (N_23861,N_23582,N_23513);
nand U23862 (N_23862,N_23076,N_22737);
xor U23863 (N_23863,N_22578,N_23504);
xor U23864 (N_23864,N_22865,N_22721);
nor U23865 (N_23865,N_23312,N_22869);
or U23866 (N_23866,N_23630,N_22550);
nor U23867 (N_23867,N_23369,N_22724);
nand U23868 (N_23868,N_22647,N_23036);
or U23869 (N_23869,N_22645,N_22999);
nor U23870 (N_23870,N_23556,N_22519);
or U23871 (N_23871,N_23284,N_23612);
or U23872 (N_23872,N_22704,N_22851);
xor U23873 (N_23873,N_22650,N_22713);
nand U23874 (N_23874,N_22986,N_22976);
nand U23875 (N_23875,N_23094,N_22560);
xnor U23876 (N_23876,N_22978,N_23669);
or U23877 (N_23877,N_23395,N_23435);
nand U23878 (N_23878,N_23472,N_23225);
nand U23879 (N_23879,N_23090,N_23073);
nor U23880 (N_23880,N_22895,N_22537);
and U23881 (N_23881,N_23112,N_23607);
and U23882 (N_23882,N_23193,N_23347);
xor U23883 (N_23883,N_23136,N_23149);
nor U23884 (N_23884,N_23162,N_23433);
nor U23885 (N_23885,N_23281,N_23022);
nand U23886 (N_23886,N_23300,N_22926);
or U23887 (N_23887,N_23332,N_22866);
nand U23888 (N_23888,N_23301,N_23494);
or U23889 (N_23889,N_23025,N_22594);
nand U23890 (N_23890,N_22690,N_22563);
xor U23891 (N_23891,N_23388,N_22994);
and U23892 (N_23892,N_22946,N_23470);
xnor U23893 (N_23893,N_23357,N_23050);
and U23894 (N_23894,N_22988,N_22676);
and U23895 (N_23895,N_22579,N_23549);
nor U23896 (N_23896,N_23637,N_22868);
nor U23897 (N_23897,N_23509,N_23054);
nand U23898 (N_23898,N_23060,N_22689);
xnor U23899 (N_23899,N_22992,N_23133);
xnor U23900 (N_23900,N_23439,N_23348);
and U23901 (N_23901,N_23010,N_22538);
and U23902 (N_23902,N_22871,N_22693);
or U23903 (N_23903,N_23092,N_22649);
xor U23904 (N_23904,N_23088,N_23084);
and U23905 (N_23905,N_23617,N_23404);
xor U23906 (N_23906,N_23604,N_23413);
xnor U23907 (N_23907,N_22932,N_23030);
or U23908 (N_23908,N_22515,N_23736);
and U23909 (N_23909,N_23401,N_23157);
xnor U23910 (N_23910,N_22827,N_22858);
and U23911 (N_23911,N_23299,N_23244);
nor U23912 (N_23912,N_22518,N_23642);
and U23913 (N_23913,N_23314,N_23720);
xnor U23914 (N_23914,N_22879,N_22933);
nor U23915 (N_23915,N_22660,N_22841);
xnor U23916 (N_23916,N_22657,N_23445);
or U23917 (N_23917,N_22964,N_23308);
or U23918 (N_23918,N_23321,N_23727);
nand U23919 (N_23919,N_22935,N_22862);
nor U23920 (N_23920,N_23070,N_22596);
or U23921 (N_23921,N_22643,N_22907);
xor U23922 (N_23922,N_22626,N_23632);
nand U23923 (N_23923,N_23375,N_23398);
nand U23924 (N_23924,N_22784,N_23098);
or U23925 (N_23925,N_22859,N_23316);
nor U23926 (N_23926,N_22717,N_22528);
nand U23927 (N_23927,N_22742,N_22891);
nor U23928 (N_23928,N_22747,N_23095);
xor U23929 (N_23929,N_23307,N_23265);
nand U23930 (N_23930,N_22983,N_23069);
nand U23931 (N_23931,N_23140,N_22821);
and U23932 (N_23932,N_23217,N_22768);
nand U23933 (N_23933,N_22663,N_23155);
or U23934 (N_23934,N_23351,N_23344);
and U23935 (N_23935,N_23440,N_23519);
or U23936 (N_23936,N_22549,N_22534);
nand U23937 (N_23937,N_23666,N_23041);
or U23938 (N_23938,N_22793,N_23599);
or U23939 (N_23939,N_23013,N_23493);
nor U23940 (N_23940,N_23263,N_23639);
or U23941 (N_23941,N_22817,N_22635);
nand U23942 (N_23942,N_23554,N_23629);
nor U23943 (N_23943,N_23732,N_23625);
and U23944 (N_23944,N_23548,N_23546);
and U23945 (N_23945,N_22605,N_23558);
xor U23946 (N_23946,N_23536,N_23449);
nor U23947 (N_23947,N_23677,N_23479);
and U23948 (N_23948,N_23644,N_22815);
xor U23949 (N_23949,N_23643,N_23109);
nand U23950 (N_23950,N_22990,N_22730);
nand U23951 (N_23951,N_22648,N_22750);
nand U23952 (N_23952,N_23738,N_22583);
nor U23953 (N_23953,N_23349,N_22658);
or U23954 (N_23954,N_23709,N_23146);
nor U23955 (N_23955,N_23636,N_22908);
xor U23956 (N_23956,N_23023,N_23083);
nor U23957 (N_23957,N_23274,N_23444);
and U23958 (N_23958,N_23606,N_22701);
xor U23959 (N_23959,N_22569,N_23613);
nand U23960 (N_23960,N_22924,N_23560);
xnor U23961 (N_23961,N_23418,N_23011);
nor U23962 (N_23962,N_23694,N_23029);
or U23963 (N_23963,N_22599,N_23327);
and U23964 (N_23964,N_23487,N_22524);
and U23965 (N_23965,N_22529,N_22826);
xor U23966 (N_23966,N_22587,N_23330);
or U23967 (N_23967,N_23743,N_23723);
or U23968 (N_23968,N_23102,N_22593);
or U23969 (N_23969,N_23206,N_22685);
or U23970 (N_23970,N_23057,N_22812);
nand U23971 (N_23971,N_23014,N_22893);
nand U23972 (N_23972,N_23729,N_23020);
or U23973 (N_23973,N_23103,N_23428);
or U23974 (N_23974,N_22957,N_23261);
xor U23975 (N_23975,N_23391,N_23724);
or U23976 (N_23976,N_23585,N_23621);
and U23977 (N_23977,N_23198,N_22877);
nor U23978 (N_23978,N_23139,N_23240);
xnor U23979 (N_23979,N_23038,N_22998);
and U23980 (N_23980,N_23695,N_23701);
and U23981 (N_23981,N_23492,N_23408);
xor U23982 (N_23982,N_23066,N_23521);
and U23983 (N_23983,N_22867,N_23600);
xor U23984 (N_23984,N_23051,N_23111);
xor U23985 (N_23985,N_23202,N_23026);
and U23986 (N_23986,N_23324,N_22546);
and U23987 (N_23987,N_23698,N_23056);
and U23988 (N_23988,N_22654,N_23411);
nor U23989 (N_23989,N_23497,N_23416);
xnor U23990 (N_23990,N_22975,N_23541);
or U23991 (N_23991,N_22834,N_23747);
xnor U23992 (N_23992,N_22852,N_22881);
or U23993 (N_23993,N_23593,N_23603);
xnor U23994 (N_23994,N_23657,N_22584);
nor U23995 (N_23995,N_22807,N_22521);
and U23996 (N_23996,N_22995,N_23682);
and U23997 (N_23997,N_22603,N_23231);
and U23998 (N_23998,N_22734,N_22516);
xnor U23999 (N_23999,N_23392,N_23460);
xnor U24000 (N_24000,N_22634,N_23230);
or U24001 (N_24001,N_23638,N_23442);
or U24002 (N_24002,N_23213,N_23336);
nand U24003 (N_24003,N_22940,N_22508);
or U24004 (N_24004,N_23352,N_23688);
nor U24005 (N_24005,N_22843,N_23242);
or U24006 (N_24006,N_23129,N_23594);
nor U24007 (N_24007,N_22513,N_22753);
and U24008 (N_24008,N_23655,N_22809);
nand U24009 (N_24009,N_22702,N_23473);
nand U24010 (N_24010,N_22971,N_23227);
xnor U24011 (N_24011,N_23239,N_23368);
or U24012 (N_24012,N_23453,N_22628);
nand U24013 (N_24013,N_23353,N_23123);
and U24014 (N_24014,N_22831,N_23735);
and U24015 (N_24015,N_23745,N_23691);
nor U24016 (N_24016,N_22695,N_23002);
xor U24017 (N_24017,N_23420,N_23226);
and U24018 (N_24018,N_22901,N_22719);
or U24019 (N_24019,N_22633,N_22928);
and U24020 (N_24020,N_23722,N_23341);
nand U24021 (N_24021,N_23627,N_23634);
xor U24022 (N_24022,N_23488,N_22853);
nand U24023 (N_24023,N_23148,N_22683);
xnor U24024 (N_24024,N_23672,N_23143);
xor U24025 (N_24025,N_22562,N_23291);
nor U24026 (N_24026,N_22845,N_22659);
xor U24027 (N_24027,N_23156,N_22898);
nand U24028 (N_24028,N_23577,N_22652);
and U24029 (N_24029,N_23702,N_23181);
and U24030 (N_24030,N_23161,N_23475);
nand U24031 (N_24031,N_23000,N_23405);
or U24032 (N_24032,N_23285,N_22706);
and U24033 (N_24033,N_23287,N_23592);
nand U24034 (N_24034,N_22525,N_22575);
or U24035 (N_24035,N_23219,N_23562);
nand U24036 (N_24036,N_23552,N_23370);
nand U24037 (N_24037,N_23431,N_23113);
or U24038 (N_24038,N_22769,N_23236);
or U24039 (N_24039,N_22646,N_23615);
and U24040 (N_24040,N_23526,N_22544);
nor U24041 (N_24041,N_23191,N_23200);
or U24042 (N_24042,N_23089,N_22510);
nand U24043 (N_24043,N_23525,N_23320);
or U24044 (N_24044,N_22839,N_23313);
and U24045 (N_24045,N_23608,N_22854);
nor U24046 (N_24046,N_23354,N_22591);
or U24047 (N_24047,N_23238,N_23616);
nor U24048 (N_24048,N_23046,N_22934);
and U24049 (N_24049,N_22577,N_23580);
nand U24050 (N_24050,N_22692,N_23186);
nor U24051 (N_24051,N_22798,N_22533);
nor U24052 (N_24052,N_22810,N_22872);
nand U24053 (N_24053,N_23421,N_22666);
or U24054 (N_24054,N_23531,N_22918);
xnor U24055 (N_24055,N_23115,N_22505);
nand U24056 (N_24056,N_23309,N_22956);
and U24057 (N_24057,N_23571,N_22697);
or U24058 (N_24058,N_23731,N_23195);
nand U24059 (N_24059,N_22776,N_23584);
or U24060 (N_24060,N_22590,N_23650);
or U24061 (N_24061,N_23520,N_22627);
or U24062 (N_24062,N_23447,N_23399);
nand U24063 (N_24063,N_23378,N_23049);
or U24064 (N_24064,N_23437,N_23619);
nor U24065 (N_24065,N_23317,N_23077);
nand U24066 (N_24066,N_22987,N_23647);
nand U24067 (N_24067,N_23180,N_22651);
nand U24068 (N_24068,N_22828,N_22963);
or U24069 (N_24069,N_23708,N_23091);
and U24070 (N_24070,N_22765,N_23124);
nand U24071 (N_24071,N_22630,N_22997);
and U24072 (N_24072,N_22875,N_22894);
xnor U24073 (N_24073,N_22523,N_23587);
xnor U24074 (N_24074,N_22746,N_23379);
xor U24075 (N_24075,N_23335,N_23371);
or U24076 (N_24076,N_22977,N_22512);
or U24077 (N_24077,N_23255,N_22761);
or U24078 (N_24078,N_23544,N_23237);
nor U24079 (N_24079,N_23631,N_22950);
nand U24080 (N_24080,N_23122,N_22699);
nor U24081 (N_24081,N_23165,N_22799);
or U24082 (N_24082,N_22849,N_23248);
and U24083 (N_24083,N_22874,N_22818);
nor U24084 (N_24084,N_22556,N_23414);
and U24085 (N_24085,N_23251,N_23559);
xor U24086 (N_24086,N_22922,N_22801);
nor U24087 (N_24087,N_23334,N_22902);
nor U24088 (N_24088,N_23052,N_22691);
xor U24089 (N_24089,N_23524,N_23082);
nand U24090 (N_24090,N_23294,N_22773);
nand U24091 (N_24091,N_22673,N_22725);
xnor U24092 (N_24092,N_23667,N_23012);
xor U24093 (N_24093,N_23063,N_23120);
nor U24094 (N_24094,N_23009,N_22927);
nor U24095 (N_24095,N_22656,N_22966);
and U24096 (N_24096,N_22755,N_22882);
and U24097 (N_24097,N_23741,N_22949);
or U24098 (N_24098,N_23482,N_23310);
nor U24099 (N_24099,N_23322,N_22638);
nor U24100 (N_24100,N_23734,N_22844);
nor U24101 (N_24101,N_23700,N_22870);
or U24102 (N_24102,N_23432,N_22567);
and U24103 (N_24103,N_23716,N_22543);
xor U24104 (N_24104,N_23469,N_23459);
nand U24105 (N_24105,N_22786,N_22887);
or U24106 (N_24106,N_22609,N_22848);
and U24107 (N_24107,N_23192,N_23522);
and U24108 (N_24108,N_22863,N_23262);
nor U24109 (N_24109,N_23706,N_23048);
and U24110 (N_24110,N_23027,N_23356);
nor U24111 (N_24111,N_23190,N_23302);
nor U24112 (N_24112,N_23015,N_23167);
or U24113 (N_24113,N_23033,N_23295);
xor U24114 (N_24114,N_23241,N_23683);
nand U24115 (N_24115,N_23376,N_22832);
nand U24116 (N_24116,N_22888,N_23480);
nor U24117 (N_24117,N_23270,N_23662);
xnor U24118 (N_24118,N_22789,N_22632);
nand U24119 (N_24119,N_23463,N_22802);
or U24120 (N_24120,N_23085,N_22714);
xor U24121 (N_24121,N_23671,N_22514);
xor U24122 (N_24122,N_23360,N_23234);
or U24123 (N_24123,N_22783,N_22621);
or U24124 (N_24124,N_23507,N_23117);
nor U24125 (N_24125,N_23635,N_23563);
xor U24126 (N_24126,N_23235,N_23675);
or U24127 (N_24127,N_23006,N_22771);
and U24128 (N_24128,N_23175,N_22745);
nor U24129 (N_24129,N_22678,N_23685);
nand U24130 (N_24130,N_22620,N_22919);
or U24131 (N_24131,N_23208,N_22527);
and U24132 (N_24132,N_23166,N_22942);
xnor U24133 (N_24133,N_22920,N_22641);
nor U24134 (N_24134,N_23481,N_23035);
or U24135 (N_24135,N_22897,N_23017);
nand U24136 (N_24136,N_23350,N_22797);
xor U24137 (N_24137,N_23712,N_22806);
and U24138 (N_24138,N_23581,N_23495);
xor U24139 (N_24139,N_23535,N_22896);
xor U24140 (N_24140,N_23288,N_23080);
nor U24141 (N_24141,N_22708,N_22985);
nand U24142 (N_24142,N_22688,N_23384);
xor U24143 (N_24143,N_23640,N_23064);
or U24144 (N_24144,N_22829,N_23256);
or U24145 (N_24145,N_23108,N_23664);
and U24146 (N_24146,N_22914,N_22857);
nor U24147 (N_24147,N_22707,N_22681);
xor U24148 (N_24148,N_22911,N_23374);
xnor U24149 (N_24149,N_22916,N_23680);
nor U24150 (N_24150,N_23311,N_23267);
and U24151 (N_24151,N_23467,N_23477);
nor U24152 (N_24152,N_22993,N_23189);
xor U24153 (N_24153,N_23114,N_23390);
nand U24154 (N_24154,N_23144,N_22906);
and U24155 (N_24155,N_23177,N_22805);
and U24156 (N_24156,N_23660,N_23164);
xor U24157 (N_24157,N_23184,N_23611);
and U24158 (N_24158,N_23512,N_23315);
and U24159 (N_24159,N_22883,N_22507);
and U24160 (N_24160,N_23283,N_22800);
nand U24161 (N_24161,N_23304,N_23365);
nand U24162 (N_24162,N_22941,N_22616);
nand U24163 (N_24163,N_23107,N_23045);
nand U24164 (N_24164,N_22787,N_22838);
nand U24165 (N_24165,N_22675,N_23649);
nand U24166 (N_24166,N_22586,N_22576);
or U24167 (N_24167,N_22640,N_22758);
or U24168 (N_24168,N_23338,N_22526);
nand U24169 (N_24169,N_23303,N_22965);
nor U24170 (N_24170,N_23053,N_22738);
or U24171 (N_24171,N_22836,N_22864);
or U24172 (N_24172,N_23361,N_22547);
nand U24173 (N_24173,N_22937,N_22878);
and U24174 (N_24174,N_23042,N_23363);
xnor U24175 (N_24175,N_22959,N_22900);
or U24176 (N_24176,N_22570,N_23500);
xnor U24177 (N_24177,N_22972,N_23417);
nor U24178 (N_24178,N_23538,N_22614);
xor U24179 (N_24179,N_23561,N_22766);
nand U24180 (N_24180,N_23610,N_23707);
nand U24181 (N_24181,N_22884,N_23205);
and U24182 (N_24182,N_23273,N_23464);
xor U24183 (N_24183,N_23062,N_23260);
xor U24184 (N_24184,N_23569,N_23018);
nand U24185 (N_24185,N_23151,N_22561);
nand U24186 (N_24186,N_22899,N_22969);
nand U24187 (N_24187,N_23253,N_23276);
nor U24188 (N_24188,N_23188,N_23160);
nor U24189 (N_24189,N_22555,N_23125);
and U24190 (N_24190,N_23289,N_22886);
or U24191 (N_24191,N_22791,N_23424);
nor U24192 (N_24192,N_22615,N_23714);
and U24193 (N_24193,N_23223,N_23407);
xnor U24194 (N_24194,N_23673,N_23153);
nand U24195 (N_24195,N_23728,N_23024);
nor U24196 (N_24196,N_23652,N_23614);
and U24197 (N_24197,N_23264,N_23196);
nand U24198 (N_24198,N_23697,N_23415);
nand U24199 (N_24199,N_23653,N_22938);
nor U24200 (N_24200,N_23529,N_22531);
or U24201 (N_24201,N_23503,N_22860);
or U24202 (N_24202,N_23483,N_23579);
nor U24203 (N_24203,N_23296,N_22530);
xnor U24204 (N_24204,N_22764,N_23620);
nand U24205 (N_24205,N_23100,N_23249);
nand U24206 (N_24206,N_23187,N_23290);
and U24207 (N_24207,N_22890,N_22566);
xor U24208 (N_24208,N_23326,N_23511);
or U24209 (N_24209,N_23491,N_22930);
and U24210 (N_24210,N_22710,N_23690);
and U24211 (N_24211,N_23106,N_22943);
and U24212 (N_24212,N_23170,N_23268);
xnor U24213 (N_24213,N_22642,N_23055);
and U24214 (N_24214,N_23171,N_22951);
xor U24215 (N_24215,N_22905,N_23568);
nand U24216 (N_24216,N_23674,N_22991);
and U24217 (N_24217,N_23623,N_22548);
xor U24218 (N_24218,N_22572,N_23329);
nor U24219 (N_24219,N_23199,N_22595);
and U24220 (N_24220,N_23699,N_22677);
nor U24221 (N_24221,N_23259,N_23131);
xor U24222 (N_24222,N_23194,N_23474);
and U24223 (N_24223,N_22804,N_23110);
and U24224 (N_24224,N_23135,N_23298);
xor U24225 (N_24225,N_22856,N_23703);
or U24226 (N_24226,N_23441,N_22611);
nand U24227 (N_24227,N_23628,N_23468);
nor U24228 (N_24228,N_23383,N_23597);
and U24229 (N_24229,N_23163,N_22644);
xor U24230 (N_24230,N_22729,N_22668);
xor U24231 (N_24231,N_23665,N_23537);
nor U24232 (N_24232,N_22698,N_23515);
and U24233 (N_24233,N_23074,N_22774);
nand U24234 (N_24234,N_23071,N_23201);
nand U24235 (N_24235,N_22778,N_23008);
xor U24236 (N_24236,N_23266,N_22925);
or U24237 (N_24237,N_23717,N_22503);
nor U24238 (N_24238,N_23746,N_22606);
or U24239 (N_24239,N_22720,N_22601);
nand U24240 (N_24240,N_22517,N_22661);
or U24241 (N_24241,N_23740,N_23277);
nand U24242 (N_24242,N_23400,N_23228);
nand U24243 (N_24243,N_22847,N_23566);
nand U24244 (N_24244,N_23419,N_23436);
nor U24245 (N_24245,N_23484,N_23272);
and U24246 (N_24246,N_22814,N_22803);
and U24247 (N_24247,N_23305,N_22726);
nor U24248 (N_24248,N_22790,N_23319);
and U24249 (N_24249,N_22948,N_22953);
nor U24250 (N_24250,N_23032,N_23725);
nand U24251 (N_24251,N_23138,N_23097);
nand U24252 (N_24252,N_22760,N_22602);
xor U24253 (N_24253,N_23358,N_22756);
or U24254 (N_24254,N_23410,N_22909);
xor U24255 (N_24255,N_22740,N_23224);
or U24256 (N_24256,N_23517,N_23142);
nor U24257 (N_24257,N_23325,N_22825);
xor U24258 (N_24258,N_22757,N_23179);
xnor U24259 (N_24259,N_23721,N_23648);
nand U24260 (N_24260,N_23214,N_23661);
and U24261 (N_24261,N_23387,N_22715);
and U24262 (N_24262,N_23403,N_23328);
nor U24263 (N_24263,N_23547,N_23121);
nand U24264 (N_24264,N_22961,N_23626);
nand U24265 (N_24265,N_23389,N_23681);
nor U24266 (N_24266,N_22722,N_22749);
xnor U24267 (N_24267,N_22780,N_22536);
nand U24268 (N_24268,N_22564,N_23397);
nor U24269 (N_24269,N_23037,N_22686);
xnor U24270 (N_24270,N_23496,N_23534);
and U24271 (N_24271,N_22520,N_23286);
nand U24272 (N_24272,N_22752,N_23402);
or U24273 (N_24273,N_23553,N_22604);
nand U24274 (N_24274,N_23532,N_23067);
nor U24275 (N_24275,N_22553,N_23297);
or U24276 (N_24276,N_22545,N_23711);
and U24277 (N_24277,N_23550,N_23586);
and U24278 (N_24278,N_22687,N_22669);
xor U24279 (N_24279,N_22830,N_23573);
nand U24280 (N_24280,N_22973,N_23168);
nor U24281 (N_24281,N_22880,N_22664);
and U24282 (N_24282,N_22835,N_22762);
nor U24283 (N_24283,N_22808,N_23622);
nor U24284 (N_24284,N_22772,N_23705);
xor U24285 (N_24285,N_22970,N_23543);
or U24286 (N_24286,N_23478,N_22712);
nor U24287 (N_24287,N_22732,N_23362);
xor U24288 (N_24288,N_22777,N_23182);
nand U24289 (N_24289,N_23668,N_23663);
nor U24290 (N_24290,N_23446,N_23169);
nor U24291 (N_24291,N_22711,N_22625);
xnor U24292 (N_24292,N_23292,N_23150);
or U24293 (N_24293,N_23075,N_22502);
xor U24294 (N_24294,N_23498,N_22974);
nor U24295 (N_24295,N_22679,N_23364);
or U24296 (N_24296,N_22703,N_23207);
xnor U24297 (N_24297,N_23072,N_22823);
and U24298 (N_24298,N_23530,N_23282);
xnor U24299 (N_24299,N_23744,N_22980);
or U24300 (N_24300,N_23704,N_23501);
xnor U24301 (N_24301,N_23452,N_23733);
nor U24302 (N_24302,N_22582,N_23718);
nand U24303 (N_24303,N_23430,N_23173);
or U24304 (N_24304,N_23247,N_23158);
and U24305 (N_24305,N_23618,N_23567);
and U24306 (N_24306,N_23748,N_23409);
and U24307 (N_24307,N_22532,N_22696);
nand U24308 (N_24308,N_22535,N_23719);
nor U24309 (N_24309,N_23141,N_23451);
xnor U24310 (N_24310,N_23605,N_23382);
xor U24311 (N_24311,N_23079,N_23222);
nand U24312 (N_24312,N_22751,N_22623);
nor U24313 (N_24313,N_23105,N_23278);
nand U24314 (N_24314,N_22541,N_22779);
or U24315 (N_24315,N_23104,N_22608);
xnor U24316 (N_24316,N_23572,N_22565);
nor U24317 (N_24317,N_23425,N_22552);
or U24318 (N_24318,N_23047,N_23034);
or U24319 (N_24319,N_23645,N_23229);
xnor U24320 (N_24320,N_22770,N_22743);
and U24321 (N_24321,N_22705,N_22723);
xnor U24322 (N_24322,N_22600,N_23539);
nand U24323 (N_24323,N_23458,N_23174);
xnor U24324 (N_24324,N_22954,N_22624);
xnor U24325 (N_24325,N_23565,N_22837);
xor U24326 (N_24326,N_23221,N_23116);
or U24327 (N_24327,N_23204,N_23185);
or U24328 (N_24328,N_23737,N_22792);
or U24329 (N_24329,N_23068,N_23506);
nand U24330 (N_24330,N_23589,N_22939);
nor U24331 (N_24331,N_23659,N_22573);
xnor U24332 (N_24332,N_23670,N_22767);
nor U24333 (N_24333,N_23448,N_23061);
nor U24334 (N_24334,N_23001,N_22540);
nand U24335 (N_24335,N_23019,N_22568);
or U24336 (N_24336,N_23007,N_23641);
nand U24337 (N_24337,N_23710,N_22846);
or U24338 (N_24338,N_22581,N_23598);
nor U24339 (N_24339,N_23028,N_23099);
nand U24340 (N_24340,N_22504,N_22785);
or U24341 (N_24341,N_22667,N_22873);
and U24342 (N_24342,N_22597,N_22571);
xnor U24343 (N_24343,N_23564,N_22588);
xnor U24344 (N_24344,N_23602,N_22718);
or U24345 (N_24345,N_23380,N_23275);
nor U24346 (N_24346,N_23505,N_23590);
nand U24347 (N_24347,N_22539,N_23693);
and U24348 (N_24348,N_22861,N_22574);
nor U24349 (N_24349,N_22506,N_22682);
nand U24350 (N_24350,N_23359,N_23381);
xnor U24351 (N_24351,N_23130,N_23377);
nand U24352 (N_24352,N_23576,N_23367);
xor U24353 (N_24353,N_22554,N_22716);
nor U24354 (N_24354,N_23218,N_23145);
nor U24355 (N_24355,N_23687,N_23059);
or U24356 (N_24356,N_23457,N_22509);
nand U24357 (N_24357,N_22636,N_23345);
nor U24358 (N_24358,N_23551,N_23438);
or U24359 (N_24359,N_22672,N_23715);
nor U24360 (N_24360,N_23742,N_23005);
nor U24361 (N_24361,N_22731,N_23318);
or U24362 (N_24362,N_23465,N_22655);
nand U24363 (N_24363,N_23462,N_23355);
nor U24364 (N_24364,N_23528,N_23172);
and U24365 (N_24365,N_22981,N_23340);
nand U24366 (N_24366,N_23609,N_22795);
and U24367 (N_24367,N_23471,N_23119);
xor U24368 (N_24368,N_23466,N_22500);
xor U24369 (N_24369,N_23271,N_23126);
xnor U24370 (N_24370,N_23279,N_23450);
nand U24371 (N_24371,N_22733,N_23257);
nor U24372 (N_24372,N_22782,N_22781);
and U24373 (N_24373,N_23596,N_23406);
nand U24374 (N_24374,N_22820,N_22522);
xor U24375 (N_24375,N_22868,N_22759);
nand U24376 (N_24376,N_22826,N_23203);
xnor U24377 (N_24377,N_23676,N_23182);
nand U24378 (N_24378,N_23393,N_22702);
xor U24379 (N_24379,N_23432,N_23430);
or U24380 (N_24380,N_22864,N_23138);
nand U24381 (N_24381,N_22931,N_22713);
or U24382 (N_24382,N_23506,N_23043);
nor U24383 (N_24383,N_22614,N_23263);
nand U24384 (N_24384,N_23281,N_23284);
xnor U24385 (N_24385,N_23034,N_23465);
nand U24386 (N_24386,N_23685,N_22721);
xor U24387 (N_24387,N_23260,N_23142);
xor U24388 (N_24388,N_22989,N_23499);
nor U24389 (N_24389,N_23285,N_23315);
and U24390 (N_24390,N_23633,N_23024);
or U24391 (N_24391,N_22916,N_23480);
nand U24392 (N_24392,N_23284,N_22606);
xor U24393 (N_24393,N_23741,N_23133);
or U24394 (N_24394,N_22744,N_23454);
xnor U24395 (N_24395,N_23561,N_22875);
nand U24396 (N_24396,N_22905,N_23099);
nand U24397 (N_24397,N_22748,N_22761);
or U24398 (N_24398,N_23444,N_23602);
and U24399 (N_24399,N_23355,N_22503);
nor U24400 (N_24400,N_23655,N_23117);
nor U24401 (N_24401,N_23584,N_22737);
xor U24402 (N_24402,N_23233,N_22797);
nand U24403 (N_24403,N_23724,N_22581);
nor U24404 (N_24404,N_22893,N_23016);
or U24405 (N_24405,N_23566,N_23049);
nor U24406 (N_24406,N_23269,N_22705);
xor U24407 (N_24407,N_23688,N_23100);
or U24408 (N_24408,N_23134,N_23383);
nand U24409 (N_24409,N_22908,N_22728);
and U24410 (N_24410,N_22988,N_23032);
xnor U24411 (N_24411,N_23092,N_22636);
nor U24412 (N_24412,N_22975,N_22870);
nor U24413 (N_24413,N_23131,N_23130);
xnor U24414 (N_24414,N_23286,N_22697);
or U24415 (N_24415,N_23733,N_23453);
or U24416 (N_24416,N_23233,N_23538);
xor U24417 (N_24417,N_23307,N_23009);
xor U24418 (N_24418,N_23129,N_23538);
and U24419 (N_24419,N_22996,N_23358);
nor U24420 (N_24420,N_22968,N_23097);
and U24421 (N_24421,N_23384,N_22881);
and U24422 (N_24422,N_23298,N_23695);
nand U24423 (N_24423,N_23697,N_22799);
nor U24424 (N_24424,N_23617,N_23283);
nand U24425 (N_24425,N_23643,N_23097);
or U24426 (N_24426,N_22532,N_22541);
nor U24427 (N_24427,N_22835,N_23740);
or U24428 (N_24428,N_22981,N_22703);
xor U24429 (N_24429,N_22578,N_23309);
nand U24430 (N_24430,N_23281,N_23327);
xnor U24431 (N_24431,N_22582,N_22811);
nand U24432 (N_24432,N_23594,N_23512);
and U24433 (N_24433,N_22650,N_23358);
nand U24434 (N_24434,N_23691,N_23015);
nor U24435 (N_24435,N_23415,N_23735);
or U24436 (N_24436,N_23493,N_23703);
or U24437 (N_24437,N_23477,N_23236);
xnor U24438 (N_24438,N_22788,N_22951);
or U24439 (N_24439,N_22584,N_23144);
nand U24440 (N_24440,N_22665,N_23681);
nor U24441 (N_24441,N_23223,N_23074);
or U24442 (N_24442,N_23130,N_23266);
nand U24443 (N_24443,N_22853,N_22790);
xor U24444 (N_24444,N_23435,N_23407);
nand U24445 (N_24445,N_23643,N_23333);
xor U24446 (N_24446,N_23478,N_23109);
xor U24447 (N_24447,N_23724,N_22626);
and U24448 (N_24448,N_22947,N_22910);
or U24449 (N_24449,N_23692,N_23432);
and U24450 (N_24450,N_23136,N_22974);
xor U24451 (N_24451,N_23053,N_23199);
xor U24452 (N_24452,N_22853,N_22906);
or U24453 (N_24453,N_22641,N_22735);
nand U24454 (N_24454,N_22739,N_23396);
xor U24455 (N_24455,N_23591,N_23128);
nand U24456 (N_24456,N_22640,N_23498);
nor U24457 (N_24457,N_23157,N_23278);
xor U24458 (N_24458,N_23545,N_23338);
xor U24459 (N_24459,N_22968,N_22882);
nor U24460 (N_24460,N_22673,N_23610);
and U24461 (N_24461,N_22835,N_22737);
nor U24462 (N_24462,N_22840,N_22985);
nor U24463 (N_24463,N_23459,N_23095);
xor U24464 (N_24464,N_22854,N_22795);
nand U24465 (N_24465,N_23458,N_22609);
nor U24466 (N_24466,N_23533,N_23157);
nor U24467 (N_24467,N_23410,N_22901);
nor U24468 (N_24468,N_22555,N_22508);
nor U24469 (N_24469,N_23062,N_23248);
nor U24470 (N_24470,N_22646,N_23308);
or U24471 (N_24471,N_23283,N_23336);
or U24472 (N_24472,N_23138,N_22733);
or U24473 (N_24473,N_23588,N_22835);
and U24474 (N_24474,N_23108,N_23404);
nand U24475 (N_24475,N_22964,N_22528);
or U24476 (N_24476,N_23738,N_22579);
nand U24477 (N_24477,N_23350,N_23065);
and U24478 (N_24478,N_23742,N_23430);
or U24479 (N_24479,N_22760,N_23125);
nor U24480 (N_24480,N_23397,N_23699);
nor U24481 (N_24481,N_23526,N_22784);
nor U24482 (N_24482,N_23150,N_22749);
and U24483 (N_24483,N_23304,N_23427);
or U24484 (N_24484,N_23630,N_23370);
xnor U24485 (N_24485,N_23199,N_23040);
and U24486 (N_24486,N_22939,N_22729);
nand U24487 (N_24487,N_22566,N_23318);
nand U24488 (N_24488,N_23215,N_22737);
xnor U24489 (N_24489,N_23441,N_22620);
nand U24490 (N_24490,N_23443,N_23006);
nand U24491 (N_24491,N_22544,N_22579);
and U24492 (N_24492,N_23498,N_23636);
or U24493 (N_24493,N_23596,N_22902);
nor U24494 (N_24494,N_23562,N_23477);
or U24495 (N_24495,N_23139,N_22500);
and U24496 (N_24496,N_22764,N_23699);
or U24497 (N_24497,N_22526,N_22894);
xnor U24498 (N_24498,N_23046,N_23630);
and U24499 (N_24499,N_22608,N_22566);
nor U24500 (N_24500,N_22558,N_22770);
nor U24501 (N_24501,N_23011,N_23216);
or U24502 (N_24502,N_22877,N_22610);
xor U24503 (N_24503,N_23530,N_22727);
and U24504 (N_24504,N_23658,N_22966);
nor U24505 (N_24505,N_23104,N_23450);
nand U24506 (N_24506,N_22992,N_23097);
xnor U24507 (N_24507,N_22836,N_23245);
or U24508 (N_24508,N_23224,N_22618);
xnor U24509 (N_24509,N_23630,N_22664);
nor U24510 (N_24510,N_23183,N_23564);
xor U24511 (N_24511,N_23058,N_22810);
xnor U24512 (N_24512,N_22622,N_23641);
or U24513 (N_24513,N_23422,N_23089);
nand U24514 (N_24514,N_23217,N_23198);
nor U24515 (N_24515,N_23260,N_23717);
nand U24516 (N_24516,N_22568,N_22958);
nand U24517 (N_24517,N_22891,N_23131);
and U24518 (N_24518,N_23182,N_22789);
and U24519 (N_24519,N_22767,N_23569);
xnor U24520 (N_24520,N_23399,N_22945);
and U24521 (N_24521,N_23152,N_23562);
nor U24522 (N_24522,N_23637,N_23716);
and U24523 (N_24523,N_23415,N_23355);
nor U24524 (N_24524,N_22627,N_22779);
nand U24525 (N_24525,N_23054,N_23015);
and U24526 (N_24526,N_23696,N_22685);
nor U24527 (N_24527,N_22766,N_22826);
nand U24528 (N_24528,N_23056,N_23519);
and U24529 (N_24529,N_22689,N_23291);
or U24530 (N_24530,N_23493,N_22833);
nand U24531 (N_24531,N_23586,N_22962);
xor U24532 (N_24532,N_22795,N_23564);
nand U24533 (N_24533,N_23710,N_22755);
nor U24534 (N_24534,N_22624,N_22694);
nor U24535 (N_24535,N_22782,N_23134);
xnor U24536 (N_24536,N_23252,N_22622);
and U24537 (N_24537,N_23052,N_22705);
nand U24538 (N_24538,N_22541,N_22727);
xor U24539 (N_24539,N_23547,N_23175);
or U24540 (N_24540,N_22778,N_22570);
nor U24541 (N_24541,N_23234,N_23357);
nor U24542 (N_24542,N_23116,N_23264);
and U24543 (N_24543,N_22675,N_22992);
and U24544 (N_24544,N_22818,N_23330);
xnor U24545 (N_24545,N_22724,N_22827);
xor U24546 (N_24546,N_23308,N_23096);
or U24547 (N_24547,N_23236,N_23638);
and U24548 (N_24548,N_22754,N_23420);
nand U24549 (N_24549,N_22847,N_22729);
or U24550 (N_24550,N_23038,N_22576);
nor U24551 (N_24551,N_23178,N_22911);
and U24552 (N_24552,N_23618,N_23739);
or U24553 (N_24553,N_23210,N_23683);
nand U24554 (N_24554,N_22503,N_23364);
xnor U24555 (N_24555,N_23605,N_23421);
nor U24556 (N_24556,N_23168,N_23217);
and U24557 (N_24557,N_23640,N_22735);
and U24558 (N_24558,N_22637,N_23388);
and U24559 (N_24559,N_22601,N_22838);
nor U24560 (N_24560,N_23151,N_23101);
or U24561 (N_24561,N_23131,N_23625);
xnor U24562 (N_24562,N_22999,N_22946);
or U24563 (N_24563,N_22588,N_22611);
xnor U24564 (N_24564,N_23253,N_23731);
and U24565 (N_24565,N_23387,N_22871);
and U24566 (N_24566,N_22751,N_22996);
nand U24567 (N_24567,N_23346,N_23322);
xor U24568 (N_24568,N_23114,N_23299);
nand U24569 (N_24569,N_22666,N_22841);
nand U24570 (N_24570,N_23604,N_23664);
and U24571 (N_24571,N_22819,N_23007);
or U24572 (N_24572,N_23249,N_23213);
nand U24573 (N_24573,N_23047,N_22643);
or U24574 (N_24574,N_22647,N_22501);
and U24575 (N_24575,N_22671,N_23154);
nand U24576 (N_24576,N_22522,N_23005);
nor U24577 (N_24577,N_22833,N_23681);
xnor U24578 (N_24578,N_23517,N_22958);
nand U24579 (N_24579,N_22710,N_23223);
or U24580 (N_24580,N_23704,N_22879);
xnor U24581 (N_24581,N_23084,N_22556);
or U24582 (N_24582,N_23626,N_23225);
xnor U24583 (N_24583,N_23558,N_22570);
and U24584 (N_24584,N_22882,N_23202);
nor U24585 (N_24585,N_22794,N_22798);
or U24586 (N_24586,N_23184,N_23330);
nand U24587 (N_24587,N_22522,N_22798);
nand U24588 (N_24588,N_23683,N_22518);
nor U24589 (N_24589,N_23647,N_23109);
and U24590 (N_24590,N_22619,N_22935);
or U24591 (N_24591,N_23264,N_22568);
xor U24592 (N_24592,N_23054,N_22967);
nand U24593 (N_24593,N_23401,N_23559);
nand U24594 (N_24594,N_23184,N_23364);
nor U24595 (N_24595,N_22659,N_23600);
nand U24596 (N_24596,N_22559,N_23489);
xnor U24597 (N_24597,N_23469,N_23184);
and U24598 (N_24598,N_23127,N_23591);
and U24599 (N_24599,N_23139,N_22842);
and U24600 (N_24600,N_23180,N_22896);
nor U24601 (N_24601,N_22524,N_22721);
nand U24602 (N_24602,N_22945,N_22957);
nand U24603 (N_24603,N_23522,N_22656);
nand U24604 (N_24604,N_22608,N_22790);
nor U24605 (N_24605,N_23506,N_23265);
and U24606 (N_24606,N_23660,N_23077);
xnor U24607 (N_24607,N_22670,N_23446);
nor U24608 (N_24608,N_23092,N_22875);
and U24609 (N_24609,N_23144,N_23149);
or U24610 (N_24610,N_23485,N_23299);
or U24611 (N_24611,N_22550,N_23626);
and U24612 (N_24612,N_23246,N_22567);
or U24613 (N_24613,N_22628,N_23700);
or U24614 (N_24614,N_23597,N_22684);
nor U24615 (N_24615,N_23520,N_23677);
nor U24616 (N_24616,N_23154,N_23126);
nor U24617 (N_24617,N_23310,N_23712);
and U24618 (N_24618,N_23735,N_22818);
or U24619 (N_24619,N_23302,N_23076);
and U24620 (N_24620,N_22952,N_22592);
nand U24621 (N_24621,N_22528,N_23359);
xor U24622 (N_24622,N_22803,N_23734);
xor U24623 (N_24623,N_22883,N_22654);
or U24624 (N_24624,N_23643,N_22970);
nor U24625 (N_24625,N_23348,N_22957);
xnor U24626 (N_24626,N_23447,N_23466);
xnor U24627 (N_24627,N_22651,N_23635);
nand U24628 (N_24628,N_23029,N_22788);
xnor U24629 (N_24629,N_22672,N_22662);
or U24630 (N_24630,N_23735,N_23343);
xor U24631 (N_24631,N_23638,N_22831);
nand U24632 (N_24632,N_23199,N_23749);
or U24633 (N_24633,N_22907,N_23204);
nand U24634 (N_24634,N_23158,N_22759);
and U24635 (N_24635,N_22578,N_23117);
xor U24636 (N_24636,N_23512,N_23327);
xor U24637 (N_24637,N_22689,N_22907);
or U24638 (N_24638,N_23648,N_23494);
xor U24639 (N_24639,N_22873,N_22682);
nor U24640 (N_24640,N_22992,N_23174);
and U24641 (N_24641,N_23286,N_23229);
nor U24642 (N_24642,N_23149,N_22747);
nor U24643 (N_24643,N_23547,N_23491);
nor U24644 (N_24644,N_23184,N_23051);
xnor U24645 (N_24645,N_22710,N_22672);
or U24646 (N_24646,N_23381,N_23319);
and U24647 (N_24647,N_23255,N_23260);
or U24648 (N_24648,N_22942,N_22643);
or U24649 (N_24649,N_23666,N_23634);
nand U24650 (N_24650,N_22879,N_23085);
or U24651 (N_24651,N_22774,N_22661);
xnor U24652 (N_24652,N_22732,N_22619);
or U24653 (N_24653,N_23685,N_22569);
nor U24654 (N_24654,N_23500,N_22569);
nor U24655 (N_24655,N_22928,N_23054);
xnor U24656 (N_24656,N_23520,N_23740);
xnor U24657 (N_24657,N_22685,N_23403);
xnor U24658 (N_24658,N_23498,N_23301);
nor U24659 (N_24659,N_22965,N_22761);
nor U24660 (N_24660,N_23466,N_23535);
or U24661 (N_24661,N_23235,N_22652);
and U24662 (N_24662,N_23193,N_23473);
and U24663 (N_24663,N_22852,N_23216);
or U24664 (N_24664,N_23532,N_22913);
xor U24665 (N_24665,N_23133,N_22722);
nor U24666 (N_24666,N_23374,N_23113);
xnor U24667 (N_24667,N_22799,N_22652);
nor U24668 (N_24668,N_23496,N_23714);
nor U24669 (N_24669,N_22500,N_23000);
or U24670 (N_24670,N_23524,N_23275);
xor U24671 (N_24671,N_23683,N_22800);
nand U24672 (N_24672,N_22762,N_23247);
xor U24673 (N_24673,N_23627,N_22682);
nor U24674 (N_24674,N_23569,N_22736);
xor U24675 (N_24675,N_23629,N_23633);
xnor U24676 (N_24676,N_23713,N_22843);
and U24677 (N_24677,N_23358,N_23142);
or U24678 (N_24678,N_23093,N_23006);
xor U24679 (N_24679,N_23573,N_22672);
xnor U24680 (N_24680,N_22526,N_22778);
nand U24681 (N_24681,N_23589,N_22733);
or U24682 (N_24682,N_23531,N_22597);
nand U24683 (N_24683,N_23562,N_23424);
nand U24684 (N_24684,N_22521,N_22893);
and U24685 (N_24685,N_22551,N_22722);
xor U24686 (N_24686,N_23269,N_23649);
or U24687 (N_24687,N_23488,N_22971);
nor U24688 (N_24688,N_23101,N_22853);
nand U24689 (N_24689,N_23081,N_23247);
nor U24690 (N_24690,N_22771,N_23011);
xor U24691 (N_24691,N_22504,N_23406);
or U24692 (N_24692,N_23602,N_22623);
xnor U24693 (N_24693,N_22695,N_23376);
nor U24694 (N_24694,N_23129,N_22661);
and U24695 (N_24695,N_23188,N_22745);
or U24696 (N_24696,N_22934,N_23390);
nor U24697 (N_24697,N_22593,N_23279);
nand U24698 (N_24698,N_22697,N_23143);
and U24699 (N_24699,N_23678,N_23615);
or U24700 (N_24700,N_22949,N_23141);
or U24701 (N_24701,N_23377,N_23127);
and U24702 (N_24702,N_22502,N_22996);
or U24703 (N_24703,N_23347,N_22879);
or U24704 (N_24704,N_22837,N_23430);
and U24705 (N_24705,N_23115,N_23603);
nand U24706 (N_24706,N_23238,N_23376);
nor U24707 (N_24707,N_23587,N_23298);
nand U24708 (N_24708,N_23547,N_23576);
or U24709 (N_24709,N_22595,N_22864);
and U24710 (N_24710,N_23740,N_22752);
xor U24711 (N_24711,N_23345,N_23488);
xnor U24712 (N_24712,N_22825,N_22732);
and U24713 (N_24713,N_22724,N_22564);
nor U24714 (N_24714,N_22942,N_22840);
nor U24715 (N_24715,N_22635,N_23588);
nor U24716 (N_24716,N_22519,N_23414);
nand U24717 (N_24717,N_23122,N_23490);
nand U24718 (N_24718,N_23652,N_22610);
and U24719 (N_24719,N_23301,N_22862);
or U24720 (N_24720,N_22587,N_22651);
and U24721 (N_24721,N_22808,N_22504);
nor U24722 (N_24722,N_23428,N_23119);
xor U24723 (N_24723,N_23727,N_22865);
and U24724 (N_24724,N_22957,N_23334);
or U24725 (N_24725,N_23097,N_23453);
xnor U24726 (N_24726,N_22650,N_23255);
nand U24727 (N_24727,N_23301,N_22715);
and U24728 (N_24728,N_23562,N_23733);
nor U24729 (N_24729,N_23207,N_23713);
nor U24730 (N_24730,N_22981,N_23461);
nand U24731 (N_24731,N_22727,N_23553);
and U24732 (N_24732,N_22747,N_23067);
and U24733 (N_24733,N_23421,N_23212);
and U24734 (N_24734,N_23682,N_23671);
nor U24735 (N_24735,N_23583,N_23632);
or U24736 (N_24736,N_22974,N_22774);
nor U24737 (N_24737,N_23463,N_22591);
nand U24738 (N_24738,N_22695,N_23109);
and U24739 (N_24739,N_23585,N_23444);
nor U24740 (N_24740,N_22519,N_22910);
xor U24741 (N_24741,N_23645,N_23169);
xor U24742 (N_24742,N_23636,N_23083);
or U24743 (N_24743,N_23206,N_23056);
and U24744 (N_24744,N_23184,N_22815);
nand U24745 (N_24745,N_23398,N_23415);
xor U24746 (N_24746,N_22711,N_23152);
or U24747 (N_24747,N_22543,N_23070);
nor U24748 (N_24748,N_23744,N_23461);
xor U24749 (N_24749,N_22714,N_22571);
and U24750 (N_24750,N_22701,N_22502);
nand U24751 (N_24751,N_23344,N_22936);
and U24752 (N_24752,N_23150,N_23644);
xnor U24753 (N_24753,N_22541,N_23100);
and U24754 (N_24754,N_23401,N_22535);
nand U24755 (N_24755,N_22586,N_22831);
xnor U24756 (N_24756,N_22796,N_22623);
xor U24757 (N_24757,N_23168,N_23581);
or U24758 (N_24758,N_22697,N_22986);
nand U24759 (N_24759,N_23733,N_23339);
and U24760 (N_24760,N_22673,N_23228);
nor U24761 (N_24761,N_22607,N_23534);
xnor U24762 (N_24762,N_22803,N_23330);
or U24763 (N_24763,N_22553,N_22697);
xor U24764 (N_24764,N_23011,N_22933);
and U24765 (N_24765,N_22778,N_23050);
and U24766 (N_24766,N_23330,N_23247);
xnor U24767 (N_24767,N_23183,N_23518);
nor U24768 (N_24768,N_23707,N_22956);
or U24769 (N_24769,N_22787,N_22565);
and U24770 (N_24770,N_22702,N_23428);
nor U24771 (N_24771,N_23693,N_23318);
xor U24772 (N_24772,N_22950,N_23481);
nand U24773 (N_24773,N_22629,N_23658);
xnor U24774 (N_24774,N_23341,N_22747);
nand U24775 (N_24775,N_23448,N_23229);
nor U24776 (N_24776,N_23116,N_23222);
and U24777 (N_24777,N_23062,N_23551);
or U24778 (N_24778,N_23619,N_22686);
or U24779 (N_24779,N_23270,N_22576);
or U24780 (N_24780,N_23575,N_22977);
and U24781 (N_24781,N_23550,N_23144);
or U24782 (N_24782,N_23479,N_23159);
xor U24783 (N_24783,N_23206,N_23654);
and U24784 (N_24784,N_23422,N_23080);
or U24785 (N_24785,N_23518,N_23745);
xnor U24786 (N_24786,N_22904,N_22757);
or U24787 (N_24787,N_22592,N_22955);
xnor U24788 (N_24788,N_22808,N_22952);
or U24789 (N_24789,N_22635,N_23645);
or U24790 (N_24790,N_23624,N_23499);
and U24791 (N_24791,N_22705,N_23110);
or U24792 (N_24792,N_23713,N_22659);
or U24793 (N_24793,N_22845,N_23328);
nand U24794 (N_24794,N_22959,N_22752);
nand U24795 (N_24795,N_23056,N_22921);
nor U24796 (N_24796,N_22663,N_23150);
nor U24797 (N_24797,N_23021,N_23385);
or U24798 (N_24798,N_22511,N_22975);
and U24799 (N_24799,N_23464,N_22915);
and U24800 (N_24800,N_22834,N_23172);
nor U24801 (N_24801,N_23665,N_22809);
or U24802 (N_24802,N_23303,N_22878);
nor U24803 (N_24803,N_23623,N_23033);
xor U24804 (N_24804,N_23249,N_23226);
xnor U24805 (N_24805,N_22849,N_23265);
nand U24806 (N_24806,N_23247,N_22571);
and U24807 (N_24807,N_23108,N_22820);
xnor U24808 (N_24808,N_22527,N_23746);
and U24809 (N_24809,N_23610,N_22767);
and U24810 (N_24810,N_22502,N_22810);
nor U24811 (N_24811,N_22596,N_22773);
xor U24812 (N_24812,N_22729,N_22606);
xnor U24813 (N_24813,N_23695,N_22686);
or U24814 (N_24814,N_23056,N_22935);
or U24815 (N_24815,N_22658,N_23563);
xor U24816 (N_24816,N_23298,N_23653);
nor U24817 (N_24817,N_23218,N_23155);
or U24818 (N_24818,N_23402,N_23367);
and U24819 (N_24819,N_23333,N_23084);
nand U24820 (N_24820,N_23384,N_22908);
or U24821 (N_24821,N_22706,N_22749);
nand U24822 (N_24822,N_22723,N_23260);
nand U24823 (N_24823,N_22627,N_22505);
nand U24824 (N_24824,N_23569,N_22535);
nand U24825 (N_24825,N_23392,N_23598);
xnor U24826 (N_24826,N_22791,N_23135);
xnor U24827 (N_24827,N_23288,N_23430);
or U24828 (N_24828,N_23518,N_22804);
or U24829 (N_24829,N_22790,N_23297);
and U24830 (N_24830,N_23398,N_23683);
or U24831 (N_24831,N_22692,N_22711);
nor U24832 (N_24832,N_23512,N_23314);
and U24833 (N_24833,N_23014,N_22628);
xnor U24834 (N_24834,N_23242,N_23451);
or U24835 (N_24835,N_22886,N_23457);
nor U24836 (N_24836,N_22977,N_23115);
and U24837 (N_24837,N_23029,N_22995);
nand U24838 (N_24838,N_22554,N_23278);
nand U24839 (N_24839,N_23478,N_23487);
or U24840 (N_24840,N_22839,N_22926);
and U24841 (N_24841,N_22865,N_23615);
xor U24842 (N_24842,N_23169,N_22673);
nor U24843 (N_24843,N_22816,N_23401);
and U24844 (N_24844,N_22905,N_22901);
or U24845 (N_24845,N_22839,N_22674);
and U24846 (N_24846,N_22943,N_22609);
and U24847 (N_24847,N_22741,N_23170);
xor U24848 (N_24848,N_23348,N_22882);
nor U24849 (N_24849,N_22640,N_22671);
xor U24850 (N_24850,N_23532,N_23324);
and U24851 (N_24851,N_22894,N_23421);
or U24852 (N_24852,N_23290,N_23529);
nand U24853 (N_24853,N_23091,N_22503);
nand U24854 (N_24854,N_23154,N_22724);
xnor U24855 (N_24855,N_23385,N_22516);
nor U24856 (N_24856,N_23143,N_23321);
nand U24857 (N_24857,N_22837,N_23701);
or U24858 (N_24858,N_22832,N_23711);
nand U24859 (N_24859,N_23001,N_23317);
nor U24860 (N_24860,N_23380,N_23355);
nor U24861 (N_24861,N_23160,N_23219);
nand U24862 (N_24862,N_23415,N_23674);
xor U24863 (N_24863,N_23644,N_23129);
xnor U24864 (N_24864,N_23709,N_23525);
or U24865 (N_24865,N_23698,N_23054);
nand U24866 (N_24866,N_22518,N_22842);
nor U24867 (N_24867,N_23710,N_22686);
or U24868 (N_24868,N_22831,N_22702);
or U24869 (N_24869,N_22604,N_22694);
and U24870 (N_24870,N_23159,N_22587);
xor U24871 (N_24871,N_23026,N_22862);
or U24872 (N_24872,N_23003,N_22708);
nand U24873 (N_24873,N_22767,N_23577);
or U24874 (N_24874,N_23177,N_23535);
nand U24875 (N_24875,N_23215,N_23197);
and U24876 (N_24876,N_22608,N_22627);
or U24877 (N_24877,N_23143,N_23331);
nand U24878 (N_24878,N_23728,N_23387);
or U24879 (N_24879,N_23326,N_22693);
xor U24880 (N_24880,N_22562,N_23003);
nor U24881 (N_24881,N_22857,N_23455);
or U24882 (N_24882,N_22585,N_22863);
and U24883 (N_24883,N_23024,N_23315);
and U24884 (N_24884,N_23307,N_22894);
nand U24885 (N_24885,N_23543,N_23509);
and U24886 (N_24886,N_22986,N_23453);
nand U24887 (N_24887,N_22919,N_23466);
and U24888 (N_24888,N_23421,N_23668);
and U24889 (N_24889,N_23182,N_23289);
nand U24890 (N_24890,N_23522,N_23163);
nand U24891 (N_24891,N_22744,N_23646);
nor U24892 (N_24892,N_22996,N_23105);
or U24893 (N_24893,N_23414,N_23043);
nand U24894 (N_24894,N_23408,N_23039);
nand U24895 (N_24895,N_23257,N_22851);
xor U24896 (N_24896,N_22782,N_23120);
and U24897 (N_24897,N_22945,N_23403);
nand U24898 (N_24898,N_22873,N_23694);
and U24899 (N_24899,N_23252,N_23123);
and U24900 (N_24900,N_22582,N_23563);
xor U24901 (N_24901,N_23739,N_23710);
nor U24902 (N_24902,N_22841,N_23540);
nor U24903 (N_24903,N_22964,N_23701);
nor U24904 (N_24904,N_23157,N_23261);
xnor U24905 (N_24905,N_23359,N_22982);
or U24906 (N_24906,N_23291,N_22832);
and U24907 (N_24907,N_23623,N_23508);
and U24908 (N_24908,N_23502,N_22733);
and U24909 (N_24909,N_23055,N_22979);
nand U24910 (N_24910,N_23223,N_23097);
nor U24911 (N_24911,N_23009,N_22738);
or U24912 (N_24912,N_22602,N_22813);
nor U24913 (N_24913,N_23156,N_23265);
xnor U24914 (N_24914,N_23085,N_23566);
nand U24915 (N_24915,N_22673,N_22714);
and U24916 (N_24916,N_23712,N_22546);
nor U24917 (N_24917,N_22918,N_23632);
xor U24918 (N_24918,N_23419,N_23287);
xnor U24919 (N_24919,N_23741,N_23135);
and U24920 (N_24920,N_22674,N_22538);
and U24921 (N_24921,N_22926,N_22835);
nor U24922 (N_24922,N_23517,N_22963);
nand U24923 (N_24923,N_23049,N_23042);
nor U24924 (N_24924,N_22774,N_23112);
and U24925 (N_24925,N_22744,N_23464);
or U24926 (N_24926,N_23308,N_23747);
and U24927 (N_24927,N_22851,N_23230);
nand U24928 (N_24928,N_23224,N_23208);
and U24929 (N_24929,N_23225,N_22991);
nor U24930 (N_24930,N_22983,N_23508);
nor U24931 (N_24931,N_22940,N_22808);
and U24932 (N_24932,N_23262,N_23294);
or U24933 (N_24933,N_23115,N_23718);
nor U24934 (N_24934,N_22632,N_23096);
or U24935 (N_24935,N_22763,N_22886);
nand U24936 (N_24936,N_23558,N_23295);
or U24937 (N_24937,N_22647,N_22898);
or U24938 (N_24938,N_22761,N_23168);
xnor U24939 (N_24939,N_23258,N_23598);
or U24940 (N_24940,N_23417,N_22508);
nor U24941 (N_24941,N_23583,N_22657);
xor U24942 (N_24942,N_23427,N_23603);
nand U24943 (N_24943,N_23624,N_23527);
and U24944 (N_24944,N_23305,N_23139);
nand U24945 (N_24945,N_22663,N_23666);
and U24946 (N_24946,N_23529,N_22857);
and U24947 (N_24947,N_23241,N_23504);
nand U24948 (N_24948,N_23723,N_23634);
and U24949 (N_24949,N_22911,N_22673);
and U24950 (N_24950,N_23370,N_22758);
xnor U24951 (N_24951,N_22795,N_23151);
and U24952 (N_24952,N_22505,N_22953);
nand U24953 (N_24953,N_23454,N_23301);
xor U24954 (N_24954,N_22979,N_22923);
nor U24955 (N_24955,N_22625,N_23389);
and U24956 (N_24956,N_23195,N_22557);
and U24957 (N_24957,N_23308,N_22773);
or U24958 (N_24958,N_23648,N_23749);
nor U24959 (N_24959,N_22969,N_22679);
and U24960 (N_24960,N_22659,N_22844);
xor U24961 (N_24961,N_23421,N_23378);
or U24962 (N_24962,N_22751,N_22589);
xor U24963 (N_24963,N_23163,N_23311);
xor U24964 (N_24964,N_22692,N_22843);
or U24965 (N_24965,N_23330,N_23230);
nand U24966 (N_24966,N_23625,N_23564);
xor U24967 (N_24967,N_23063,N_22686);
nor U24968 (N_24968,N_23147,N_23437);
nor U24969 (N_24969,N_22853,N_23147);
nor U24970 (N_24970,N_23058,N_23052);
xnor U24971 (N_24971,N_23185,N_22627);
nor U24972 (N_24972,N_23445,N_23360);
nand U24973 (N_24973,N_22865,N_22708);
and U24974 (N_24974,N_22936,N_22921);
nand U24975 (N_24975,N_22830,N_23525);
nand U24976 (N_24976,N_23077,N_22829);
xor U24977 (N_24977,N_22954,N_23373);
nand U24978 (N_24978,N_23449,N_23663);
nand U24979 (N_24979,N_23364,N_22540);
and U24980 (N_24980,N_23701,N_23186);
nor U24981 (N_24981,N_23422,N_22804);
nand U24982 (N_24982,N_23706,N_23542);
and U24983 (N_24983,N_23600,N_23189);
nor U24984 (N_24984,N_23125,N_23455);
and U24985 (N_24985,N_23155,N_23039);
xnor U24986 (N_24986,N_23400,N_22503);
and U24987 (N_24987,N_22558,N_23453);
or U24988 (N_24988,N_23666,N_23157);
or U24989 (N_24989,N_22965,N_22858);
xnor U24990 (N_24990,N_22759,N_23651);
nor U24991 (N_24991,N_23299,N_22770);
xnor U24992 (N_24992,N_23560,N_23168);
xnor U24993 (N_24993,N_23510,N_22608);
nor U24994 (N_24994,N_22504,N_23228);
nor U24995 (N_24995,N_23578,N_23739);
nand U24996 (N_24996,N_22955,N_23702);
nor U24997 (N_24997,N_23733,N_22672);
xnor U24998 (N_24998,N_23064,N_23326);
xnor U24999 (N_24999,N_23559,N_22968);
xnor UO_0 (O_0,N_24935,N_24319);
nor UO_1 (O_1,N_24544,N_23893);
xor UO_2 (O_2,N_24498,N_24385);
nand UO_3 (O_3,N_24764,N_24595);
or UO_4 (O_4,N_24482,N_24535);
or UO_5 (O_5,N_24077,N_24342);
and UO_6 (O_6,N_24897,N_24219);
nor UO_7 (O_7,N_24218,N_24555);
or UO_8 (O_8,N_24287,N_24628);
xor UO_9 (O_9,N_24979,N_24837);
and UO_10 (O_10,N_24965,N_24552);
or UO_11 (O_11,N_24075,N_24759);
xor UO_12 (O_12,N_23826,N_24952);
xor UO_13 (O_13,N_23852,N_23933);
xnor UO_14 (O_14,N_24557,N_23832);
xor UO_15 (O_15,N_24048,N_24084);
and UO_16 (O_16,N_23869,N_24254);
nand UO_17 (O_17,N_24514,N_24991);
or UO_18 (O_18,N_24869,N_24120);
nor UO_19 (O_19,N_24808,N_24064);
nor UO_20 (O_20,N_24594,N_24384);
nor UO_21 (O_21,N_23836,N_23866);
and UO_22 (O_22,N_24237,N_24839);
or UO_23 (O_23,N_24743,N_24649);
nor UO_24 (O_24,N_24549,N_24210);
xor UO_25 (O_25,N_24370,N_24556);
or UO_26 (O_26,N_24195,N_23990);
nor UO_27 (O_27,N_24000,N_24426);
or UO_28 (O_28,N_24113,N_24209);
nand UO_29 (O_29,N_24014,N_24564);
xnor UO_30 (O_30,N_24034,N_24081);
or UO_31 (O_31,N_24510,N_24019);
nor UO_32 (O_32,N_24364,N_24223);
or UO_33 (O_33,N_23850,N_23879);
and UO_34 (O_34,N_24292,N_24154);
and UO_35 (O_35,N_24003,N_24485);
and UO_36 (O_36,N_24422,N_23795);
nand UO_37 (O_37,N_24948,N_24133);
and UO_38 (O_38,N_24005,N_24169);
and UO_39 (O_39,N_23759,N_23931);
nor UO_40 (O_40,N_23958,N_24134);
and UO_41 (O_41,N_24647,N_24363);
nor UO_42 (O_42,N_24990,N_24011);
xnor UO_43 (O_43,N_23767,N_24956);
xnor UO_44 (O_44,N_24761,N_24311);
nor UO_45 (O_45,N_23975,N_24314);
or UO_46 (O_46,N_24610,N_24813);
nor UO_47 (O_47,N_24528,N_24155);
nor UO_48 (O_48,N_24161,N_24700);
nor UO_49 (O_49,N_24088,N_24351);
nand UO_50 (O_50,N_23865,N_24253);
and UO_51 (O_51,N_24864,N_23860);
or UO_52 (O_52,N_24454,N_24442);
nor UO_53 (O_53,N_24309,N_24726);
nor UO_54 (O_54,N_24644,N_23983);
xnor UO_55 (O_55,N_24488,N_24909);
xnor UO_56 (O_56,N_24786,N_24248);
or UO_57 (O_57,N_23867,N_23964);
or UO_58 (O_58,N_24770,N_24435);
xnor UO_59 (O_59,N_24554,N_24350);
nand UO_60 (O_60,N_23984,N_23912);
xor UO_61 (O_61,N_24741,N_24211);
and UO_62 (O_62,N_23907,N_24086);
nand UO_63 (O_63,N_24208,N_24879);
xor UO_64 (O_64,N_24505,N_23946);
nor UO_65 (O_65,N_24190,N_24410);
nand UO_66 (O_66,N_24188,N_24280);
nand UO_67 (O_67,N_24724,N_23878);
xnor UO_68 (O_68,N_24380,N_24127);
or UO_69 (O_69,N_24082,N_23947);
nor UO_70 (O_70,N_24964,N_24899);
and UO_71 (O_71,N_23972,N_24407);
xnor UO_72 (O_72,N_24215,N_24260);
nor UO_73 (O_73,N_24334,N_24492);
xor UO_74 (O_74,N_23848,N_24579);
and UO_75 (O_75,N_24642,N_24719);
or UO_76 (O_76,N_23986,N_24933);
or UO_77 (O_77,N_23856,N_24372);
xor UO_78 (O_78,N_23837,N_23903);
nor UO_79 (O_79,N_23979,N_23757);
nor UO_80 (O_80,N_24887,N_24315);
nor UO_81 (O_81,N_24341,N_24698);
or UO_82 (O_82,N_23835,N_24721);
xor UO_83 (O_83,N_24227,N_24776);
and UO_84 (O_84,N_24553,N_24112);
and UO_85 (O_85,N_24947,N_24576);
nor UO_86 (O_86,N_24852,N_23922);
or UO_87 (O_87,N_24335,N_23918);
and UO_88 (O_88,N_24284,N_24123);
nand UO_89 (O_89,N_24636,N_24397);
or UO_90 (O_90,N_24916,N_24265);
nor UO_91 (O_91,N_24274,N_24078);
xor UO_92 (O_92,N_24402,N_24691);
nor UO_93 (O_93,N_24129,N_24865);
xnor UO_94 (O_94,N_24033,N_24163);
xnor UO_95 (O_95,N_23994,N_24373);
nor UO_96 (O_96,N_24160,N_24906);
and UO_97 (O_97,N_24558,N_24794);
or UO_98 (O_98,N_24712,N_23809);
or UO_99 (O_99,N_24749,N_24360);
xor UO_100 (O_100,N_23960,N_23894);
nor UO_101 (O_101,N_24667,N_24295);
xor UO_102 (O_102,N_24357,N_24122);
nor UO_103 (O_103,N_23909,N_24844);
xor UO_104 (O_104,N_24585,N_24944);
nand UO_105 (O_105,N_24547,N_24496);
nand UO_106 (O_106,N_23873,N_23805);
xor UO_107 (O_107,N_24306,N_24013);
and UO_108 (O_108,N_24408,N_24308);
nand UO_109 (O_109,N_24942,N_23899);
and UO_110 (O_110,N_23940,N_24792);
nand UO_111 (O_111,N_24300,N_24670);
xnor UO_112 (O_112,N_24074,N_24103);
nand UO_113 (O_113,N_24149,N_24238);
nor UO_114 (O_114,N_24838,N_24597);
nand UO_115 (O_115,N_24958,N_24400);
nor UO_116 (O_116,N_24136,N_24425);
and UO_117 (O_117,N_24204,N_24125);
nor UO_118 (O_118,N_24520,N_24391);
nor UO_119 (O_119,N_24665,N_24497);
and UO_120 (O_120,N_24730,N_24060);
and UO_121 (O_121,N_24489,N_24825);
and UO_122 (O_122,N_24530,N_24340);
xor UO_123 (O_123,N_23913,N_24929);
xor UO_124 (O_124,N_24509,N_24826);
and UO_125 (O_125,N_24703,N_24932);
xnor UO_126 (O_126,N_24087,N_24023);
and UO_127 (O_127,N_24707,N_24881);
or UO_128 (O_128,N_23791,N_24867);
nand UO_129 (O_129,N_24258,N_24563);
and UO_130 (O_130,N_23987,N_23801);
or UO_131 (O_131,N_24212,N_24059);
or UO_132 (O_132,N_24091,N_23895);
or UO_133 (O_133,N_24255,N_24612);
nand UO_134 (O_134,N_24409,N_24207);
xor UO_135 (O_135,N_23838,N_24574);
nor UO_136 (O_136,N_24620,N_23849);
nor UO_137 (O_137,N_24898,N_24302);
or UO_138 (O_138,N_24429,N_24953);
or UO_139 (O_139,N_24616,N_23956);
or UO_140 (O_140,N_23788,N_24511);
and UO_141 (O_141,N_24097,N_24857);
nand UO_142 (O_142,N_24111,N_24889);
and UO_143 (O_143,N_24247,N_24180);
nor UO_144 (O_144,N_24008,N_23770);
xor UO_145 (O_145,N_24720,N_24821);
nand UO_146 (O_146,N_24239,N_24756);
or UO_147 (O_147,N_24690,N_24875);
or UO_148 (O_148,N_24971,N_24320);
or UO_149 (O_149,N_24571,N_24096);
nor UO_150 (O_150,N_24469,N_24467);
or UO_151 (O_151,N_24781,N_24949);
and UO_152 (O_152,N_24550,N_23973);
xor UO_153 (O_153,N_24045,N_23962);
nor UO_154 (O_154,N_24433,N_24858);
and UO_155 (O_155,N_24099,N_24827);
nand UO_156 (O_156,N_24962,N_24104);
nand UO_157 (O_157,N_24851,N_24181);
xor UO_158 (O_158,N_24465,N_24069);
xor UO_159 (O_159,N_24142,N_24184);
or UO_160 (O_160,N_24029,N_24974);
nor UO_161 (O_161,N_24891,N_24450);
xnor UO_162 (O_162,N_24714,N_24600);
xnor UO_163 (O_163,N_24472,N_23941);
nor UO_164 (O_164,N_24685,N_23910);
and UO_165 (O_165,N_24191,N_23796);
nand UO_166 (O_166,N_24533,N_23923);
or UO_167 (O_167,N_24683,N_23934);
xnor UO_168 (O_168,N_24396,N_24307);
nand UO_169 (O_169,N_24999,N_24829);
nor UO_170 (O_170,N_24645,N_24158);
nand UO_171 (O_171,N_24313,N_24710);
and UO_172 (O_172,N_24519,N_23814);
or UO_173 (O_173,N_24273,N_24796);
nor UO_174 (O_174,N_24785,N_24382);
nor UO_175 (O_175,N_23804,N_24871);
and UO_176 (O_176,N_24268,N_23874);
or UO_177 (O_177,N_24413,N_24592);
xor UO_178 (O_178,N_24083,N_23845);
nand UO_179 (O_179,N_24537,N_24298);
nand UO_180 (O_180,N_24684,N_24903);
nor UO_181 (O_181,N_24346,N_23891);
nand UO_182 (O_182,N_23995,N_23982);
xor UO_183 (O_183,N_23834,N_24961);
and UO_184 (O_184,N_24114,N_24568);
nand UO_185 (O_185,N_24596,N_24419);
xor UO_186 (O_186,N_24232,N_24850);
xnor UO_187 (O_187,N_23810,N_24922);
xor UO_188 (O_188,N_23752,N_24186);
xnor UO_189 (O_189,N_24175,N_24809);
or UO_190 (O_190,N_24228,N_24768);
nor UO_191 (O_191,N_24374,N_24878);
xnor UO_192 (O_192,N_24279,N_23840);
and UO_193 (O_193,N_24806,N_24230);
nand UO_194 (O_194,N_24805,N_24696);
or UO_195 (O_195,N_24404,N_24109);
nand UO_196 (O_196,N_24143,N_24895);
nand UO_197 (O_197,N_24460,N_24718);
nand UO_198 (O_198,N_24689,N_24742);
nand UO_199 (O_199,N_24976,N_24371);
or UO_200 (O_200,N_23883,N_24057);
or UO_201 (O_201,N_23841,N_23799);
nor UO_202 (O_202,N_24739,N_24412);
xor UO_203 (O_203,N_23925,N_24093);
or UO_204 (O_204,N_24967,N_23821);
and UO_205 (O_205,N_24673,N_24859);
and UO_206 (O_206,N_24441,N_24783);
nand UO_207 (O_207,N_24807,N_24729);
nor UO_208 (O_208,N_24733,N_23800);
xor UO_209 (O_209,N_24330,N_24249);
nand UO_210 (O_210,N_24527,N_24732);
or UO_211 (O_211,N_24836,N_24146);
or UO_212 (O_212,N_24677,N_24766);
nor UO_213 (O_213,N_24815,N_24312);
or UO_214 (O_214,N_24516,N_24686);
nand UO_215 (O_215,N_24892,N_24148);
nand UO_216 (O_216,N_24814,N_23996);
or UO_217 (O_217,N_24581,N_24010);
and UO_218 (O_218,N_24070,N_24561);
xor UO_219 (O_219,N_24572,N_23951);
nand UO_220 (O_220,N_24233,N_24092);
nand UO_221 (O_221,N_24451,N_24437);
xor UO_222 (O_222,N_24855,N_23900);
or UO_223 (O_223,N_24966,N_24376);
nor UO_224 (O_224,N_24995,N_24463);
or UO_225 (O_225,N_24760,N_24183);
and UO_226 (O_226,N_24235,N_24027);
or UO_227 (O_227,N_23785,N_24675);
and UO_228 (O_228,N_24316,N_24694);
nand UO_229 (O_229,N_23762,N_24073);
nor UO_230 (O_230,N_24757,N_24586);
nor UO_231 (O_231,N_24153,N_24926);
nor UO_232 (O_232,N_24882,N_24512);
or UO_233 (O_233,N_23977,N_24115);
nand UO_234 (O_234,N_24824,N_24353);
xnor UO_235 (O_235,N_24669,N_24870);
xnor UO_236 (O_236,N_24752,N_23875);
xnor UO_237 (O_237,N_24641,N_24007);
nand UO_238 (O_238,N_24750,N_24056);
nand UO_239 (O_239,N_24894,N_24477);
or UO_240 (O_240,N_24790,N_24840);
nand UO_241 (O_241,N_24399,N_23773);
nand UO_242 (O_242,N_24754,N_23755);
or UO_243 (O_243,N_24795,N_24793);
nand UO_244 (O_244,N_24480,N_24338);
nor UO_245 (O_245,N_23985,N_24635);
nand UO_246 (O_246,N_24196,N_23970);
xnor UO_247 (O_247,N_24668,N_24765);
and UO_248 (O_248,N_24189,N_23794);
and UO_249 (O_249,N_24993,N_24985);
and UO_250 (O_250,N_24379,N_24524);
nor UO_251 (O_251,N_24693,N_24411);
nor UO_252 (O_252,N_24621,N_24911);
nor UO_253 (O_253,N_24622,N_24919);
and UO_254 (O_254,N_23815,N_24333);
xnor UO_255 (O_255,N_24938,N_24748);
nand UO_256 (O_256,N_24130,N_23932);
and UO_257 (O_257,N_24646,N_24165);
xor UO_258 (O_258,N_24615,N_24521);
xnor UO_259 (O_259,N_23780,N_24883);
nand UO_260 (O_260,N_24625,N_24769);
and UO_261 (O_261,N_24475,N_23844);
and UO_262 (O_262,N_24992,N_24860);
xor UO_263 (O_263,N_24978,N_24963);
nor UO_264 (O_264,N_24630,N_23976);
nor UO_265 (O_265,N_24988,N_24174);
nand UO_266 (O_266,N_24162,N_24704);
nor UO_267 (O_267,N_24831,N_24406);
nor UO_268 (O_268,N_23974,N_24832);
nor UO_269 (O_269,N_24026,N_24224);
or UO_270 (O_270,N_24015,N_24303);
and UO_271 (O_271,N_24427,N_23811);
nand UO_272 (O_272,N_24043,N_24041);
xor UO_273 (O_273,N_24500,N_23766);
or UO_274 (O_274,N_24448,N_24318);
and UO_275 (O_275,N_24713,N_24588);
xor UO_276 (O_276,N_24727,N_24570);
and UO_277 (O_277,N_24278,N_24317);
or UO_278 (O_278,N_24659,N_24331);
and UO_279 (O_279,N_24434,N_24501);
xnor UO_280 (O_280,N_24355,N_24671);
nor UO_281 (O_281,N_24166,N_24002);
nor UO_282 (O_282,N_24305,N_24657);
nand UO_283 (O_283,N_24950,N_24022);
and UO_284 (O_284,N_24969,N_24904);
nor UO_285 (O_285,N_23786,N_24301);
or UO_286 (O_286,N_24167,N_23914);
nand UO_287 (O_287,N_24676,N_24152);
nand UO_288 (O_288,N_24359,N_24589);
nor UO_289 (O_289,N_23916,N_23959);
or UO_290 (O_290,N_24885,N_24050);
nand UO_291 (O_291,N_23955,N_24639);
nor UO_292 (O_292,N_24416,N_24325);
nand UO_293 (O_293,N_24150,N_23813);
nor UO_294 (O_294,N_24377,N_23760);
xnor UO_295 (O_295,N_24717,N_24737);
or UO_296 (O_296,N_23901,N_24170);
xnor UO_297 (O_297,N_24841,N_24297);
xor UO_298 (O_298,N_24495,N_24243);
nand UO_299 (O_299,N_24893,N_24140);
xnor UO_300 (O_300,N_24276,N_24066);
nor UO_301 (O_301,N_24951,N_23787);
and UO_302 (O_302,N_23858,N_23981);
nor UO_303 (O_303,N_24328,N_24734);
xor UO_304 (O_304,N_23846,N_24229);
and UO_305 (O_305,N_24605,N_24623);
and UO_306 (O_306,N_24632,N_24736);
nand UO_307 (O_307,N_24791,N_24819);
xnor UO_308 (O_308,N_24517,N_23870);
nor UO_309 (O_309,N_23950,N_24362);
xor UO_310 (O_310,N_24336,N_24924);
or UO_311 (O_311,N_24455,N_23880);
and UO_312 (O_312,N_24137,N_24456);
nand UO_313 (O_313,N_24823,N_24912);
or UO_314 (O_314,N_23953,N_24848);
nor UO_315 (O_315,N_23942,N_24051);
nand UO_316 (O_316,N_24337,N_24105);
nor UO_317 (O_317,N_24473,N_24423);
nor UO_318 (O_318,N_23831,N_24420);
nor UO_319 (O_319,N_23790,N_24004);
nand UO_320 (O_320,N_24271,N_24567);
and UO_321 (O_321,N_23871,N_24834);
nand UO_322 (O_322,N_24187,N_23864);
nand UO_323 (O_323,N_24666,N_24028);
or UO_324 (O_324,N_24250,N_24536);
xor UO_325 (O_325,N_24680,N_24076);
nand UO_326 (O_326,N_23756,N_24221);
nor UO_327 (O_327,N_24856,N_24296);
or UO_328 (O_328,N_24164,N_24144);
and UO_329 (O_329,N_24062,N_24545);
nand UO_330 (O_330,N_23969,N_24388);
or UO_331 (O_331,N_24812,N_24348);
and UO_332 (O_332,N_24529,N_24256);
xnor UO_333 (O_333,N_23993,N_24582);
or UO_334 (O_334,N_23827,N_24880);
nand UO_335 (O_335,N_24277,N_23989);
nor UO_336 (O_336,N_24876,N_24378);
nand UO_337 (O_337,N_24018,N_23847);
and UO_338 (O_338,N_24040,N_24468);
or UO_339 (O_339,N_24067,N_24058);
xnor UO_340 (O_340,N_23818,N_24987);
and UO_341 (O_341,N_24888,N_24257);
nand UO_342 (O_342,N_23798,N_23952);
xor UO_343 (O_343,N_24902,N_23954);
xor UO_344 (O_344,N_24656,N_23967);
xnor UO_345 (O_345,N_24798,N_24132);
xnor UO_346 (O_346,N_24282,N_24361);
nand UO_347 (O_347,N_24811,N_24598);
nand UO_348 (O_348,N_24868,N_24168);
and UO_349 (O_349,N_24936,N_24053);
and UO_350 (O_350,N_23884,N_24012);
and UO_351 (O_351,N_23877,N_23777);
or UO_352 (O_352,N_24415,N_24651);
and UO_353 (O_353,N_24095,N_24443);
nand UO_354 (O_354,N_24996,N_24593);
and UO_355 (O_355,N_24339,N_23781);
nand UO_356 (O_356,N_24231,N_24584);
xor UO_357 (O_357,N_24151,N_24205);
nor UO_358 (O_358,N_24159,N_24172);
or UO_359 (O_359,N_24395,N_23938);
or UO_360 (O_360,N_24513,N_24121);
nor UO_361 (O_361,N_24577,N_24197);
nor UO_362 (O_362,N_24998,N_24431);
and UO_363 (O_363,N_23802,N_24901);
nand UO_364 (O_364,N_24021,N_23862);
and UO_365 (O_365,N_24853,N_24539);
xnor UO_366 (O_366,N_23991,N_23929);
and UO_367 (O_367,N_24661,N_24835);
nand UO_368 (O_368,N_23764,N_24744);
xnor UO_369 (O_369,N_23758,N_24927);
nor UO_370 (O_370,N_23753,N_23876);
or UO_371 (O_371,N_23924,N_24886);
or UO_372 (O_372,N_24955,N_23926);
nand UO_373 (O_373,N_24462,N_24611);
nor UO_374 (O_374,N_24182,N_24507);
nand UO_375 (O_375,N_23763,N_24787);
and UO_376 (O_376,N_24128,N_24080);
or UO_377 (O_377,N_24525,N_23971);
xnor UO_378 (O_378,N_24063,N_24715);
or UO_379 (O_379,N_24695,N_24777);
nor UO_380 (O_380,N_23965,N_24913);
nand UO_381 (O_381,N_24367,N_23750);
nor UO_382 (O_382,N_24236,N_24025);
xnor UO_383 (O_383,N_24368,N_24432);
and UO_384 (O_384,N_23908,N_24483);
and UO_385 (O_385,N_24071,N_24046);
xnor UO_386 (O_386,N_24728,N_23920);
nor UO_387 (O_387,N_24173,N_24687);
nand UO_388 (O_388,N_24650,N_24800);
nand UO_389 (O_389,N_24458,N_24398);
or UO_390 (O_390,N_24716,N_24917);
or UO_391 (O_391,N_24030,N_24590);
and UO_392 (O_392,N_24818,N_23935);
nand UO_393 (O_393,N_23968,N_24405);
nor UO_394 (O_394,N_24846,N_24089);
nor UO_395 (O_395,N_23919,N_24440);
nand UO_396 (O_396,N_24799,N_24006);
and UO_397 (O_397,N_24107,N_23839);
nor UO_398 (O_398,N_24466,N_24873);
xnor UO_399 (O_399,N_24702,N_24643);
nor UO_400 (O_400,N_24481,N_23863);
nor UO_401 (O_401,N_23797,N_24038);
xnor UO_402 (O_402,N_24179,N_24141);
and UO_403 (O_403,N_24663,N_23754);
and UO_404 (O_404,N_24634,N_24609);
nor UO_405 (O_405,N_24679,N_24866);
nand UO_406 (O_406,N_24531,N_23775);
xor UO_407 (O_407,N_24775,N_24915);
nor UO_408 (O_408,N_24890,N_24241);
nand UO_409 (O_409,N_23896,N_23906);
xor UO_410 (O_410,N_24753,N_23782);
and UO_411 (O_411,N_24607,N_24709);
or UO_412 (O_412,N_24266,N_24220);
or UO_413 (O_413,N_24193,N_23779);
nand UO_414 (O_414,N_24997,N_24185);
and UO_415 (O_415,N_24072,N_24110);
nand UO_416 (O_416,N_23817,N_23886);
and UO_417 (O_417,N_23905,N_24036);
nor UO_418 (O_418,N_24655,N_24272);
nor UO_419 (O_419,N_23825,N_24242);
and UO_420 (O_420,N_24706,N_23793);
xnor UO_421 (O_421,N_24773,N_24941);
nor UO_422 (O_422,N_24559,N_24560);
nand UO_423 (O_423,N_24569,N_23768);
xnor UO_424 (O_424,N_24578,N_24608);
or UO_425 (O_425,N_24619,N_24986);
and UO_426 (O_426,N_24200,N_24270);
nor UO_427 (O_427,N_24478,N_24872);
nand UO_428 (O_428,N_24024,N_23928);
xnor UO_429 (O_429,N_23751,N_24214);
xor UO_430 (O_430,N_24293,N_24614);
nor UO_431 (O_431,N_24541,N_24369);
nand UO_432 (O_432,N_24863,N_24366);
nor UO_433 (O_433,N_24401,N_24439);
and UO_434 (O_434,N_24711,N_23892);
nor UO_435 (O_435,N_24387,N_24327);
nand UO_436 (O_436,N_24534,N_24065);
or UO_437 (O_437,N_24329,N_24445);
or UO_438 (O_438,N_23859,N_24980);
or UO_439 (O_439,N_24658,N_24213);
nor UO_440 (O_440,N_24383,N_23853);
or UO_441 (O_441,N_24147,N_24830);
and UO_442 (O_442,N_24772,N_23784);
and UO_443 (O_443,N_24470,N_24349);
or UO_444 (O_444,N_24847,N_24090);
and UO_445 (O_445,N_24874,N_24526);
nand UO_446 (O_446,N_24506,N_24820);
nand UO_447 (O_447,N_24626,N_24983);
or UO_448 (O_448,N_24989,N_24583);
xor UO_449 (O_449,N_24119,N_24202);
nand UO_450 (O_450,N_23819,N_24833);
nand UO_451 (O_451,N_24801,N_24203);
nand UO_452 (O_452,N_23854,N_24251);
nand UO_453 (O_453,N_24810,N_24900);
or UO_454 (O_454,N_24587,N_24491);
and UO_455 (O_455,N_24981,N_23812);
or UO_456 (O_456,N_24921,N_24476);
xnor UO_457 (O_457,N_24637,N_23963);
nand UO_458 (O_458,N_24975,N_23930);
nor UO_459 (O_459,N_24323,N_24288);
xor UO_460 (O_460,N_23937,N_24779);
and UO_461 (O_461,N_24457,N_24939);
or UO_462 (O_462,N_24972,N_24740);
xnor UO_463 (O_463,N_23915,N_24016);
nand UO_464 (O_464,N_24931,N_24861);
xor UO_465 (O_465,N_24156,N_24290);
or UO_466 (O_466,N_23792,N_24375);
nand UO_467 (O_467,N_24201,N_24106);
nor UO_468 (O_468,N_23774,N_24660);
nor UO_469 (O_469,N_24640,N_24421);
xnor UO_470 (O_470,N_24042,N_24862);
xor UO_471 (O_471,N_24662,N_23889);
xnor UO_472 (O_472,N_23778,N_24751);
nor UO_473 (O_473,N_23921,N_24782);
xor UO_474 (O_474,N_24108,N_24049);
or UO_475 (O_475,N_23961,N_24653);
or UO_476 (O_476,N_23997,N_24784);
nor UO_477 (O_477,N_23917,N_24177);
xor UO_478 (O_478,N_24322,N_24192);
or UO_479 (O_479,N_24055,N_24735);
nand UO_480 (O_480,N_24244,N_24816);
xor UO_481 (O_481,N_24044,N_24849);
and UO_482 (O_482,N_24746,N_24347);
xnor UO_483 (O_483,N_24697,N_24682);
nor UO_484 (O_484,N_23868,N_24326);
or UO_485 (O_485,N_23887,N_24543);
nor UO_486 (O_486,N_24771,N_23936);
nor UO_487 (O_487,N_24145,N_24471);
nor UO_488 (O_488,N_24094,N_24701);
nor UO_489 (O_489,N_24068,N_24788);
xnor UO_490 (O_490,N_24914,N_24438);
or UO_491 (O_491,N_24286,N_24358);
or UO_492 (O_492,N_24960,N_24452);
nand UO_493 (O_493,N_24424,N_24907);
xor UO_494 (O_494,N_24523,N_24310);
xor UO_495 (O_495,N_23833,N_24101);
or UO_496 (O_496,N_24386,N_24100);
and UO_497 (O_497,N_24403,N_23882);
nand UO_498 (O_498,N_24479,N_24522);
and UO_499 (O_499,N_24722,N_24356);
and UO_500 (O_500,N_24896,N_24035);
xor UO_501 (O_501,N_23992,N_24446);
nand UO_502 (O_502,N_24264,N_24780);
and UO_503 (O_503,N_24447,N_23949);
xor UO_504 (O_504,N_24240,N_24603);
nand UO_505 (O_505,N_24344,N_24925);
and UO_506 (O_506,N_24994,N_24117);
nor UO_507 (O_507,N_24393,N_24131);
and UO_508 (O_508,N_24490,N_24171);
nor UO_509 (O_509,N_24606,N_24803);
or UO_510 (O_510,N_24032,N_24453);
or UO_511 (O_511,N_24428,N_24854);
or UO_512 (O_512,N_24817,N_24345);
xor UO_513 (O_513,N_23888,N_24705);
nand UO_514 (O_514,N_23771,N_24943);
or UO_515 (O_515,N_24102,N_23904);
and UO_516 (O_516,N_24575,N_24654);
xor UO_517 (O_517,N_24194,N_24503);
nand UO_518 (O_518,N_24139,N_24098);
nor UO_519 (O_519,N_24459,N_24381);
nand UO_520 (O_520,N_24802,N_24804);
nand UO_521 (O_521,N_23944,N_24085);
nand UO_522 (O_522,N_23822,N_24017);
and UO_523 (O_523,N_24499,N_24540);
nor UO_524 (O_524,N_24842,N_24267);
nand UO_525 (O_525,N_23806,N_24681);
nor UO_526 (O_526,N_24047,N_23872);
or UO_527 (O_527,N_23808,N_24283);
nor UO_528 (O_528,N_24299,N_24052);
nand UO_529 (O_529,N_24157,N_24672);
nand UO_530 (O_530,N_23828,N_24877);
nand UO_531 (O_531,N_24474,N_24464);
xnor UO_532 (O_532,N_24580,N_24920);
nand UO_533 (O_533,N_24226,N_24738);
xor UO_534 (O_534,N_23776,N_24225);
and UO_535 (O_535,N_24518,N_23898);
nor UO_536 (O_536,N_23851,N_24054);
and UO_537 (O_537,N_24390,N_24745);
nor UO_538 (O_538,N_24602,N_24648);
or UO_539 (O_539,N_24269,N_23939);
nand UO_540 (O_540,N_23966,N_24430);
nor UO_541 (O_541,N_24332,N_23761);
nor UO_542 (O_542,N_24449,N_24486);
and UO_543 (O_543,N_24797,N_23957);
nand UO_544 (O_544,N_24725,N_24343);
xor UO_545 (O_545,N_24285,N_24199);
nand UO_546 (O_546,N_24928,N_23945);
nand UO_547 (O_547,N_24222,N_24542);
and UO_548 (O_548,N_24418,N_24638);
and UO_549 (O_549,N_24982,N_24918);
nand UO_550 (O_550,N_24444,N_24905);
xnor UO_551 (O_551,N_23927,N_23861);
and UO_552 (O_552,N_24674,N_24234);
or UO_553 (O_553,N_24217,N_24262);
nor UO_554 (O_554,N_23807,N_24352);
and UO_555 (O_555,N_24354,N_24394);
and UO_556 (O_556,N_24259,N_24763);
xnor UO_557 (O_557,N_23911,N_24246);
and UO_558 (O_558,N_24789,N_24261);
and UO_559 (O_559,N_24774,N_24977);
xor UO_560 (O_560,N_23783,N_24532);
and UO_561 (O_561,N_23843,N_24546);
nor UO_562 (O_562,N_24116,N_24688);
nand UO_563 (O_563,N_24389,N_24664);
and UO_564 (O_564,N_24778,N_24624);
nor UO_565 (O_565,N_23842,N_24039);
nor UO_566 (O_566,N_24216,N_24617);
xor UO_567 (O_567,N_24959,N_24138);
nor UO_568 (O_568,N_24828,N_24484);
xor UO_569 (O_569,N_24954,N_24631);
or UO_570 (O_570,N_23897,N_23999);
and UO_571 (O_571,N_24291,N_24627);
xnor UO_572 (O_572,N_24591,N_24945);
nand UO_573 (O_573,N_24946,N_24822);
xor UO_574 (O_574,N_23943,N_24417);
xnor UO_575 (O_575,N_24613,N_24762);
or UO_576 (O_576,N_24079,N_23857);
or UO_577 (O_577,N_24884,N_24599);
or UO_578 (O_578,N_23881,N_23772);
and UO_579 (O_579,N_24263,N_24304);
nor UO_580 (O_580,N_24061,N_24562);
nor UO_581 (O_581,N_24678,N_24124);
xnor UO_582 (O_582,N_23816,N_24487);
xnor UO_583 (O_583,N_24135,N_24984);
xor UO_584 (O_584,N_24494,N_24321);
nand UO_585 (O_585,N_24940,N_24566);
nor UO_586 (O_586,N_24843,N_24565);
xnor UO_587 (O_587,N_23823,N_24031);
and UO_588 (O_588,N_23824,N_24957);
nand UO_589 (O_589,N_24910,N_24198);
or UO_590 (O_590,N_24731,N_23885);
nand UO_591 (O_591,N_24289,N_24118);
nand UO_592 (O_592,N_24037,N_23980);
or UO_593 (O_593,N_23820,N_23830);
or UO_594 (O_594,N_23988,N_24502);
or UO_595 (O_595,N_24206,N_24923);
xnor UO_596 (O_596,N_23789,N_24508);
and UO_597 (O_597,N_24414,N_24324);
nor UO_598 (O_598,N_24767,N_24937);
nor UO_599 (O_599,N_24845,N_23890);
and UO_600 (O_600,N_24281,N_24758);
xor UO_601 (O_601,N_24020,N_24436);
xor UO_602 (O_602,N_24548,N_24493);
nand UO_603 (O_603,N_24392,N_23829);
and UO_604 (O_604,N_24934,N_24755);
nand UO_605 (O_605,N_24461,N_24633);
and UO_606 (O_606,N_24275,N_24968);
nor UO_607 (O_607,N_24699,N_24629);
nand UO_608 (O_608,N_23803,N_24604);
and UO_609 (O_609,N_24176,N_24652);
and UO_610 (O_610,N_24970,N_24365);
nand UO_611 (O_611,N_24504,N_24708);
xor UO_612 (O_612,N_24973,N_24538);
nor UO_613 (O_613,N_24551,N_24252);
nand UO_614 (O_614,N_23902,N_24573);
nand UO_615 (O_615,N_24747,N_24009);
xnor UO_616 (O_616,N_24126,N_24692);
or UO_617 (O_617,N_23998,N_24245);
xor UO_618 (O_618,N_24178,N_23948);
or UO_619 (O_619,N_23765,N_24908);
nor UO_620 (O_620,N_24723,N_23769);
xnor UO_621 (O_621,N_24930,N_23855);
xor UO_622 (O_622,N_24294,N_24515);
xnor UO_623 (O_623,N_24618,N_24601);
xor UO_624 (O_624,N_24001,N_23978);
or UO_625 (O_625,N_24440,N_24469);
xor UO_626 (O_626,N_24759,N_24195);
nor UO_627 (O_627,N_24416,N_24816);
nand UO_628 (O_628,N_24140,N_24317);
and UO_629 (O_629,N_23976,N_24606);
and UO_630 (O_630,N_24286,N_24161);
nor UO_631 (O_631,N_24501,N_24517);
nor UO_632 (O_632,N_24552,N_23928);
or UO_633 (O_633,N_24585,N_23987);
or UO_634 (O_634,N_24544,N_23801);
nand UO_635 (O_635,N_24021,N_24353);
xnor UO_636 (O_636,N_24788,N_24018);
nor UO_637 (O_637,N_24839,N_24683);
or UO_638 (O_638,N_24593,N_24096);
or UO_639 (O_639,N_23856,N_23913);
nor UO_640 (O_640,N_24640,N_24113);
and UO_641 (O_641,N_24623,N_24019);
nand UO_642 (O_642,N_24958,N_23782);
nand UO_643 (O_643,N_24837,N_24188);
and UO_644 (O_644,N_23807,N_24748);
xor UO_645 (O_645,N_24365,N_23759);
and UO_646 (O_646,N_24350,N_24979);
nor UO_647 (O_647,N_24662,N_23877);
and UO_648 (O_648,N_24292,N_24342);
and UO_649 (O_649,N_24209,N_24151);
and UO_650 (O_650,N_23845,N_23841);
or UO_651 (O_651,N_24720,N_23846);
nor UO_652 (O_652,N_24700,N_24220);
or UO_653 (O_653,N_24217,N_24673);
nor UO_654 (O_654,N_24663,N_24389);
or UO_655 (O_655,N_24703,N_24228);
nor UO_656 (O_656,N_24697,N_24034);
nand UO_657 (O_657,N_24404,N_24767);
xor UO_658 (O_658,N_24904,N_24570);
xor UO_659 (O_659,N_24645,N_24948);
xnor UO_660 (O_660,N_24557,N_24189);
nor UO_661 (O_661,N_24388,N_24719);
or UO_662 (O_662,N_24671,N_23970);
and UO_663 (O_663,N_24759,N_24910);
or UO_664 (O_664,N_24428,N_24170);
nor UO_665 (O_665,N_24755,N_24861);
or UO_666 (O_666,N_24732,N_23764);
or UO_667 (O_667,N_24043,N_23805);
nand UO_668 (O_668,N_24051,N_24886);
or UO_669 (O_669,N_24617,N_24858);
and UO_670 (O_670,N_23751,N_24381);
nor UO_671 (O_671,N_24222,N_24178);
nand UO_672 (O_672,N_24854,N_23997);
nand UO_673 (O_673,N_23996,N_24233);
xor UO_674 (O_674,N_24609,N_23964);
nand UO_675 (O_675,N_24384,N_23888);
nor UO_676 (O_676,N_24849,N_24299);
xnor UO_677 (O_677,N_23975,N_24056);
nor UO_678 (O_678,N_24894,N_24920);
nand UO_679 (O_679,N_24581,N_24262);
xor UO_680 (O_680,N_24217,N_24115);
xor UO_681 (O_681,N_24414,N_24235);
or UO_682 (O_682,N_24066,N_24414);
xnor UO_683 (O_683,N_24148,N_24678);
or UO_684 (O_684,N_24519,N_24308);
and UO_685 (O_685,N_23830,N_24729);
and UO_686 (O_686,N_24166,N_24018);
xor UO_687 (O_687,N_24497,N_23756);
or UO_688 (O_688,N_24634,N_23764);
nor UO_689 (O_689,N_24900,N_24685);
nand UO_690 (O_690,N_24665,N_24760);
nor UO_691 (O_691,N_23908,N_24427);
or UO_692 (O_692,N_24259,N_24616);
xor UO_693 (O_693,N_24627,N_24876);
or UO_694 (O_694,N_24632,N_24100);
xnor UO_695 (O_695,N_24221,N_24041);
or UO_696 (O_696,N_24522,N_24974);
nand UO_697 (O_697,N_24065,N_24121);
nand UO_698 (O_698,N_24884,N_24410);
nand UO_699 (O_699,N_24396,N_24039);
nand UO_700 (O_700,N_24740,N_24394);
or UO_701 (O_701,N_23785,N_24039);
or UO_702 (O_702,N_24534,N_23795);
nand UO_703 (O_703,N_24179,N_24774);
nor UO_704 (O_704,N_24714,N_24532);
nor UO_705 (O_705,N_24335,N_23997);
or UO_706 (O_706,N_24057,N_24847);
nor UO_707 (O_707,N_24799,N_24372);
and UO_708 (O_708,N_24910,N_24474);
and UO_709 (O_709,N_24463,N_24092);
nor UO_710 (O_710,N_23956,N_23929);
nand UO_711 (O_711,N_24255,N_23989);
or UO_712 (O_712,N_24429,N_23921);
nor UO_713 (O_713,N_24653,N_24493);
xnor UO_714 (O_714,N_23955,N_24335);
and UO_715 (O_715,N_24565,N_24331);
and UO_716 (O_716,N_24949,N_24137);
xor UO_717 (O_717,N_24849,N_24964);
and UO_718 (O_718,N_24346,N_24462);
and UO_719 (O_719,N_23837,N_24581);
or UO_720 (O_720,N_24728,N_24277);
and UO_721 (O_721,N_24912,N_24636);
and UO_722 (O_722,N_23970,N_23973);
nor UO_723 (O_723,N_24438,N_24743);
or UO_724 (O_724,N_24941,N_24004);
xnor UO_725 (O_725,N_24740,N_24032);
nand UO_726 (O_726,N_23867,N_24447);
and UO_727 (O_727,N_23795,N_24795);
nand UO_728 (O_728,N_24284,N_23786);
or UO_729 (O_729,N_24506,N_23958);
or UO_730 (O_730,N_23770,N_24697);
and UO_731 (O_731,N_23964,N_24161);
and UO_732 (O_732,N_24359,N_24895);
and UO_733 (O_733,N_24020,N_24078);
or UO_734 (O_734,N_24192,N_24019);
or UO_735 (O_735,N_24723,N_24892);
xor UO_736 (O_736,N_23817,N_23786);
nor UO_737 (O_737,N_24864,N_24484);
xnor UO_738 (O_738,N_23835,N_23977);
nor UO_739 (O_739,N_24549,N_24860);
and UO_740 (O_740,N_23961,N_24230);
xnor UO_741 (O_741,N_24374,N_24873);
and UO_742 (O_742,N_24419,N_24005);
nand UO_743 (O_743,N_24593,N_24734);
nand UO_744 (O_744,N_24815,N_24270);
xnor UO_745 (O_745,N_24617,N_24370);
nor UO_746 (O_746,N_24113,N_24641);
nor UO_747 (O_747,N_24227,N_24306);
and UO_748 (O_748,N_23925,N_24806);
and UO_749 (O_749,N_24392,N_24352);
nor UO_750 (O_750,N_24474,N_24456);
nand UO_751 (O_751,N_23857,N_24649);
nand UO_752 (O_752,N_24819,N_24696);
or UO_753 (O_753,N_24512,N_24953);
and UO_754 (O_754,N_24989,N_24312);
and UO_755 (O_755,N_24822,N_24597);
and UO_756 (O_756,N_24614,N_23802);
nor UO_757 (O_757,N_23989,N_24437);
or UO_758 (O_758,N_23858,N_24897);
nor UO_759 (O_759,N_24956,N_23885);
or UO_760 (O_760,N_24727,N_24018);
and UO_761 (O_761,N_23826,N_24614);
nand UO_762 (O_762,N_23949,N_24298);
xnor UO_763 (O_763,N_24850,N_24784);
xnor UO_764 (O_764,N_24103,N_24652);
and UO_765 (O_765,N_24209,N_24382);
nand UO_766 (O_766,N_23798,N_24878);
nand UO_767 (O_767,N_24510,N_24238);
nor UO_768 (O_768,N_24521,N_24023);
nor UO_769 (O_769,N_24240,N_24385);
and UO_770 (O_770,N_24159,N_24102);
and UO_771 (O_771,N_24816,N_24318);
nor UO_772 (O_772,N_24780,N_24011);
nor UO_773 (O_773,N_24569,N_24818);
nor UO_774 (O_774,N_24378,N_24971);
nand UO_775 (O_775,N_24418,N_24788);
or UO_776 (O_776,N_24959,N_24716);
nor UO_777 (O_777,N_24457,N_24896);
and UO_778 (O_778,N_24632,N_24403);
or UO_779 (O_779,N_24093,N_24344);
and UO_780 (O_780,N_24035,N_24549);
xnor UO_781 (O_781,N_24890,N_24402);
and UO_782 (O_782,N_24812,N_24250);
nand UO_783 (O_783,N_24198,N_24732);
or UO_784 (O_784,N_24500,N_24167);
xor UO_785 (O_785,N_24559,N_24600);
xnor UO_786 (O_786,N_23959,N_24735);
xnor UO_787 (O_787,N_24320,N_24155);
xor UO_788 (O_788,N_24753,N_24934);
nor UO_789 (O_789,N_24008,N_24572);
xnor UO_790 (O_790,N_24989,N_24147);
xor UO_791 (O_791,N_23839,N_23921);
or UO_792 (O_792,N_24367,N_24910);
xnor UO_793 (O_793,N_24110,N_24631);
or UO_794 (O_794,N_24629,N_24435);
nand UO_795 (O_795,N_24800,N_23872);
nand UO_796 (O_796,N_23899,N_24232);
and UO_797 (O_797,N_24974,N_24741);
nor UO_798 (O_798,N_24831,N_24324);
nand UO_799 (O_799,N_23788,N_24115);
xnor UO_800 (O_800,N_24698,N_24577);
xnor UO_801 (O_801,N_24249,N_24851);
and UO_802 (O_802,N_24258,N_24171);
xnor UO_803 (O_803,N_24436,N_24303);
and UO_804 (O_804,N_24311,N_24390);
xnor UO_805 (O_805,N_23869,N_24684);
and UO_806 (O_806,N_24871,N_23911);
nand UO_807 (O_807,N_24158,N_24025);
and UO_808 (O_808,N_24783,N_23943);
nand UO_809 (O_809,N_24579,N_24046);
nor UO_810 (O_810,N_23999,N_24640);
nand UO_811 (O_811,N_24744,N_24713);
xor UO_812 (O_812,N_24503,N_24013);
nor UO_813 (O_813,N_24690,N_23983);
xor UO_814 (O_814,N_24256,N_24139);
and UO_815 (O_815,N_24757,N_24688);
nand UO_816 (O_816,N_23907,N_24335);
or UO_817 (O_817,N_23772,N_24113);
or UO_818 (O_818,N_24432,N_23931);
nor UO_819 (O_819,N_24116,N_24833);
nand UO_820 (O_820,N_24097,N_23769);
nor UO_821 (O_821,N_24566,N_24810);
nor UO_822 (O_822,N_23941,N_24314);
nand UO_823 (O_823,N_24766,N_23776);
and UO_824 (O_824,N_24118,N_24866);
nor UO_825 (O_825,N_24181,N_23791);
and UO_826 (O_826,N_24269,N_24723);
nand UO_827 (O_827,N_23967,N_23804);
xnor UO_828 (O_828,N_24695,N_23963);
and UO_829 (O_829,N_23793,N_24548);
nor UO_830 (O_830,N_24497,N_24596);
and UO_831 (O_831,N_23918,N_24008);
nand UO_832 (O_832,N_24094,N_23752);
nand UO_833 (O_833,N_23888,N_24700);
nor UO_834 (O_834,N_24144,N_24495);
nor UO_835 (O_835,N_24521,N_23853);
xor UO_836 (O_836,N_23968,N_23826);
nor UO_837 (O_837,N_24534,N_24419);
or UO_838 (O_838,N_24990,N_24938);
or UO_839 (O_839,N_24546,N_24040);
or UO_840 (O_840,N_24029,N_24850);
and UO_841 (O_841,N_24698,N_24193);
nand UO_842 (O_842,N_24883,N_24754);
xnor UO_843 (O_843,N_24092,N_23766);
nand UO_844 (O_844,N_23816,N_24780);
xor UO_845 (O_845,N_23931,N_24124);
nor UO_846 (O_846,N_24129,N_24334);
xor UO_847 (O_847,N_24371,N_24110);
and UO_848 (O_848,N_24738,N_23991);
xnor UO_849 (O_849,N_24828,N_23910);
or UO_850 (O_850,N_23872,N_24079);
xnor UO_851 (O_851,N_24163,N_24319);
nor UO_852 (O_852,N_23955,N_24822);
nand UO_853 (O_853,N_24826,N_24722);
nor UO_854 (O_854,N_24801,N_24145);
and UO_855 (O_855,N_24551,N_24799);
xor UO_856 (O_856,N_24327,N_24602);
and UO_857 (O_857,N_24497,N_23800);
xor UO_858 (O_858,N_24713,N_24928);
xnor UO_859 (O_859,N_24683,N_24778);
nor UO_860 (O_860,N_23850,N_23792);
or UO_861 (O_861,N_24208,N_24125);
xnor UO_862 (O_862,N_24378,N_24036);
or UO_863 (O_863,N_24007,N_24280);
xor UO_864 (O_864,N_24367,N_24439);
nand UO_865 (O_865,N_23911,N_24718);
or UO_866 (O_866,N_24354,N_24382);
nand UO_867 (O_867,N_24428,N_23993);
nand UO_868 (O_868,N_24405,N_24956);
nand UO_869 (O_869,N_23813,N_23795);
and UO_870 (O_870,N_24790,N_24223);
nor UO_871 (O_871,N_23963,N_24368);
and UO_872 (O_872,N_23859,N_24846);
nor UO_873 (O_873,N_24184,N_24965);
nand UO_874 (O_874,N_23936,N_24503);
nand UO_875 (O_875,N_24780,N_23814);
xor UO_876 (O_876,N_23927,N_24925);
and UO_877 (O_877,N_23839,N_24257);
nand UO_878 (O_878,N_24963,N_24932);
xor UO_879 (O_879,N_24496,N_24155);
nand UO_880 (O_880,N_23799,N_24696);
nand UO_881 (O_881,N_24118,N_23862);
xor UO_882 (O_882,N_24730,N_23767);
or UO_883 (O_883,N_24014,N_24786);
and UO_884 (O_884,N_24710,N_23777);
xor UO_885 (O_885,N_24879,N_24655);
nor UO_886 (O_886,N_24982,N_24995);
xor UO_887 (O_887,N_23773,N_24487);
xnor UO_888 (O_888,N_24447,N_24727);
and UO_889 (O_889,N_24397,N_23815);
xnor UO_890 (O_890,N_24275,N_24075);
xnor UO_891 (O_891,N_24353,N_24375);
and UO_892 (O_892,N_24963,N_24838);
or UO_893 (O_893,N_24016,N_23971);
nand UO_894 (O_894,N_24147,N_24062);
nor UO_895 (O_895,N_24887,N_24297);
and UO_896 (O_896,N_23913,N_24867);
and UO_897 (O_897,N_24087,N_24500);
or UO_898 (O_898,N_24316,N_24928);
nand UO_899 (O_899,N_24930,N_24692);
nor UO_900 (O_900,N_24598,N_24099);
nor UO_901 (O_901,N_23933,N_24539);
nand UO_902 (O_902,N_24167,N_24427);
nand UO_903 (O_903,N_24015,N_24120);
and UO_904 (O_904,N_24830,N_24708);
nand UO_905 (O_905,N_24111,N_24235);
nor UO_906 (O_906,N_24203,N_24022);
nor UO_907 (O_907,N_24525,N_24004);
nor UO_908 (O_908,N_24259,N_24385);
nor UO_909 (O_909,N_24132,N_23941);
nor UO_910 (O_910,N_24918,N_24602);
xnor UO_911 (O_911,N_24660,N_24320);
or UO_912 (O_912,N_23883,N_23893);
nor UO_913 (O_913,N_24984,N_24447);
xor UO_914 (O_914,N_24978,N_24576);
xnor UO_915 (O_915,N_24412,N_24012);
and UO_916 (O_916,N_24434,N_24795);
or UO_917 (O_917,N_24159,N_23954);
nand UO_918 (O_918,N_24855,N_24652);
nor UO_919 (O_919,N_23832,N_23792);
and UO_920 (O_920,N_24498,N_24547);
nand UO_921 (O_921,N_24686,N_24867);
nor UO_922 (O_922,N_23902,N_24937);
xor UO_923 (O_923,N_24285,N_24621);
xnor UO_924 (O_924,N_24125,N_24680);
nor UO_925 (O_925,N_24735,N_24426);
or UO_926 (O_926,N_24138,N_24333);
or UO_927 (O_927,N_24242,N_24639);
xnor UO_928 (O_928,N_24439,N_24060);
and UO_929 (O_929,N_24674,N_23907);
or UO_930 (O_930,N_24666,N_24826);
and UO_931 (O_931,N_24040,N_24985);
xor UO_932 (O_932,N_23758,N_23765);
nand UO_933 (O_933,N_24922,N_23863);
xor UO_934 (O_934,N_24316,N_24945);
and UO_935 (O_935,N_24956,N_24545);
and UO_936 (O_936,N_24759,N_24261);
and UO_937 (O_937,N_24974,N_24435);
and UO_938 (O_938,N_23851,N_24627);
nor UO_939 (O_939,N_24889,N_23829);
and UO_940 (O_940,N_24436,N_24471);
xor UO_941 (O_941,N_24518,N_23961);
or UO_942 (O_942,N_23969,N_24912);
nor UO_943 (O_943,N_24978,N_23853);
nand UO_944 (O_944,N_24562,N_24822);
or UO_945 (O_945,N_24758,N_23860);
and UO_946 (O_946,N_23961,N_24014);
nor UO_947 (O_947,N_24182,N_24847);
and UO_948 (O_948,N_23895,N_23782);
or UO_949 (O_949,N_24093,N_23962);
xor UO_950 (O_950,N_24241,N_23980);
or UO_951 (O_951,N_24278,N_24877);
nor UO_952 (O_952,N_24384,N_23892);
xnor UO_953 (O_953,N_24336,N_24677);
or UO_954 (O_954,N_23837,N_24221);
and UO_955 (O_955,N_24107,N_24321);
nand UO_956 (O_956,N_24599,N_24796);
nand UO_957 (O_957,N_24739,N_24308);
and UO_958 (O_958,N_24947,N_24156);
or UO_959 (O_959,N_24740,N_24755);
and UO_960 (O_960,N_24490,N_24924);
nand UO_961 (O_961,N_24257,N_24602);
or UO_962 (O_962,N_23879,N_24102);
nor UO_963 (O_963,N_24459,N_24460);
nand UO_964 (O_964,N_24999,N_24124);
and UO_965 (O_965,N_24952,N_24198);
and UO_966 (O_966,N_24774,N_23919);
nor UO_967 (O_967,N_23929,N_24786);
nor UO_968 (O_968,N_24492,N_24199);
nor UO_969 (O_969,N_24140,N_24974);
or UO_970 (O_970,N_24497,N_24534);
or UO_971 (O_971,N_24188,N_24786);
or UO_972 (O_972,N_24721,N_24148);
xor UO_973 (O_973,N_24383,N_23796);
or UO_974 (O_974,N_24689,N_24113);
nor UO_975 (O_975,N_24216,N_24951);
and UO_976 (O_976,N_24352,N_24308);
or UO_977 (O_977,N_24222,N_23902);
and UO_978 (O_978,N_23870,N_24407);
nand UO_979 (O_979,N_24780,N_24248);
nand UO_980 (O_980,N_24052,N_24335);
or UO_981 (O_981,N_23975,N_24855);
nand UO_982 (O_982,N_23967,N_24635);
or UO_983 (O_983,N_24425,N_24148);
and UO_984 (O_984,N_23772,N_24238);
and UO_985 (O_985,N_24404,N_23798);
xor UO_986 (O_986,N_24013,N_24750);
nor UO_987 (O_987,N_24919,N_24560);
and UO_988 (O_988,N_24574,N_24873);
or UO_989 (O_989,N_24780,N_24465);
and UO_990 (O_990,N_24031,N_24589);
and UO_991 (O_991,N_23818,N_24369);
and UO_992 (O_992,N_24124,N_24624);
and UO_993 (O_993,N_24719,N_23937);
and UO_994 (O_994,N_23790,N_24918);
xnor UO_995 (O_995,N_24967,N_24137);
xnor UO_996 (O_996,N_24425,N_24233);
and UO_997 (O_997,N_24741,N_24147);
nand UO_998 (O_998,N_24426,N_24558);
or UO_999 (O_999,N_24906,N_23908);
xnor UO_1000 (O_1000,N_23807,N_24092);
or UO_1001 (O_1001,N_24321,N_24813);
xnor UO_1002 (O_1002,N_24591,N_24573);
xnor UO_1003 (O_1003,N_23942,N_23937);
or UO_1004 (O_1004,N_23866,N_24623);
and UO_1005 (O_1005,N_24198,N_24875);
nand UO_1006 (O_1006,N_23950,N_24472);
nand UO_1007 (O_1007,N_23853,N_24999);
nand UO_1008 (O_1008,N_24326,N_24879);
nand UO_1009 (O_1009,N_24496,N_24162);
or UO_1010 (O_1010,N_24319,N_24272);
nand UO_1011 (O_1011,N_24712,N_24730);
or UO_1012 (O_1012,N_24891,N_24790);
and UO_1013 (O_1013,N_24175,N_24042);
or UO_1014 (O_1014,N_23940,N_24460);
xnor UO_1015 (O_1015,N_24186,N_24433);
and UO_1016 (O_1016,N_24640,N_23969);
and UO_1017 (O_1017,N_24415,N_24034);
nand UO_1018 (O_1018,N_24358,N_24580);
nor UO_1019 (O_1019,N_23814,N_24643);
xor UO_1020 (O_1020,N_24487,N_24888);
and UO_1021 (O_1021,N_24770,N_23886);
xnor UO_1022 (O_1022,N_24771,N_24896);
nand UO_1023 (O_1023,N_24963,N_24933);
or UO_1024 (O_1024,N_24322,N_24197);
and UO_1025 (O_1025,N_24957,N_23922);
and UO_1026 (O_1026,N_24270,N_24450);
xnor UO_1027 (O_1027,N_24394,N_24196);
and UO_1028 (O_1028,N_24030,N_24279);
nor UO_1029 (O_1029,N_24675,N_24031);
nor UO_1030 (O_1030,N_24954,N_24495);
or UO_1031 (O_1031,N_24314,N_24524);
or UO_1032 (O_1032,N_24977,N_24217);
nand UO_1033 (O_1033,N_24169,N_24650);
xor UO_1034 (O_1034,N_23774,N_24418);
and UO_1035 (O_1035,N_24452,N_24629);
xnor UO_1036 (O_1036,N_24992,N_23879);
or UO_1037 (O_1037,N_24882,N_23823);
xor UO_1038 (O_1038,N_24437,N_24501);
nand UO_1039 (O_1039,N_24329,N_24223);
nand UO_1040 (O_1040,N_24015,N_24135);
xnor UO_1041 (O_1041,N_24893,N_23969);
xor UO_1042 (O_1042,N_24461,N_24067);
and UO_1043 (O_1043,N_24494,N_23774);
nand UO_1044 (O_1044,N_24412,N_23812);
and UO_1045 (O_1045,N_24118,N_24814);
and UO_1046 (O_1046,N_24812,N_24751);
nor UO_1047 (O_1047,N_23767,N_24390);
and UO_1048 (O_1048,N_24228,N_24362);
nand UO_1049 (O_1049,N_24748,N_24899);
and UO_1050 (O_1050,N_24697,N_23835);
xnor UO_1051 (O_1051,N_24481,N_24672);
nor UO_1052 (O_1052,N_24477,N_24628);
or UO_1053 (O_1053,N_24977,N_23812);
or UO_1054 (O_1054,N_23919,N_24769);
nor UO_1055 (O_1055,N_23899,N_24451);
and UO_1056 (O_1056,N_24564,N_24839);
xnor UO_1057 (O_1057,N_23904,N_24947);
nor UO_1058 (O_1058,N_24109,N_24727);
and UO_1059 (O_1059,N_24933,N_24483);
nand UO_1060 (O_1060,N_24644,N_23865);
and UO_1061 (O_1061,N_23812,N_24408);
and UO_1062 (O_1062,N_23876,N_24612);
and UO_1063 (O_1063,N_24561,N_24222);
nand UO_1064 (O_1064,N_23821,N_24535);
or UO_1065 (O_1065,N_23759,N_23764);
and UO_1066 (O_1066,N_23947,N_24325);
nor UO_1067 (O_1067,N_24057,N_24163);
or UO_1068 (O_1068,N_24021,N_24827);
nand UO_1069 (O_1069,N_23798,N_24534);
and UO_1070 (O_1070,N_24994,N_24154);
nor UO_1071 (O_1071,N_24017,N_24595);
nor UO_1072 (O_1072,N_24402,N_24575);
or UO_1073 (O_1073,N_24754,N_24057);
xnor UO_1074 (O_1074,N_24526,N_24329);
xnor UO_1075 (O_1075,N_24570,N_24671);
nor UO_1076 (O_1076,N_23771,N_24461);
xnor UO_1077 (O_1077,N_24342,N_24257);
or UO_1078 (O_1078,N_24730,N_24464);
nand UO_1079 (O_1079,N_24025,N_24073);
nand UO_1080 (O_1080,N_23862,N_23823);
and UO_1081 (O_1081,N_24432,N_23792);
xor UO_1082 (O_1082,N_24924,N_24867);
xor UO_1083 (O_1083,N_23953,N_24223);
and UO_1084 (O_1084,N_24815,N_24688);
nand UO_1085 (O_1085,N_24459,N_24908);
and UO_1086 (O_1086,N_24862,N_24158);
nand UO_1087 (O_1087,N_23853,N_24313);
or UO_1088 (O_1088,N_23794,N_23755);
or UO_1089 (O_1089,N_24824,N_23843);
nand UO_1090 (O_1090,N_23918,N_24634);
and UO_1091 (O_1091,N_24758,N_24672);
nor UO_1092 (O_1092,N_24658,N_24062);
or UO_1093 (O_1093,N_24599,N_24591);
nand UO_1094 (O_1094,N_23944,N_23804);
or UO_1095 (O_1095,N_24207,N_23774);
and UO_1096 (O_1096,N_24183,N_24578);
xnor UO_1097 (O_1097,N_24352,N_24690);
or UO_1098 (O_1098,N_23932,N_24546);
nor UO_1099 (O_1099,N_24969,N_24077);
nand UO_1100 (O_1100,N_24394,N_24626);
nor UO_1101 (O_1101,N_23807,N_23770);
nand UO_1102 (O_1102,N_24625,N_24866);
or UO_1103 (O_1103,N_24093,N_24352);
nand UO_1104 (O_1104,N_23754,N_24415);
and UO_1105 (O_1105,N_23855,N_24644);
and UO_1106 (O_1106,N_23822,N_24592);
or UO_1107 (O_1107,N_24590,N_23755);
and UO_1108 (O_1108,N_24106,N_24958);
and UO_1109 (O_1109,N_24569,N_24957);
nor UO_1110 (O_1110,N_24909,N_23868);
or UO_1111 (O_1111,N_24387,N_24730);
xnor UO_1112 (O_1112,N_24310,N_24468);
nor UO_1113 (O_1113,N_24862,N_24324);
nand UO_1114 (O_1114,N_23772,N_23789);
or UO_1115 (O_1115,N_24513,N_24637);
xnor UO_1116 (O_1116,N_24236,N_23802);
nor UO_1117 (O_1117,N_24192,N_24223);
nand UO_1118 (O_1118,N_24777,N_24735);
nand UO_1119 (O_1119,N_24948,N_24196);
xor UO_1120 (O_1120,N_24026,N_24529);
or UO_1121 (O_1121,N_24465,N_24995);
or UO_1122 (O_1122,N_23842,N_24406);
xor UO_1123 (O_1123,N_24056,N_23810);
xnor UO_1124 (O_1124,N_24827,N_24024);
nor UO_1125 (O_1125,N_24070,N_24109);
or UO_1126 (O_1126,N_24188,N_23917);
xnor UO_1127 (O_1127,N_24450,N_23891);
nor UO_1128 (O_1128,N_23802,N_24342);
xnor UO_1129 (O_1129,N_24166,N_24252);
nand UO_1130 (O_1130,N_24922,N_24859);
xor UO_1131 (O_1131,N_24236,N_23952);
and UO_1132 (O_1132,N_24413,N_24458);
xor UO_1133 (O_1133,N_24721,N_24357);
nand UO_1134 (O_1134,N_24035,N_24602);
nor UO_1135 (O_1135,N_24054,N_24079);
xor UO_1136 (O_1136,N_24938,N_24905);
nor UO_1137 (O_1137,N_24379,N_24740);
nor UO_1138 (O_1138,N_24617,N_24968);
nand UO_1139 (O_1139,N_23802,N_24241);
nor UO_1140 (O_1140,N_24174,N_24259);
and UO_1141 (O_1141,N_23912,N_24623);
nor UO_1142 (O_1142,N_24868,N_24720);
and UO_1143 (O_1143,N_24962,N_24706);
and UO_1144 (O_1144,N_23982,N_23768);
nor UO_1145 (O_1145,N_23754,N_24812);
nand UO_1146 (O_1146,N_24789,N_24464);
and UO_1147 (O_1147,N_23869,N_24465);
xor UO_1148 (O_1148,N_24138,N_23997);
or UO_1149 (O_1149,N_24302,N_23943);
or UO_1150 (O_1150,N_23893,N_24257);
nor UO_1151 (O_1151,N_24898,N_23770);
and UO_1152 (O_1152,N_24193,N_24587);
xnor UO_1153 (O_1153,N_24323,N_23901);
or UO_1154 (O_1154,N_24128,N_24550);
xor UO_1155 (O_1155,N_23891,N_24581);
or UO_1156 (O_1156,N_24880,N_24528);
and UO_1157 (O_1157,N_24641,N_24858);
nor UO_1158 (O_1158,N_24647,N_23846);
xor UO_1159 (O_1159,N_23900,N_23914);
or UO_1160 (O_1160,N_24545,N_24427);
or UO_1161 (O_1161,N_24997,N_24724);
or UO_1162 (O_1162,N_24194,N_24739);
nor UO_1163 (O_1163,N_23825,N_24830);
xor UO_1164 (O_1164,N_23800,N_24812);
or UO_1165 (O_1165,N_24831,N_23810);
nor UO_1166 (O_1166,N_24060,N_24319);
nand UO_1167 (O_1167,N_24376,N_24545);
nand UO_1168 (O_1168,N_24061,N_23887);
xor UO_1169 (O_1169,N_24691,N_24909);
or UO_1170 (O_1170,N_24793,N_23766);
nor UO_1171 (O_1171,N_24295,N_24234);
xnor UO_1172 (O_1172,N_24618,N_24316);
and UO_1173 (O_1173,N_23961,N_23996);
and UO_1174 (O_1174,N_24493,N_24042);
xor UO_1175 (O_1175,N_24166,N_24664);
and UO_1176 (O_1176,N_24613,N_23944);
xnor UO_1177 (O_1177,N_24244,N_24022);
nand UO_1178 (O_1178,N_24355,N_24533);
nand UO_1179 (O_1179,N_24846,N_24032);
nor UO_1180 (O_1180,N_24972,N_24056);
nor UO_1181 (O_1181,N_23884,N_24306);
or UO_1182 (O_1182,N_23910,N_24434);
and UO_1183 (O_1183,N_23772,N_24673);
nand UO_1184 (O_1184,N_24075,N_23792);
nor UO_1185 (O_1185,N_24463,N_24504);
and UO_1186 (O_1186,N_24909,N_23834);
and UO_1187 (O_1187,N_24204,N_24402);
or UO_1188 (O_1188,N_24193,N_24489);
or UO_1189 (O_1189,N_24036,N_24369);
nor UO_1190 (O_1190,N_23883,N_24135);
nor UO_1191 (O_1191,N_24895,N_24814);
nand UO_1192 (O_1192,N_23895,N_24036);
or UO_1193 (O_1193,N_24028,N_24357);
and UO_1194 (O_1194,N_24459,N_24536);
and UO_1195 (O_1195,N_24280,N_24683);
or UO_1196 (O_1196,N_23842,N_24706);
nand UO_1197 (O_1197,N_24967,N_24944);
and UO_1198 (O_1198,N_24977,N_23882);
or UO_1199 (O_1199,N_24608,N_24375);
xor UO_1200 (O_1200,N_24530,N_24690);
nor UO_1201 (O_1201,N_23995,N_23890);
nor UO_1202 (O_1202,N_23834,N_24789);
and UO_1203 (O_1203,N_24317,N_23891);
or UO_1204 (O_1204,N_24586,N_23778);
and UO_1205 (O_1205,N_24160,N_24091);
nor UO_1206 (O_1206,N_24421,N_24061);
and UO_1207 (O_1207,N_24161,N_24844);
nand UO_1208 (O_1208,N_24661,N_24482);
nor UO_1209 (O_1209,N_24821,N_24170);
nand UO_1210 (O_1210,N_24698,N_23894);
nor UO_1211 (O_1211,N_24552,N_24631);
and UO_1212 (O_1212,N_23874,N_24656);
nor UO_1213 (O_1213,N_24827,N_24437);
nor UO_1214 (O_1214,N_24060,N_24752);
nand UO_1215 (O_1215,N_24523,N_24988);
or UO_1216 (O_1216,N_24310,N_24144);
and UO_1217 (O_1217,N_24537,N_24927);
xnor UO_1218 (O_1218,N_23778,N_24707);
or UO_1219 (O_1219,N_24046,N_24999);
or UO_1220 (O_1220,N_24452,N_24120);
nand UO_1221 (O_1221,N_24514,N_24865);
nor UO_1222 (O_1222,N_24122,N_24126);
nand UO_1223 (O_1223,N_24903,N_24077);
nand UO_1224 (O_1224,N_24578,N_24195);
or UO_1225 (O_1225,N_24563,N_24404);
nor UO_1226 (O_1226,N_24719,N_24929);
nand UO_1227 (O_1227,N_24688,N_23890);
nand UO_1228 (O_1228,N_24771,N_24832);
nand UO_1229 (O_1229,N_23935,N_24172);
nand UO_1230 (O_1230,N_24840,N_24298);
xnor UO_1231 (O_1231,N_23969,N_23835);
and UO_1232 (O_1232,N_24701,N_24499);
nand UO_1233 (O_1233,N_24572,N_23794);
or UO_1234 (O_1234,N_24885,N_24661);
and UO_1235 (O_1235,N_23884,N_24090);
nor UO_1236 (O_1236,N_24017,N_24584);
nor UO_1237 (O_1237,N_24080,N_24909);
nand UO_1238 (O_1238,N_24039,N_24736);
or UO_1239 (O_1239,N_23825,N_24343);
xor UO_1240 (O_1240,N_24612,N_24966);
nand UO_1241 (O_1241,N_23912,N_24982);
nor UO_1242 (O_1242,N_24281,N_24538);
or UO_1243 (O_1243,N_23958,N_23798);
nor UO_1244 (O_1244,N_23932,N_23836);
or UO_1245 (O_1245,N_23864,N_24537);
and UO_1246 (O_1246,N_24187,N_24176);
xnor UO_1247 (O_1247,N_24011,N_24491);
and UO_1248 (O_1248,N_24786,N_23844);
nand UO_1249 (O_1249,N_23840,N_23871);
and UO_1250 (O_1250,N_24995,N_24941);
nor UO_1251 (O_1251,N_23865,N_23955);
or UO_1252 (O_1252,N_24496,N_23901);
or UO_1253 (O_1253,N_23798,N_24472);
or UO_1254 (O_1254,N_24670,N_23935);
xor UO_1255 (O_1255,N_24062,N_24554);
or UO_1256 (O_1256,N_23966,N_24745);
xor UO_1257 (O_1257,N_24981,N_24294);
nand UO_1258 (O_1258,N_24215,N_24899);
or UO_1259 (O_1259,N_24798,N_24639);
xor UO_1260 (O_1260,N_24102,N_23913);
nor UO_1261 (O_1261,N_23925,N_23902);
or UO_1262 (O_1262,N_24815,N_24028);
and UO_1263 (O_1263,N_23861,N_24709);
nor UO_1264 (O_1264,N_23955,N_24366);
xor UO_1265 (O_1265,N_24621,N_23760);
or UO_1266 (O_1266,N_23994,N_23788);
nor UO_1267 (O_1267,N_24187,N_24297);
nand UO_1268 (O_1268,N_23852,N_23819);
xor UO_1269 (O_1269,N_24186,N_24059);
and UO_1270 (O_1270,N_24648,N_24432);
nor UO_1271 (O_1271,N_23821,N_23765);
nand UO_1272 (O_1272,N_24596,N_23838);
or UO_1273 (O_1273,N_24092,N_24038);
nand UO_1274 (O_1274,N_24530,N_24445);
or UO_1275 (O_1275,N_23876,N_24115);
nor UO_1276 (O_1276,N_24322,N_23931);
nor UO_1277 (O_1277,N_23766,N_24203);
and UO_1278 (O_1278,N_24224,N_24955);
nor UO_1279 (O_1279,N_23942,N_23874);
xnor UO_1280 (O_1280,N_24046,N_24401);
and UO_1281 (O_1281,N_24270,N_23862);
nand UO_1282 (O_1282,N_24517,N_24813);
nand UO_1283 (O_1283,N_24017,N_23893);
xor UO_1284 (O_1284,N_23925,N_24272);
nand UO_1285 (O_1285,N_24630,N_24098);
nor UO_1286 (O_1286,N_24642,N_24389);
nand UO_1287 (O_1287,N_24091,N_23851);
xor UO_1288 (O_1288,N_23803,N_24303);
or UO_1289 (O_1289,N_24512,N_24559);
xnor UO_1290 (O_1290,N_24412,N_23803);
or UO_1291 (O_1291,N_24776,N_24189);
or UO_1292 (O_1292,N_24782,N_24533);
xnor UO_1293 (O_1293,N_24800,N_24697);
nand UO_1294 (O_1294,N_24072,N_24624);
nand UO_1295 (O_1295,N_23968,N_23754);
nor UO_1296 (O_1296,N_24052,N_24463);
nor UO_1297 (O_1297,N_24041,N_24477);
or UO_1298 (O_1298,N_24741,N_24334);
xor UO_1299 (O_1299,N_24052,N_24275);
xnor UO_1300 (O_1300,N_23753,N_24467);
nor UO_1301 (O_1301,N_24165,N_24899);
nor UO_1302 (O_1302,N_24015,N_23764);
and UO_1303 (O_1303,N_24531,N_24831);
nor UO_1304 (O_1304,N_24886,N_24993);
or UO_1305 (O_1305,N_24360,N_24482);
or UO_1306 (O_1306,N_24301,N_24552);
nor UO_1307 (O_1307,N_24180,N_24861);
nand UO_1308 (O_1308,N_23804,N_24875);
or UO_1309 (O_1309,N_24867,N_24285);
and UO_1310 (O_1310,N_23894,N_24190);
nor UO_1311 (O_1311,N_24431,N_23815);
nand UO_1312 (O_1312,N_24247,N_24139);
nor UO_1313 (O_1313,N_24229,N_24841);
nand UO_1314 (O_1314,N_24208,N_24295);
nand UO_1315 (O_1315,N_24945,N_24434);
xor UO_1316 (O_1316,N_23872,N_23899);
and UO_1317 (O_1317,N_24236,N_24764);
nand UO_1318 (O_1318,N_24957,N_24130);
or UO_1319 (O_1319,N_24239,N_24968);
nand UO_1320 (O_1320,N_24053,N_24366);
nor UO_1321 (O_1321,N_24290,N_24380);
and UO_1322 (O_1322,N_24324,N_24215);
nor UO_1323 (O_1323,N_24384,N_24859);
xor UO_1324 (O_1324,N_23861,N_23956);
and UO_1325 (O_1325,N_24153,N_24618);
nand UO_1326 (O_1326,N_24920,N_24753);
nand UO_1327 (O_1327,N_23991,N_24523);
xnor UO_1328 (O_1328,N_23881,N_23963);
xor UO_1329 (O_1329,N_24018,N_24055);
nor UO_1330 (O_1330,N_24692,N_24093);
nor UO_1331 (O_1331,N_24039,N_24210);
xnor UO_1332 (O_1332,N_24146,N_23823);
nand UO_1333 (O_1333,N_24560,N_24211);
nand UO_1334 (O_1334,N_23902,N_24671);
or UO_1335 (O_1335,N_24233,N_24807);
or UO_1336 (O_1336,N_24798,N_24818);
and UO_1337 (O_1337,N_24659,N_24285);
and UO_1338 (O_1338,N_24355,N_23842);
nor UO_1339 (O_1339,N_24902,N_24444);
nor UO_1340 (O_1340,N_24911,N_23891);
xnor UO_1341 (O_1341,N_24477,N_24525);
nor UO_1342 (O_1342,N_24012,N_24972);
and UO_1343 (O_1343,N_24783,N_24149);
nor UO_1344 (O_1344,N_24196,N_24313);
or UO_1345 (O_1345,N_23906,N_24610);
and UO_1346 (O_1346,N_24298,N_24382);
nor UO_1347 (O_1347,N_23849,N_24986);
nand UO_1348 (O_1348,N_24743,N_24915);
xor UO_1349 (O_1349,N_23998,N_24806);
nor UO_1350 (O_1350,N_24044,N_24713);
nand UO_1351 (O_1351,N_24833,N_24452);
nand UO_1352 (O_1352,N_24084,N_24634);
or UO_1353 (O_1353,N_24443,N_24899);
and UO_1354 (O_1354,N_24578,N_24444);
or UO_1355 (O_1355,N_23891,N_24580);
nand UO_1356 (O_1356,N_24483,N_24340);
nand UO_1357 (O_1357,N_24655,N_24103);
and UO_1358 (O_1358,N_24503,N_24103);
nand UO_1359 (O_1359,N_24593,N_24780);
nand UO_1360 (O_1360,N_24017,N_24727);
xnor UO_1361 (O_1361,N_23960,N_24812);
xnor UO_1362 (O_1362,N_24162,N_24303);
or UO_1363 (O_1363,N_24627,N_24016);
or UO_1364 (O_1364,N_24753,N_24081);
and UO_1365 (O_1365,N_24921,N_24698);
and UO_1366 (O_1366,N_23787,N_24493);
nand UO_1367 (O_1367,N_24869,N_24426);
and UO_1368 (O_1368,N_24761,N_24565);
nor UO_1369 (O_1369,N_24827,N_23919);
and UO_1370 (O_1370,N_23896,N_24158);
and UO_1371 (O_1371,N_23954,N_24323);
nor UO_1372 (O_1372,N_24795,N_24598);
xnor UO_1373 (O_1373,N_24069,N_24431);
nor UO_1374 (O_1374,N_24426,N_24575);
xor UO_1375 (O_1375,N_23760,N_24783);
xnor UO_1376 (O_1376,N_24636,N_23825);
or UO_1377 (O_1377,N_24582,N_24307);
nor UO_1378 (O_1378,N_24422,N_24781);
or UO_1379 (O_1379,N_24218,N_24814);
and UO_1380 (O_1380,N_24803,N_24403);
and UO_1381 (O_1381,N_24277,N_24107);
xor UO_1382 (O_1382,N_23780,N_24420);
nor UO_1383 (O_1383,N_24814,N_24046);
nor UO_1384 (O_1384,N_23841,N_24502);
and UO_1385 (O_1385,N_24500,N_24634);
xor UO_1386 (O_1386,N_24186,N_23892);
and UO_1387 (O_1387,N_24337,N_24049);
xor UO_1388 (O_1388,N_24091,N_24322);
nor UO_1389 (O_1389,N_24738,N_24713);
and UO_1390 (O_1390,N_24600,N_24478);
nor UO_1391 (O_1391,N_24583,N_24794);
nand UO_1392 (O_1392,N_24436,N_23928);
nor UO_1393 (O_1393,N_24331,N_23874);
and UO_1394 (O_1394,N_24455,N_24949);
or UO_1395 (O_1395,N_23890,N_24725);
or UO_1396 (O_1396,N_24856,N_24912);
or UO_1397 (O_1397,N_24281,N_24455);
nor UO_1398 (O_1398,N_24236,N_24650);
nand UO_1399 (O_1399,N_24006,N_24619);
nand UO_1400 (O_1400,N_24217,N_24429);
nand UO_1401 (O_1401,N_23757,N_24682);
nor UO_1402 (O_1402,N_24169,N_24818);
xnor UO_1403 (O_1403,N_24573,N_23981);
or UO_1404 (O_1404,N_24643,N_24162);
or UO_1405 (O_1405,N_24478,N_23803);
or UO_1406 (O_1406,N_24031,N_24922);
xor UO_1407 (O_1407,N_24685,N_24383);
or UO_1408 (O_1408,N_24729,N_24878);
nor UO_1409 (O_1409,N_24688,N_24431);
nand UO_1410 (O_1410,N_23891,N_23802);
nand UO_1411 (O_1411,N_24401,N_23822);
xor UO_1412 (O_1412,N_24689,N_24218);
xor UO_1413 (O_1413,N_24163,N_24591);
xor UO_1414 (O_1414,N_23896,N_24036);
nand UO_1415 (O_1415,N_24977,N_24024);
nand UO_1416 (O_1416,N_24999,N_24804);
and UO_1417 (O_1417,N_23975,N_24621);
and UO_1418 (O_1418,N_24452,N_24596);
xnor UO_1419 (O_1419,N_23831,N_23977);
or UO_1420 (O_1420,N_24704,N_24339);
xor UO_1421 (O_1421,N_24526,N_24501);
or UO_1422 (O_1422,N_24539,N_24468);
nand UO_1423 (O_1423,N_23799,N_24701);
xnor UO_1424 (O_1424,N_24812,N_24188);
xor UO_1425 (O_1425,N_23882,N_24537);
xnor UO_1426 (O_1426,N_24318,N_24747);
nand UO_1427 (O_1427,N_24003,N_24915);
and UO_1428 (O_1428,N_24464,N_24386);
xnor UO_1429 (O_1429,N_24260,N_24195);
xor UO_1430 (O_1430,N_24633,N_24162);
xnor UO_1431 (O_1431,N_24466,N_24037);
and UO_1432 (O_1432,N_24300,N_24682);
nand UO_1433 (O_1433,N_24284,N_23929);
nand UO_1434 (O_1434,N_24229,N_24210);
xnor UO_1435 (O_1435,N_24065,N_24506);
or UO_1436 (O_1436,N_24449,N_24891);
nor UO_1437 (O_1437,N_24253,N_23892);
nand UO_1438 (O_1438,N_24841,N_23952);
nor UO_1439 (O_1439,N_24030,N_24538);
xnor UO_1440 (O_1440,N_24850,N_23811);
nor UO_1441 (O_1441,N_24706,N_24496);
nand UO_1442 (O_1442,N_23931,N_24258);
nor UO_1443 (O_1443,N_24772,N_24892);
nor UO_1444 (O_1444,N_24977,N_24378);
and UO_1445 (O_1445,N_24653,N_24816);
and UO_1446 (O_1446,N_24403,N_24279);
xor UO_1447 (O_1447,N_24902,N_24084);
nor UO_1448 (O_1448,N_23963,N_24213);
and UO_1449 (O_1449,N_24651,N_24704);
nand UO_1450 (O_1450,N_24748,N_24389);
nor UO_1451 (O_1451,N_24366,N_23822);
and UO_1452 (O_1452,N_24961,N_24859);
nand UO_1453 (O_1453,N_24095,N_24990);
nor UO_1454 (O_1454,N_24456,N_24545);
nor UO_1455 (O_1455,N_24428,N_23867);
xnor UO_1456 (O_1456,N_24428,N_24274);
nand UO_1457 (O_1457,N_24842,N_24777);
xor UO_1458 (O_1458,N_24912,N_24210);
xor UO_1459 (O_1459,N_24430,N_24563);
and UO_1460 (O_1460,N_24259,N_23814);
or UO_1461 (O_1461,N_24787,N_24615);
nand UO_1462 (O_1462,N_24148,N_24008);
and UO_1463 (O_1463,N_24713,N_24986);
nor UO_1464 (O_1464,N_23949,N_24264);
or UO_1465 (O_1465,N_23812,N_23750);
and UO_1466 (O_1466,N_24940,N_24843);
or UO_1467 (O_1467,N_23802,N_24415);
and UO_1468 (O_1468,N_23984,N_24662);
nor UO_1469 (O_1469,N_24497,N_24340);
or UO_1470 (O_1470,N_24379,N_24714);
nand UO_1471 (O_1471,N_24753,N_24543);
or UO_1472 (O_1472,N_23840,N_23760);
and UO_1473 (O_1473,N_24652,N_24392);
nor UO_1474 (O_1474,N_23856,N_24105);
nor UO_1475 (O_1475,N_24552,N_24759);
xnor UO_1476 (O_1476,N_24417,N_23952);
or UO_1477 (O_1477,N_24318,N_24180);
nand UO_1478 (O_1478,N_24556,N_23871);
nand UO_1479 (O_1479,N_24393,N_24289);
nor UO_1480 (O_1480,N_24480,N_24943);
xor UO_1481 (O_1481,N_24553,N_24646);
xor UO_1482 (O_1482,N_24687,N_23795);
nor UO_1483 (O_1483,N_24561,N_24775);
nand UO_1484 (O_1484,N_24546,N_24535);
or UO_1485 (O_1485,N_23824,N_23943);
nor UO_1486 (O_1486,N_24102,N_23884);
nand UO_1487 (O_1487,N_24364,N_24933);
xnor UO_1488 (O_1488,N_24563,N_23891);
and UO_1489 (O_1489,N_24127,N_24816);
and UO_1490 (O_1490,N_23770,N_24377);
xor UO_1491 (O_1491,N_24282,N_24684);
or UO_1492 (O_1492,N_24228,N_24663);
nand UO_1493 (O_1493,N_24792,N_23886);
xor UO_1494 (O_1494,N_24996,N_24463);
xnor UO_1495 (O_1495,N_24412,N_24770);
nor UO_1496 (O_1496,N_24137,N_23925);
and UO_1497 (O_1497,N_23918,N_24496);
and UO_1498 (O_1498,N_23874,N_24228);
or UO_1499 (O_1499,N_24761,N_24110);
nand UO_1500 (O_1500,N_24933,N_24430);
xnor UO_1501 (O_1501,N_23797,N_24003);
nand UO_1502 (O_1502,N_24239,N_24335);
and UO_1503 (O_1503,N_23826,N_24492);
or UO_1504 (O_1504,N_24860,N_24006);
nand UO_1505 (O_1505,N_24258,N_24981);
nand UO_1506 (O_1506,N_24538,N_23977);
nand UO_1507 (O_1507,N_23875,N_24338);
nor UO_1508 (O_1508,N_24252,N_24940);
nand UO_1509 (O_1509,N_24926,N_24781);
nand UO_1510 (O_1510,N_23950,N_24317);
nor UO_1511 (O_1511,N_24796,N_23947);
xnor UO_1512 (O_1512,N_24249,N_23858);
nand UO_1513 (O_1513,N_24033,N_24887);
and UO_1514 (O_1514,N_24894,N_24328);
nor UO_1515 (O_1515,N_24294,N_24385);
and UO_1516 (O_1516,N_24818,N_24180);
and UO_1517 (O_1517,N_24097,N_24745);
nand UO_1518 (O_1518,N_24903,N_23806);
nand UO_1519 (O_1519,N_24674,N_24454);
and UO_1520 (O_1520,N_24986,N_24975);
or UO_1521 (O_1521,N_23975,N_24337);
or UO_1522 (O_1522,N_24786,N_24503);
nor UO_1523 (O_1523,N_24082,N_23994);
and UO_1524 (O_1524,N_23771,N_24341);
xnor UO_1525 (O_1525,N_24877,N_24759);
and UO_1526 (O_1526,N_24276,N_23877);
nand UO_1527 (O_1527,N_24759,N_24397);
xnor UO_1528 (O_1528,N_24525,N_24834);
and UO_1529 (O_1529,N_24117,N_23789);
or UO_1530 (O_1530,N_24816,N_24021);
nor UO_1531 (O_1531,N_24316,N_24759);
and UO_1532 (O_1532,N_24930,N_23929);
and UO_1533 (O_1533,N_23900,N_24919);
nor UO_1534 (O_1534,N_24046,N_23981);
nand UO_1535 (O_1535,N_24895,N_24955);
nand UO_1536 (O_1536,N_24417,N_24774);
nor UO_1537 (O_1537,N_23895,N_23790);
nand UO_1538 (O_1538,N_23886,N_24663);
nor UO_1539 (O_1539,N_23793,N_24624);
or UO_1540 (O_1540,N_24522,N_24041);
and UO_1541 (O_1541,N_24584,N_24293);
and UO_1542 (O_1542,N_24044,N_23844);
and UO_1543 (O_1543,N_24885,N_24733);
xnor UO_1544 (O_1544,N_23896,N_24807);
nor UO_1545 (O_1545,N_24789,N_24466);
nor UO_1546 (O_1546,N_24713,N_24015);
and UO_1547 (O_1547,N_24401,N_24047);
nand UO_1548 (O_1548,N_24656,N_24817);
nand UO_1549 (O_1549,N_24103,N_24665);
or UO_1550 (O_1550,N_24694,N_23758);
nand UO_1551 (O_1551,N_23881,N_23832);
or UO_1552 (O_1552,N_24072,N_24040);
or UO_1553 (O_1553,N_24017,N_23865);
or UO_1554 (O_1554,N_24317,N_23810);
and UO_1555 (O_1555,N_24948,N_24602);
nand UO_1556 (O_1556,N_24930,N_23986);
xnor UO_1557 (O_1557,N_24229,N_24460);
xor UO_1558 (O_1558,N_23820,N_24260);
nand UO_1559 (O_1559,N_24425,N_24448);
xor UO_1560 (O_1560,N_24837,N_24660);
nand UO_1561 (O_1561,N_24599,N_24340);
or UO_1562 (O_1562,N_23846,N_24604);
nor UO_1563 (O_1563,N_24743,N_24170);
and UO_1564 (O_1564,N_23776,N_24428);
xnor UO_1565 (O_1565,N_23758,N_23955);
xnor UO_1566 (O_1566,N_24237,N_23968);
or UO_1567 (O_1567,N_24250,N_24023);
nand UO_1568 (O_1568,N_24652,N_23966);
or UO_1569 (O_1569,N_23824,N_24332);
xnor UO_1570 (O_1570,N_24283,N_23860);
nand UO_1571 (O_1571,N_24065,N_24501);
nor UO_1572 (O_1572,N_23892,N_23886);
nor UO_1573 (O_1573,N_24886,N_24125);
or UO_1574 (O_1574,N_24880,N_24630);
nor UO_1575 (O_1575,N_24723,N_24758);
and UO_1576 (O_1576,N_23761,N_24365);
nor UO_1577 (O_1577,N_24958,N_24616);
xnor UO_1578 (O_1578,N_24446,N_24463);
xnor UO_1579 (O_1579,N_24172,N_24540);
nand UO_1580 (O_1580,N_24183,N_24340);
and UO_1581 (O_1581,N_24575,N_23812);
and UO_1582 (O_1582,N_24805,N_24108);
xnor UO_1583 (O_1583,N_23861,N_24839);
and UO_1584 (O_1584,N_24693,N_24073);
and UO_1585 (O_1585,N_23947,N_24707);
xor UO_1586 (O_1586,N_23751,N_24690);
and UO_1587 (O_1587,N_23763,N_24038);
or UO_1588 (O_1588,N_24721,N_23769);
xor UO_1589 (O_1589,N_24754,N_24969);
or UO_1590 (O_1590,N_24403,N_24972);
or UO_1591 (O_1591,N_24468,N_24926);
and UO_1592 (O_1592,N_23794,N_24973);
nand UO_1593 (O_1593,N_24007,N_23759);
nor UO_1594 (O_1594,N_24175,N_23780);
xnor UO_1595 (O_1595,N_24830,N_24472);
nand UO_1596 (O_1596,N_24599,N_24823);
or UO_1597 (O_1597,N_24373,N_24275);
and UO_1598 (O_1598,N_24385,N_24451);
or UO_1599 (O_1599,N_24586,N_24442);
nor UO_1600 (O_1600,N_23829,N_23953);
xor UO_1601 (O_1601,N_23911,N_24202);
nand UO_1602 (O_1602,N_23759,N_24466);
xor UO_1603 (O_1603,N_24239,N_23984);
and UO_1604 (O_1604,N_23992,N_24562);
and UO_1605 (O_1605,N_24049,N_24863);
nand UO_1606 (O_1606,N_24746,N_24522);
nor UO_1607 (O_1607,N_24765,N_24060);
nor UO_1608 (O_1608,N_24726,N_24959);
xnor UO_1609 (O_1609,N_23883,N_24279);
or UO_1610 (O_1610,N_24855,N_24635);
or UO_1611 (O_1611,N_23793,N_24970);
and UO_1612 (O_1612,N_24613,N_24699);
or UO_1613 (O_1613,N_24385,N_24474);
nand UO_1614 (O_1614,N_24807,N_24273);
and UO_1615 (O_1615,N_24696,N_24711);
or UO_1616 (O_1616,N_24864,N_24627);
or UO_1617 (O_1617,N_24566,N_24241);
or UO_1618 (O_1618,N_24782,N_23811);
and UO_1619 (O_1619,N_24246,N_24430);
xor UO_1620 (O_1620,N_24724,N_24468);
nor UO_1621 (O_1621,N_23993,N_24695);
or UO_1622 (O_1622,N_23944,N_24154);
nor UO_1623 (O_1623,N_23958,N_24479);
and UO_1624 (O_1624,N_24765,N_24940);
or UO_1625 (O_1625,N_24759,N_24851);
nor UO_1626 (O_1626,N_23832,N_23904);
or UO_1627 (O_1627,N_24445,N_23811);
and UO_1628 (O_1628,N_23879,N_24794);
or UO_1629 (O_1629,N_23771,N_24654);
and UO_1630 (O_1630,N_23934,N_24712);
xnor UO_1631 (O_1631,N_24699,N_24826);
and UO_1632 (O_1632,N_24959,N_24264);
xor UO_1633 (O_1633,N_24489,N_23770);
or UO_1634 (O_1634,N_24222,N_24463);
xnor UO_1635 (O_1635,N_23803,N_24794);
or UO_1636 (O_1636,N_24933,N_24744);
or UO_1637 (O_1637,N_24482,N_23765);
nand UO_1638 (O_1638,N_24655,N_24333);
xor UO_1639 (O_1639,N_24914,N_23973);
nand UO_1640 (O_1640,N_23882,N_23832);
xor UO_1641 (O_1641,N_24077,N_24622);
nor UO_1642 (O_1642,N_23754,N_24367);
xor UO_1643 (O_1643,N_24226,N_24408);
nand UO_1644 (O_1644,N_24947,N_24391);
or UO_1645 (O_1645,N_24671,N_24864);
or UO_1646 (O_1646,N_24222,N_24545);
nand UO_1647 (O_1647,N_23880,N_24518);
or UO_1648 (O_1648,N_24433,N_24779);
nand UO_1649 (O_1649,N_23864,N_24318);
xor UO_1650 (O_1650,N_24099,N_24500);
nand UO_1651 (O_1651,N_24910,N_23986);
and UO_1652 (O_1652,N_24459,N_24091);
xor UO_1653 (O_1653,N_24812,N_24358);
nand UO_1654 (O_1654,N_23963,N_24545);
nand UO_1655 (O_1655,N_24527,N_23805);
nand UO_1656 (O_1656,N_24853,N_24863);
and UO_1657 (O_1657,N_24033,N_24838);
and UO_1658 (O_1658,N_24767,N_23765);
or UO_1659 (O_1659,N_24105,N_23931);
nand UO_1660 (O_1660,N_24286,N_24114);
nor UO_1661 (O_1661,N_24067,N_24623);
xnor UO_1662 (O_1662,N_23911,N_24385);
and UO_1663 (O_1663,N_24591,N_24153);
nor UO_1664 (O_1664,N_24099,N_23854);
or UO_1665 (O_1665,N_23997,N_24618);
xor UO_1666 (O_1666,N_24004,N_24986);
and UO_1667 (O_1667,N_24039,N_24845);
nand UO_1668 (O_1668,N_24799,N_24015);
xnor UO_1669 (O_1669,N_24154,N_24656);
or UO_1670 (O_1670,N_23958,N_24049);
xor UO_1671 (O_1671,N_24256,N_23975);
nor UO_1672 (O_1672,N_24981,N_24863);
nor UO_1673 (O_1673,N_24135,N_24235);
nor UO_1674 (O_1674,N_24936,N_24578);
nor UO_1675 (O_1675,N_24342,N_24239);
and UO_1676 (O_1676,N_24477,N_24150);
nor UO_1677 (O_1677,N_24713,N_24519);
or UO_1678 (O_1678,N_23880,N_24266);
nand UO_1679 (O_1679,N_24470,N_24250);
nor UO_1680 (O_1680,N_24910,N_23934);
or UO_1681 (O_1681,N_24818,N_24381);
or UO_1682 (O_1682,N_23931,N_24845);
and UO_1683 (O_1683,N_24662,N_24506);
xnor UO_1684 (O_1684,N_24577,N_23879);
and UO_1685 (O_1685,N_24846,N_24002);
nor UO_1686 (O_1686,N_24465,N_24901);
xnor UO_1687 (O_1687,N_24862,N_23768);
xnor UO_1688 (O_1688,N_24941,N_24619);
xnor UO_1689 (O_1689,N_24129,N_23782);
nor UO_1690 (O_1690,N_23861,N_24489);
and UO_1691 (O_1691,N_24051,N_24284);
xnor UO_1692 (O_1692,N_23926,N_24690);
nor UO_1693 (O_1693,N_23885,N_24504);
and UO_1694 (O_1694,N_24608,N_24644);
nor UO_1695 (O_1695,N_24742,N_23795);
nor UO_1696 (O_1696,N_24223,N_24919);
xor UO_1697 (O_1697,N_24152,N_24952);
and UO_1698 (O_1698,N_23761,N_23799);
or UO_1699 (O_1699,N_23904,N_24486);
and UO_1700 (O_1700,N_24928,N_23829);
xnor UO_1701 (O_1701,N_24517,N_24569);
or UO_1702 (O_1702,N_24927,N_24337);
xor UO_1703 (O_1703,N_23979,N_24511);
nand UO_1704 (O_1704,N_23982,N_23893);
xnor UO_1705 (O_1705,N_24086,N_24638);
nor UO_1706 (O_1706,N_23865,N_24973);
nand UO_1707 (O_1707,N_23848,N_24576);
or UO_1708 (O_1708,N_24227,N_24697);
nor UO_1709 (O_1709,N_24086,N_24761);
nor UO_1710 (O_1710,N_23825,N_24486);
and UO_1711 (O_1711,N_23784,N_24440);
and UO_1712 (O_1712,N_24953,N_24886);
or UO_1713 (O_1713,N_24490,N_24085);
and UO_1714 (O_1714,N_24145,N_24422);
or UO_1715 (O_1715,N_24724,N_24172);
or UO_1716 (O_1716,N_24302,N_24364);
or UO_1717 (O_1717,N_24382,N_24544);
xor UO_1718 (O_1718,N_24806,N_23937);
and UO_1719 (O_1719,N_24313,N_24460);
or UO_1720 (O_1720,N_24148,N_23955);
nand UO_1721 (O_1721,N_24351,N_24875);
xnor UO_1722 (O_1722,N_24269,N_23889);
nand UO_1723 (O_1723,N_24300,N_23887);
and UO_1724 (O_1724,N_23868,N_23953);
or UO_1725 (O_1725,N_24391,N_23801);
and UO_1726 (O_1726,N_24818,N_23796);
nor UO_1727 (O_1727,N_24173,N_24273);
nand UO_1728 (O_1728,N_24139,N_23995);
nor UO_1729 (O_1729,N_23901,N_24681);
nor UO_1730 (O_1730,N_24429,N_24151);
xnor UO_1731 (O_1731,N_24232,N_24719);
and UO_1732 (O_1732,N_24449,N_24308);
or UO_1733 (O_1733,N_24929,N_24326);
nor UO_1734 (O_1734,N_24220,N_24250);
or UO_1735 (O_1735,N_23857,N_23806);
and UO_1736 (O_1736,N_24422,N_24976);
and UO_1737 (O_1737,N_24638,N_24088);
nor UO_1738 (O_1738,N_24167,N_24377);
xor UO_1739 (O_1739,N_24869,N_24990);
or UO_1740 (O_1740,N_24629,N_24969);
nor UO_1741 (O_1741,N_24821,N_24348);
nand UO_1742 (O_1742,N_24836,N_24125);
and UO_1743 (O_1743,N_24238,N_24083);
or UO_1744 (O_1744,N_24676,N_24228);
nand UO_1745 (O_1745,N_24261,N_24980);
and UO_1746 (O_1746,N_24063,N_24529);
nor UO_1747 (O_1747,N_24833,N_24752);
and UO_1748 (O_1748,N_24747,N_24023);
and UO_1749 (O_1749,N_24110,N_24861);
xor UO_1750 (O_1750,N_24708,N_24432);
nand UO_1751 (O_1751,N_23786,N_23886);
or UO_1752 (O_1752,N_24177,N_24602);
xor UO_1753 (O_1753,N_23961,N_24448);
nand UO_1754 (O_1754,N_24177,N_23961);
xnor UO_1755 (O_1755,N_24688,N_23874);
xor UO_1756 (O_1756,N_23775,N_24543);
nor UO_1757 (O_1757,N_23792,N_24517);
nand UO_1758 (O_1758,N_24748,N_24939);
xor UO_1759 (O_1759,N_24473,N_24681);
xnor UO_1760 (O_1760,N_24444,N_23933);
or UO_1761 (O_1761,N_24221,N_24540);
nor UO_1762 (O_1762,N_24395,N_24757);
nor UO_1763 (O_1763,N_23785,N_24053);
and UO_1764 (O_1764,N_24971,N_24817);
and UO_1765 (O_1765,N_24424,N_23810);
xnor UO_1766 (O_1766,N_23786,N_24809);
and UO_1767 (O_1767,N_24699,N_23838);
or UO_1768 (O_1768,N_23854,N_24450);
or UO_1769 (O_1769,N_24966,N_24548);
or UO_1770 (O_1770,N_24159,N_24156);
and UO_1771 (O_1771,N_24235,N_24383);
nand UO_1772 (O_1772,N_24825,N_23799);
nand UO_1773 (O_1773,N_23754,N_24648);
or UO_1774 (O_1774,N_24032,N_24784);
or UO_1775 (O_1775,N_24934,N_24118);
and UO_1776 (O_1776,N_24463,N_24510);
xor UO_1777 (O_1777,N_24873,N_24246);
nor UO_1778 (O_1778,N_24461,N_24715);
and UO_1779 (O_1779,N_24516,N_23903);
and UO_1780 (O_1780,N_24434,N_24753);
nor UO_1781 (O_1781,N_24674,N_24135);
nor UO_1782 (O_1782,N_24484,N_24014);
or UO_1783 (O_1783,N_24975,N_24930);
nor UO_1784 (O_1784,N_23762,N_24929);
or UO_1785 (O_1785,N_24732,N_24470);
and UO_1786 (O_1786,N_24012,N_24879);
nor UO_1787 (O_1787,N_24031,N_24471);
xnor UO_1788 (O_1788,N_24865,N_24863);
nor UO_1789 (O_1789,N_23848,N_24516);
nor UO_1790 (O_1790,N_24153,N_24175);
xnor UO_1791 (O_1791,N_24758,N_24981);
xnor UO_1792 (O_1792,N_24727,N_24535);
and UO_1793 (O_1793,N_24662,N_24056);
nand UO_1794 (O_1794,N_24152,N_24420);
and UO_1795 (O_1795,N_24613,N_24639);
and UO_1796 (O_1796,N_23793,N_24375);
xor UO_1797 (O_1797,N_24623,N_24905);
nand UO_1798 (O_1798,N_24058,N_23843);
or UO_1799 (O_1799,N_24224,N_24032);
and UO_1800 (O_1800,N_24271,N_24706);
and UO_1801 (O_1801,N_24461,N_23967);
xor UO_1802 (O_1802,N_23752,N_24945);
and UO_1803 (O_1803,N_24470,N_24138);
nand UO_1804 (O_1804,N_24239,N_24901);
and UO_1805 (O_1805,N_23797,N_24933);
or UO_1806 (O_1806,N_23940,N_24692);
nand UO_1807 (O_1807,N_23858,N_24382);
and UO_1808 (O_1808,N_24913,N_24427);
nor UO_1809 (O_1809,N_24201,N_24992);
and UO_1810 (O_1810,N_24023,N_24537);
nor UO_1811 (O_1811,N_24803,N_24139);
nor UO_1812 (O_1812,N_24092,N_24423);
or UO_1813 (O_1813,N_24604,N_24905);
nor UO_1814 (O_1814,N_24365,N_24772);
nor UO_1815 (O_1815,N_24134,N_23770);
or UO_1816 (O_1816,N_23974,N_24422);
nor UO_1817 (O_1817,N_24440,N_24404);
nand UO_1818 (O_1818,N_24116,N_24764);
nor UO_1819 (O_1819,N_24771,N_24395);
nor UO_1820 (O_1820,N_23953,N_24221);
or UO_1821 (O_1821,N_24076,N_24172);
nor UO_1822 (O_1822,N_24397,N_24964);
nor UO_1823 (O_1823,N_23824,N_24512);
nor UO_1824 (O_1824,N_24688,N_24598);
nor UO_1825 (O_1825,N_24688,N_24653);
nand UO_1826 (O_1826,N_24501,N_24538);
xnor UO_1827 (O_1827,N_24770,N_24565);
or UO_1828 (O_1828,N_23812,N_24537);
and UO_1829 (O_1829,N_24506,N_24280);
and UO_1830 (O_1830,N_24713,N_24817);
xnor UO_1831 (O_1831,N_24392,N_24251);
or UO_1832 (O_1832,N_24595,N_24290);
nand UO_1833 (O_1833,N_24109,N_24346);
nor UO_1834 (O_1834,N_24347,N_24406);
and UO_1835 (O_1835,N_23784,N_24616);
nand UO_1836 (O_1836,N_24127,N_24357);
and UO_1837 (O_1837,N_24961,N_24127);
and UO_1838 (O_1838,N_24408,N_23862);
xor UO_1839 (O_1839,N_23788,N_24716);
and UO_1840 (O_1840,N_24943,N_24416);
nor UO_1841 (O_1841,N_24026,N_24143);
nor UO_1842 (O_1842,N_24677,N_24106);
xnor UO_1843 (O_1843,N_23938,N_24650);
and UO_1844 (O_1844,N_24239,N_23781);
xnor UO_1845 (O_1845,N_24080,N_24557);
and UO_1846 (O_1846,N_24766,N_24961);
xnor UO_1847 (O_1847,N_24046,N_24606);
nor UO_1848 (O_1848,N_24880,N_24072);
or UO_1849 (O_1849,N_23827,N_24242);
nor UO_1850 (O_1850,N_24270,N_24282);
nand UO_1851 (O_1851,N_24780,N_24794);
and UO_1852 (O_1852,N_24170,N_24523);
nand UO_1853 (O_1853,N_24211,N_23796);
and UO_1854 (O_1854,N_24839,N_24486);
nor UO_1855 (O_1855,N_23917,N_24386);
nand UO_1856 (O_1856,N_24476,N_24902);
nand UO_1857 (O_1857,N_23778,N_23922);
and UO_1858 (O_1858,N_24298,N_24316);
or UO_1859 (O_1859,N_23928,N_24902);
and UO_1860 (O_1860,N_23837,N_24177);
and UO_1861 (O_1861,N_24010,N_24068);
xor UO_1862 (O_1862,N_24742,N_24096);
xor UO_1863 (O_1863,N_24203,N_24260);
nand UO_1864 (O_1864,N_24163,N_24326);
nor UO_1865 (O_1865,N_24544,N_24837);
nand UO_1866 (O_1866,N_24771,N_24374);
nand UO_1867 (O_1867,N_24782,N_24066);
nor UO_1868 (O_1868,N_24014,N_24133);
xor UO_1869 (O_1869,N_24385,N_24031);
nand UO_1870 (O_1870,N_24805,N_24452);
and UO_1871 (O_1871,N_24722,N_24069);
nor UO_1872 (O_1872,N_23896,N_23750);
or UO_1873 (O_1873,N_24447,N_24455);
nor UO_1874 (O_1874,N_24626,N_23913);
and UO_1875 (O_1875,N_24296,N_24027);
or UO_1876 (O_1876,N_24959,N_24450);
or UO_1877 (O_1877,N_24442,N_23971);
nor UO_1878 (O_1878,N_24416,N_24931);
or UO_1879 (O_1879,N_24109,N_24473);
or UO_1880 (O_1880,N_24168,N_24783);
and UO_1881 (O_1881,N_24992,N_24655);
xnor UO_1882 (O_1882,N_24765,N_24486);
or UO_1883 (O_1883,N_24556,N_24553);
xor UO_1884 (O_1884,N_24090,N_23915);
nor UO_1885 (O_1885,N_23973,N_24038);
or UO_1886 (O_1886,N_24630,N_23870);
or UO_1887 (O_1887,N_23970,N_24115);
xnor UO_1888 (O_1888,N_24844,N_24101);
or UO_1889 (O_1889,N_24960,N_23784);
nor UO_1890 (O_1890,N_24738,N_23939);
and UO_1891 (O_1891,N_23997,N_23821);
nand UO_1892 (O_1892,N_24140,N_24255);
nor UO_1893 (O_1893,N_24088,N_24255);
or UO_1894 (O_1894,N_24093,N_24402);
or UO_1895 (O_1895,N_24894,N_24659);
and UO_1896 (O_1896,N_24036,N_24467);
xnor UO_1897 (O_1897,N_24081,N_24812);
and UO_1898 (O_1898,N_24766,N_23979);
nand UO_1899 (O_1899,N_24550,N_24839);
nor UO_1900 (O_1900,N_24003,N_23781);
or UO_1901 (O_1901,N_24531,N_24078);
or UO_1902 (O_1902,N_23847,N_24258);
and UO_1903 (O_1903,N_24059,N_24064);
nor UO_1904 (O_1904,N_24217,N_24252);
and UO_1905 (O_1905,N_23794,N_24385);
nand UO_1906 (O_1906,N_24915,N_24124);
xnor UO_1907 (O_1907,N_23799,N_24933);
nand UO_1908 (O_1908,N_23766,N_23847);
xnor UO_1909 (O_1909,N_24263,N_24997);
and UO_1910 (O_1910,N_24664,N_24334);
or UO_1911 (O_1911,N_24934,N_24914);
nor UO_1912 (O_1912,N_24239,N_24104);
and UO_1913 (O_1913,N_24060,N_24881);
xor UO_1914 (O_1914,N_23922,N_24265);
nand UO_1915 (O_1915,N_24219,N_24171);
or UO_1916 (O_1916,N_24628,N_23797);
nor UO_1917 (O_1917,N_24643,N_24813);
nand UO_1918 (O_1918,N_24666,N_23976);
or UO_1919 (O_1919,N_24014,N_24368);
and UO_1920 (O_1920,N_24786,N_24662);
and UO_1921 (O_1921,N_23758,N_24189);
and UO_1922 (O_1922,N_24714,N_23963);
nor UO_1923 (O_1923,N_24570,N_24073);
nor UO_1924 (O_1924,N_24955,N_24367);
or UO_1925 (O_1925,N_24729,N_24590);
nor UO_1926 (O_1926,N_24141,N_24892);
xor UO_1927 (O_1927,N_24855,N_24174);
nor UO_1928 (O_1928,N_24712,N_24368);
nor UO_1929 (O_1929,N_24225,N_23987);
nor UO_1930 (O_1930,N_24327,N_24817);
and UO_1931 (O_1931,N_23804,N_24253);
nor UO_1932 (O_1932,N_24135,N_23870);
nand UO_1933 (O_1933,N_24323,N_24049);
or UO_1934 (O_1934,N_24434,N_24594);
nor UO_1935 (O_1935,N_24881,N_24629);
xnor UO_1936 (O_1936,N_23997,N_24076);
nand UO_1937 (O_1937,N_24960,N_24829);
and UO_1938 (O_1938,N_24756,N_23920);
nand UO_1939 (O_1939,N_24189,N_24088);
xor UO_1940 (O_1940,N_24612,N_24971);
or UO_1941 (O_1941,N_24141,N_24803);
xor UO_1942 (O_1942,N_24501,N_24431);
nand UO_1943 (O_1943,N_24659,N_23780);
nand UO_1944 (O_1944,N_24684,N_23868);
and UO_1945 (O_1945,N_24292,N_24446);
nand UO_1946 (O_1946,N_24788,N_24991);
and UO_1947 (O_1947,N_24838,N_24596);
nand UO_1948 (O_1948,N_23791,N_23873);
nand UO_1949 (O_1949,N_24808,N_23866);
nor UO_1950 (O_1950,N_24327,N_24470);
or UO_1951 (O_1951,N_24958,N_24929);
nor UO_1952 (O_1952,N_24080,N_23838);
nor UO_1953 (O_1953,N_24856,N_23910);
nand UO_1954 (O_1954,N_24478,N_24811);
or UO_1955 (O_1955,N_24008,N_24738);
and UO_1956 (O_1956,N_24818,N_24637);
nand UO_1957 (O_1957,N_24096,N_23869);
nor UO_1958 (O_1958,N_23851,N_24117);
and UO_1959 (O_1959,N_24284,N_24590);
or UO_1960 (O_1960,N_24657,N_23824);
or UO_1961 (O_1961,N_24618,N_24370);
or UO_1962 (O_1962,N_24268,N_24786);
and UO_1963 (O_1963,N_24205,N_23918);
nor UO_1964 (O_1964,N_24519,N_24878);
xnor UO_1965 (O_1965,N_24231,N_24259);
and UO_1966 (O_1966,N_24399,N_23844);
nand UO_1967 (O_1967,N_24499,N_24752);
nand UO_1968 (O_1968,N_24611,N_24293);
or UO_1969 (O_1969,N_24920,N_23762);
xnor UO_1970 (O_1970,N_24169,N_23798);
nor UO_1971 (O_1971,N_24063,N_24744);
nor UO_1972 (O_1972,N_24346,N_23790);
nor UO_1973 (O_1973,N_24053,N_24449);
or UO_1974 (O_1974,N_24755,N_24339);
nand UO_1975 (O_1975,N_24679,N_24212);
nand UO_1976 (O_1976,N_24385,N_24994);
or UO_1977 (O_1977,N_23800,N_23874);
and UO_1978 (O_1978,N_23796,N_24756);
nand UO_1979 (O_1979,N_24877,N_24918);
nor UO_1980 (O_1980,N_24279,N_24015);
and UO_1981 (O_1981,N_24393,N_23961);
nor UO_1982 (O_1982,N_24083,N_24032);
and UO_1983 (O_1983,N_24665,N_24415);
and UO_1984 (O_1984,N_24949,N_24012);
xnor UO_1985 (O_1985,N_24920,N_24572);
xnor UO_1986 (O_1986,N_23817,N_24146);
or UO_1987 (O_1987,N_24141,N_23887);
nor UO_1988 (O_1988,N_24557,N_24904);
nor UO_1989 (O_1989,N_24474,N_24502);
nand UO_1990 (O_1990,N_24498,N_24785);
or UO_1991 (O_1991,N_23828,N_24596);
xor UO_1992 (O_1992,N_24118,N_24746);
nand UO_1993 (O_1993,N_24033,N_23910);
xnor UO_1994 (O_1994,N_24872,N_24032);
nand UO_1995 (O_1995,N_24218,N_24160);
or UO_1996 (O_1996,N_24500,N_23892);
and UO_1997 (O_1997,N_24553,N_24950);
xnor UO_1998 (O_1998,N_24340,N_24235);
and UO_1999 (O_1999,N_24005,N_24903);
nor UO_2000 (O_2000,N_23941,N_23994);
or UO_2001 (O_2001,N_23893,N_24386);
xor UO_2002 (O_2002,N_24040,N_24262);
xor UO_2003 (O_2003,N_24293,N_24662);
nor UO_2004 (O_2004,N_24426,N_24243);
xnor UO_2005 (O_2005,N_24680,N_24561);
or UO_2006 (O_2006,N_24730,N_24924);
or UO_2007 (O_2007,N_24742,N_24154);
or UO_2008 (O_2008,N_23791,N_23949);
and UO_2009 (O_2009,N_23872,N_23926);
or UO_2010 (O_2010,N_24428,N_24934);
and UO_2011 (O_2011,N_24445,N_24903);
nand UO_2012 (O_2012,N_24338,N_23855);
xnor UO_2013 (O_2013,N_24824,N_24583);
nor UO_2014 (O_2014,N_23926,N_24774);
xor UO_2015 (O_2015,N_24854,N_24650);
nor UO_2016 (O_2016,N_24164,N_24479);
nand UO_2017 (O_2017,N_23999,N_24279);
xnor UO_2018 (O_2018,N_24188,N_23851);
xnor UO_2019 (O_2019,N_23908,N_24371);
or UO_2020 (O_2020,N_23750,N_24335);
and UO_2021 (O_2021,N_24199,N_24793);
nor UO_2022 (O_2022,N_24705,N_24355);
xor UO_2023 (O_2023,N_24103,N_23919);
and UO_2024 (O_2024,N_24104,N_24295);
or UO_2025 (O_2025,N_24804,N_24447);
xnor UO_2026 (O_2026,N_24770,N_23885);
nor UO_2027 (O_2027,N_24204,N_24038);
nor UO_2028 (O_2028,N_24520,N_23765);
xor UO_2029 (O_2029,N_24455,N_24418);
nor UO_2030 (O_2030,N_24530,N_24587);
xor UO_2031 (O_2031,N_24830,N_24672);
nand UO_2032 (O_2032,N_24429,N_24934);
nor UO_2033 (O_2033,N_24332,N_24571);
nor UO_2034 (O_2034,N_23991,N_24558);
nor UO_2035 (O_2035,N_24613,N_24879);
xor UO_2036 (O_2036,N_24896,N_23802);
xnor UO_2037 (O_2037,N_24198,N_24152);
xor UO_2038 (O_2038,N_24946,N_24723);
nand UO_2039 (O_2039,N_24700,N_23898);
nor UO_2040 (O_2040,N_24746,N_24680);
xnor UO_2041 (O_2041,N_23838,N_24243);
nand UO_2042 (O_2042,N_24182,N_24974);
and UO_2043 (O_2043,N_24790,N_24750);
nand UO_2044 (O_2044,N_24647,N_24461);
or UO_2045 (O_2045,N_24431,N_24587);
nor UO_2046 (O_2046,N_24139,N_24712);
nand UO_2047 (O_2047,N_24385,N_24485);
and UO_2048 (O_2048,N_24879,N_23867);
or UO_2049 (O_2049,N_24525,N_24334);
nand UO_2050 (O_2050,N_24524,N_24521);
or UO_2051 (O_2051,N_23838,N_24905);
xnor UO_2052 (O_2052,N_24429,N_24762);
xnor UO_2053 (O_2053,N_24632,N_23849);
and UO_2054 (O_2054,N_24737,N_24460);
xor UO_2055 (O_2055,N_24025,N_24075);
xor UO_2056 (O_2056,N_23864,N_24018);
and UO_2057 (O_2057,N_24085,N_24593);
and UO_2058 (O_2058,N_24839,N_24671);
nor UO_2059 (O_2059,N_23834,N_23855);
xor UO_2060 (O_2060,N_24207,N_24139);
xor UO_2061 (O_2061,N_24609,N_24073);
and UO_2062 (O_2062,N_24951,N_24419);
nand UO_2063 (O_2063,N_24148,N_24865);
xor UO_2064 (O_2064,N_24979,N_24424);
nor UO_2065 (O_2065,N_24363,N_23955);
nand UO_2066 (O_2066,N_24629,N_24612);
nor UO_2067 (O_2067,N_24339,N_23941);
nor UO_2068 (O_2068,N_23811,N_24967);
nand UO_2069 (O_2069,N_24045,N_23935);
nor UO_2070 (O_2070,N_24065,N_24553);
nand UO_2071 (O_2071,N_23818,N_24922);
xnor UO_2072 (O_2072,N_24109,N_24776);
xor UO_2073 (O_2073,N_24170,N_24409);
nand UO_2074 (O_2074,N_23858,N_24766);
nand UO_2075 (O_2075,N_23829,N_24803);
xor UO_2076 (O_2076,N_23835,N_23848);
or UO_2077 (O_2077,N_24059,N_24774);
or UO_2078 (O_2078,N_24645,N_24408);
nand UO_2079 (O_2079,N_24639,N_24028);
or UO_2080 (O_2080,N_24716,N_24552);
nor UO_2081 (O_2081,N_24662,N_24209);
or UO_2082 (O_2082,N_24945,N_24390);
and UO_2083 (O_2083,N_23992,N_23761);
xor UO_2084 (O_2084,N_23756,N_24525);
and UO_2085 (O_2085,N_24154,N_24253);
nor UO_2086 (O_2086,N_24846,N_24595);
xnor UO_2087 (O_2087,N_24461,N_24535);
or UO_2088 (O_2088,N_24333,N_23993);
xor UO_2089 (O_2089,N_24350,N_24128);
xor UO_2090 (O_2090,N_24135,N_23888);
xor UO_2091 (O_2091,N_24867,N_24881);
nor UO_2092 (O_2092,N_24480,N_23885);
nand UO_2093 (O_2093,N_24766,N_24711);
or UO_2094 (O_2094,N_23953,N_24929);
nor UO_2095 (O_2095,N_24330,N_23917);
or UO_2096 (O_2096,N_24088,N_24077);
and UO_2097 (O_2097,N_24529,N_24470);
xor UO_2098 (O_2098,N_24763,N_24449);
nand UO_2099 (O_2099,N_24429,N_23922);
and UO_2100 (O_2100,N_24004,N_23755);
and UO_2101 (O_2101,N_24106,N_24797);
nand UO_2102 (O_2102,N_24166,N_24271);
nand UO_2103 (O_2103,N_24215,N_24168);
or UO_2104 (O_2104,N_23838,N_23762);
or UO_2105 (O_2105,N_24030,N_24760);
and UO_2106 (O_2106,N_24716,N_24820);
xor UO_2107 (O_2107,N_24494,N_24407);
or UO_2108 (O_2108,N_24456,N_24336);
xor UO_2109 (O_2109,N_24550,N_24210);
and UO_2110 (O_2110,N_24415,N_23915);
or UO_2111 (O_2111,N_24642,N_24462);
or UO_2112 (O_2112,N_24623,N_24064);
nand UO_2113 (O_2113,N_24098,N_24414);
and UO_2114 (O_2114,N_24818,N_24975);
and UO_2115 (O_2115,N_24292,N_24139);
xnor UO_2116 (O_2116,N_24807,N_24337);
and UO_2117 (O_2117,N_24514,N_24145);
nand UO_2118 (O_2118,N_23982,N_24630);
xor UO_2119 (O_2119,N_24651,N_24181);
nor UO_2120 (O_2120,N_24259,N_24939);
xnor UO_2121 (O_2121,N_24193,N_24396);
xor UO_2122 (O_2122,N_24601,N_24393);
and UO_2123 (O_2123,N_24223,N_24180);
xnor UO_2124 (O_2124,N_24214,N_24289);
nand UO_2125 (O_2125,N_24218,N_24923);
xor UO_2126 (O_2126,N_24848,N_24156);
nand UO_2127 (O_2127,N_24569,N_23874);
xor UO_2128 (O_2128,N_24630,N_24913);
nand UO_2129 (O_2129,N_24972,N_23919);
and UO_2130 (O_2130,N_24860,N_23837);
or UO_2131 (O_2131,N_24105,N_24224);
nand UO_2132 (O_2132,N_23859,N_24298);
xnor UO_2133 (O_2133,N_24372,N_23773);
nor UO_2134 (O_2134,N_24168,N_23759);
and UO_2135 (O_2135,N_24432,N_24825);
nand UO_2136 (O_2136,N_23864,N_24776);
xnor UO_2137 (O_2137,N_24337,N_24720);
nor UO_2138 (O_2138,N_24033,N_23784);
and UO_2139 (O_2139,N_24227,N_23759);
and UO_2140 (O_2140,N_24507,N_24200);
and UO_2141 (O_2141,N_24239,N_24021);
nand UO_2142 (O_2142,N_23910,N_24047);
xor UO_2143 (O_2143,N_23903,N_24181);
or UO_2144 (O_2144,N_24615,N_24918);
nor UO_2145 (O_2145,N_23877,N_24755);
and UO_2146 (O_2146,N_24024,N_24226);
and UO_2147 (O_2147,N_24663,N_24156);
xnor UO_2148 (O_2148,N_24502,N_23930);
or UO_2149 (O_2149,N_24324,N_24780);
nand UO_2150 (O_2150,N_24725,N_24406);
or UO_2151 (O_2151,N_24700,N_24297);
or UO_2152 (O_2152,N_23819,N_24034);
or UO_2153 (O_2153,N_24138,N_24405);
or UO_2154 (O_2154,N_24947,N_24297);
nand UO_2155 (O_2155,N_24280,N_24458);
nor UO_2156 (O_2156,N_24212,N_24296);
nor UO_2157 (O_2157,N_24281,N_24753);
or UO_2158 (O_2158,N_24319,N_24494);
nor UO_2159 (O_2159,N_24596,N_24350);
and UO_2160 (O_2160,N_24093,N_24909);
and UO_2161 (O_2161,N_24280,N_24085);
xor UO_2162 (O_2162,N_24233,N_24265);
or UO_2163 (O_2163,N_24954,N_24266);
xnor UO_2164 (O_2164,N_24171,N_24140);
and UO_2165 (O_2165,N_23998,N_24430);
and UO_2166 (O_2166,N_24926,N_24849);
nor UO_2167 (O_2167,N_24138,N_24126);
nand UO_2168 (O_2168,N_24796,N_24584);
xor UO_2169 (O_2169,N_24515,N_23945);
nand UO_2170 (O_2170,N_24089,N_24966);
and UO_2171 (O_2171,N_24043,N_24399);
nand UO_2172 (O_2172,N_24169,N_24117);
nand UO_2173 (O_2173,N_23812,N_23937);
xor UO_2174 (O_2174,N_23941,N_24460);
and UO_2175 (O_2175,N_24535,N_24282);
xnor UO_2176 (O_2176,N_24216,N_24439);
or UO_2177 (O_2177,N_24541,N_24199);
xor UO_2178 (O_2178,N_24223,N_23973);
or UO_2179 (O_2179,N_24974,N_24559);
nor UO_2180 (O_2180,N_24214,N_23973);
nand UO_2181 (O_2181,N_24472,N_24245);
xor UO_2182 (O_2182,N_24840,N_24991);
and UO_2183 (O_2183,N_23910,N_23992);
nand UO_2184 (O_2184,N_24080,N_24764);
and UO_2185 (O_2185,N_23912,N_24063);
nor UO_2186 (O_2186,N_23826,N_24533);
nor UO_2187 (O_2187,N_23965,N_24198);
xnor UO_2188 (O_2188,N_23971,N_24480);
nor UO_2189 (O_2189,N_24719,N_24749);
or UO_2190 (O_2190,N_24004,N_23771);
nand UO_2191 (O_2191,N_24297,N_23786);
nor UO_2192 (O_2192,N_23995,N_24846);
and UO_2193 (O_2193,N_24716,N_23981);
nand UO_2194 (O_2194,N_24422,N_24345);
nor UO_2195 (O_2195,N_24152,N_24041);
xor UO_2196 (O_2196,N_24455,N_24265);
or UO_2197 (O_2197,N_23846,N_24277);
nand UO_2198 (O_2198,N_24766,N_23874);
and UO_2199 (O_2199,N_24090,N_24647);
and UO_2200 (O_2200,N_23851,N_24562);
nand UO_2201 (O_2201,N_24153,N_24149);
or UO_2202 (O_2202,N_24459,N_24292);
nor UO_2203 (O_2203,N_24545,N_24528);
xnor UO_2204 (O_2204,N_24222,N_23858);
xor UO_2205 (O_2205,N_24037,N_24238);
and UO_2206 (O_2206,N_24726,N_24669);
or UO_2207 (O_2207,N_24759,N_23979);
xnor UO_2208 (O_2208,N_23897,N_24723);
and UO_2209 (O_2209,N_24361,N_24800);
nor UO_2210 (O_2210,N_24428,N_24780);
xnor UO_2211 (O_2211,N_24446,N_24622);
or UO_2212 (O_2212,N_24826,N_24560);
nor UO_2213 (O_2213,N_24366,N_24720);
nor UO_2214 (O_2214,N_23825,N_24491);
nor UO_2215 (O_2215,N_24498,N_23778);
xor UO_2216 (O_2216,N_24238,N_23858);
and UO_2217 (O_2217,N_24653,N_24623);
or UO_2218 (O_2218,N_24789,N_24393);
nand UO_2219 (O_2219,N_24748,N_24571);
xnor UO_2220 (O_2220,N_23790,N_23872);
nor UO_2221 (O_2221,N_24759,N_24888);
nor UO_2222 (O_2222,N_24214,N_24204);
xor UO_2223 (O_2223,N_24967,N_23909);
or UO_2224 (O_2224,N_24393,N_24962);
xnor UO_2225 (O_2225,N_24703,N_24704);
or UO_2226 (O_2226,N_24973,N_24535);
xor UO_2227 (O_2227,N_23820,N_23888);
nand UO_2228 (O_2228,N_24791,N_24331);
xor UO_2229 (O_2229,N_23775,N_23924);
nor UO_2230 (O_2230,N_24990,N_24981);
nand UO_2231 (O_2231,N_24348,N_24265);
and UO_2232 (O_2232,N_24058,N_24060);
nor UO_2233 (O_2233,N_24552,N_24906);
nor UO_2234 (O_2234,N_24768,N_24025);
nand UO_2235 (O_2235,N_24599,N_23896);
and UO_2236 (O_2236,N_24118,N_24043);
and UO_2237 (O_2237,N_24524,N_24325);
and UO_2238 (O_2238,N_24143,N_24782);
nor UO_2239 (O_2239,N_24917,N_24381);
xor UO_2240 (O_2240,N_24429,N_24382);
nor UO_2241 (O_2241,N_24373,N_24708);
or UO_2242 (O_2242,N_23992,N_23771);
and UO_2243 (O_2243,N_23791,N_24890);
and UO_2244 (O_2244,N_24145,N_24772);
nand UO_2245 (O_2245,N_24288,N_23867);
nor UO_2246 (O_2246,N_23804,N_24950);
nor UO_2247 (O_2247,N_23753,N_23841);
nand UO_2248 (O_2248,N_24905,N_24205);
or UO_2249 (O_2249,N_23754,N_24023);
or UO_2250 (O_2250,N_24502,N_24783);
or UO_2251 (O_2251,N_24274,N_24467);
or UO_2252 (O_2252,N_23814,N_24109);
nand UO_2253 (O_2253,N_24392,N_24798);
nand UO_2254 (O_2254,N_24016,N_23862);
and UO_2255 (O_2255,N_24525,N_24206);
nor UO_2256 (O_2256,N_23953,N_24548);
nor UO_2257 (O_2257,N_24513,N_24967);
and UO_2258 (O_2258,N_24800,N_24006);
nand UO_2259 (O_2259,N_24577,N_24508);
nand UO_2260 (O_2260,N_23907,N_24855);
nand UO_2261 (O_2261,N_24063,N_24275);
or UO_2262 (O_2262,N_24517,N_24086);
and UO_2263 (O_2263,N_24192,N_24103);
nand UO_2264 (O_2264,N_24338,N_24512);
and UO_2265 (O_2265,N_24650,N_24222);
and UO_2266 (O_2266,N_23921,N_24122);
nand UO_2267 (O_2267,N_23834,N_24003);
and UO_2268 (O_2268,N_23755,N_24845);
and UO_2269 (O_2269,N_23807,N_24128);
and UO_2270 (O_2270,N_24767,N_24656);
or UO_2271 (O_2271,N_24091,N_23917);
and UO_2272 (O_2272,N_24956,N_24389);
nor UO_2273 (O_2273,N_24148,N_24618);
or UO_2274 (O_2274,N_24254,N_24097);
nand UO_2275 (O_2275,N_24943,N_24885);
or UO_2276 (O_2276,N_24129,N_23993);
or UO_2277 (O_2277,N_24348,N_24900);
and UO_2278 (O_2278,N_24371,N_24836);
nor UO_2279 (O_2279,N_24480,N_24094);
nor UO_2280 (O_2280,N_24728,N_23878);
nand UO_2281 (O_2281,N_23981,N_24401);
nand UO_2282 (O_2282,N_24195,N_24995);
or UO_2283 (O_2283,N_23773,N_24896);
or UO_2284 (O_2284,N_24247,N_24476);
or UO_2285 (O_2285,N_24666,N_24373);
nor UO_2286 (O_2286,N_23883,N_24691);
xnor UO_2287 (O_2287,N_24323,N_24593);
xor UO_2288 (O_2288,N_23999,N_23781);
nor UO_2289 (O_2289,N_24656,N_23843);
and UO_2290 (O_2290,N_23899,N_24935);
xor UO_2291 (O_2291,N_24540,N_24028);
and UO_2292 (O_2292,N_24658,N_24504);
xnor UO_2293 (O_2293,N_24654,N_24545);
xnor UO_2294 (O_2294,N_24585,N_24741);
nor UO_2295 (O_2295,N_24306,N_24655);
or UO_2296 (O_2296,N_24011,N_23763);
and UO_2297 (O_2297,N_23929,N_24893);
nand UO_2298 (O_2298,N_24401,N_23883);
and UO_2299 (O_2299,N_23846,N_24022);
and UO_2300 (O_2300,N_24037,N_23871);
nor UO_2301 (O_2301,N_24407,N_24641);
or UO_2302 (O_2302,N_24275,N_24697);
or UO_2303 (O_2303,N_24149,N_24407);
nand UO_2304 (O_2304,N_24330,N_24134);
nor UO_2305 (O_2305,N_24046,N_23998);
nand UO_2306 (O_2306,N_24046,N_24902);
and UO_2307 (O_2307,N_24522,N_24560);
nor UO_2308 (O_2308,N_24580,N_24636);
nor UO_2309 (O_2309,N_24202,N_24674);
xnor UO_2310 (O_2310,N_24882,N_24569);
nand UO_2311 (O_2311,N_24135,N_24563);
or UO_2312 (O_2312,N_24172,N_24622);
nand UO_2313 (O_2313,N_24499,N_24656);
xor UO_2314 (O_2314,N_24038,N_24706);
nor UO_2315 (O_2315,N_23888,N_24637);
nand UO_2316 (O_2316,N_24871,N_24810);
and UO_2317 (O_2317,N_24734,N_23982);
nand UO_2318 (O_2318,N_24551,N_24265);
and UO_2319 (O_2319,N_24471,N_24546);
nor UO_2320 (O_2320,N_24573,N_24736);
nand UO_2321 (O_2321,N_24951,N_24186);
nand UO_2322 (O_2322,N_24971,N_24788);
and UO_2323 (O_2323,N_24061,N_24996);
nor UO_2324 (O_2324,N_24232,N_23931);
xnor UO_2325 (O_2325,N_24983,N_23934);
nand UO_2326 (O_2326,N_24846,N_23948);
xor UO_2327 (O_2327,N_24405,N_24587);
and UO_2328 (O_2328,N_23794,N_24302);
or UO_2329 (O_2329,N_24779,N_24006);
and UO_2330 (O_2330,N_24659,N_24673);
nand UO_2331 (O_2331,N_24666,N_24007);
and UO_2332 (O_2332,N_24493,N_24838);
or UO_2333 (O_2333,N_24149,N_24907);
xor UO_2334 (O_2334,N_24460,N_24645);
or UO_2335 (O_2335,N_24478,N_23928);
or UO_2336 (O_2336,N_23906,N_24706);
nand UO_2337 (O_2337,N_24685,N_23990);
or UO_2338 (O_2338,N_24133,N_24714);
xor UO_2339 (O_2339,N_23935,N_23878);
nand UO_2340 (O_2340,N_24705,N_24458);
and UO_2341 (O_2341,N_24892,N_24461);
and UO_2342 (O_2342,N_24891,N_24216);
nand UO_2343 (O_2343,N_24346,N_24396);
xor UO_2344 (O_2344,N_24996,N_24127);
or UO_2345 (O_2345,N_24018,N_24791);
nor UO_2346 (O_2346,N_24144,N_23952);
nor UO_2347 (O_2347,N_24653,N_24027);
and UO_2348 (O_2348,N_24766,N_24155);
or UO_2349 (O_2349,N_24082,N_24140);
nand UO_2350 (O_2350,N_24087,N_23991);
and UO_2351 (O_2351,N_24435,N_23879);
xnor UO_2352 (O_2352,N_24071,N_23944);
or UO_2353 (O_2353,N_24824,N_24595);
and UO_2354 (O_2354,N_24835,N_24224);
nor UO_2355 (O_2355,N_24348,N_24754);
nand UO_2356 (O_2356,N_24375,N_24880);
or UO_2357 (O_2357,N_24487,N_24341);
or UO_2358 (O_2358,N_24259,N_24625);
or UO_2359 (O_2359,N_24568,N_23966);
or UO_2360 (O_2360,N_23781,N_23981);
nor UO_2361 (O_2361,N_24779,N_24539);
or UO_2362 (O_2362,N_24085,N_23857);
or UO_2363 (O_2363,N_24327,N_24737);
or UO_2364 (O_2364,N_24794,N_24305);
xor UO_2365 (O_2365,N_24829,N_24410);
nand UO_2366 (O_2366,N_24747,N_24076);
and UO_2367 (O_2367,N_24575,N_24289);
xnor UO_2368 (O_2368,N_24645,N_23774);
or UO_2369 (O_2369,N_24326,N_24351);
nand UO_2370 (O_2370,N_23796,N_24212);
nand UO_2371 (O_2371,N_24571,N_24383);
and UO_2372 (O_2372,N_24577,N_24475);
nand UO_2373 (O_2373,N_24479,N_24380);
nor UO_2374 (O_2374,N_24831,N_24874);
xnor UO_2375 (O_2375,N_24592,N_24326);
nand UO_2376 (O_2376,N_24037,N_24795);
and UO_2377 (O_2377,N_24593,N_24826);
and UO_2378 (O_2378,N_24375,N_24234);
nand UO_2379 (O_2379,N_24905,N_23928);
xnor UO_2380 (O_2380,N_24303,N_24731);
nand UO_2381 (O_2381,N_24868,N_24903);
xor UO_2382 (O_2382,N_24207,N_23843);
nand UO_2383 (O_2383,N_24031,N_23825);
xor UO_2384 (O_2384,N_24472,N_24322);
nand UO_2385 (O_2385,N_24350,N_24922);
nand UO_2386 (O_2386,N_23914,N_23840);
and UO_2387 (O_2387,N_23942,N_24287);
nand UO_2388 (O_2388,N_24094,N_24888);
xor UO_2389 (O_2389,N_24067,N_24004);
nor UO_2390 (O_2390,N_24520,N_23753);
xnor UO_2391 (O_2391,N_24741,N_24397);
nand UO_2392 (O_2392,N_24448,N_24626);
and UO_2393 (O_2393,N_23904,N_24410);
nand UO_2394 (O_2394,N_23920,N_24400);
nor UO_2395 (O_2395,N_24665,N_24072);
or UO_2396 (O_2396,N_23952,N_24102);
nand UO_2397 (O_2397,N_23825,N_24237);
or UO_2398 (O_2398,N_24776,N_24366);
and UO_2399 (O_2399,N_24830,N_24699);
or UO_2400 (O_2400,N_24183,N_23771);
xor UO_2401 (O_2401,N_23967,N_24000);
nand UO_2402 (O_2402,N_24666,N_24457);
nand UO_2403 (O_2403,N_24497,N_23889);
xor UO_2404 (O_2404,N_23944,N_24862);
nor UO_2405 (O_2405,N_24268,N_24973);
nor UO_2406 (O_2406,N_24954,N_24854);
and UO_2407 (O_2407,N_24142,N_24506);
nand UO_2408 (O_2408,N_24177,N_24275);
or UO_2409 (O_2409,N_24242,N_24892);
and UO_2410 (O_2410,N_24253,N_24408);
and UO_2411 (O_2411,N_24614,N_23806);
nand UO_2412 (O_2412,N_24529,N_24658);
nor UO_2413 (O_2413,N_24551,N_23827);
and UO_2414 (O_2414,N_24546,N_24339);
nand UO_2415 (O_2415,N_24530,N_24202);
and UO_2416 (O_2416,N_23963,N_23916);
xor UO_2417 (O_2417,N_24030,N_24723);
nand UO_2418 (O_2418,N_24179,N_24507);
xnor UO_2419 (O_2419,N_24809,N_24007);
and UO_2420 (O_2420,N_24509,N_23776);
nand UO_2421 (O_2421,N_24883,N_24834);
nand UO_2422 (O_2422,N_24054,N_24473);
nand UO_2423 (O_2423,N_24614,N_23771);
xnor UO_2424 (O_2424,N_24792,N_24697);
nor UO_2425 (O_2425,N_23888,N_23773);
nand UO_2426 (O_2426,N_24969,N_24804);
xnor UO_2427 (O_2427,N_24006,N_23843);
nor UO_2428 (O_2428,N_23919,N_24450);
nor UO_2429 (O_2429,N_24484,N_23829);
nor UO_2430 (O_2430,N_24103,N_24828);
xor UO_2431 (O_2431,N_23875,N_24082);
nor UO_2432 (O_2432,N_23775,N_24817);
nor UO_2433 (O_2433,N_24800,N_24923);
or UO_2434 (O_2434,N_24323,N_23772);
and UO_2435 (O_2435,N_24359,N_24122);
or UO_2436 (O_2436,N_24527,N_24191);
xnor UO_2437 (O_2437,N_23974,N_24509);
and UO_2438 (O_2438,N_24361,N_24197);
nand UO_2439 (O_2439,N_24686,N_24662);
and UO_2440 (O_2440,N_24529,N_24176);
xor UO_2441 (O_2441,N_24750,N_24986);
or UO_2442 (O_2442,N_24315,N_23806);
and UO_2443 (O_2443,N_24992,N_24570);
xor UO_2444 (O_2444,N_24209,N_24668);
or UO_2445 (O_2445,N_24150,N_24880);
and UO_2446 (O_2446,N_24783,N_24293);
or UO_2447 (O_2447,N_24856,N_23992);
or UO_2448 (O_2448,N_24873,N_24626);
or UO_2449 (O_2449,N_24977,N_23878);
nand UO_2450 (O_2450,N_24556,N_24846);
and UO_2451 (O_2451,N_24066,N_24537);
or UO_2452 (O_2452,N_24691,N_24003);
nor UO_2453 (O_2453,N_24586,N_24965);
and UO_2454 (O_2454,N_24238,N_24645);
xnor UO_2455 (O_2455,N_24950,N_24964);
or UO_2456 (O_2456,N_24819,N_24923);
or UO_2457 (O_2457,N_24336,N_24096);
and UO_2458 (O_2458,N_24529,N_23776);
and UO_2459 (O_2459,N_23808,N_24703);
nand UO_2460 (O_2460,N_23802,N_23755);
or UO_2461 (O_2461,N_24072,N_23789);
or UO_2462 (O_2462,N_23845,N_23943);
or UO_2463 (O_2463,N_24824,N_24087);
and UO_2464 (O_2464,N_24122,N_24872);
nor UO_2465 (O_2465,N_24750,N_24974);
nor UO_2466 (O_2466,N_23752,N_24948);
and UO_2467 (O_2467,N_23938,N_24950);
xor UO_2468 (O_2468,N_24255,N_24044);
or UO_2469 (O_2469,N_24710,N_24719);
nor UO_2470 (O_2470,N_23888,N_23777);
xor UO_2471 (O_2471,N_24281,N_24320);
or UO_2472 (O_2472,N_24070,N_24349);
nand UO_2473 (O_2473,N_24668,N_24060);
and UO_2474 (O_2474,N_24553,N_24786);
or UO_2475 (O_2475,N_24824,N_24249);
and UO_2476 (O_2476,N_23864,N_24912);
nor UO_2477 (O_2477,N_24525,N_24897);
nand UO_2478 (O_2478,N_23890,N_24887);
nand UO_2479 (O_2479,N_24553,N_24974);
and UO_2480 (O_2480,N_24221,N_24519);
nand UO_2481 (O_2481,N_24493,N_23821);
xor UO_2482 (O_2482,N_24413,N_24998);
and UO_2483 (O_2483,N_23877,N_24588);
or UO_2484 (O_2484,N_24338,N_24619);
nand UO_2485 (O_2485,N_23949,N_24350);
xnor UO_2486 (O_2486,N_24459,N_24524);
or UO_2487 (O_2487,N_24556,N_24001);
and UO_2488 (O_2488,N_24063,N_24856);
and UO_2489 (O_2489,N_24238,N_24986);
and UO_2490 (O_2490,N_23931,N_24936);
xor UO_2491 (O_2491,N_23797,N_24455);
nor UO_2492 (O_2492,N_23904,N_23984);
xnor UO_2493 (O_2493,N_24526,N_23981);
nand UO_2494 (O_2494,N_24895,N_23905);
or UO_2495 (O_2495,N_24376,N_24479);
or UO_2496 (O_2496,N_24345,N_23767);
or UO_2497 (O_2497,N_23819,N_24582);
nand UO_2498 (O_2498,N_24337,N_24061);
or UO_2499 (O_2499,N_24338,N_24902);
xnor UO_2500 (O_2500,N_23848,N_24238);
and UO_2501 (O_2501,N_24958,N_24734);
nand UO_2502 (O_2502,N_24699,N_24281);
nor UO_2503 (O_2503,N_24483,N_24084);
nand UO_2504 (O_2504,N_24689,N_23855);
nor UO_2505 (O_2505,N_24752,N_24400);
nor UO_2506 (O_2506,N_24209,N_24264);
xnor UO_2507 (O_2507,N_24736,N_24975);
xor UO_2508 (O_2508,N_23899,N_24810);
and UO_2509 (O_2509,N_24403,N_24372);
and UO_2510 (O_2510,N_24532,N_24248);
xor UO_2511 (O_2511,N_24580,N_24285);
and UO_2512 (O_2512,N_24038,N_24676);
or UO_2513 (O_2513,N_24402,N_24640);
nand UO_2514 (O_2514,N_23804,N_23987);
or UO_2515 (O_2515,N_23759,N_24038);
or UO_2516 (O_2516,N_24620,N_24826);
nor UO_2517 (O_2517,N_23948,N_24858);
nand UO_2518 (O_2518,N_24923,N_24687);
or UO_2519 (O_2519,N_24841,N_24354);
and UO_2520 (O_2520,N_23863,N_24865);
nand UO_2521 (O_2521,N_24363,N_24317);
and UO_2522 (O_2522,N_23825,N_24004);
and UO_2523 (O_2523,N_24977,N_24489);
and UO_2524 (O_2524,N_23996,N_24510);
nor UO_2525 (O_2525,N_24470,N_23934);
and UO_2526 (O_2526,N_24948,N_24339);
or UO_2527 (O_2527,N_24339,N_24353);
nor UO_2528 (O_2528,N_23968,N_24888);
or UO_2529 (O_2529,N_24679,N_24122);
and UO_2530 (O_2530,N_24332,N_23800);
and UO_2531 (O_2531,N_24999,N_24346);
nand UO_2532 (O_2532,N_24612,N_24722);
nor UO_2533 (O_2533,N_23962,N_24604);
or UO_2534 (O_2534,N_24057,N_24401);
nand UO_2535 (O_2535,N_24831,N_24919);
xor UO_2536 (O_2536,N_24943,N_24836);
xnor UO_2537 (O_2537,N_24182,N_24030);
nor UO_2538 (O_2538,N_24780,N_24576);
nand UO_2539 (O_2539,N_24148,N_24464);
xnor UO_2540 (O_2540,N_24139,N_24271);
and UO_2541 (O_2541,N_24300,N_23837);
nand UO_2542 (O_2542,N_24522,N_24251);
and UO_2543 (O_2543,N_23984,N_24049);
nor UO_2544 (O_2544,N_24356,N_24588);
and UO_2545 (O_2545,N_23899,N_24353);
xnor UO_2546 (O_2546,N_24433,N_23759);
xor UO_2547 (O_2547,N_24699,N_24997);
and UO_2548 (O_2548,N_24397,N_24010);
nand UO_2549 (O_2549,N_24455,N_23872);
or UO_2550 (O_2550,N_24333,N_24510);
and UO_2551 (O_2551,N_24356,N_24455);
xor UO_2552 (O_2552,N_24107,N_24810);
or UO_2553 (O_2553,N_24984,N_24778);
xnor UO_2554 (O_2554,N_23784,N_24225);
xor UO_2555 (O_2555,N_23782,N_24483);
nand UO_2556 (O_2556,N_24922,N_24782);
nor UO_2557 (O_2557,N_24427,N_23914);
xnor UO_2558 (O_2558,N_24930,N_24466);
nand UO_2559 (O_2559,N_24666,N_24937);
xor UO_2560 (O_2560,N_24691,N_24399);
nand UO_2561 (O_2561,N_24052,N_24359);
nand UO_2562 (O_2562,N_24639,N_24160);
nand UO_2563 (O_2563,N_23843,N_24977);
or UO_2564 (O_2564,N_24109,N_23842);
nor UO_2565 (O_2565,N_24887,N_24810);
nor UO_2566 (O_2566,N_24968,N_24839);
or UO_2567 (O_2567,N_24975,N_23842);
nand UO_2568 (O_2568,N_24884,N_24477);
xnor UO_2569 (O_2569,N_24225,N_24152);
xor UO_2570 (O_2570,N_24432,N_24017);
nor UO_2571 (O_2571,N_24895,N_24186);
xnor UO_2572 (O_2572,N_24551,N_24986);
xor UO_2573 (O_2573,N_24579,N_24494);
and UO_2574 (O_2574,N_24975,N_24680);
or UO_2575 (O_2575,N_23758,N_24789);
or UO_2576 (O_2576,N_24722,N_24752);
nor UO_2577 (O_2577,N_24150,N_24090);
or UO_2578 (O_2578,N_23929,N_24425);
nand UO_2579 (O_2579,N_24047,N_24515);
and UO_2580 (O_2580,N_24989,N_24244);
or UO_2581 (O_2581,N_24846,N_24819);
nand UO_2582 (O_2582,N_24977,N_23844);
xor UO_2583 (O_2583,N_24448,N_23920);
and UO_2584 (O_2584,N_24279,N_24373);
or UO_2585 (O_2585,N_24343,N_24804);
nor UO_2586 (O_2586,N_23859,N_24346);
nand UO_2587 (O_2587,N_24685,N_24097);
or UO_2588 (O_2588,N_24009,N_24079);
or UO_2589 (O_2589,N_23988,N_23832);
and UO_2590 (O_2590,N_24984,N_24956);
or UO_2591 (O_2591,N_24602,N_23903);
xor UO_2592 (O_2592,N_23973,N_24611);
or UO_2593 (O_2593,N_23852,N_24632);
and UO_2594 (O_2594,N_23993,N_24925);
xor UO_2595 (O_2595,N_24881,N_24828);
nand UO_2596 (O_2596,N_24685,N_24756);
nand UO_2597 (O_2597,N_24922,N_23956);
or UO_2598 (O_2598,N_24834,N_24726);
nor UO_2599 (O_2599,N_24001,N_24640);
nor UO_2600 (O_2600,N_23867,N_24186);
nand UO_2601 (O_2601,N_24821,N_24198);
or UO_2602 (O_2602,N_23963,N_24129);
xnor UO_2603 (O_2603,N_24866,N_24257);
xor UO_2604 (O_2604,N_24169,N_24951);
nand UO_2605 (O_2605,N_23810,N_24721);
nand UO_2606 (O_2606,N_23947,N_24146);
nor UO_2607 (O_2607,N_24340,N_24133);
nand UO_2608 (O_2608,N_24569,N_23935);
nand UO_2609 (O_2609,N_23789,N_24181);
nand UO_2610 (O_2610,N_23972,N_24467);
and UO_2611 (O_2611,N_23941,N_24748);
nor UO_2612 (O_2612,N_24004,N_24364);
nand UO_2613 (O_2613,N_24761,N_24721);
nand UO_2614 (O_2614,N_24534,N_24151);
and UO_2615 (O_2615,N_23991,N_24816);
or UO_2616 (O_2616,N_24237,N_24134);
nor UO_2617 (O_2617,N_24808,N_24208);
nand UO_2618 (O_2618,N_24167,N_24074);
xor UO_2619 (O_2619,N_24999,N_23775);
nand UO_2620 (O_2620,N_24698,N_24221);
nor UO_2621 (O_2621,N_23881,N_23942);
xnor UO_2622 (O_2622,N_23952,N_23806);
and UO_2623 (O_2623,N_24110,N_24466);
or UO_2624 (O_2624,N_23985,N_24389);
xor UO_2625 (O_2625,N_23833,N_24586);
or UO_2626 (O_2626,N_24910,N_24922);
and UO_2627 (O_2627,N_23752,N_23976);
nand UO_2628 (O_2628,N_23821,N_23848);
nor UO_2629 (O_2629,N_24481,N_24523);
and UO_2630 (O_2630,N_24200,N_24312);
nand UO_2631 (O_2631,N_24428,N_23817);
nor UO_2632 (O_2632,N_24725,N_24861);
or UO_2633 (O_2633,N_24879,N_24575);
nand UO_2634 (O_2634,N_24907,N_24100);
or UO_2635 (O_2635,N_24574,N_24998);
xnor UO_2636 (O_2636,N_24240,N_23764);
or UO_2637 (O_2637,N_24001,N_24173);
or UO_2638 (O_2638,N_24976,N_24022);
nor UO_2639 (O_2639,N_24930,N_24264);
nor UO_2640 (O_2640,N_23842,N_24800);
nor UO_2641 (O_2641,N_24540,N_24283);
and UO_2642 (O_2642,N_24074,N_23777);
and UO_2643 (O_2643,N_24575,N_24111);
nand UO_2644 (O_2644,N_24037,N_24621);
xor UO_2645 (O_2645,N_24103,N_24464);
nand UO_2646 (O_2646,N_24085,N_24094);
or UO_2647 (O_2647,N_24249,N_24539);
nand UO_2648 (O_2648,N_23925,N_24366);
nand UO_2649 (O_2649,N_24998,N_23908);
and UO_2650 (O_2650,N_24955,N_24199);
xnor UO_2651 (O_2651,N_23874,N_24197);
nand UO_2652 (O_2652,N_24152,N_24071);
nand UO_2653 (O_2653,N_23981,N_24815);
or UO_2654 (O_2654,N_24978,N_24251);
xor UO_2655 (O_2655,N_24121,N_24329);
nand UO_2656 (O_2656,N_24440,N_24899);
nand UO_2657 (O_2657,N_23928,N_24680);
nor UO_2658 (O_2658,N_23829,N_24958);
or UO_2659 (O_2659,N_24129,N_24011);
nor UO_2660 (O_2660,N_23763,N_24833);
nor UO_2661 (O_2661,N_24652,N_24127);
and UO_2662 (O_2662,N_24346,N_24637);
and UO_2663 (O_2663,N_24011,N_23845);
nor UO_2664 (O_2664,N_23801,N_24006);
or UO_2665 (O_2665,N_24617,N_24791);
xor UO_2666 (O_2666,N_23877,N_23792);
nor UO_2667 (O_2667,N_24735,N_24200);
xnor UO_2668 (O_2668,N_24826,N_24438);
nand UO_2669 (O_2669,N_24062,N_24012);
nor UO_2670 (O_2670,N_24812,N_24089);
or UO_2671 (O_2671,N_24501,N_24988);
nor UO_2672 (O_2672,N_24550,N_24253);
nor UO_2673 (O_2673,N_24580,N_24003);
nor UO_2674 (O_2674,N_24961,N_24900);
and UO_2675 (O_2675,N_24650,N_24728);
xor UO_2676 (O_2676,N_23936,N_23961);
xor UO_2677 (O_2677,N_24428,N_24340);
nor UO_2678 (O_2678,N_24503,N_24062);
xor UO_2679 (O_2679,N_24492,N_24859);
nand UO_2680 (O_2680,N_24867,N_24771);
xor UO_2681 (O_2681,N_23947,N_24460);
or UO_2682 (O_2682,N_24172,N_23951);
and UO_2683 (O_2683,N_23898,N_24038);
nand UO_2684 (O_2684,N_24996,N_24168);
and UO_2685 (O_2685,N_24879,N_24420);
or UO_2686 (O_2686,N_23888,N_24947);
and UO_2687 (O_2687,N_23769,N_24459);
and UO_2688 (O_2688,N_24420,N_24014);
xnor UO_2689 (O_2689,N_24722,N_24874);
or UO_2690 (O_2690,N_24071,N_23915);
or UO_2691 (O_2691,N_24218,N_24323);
xnor UO_2692 (O_2692,N_24807,N_24545);
nand UO_2693 (O_2693,N_24429,N_24523);
nor UO_2694 (O_2694,N_24037,N_24642);
nand UO_2695 (O_2695,N_24587,N_24816);
nor UO_2696 (O_2696,N_24644,N_24429);
nor UO_2697 (O_2697,N_24289,N_24380);
xor UO_2698 (O_2698,N_24176,N_24995);
or UO_2699 (O_2699,N_24851,N_24171);
and UO_2700 (O_2700,N_23813,N_24373);
nand UO_2701 (O_2701,N_23817,N_24673);
nand UO_2702 (O_2702,N_24755,N_24347);
or UO_2703 (O_2703,N_24084,N_24509);
and UO_2704 (O_2704,N_24288,N_24086);
and UO_2705 (O_2705,N_24777,N_24430);
and UO_2706 (O_2706,N_24767,N_24136);
nand UO_2707 (O_2707,N_24492,N_24965);
nand UO_2708 (O_2708,N_24305,N_24808);
nor UO_2709 (O_2709,N_24346,N_24503);
nand UO_2710 (O_2710,N_24091,N_24918);
nand UO_2711 (O_2711,N_24001,N_24153);
or UO_2712 (O_2712,N_24774,N_23936);
nor UO_2713 (O_2713,N_24118,N_24121);
nor UO_2714 (O_2714,N_24536,N_24036);
and UO_2715 (O_2715,N_24829,N_23804);
nor UO_2716 (O_2716,N_24484,N_24491);
and UO_2717 (O_2717,N_23775,N_24441);
xor UO_2718 (O_2718,N_24444,N_24629);
xor UO_2719 (O_2719,N_24998,N_24674);
nand UO_2720 (O_2720,N_24886,N_23800);
nand UO_2721 (O_2721,N_24738,N_24923);
and UO_2722 (O_2722,N_24586,N_24576);
or UO_2723 (O_2723,N_24789,N_24615);
nand UO_2724 (O_2724,N_24063,N_24902);
and UO_2725 (O_2725,N_24912,N_24182);
xnor UO_2726 (O_2726,N_24277,N_24154);
and UO_2727 (O_2727,N_24534,N_24399);
nand UO_2728 (O_2728,N_24432,N_24180);
and UO_2729 (O_2729,N_24386,N_24688);
nor UO_2730 (O_2730,N_24068,N_24194);
xnor UO_2731 (O_2731,N_24369,N_24452);
xnor UO_2732 (O_2732,N_24754,N_23912);
or UO_2733 (O_2733,N_24518,N_24414);
or UO_2734 (O_2734,N_24738,N_24974);
or UO_2735 (O_2735,N_24883,N_24680);
xnor UO_2736 (O_2736,N_23875,N_24136);
nor UO_2737 (O_2737,N_24075,N_24648);
nand UO_2738 (O_2738,N_24137,N_23931);
or UO_2739 (O_2739,N_24459,N_24976);
nand UO_2740 (O_2740,N_23889,N_24086);
and UO_2741 (O_2741,N_24241,N_24877);
nand UO_2742 (O_2742,N_24387,N_24839);
nand UO_2743 (O_2743,N_24831,N_23877);
xor UO_2744 (O_2744,N_24712,N_24690);
nor UO_2745 (O_2745,N_24531,N_24376);
xnor UO_2746 (O_2746,N_24708,N_23890);
and UO_2747 (O_2747,N_24204,N_24241);
nand UO_2748 (O_2748,N_24000,N_23869);
nand UO_2749 (O_2749,N_24382,N_24646);
nor UO_2750 (O_2750,N_24816,N_24829);
nand UO_2751 (O_2751,N_24040,N_24861);
nand UO_2752 (O_2752,N_24219,N_24716);
xnor UO_2753 (O_2753,N_24854,N_24028);
or UO_2754 (O_2754,N_24142,N_23784);
or UO_2755 (O_2755,N_24431,N_24343);
or UO_2756 (O_2756,N_24255,N_24929);
or UO_2757 (O_2757,N_23817,N_24993);
nor UO_2758 (O_2758,N_24728,N_24910);
or UO_2759 (O_2759,N_24271,N_24789);
xor UO_2760 (O_2760,N_24554,N_23753);
nor UO_2761 (O_2761,N_24024,N_24386);
nand UO_2762 (O_2762,N_24921,N_23872);
nand UO_2763 (O_2763,N_24324,N_24370);
or UO_2764 (O_2764,N_24634,N_24088);
and UO_2765 (O_2765,N_24548,N_24608);
and UO_2766 (O_2766,N_24895,N_24343);
nor UO_2767 (O_2767,N_24311,N_24377);
nor UO_2768 (O_2768,N_24161,N_24397);
or UO_2769 (O_2769,N_24269,N_24566);
nor UO_2770 (O_2770,N_24572,N_24974);
or UO_2771 (O_2771,N_24588,N_24362);
or UO_2772 (O_2772,N_24993,N_23985);
nand UO_2773 (O_2773,N_24202,N_24549);
xor UO_2774 (O_2774,N_24425,N_24719);
xnor UO_2775 (O_2775,N_23939,N_24581);
nand UO_2776 (O_2776,N_23854,N_24690);
or UO_2777 (O_2777,N_24010,N_23785);
nor UO_2778 (O_2778,N_24933,N_24682);
nor UO_2779 (O_2779,N_24460,N_23878);
nor UO_2780 (O_2780,N_23908,N_24892);
xor UO_2781 (O_2781,N_24377,N_24390);
nor UO_2782 (O_2782,N_24704,N_24663);
nor UO_2783 (O_2783,N_24135,N_24976);
nand UO_2784 (O_2784,N_24596,N_23948);
or UO_2785 (O_2785,N_24607,N_23904);
nand UO_2786 (O_2786,N_24649,N_24493);
or UO_2787 (O_2787,N_24201,N_24342);
nor UO_2788 (O_2788,N_24031,N_23887);
xnor UO_2789 (O_2789,N_24849,N_23946);
xnor UO_2790 (O_2790,N_23905,N_24906);
or UO_2791 (O_2791,N_24114,N_24842);
xnor UO_2792 (O_2792,N_24242,N_24327);
or UO_2793 (O_2793,N_24066,N_24387);
nor UO_2794 (O_2794,N_24107,N_24732);
and UO_2795 (O_2795,N_24994,N_24361);
and UO_2796 (O_2796,N_23983,N_24662);
nor UO_2797 (O_2797,N_24552,N_24545);
nor UO_2798 (O_2798,N_24521,N_23912);
nor UO_2799 (O_2799,N_24186,N_24890);
and UO_2800 (O_2800,N_24391,N_24282);
or UO_2801 (O_2801,N_24904,N_23879);
or UO_2802 (O_2802,N_24627,N_24230);
nor UO_2803 (O_2803,N_24667,N_23850);
or UO_2804 (O_2804,N_24443,N_24218);
xnor UO_2805 (O_2805,N_24017,N_24556);
and UO_2806 (O_2806,N_24902,N_24707);
and UO_2807 (O_2807,N_24929,N_24112);
nor UO_2808 (O_2808,N_24099,N_23994);
nand UO_2809 (O_2809,N_24267,N_24850);
or UO_2810 (O_2810,N_24802,N_24588);
nand UO_2811 (O_2811,N_24445,N_24402);
or UO_2812 (O_2812,N_24824,N_24106);
nand UO_2813 (O_2813,N_24952,N_24324);
nor UO_2814 (O_2814,N_24488,N_24977);
and UO_2815 (O_2815,N_23841,N_24149);
nand UO_2816 (O_2816,N_24816,N_24218);
xor UO_2817 (O_2817,N_24506,N_23898);
or UO_2818 (O_2818,N_24048,N_24246);
and UO_2819 (O_2819,N_24052,N_24426);
nor UO_2820 (O_2820,N_24503,N_24925);
or UO_2821 (O_2821,N_24552,N_23945);
xnor UO_2822 (O_2822,N_24093,N_24457);
xnor UO_2823 (O_2823,N_24554,N_24710);
nor UO_2824 (O_2824,N_23754,N_23886);
nand UO_2825 (O_2825,N_23820,N_23860);
and UO_2826 (O_2826,N_24410,N_24754);
and UO_2827 (O_2827,N_24828,N_24410);
nor UO_2828 (O_2828,N_24801,N_24462);
xor UO_2829 (O_2829,N_24262,N_24665);
nor UO_2830 (O_2830,N_24800,N_24503);
and UO_2831 (O_2831,N_24164,N_24042);
or UO_2832 (O_2832,N_24542,N_24528);
and UO_2833 (O_2833,N_24281,N_24810);
or UO_2834 (O_2834,N_24725,N_24439);
nor UO_2835 (O_2835,N_24491,N_24647);
nand UO_2836 (O_2836,N_24667,N_24725);
nand UO_2837 (O_2837,N_24357,N_24257);
xor UO_2838 (O_2838,N_24588,N_23801);
or UO_2839 (O_2839,N_24432,N_24454);
and UO_2840 (O_2840,N_24043,N_24381);
nand UO_2841 (O_2841,N_24630,N_24095);
nand UO_2842 (O_2842,N_23950,N_24396);
xor UO_2843 (O_2843,N_23805,N_23995);
nor UO_2844 (O_2844,N_24499,N_24786);
xnor UO_2845 (O_2845,N_24516,N_23796);
nor UO_2846 (O_2846,N_24003,N_24896);
and UO_2847 (O_2847,N_24385,N_24696);
nand UO_2848 (O_2848,N_24293,N_24588);
nor UO_2849 (O_2849,N_24193,N_24680);
xor UO_2850 (O_2850,N_24406,N_24945);
nand UO_2851 (O_2851,N_24030,N_23942);
and UO_2852 (O_2852,N_24765,N_24282);
and UO_2853 (O_2853,N_24056,N_24672);
nand UO_2854 (O_2854,N_24047,N_23975);
nand UO_2855 (O_2855,N_24755,N_24679);
and UO_2856 (O_2856,N_24877,N_24803);
xnor UO_2857 (O_2857,N_24962,N_24684);
nor UO_2858 (O_2858,N_24603,N_24637);
or UO_2859 (O_2859,N_24233,N_24089);
xnor UO_2860 (O_2860,N_24219,N_24300);
nand UO_2861 (O_2861,N_23828,N_23930);
and UO_2862 (O_2862,N_24650,N_24906);
nand UO_2863 (O_2863,N_24061,N_24223);
nand UO_2864 (O_2864,N_24474,N_24340);
nand UO_2865 (O_2865,N_24563,N_24790);
xor UO_2866 (O_2866,N_23809,N_23888);
and UO_2867 (O_2867,N_24092,N_24009);
nor UO_2868 (O_2868,N_24820,N_23949);
nor UO_2869 (O_2869,N_24281,N_24037);
or UO_2870 (O_2870,N_23940,N_24391);
and UO_2871 (O_2871,N_24599,N_24635);
and UO_2872 (O_2872,N_24196,N_24672);
or UO_2873 (O_2873,N_24226,N_24914);
nand UO_2874 (O_2874,N_24904,N_24271);
xor UO_2875 (O_2875,N_24452,N_24924);
or UO_2876 (O_2876,N_23881,N_24415);
nor UO_2877 (O_2877,N_24511,N_24828);
or UO_2878 (O_2878,N_24615,N_24287);
or UO_2879 (O_2879,N_24180,N_24498);
xor UO_2880 (O_2880,N_24522,N_24949);
xnor UO_2881 (O_2881,N_24228,N_24918);
xnor UO_2882 (O_2882,N_23989,N_24473);
nand UO_2883 (O_2883,N_24281,N_24528);
nand UO_2884 (O_2884,N_24597,N_23911);
xor UO_2885 (O_2885,N_24538,N_23900);
and UO_2886 (O_2886,N_24833,N_24247);
xnor UO_2887 (O_2887,N_24079,N_24402);
nor UO_2888 (O_2888,N_24853,N_24574);
xor UO_2889 (O_2889,N_24124,N_24134);
nand UO_2890 (O_2890,N_24154,N_24619);
xnor UO_2891 (O_2891,N_24634,N_24239);
and UO_2892 (O_2892,N_24300,N_24057);
or UO_2893 (O_2893,N_23879,N_24601);
nor UO_2894 (O_2894,N_24778,N_24480);
xnor UO_2895 (O_2895,N_24629,N_24961);
xnor UO_2896 (O_2896,N_24951,N_24784);
or UO_2897 (O_2897,N_24331,N_24037);
and UO_2898 (O_2898,N_23798,N_23976);
xnor UO_2899 (O_2899,N_24176,N_23942);
xnor UO_2900 (O_2900,N_24108,N_23921);
and UO_2901 (O_2901,N_24725,N_24411);
xor UO_2902 (O_2902,N_24907,N_23992);
nor UO_2903 (O_2903,N_24350,N_24491);
xor UO_2904 (O_2904,N_24401,N_24777);
nor UO_2905 (O_2905,N_24393,N_23994);
xnor UO_2906 (O_2906,N_24066,N_24699);
nand UO_2907 (O_2907,N_23968,N_23819);
or UO_2908 (O_2908,N_24446,N_24271);
and UO_2909 (O_2909,N_23850,N_23857);
or UO_2910 (O_2910,N_23784,N_24431);
xor UO_2911 (O_2911,N_24379,N_23832);
xor UO_2912 (O_2912,N_24274,N_24336);
nor UO_2913 (O_2913,N_24352,N_24222);
nand UO_2914 (O_2914,N_24078,N_24552);
nand UO_2915 (O_2915,N_24926,N_24377);
and UO_2916 (O_2916,N_24556,N_24162);
nor UO_2917 (O_2917,N_24619,N_24756);
xor UO_2918 (O_2918,N_24854,N_23852);
or UO_2919 (O_2919,N_23938,N_24214);
nand UO_2920 (O_2920,N_24776,N_24535);
xor UO_2921 (O_2921,N_24709,N_23947);
nand UO_2922 (O_2922,N_24984,N_24564);
or UO_2923 (O_2923,N_24367,N_24874);
xnor UO_2924 (O_2924,N_24722,N_24272);
nor UO_2925 (O_2925,N_23811,N_24726);
xnor UO_2926 (O_2926,N_23969,N_24796);
xor UO_2927 (O_2927,N_23821,N_24183);
xnor UO_2928 (O_2928,N_24254,N_24117);
nand UO_2929 (O_2929,N_23924,N_24061);
nand UO_2930 (O_2930,N_24439,N_24871);
xnor UO_2931 (O_2931,N_24042,N_23911);
xnor UO_2932 (O_2932,N_24050,N_24332);
or UO_2933 (O_2933,N_24890,N_24784);
xor UO_2934 (O_2934,N_23891,N_24227);
nand UO_2935 (O_2935,N_24768,N_24200);
nand UO_2936 (O_2936,N_24664,N_24006);
nor UO_2937 (O_2937,N_24099,N_24961);
or UO_2938 (O_2938,N_23857,N_23825);
xor UO_2939 (O_2939,N_24467,N_24108);
and UO_2940 (O_2940,N_24328,N_24355);
xnor UO_2941 (O_2941,N_24168,N_24241);
nor UO_2942 (O_2942,N_24213,N_24618);
nor UO_2943 (O_2943,N_24994,N_24173);
and UO_2944 (O_2944,N_24426,N_24141);
nand UO_2945 (O_2945,N_24557,N_24254);
xor UO_2946 (O_2946,N_24303,N_24068);
or UO_2947 (O_2947,N_24175,N_24808);
and UO_2948 (O_2948,N_24760,N_24691);
or UO_2949 (O_2949,N_23840,N_24820);
and UO_2950 (O_2950,N_24365,N_24097);
or UO_2951 (O_2951,N_24545,N_23810);
nand UO_2952 (O_2952,N_24839,N_24893);
xnor UO_2953 (O_2953,N_24824,N_24196);
nand UO_2954 (O_2954,N_24267,N_24430);
and UO_2955 (O_2955,N_23804,N_24083);
and UO_2956 (O_2956,N_24161,N_23940);
nor UO_2957 (O_2957,N_24791,N_24280);
nor UO_2958 (O_2958,N_23789,N_24807);
nor UO_2959 (O_2959,N_24252,N_24112);
nand UO_2960 (O_2960,N_24794,N_24462);
nor UO_2961 (O_2961,N_24062,N_24223);
xnor UO_2962 (O_2962,N_24741,N_23944);
or UO_2963 (O_2963,N_24793,N_24553);
nor UO_2964 (O_2964,N_23882,N_24327);
xor UO_2965 (O_2965,N_24804,N_24454);
and UO_2966 (O_2966,N_24336,N_24549);
nor UO_2967 (O_2967,N_24631,N_24724);
xnor UO_2968 (O_2968,N_23977,N_24459);
or UO_2969 (O_2969,N_24015,N_24595);
nor UO_2970 (O_2970,N_24201,N_24868);
nor UO_2971 (O_2971,N_24869,N_24749);
nor UO_2972 (O_2972,N_24491,N_23814);
or UO_2973 (O_2973,N_24252,N_24132);
nand UO_2974 (O_2974,N_24621,N_24460);
and UO_2975 (O_2975,N_24222,N_24399);
nand UO_2976 (O_2976,N_24726,N_24316);
xor UO_2977 (O_2977,N_23834,N_24751);
nand UO_2978 (O_2978,N_24634,N_24317);
or UO_2979 (O_2979,N_23824,N_23750);
or UO_2980 (O_2980,N_23817,N_24698);
xor UO_2981 (O_2981,N_24892,N_23958);
xor UO_2982 (O_2982,N_24776,N_24823);
and UO_2983 (O_2983,N_24883,N_24850);
xor UO_2984 (O_2984,N_24032,N_24601);
xnor UO_2985 (O_2985,N_24219,N_24038);
and UO_2986 (O_2986,N_23890,N_24143);
and UO_2987 (O_2987,N_24943,N_24441);
nor UO_2988 (O_2988,N_24061,N_24744);
xor UO_2989 (O_2989,N_24890,N_24079);
and UO_2990 (O_2990,N_24978,N_24109);
nor UO_2991 (O_2991,N_24651,N_24051);
nand UO_2992 (O_2992,N_24632,N_24299);
or UO_2993 (O_2993,N_23813,N_24749);
xor UO_2994 (O_2994,N_23908,N_24730);
or UO_2995 (O_2995,N_23962,N_24783);
or UO_2996 (O_2996,N_23914,N_24045);
nand UO_2997 (O_2997,N_23885,N_24081);
xor UO_2998 (O_2998,N_24856,N_24477);
nand UO_2999 (O_2999,N_24642,N_24711);
endmodule