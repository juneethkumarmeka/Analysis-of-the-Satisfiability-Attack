module basic_1500_15000_2000_3_levels_1xor_3(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10003,N_10005,N_10007,N_10008,N_10010,N_10011,N_10012,N_10014,N_10015,N_10016,N_10017,N_10018,N_10020,N_10022,N_10023,N_10025,N_10027,N_10028,N_10029,N_10031,N_10032,N_10033,N_10034,N_10036,N_10037,N_10039,N_10040,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10051,N_10053,N_10054,N_10056,N_10060,N_10062,N_10063,N_10064,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10078,N_10079,N_10080,N_10082,N_10084,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10109,N_10111,N_10112,N_10113,N_10115,N_10116,N_10117,N_10118,N_10119,N_10121,N_10122,N_10123,N_10124,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10154,N_10155,N_10156,N_10157,N_10158,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10169,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10178,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10201,N_10203,N_10204,N_10205,N_10206,N_10208,N_10209,N_10211,N_10212,N_10213,N_10215,N_10216,N_10217,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10230,N_10231,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10241,N_10242,N_10243,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10254,N_10255,N_10257,N_10258,N_10259,N_10260,N_10261,N_10263,N_10264,N_10266,N_10269,N_10271,N_10272,N_10273,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10290,N_10291,N_10292,N_10294,N_10295,N_10297,N_10298,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10309,N_10310,N_10311,N_10312,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10321,N_10322,N_10323,N_10324,N_10325,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10348,N_10349,N_10351,N_10352,N_10353,N_10354,N_10356,N_10357,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10397,N_10398,N_10399,N_10401,N_10402,N_10404,N_10405,N_10406,N_10408,N_10410,N_10411,N_10412,N_10413,N_10414,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10424,N_10425,N_10426,N_10427,N_10428,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10439,N_10440,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10450,N_10451,N_10452,N_10453,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10464,N_10465,N_10467,N_10470,N_10471,N_10472,N_10474,N_10475,N_10477,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10518,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10529,N_10530,N_10531,N_10532,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10561,N_10562,N_10564,N_10566,N_10567,N_10568,N_10571,N_10572,N_10574,N_10575,N_10577,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10612,N_10614,N_10615,N_10616,N_10617,N_10619,N_10620,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10652,N_10654,N_10655,N_10656,N_10659,N_10661,N_10664,N_10666,N_10667,N_10668,N_10669,N_10670,N_10673,N_10674,N_10676,N_10677,N_10678,N_10679,N_10681,N_10683,N_10684,N_10685,N_10686,N_10687,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10717,N_10721,N_10722,N_10723,N_10724,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10737,N_10738,N_10739,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10771,N_10772,N_10774,N_10776,N_10778,N_10779,N_10780,N_10781,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10801,N_10803,N_10804,N_10805,N_10806,N_10808,N_10810,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10820,N_10821,N_10822,N_10823,N_10827,N_10831,N_10832,N_10833,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10844,N_10846,N_10847,N_10848,N_10849,N_10850,N_10852,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10862,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10871,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10893,N_10894,N_10895,N_10896,N_10897,N_10900,N_10901,N_10903,N_10904,N_10905,N_10907,N_10908,N_10909,N_10911,N_10912,N_10913,N_10914,N_10915,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10924,N_10925,N_10926,N_10929,N_10930,N_10932,N_10933,N_10934,N_10935,N_10936,N_10938,N_10941,N_10942,N_10944,N_10945,N_10947,N_10948,N_10949,N_10950,N_10952,N_10953,N_10955,N_10956,N_10957,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10968,N_10969,N_10970,N_10971,N_10972,N_10975,N_10976,N_10977,N_10978,N_10980,N_10981,N_10982,N_10983,N_10984,N_10988,N_10989,N_10991,N_10992,N_10993,N_10995,N_10996,N_10997,N_10998,N_10999,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11047,N_11048,N_11050,N_11051,N_11052,N_11053,N_11054,N_11056,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11077,N_11078,N_11079,N_11080,N_11086,N_11087,N_11089,N_11090,N_11093,N_11094,N_11096,N_11097,N_11098,N_11099,N_11100,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11110,N_11112,N_11114,N_11116,N_11117,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11131,N_11132,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11162,N_11165,N_11166,N_11167,N_11169,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11190,N_11191,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11202,N_11203,N_11204,N_11206,N_11208,N_11210,N_11211,N_11212,N_11213,N_11215,N_11216,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11230,N_11231,N_11232,N_11233,N_11234,N_11237,N_11239,N_11240,N_11241,N_11243,N_11244,N_11246,N_11247,N_11249,N_11251,N_11252,N_11253,N_11254,N_11256,N_11257,N_11258,N_11259,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11291,N_11292,N_11293,N_11294,N_11296,N_11297,N_11298,N_11299,N_11300,N_11302,N_11303,N_11304,N_11305,N_11306,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11331,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11356,N_11357,N_11358,N_11359,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11387,N_11388,N_11389,N_11391,N_11392,N_11394,N_11395,N_11396,N_11397,N_11398,N_11400,N_11402,N_11403,N_11404,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11420,N_11421,N_11422,N_11423,N_11427,N_11428,N_11430,N_11431,N_11432,N_11433,N_11434,N_11437,N_11438,N_11439,N_11440,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11454,N_11456,N_11457,N_11459,N_11460,N_11461,N_11462,N_11463,N_11465,N_11466,N_11467,N_11470,N_11472,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11483,N_11484,N_11486,N_11488,N_11489,N_11490,N_11493,N_11494,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11515,N_11516,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11540,N_11541,N_11542,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11563,N_11564,N_11565,N_11566,N_11567,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11592,N_11594,N_11595,N_11596,N_11597,N_11599,N_11600,N_11601,N_11604,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11645,N_11646,N_11647,N_11648,N_11649,N_11651,N_11652,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11673,N_11674,N_11675,N_11676,N_11678,N_11679,N_11680,N_11681,N_11682,N_11686,N_11687,N_11688,N_11691,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11701,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11722,N_11726,N_11727,N_11731,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11742,N_11743,N_11744,N_11745,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11762,N_11763,N_11764,N_11765,N_11766,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11786,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11820,N_11821,N_11823,N_11824,N_11825,N_11826,N_11829,N_11830,N_11832,N_11833,N_11835,N_11836,N_11837,N_11838,N_11839,N_11842,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11894,N_11895,N_11897,N_11898,N_11900,N_11901,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11916,N_11917,N_11918,N_11920,N_11922,N_11923,N_11924,N_11926,N_11928,N_11930,N_11931,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11942,N_11944,N_11945,N_11946,N_11948,N_11949,N_11950,N_11954,N_11955,N_11956,N_11957,N_11959,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11970,N_11971,N_11972,N_11974,N_11976,N_11977,N_11978,N_11979,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11990,N_11991,N_11992,N_11994,N_11995,N_11996,N_11998,N_11999,N_12000,N_12002,N_12003,N_12004,N_12006,N_12007,N_12008,N_12009,N_12010,N_12012,N_12013,N_12014,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12041,N_12042,N_12043,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12069,N_12070,N_12071,N_12073,N_12074,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12087,N_12088,N_12089,N_12091,N_12092,N_12093,N_12094,N_12095,N_12097,N_12098,N_12099,N_12101,N_12102,N_12103,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12113,N_12114,N_12118,N_12119,N_12120,N_12121,N_12122,N_12124,N_12125,N_12126,N_12128,N_12129,N_12130,N_12132,N_12133,N_12134,N_12135,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12149,N_12150,N_12151,N_12152,N_12153,N_12155,N_12156,N_12157,N_12159,N_12160,N_12161,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12191,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12200,N_12201,N_12203,N_12205,N_12206,N_12207,N_12209,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12219,N_12220,N_12221,N_12223,N_12225,N_12226,N_12227,N_12228,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12238,N_12239,N_12240,N_12241,N_12243,N_12245,N_12246,N_12247,N_12248,N_12250,N_12251,N_12253,N_12254,N_12255,N_12256,N_12257,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12269,N_12270,N_12272,N_12273,N_12274,N_12275,N_12276,N_12278,N_12280,N_12281,N_12282,N_12285,N_12286,N_12288,N_12289,N_12290,N_12291,N_12292,N_12294,N_12296,N_12297,N_12298,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12307,N_12308,N_12309,N_12310,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12319,N_12320,N_12322,N_12323,N_12324,N_12325,N_12326,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12339,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12373,N_12375,N_12377,N_12380,N_12381,N_12382,N_12383,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12396,N_12397,N_12398,N_12399,N_12401,N_12402,N_12403,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12435,N_12436,N_12438,N_12439,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12450,N_12451,N_12452,N_12453,N_12454,N_12456,N_12457,N_12459,N_12460,N_12461,N_12462,N_12464,N_12465,N_12466,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12479,N_12480,N_12481,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12490,N_12491,N_12492,N_12494,N_12495,N_12496,N_12497,N_12500,N_12502,N_12503,N_12504,N_12505,N_12506,N_12508,N_12510,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12528,N_12529,N_12530,N_12531,N_12533,N_12535,N_12536,N_12537,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12552,N_12553,N_12555,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12568,N_12569,N_12570,N_12571,N_12572,N_12574,N_12576,N_12579,N_12582,N_12583,N_12584,N_12585,N_12587,N_12588,N_12589,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12606,N_12607,N_12609,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12635,N_12636,N_12638,N_12639,N_12641,N_12642,N_12643,N_12644,N_12645,N_12647,N_12649,N_12650,N_12651,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12673,N_12674,N_12675,N_12676,N_12679,N_12680,N_12681,N_12683,N_12686,N_12687,N_12688,N_12689,N_12691,N_12693,N_12694,N_12695,N_12696,N_12698,N_12699,N_12701,N_12702,N_12704,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12716,N_12717,N_12718,N_12720,N_12724,N_12725,N_12726,N_12727,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12767,N_12768,N_12770,N_12771,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12790,N_12791,N_12792,N_12794,N_12796,N_12797,N_12799,N_12800,N_12802,N_12803,N_12804,N_12805,N_12806,N_12808,N_12810,N_12811,N_12812,N_12813,N_12814,N_12816,N_12817,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12839,N_12840,N_12841,N_12842,N_12844,N_12845,N_12846,N_12847,N_12848,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12865,N_12866,N_12868,N_12870,N_12872,N_12873,N_12874,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12888,N_12889,N_12891,N_12892,N_12893,N_12896,N_12897,N_12900,N_12901,N_12902,N_12903,N_12905,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12925,N_12926,N_12927,N_12928,N_12930,N_12932,N_12933,N_12934,N_12938,N_12939,N_12940,N_12942,N_12943,N_12944,N_12945,N_12947,N_12948,N_12949,N_12950,N_12952,N_12953,N_12954,N_12955,N_12956,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12966,N_12967,N_12968,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12979,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12994,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13011,N_13012,N_13013,N_13015,N_13016,N_13017,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13036,N_13037,N_13039,N_13040,N_13041,N_13042,N_13044,N_13045,N_13047,N_13048,N_13050,N_13052,N_13053,N_13054,N_13056,N_13057,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13067,N_13068,N_13069,N_13070,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13087,N_13089,N_13090,N_13091,N_13093,N_13097,N_13098,N_13099,N_13100,N_13101,N_13103,N_13104,N_13105,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13141,N_13142,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13162,N_13163,N_13164,N_13165,N_13168,N_13170,N_13171,N_13173,N_13174,N_13175,N_13177,N_13179,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13208,N_13210,N_13212,N_13213,N_13214,N_13216,N_13218,N_13220,N_13226,N_13227,N_13228,N_13229,N_13231,N_13232,N_13233,N_13235,N_13236,N_13238,N_13239,N_13241,N_13243,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13261,N_13263,N_13264,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13276,N_13278,N_13279,N_13280,N_13281,N_13282,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13297,N_13298,N_13299,N_13300,N_13302,N_13303,N_13304,N_13308,N_13310,N_13312,N_13314,N_13316,N_13317,N_13318,N_13319,N_13321,N_13322,N_13323,N_13325,N_13327,N_13328,N_13329,N_13330,N_13331,N_13335,N_13336,N_13337,N_13338,N_13340,N_13342,N_13343,N_13345,N_13346,N_13347,N_13349,N_13350,N_13351,N_13353,N_13354,N_13355,N_13356,N_13357,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13373,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13384,N_13385,N_13386,N_13387,N_13389,N_13390,N_13391,N_13392,N_13395,N_13399,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13436,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13450,N_13451,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13480,N_13482,N_13483,N_13485,N_13487,N_13488,N_13489,N_13490,N_13491,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13517,N_13518,N_13519,N_13521,N_13522,N_13523,N_13524,N_13525,N_13527,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13536,N_13538,N_13540,N_13544,N_13545,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13580,N_13581,N_13584,N_13587,N_13588,N_13589,N_13590,N_13592,N_13593,N_13594,N_13595,N_13597,N_13601,N_13602,N_13603,N_13604,N_13605,N_13608,N_13609,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13632,N_13633,N_13636,N_13637,N_13638,N_13639,N_13640,N_13642,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13651,N_13652,N_13653,N_13654,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13678,N_13680,N_13681,N_13682,N_13683,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13694,N_13695,N_13697,N_13698,N_13699,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13713,N_13714,N_13715,N_13718,N_13719,N_13720,N_13721,N_13722,N_13725,N_13726,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13753,N_13754,N_13755,N_13756,N_13757,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13770,N_13771,N_13772,N_13774,N_13775,N_13778,N_13779,N_13781,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13792,N_13795,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13816,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13849,N_13851,N_13852,N_13853,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13867,N_13868,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13894,N_13895,N_13896,N_13897,N_13899,N_13901,N_13902,N_13903,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13958,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13971,N_13972,N_13973,N_13975,N_13976,N_13977,N_13979,N_13980,N_13981,N_13982,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13991,N_13993,N_13994,N_13996,N_13997,N_13998,N_13999,N_14000,N_14002,N_14003,N_14004,N_14005,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14041,N_14042,N_14043,N_14044,N_14046,N_14047,N_14048,N_14050,N_14052,N_14053,N_14054,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14063,N_14065,N_14066,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14079,N_14080,N_14081,N_14082,N_14084,N_14085,N_14086,N_14087,N_14088,N_14090,N_14092,N_14094,N_14095,N_14096,N_14097,N_14099,N_14100,N_14102,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14125,N_14126,N_14127,N_14128,N_14130,N_14131,N_14133,N_14134,N_14137,N_14138,N_14140,N_14142,N_14144,N_14145,N_14146,N_14148,N_14149,N_14151,N_14152,N_14153,N_14155,N_14156,N_14157,N_14159,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14170,N_14171,N_14173,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14187,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14231,N_14232,N_14233,N_14234,N_14236,N_14237,N_14238,N_14239,N_14241,N_14242,N_14243,N_14244,N_14245,N_14247,N_14248,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14266,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14283,N_14284,N_14285,N_14286,N_14288,N_14289,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14298,N_14299,N_14300,N_14301,N_14303,N_14304,N_14305,N_14306,N_14307,N_14309,N_14310,N_14311,N_14312,N_14313,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14327,N_14328,N_14329,N_14330,N_14332,N_14333,N_14335,N_14337,N_14339,N_14340,N_14341,N_14343,N_14344,N_14345,N_14346,N_14348,N_14350,N_14351,N_14352,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14387,N_14388,N_14389,N_14391,N_14392,N_14394,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14455,N_14456,N_14457,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14502,N_14503,N_14504,N_14506,N_14507,N_14508,N_14511,N_14512,N_14515,N_14516,N_14517,N_14518,N_14521,N_14522,N_14523,N_14525,N_14526,N_14527,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14539,N_14540,N_14542,N_14543,N_14545,N_14546,N_14547,N_14548,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14559,N_14561,N_14563,N_14564,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14584,N_14586,N_14587,N_14588,N_14590,N_14592,N_14594,N_14595,N_14596,N_14597,N_14599,N_14600,N_14602,N_14603,N_14605,N_14606,N_14607,N_14609,N_14610,N_14611,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14621,N_14622,N_14624,N_14625,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14642,N_14644,N_14645,N_14646,N_14647,N_14648,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14659,N_14660,N_14661,N_14663,N_14664,N_14665,N_14667,N_14669,N_14670,N_14672,N_14673,N_14674,N_14675,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14717,N_14718,N_14719,N_14720,N_14721,N_14723,N_14724,N_14725,N_14727,N_14728,N_14729,N_14730,N_14732,N_14734,N_14737,N_14738,N_14741,N_14742,N_14743,N_14745,N_14746,N_14748,N_14749,N_14750,N_14752,N_14753,N_14754,N_14758,N_14759,N_14760,N_14761,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14771,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14789,N_14790,N_14791,N_14792,N_14794,N_14795,N_14796,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14807,N_14808,N_14809,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14818,N_14819,N_14820,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14854,N_14855,N_14857,N_14858,N_14860,N_14861,N_14862,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14878,N_14879,N_14881,N_14882,N_14885,N_14886,N_14887,N_14888,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14924,N_14925,N_14926,N_14927,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14940,N_14942,N_14943,N_14946,N_14947,N_14948,N_14949,N_14950,N_14952,N_14953,N_14956,N_14957,N_14958,N_14959,N_14961,N_14962,N_14965,N_14966,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14987,N_14988,N_14989,N_14990,N_14991,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999;
or U0 (N_0,In_1315,In_895);
or U1 (N_1,In_1041,In_1300);
nand U2 (N_2,In_1326,In_664);
or U3 (N_3,In_260,In_598);
and U4 (N_4,In_1174,In_763);
nor U5 (N_5,In_175,In_819);
and U6 (N_6,In_428,In_1153);
and U7 (N_7,In_1022,In_731);
nand U8 (N_8,In_959,In_810);
nor U9 (N_9,In_513,In_347);
nor U10 (N_10,In_764,In_159);
or U11 (N_11,In_1206,In_683);
xor U12 (N_12,In_267,In_326);
and U13 (N_13,In_775,In_935);
xnor U14 (N_14,In_710,In_1016);
or U15 (N_15,In_658,In_135);
nand U16 (N_16,In_1230,In_336);
nand U17 (N_17,In_491,In_1444);
nor U18 (N_18,In_1056,In_1098);
nor U19 (N_19,In_863,In_765);
nand U20 (N_20,In_1448,In_784);
and U21 (N_21,In_606,In_1467);
or U22 (N_22,In_1148,In_484);
and U23 (N_23,In_264,In_91);
or U24 (N_24,In_348,In_406);
or U25 (N_25,In_463,In_649);
or U26 (N_26,In_1301,In_704);
nand U27 (N_27,In_1078,In_1119);
or U28 (N_28,In_1049,In_423);
or U29 (N_29,In_609,In_651);
nand U30 (N_30,In_201,In_1442);
nand U31 (N_31,In_542,In_750);
or U32 (N_32,In_377,In_431);
and U33 (N_33,In_1297,In_565);
or U34 (N_34,In_562,In_953);
and U35 (N_35,In_945,In_1062);
nor U36 (N_36,In_320,In_1152);
and U37 (N_37,In_602,In_1325);
or U38 (N_38,In_1479,In_712);
and U39 (N_39,In_1350,In_174);
nor U40 (N_40,In_1238,In_772);
and U41 (N_41,In_1047,In_1172);
nor U42 (N_42,In_1007,In_1169);
or U43 (N_43,In_982,In_586);
and U44 (N_44,In_1494,In_939);
and U45 (N_45,In_1406,In_1284);
and U46 (N_46,In_1142,In_70);
or U47 (N_47,In_1242,In_405);
nand U48 (N_48,In_902,In_655);
and U49 (N_49,In_448,In_202);
nand U50 (N_50,In_900,In_1082);
nor U51 (N_51,In_497,In_854);
nand U52 (N_52,In_725,In_891);
nor U53 (N_53,In_908,In_1211);
and U54 (N_54,In_1304,In_340);
and U55 (N_55,In_873,In_862);
nand U56 (N_56,In_691,In_1313);
nor U57 (N_57,In_1283,In_1031);
or U58 (N_58,In_138,In_1351);
nand U59 (N_59,In_1255,In_1194);
nand U60 (N_60,In_250,In_384);
nand U61 (N_61,In_673,In_608);
or U62 (N_62,In_830,In_1394);
and U63 (N_63,In_1055,In_7);
and U64 (N_64,In_1319,In_1088);
and U65 (N_65,In_86,In_870);
or U66 (N_66,In_590,In_1190);
nor U67 (N_67,In_112,In_919);
or U68 (N_68,In_997,In_697);
and U69 (N_69,In_514,In_989);
or U70 (N_70,In_1435,In_426);
nand U71 (N_71,In_196,In_748);
xor U72 (N_72,In_753,In_1258);
nor U73 (N_73,In_1265,In_1376);
nor U74 (N_74,In_285,In_1468);
or U75 (N_75,In_479,In_1495);
or U76 (N_76,In_550,In_1220);
and U77 (N_77,In_367,In_469);
and U78 (N_78,In_686,In_1015);
or U79 (N_79,In_1484,In_1424);
and U80 (N_80,In_946,In_1187);
and U81 (N_81,In_847,In_1084);
xor U82 (N_82,In_852,In_1359);
nand U83 (N_83,In_229,In_1093);
nand U84 (N_84,In_1491,In_493);
nor U85 (N_85,In_918,In_478);
or U86 (N_86,In_409,In_780);
nor U87 (N_87,In_523,In_95);
and U88 (N_88,In_884,In_587);
and U89 (N_89,In_1048,In_848);
and U90 (N_90,In_793,In_975);
nor U91 (N_91,In_1485,In_1438);
or U92 (N_92,In_886,In_318);
nor U93 (N_93,In_172,In_818);
or U94 (N_94,In_1369,In_752);
or U95 (N_95,In_857,In_948);
nor U96 (N_96,In_841,In_532);
nand U97 (N_97,In_16,In_932);
nor U98 (N_98,In_619,In_165);
nand U99 (N_99,In_1458,In_443);
and U100 (N_100,In_1499,In_1449);
nor U101 (N_101,In_199,In_114);
or U102 (N_102,In_694,In_218);
nand U103 (N_103,In_1223,In_677);
and U104 (N_104,In_999,In_1289);
and U105 (N_105,In_287,In_966);
nand U106 (N_106,In_1009,In_432);
or U107 (N_107,In_226,In_351);
nor U108 (N_108,In_1116,In_998);
or U109 (N_109,In_223,In_526);
nor U110 (N_110,In_552,In_8);
nor U111 (N_111,In_976,In_450);
nor U112 (N_112,In_1236,In_1332);
nor U113 (N_113,In_1307,In_1488);
and U114 (N_114,In_692,In_158);
nor U115 (N_115,In_518,In_113);
nand U116 (N_116,In_99,In_599);
or U117 (N_117,In_420,In_482);
nor U118 (N_118,In_75,In_1147);
and U119 (N_119,In_54,In_1276);
xnor U120 (N_120,In_1034,In_881);
nor U121 (N_121,In_1447,In_3);
or U122 (N_122,In_1043,In_715);
and U123 (N_123,In_1375,In_4);
nand U124 (N_124,In_992,In_475);
nand U125 (N_125,In_883,In_719);
nor U126 (N_126,In_676,In_1004);
nor U127 (N_127,In_1161,In_1033);
nand U128 (N_128,In_500,In_706);
nand U129 (N_129,In_191,In_477);
xnor U130 (N_130,In_1329,In_779);
nor U131 (N_131,In_689,In_42);
or U132 (N_132,In_567,In_111);
or U133 (N_133,In_885,In_427);
nand U134 (N_134,In_417,In_1419);
and U135 (N_135,In_1186,In_1097);
or U136 (N_136,In_397,In_1069);
and U137 (N_137,In_1261,In_462);
nand U138 (N_138,In_290,In_211);
nor U139 (N_139,In_1165,In_1498);
or U140 (N_140,In_9,In_395);
and U141 (N_141,In_124,In_796);
or U142 (N_142,In_1130,In_659);
nand U143 (N_143,In_508,In_101);
and U144 (N_144,In_474,In_815);
nand U145 (N_145,In_1475,In_392);
xor U146 (N_146,In_802,In_820);
nor U147 (N_147,In_422,In_1270);
nand U148 (N_148,In_104,In_1094);
nor U149 (N_149,In_1331,In_528);
nor U150 (N_150,In_178,In_964);
and U151 (N_151,In_1286,In_566);
or U152 (N_152,In_1366,In_382);
or U153 (N_153,In_149,In_519);
or U154 (N_154,In_1459,In_315);
and U155 (N_155,In_1074,In_1476);
nand U156 (N_156,In_806,In_281);
and U157 (N_157,In_1020,In_321);
or U158 (N_158,In_1358,In_180);
or U159 (N_159,In_913,In_49);
nor U160 (N_160,In_1210,In_1387);
nor U161 (N_161,In_1235,In_546);
nor U162 (N_162,In_665,In_1149);
nand U163 (N_163,In_237,In_127);
and U164 (N_164,In_1285,In_17);
or U165 (N_165,In_301,In_1102);
and U166 (N_166,In_1288,In_132);
nand U167 (N_167,In_146,In_768);
nor U168 (N_168,In_615,In_632);
nor U169 (N_169,In_524,In_593);
and U170 (N_170,In_179,In_20);
nor U171 (N_171,In_440,In_205);
or U172 (N_172,In_912,In_1399);
nand U173 (N_173,In_574,In_1024);
or U174 (N_174,In_1477,In_369);
and U175 (N_175,In_208,In_1036);
nor U176 (N_176,In_152,In_168);
and U177 (N_177,In_1189,In_822);
or U178 (N_178,In_222,In_410);
or U179 (N_179,In_718,In_15);
nand U180 (N_180,In_1081,In_682);
or U181 (N_181,In_742,In_1170);
and U182 (N_182,In_960,In_693);
nand U183 (N_183,In_700,In_1405);
and U184 (N_184,In_72,In_483);
or U185 (N_185,In_1196,In_1341);
and U186 (N_186,In_1393,In_1143);
nand U187 (N_187,In_1002,In_594);
or U188 (N_188,In_128,In_404);
nand U189 (N_189,In_1386,In_1180);
nand U190 (N_190,In_849,In_1339);
nor U191 (N_191,In_961,In_769);
and U192 (N_192,In_639,In_995);
nor U193 (N_193,In_618,In_1355);
xor U194 (N_194,In_842,In_545);
nor U195 (N_195,In_327,In_65);
nor U196 (N_196,In_123,In_936);
or U197 (N_197,In_1374,In_538);
nor U198 (N_198,In_875,In_1079);
nand U199 (N_199,In_1184,In_286);
and U200 (N_200,In_1384,In_557);
nor U201 (N_201,In_248,In_1425);
and U202 (N_202,In_1185,In_931);
nor U203 (N_203,In_81,In_68);
and U204 (N_204,In_1240,In_1029);
and U205 (N_205,In_987,In_46);
nand U206 (N_206,In_2,In_1478);
nor U207 (N_207,In_84,In_1133);
and U208 (N_208,In_372,In_258);
nand U209 (N_209,In_511,In_1065);
nor U210 (N_210,In_1232,In_654);
nand U211 (N_211,In_1316,In_628);
or U212 (N_212,In_901,In_906);
nand U213 (N_213,In_687,In_343);
nor U214 (N_214,In_1416,In_394);
or U215 (N_215,In_838,In_1303);
or U216 (N_216,In_1352,In_1299);
nand U217 (N_217,In_192,In_1277);
or U218 (N_218,In_1112,In_1395);
and U219 (N_219,In_774,In_1431);
nand U220 (N_220,In_282,In_1259);
nand U221 (N_221,In_726,In_1001);
nand U222 (N_222,In_1204,In_636);
or U223 (N_223,In_588,In_487);
or U224 (N_224,In_176,In_798);
or U225 (N_225,In_903,In_579);
nand U226 (N_226,In_1076,In_1171);
nand U227 (N_227,In_1305,In_140);
nor U228 (N_228,In_302,In_1249);
or U229 (N_229,In_1096,In_1208);
and U230 (N_230,In_630,In_1377);
and U231 (N_231,In_207,In_121);
and U232 (N_232,In_454,In_1177);
or U233 (N_233,In_1492,In_1317);
xnor U234 (N_234,In_759,In_445);
nor U235 (N_235,In_845,In_306);
nand U236 (N_236,In_1335,In_1275);
nand U237 (N_237,In_537,In_74);
nor U238 (N_238,In_144,In_419);
and U239 (N_239,In_878,In_790);
nor U240 (N_240,In_1120,In_648);
or U241 (N_241,In_942,In_1465);
nor U242 (N_242,In_391,In_489);
and U243 (N_243,In_230,In_657);
xor U244 (N_244,In_1434,In_244);
nor U245 (N_245,In_224,In_283);
or U246 (N_246,In_332,In_106);
nor U247 (N_247,In_1136,In_5);
and U248 (N_248,In_621,In_671);
nor U249 (N_249,In_754,In_1163);
nand U250 (N_250,In_398,In_119);
and U251 (N_251,In_115,In_1312);
or U252 (N_252,In_167,In_596);
or U253 (N_253,In_293,In_559);
or U254 (N_254,In_696,In_1396);
or U255 (N_255,In_957,In_62);
and U256 (N_256,In_379,In_1080);
and U257 (N_257,In_1401,In_1101);
and U258 (N_258,In_52,In_241);
and U259 (N_259,In_698,In_1346);
or U260 (N_260,In_1349,In_929);
and U261 (N_261,In_1214,In_702);
and U262 (N_262,In_77,In_107);
nand U263 (N_263,In_368,In_1215);
and U264 (N_264,In_905,In_721);
nor U265 (N_265,In_217,In_766);
or U266 (N_266,In_613,In_699);
or U267 (N_267,In_1121,In_1390);
and U268 (N_268,In_642,In_187);
nand U269 (N_269,In_346,In_76);
or U270 (N_270,In_1450,In_751);
or U271 (N_271,In_154,In_1379);
or U272 (N_272,In_788,In_371);
nand U273 (N_273,In_451,In_564);
and U274 (N_274,In_303,In_43);
nor U275 (N_275,In_1113,In_1203);
and U276 (N_276,In_958,In_90);
nand U277 (N_277,In_1226,In_733);
or U278 (N_278,In_1432,In_344);
and U279 (N_279,In_1027,In_1042);
nor U280 (N_280,In_1179,In_341);
xnor U281 (N_281,In_360,In_1362);
nand U282 (N_282,In_1292,In_125);
or U283 (N_283,In_1426,In_1008);
nor U284 (N_284,In_446,In_47);
or U285 (N_285,In_1260,In_193);
nor U286 (N_286,In_517,In_109);
nand U287 (N_287,In_437,In_10);
nor U288 (N_288,In_416,In_1414);
nor U289 (N_289,In_380,In_1314);
nor U290 (N_290,In_1117,In_1252);
or U291 (N_291,In_1291,In_44);
and U292 (N_292,In_364,In_261);
or U293 (N_293,In_310,In_529);
or U294 (N_294,In_672,In_485);
or U295 (N_295,In_69,In_1181);
and U296 (N_296,In_79,In_1075);
or U297 (N_297,In_277,In_894);
and U298 (N_298,In_82,In_1445);
and U299 (N_299,In_582,In_1044);
nand U300 (N_300,In_108,In_746);
nor U301 (N_301,In_59,In_255);
and U302 (N_302,In_383,In_438);
nor U303 (N_303,In_647,In_19);
or U304 (N_304,In_269,In_137);
and U305 (N_305,In_316,In_745);
nand U306 (N_306,In_926,In_130);
nand U307 (N_307,In_743,In_401);
or U308 (N_308,In_1061,In_872);
nor U309 (N_309,In_661,In_840);
nand U310 (N_310,In_776,In_28);
nand U311 (N_311,In_1373,In_225);
nor U312 (N_312,In_1483,In_943);
nor U313 (N_313,In_257,In_203);
and U314 (N_314,In_24,In_947);
nor U315 (N_315,In_548,In_1493);
and U316 (N_316,In_359,In_1229);
or U317 (N_317,In_907,In_889);
nor U318 (N_318,In_1122,In_139);
and U319 (N_319,In_1473,In_50);
and U320 (N_320,In_853,In_1338);
and U321 (N_321,In_1237,In_956);
nand U322 (N_322,In_506,In_27);
and U323 (N_323,In_442,In_551);
or U324 (N_324,In_418,In_965);
and U325 (N_325,In_300,In_276);
or U326 (N_326,In_1057,In_1423);
and U327 (N_327,In_403,In_435);
or U328 (N_328,In_601,In_778);
nand U329 (N_329,In_861,In_89);
nor U330 (N_330,In_1248,In_415);
and U331 (N_331,In_399,In_805);
or U332 (N_332,In_262,In_323);
and U333 (N_333,In_85,In_324);
nand U334 (N_334,In_1410,In_1323);
nor U335 (N_335,In_543,In_1269);
and U336 (N_336,In_1453,In_1175);
or U337 (N_337,In_1137,In_195);
and U338 (N_338,In_1262,In_206);
nand U339 (N_339,In_1440,In_1274);
nor U340 (N_340,In_569,In_1404);
or U341 (N_341,In_1470,In_864);
and U342 (N_342,In_1272,In_735);
or U343 (N_343,In_337,In_298);
or U344 (N_344,In_429,In_1412);
and U345 (N_345,In_1216,In_614);
nand U346 (N_346,In_634,In_1217);
and U347 (N_347,In_1273,In_626);
and U348 (N_348,In_1000,In_339);
nor U349 (N_349,In_1134,In_1039);
nand U350 (N_350,In_539,In_1382);
and U351 (N_351,In_867,In_288);
nor U352 (N_352,In_1018,In_1025);
or U353 (N_353,In_1191,In_595);
or U354 (N_354,In_678,In_1253);
or U355 (N_355,In_194,In_1480);
or U356 (N_356,In_732,In_374);
or U357 (N_357,In_312,In_533);
nor U358 (N_358,In_877,In_1322);
and U359 (N_359,In_170,In_1158);
nor U360 (N_360,In_177,In_496);
or U361 (N_361,In_844,In_1132);
and U362 (N_362,In_684,In_1464);
and U363 (N_363,In_1234,In_1280);
or U364 (N_364,In_663,In_1095);
nor U365 (N_365,In_1392,In_461);
nand U366 (N_366,In_734,In_879);
and U367 (N_367,In_1462,In_204);
nand U368 (N_368,In_993,In_1363);
nand U369 (N_369,In_1115,In_994);
nand U370 (N_370,In_182,In_527);
and U371 (N_371,In_685,In_1348);
nand U372 (N_372,In_1228,In_279);
nor U373 (N_373,In_827,In_917);
nand U374 (N_374,In_974,In_1068);
nor U375 (N_375,In_826,In_728);
nand U376 (N_376,In_1311,In_30);
nand U377 (N_377,In_1037,In_1302);
xnor U378 (N_378,In_973,In_1193);
nand U379 (N_379,In_701,In_80);
and U380 (N_380,In_1360,In_717);
nand U381 (N_381,In_761,In_501);
and U382 (N_382,In_319,In_22);
or U383 (N_383,In_835,In_851);
or U384 (N_384,In_1114,In_888);
and U385 (N_385,In_629,In_1106);
and U386 (N_386,In_1086,In_812);
nand U387 (N_387,In_695,In_63);
nand U388 (N_388,In_858,In_307);
and U389 (N_389,In_39,In_892);
or U390 (N_390,In_755,In_235);
and U391 (N_391,In_280,In_171);
nand U392 (N_392,In_433,In_771);
nor U393 (N_393,In_1160,In_1298);
or U394 (N_394,In_57,In_60);
and U395 (N_395,In_295,In_1407);
and U396 (N_396,In_984,In_1245);
and U397 (N_397,In_985,In_1131);
or U398 (N_398,In_1013,In_591);
nand U399 (N_399,In_1053,In_1125);
or U400 (N_400,In_1365,In_83);
nor U401 (N_401,In_116,In_580);
nor U402 (N_402,In_14,In_928);
and U403 (N_403,In_762,In_21);
nand U404 (N_404,In_1085,In_1361);
or U405 (N_405,In_915,In_1135);
nand U406 (N_406,In_1466,In_1408);
and U407 (N_407,In_342,In_1012);
and U408 (N_408,In_1213,In_813);
nand U409 (N_409,In_1337,In_1422);
or U410 (N_410,In_744,In_1073);
nand U411 (N_411,In_1207,In_197);
or U412 (N_412,In_604,In_767);
xnor U413 (N_413,In_644,In_736);
nor U414 (N_414,In_625,In_273);
nor U415 (N_415,In_29,In_1231);
or U416 (N_416,In_713,In_944);
and U417 (N_417,In_1254,In_723);
nor U418 (N_418,In_716,In_373);
nor U419 (N_419,In_592,In_1188);
nor U420 (N_420,In_1345,In_93);
nor U421 (N_421,In_234,In_1411);
and U422 (N_422,In_708,In_1437);
nand U423 (N_423,In_1430,In_186);
or U424 (N_424,In_801,In_1328);
nor U425 (N_425,In_314,In_610);
or U426 (N_426,In_45,In_471);
nand U427 (N_427,In_979,In_617);
nand U428 (N_428,In_110,In_1105);
nor U429 (N_429,In_510,In_1138);
nand U430 (N_430,In_1461,In_652);
or U431 (N_431,In_183,In_345);
and U432 (N_432,In_1489,In_1308);
nand U433 (N_433,In_1107,In_1032);
nor U434 (N_434,In_1064,In_674);
or U435 (N_435,In_1343,In_646);
nand U436 (N_436,In_1071,In_834);
nor U437 (N_437,In_1296,In_624);
nor U438 (N_438,In_1318,In_898);
nor U439 (N_439,In_856,In_155);
nand U440 (N_440,In_690,In_758);
nand U441 (N_441,In_1388,In_335);
nor U442 (N_442,In_578,In_924);
nor U443 (N_443,In_773,In_583);
or U444 (N_444,In_232,In_536);
and U445 (N_445,In_738,In_737);
nor U446 (N_446,In_492,In_1336);
nor U447 (N_447,In_381,In_1221);
nand U448 (N_448,In_680,In_221);
and U449 (N_449,In_777,In_227);
or U450 (N_450,In_968,In_670);
or U451 (N_451,In_534,In_352);
and U452 (N_452,In_572,In_228);
and U453 (N_453,In_102,In_325);
nor U454 (N_454,In_933,In_893);
nand U455 (N_455,In_1108,In_1455);
nand U456 (N_456,In_741,In_1239);
nor U457 (N_457,In_498,In_328);
nor U458 (N_458,In_1290,In_874);
nand U459 (N_459,In_212,In_855);
nor U460 (N_460,In_272,In_1321);
nor U461 (N_461,In_505,In_268);
and U462 (N_462,In_525,In_430);
nor U463 (N_463,In_1327,In_794);
or U464 (N_464,In_1222,In_747);
and U465 (N_465,In_904,In_67);
nand U466 (N_466,In_486,In_923);
nor U467 (N_467,In_850,In_233);
nand U468 (N_468,In_1371,In_129);
or U469 (N_469,In_349,In_1278);
and U470 (N_470,In_955,In_407);
or U471 (N_471,In_464,In_434);
and U472 (N_472,In_64,In_1089);
nand U473 (N_473,In_720,In_58);
or U474 (N_474,In_876,In_1111);
nand U475 (N_475,In_1271,In_711);
or U476 (N_476,In_729,In_996);
nand U477 (N_477,In_1247,In_1168);
nand U478 (N_478,In_584,In_389);
nor U479 (N_479,In_1436,In_1486);
nand U480 (N_480,In_363,In_1159);
nand U481 (N_481,In_757,In_117);
nor U482 (N_482,In_236,In_1452);
or U483 (N_483,In_169,In_1287);
nand U484 (N_484,In_978,In_951);
nor U485 (N_485,In_843,In_1126);
nand U486 (N_486,In_357,In_504);
nor U487 (N_487,In_210,In_1209);
or U488 (N_488,In_916,In_1398);
or U489 (N_489,In_860,In_1167);
nand U490 (N_490,In_623,In_972);
or U491 (N_491,In_166,In_313);
or U492 (N_492,In_714,In_1344);
and U493 (N_493,In_1192,In_161);
or U494 (N_494,In_338,In_1118);
nand U495 (N_495,In_547,In_411);
nand U496 (N_496,In_1487,In_1205);
nand U497 (N_497,In_333,In_631);
nor U498 (N_498,In_162,In_88);
nor U499 (N_499,In_156,In_388);
and U500 (N_500,In_386,In_453);
or U501 (N_501,In_600,In_331);
nand U502 (N_502,In_760,In_322);
nand U503 (N_503,In_817,In_1026);
nand U504 (N_504,In_304,In_256);
nand U505 (N_505,In_105,In_1417);
nor U506 (N_506,In_25,In_950);
nor U507 (N_507,In_35,In_824);
nor U508 (N_508,In_378,In_914);
nor U509 (N_509,In_570,In_1282);
nand U510 (N_510,In_457,In_1166);
or U511 (N_511,In_266,In_96);
nand U512 (N_512,In_353,In_92);
nand U513 (N_513,In_553,In_456);
nor U514 (N_514,In_1257,In_1402);
and U515 (N_515,In_576,In_184);
nor U516 (N_516,In_531,In_1046);
or U517 (N_517,In_263,In_56);
nor U518 (N_518,In_274,In_589);
nor U519 (N_519,In_458,In_136);
and U520 (N_520,In_1227,In_18);
or U521 (N_521,In_1003,In_375);
nor U522 (N_522,In_153,In_1334);
nor U523 (N_523,In_560,In_1212);
nand U524 (N_524,In_781,In_78);
nor U525 (N_525,In_828,In_32);
nand U526 (N_526,In_616,In_1441);
nor U527 (N_527,In_1496,In_97);
nand U528 (N_528,In_1154,In_495);
or U529 (N_529,In_134,In_1266);
and U530 (N_530,In_1010,In_1145);
and U531 (N_531,In_882,In_33);
or U532 (N_532,In_688,In_521);
and U533 (N_533,In_488,In_1139);
and U534 (N_534,In_1040,In_627);
nor U535 (N_535,In_577,In_814);
nor U536 (N_536,In_413,In_436);
nor U537 (N_537,In_568,In_455);
nor U538 (N_538,In_656,In_660);
and U539 (N_539,In_512,In_466);
or U540 (N_540,In_927,In_289);
and U541 (N_541,In_1173,In_393);
nor U542 (N_542,In_1127,In_823);
nor U543 (N_543,In_308,In_1263);
and U544 (N_544,In_977,In_703);
nor U545 (N_545,In_270,In_246);
nand U546 (N_546,In_1295,In_622);
nor U547 (N_547,In_980,In_581);
nor U548 (N_548,In_334,In_866);
nor U549 (N_549,In_51,In_503);
and U550 (N_550,In_509,In_400);
or U551 (N_551,In_833,In_1427);
nand U552 (N_552,In_522,In_147);
nor U553 (N_553,In_1389,In_549);
nor U554 (N_554,In_34,In_573);
and U555 (N_555,In_1157,In_799);
or U556 (N_556,In_385,In_311);
nor U557 (N_557,In_1456,In_1457);
nor U558 (N_558,In_1347,In_23);
and U559 (N_559,In_259,In_150);
or U560 (N_560,In_1324,In_6);
and U561 (N_561,In_681,In_887);
nand U562 (N_562,In_837,In_36);
nand U563 (N_563,In_470,In_48);
nor U564 (N_564,In_1146,In_1129);
or U565 (N_565,In_666,In_1383);
nor U566 (N_566,In_662,In_1370);
nand U567 (N_567,In_653,In_1281);
nand U568 (N_568,In_846,In_1400);
nand U569 (N_569,In_252,In_275);
nand U570 (N_570,In_1474,In_1005);
and U571 (N_571,In_387,In_189);
and U572 (N_572,In_645,In_981);
nand U573 (N_573,In_1199,In_1385);
and U574 (N_574,In_1356,In_145);
nor U575 (N_575,In_880,In_983);
or U576 (N_576,In_520,In_1045);
and U577 (N_577,In_971,In_1077);
and U578 (N_578,In_920,In_292);
or U579 (N_579,In_53,In_783);
nor U580 (N_580,In_1268,In_476);
nand U581 (N_581,In_1415,In_317);
and U582 (N_582,In_1397,In_240);
and U583 (N_583,In_808,In_785);
or U584 (N_584,In_245,In_1017);
or U585 (N_585,In_188,In_1368);
nand U586 (N_586,In_354,In_209);
nand U587 (N_587,In_1066,In_494);
or U588 (N_588,In_1225,In_249);
and U589 (N_589,In_151,In_540);
nand U590 (N_590,In_940,In_1035);
nand U591 (N_591,In_190,In_1354);
nor U592 (N_592,In_120,In_804);
nand U593 (N_593,In_1357,In_390);
nor U594 (N_594,In_1091,In_185);
nand U595 (N_595,In_231,In_1497);
and U596 (N_596,In_1201,In_142);
nand U597 (N_597,In_641,In_1162);
and U598 (N_598,In_412,In_198);
or U599 (N_599,In_967,In_792);
or U600 (N_600,In_1413,In_473);
or U601 (N_601,In_490,In_131);
and U602 (N_602,In_1038,In_499);
and U603 (N_603,In_597,In_309);
or U604 (N_604,In_1420,In_1330);
and U605 (N_605,In_424,In_1083);
nor U606 (N_606,In_899,In_284);
or U607 (N_607,In_181,In_1155);
nor U608 (N_608,In_100,In_1103);
nor U609 (N_609,In_37,In_1023);
or U610 (N_610,In_890,In_239);
or U611 (N_611,In_1198,In_770);
and U612 (N_612,In_160,In_1128);
or U613 (N_613,In_350,In_640);
and U614 (N_614,In_94,In_571);
nor U615 (N_615,In_740,In_925);
nand U616 (N_616,In_447,In_724);
nand U617 (N_617,In_40,In_739);
or U618 (N_618,In_990,In_865);
nand U619 (N_619,In_1243,In_669);
nor U620 (N_620,In_396,In_722);
or U621 (N_621,In_515,In_459);
nand U622 (N_622,In_516,In_1197);
and U623 (N_623,In_668,In_1418);
nand U624 (N_624,In_1151,In_1183);
or U625 (N_625,In_87,In_1233);
nand U626 (N_626,In_12,In_937);
or U627 (N_627,In_1251,In_1100);
nand U628 (N_628,In_1059,In_1072);
and U629 (N_629,In_200,In_1051);
or U630 (N_630,In_1195,In_414);
and U631 (N_631,In_611,In_637);
xor U632 (N_632,In_869,In_1021);
nand U633 (N_633,In_98,In_962);
or U634 (N_634,In_11,In_1372);
nor U635 (N_635,In_254,In_1110);
nand U636 (N_636,In_556,In_1052);
nor U637 (N_637,In_247,In_253);
and U638 (N_638,In_1,In_1156);
nor U639 (N_639,In_1176,In_465);
or U640 (N_640,In_1244,In_1293);
nand U641 (N_641,In_909,In_1140);
nand U642 (N_642,In_38,In_1482);
and U643 (N_643,In_797,In_1367);
nand U644 (N_644,In_633,In_756);
nand U645 (N_645,In_1090,In_71);
nand U646 (N_646,In_1063,In_122);
nand U647 (N_647,In_143,In_795);
nand U648 (N_648,In_1202,In_163);
nor U649 (N_649,In_836,In_1309);
or U650 (N_650,In_220,In_1099);
nand U651 (N_651,In_402,In_563);
or U652 (N_652,In_541,In_118);
nor U653 (N_653,In_1150,In_859);
nand U654 (N_654,In_1141,In_1471);
and U655 (N_655,In_358,In_305);
and U656 (N_656,In_679,In_452);
or U657 (N_657,In_1054,In_61);
or U658 (N_658,In_1109,In_1481);
nor U659 (N_659,In_829,In_787);
and U660 (N_660,In_897,In_219);
xnor U661 (N_661,In_251,In_1294);
or U662 (N_662,In_1028,In_991);
and U663 (N_663,In_544,In_803);
nand U664 (N_664,In_271,In_1092);
or U665 (N_665,In_444,In_809);
nor U666 (N_666,In_238,In_480);
nand U667 (N_667,In_1409,In_365);
and U668 (N_668,In_871,In_635);
or U669 (N_669,In_296,In_1320);
nand U670 (N_670,In_667,In_265);
nand U671 (N_671,In_1433,In_507);
and U672 (N_672,In_1256,In_1446);
nand U673 (N_673,In_816,In_213);
nor U674 (N_674,In_472,In_963);
and U675 (N_675,In_449,In_164);
or U676 (N_676,In_1014,In_821);
nor U677 (N_677,In_607,In_868);
nor U678 (N_678,In_1124,In_215);
or U679 (N_679,In_1060,In_0);
or U680 (N_680,In_1019,In_555);
or U681 (N_681,In_1182,In_954);
nand U682 (N_682,In_675,In_1011);
or U683 (N_683,In_1144,In_709);
or U684 (N_684,In_1087,In_558);
nor U685 (N_685,In_643,In_1342);
nand U686 (N_686,In_831,In_1490);
nand U687 (N_687,In_467,In_362);
nand U688 (N_688,In_1104,In_1224);
nor U689 (N_689,In_157,In_1279);
and U690 (N_690,In_1381,In_561);
nand U691 (N_691,In_969,In_243);
or U692 (N_692,In_356,In_291);
and U693 (N_693,In_585,In_921);
nor U694 (N_694,In_789,In_66);
nor U695 (N_695,In_705,In_930);
or U696 (N_696,In_1310,In_1451);
or U697 (N_697,In_970,In_1460);
nor U698 (N_698,In_941,In_148);
and U699 (N_699,In_1469,In_441);
nand U700 (N_700,In_791,In_612);
and U701 (N_701,In_811,In_26);
and U702 (N_702,In_1378,In_1443);
or U703 (N_703,In_934,In_1421);
or U704 (N_704,In_749,In_707);
nor U705 (N_705,In_575,In_1178);
and U706 (N_706,In_910,In_554);
nor U707 (N_707,In_468,In_370);
or U708 (N_708,In_366,In_1472);
nand U709 (N_709,In_1264,In_952);
or U710 (N_710,In_1241,In_911);
or U711 (N_711,In_535,In_126);
and U712 (N_712,In_294,In_1428);
and U713 (N_713,In_216,In_638);
or U714 (N_714,In_832,In_1164);
and U715 (N_715,In_730,In_1353);
nand U716 (N_716,In_1123,In_242);
nor U717 (N_717,In_1219,In_1403);
nor U718 (N_718,In_896,In_31);
nand U719 (N_719,In_825,In_330);
nor U720 (N_720,In_1429,In_408);
nand U721 (N_721,In_329,In_297);
and U722 (N_722,In_938,In_173);
nor U723 (N_723,In_55,In_1246);
nor U724 (N_724,In_1454,In_786);
and U725 (N_725,In_839,In_103);
nand U726 (N_726,In_73,In_1306);
nor U727 (N_727,In_1058,In_1218);
or U728 (N_728,In_355,In_1006);
and U729 (N_729,In_1267,In_460);
nor U730 (N_730,In_1463,In_1364);
or U731 (N_731,In_1067,In_299);
or U732 (N_732,In_949,In_1250);
nor U733 (N_733,In_988,In_1333);
or U734 (N_734,In_800,In_1380);
and U735 (N_735,In_133,In_214);
nor U736 (N_736,In_782,In_922);
nor U737 (N_737,In_530,In_502);
nand U738 (N_738,In_1070,In_727);
nor U739 (N_739,In_605,In_13);
or U740 (N_740,In_361,In_603);
and U741 (N_741,In_1340,In_376);
or U742 (N_742,In_1439,In_1391);
and U743 (N_743,In_278,In_650);
nand U744 (N_744,In_425,In_421);
nor U745 (N_745,In_620,In_986);
and U746 (N_746,In_141,In_41);
nor U747 (N_747,In_1030,In_1050);
or U748 (N_748,In_481,In_807);
and U749 (N_749,In_439,In_1200);
xnor U750 (N_750,In_479,In_623);
and U751 (N_751,In_418,In_718);
or U752 (N_752,In_1458,In_135);
nor U753 (N_753,In_226,In_1455);
or U754 (N_754,In_1062,In_954);
nor U755 (N_755,In_1089,In_1051);
xnor U756 (N_756,In_410,In_347);
nor U757 (N_757,In_700,In_353);
or U758 (N_758,In_1003,In_319);
nor U759 (N_759,In_815,In_1288);
and U760 (N_760,In_72,In_1034);
and U761 (N_761,In_243,In_9);
or U762 (N_762,In_1234,In_1232);
or U763 (N_763,In_910,In_17);
and U764 (N_764,In_1346,In_129);
or U765 (N_765,In_1166,In_701);
nor U766 (N_766,In_158,In_1400);
nand U767 (N_767,In_469,In_923);
nand U768 (N_768,In_1057,In_80);
and U769 (N_769,In_994,In_1493);
and U770 (N_770,In_309,In_604);
or U771 (N_771,In_563,In_962);
nor U772 (N_772,In_418,In_646);
nand U773 (N_773,In_1248,In_1223);
or U774 (N_774,In_752,In_539);
nor U775 (N_775,In_1246,In_1273);
and U776 (N_776,In_393,In_1392);
nor U777 (N_777,In_624,In_161);
and U778 (N_778,In_734,In_1191);
nor U779 (N_779,In_135,In_1241);
or U780 (N_780,In_568,In_359);
and U781 (N_781,In_1093,In_1367);
or U782 (N_782,In_143,In_861);
and U783 (N_783,In_194,In_941);
and U784 (N_784,In_1207,In_890);
or U785 (N_785,In_646,In_812);
nand U786 (N_786,In_285,In_240);
or U787 (N_787,In_139,In_840);
nand U788 (N_788,In_869,In_1460);
nand U789 (N_789,In_742,In_1403);
nor U790 (N_790,In_1355,In_43);
nor U791 (N_791,In_1339,In_490);
nor U792 (N_792,In_555,In_545);
or U793 (N_793,In_1211,In_704);
nand U794 (N_794,In_379,In_967);
nand U795 (N_795,In_1370,In_27);
or U796 (N_796,In_950,In_733);
nand U797 (N_797,In_1204,In_1299);
nor U798 (N_798,In_528,In_424);
or U799 (N_799,In_1302,In_1111);
and U800 (N_800,In_1307,In_1475);
nand U801 (N_801,In_82,In_319);
nor U802 (N_802,In_473,In_520);
and U803 (N_803,In_1236,In_1195);
or U804 (N_804,In_775,In_842);
nor U805 (N_805,In_750,In_932);
nor U806 (N_806,In_874,In_362);
nand U807 (N_807,In_110,In_901);
nor U808 (N_808,In_451,In_1409);
nor U809 (N_809,In_830,In_552);
nand U810 (N_810,In_1149,In_523);
nor U811 (N_811,In_821,In_339);
nor U812 (N_812,In_34,In_1090);
nor U813 (N_813,In_957,In_1467);
or U814 (N_814,In_657,In_408);
nand U815 (N_815,In_759,In_110);
or U816 (N_816,In_1165,In_906);
nor U817 (N_817,In_142,In_911);
nand U818 (N_818,In_514,In_40);
or U819 (N_819,In_1089,In_880);
nand U820 (N_820,In_738,In_654);
nand U821 (N_821,In_218,In_1142);
or U822 (N_822,In_1199,In_931);
nand U823 (N_823,In_1376,In_835);
or U824 (N_824,In_1080,In_579);
and U825 (N_825,In_789,In_1428);
nand U826 (N_826,In_1061,In_232);
nand U827 (N_827,In_23,In_1273);
nand U828 (N_828,In_1298,In_925);
or U829 (N_829,In_671,In_745);
nor U830 (N_830,In_1234,In_399);
nor U831 (N_831,In_922,In_933);
nor U832 (N_832,In_618,In_1466);
or U833 (N_833,In_771,In_1304);
nand U834 (N_834,In_314,In_659);
and U835 (N_835,In_1257,In_1166);
and U836 (N_836,In_1163,In_512);
or U837 (N_837,In_84,In_570);
nor U838 (N_838,In_561,In_1326);
and U839 (N_839,In_1098,In_41);
and U840 (N_840,In_989,In_720);
nand U841 (N_841,In_1308,In_21);
nor U842 (N_842,In_218,In_283);
nor U843 (N_843,In_75,In_945);
nor U844 (N_844,In_991,In_189);
or U845 (N_845,In_681,In_1106);
nor U846 (N_846,In_228,In_1154);
nand U847 (N_847,In_169,In_51);
or U848 (N_848,In_832,In_289);
and U849 (N_849,In_204,In_1160);
or U850 (N_850,In_1369,In_1050);
nor U851 (N_851,In_834,In_1229);
nand U852 (N_852,In_335,In_741);
nor U853 (N_853,In_1180,In_896);
and U854 (N_854,In_1475,In_740);
nand U855 (N_855,In_1418,In_1476);
or U856 (N_856,In_370,In_710);
nor U857 (N_857,In_1099,In_111);
or U858 (N_858,In_667,In_1397);
nor U859 (N_859,In_1456,In_1291);
or U860 (N_860,In_1173,In_666);
nor U861 (N_861,In_853,In_723);
or U862 (N_862,In_503,In_578);
nor U863 (N_863,In_747,In_86);
and U864 (N_864,In_994,In_66);
xor U865 (N_865,In_617,In_1486);
nand U866 (N_866,In_1117,In_861);
nand U867 (N_867,In_932,In_981);
or U868 (N_868,In_340,In_84);
nor U869 (N_869,In_1013,In_106);
or U870 (N_870,In_303,In_406);
nand U871 (N_871,In_552,In_1003);
nor U872 (N_872,In_1066,In_1257);
nand U873 (N_873,In_957,In_1080);
nand U874 (N_874,In_1201,In_1075);
and U875 (N_875,In_922,In_1034);
nand U876 (N_876,In_1256,In_1092);
nand U877 (N_877,In_594,In_359);
nand U878 (N_878,In_1031,In_372);
or U879 (N_879,In_1390,In_86);
or U880 (N_880,In_883,In_131);
nor U881 (N_881,In_200,In_60);
or U882 (N_882,In_610,In_262);
nand U883 (N_883,In_960,In_1489);
nand U884 (N_884,In_690,In_450);
nand U885 (N_885,In_1186,In_0);
nand U886 (N_886,In_1445,In_927);
nand U887 (N_887,In_463,In_313);
and U888 (N_888,In_899,In_1334);
nor U889 (N_889,In_456,In_307);
and U890 (N_890,In_250,In_687);
nor U891 (N_891,In_668,In_1189);
or U892 (N_892,In_1411,In_88);
nor U893 (N_893,In_1211,In_627);
nor U894 (N_894,In_1132,In_1229);
nand U895 (N_895,In_995,In_65);
or U896 (N_896,In_1250,In_357);
nand U897 (N_897,In_152,In_986);
or U898 (N_898,In_231,In_837);
nand U899 (N_899,In_90,In_1248);
xor U900 (N_900,In_719,In_881);
or U901 (N_901,In_1175,In_354);
nand U902 (N_902,In_594,In_36);
nand U903 (N_903,In_411,In_99);
or U904 (N_904,In_1259,In_125);
or U905 (N_905,In_1232,In_36);
nand U906 (N_906,In_454,In_1367);
and U907 (N_907,In_133,In_749);
nor U908 (N_908,In_314,In_160);
nand U909 (N_909,In_586,In_59);
and U910 (N_910,In_1097,In_412);
or U911 (N_911,In_1172,In_568);
or U912 (N_912,In_329,In_1386);
or U913 (N_913,In_526,In_1152);
and U914 (N_914,In_1312,In_540);
nor U915 (N_915,In_1243,In_94);
and U916 (N_916,In_972,In_29);
or U917 (N_917,In_1127,In_1232);
or U918 (N_918,In_886,In_415);
and U919 (N_919,In_1378,In_966);
or U920 (N_920,In_1400,In_715);
or U921 (N_921,In_321,In_1022);
and U922 (N_922,In_537,In_1296);
nor U923 (N_923,In_1206,In_351);
and U924 (N_924,In_480,In_846);
or U925 (N_925,In_134,In_1319);
nor U926 (N_926,In_435,In_1432);
nor U927 (N_927,In_349,In_708);
nand U928 (N_928,In_162,In_279);
or U929 (N_929,In_580,In_964);
and U930 (N_930,In_1347,In_1178);
or U931 (N_931,In_925,In_945);
or U932 (N_932,In_904,In_534);
nor U933 (N_933,In_64,In_315);
nor U934 (N_934,In_1478,In_1056);
nor U935 (N_935,In_1439,In_502);
or U936 (N_936,In_889,In_721);
and U937 (N_937,In_273,In_1477);
and U938 (N_938,In_1464,In_847);
or U939 (N_939,In_146,In_75);
and U940 (N_940,In_1286,In_181);
nor U941 (N_941,In_1496,In_454);
or U942 (N_942,In_266,In_989);
nor U943 (N_943,In_862,In_849);
and U944 (N_944,In_836,In_1186);
and U945 (N_945,In_291,In_414);
or U946 (N_946,In_862,In_25);
or U947 (N_947,In_490,In_79);
and U948 (N_948,In_424,In_1392);
or U949 (N_949,In_858,In_1029);
or U950 (N_950,In_409,In_67);
nand U951 (N_951,In_1337,In_15);
nand U952 (N_952,In_1247,In_1222);
nand U953 (N_953,In_236,In_1124);
or U954 (N_954,In_54,In_647);
and U955 (N_955,In_1020,In_541);
or U956 (N_956,In_1000,In_1471);
nor U957 (N_957,In_738,In_547);
nand U958 (N_958,In_401,In_319);
and U959 (N_959,In_313,In_76);
nand U960 (N_960,In_1193,In_848);
and U961 (N_961,In_408,In_1011);
nand U962 (N_962,In_1224,In_826);
nor U963 (N_963,In_1272,In_263);
nor U964 (N_964,In_396,In_91);
and U965 (N_965,In_512,In_365);
nor U966 (N_966,In_764,In_1253);
or U967 (N_967,In_1253,In_1030);
or U968 (N_968,In_979,In_220);
and U969 (N_969,In_589,In_817);
xor U970 (N_970,In_876,In_1218);
or U971 (N_971,In_487,In_263);
and U972 (N_972,In_709,In_74);
and U973 (N_973,In_553,In_891);
or U974 (N_974,In_859,In_478);
nand U975 (N_975,In_417,In_660);
nand U976 (N_976,In_304,In_470);
or U977 (N_977,In_537,In_1435);
or U978 (N_978,In_802,In_1377);
or U979 (N_979,In_65,In_1028);
nor U980 (N_980,In_1424,In_647);
nor U981 (N_981,In_367,In_129);
xnor U982 (N_982,In_1014,In_1136);
nor U983 (N_983,In_1077,In_995);
and U984 (N_984,In_439,In_221);
or U985 (N_985,In_922,In_172);
nor U986 (N_986,In_299,In_792);
and U987 (N_987,In_276,In_1038);
and U988 (N_988,In_1215,In_927);
nor U989 (N_989,In_1115,In_809);
nand U990 (N_990,In_852,In_383);
nor U991 (N_991,In_1446,In_987);
nand U992 (N_992,In_896,In_738);
or U993 (N_993,In_1429,In_1315);
nor U994 (N_994,In_63,In_388);
nand U995 (N_995,In_35,In_875);
and U996 (N_996,In_631,In_136);
nor U997 (N_997,In_1365,In_362);
nor U998 (N_998,In_72,In_1255);
nor U999 (N_999,In_29,In_218);
nand U1000 (N_1000,In_1213,In_175);
and U1001 (N_1001,In_1079,In_919);
nand U1002 (N_1002,In_597,In_64);
nor U1003 (N_1003,In_569,In_1209);
nor U1004 (N_1004,In_462,In_848);
or U1005 (N_1005,In_464,In_89);
and U1006 (N_1006,In_704,In_297);
or U1007 (N_1007,In_751,In_293);
nand U1008 (N_1008,In_29,In_755);
or U1009 (N_1009,In_433,In_814);
or U1010 (N_1010,In_670,In_969);
and U1011 (N_1011,In_167,In_924);
and U1012 (N_1012,In_504,In_410);
nor U1013 (N_1013,In_1384,In_377);
nor U1014 (N_1014,In_175,In_878);
or U1015 (N_1015,In_327,In_942);
or U1016 (N_1016,In_616,In_873);
and U1017 (N_1017,In_840,In_825);
and U1018 (N_1018,In_267,In_1343);
nand U1019 (N_1019,In_84,In_842);
nand U1020 (N_1020,In_31,In_477);
and U1021 (N_1021,In_1049,In_1342);
or U1022 (N_1022,In_622,In_460);
nor U1023 (N_1023,In_123,In_229);
nor U1024 (N_1024,In_1483,In_1400);
xnor U1025 (N_1025,In_1372,In_1154);
nand U1026 (N_1026,In_1173,In_449);
nand U1027 (N_1027,In_1203,In_230);
and U1028 (N_1028,In_204,In_915);
or U1029 (N_1029,In_225,In_494);
nor U1030 (N_1030,In_1143,In_1182);
or U1031 (N_1031,In_838,In_1296);
and U1032 (N_1032,In_156,In_482);
or U1033 (N_1033,In_1315,In_1100);
nand U1034 (N_1034,In_1179,In_735);
nor U1035 (N_1035,In_995,In_754);
and U1036 (N_1036,In_1368,In_936);
or U1037 (N_1037,In_386,In_520);
and U1038 (N_1038,In_666,In_931);
and U1039 (N_1039,In_892,In_1432);
and U1040 (N_1040,In_1416,In_931);
nor U1041 (N_1041,In_980,In_489);
or U1042 (N_1042,In_1417,In_385);
or U1043 (N_1043,In_1368,In_952);
nand U1044 (N_1044,In_1234,In_671);
and U1045 (N_1045,In_1017,In_737);
nor U1046 (N_1046,In_1155,In_1157);
or U1047 (N_1047,In_832,In_628);
or U1048 (N_1048,In_347,In_400);
and U1049 (N_1049,In_310,In_108);
and U1050 (N_1050,In_148,In_740);
nor U1051 (N_1051,In_65,In_1172);
and U1052 (N_1052,In_73,In_1190);
or U1053 (N_1053,In_225,In_1077);
nand U1054 (N_1054,In_1171,In_1179);
and U1055 (N_1055,In_1457,In_1367);
nor U1056 (N_1056,In_152,In_93);
or U1057 (N_1057,In_1472,In_1461);
nor U1058 (N_1058,In_474,In_1326);
nor U1059 (N_1059,In_875,In_124);
or U1060 (N_1060,In_274,In_405);
or U1061 (N_1061,In_996,In_318);
nor U1062 (N_1062,In_752,In_1272);
nand U1063 (N_1063,In_1439,In_636);
and U1064 (N_1064,In_1331,In_588);
nand U1065 (N_1065,In_211,In_1291);
nand U1066 (N_1066,In_515,In_1429);
or U1067 (N_1067,In_79,In_661);
and U1068 (N_1068,In_1428,In_1138);
or U1069 (N_1069,In_651,In_807);
nand U1070 (N_1070,In_209,In_1353);
nor U1071 (N_1071,In_986,In_1290);
nor U1072 (N_1072,In_1462,In_739);
nor U1073 (N_1073,In_763,In_1492);
nor U1074 (N_1074,In_724,In_1108);
nor U1075 (N_1075,In_1397,In_388);
or U1076 (N_1076,In_137,In_1389);
or U1077 (N_1077,In_1013,In_992);
or U1078 (N_1078,In_229,In_1253);
nor U1079 (N_1079,In_303,In_644);
and U1080 (N_1080,In_770,In_294);
nor U1081 (N_1081,In_786,In_1194);
nor U1082 (N_1082,In_604,In_730);
xor U1083 (N_1083,In_709,In_495);
and U1084 (N_1084,In_143,In_515);
and U1085 (N_1085,In_434,In_794);
or U1086 (N_1086,In_469,In_42);
or U1087 (N_1087,In_1050,In_555);
and U1088 (N_1088,In_247,In_1285);
or U1089 (N_1089,In_290,In_1182);
and U1090 (N_1090,In_849,In_765);
nor U1091 (N_1091,In_266,In_1005);
nor U1092 (N_1092,In_540,In_990);
or U1093 (N_1093,In_240,In_55);
nor U1094 (N_1094,In_650,In_205);
and U1095 (N_1095,In_780,In_523);
or U1096 (N_1096,In_1100,In_1114);
or U1097 (N_1097,In_711,In_276);
or U1098 (N_1098,In_1290,In_563);
or U1099 (N_1099,In_1126,In_1275);
nor U1100 (N_1100,In_609,In_1029);
and U1101 (N_1101,In_1324,In_1335);
nor U1102 (N_1102,In_72,In_442);
nor U1103 (N_1103,In_437,In_1101);
nand U1104 (N_1104,In_297,In_950);
nor U1105 (N_1105,In_1253,In_846);
xnor U1106 (N_1106,In_453,In_708);
nor U1107 (N_1107,In_711,In_1150);
and U1108 (N_1108,In_671,In_188);
or U1109 (N_1109,In_1080,In_439);
or U1110 (N_1110,In_354,In_198);
and U1111 (N_1111,In_665,In_1233);
nand U1112 (N_1112,In_665,In_1045);
or U1113 (N_1113,In_217,In_287);
nand U1114 (N_1114,In_1276,In_1040);
nand U1115 (N_1115,In_1012,In_854);
nand U1116 (N_1116,In_72,In_1413);
nor U1117 (N_1117,In_582,In_1038);
nand U1118 (N_1118,In_989,In_1342);
nand U1119 (N_1119,In_386,In_356);
and U1120 (N_1120,In_545,In_560);
nor U1121 (N_1121,In_301,In_528);
nand U1122 (N_1122,In_1206,In_116);
and U1123 (N_1123,In_496,In_369);
or U1124 (N_1124,In_270,In_1210);
and U1125 (N_1125,In_870,In_177);
nand U1126 (N_1126,In_1345,In_1326);
nand U1127 (N_1127,In_1171,In_1105);
or U1128 (N_1128,In_869,In_46);
nor U1129 (N_1129,In_567,In_747);
or U1130 (N_1130,In_383,In_615);
and U1131 (N_1131,In_367,In_1021);
nand U1132 (N_1132,In_108,In_865);
xor U1133 (N_1133,In_600,In_936);
nand U1134 (N_1134,In_622,In_230);
and U1135 (N_1135,In_527,In_1007);
or U1136 (N_1136,In_24,In_1441);
or U1137 (N_1137,In_549,In_795);
and U1138 (N_1138,In_916,In_357);
or U1139 (N_1139,In_122,In_20);
or U1140 (N_1140,In_1036,In_1100);
or U1141 (N_1141,In_1393,In_1444);
or U1142 (N_1142,In_1192,In_658);
and U1143 (N_1143,In_166,In_238);
nor U1144 (N_1144,In_900,In_166);
or U1145 (N_1145,In_1085,In_1233);
nor U1146 (N_1146,In_514,In_308);
nor U1147 (N_1147,In_1330,In_735);
nand U1148 (N_1148,In_1289,In_1310);
and U1149 (N_1149,In_1470,In_1410);
and U1150 (N_1150,In_118,In_348);
or U1151 (N_1151,In_3,In_126);
nand U1152 (N_1152,In_1361,In_315);
and U1153 (N_1153,In_1040,In_379);
nand U1154 (N_1154,In_723,In_347);
and U1155 (N_1155,In_1283,In_71);
and U1156 (N_1156,In_1186,In_351);
and U1157 (N_1157,In_1022,In_495);
or U1158 (N_1158,In_959,In_1182);
or U1159 (N_1159,In_1429,In_1017);
xor U1160 (N_1160,In_987,In_244);
and U1161 (N_1161,In_225,In_128);
or U1162 (N_1162,In_1029,In_383);
nand U1163 (N_1163,In_156,In_995);
and U1164 (N_1164,In_1409,In_890);
and U1165 (N_1165,In_285,In_268);
nor U1166 (N_1166,In_131,In_140);
nand U1167 (N_1167,In_1411,In_12);
nand U1168 (N_1168,In_975,In_298);
or U1169 (N_1169,In_129,In_391);
nor U1170 (N_1170,In_38,In_761);
nand U1171 (N_1171,In_274,In_1466);
nor U1172 (N_1172,In_189,In_610);
or U1173 (N_1173,In_1111,In_1181);
nor U1174 (N_1174,In_206,In_113);
or U1175 (N_1175,In_261,In_1093);
nand U1176 (N_1176,In_484,In_164);
nand U1177 (N_1177,In_23,In_310);
nor U1178 (N_1178,In_1027,In_1468);
or U1179 (N_1179,In_1155,In_1400);
nor U1180 (N_1180,In_1144,In_1247);
and U1181 (N_1181,In_828,In_1107);
nor U1182 (N_1182,In_1084,In_392);
nor U1183 (N_1183,In_616,In_1057);
nand U1184 (N_1184,In_325,In_1249);
or U1185 (N_1185,In_25,In_1110);
or U1186 (N_1186,In_1000,In_766);
nand U1187 (N_1187,In_421,In_57);
nor U1188 (N_1188,In_1365,In_381);
and U1189 (N_1189,In_512,In_127);
nand U1190 (N_1190,In_645,In_26);
nand U1191 (N_1191,In_184,In_160);
nor U1192 (N_1192,In_149,In_1274);
or U1193 (N_1193,In_555,In_94);
nor U1194 (N_1194,In_958,In_143);
nand U1195 (N_1195,In_365,In_1229);
and U1196 (N_1196,In_1209,In_527);
or U1197 (N_1197,In_1321,In_275);
nand U1198 (N_1198,In_1140,In_1036);
or U1199 (N_1199,In_1131,In_537);
and U1200 (N_1200,In_858,In_335);
and U1201 (N_1201,In_1300,In_1211);
or U1202 (N_1202,In_839,In_1097);
or U1203 (N_1203,In_860,In_1184);
or U1204 (N_1204,In_236,In_706);
nor U1205 (N_1205,In_843,In_61);
nor U1206 (N_1206,In_1080,In_1071);
or U1207 (N_1207,In_948,In_662);
nor U1208 (N_1208,In_77,In_1396);
nand U1209 (N_1209,In_304,In_709);
nor U1210 (N_1210,In_389,In_268);
nor U1211 (N_1211,In_853,In_964);
nand U1212 (N_1212,In_77,In_284);
nand U1213 (N_1213,In_960,In_895);
nor U1214 (N_1214,In_318,In_380);
and U1215 (N_1215,In_1148,In_1099);
nand U1216 (N_1216,In_339,In_791);
nand U1217 (N_1217,In_803,In_117);
nor U1218 (N_1218,In_57,In_1199);
or U1219 (N_1219,In_286,In_204);
nand U1220 (N_1220,In_922,In_1230);
nand U1221 (N_1221,In_952,In_1017);
nor U1222 (N_1222,In_1330,In_928);
nand U1223 (N_1223,In_180,In_1263);
and U1224 (N_1224,In_591,In_940);
nor U1225 (N_1225,In_1037,In_270);
nor U1226 (N_1226,In_137,In_1002);
or U1227 (N_1227,In_581,In_919);
and U1228 (N_1228,In_420,In_396);
or U1229 (N_1229,In_1120,In_456);
or U1230 (N_1230,In_388,In_440);
or U1231 (N_1231,In_328,In_873);
or U1232 (N_1232,In_160,In_1131);
nor U1233 (N_1233,In_1078,In_557);
nand U1234 (N_1234,In_737,In_447);
nand U1235 (N_1235,In_1301,In_769);
nor U1236 (N_1236,In_172,In_777);
or U1237 (N_1237,In_277,In_847);
nand U1238 (N_1238,In_701,In_1475);
and U1239 (N_1239,In_694,In_1161);
or U1240 (N_1240,In_372,In_119);
nand U1241 (N_1241,In_422,In_923);
nand U1242 (N_1242,In_1069,In_692);
nor U1243 (N_1243,In_179,In_98);
nor U1244 (N_1244,In_1429,In_470);
or U1245 (N_1245,In_31,In_1244);
and U1246 (N_1246,In_163,In_1476);
nand U1247 (N_1247,In_1232,In_303);
and U1248 (N_1248,In_1060,In_109);
nor U1249 (N_1249,In_771,In_326);
and U1250 (N_1250,In_38,In_625);
xnor U1251 (N_1251,In_153,In_104);
nor U1252 (N_1252,In_1238,In_1042);
and U1253 (N_1253,In_1349,In_1082);
nand U1254 (N_1254,In_1455,In_1122);
and U1255 (N_1255,In_1045,In_710);
and U1256 (N_1256,In_1119,In_1135);
and U1257 (N_1257,In_1282,In_1467);
and U1258 (N_1258,In_1463,In_1009);
and U1259 (N_1259,In_558,In_793);
nor U1260 (N_1260,In_1213,In_1263);
nand U1261 (N_1261,In_457,In_864);
or U1262 (N_1262,In_278,In_1144);
nand U1263 (N_1263,In_365,In_448);
nor U1264 (N_1264,In_587,In_1179);
and U1265 (N_1265,In_505,In_1274);
nor U1266 (N_1266,In_92,In_1307);
and U1267 (N_1267,In_846,In_1345);
and U1268 (N_1268,In_519,In_1462);
and U1269 (N_1269,In_430,In_746);
nand U1270 (N_1270,In_492,In_976);
and U1271 (N_1271,In_1085,In_1170);
or U1272 (N_1272,In_989,In_1264);
and U1273 (N_1273,In_565,In_710);
and U1274 (N_1274,In_128,In_31);
nor U1275 (N_1275,In_1313,In_603);
and U1276 (N_1276,In_176,In_268);
or U1277 (N_1277,In_799,In_426);
nor U1278 (N_1278,In_988,In_372);
or U1279 (N_1279,In_1344,In_663);
and U1280 (N_1280,In_549,In_965);
or U1281 (N_1281,In_385,In_269);
or U1282 (N_1282,In_452,In_1056);
nor U1283 (N_1283,In_475,In_71);
or U1284 (N_1284,In_647,In_499);
or U1285 (N_1285,In_124,In_1100);
nand U1286 (N_1286,In_61,In_948);
nor U1287 (N_1287,In_466,In_1151);
and U1288 (N_1288,In_847,In_1324);
nand U1289 (N_1289,In_270,In_549);
nand U1290 (N_1290,In_945,In_589);
and U1291 (N_1291,In_1346,In_594);
nor U1292 (N_1292,In_433,In_828);
and U1293 (N_1293,In_806,In_353);
and U1294 (N_1294,In_584,In_1168);
nor U1295 (N_1295,In_1271,In_289);
nand U1296 (N_1296,In_468,In_934);
nand U1297 (N_1297,In_1399,In_329);
and U1298 (N_1298,In_1260,In_1271);
and U1299 (N_1299,In_161,In_1);
or U1300 (N_1300,In_107,In_530);
nor U1301 (N_1301,In_1460,In_547);
nand U1302 (N_1302,In_678,In_417);
and U1303 (N_1303,In_101,In_970);
or U1304 (N_1304,In_1096,In_301);
or U1305 (N_1305,In_1293,In_788);
nor U1306 (N_1306,In_442,In_248);
nor U1307 (N_1307,In_77,In_1463);
nor U1308 (N_1308,In_232,In_979);
and U1309 (N_1309,In_1315,In_53);
nor U1310 (N_1310,In_177,In_1016);
and U1311 (N_1311,In_825,In_1404);
nand U1312 (N_1312,In_296,In_964);
and U1313 (N_1313,In_72,In_1130);
or U1314 (N_1314,In_862,In_1409);
or U1315 (N_1315,In_1018,In_805);
nand U1316 (N_1316,In_682,In_34);
or U1317 (N_1317,In_1175,In_1354);
or U1318 (N_1318,In_1484,In_53);
nand U1319 (N_1319,In_817,In_1369);
nand U1320 (N_1320,In_24,In_330);
nor U1321 (N_1321,In_1060,In_349);
nand U1322 (N_1322,In_271,In_1341);
nand U1323 (N_1323,In_709,In_368);
or U1324 (N_1324,In_719,In_1229);
and U1325 (N_1325,In_1067,In_914);
nand U1326 (N_1326,In_103,In_342);
xnor U1327 (N_1327,In_1140,In_76);
and U1328 (N_1328,In_316,In_1116);
and U1329 (N_1329,In_760,In_31);
nand U1330 (N_1330,In_794,In_1218);
nand U1331 (N_1331,In_738,In_1317);
or U1332 (N_1332,In_167,In_867);
nor U1333 (N_1333,In_585,In_1362);
and U1334 (N_1334,In_382,In_1206);
nor U1335 (N_1335,In_1285,In_520);
nand U1336 (N_1336,In_654,In_1143);
nand U1337 (N_1337,In_357,In_543);
nand U1338 (N_1338,In_1068,In_514);
nand U1339 (N_1339,In_749,In_96);
nand U1340 (N_1340,In_1188,In_837);
or U1341 (N_1341,In_893,In_835);
nor U1342 (N_1342,In_1181,In_423);
nor U1343 (N_1343,In_175,In_1204);
and U1344 (N_1344,In_225,In_903);
nor U1345 (N_1345,In_1285,In_1310);
or U1346 (N_1346,In_20,In_1094);
nand U1347 (N_1347,In_325,In_789);
nand U1348 (N_1348,In_854,In_853);
or U1349 (N_1349,In_283,In_885);
nor U1350 (N_1350,In_368,In_699);
and U1351 (N_1351,In_1121,In_36);
or U1352 (N_1352,In_1204,In_765);
nor U1353 (N_1353,In_436,In_1453);
nand U1354 (N_1354,In_397,In_782);
nor U1355 (N_1355,In_881,In_189);
nand U1356 (N_1356,In_318,In_243);
nor U1357 (N_1357,In_624,In_1154);
or U1358 (N_1358,In_183,In_421);
or U1359 (N_1359,In_1037,In_1369);
and U1360 (N_1360,In_115,In_692);
nor U1361 (N_1361,In_894,In_248);
nand U1362 (N_1362,In_1397,In_943);
nand U1363 (N_1363,In_305,In_801);
and U1364 (N_1364,In_1298,In_1295);
or U1365 (N_1365,In_1114,In_962);
or U1366 (N_1366,In_165,In_183);
nand U1367 (N_1367,In_546,In_1165);
and U1368 (N_1368,In_927,In_310);
or U1369 (N_1369,In_600,In_1171);
or U1370 (N_1370,In_1221,In_1411);
nand U1371 (N_1371,In_1000,In_249);
nand U1372 (N_1372,In_597,In_1394);
nand U1373 (N_1373,In_676,In_854);
or U1374 (N_1374,In_1318,In_874);
xnor U1375 (N_1375,In_972,In_967);
and U1376 (N_1376,In_1104,In_850);
or U1377 (N_1377,In_954,In_875);
or U1378 (N_1378,In_166,In_967);
or U1379 (N_1379,In_784,In_1411);
nor U1380 (N_1380,In_5,In_1114);
xnor U1381 (N_1381,In_796,In_1174);
nor U1382 (N_1382,In_1305,In_619);
or U1383 (N_1383,In_746,In_894);
nand U1384 (N_1384,In_1205,In_669);
or U1385 (N_1385,In_738,In_391);
nor U1386 (N_1386,In_522,In_766);
or U1387 (N_1387,In_821,In_39);
nor U1388 (N_1388,In_691,In_938);
nand U1389 (N_1389,In_975,In_85);
nor U1390 (N_1390,In_799,In_588);
or U1391 (N_1391,In_1498,In_289);
and U1392 (N_1392,In_618,In_1221);
nand U1393 (N_1393,In_1180,In_1020);
or U1394 (N_1394,In_1361,In_627);
or U1395 (N_1395,In_582,In_1300);
and U1396 (N_1396,In_1003,In_754);
and U1397 (N_1397,In_303,In_683);
nand U1398 (N_1398,In_797,In_1090);
nor U1399 (N_1399,In_460,In_546);
nand U1400 (N_1400,In_305,In_698);
and U1401 (N_1401,In_845,In_562);
or U1402 (N_1402,In_800,In_1136);
and U1403 (N_1403,In_864,In_253);
and U1404 (N_1404,In_823,In_996);
or U1405 (N_1405,In_486,In_817);
nor U1406 (N_1406,In_244,In_682);
nor U1407 (N_1407,In_708,In_1255);
nand U1408 (N_1408,In_336,In_1044);
nand U1409 (N_1409,In_613,In_35);
nor U1410 (N_1410,In_379,In_10);
nand U1411 (N_1411,In_975,In_1367);
and U1412 (N_1412,In_1026,In_383);
or U1413 (N_1413,In_349,In_503);
nand U1414 (N_1414,In_775,In_1324);
nand U1415 (N_1415,In_85,In_905);
and U1416 (N_1416,In_1084,In_415);
nand U1417 (N_1417,In_1063,In_64);
nand U1418 (N_1418,In_676,In_123);
nand U1419 (N_1419,In_1251,In_1288);
or U1420 (N_1420,In_1009,In_905);
or U1421 (N_1421,In_906,In_987);
or U1422 (N_1422,In_381,In_968);
or U1423 (N_1423,In_1034,In_376);
nand U1424 (N_1424,In_358,In_617);
and U1425 (N_1425,In_536,In_494);
nor U1426 (N_1426,In_264,In_1202);
or U1427 (N_1427,In_373,In_557);
or U1428 (N_1428,In_1105,In_683);
and U1429 (N_1429,In_916,In_673);
nor U1430 (N_1430,In_1132,In_951);
nand U1431 (N_1431,In_1024,In_1300);
or U1432 (N_1432,In_1088,In_1452);
and U1433 (N_1433,In_1335,In_1227);
nor U1434 (N_1434,In_847,In_333);
or U1435 (N_1435,In_396,In_428);
nand U1436 (N_1436,In_728,In_711);
nand U1437 (N_1437,In_670,In_213);
and U1438 (N_1438,In_222,In_968);
and U1439 (N_1439,In_1010,In_666);
nand U1440 (N_1440,In_664,In_1361);
nand U1441 (N_1441,In_470,In_1460);
nor U1442 (N_1442,In_1080,In_787);
nand U1443 (N_1443,In_1438,In_324);
or U1444 (N_1444,In_534,In_1377);
or U1445 (N_1445,In_1261,In_20);
or U1446 (N_1446,In_819,In_101);
or U1447 (N_1447,In_317,In_1236);
nor U1448 (N_1448,In_903,In_524);
nand U1449 (N_1449,In_866,In_790);
or U1450 (N_1450,In_901,In_133);
or U1451 (N_1451,In_111,In_256);
nand U1452 (N_1452,In_841,In_1373);
and U1453 (N_1453,In_1322,In_880);
and U1454 (N_1454,In_120,In_707);
nand U1455 (N_1455,In_1068,In_1225);
and U1456 (N_1456,In_1260,In_964);
nand U1457 (N_1457,In_974,In_1204);
nand U1458 (N_1458,In_530,In_316);
nor U1459 (N_1459,In_1457,In_1381);
nand U1460 (N_1460,In_632,In_43);
or U1461 (N_1461,In_1126,In_49);
or U1462 (N_1462,In_957,In_172);
nand U1463 (N_1463,In_660,In_201);
or U1464 (N_1464,In_1217,In_105);
and U1465 (N_1465,In_440,In_1364);
nand U1466 (N_1466,In_53,In_250);
and U1467 (N_1467,In_916,In_934);
nand U1468 (N_1468,In_1166,In_64);
and U1469 (N_1469,In_1114,In_1000);
nor U1470 (N_1470,In_526,In_1181);
or U1471 (N_1471,In_101,In_402);
nor U1472 (N_1472,In_1216,In_1452);
and U1473 (N_1473,In_683,In_1441);
nand U1474 (N_1474,In_373,In_192);
or U1475 (N_1475,In_1484,In_737);
and U1476 (N_1476,In_1368,In_917);
nor U1477 (N_1477,In_1478,In_1215);
nor U1478 (N_1478,In_1475,In_397);
or U1479 (N_1479,In_475,In_263);
or U1480 (N_1480,In_911,In_1055);
or U1481 (N_1481,In_485,In_1146);
nor U1482 (N_1482,In_323,In_164);
or U1483 (N_1483,In_775,In_1164);
nand U1484 (N_1484,In_1050,In_424);
nor U1485 (N_1485,In_1049,In_342);
nand U1486 (N_1486,In_285,In_776);
and U1487 (N_1487,In_135,In_345);
or U1488 (N_1488,In_1487,In_1141);
and U1489 (N_1489,In_556,In_318);
nand U1490 (N_1490,In_474,In_224);
and U1491 (N_1491,In_1493,In_1105);
nor U1492 (N_1492,In_623,In_1063);
nor U1493 (N_1493,In_129,In_1225);
nand U1494 (N_1494,In_1058,In_1195);
nand U1495 (N_1495,In_163,In_1436);
and U1496 (N_1496,In_268,In_910);
nand U1497 (N_1497,In_112,In_1259);
or U1498 (N_1498,In_1048,In_775);
or U1499 (N_1499,In_1034,In_652);
and U1500 (N_1500,In_194,In_956);
or U1501 (N_1501,In_58,In_259);
or U1502 (N_1502,In_1099,In_1145);
nor U1503 (N_1503,In_1001,In_422);
and U1504 (N_1504,In_1444,In_1104);
or U1505 (N_1505,In_169,In_1147);
and U1506 (N_1506,In_413,In_885);
nand U1507 (N_1507,In_88,In_343);
or U1508 (N_1508,In_696,In_1392);
nor U1509 (N_1509,In_546,In_1275);
nor U1510 (N_1510,In_1151,In_1412);
or U1511 (N_1511,In_877,In_337);
nand U1512 (N_1512,In_281,In_1478);
or U1513 (N_1513,In_50,In_520);
or U1514 (N_1514,In_428,In_1456);
nand U1515 (N_1515,In_753,In_1325);
and U1516 (N_1516,In_905,In_1072);
and U1517 (N_1517,In_1312,In_84);
xor U1518 (N_1518,In_120,In_993);
nor U1519 (N_1519,In_1376,In_1493);
nand U1520 (N_1520,In_572,In_163);
or U1521 (N_1521,In_572,In_214);
or U1522 (N_1522,In_334,In_710);
nor U1523 (N_1523,In_70,In_1091);
nor U1524 (N_1524,In_333,In_1312);
and U1525 (N_1525,In_1398,In_615);
nor U1526 (N_1526,In_954,In_1016);
and U1527 (N_1527,In_341,In_645);
nor U1528 (N_1528,In_525,In_607);
nor U1529 (N_1529,In_302,In_1449);
nand U1530 (N_1530,In_392,In_1083);
nand U1531 (N_1531,In_351,In_1120);
nor U1532 (N_1532,In_1449,In_1000);
or U1533 (N_1533,In_1292,In_213);
nor U1534 (N_1534,In_390,In_890);
nand U1535 (N_1535,In_497,In_1358);
or U1536 (N_1536,In_743,In_502);
nor U1537 (N_1537,In_526,In_382);
nand U1538 (N_1538,In_337,In_501);
and U1539 (N_1539,In_100,In_1096);
and U1540 (N_1540,In_1017,In_578);
and U1541 (N_1541,In_50,In_626);
or U1542 (N_1542,In_893,In_1073);
or U1543 (N_1543,In_799,In_1091);
nor U1544 (N_1544,In_1425,In_1325);
and U1545 (N_1545,In_1112,In_485);
nand U1546 (N_1546,In_483,In_454);
or U1547 (N_1547,In_986,In_854);
nor U1548 (N_1548,In_404,In_1320);
nor U1549 (N_1549,In_815,In_937);
nor U1550 (N_1550,In_1095,In_284);
or U1551 (N_1551,In_1185,In_548);
or U1552 (N_1552,In_816,In_1335);
or U1553 (N_1553,In_137,In_1454);
or U1554 (N_1554,In_9,In_1402);
nand U1555 (N_1555,In_855,In_529);
nor U1556 (N_1556,In_1248,In_783);
or U1557 (N_1557,In_284,In_116);
and U1558 (N_1558,In_1470,In_317);
nand U1559 (N_1559,In_1206,In_376);
nor U1560 (N_1560,In_219,In_736);
or U1561 (N_1561,In_690,In_1200);
or U1562 (N_1562,In_167,In_1252);
and U1563 (N_1563,In_243,In_460);
nand U1564 (N_1564,In_1108,In_1296);
and U1565 (N_1565,In_849,In_141);
or U1566 (N_1566,In_539,In_681);
and U1567 (N_1567,In_1368,In_167);
or U1568 (N_1568,In_391,In_300);
or U1569 (N_1569,In_185,In_384);
nor U1570 (N_1570,In_1392,In_1150);
and U1571 (N_1571,In_850,In_941);
and U1572 (N_1572,In_1302,In_1150);
and U1573 (N_1573,In_651,In_1482);
nor U1574 (N_1574,In_1203,In_433);
and U1575 (N_1575,In_859,In_56);
and U1576 (N_1576,In_723,In_4);
nand U1577 (N_1577,In_155,In_968);
nand U1578 (N_1578,In_1054,In_1407);
nor U1579 (N_1579,In_386,In_784);
nor U1580 (N_1580,In_849,In_848);
and U1581 (N_1581,In_478,In_54);
or U1582 (N_1582,In_1077,In_659);
nor U1583 (N_1583,In_595,In_1104);
or U1584 (N_1584,In_952,In_773);
nand U1585 (N_1585,In_1225,In_885);
nor U1586 (N_1586,In_1327,In_1322);
nand U1587 (N_1587,In_200,In_1052);
nand U1588 (N_1588,In_750,In_1358);
or U1589 (N_1589,In_562,In_94);
nor U1590 (N_1590,In_82,In_1126);
nor U1591 (N_1591,In_739,In_749);
nand U1592 (N_1592,In_602,In_1415);
or U1593 (N_1593,In_173,In_1084);
or U1594 (N_1594,In_1161,In_631);
nor U1595 (N_1595,In_480,In_555);
or U1596 (N_1596,In_1193,In_426);
or U1597 (N_1597,In_1338,In_965);
and U1598 (N_1598,In_303,In_1324);
and U1599 (N_1599,In_903,In_829);
nor U1600 (N_1600,In_1,In_374);
and U1601 (N_1601,In_654,In_386);
and U1602 (N_1602,In_73,In_1356);
xor U1603 (N_1603,In_1440,In_803);
and U1604 (N_1604,In_56,In_388);
or U1605 (N_1605,In_129,In_412);
or U1606 (N_1606,In_239,In_880);
and U1607 (N_1607,In_1474,In_1043);
and U1608 (N_1608,In_1297,In_1205);
nand U1609 (N_1609,In_650,In_1344);
and U1610 (N_1610,In_1075,In_802);
and U1611 (N_1611,In_916,In_1132);
nor U1612 (N_1612,In_1212,In_1186);
and U1613 (N_1613,In_490,In_390);
nor U1614 (N_1614,In_409,In_280);
nor U1615 (N_1615,In_848,In_305);
and U1616 (N_1616,In_1468,In_601);
and U1617 (N_1617,In_1476,In_213);
or U1618 (N_1618,In_555,In_128);
nand U1619 (N_1619,In_347,In_289);
and U1620 (N_1620,In_494,In_465);
nand U1621 (N_1621,In_119,In_591);
nand U1622 (N_1622,In_883,In_912);
nor U1623 (N_1623,In_228,In_1386);
or U1624 (N_1624,In_1482,In_625);
nor U1625 (N_1625,In_580,In_1002);
nor U1626 (N_1626,In_45,In_608);
or U1627 (N_1627,In_1056,In_135);
or U1628 (N_1628,In_132,In_647);
and U1629 (N_1629,In_1089,In_272);
and U1630 (N_1630,In_967,In_832);
nor U1631 (N_1631,In_775,In_640);
and U1632 (N_1632,In_1017,In_101);
and U1633 (N_1633,In_762,In_1229);
or U1634 (N_1634,In_927,In_1455);
or U1635 (N_1635,In_606,In_1077);
nand U1636 (N_1636,In_1044,In_147);
nor U1637 (N_1637,In_457,In_616);
nor U1638 (N_1638,In_116,In_441);
and U1639 (N_1639,In_1151,In_858);
nor U1640 (N_1640,In_1108,In_817);
nand U1641 (N_1641,In_356,In_7);
nand U1642 (N_1642,In_701,In_1226);
or U1643 (N_1643,In_904,In_224);
and U1644 (N_1644,In_129,In_1368);
nor U1645 (N_1645,In_67,In_336);
nor U1646 (N_1646,In_382,In_1135);
nand U1647 (N_1647,In_626,In_290);
or U1648 (N_1648,In_1291,In_1014);
nand U1649 (N_1649,In_777,In_1285);
or U1650 (N_1650,In_913,In_172);
nand U1651 (N_1651,In_661,In_869);
xnor U1652 (N_1652,In_1123,In_881);
and U1653 (N_1653,In_273,In_1469);
nand U1654 (N_1654,In_1425,In_626);
or U1655 (N_1655,In_179,In_837);
nor U1656 (N_1656,In_627,In_1216);
or U1657 (N_1657,In_132,In_835);
and U1658 (N_1658,In_544,In_312);
and U1659 (N_1659,In_683,In_887);
or U1660 (N_1660,In_236,In_820);
nand U1661 (N_1661,In_596,In_1093);
nand U1662 (N_1662,In_1147,In_501);
nor U1663 (N_1663,In_1433,In_1200);
nor U1664 (N_1664,In_328,In_1255);
or U1665 (N_1665,In_138,In_1358);
nand U1666 (N_1666,In_415,In_933);
or U1667 (N_1667,In_870,In_195);
or U1668 (N_1668,In_978,In_691);
or U1669 (N_1669,In_1438,In_175);
nor U1670 (N_1670,In_1077,In_644);
or U1671 (N_1671,In_1131,In_355);
nor U1672 (N_1672,In_666,In_1416);
nor U1673 (N_1673,In_908,In_444);
or U1674 (N_1674,In_1023,In_1401);
and U1675 (N_1675,In_850,In_159);
and U1676 (N_1676,In_182,In_222);
nor U1677 (N_1677,In_606,In_1401);
or U1678 (N_1678,In_1270,In_578);
nor U1679 (N_1679,In_330,In_1142);
and U1680 (N_1680,In_333,In_825);
nand U1681 (N_1681,In_1247,In_688);
nor U1682 (N_1682,In_986,In_984);
nor U1683 (N_1683,In_714,In_1253);
nand U1684 (N_1684,In_934,In_58);
nand U1685 (N_1685,In_153,In_42);
and U1686 (N_1686,In_816,In_57);
and U1687 (N_1687,In_357,In_825);
or U1688 (N_1688,In_741,In_1125);
nand U1689 (N_1689,In_20,In_314);
and U1690 (N_1690,In_1336,In_826);
nand U1691 (N_1691,In_451,In_223);
nand U1692 (N_1692,In_754,In_554);
nor U1693 (N_1693,In_784,In_22);
or U1694 (N_1694,In_402,In_1258);
nand U1695 (N_1695,In_679,In_152);
nand U1696 (N_1696,In_1013,In_1415);
or U1697 (N_1697,In_1431,In_1426);
and U1698 (N_1698,In_564,In_1483);
and U1699 (N_1699,In_711,In_298);
or U1700 (N_1700,In_1070,In_768);
and U1701 (N_1701,In_32,In_1156);
nand U1702 (N_1702,In_734,In_953);
nand U1703 (N_1703,In_956,In_478);
and U1704 (N_1704,In_405,In_909);
or U1705 (N_1705,In_827,In_162);
nor U1706 (N_1706,In_293,In_1332);
nand U1707 (N_1707,In_231,In_599);
and U1708 (N_1708,In_1216,In_213);
or U1709 (N_1709,In_1348,In_366);
or U1710 (N_1710,In_1002,In_401);
and U1711 (N_1711,In_1045,In_1344);
or U1712 (N_1712,In_1162,In_525);
and U1713 (N_1713,In_26,In_823);
or U1714 (N_1714,In_630,In_92);
nand U1715 (N_1715,In_1098,In_3);
or U1716 (N_1716,In_651,In_942);
nand U1717 (N_1717,In_1193,In_1343);
and U1718 (N_1718,In_467,In_1285);
nand U1719 (N_1719,In_1029,In_1352);
nand U1720 (N_1720,In_1296,In_1136);
and U1721 (N_1721,In_1186,In_1315);
and U1722 (N_1722,In_355,In_911);
nor U1723 (N_1723,In_662,In_412);
nor U1724 (N_1724,In_1415,In_646);
nor U1725 (N_1725,In_789,In_402);
or U1726 (N_1726,In_1130,In_1172);
nor U1727 (N_1727,In_1481,In_634);
nor U1728 (N_1728,In_927,In_558);
nor U1729 (N_1729,In_1153,In_842);
or U1730 (N_1730,In_1059,In_444);
or U1731 (N_1731,In_1383,In_379);
nor U1732 (N_1732,In_1374,In_1477);
nand U1733 (N_1733,In_1233,In_386);
nand U1734 (N_1734,In_824,In_1397);
nand U1735 (N_1735,In_1037,In_1157);
nand U1736 (N_1736,In_1356,In_868);
nor U1737 (N_1737,In_117,In_629);
and U1738 (N_1738,In_632,In_479);
or U1739 (N_1739,In_299,In_1110);
nand U1740 (N_1740,In_799,In_1296);
nand U1741 (N_1741,In_555,In_56);
and U1742 (N_1742,In_1130,In_973);
nand U1743 (N_1743,In_1054,In_1486);
nand U1744 (N_1744,In_209,In_1094);
and U1745 (N_1745,In_989,In_1111);
nor U1746 (N_1746,In_997,In_876);
nand U1747 (N_1747,In_454,In_717);
nor U1748 (N_1748,In_653,In_456);
or U1749 (N_1749,In_111,In_247);
or U1750 (N_1750,In_1459,In_828);
and U1751 (N_1751,In_259,In_475);
and U1752 (N_1752,In_1140,In_1127);
nand U1753 (N_1753,In_981,In_3);
nand U1754 (N_1754,In_1250,In_1417);
and U1755 (N_1755,In_1297,In_1462);
and U1756 (N_1756,In_869,In_1268);
or U1757 (N_1757,In_279,In_506);
nor U1758 (N_1758,In_917,In_1202);
or U1759 (N_1759,In_329,In_85);
and U1760 (N_1760,In_371,In_26);
or U1761 (N_1761,In_1085,In_1356);
or U1762 (N_1762,In_207,In_324);
or U1763 (N_1763,In_37,In_892);
nand U1764 (N_1764,In_116,In_591);
nand U1765 (N_1765,In_1473,In_241);
and U1766 (N_1766,In_55,In_588);
nand U1767 (N_1767,In_21,In_563);
nor U1768 (N_1768,In_181,In_388);
nand U1769 (N_1769,In_457,In_128);
and U1770 (N_1770,In_292,In_1200);
nor U1771 (N_1771,In_1063,In_5);
or U1772 (N_1772,In_85,In_767);
nor U1773 (N_1773,In_1491,In_157);
nand U1774 (N_1774,In_589,In_574);
nor U1775 (N_1775,In_102,In_515);
or U1776 (N_1776,In_1417,In_1482);
and U1777 (N_1777,In_803,In_346);
and U1778 (N_1778,In_1466,In_1208);
nand U1779 (N_1779,In_1352,In_703);
and U1780 (N_1780,In_90,In_1433);
or U1781 (N_1781,In_1170,In_1300);
and U1782 (N_1782,In_340,In_748);
nor U1783 (N_1783,In_1452,In_774);
or U1784 (N_1784,In_184,In_1051);
nor U1785 (N_1785,In_273,In_1394);
and U1786 (N_1786,In_403,In_247);
and U1787 (N_1787,In_541,In_1085);
nand U1788 (N_1788,In_1044,In_414);
nor U1789 (N_1789,In_1192,In_1096);
and U1790 (N_1790,In_345,In_1036);
nor U1791 (N_1791,In_164,In_1092);
xor U1792 (N_1792,In_399,In_900);
and U1793 (N_1793,In_461,In_1136);
nor U1794 (N_1794,In_976,In_88);
nand U1795 (N_1795,In_408,In_1358);
nand U1796 (N_1796,In_835,In_844);
nor U1797 (N_1797,In_752,In_457);
nand U1798 (N_1798,In_404,In_817);
and U1799 (N_1799,In_661,In_1335);
or U1800 (N_1800,In_130,In_1366);
and U1801 (N_1801,In_1101,In_276);
or U1802 (N_1802,In_1137,In_856);
and U1803 (N_1803,In_1095,In_540);
nor U1804 (N_1804,In_406,In_617);
and U1805 (N_1805,In_1475,In_519);
nand U1806 (N_1806,In_1463,In_689);
and U1807 (N_1807,In_935,In_1103);
and U1808 (N_1808,In_647,In_799);
or U1809 (N_1809,In_1179,In_1017);
nor U1810 (N_1810,In_95,In_69);
or U1811 (N_1811,In_1407,In_155);
or U1812 (N_1812,In_920,In_1481);
and U1813 (N_1813,In_849,In_183);
nor U1814 (N_1814,In_1200,In_1396);
or U1815 (N_1815,In_364,In_311);
nor U1816 (N_1816,In_673,In_808);
and U1817 (N_1817,In_113,In_37);
and U1818 (N_1818,In_866,In_1236);
nor U1819 (N_1819,In_1003,In_1192);
nor U1820 (N_1820,In_1060,In_509);
and U1821 (N_1821,In_336,In_1259);
or U1822 (N_1822,In_1187,In_954);
or U1823 (N_1823,In_1269,In_2);
or U1824 (N_1824,In_470,In_516);
or U1825 (N_1825,In_703,In_84);
nor U1826 (N_1826,In_107,In_820);
nor U1827 (N_1827,In_277,In_598);
nor U1828 (N_1828,In_1450,In_810);
nor U1829 (N_1829,In_1349,In_1204);
and U1830 (N_1830,In_574,In_444);
or U1831 (N_1831,In_454,In_16);
or U1832 (N_1832,In_891,In_376);
or U1833 (N_1833,In_365,In_1010);
nor U1834 (N_1834,In_1430,In_1472);
nand U1835 (N_1835,In_1302,In_291);
or U1836 (N_1836,In_1049,In_1130);
nand U1837 (N_1837,In_160,In_880);
nand U1838 (N_1838,In_631,In_638);
or U1839 (N_1839,In_1374,In_90);
nand U1840 (N_1840,In_1304,In_826);
nor U1841 (N_1841,In_1145,In_717);
nand U1842 (N_1842,In_964,In_1252);
or U1843 (N_1843,In_1127,In_530);
and U1844 (N_1844,In_96,In_888);
nor U1845 (N_1845,In_1395,In_491);
or U1846 (N_1846,In_994,In_728);
and U1847 (N_1847,In_428,In_468);
and U1848 (N_1848,In_139,In_60);
or U1849 (N_1849,In_1237,In_1154);
nor U1850 (N_1850,In_137,In_140);
nor U1851 (N_1851,In_1316,In_396);
nor U1852 (N_1852,In_1179,In_990);
nor U1853 (N_1853,In_407,In_1476);
nand U1854 (N_1854,In_551,In_93);
nand U1855 (N_1855,In_1485,In_889);
nor U1856 (N_1856,In_734,In_458);
nand U1857 (N_1857,In_48,In_322);
or U1858 (N_1858,In_1011,In_146);
or U1859 (N_1859,In_336,In_515);
nor U1860 (N_1860,In_434,In_132);
nor U1861 (N_1861,In_820,In_339);
nor U1862 (N_1862,In_540,In_29);
and U1863 (N_1863,In_921,In_71);
nor U1864 (N_1864,In_201,In_449);
xor U1865 (N_1865,In_763,In_10);
nand U1866 (N_1866,In_1204,In_1373);
or U1867 (N_1867,In_1044,In_347);
or U1868 (N_1868,In_142,In_788);
and U1869 (N_1869,In_397,In_1176);
nor U1870 (N_1870,In_175,In_1182);
or U1871 (N_1871,In_1060,In_323);
or U1872 (N_1872,In_931,In_67);
nor U1873 (N_1873,In_374,In_587);
nand U1874 (N_1874,In_824,In_978);
and U1875 (N_1875,In_1011,In_628);
nand U1876 (N_1876,In_645,In_1351);
nand U1877 (N_1877,In_1374,In_1145);
or U1878 (N_1878,In_630,In_1427);
nor U1879 (N_1879,In_1431,In_752);
and U1880 (N_1880,In_150,In_760);
and U1881 (N_1881,In_1005,In_671);
or U1882 (N_1882,In_1290,In_1218);
nand U1883 (N_1883,In_1330,In_1417);
nor U1884 (N_1884,In_725,In_264);
and U1885 (N_1885,In_630,In_457);
nand U1886 (N_1886,In_436,In_974);
nor U1887 (N_1887,In_572,In_815);
nand U1888 (N_1888,In_685,In_1158);
and U1889 (N_1889,In_857,In_1496);
nand U1890 (N_1890,In_281,In_1429);
nor U1891 (N_1891,In_722,In_296);
nand U1892 (N_1892,In_225,In_134);
or U1893 (N_1893,In_1200,In_1355);
and U1894 (N_1894,In_547,In_419);
and U1895 (N_1895,In_1346,In_1275);
and U1896 (N_1896,In_410,In_821);
or U1897 (N_1897,In_778,In_528);
or U1898 (N_1898,In_1254,In_753);
or U1899 (N_1899,In_272,In_257);
or U1900 (N_1900,In_1362,In_270);
or U1901 (N_1901,In_1115,In_1077);
or U1902 (N_1902,In_1050,In_1024);
or U1903 (N_1903,In_597,In_719);
and U1904 (N_1904,In_604,In_129);
and U1905 (N_1905,In_797,In_1414);
and U1906 (N_1906,In_314,In_360);
nand U1907 (N_1907,In_1494,In_1456);
or U1908 (N_1908,In_1184,In_683);
or U1909 (N_1909,In_350,In_998);
nand U1910 (N_1910,In_1338,In_1359);
nor U1911 (N_1911,In_227,In_455);
and U1912 (N_1912,In_934,In_1420);
nor U1913 (N_1913,In_421,In_412);
nand U1914 (N_1914,In_1247,In_1359);
nand U1915 (N_1915,In_454,In_848);
nor U1916 (N_1916,In_999,In_184);
nand U1917 (N_1917,In_11,In_541);
nand U1918 (N_1918,In_1392,In_386);
and U1919 (N_1919,In_538,In_89);
or U1920 (N_1920,In_582,In_486);
or U1921 (N_1921,In_1123,In_1149);
and U1922 (N_1922,In_553,In_1398);
nand U1923 (N_1923,In_329,In_1284);
nor U1924 (N_1924,In_766,In_158);
and U1925 (N_1925,In_634,In_1340);
nor U1926 (N_1926,In_316,In_1425);
nor U1927 (N_1927,In_447,In_33);
nor U1928 (N_1928,In_102,In_444);
or U1929 (N_1929,In_224,In_655);
and U1930 (N_1930,In_726,In_1155);
nand U1931 (N_1931,In_568,In_1430);
nand U1932 (N_1932,In_743,In_957);
nor U1933 (N_1933,In_445,In_1181);
nor U1934 (N_1934,In_1285,In_1307);
or U1935 (N_1935,In_1205,In_456);
and U1936 (N_1936,In_681,In_8);
nand U1937 (N_1937,In_1264,In_813);
or U1938 (N_1938,In_907,In_218);
or U1939 (N_1939,In_868,In_387);
and U1940 (N_1940,In_59,In_717);
and U1941 (N_1941,In_550,In_1386);
nor U1942 (N_1942,In_1078,In_69);
and U1943 (N_1943,In_811,In_45);
nand U1944 (N_1944,In_17,In_687);
and U1945 (N_1945,In_509,In_1108);
or U1946 (N_1946,In_718,In_285);
or U1947 (N_1947,In_1330,In_1389);
nand U1948 (N_1948,In_312,In_1054);
nand U1949 (N_1949,In_870,In_1038);
and U1950 (N_1950,In_161,In_18);
and U1951 (N_1951,In_551,In_1361);
and U1952 (N_1952,In_325,In_195);
xnor U1953 (N_1953,In_744,In_732);
and U1954 (N_1954,In_1373,In_865);
or U1955 (N_1955,In_684,In_449);
nor U1956 (N_1956,In_331,In_133);
nor U1957 (N_1957,In_745,In_1017);
or U1958 (N_1958,In_1147,In_750);
and U1959 (N_1959,In_685,In_53);
or U1960 (N_1960,In_784,In_148);
nor U1961 (N_1961,In_1088,In_192);
or U1962 (N_1962,In_1106,In_999);
or U1963 (N_1963,In_490,In_983);
or U1964 (N_1964,In_1371,In_1064);
nand U1965 (N_1965,In_306,In_614);
or U1966 (N_1966,In_714,In_277);
and U1967 (N_1967,In_98,In_1321);
nand U1968 (N_1968,In_1000,In_606);
or U1969 (N_1969,In_81,In_1233);
or U1970 (N_1970,In_1434,In_1211);
xor U1971 (N_1971,In_1164,In_835);
and U1972 (N_1972,In_463,In_861);
nand U1973 (N_1973,In_1399,In_524);
nand U1974 (N_1974,In_671,In_194);
nand U1975 (N_1975,In_744,In_1221);
nand U1976 (N_1976,In_948,In_318);
or U1977 (N_1977,In_1073,In_673);
and U1978 (N_1978,In_685,In_459);
nor U1979 (N_1979,In_287,In_310);
nand U1980 (N_1980,In_793,In_1146);
nand U1981 (N_1981,In_1239,In_861);
nor U1982 (N_1982,In_1125,In_248);
nor U1983 (N_1983,In_336,In_799);
or U1984 (N_1984,In_812,In_352);
nor U1985 (N_1985,In_1477,In_807);
nor U1986 (N_1986,In_1195,In_1249);
nor U1987 (N_1987,In_565,In_711);
and U1988 (N_1988,In_1191,In_722);
nand U1989 (N_1989,In_845,In_452);
or U1990 (N_1990,In_884,In_20);
nor U1991 (N_1991,In_35,In_1072);
nand U1992 (N_1992,In_592,In_1145);
nand U1993 (N_1993,In_808,In_775);
nor U1994 (N_1994,In_905,In_284);
nand U1995 (N_1995,In_453,In_422);
and U1996 (N_1996,In_153,In_162);
nor U1997 (N_1997,In_79,In_404);
and U1998 (N_1998,In_1038,In_284);
nor U1999 (N_1999,In_526,In_760);
or U2000 (N_2000,In_130,In_61);
nor U2001 (N_2001,In_1000,In_219);
and U2002 (N_2002,In_1127,In_155);
nor U2003 (N_2003,In_18,In_17);
nor U2004 (N_2004,In_1417,In_1096);
nand U2005 (N_2005,In_527,In_1258);
xnor U2006 (N_2006,In_1165,In_765);
or U2007 (N_2007,In_459,In_1083);
and U2008 (N_2008,In_464,In_821);
nand U2009 (N_2009,In_54,In_980);
and U2010 (N_2010,In_1487,In_240);
nand U2011 (N_2011,In_365,In_559);
and U2012 (N_2012,In_672,In_230);
nand U2013 (N_2013,In_99,In_507);
nand U2014 (N_2014,In_1023,In_785);
and U2015 (N_2015,In_354,In_1081);
nor U2016 (N_2016,In_671,In_260);
or U2017 (N_2017,In_936,In_843);
nor U2018 (N_2018,In_655,In_660);
nand U2019 (N_2019,In_1256,In_1184);
or U2020 (N_2020,In_264,In_1250);
nand U2021 (N_2021,In_1253,In_596);
nand U2022 (N_2022,In_993,In_1152);
and U2023 (N_2023,In_1438,In_240);
nand U2024 (N_2024,In_1039,In_863);
nor U2025 (N_2025,In_443,In_571);
or U2026 (N_2026,In_626,In_1299);
and U2027 (N_2027,In_885,In_1442);
xor U2028 (N_2028,In_987,In_533);
or U2029 (N_2029,In_96,In_220);
or U2030 (N_2030,In_1033,In_1489);
and U2031 (N_2031,In_4,In_1044);
or U2032 (N_2032,In_54,In_1213);
or U2033 (N_2033,In_768,In_1428);
nor U2034 (N_2034,In_129,In_120);
nor U2035 (N_2035,In_486,In_1481);
nand U2036 (N_2036,In_868,In_927);
and U2037 (N_2037,In_36,In_60);
nor U2038 (N_2038,In_1341,In_1007);
and U2039 (N_2039,In_1194,In_13);
and U2040 (N_2040,In_1488,In_1044);
and U2041 (N_2041,In_968,In_749);
or U2042 (N_2042,In_316,In_1306);
nor U2043 (N_2043,In_891,In_1251);
nor U2044 (N_2044,In_652,In_107);
nand U2045 (N_2045,In_817,In_352);
nand U2046 (N_2046,In_677,In_169);
nand U2047 (N_2047,In_314,In_92);
or U2048 (N_2048,In_444,In_168);
nand U2049 (N_2049,In_67,In_709);
nand U2050 (N_2050,In_1173,In_1451);
and U2051 (N_2051,In_929,In_1114);
nand U2052 (N_2052,In_417,In_799);
or U2053 (N_2053,In_1026,In_156);
and U2054 (N_2054,In_387,In_79);
and U2055 (N_2055,In_581,In_484);
nand U2056 (N_2056,In_1120,In_256);
nand U2057 (N_2057,In_628,In_281);
nor U2058 (N_2058,In_554,In_726);
or U2059 (N_2059,In_1333,In_206);
nor U2060 (N_2060,In_1245,In_1084);
nor U2061 (N_2061,In_1065,In_121);
and U2062 (N_2062,In_597,In_729);
and U2063 (N_2063,In_561,In_1492);
and U2064 (N_2064,In_400,In_337);
or U2065 (N_2065,In_346,In_873);
nor U2066 (N_2066,In_862,In_468);
or U2067 (N_2067,In_1487,In_502);
and U2068 (N_2068,In_703,In_43);
nor U2069 (N_2069,In_859,In_520);
or U2070 (N_2070,In_1181,In_845);
nor U2071 (N_2071,In_114,In_932);
and U2072 (N_2072,In_1456,In_311);
or U2073 (N_2073,In_1433,In_1491);
nand U2074 (N_2074,In_210,In_1311);
or U2075 (N_2075,In_472,In_1078);
and U2076 (N_2076,In_248,In_1077);
or U2077 (N_2077,In_281,In_1018);
xnor U2078 (N_2078,In_1106,In_292);
or U2079 (N_2079,In_732,In_88);
nand U2080 (N_2080,In_1035,In_472);
and U2081 (N_2081,In_313,In_662);
or U2082 (N_2082,In_548,In_899);
or U2083 (N_2083,In_1006,In_1189);
nand U2084 (N_2084,In_487,In_920);
and U2085 (N_2085,In_1455,In_596);
or U2086 (N_2086,In_1257,In_754);
or U2087 (N_2087,In_430,In_1229);
or U2088 (N_2088,In_1045,In_788);
and U2089 (N_2089,In_362,In_564);
and U2090 (N_2090,In_551,In_1163);
nor U2091 (N_2091,In_1252,In_741);
or U2092 (N_2092,In_349,In_690);
nand U2093 (N_2093,In_104,In_1063);
and U2094 (N_2094,In_246,In_1081);
and U2095 (N_2095,In_334,In_206);
nor U2096 (N_2096,In_555,In_810);
nand U2097 (N_2097,In_733,In_1005);
nor U2098 (N_2098,In_1394,In_1440);
nand U2099 (N_2099,In_1474,In_45);
and U2100 (N_2100,In_553,In_223);
nor U2101 (N_2101,In_89,In_1057);
nand U2102 (N_2102,In_928,In_250);
and U2103 (N_2103,In_45,In_787);
nor U2104 (N_2104,In_802,In_132);
nor U2105 (N_2105,In_1463,In_12);
nor U2106 (N_2106,In_379,In_975);
nand U2107 (N_2107,In_52,In_911);
nor U2108 (N_2108,In_1368,In_300);
nor U2109 (N_2109,In_818,In_489);
nor U2110 (N_2110,In_1490,In_363);
nand U2111 (N_2111,In_520,In_1228);
and U2112 (N_2112,In_468,In_654);
or U2113 (N_2113,In_482,In_874);
or U2114 (N_2114,In_738,In_650);
nor U2115 (N_2115,In_124,In_293);
nor U2116 (N_2116,In_973,In_726);
nand U2117 (N_2117,In_1145,In_412);
and U2118 (N_2118,In_26,In_1443);
nand U2119 (N_2119,In_197,In_1452);
nand U2120 (N_2120,In_1078,In_712);
or U2121 (N_2121,In_1448,In_642);
and U2122 (N_2122,In_1267,In_1069);
nor U2123 (N_2123,In_1083,In_397);
nor U2124 (N_2124,In_696,In_562);
or U2125 (N_2125,In_1281,In_348);
and U2126 (N_2126,In_986,In_800);
and U2127 (N_2127,In_247,In_54);
nand U2128 (N_2128,In_149,In_1436);
or U2129 (N_2129,In_1376,In_980);
or U2130 (N_2130,In_575,In_651);
nand U2131 (N_2131,In_1487,In_567);
or U2132 (N_2132,In_1178,In_484);
xnor U2133 (N_2133,In_74,In_797);
and U2134 (N_2134,In_240,In_319);
and U2135 (N_2135,In_989,In_378);
nand U2136 (N_2136,In_724,In_407);
nor U2137 (N_2137,In_1211,In_1495);
nand U2138 (N_2138,In_1283,In_28);
or U2139 (N_2139,In_1125,In_1225);
nand U2140 (N_2140,In_154,In_1180);
or U2141 (N_2141,In_1289,In_948);
nor U2142 (N_2142,In_246,In_1061);
nand U2143 (N_2143,In_566,In_1417);
nor U2144 (N_2144,In_546,In_39);
nor U2145 (N_2145,In_1352,In_1201);
nor U2146 (N_2146,In_1165,In_545);
nor U2147 (N_2147,In_451,In_514);
and U2148 (N_2148,In_59,In_669);
and U2149 (N_2149,In_6,In_555);
nand U2150 (N_2150,In_325,In_1027);
and U2151 (N_2151,In_1077,In_396);
and U2152 (N_2152,In_912,In_1123);
nor U2153 (N_2153,In_113,In_1059);
or U2154 (N_2154,In_157,In_976);
xor U2155 (N_2155,In_62,In_1143);
nand U2156 (N_2156,In_859,In_394);
or U2157 (N_2157,In_1212,In_615);
nand U2158 (N_2158,In_790,In_1204);
and U2159 (N_2159,In_41,In_334);
nand U2160 (N_2160,In_371,In_1344);
and U2161 (N_2161,In_435,In_514);
nand U2162 (N_2162,In_1299,In_1390);
and U2163 (N_2163,In_604,In_444);
nand U2164 (N_2164,In_747,In_491);
or U2165 (N_2165,In_90,In_634);
nor U2166 (N_2166,In_1492,In_621);
or U2167 (N_2167,In_374,In_910);
and U2168 (N_2168,In_591,In_1303);
xor U2169 (N_2169,In_70,In_678);
nor U2170 (N_2170,In_739,In_1238);
nor U2171 (N_2171,In_1136,In_399);
and U2172 (N_2172,In_1388,In_479);
and U2173 (N_2173,In_616,In_537);
and U2174 (N_2174,In_1025,In_724);
nor U2175 (N_2175,In_397,In_904);
nor U2176 (N_2176,In_471,In_1312);
or U2177 (N_2177,In_46,In_379);
and U2178 (N_2178,In_921,In_1238);
xnor U2179 (N_2179,In_1468,In_138);
and U2180 (N_2180,In_795,In_373);
nand U2181 (N_2181,In_1059,In_1394);
xnor U2182 (N_2182,In_352,In_1201);
or U2183 (N_2183,In_21,In_1305);
nand U2184 (N_2184,In_1492,In_338);
and U2185 (N_2185,In_177,In_415);
and U2186 (N_2186,In_609,In_361);
and U2187 (N_2187,In_1194,In_1061);
and U2188 (N_2188,In_452,In_210);
or U2189 (N_2189,In_1012,In_692);
or U2190 (N_2190,In_1326,In_129);
nand U2191 (N_2191,In_1040,In_388);
xnor U2192 (N_2192,In_339,In_424);
or U2193 (N_2193,In_893,In_48);
and U2194 (N_2194,In_1215,In_918);
nor U2195 (N_2195,In_953,In_838);
and U2196 (N_2196,In_417,In_621);
and U2197 (N_2197,In_1263,In_885);
or U2198 (N_2198,In_341,In_1050);
or U2199 (N_2199,In_1226,In_1264);
nor U2200 (N_2200,In_757,In_43);
and U2201 (N_2201,In_1387,In_864);
and U2202 (N_2202,In_355,In_479);
and U2203 (N_2203,In_415,In_1076);
and U2204 (N_2204,In_1429,In_769);
and U2205 (N_2205,In_1155,In_1067);
or U2206 (N_2206,In_495,In_1216);
or U2207 (N_2207,In_876,In_177);
nor U2208 (N_2208,In_123,In_1076);
or U2209 (N_2209,In_475,In_533);
or U2210 (N_2210,In_823,In_413);
and U2211 (N_2211,In_571,In_568);
nand U2212 (N_2212,In_1386,In_695);
nor U2213 (N_2213,In_117,In_699);
and U2214 (N_2214,In_33,In_1003);
and U2215 (N_2215,In_375,In_1087);
nand U2216 (N_2216,In_93,In_1146);
or U2217 (N_2217,In_72,In_839);
and U2218 (N_2218,In_1235,In_1021);
nor U2219 (N_2219,In_1176,In_1006);
nand U2220 (N_2220,In_1472,In_798);
or U2221 (N_2221,In_936,In_183);
or U2222 (N_2222,In_1289,In_228);
nor U2223 (N_2223,In_835,In_336);
and U2224 (N_2224,In_832,In_1288);
or U2225 (N_2225,In_854,In_390);
and U2226 (N_2226,In_1197,In_681);
and U2227 (N_2227,In_287,In_770);
or U2228 (N_2228,In_1160,In_727);
nand U2229 (N_2229,In_764,In_629);
and U2230 (N_2230,In_143,In_713);
or U2231 (N_2231,In_852,In_1081);
nor U2232 (N_2232,In_361,In_315);
or U2233 (N_2233,In_542,In_1063);
nand U2234 (N_2234,In_493,In_783);
nand U2235 (N_2235,In_756,In_1113);
and U2236 (N_2236,In_72,In_1488);
nor U2237 (N_2237,In_834,In_806);
nand U2238 (N_2238,In_1191,In_384);
or U2239 (N_2239,In_626,In_995);
and U2240 (N_2240,In_918,In_652);
and U2241 (N_2241,In_1059,In_431);
or U2242 (N_2242,In_1345,In_1149);
nor U2243 (N_2243,In_351,In_449);
nor U2244 (N_2244,In_73,In_1137);
nand U2245 (N_2245,In_1036,In_128);
nor U2246 (N_2246,In_897,In_1490);
or U2247 (N_2247,In_311,In_1103);
or U2248 (N_2248,In_876,In_634);
nand U2249 (N_2249,In_527,In_631);
or U2250 (N_2250,In_38,In_268);
and U2251 (N_2251,In_493,In_1160);
and U2252 (N_2252,In_791,In_624);
and U2253 (N_2253,In_1478,In_546);
nand U2254 (N_2254,In_316,In_730);
and U2255 (N_2255,In_956,In_757);
or U2256 (N_2256,In_908,In_704);
nand U2257 (N_2257,In_785,In_1450);
nor U2258 (N_2258,In_1394,In_106);
xor U2259 (N_2259,In_177,In_784);
and U2260 (N_2260,In_1287,In_1474);
and U2261 (N_2261,In_1433,In_686);
nand U2262 (N_2262,In_256,In_57);
nand U2263 (N_2263,In_1122,In_294);
nand U2264 (N_2264,In_1108,In_1493);
or U2265 (N_2265,In_370,In_210);
and U2266 (N_2266,In_366,In_479);
and U2267 (N_2267,In_1179,In_1411);
nor U2268 (N_2268,In_1043,In_922);
or U2269 (N_2269,In_666,In_150);
nand U2270 (N_2270,In_212,In_1209);
or U2271 (N_2271,In_938,In_1160);
nor U2272 (N_2272,In_1138,In_204);
xor U2273 (N_2273,In_1457,In_1364);
nor U2274 (N_2274,In_190,In_733);
or U2275 (N_2275,In_1363,In_1199);
nand U2276 (N_2276,In_690,In_900);
and U2277 (N_2277,In_997,In_417);
nand U2278 (N_2278,In_731,In_341);
nor U2279 (N_2279,In_299,In_857);
nand U2280 (N_2280,In_255,In_1477);
nand U2281 (N_2281,In_746,In_616);
xnor U2282 (N_2282,In_1319,In_594);
or U2283 (N_2283,In_188,In_303);
and U2284 (N_2284,In_1429,In_278);
and U2285 (N_2285,In_397,In_465);
or U2286 (N_2286,In_566,In_1432);
or U2287 (N_2287,In_726,In_1278);
and U2288 (N_2288,In_1085,In_1367);
or U2289 (N_2289,In_776,In_202);
nor U2290 (N_2290,In_794,In_366);
nor U2291 (N_2291,In_1151,In_761);
nor U2292 (N_2292,In_688,In_1393);
or U2293 (N_2293,In_1313,In_1372);
nor U2294 (N_2294,In_113,In_353);
or U2295 (N_2295,In_847,In_92);
or U2296 (N_2296,In_1372,In_495);
and U2297 (N_2297,In_744,In_594);
or U2298 (N_2298,In_1155,In_430);
nor U2299 (N_2299,In_743,In_1274);
nor U2300 (N_2300,In_472,In_62);
nand U2301 (N_2301,In_191,In_102);
and U2302 (N_2302,In_1468,In_1308);
or U2303 (N_2303,In_1358,In_263);
or U2304 (N_2304,In_250,In_1339);
and U2305 (N_2305,In_430,In_684);
nand U2306 (N_2306,In_1095,In_1441);
nand U2307 (N_2307,In_1153,In_49);
nand U2308 (N_2308,In_1314,In_252);
nor U2309 (N_2309,In_338,In_289);
nor U2310 (N_2310,In_1342,In_840);
nand U2311 (N_2311,In_1175,In_1229);
nor U2312 (N_2312,In_81,In_1443);
or U2313 (N_2313,In_717,In_947);
and U2314 (N_2314,In_69,In_405);
or U2315 (N_2315,In_750,In_1155);
nand U2316 (N_2316,In_1425,In_1227);
xnor U2317 (N_2317,In_900,In_1451);
and U2318 (N_2318,In_660,In_1004);
nor U2319 (N_2319,In_1118,In_74);
or U2320 (N_2320,In_1440,In_54);
and U2321 (N_2321,In_927,In_972);
and U2322 (N_2322,In_1492,In_1291);
nor U2323 (N_2323,In_1371,In_533);
or U2324 (N_2324,In_271,In_1041);
and U2325 (N_2325,In_626,In_569);
xnor U2326 (N_2326,In_925,In_335);
nand U2327 (N_2327,In_93,In_300);
and U2328 (N_2328,In_1309,In_704);
and U2329 (N_2329,In_1218,In_682);
nor U2330 (N_2330,In_1044,In_423);
xor U2331 (N_2331,In_148,In_1449);
nand U2332 (N_2332,In_744,In_1425);
or U2333 (N_2333,In_1319,In_1135);
nor U2334 (N_2334,In_1064,In_1197);
and U2335 (N_2335,In_8,In_1414);
nor U2336 (N_2336,In_32,In_398);
nand U2337 (N_2337,In_798,In_833);
and U2338 (N_2338,In_891,In_1346);
and U2339 (N_2339,In_351,In_1011);
or U2340 (N_2340,In_519,In_295);
nor U2341 (N_2341,In_309,In_156);
nand U2342 (N_2342,In_897,In_978);
nand U2343 (N_2343,In_168,In_745);
or U2344 (N_2344,In_279,In_249);
and U2345 (N_2345,In_552,In_763);
nor U2346 (N_2346,In_160,In_115);
and U2347 (N_2347,In_1424,In_1361);
nand U2348 (N_2348,In_353,In_1477);
and U2349 (N_2349,In_245,In_1440);
or U2350 (N_2350,In_127,In_1410);
and U2351 (N_2351,In_1078,In_35);
or U2352 (N_2352,In_1309,In_698);
nand U2353 (N_2353,In_849,In_1088);
nor U2354 (N_2354,In_902,In_1166);
nor U2355 (N_2355,In_1173,In_759);
nand U2356 (N_2356,In_357,In_553);
nand U2357 (N_2357,In_350,In_1047);
nor U2358 (N_2358,In_663,In_593);
or U2359 (N_2359,In_19,In_858);
or U2360 (N_2360,In_498,In_153);
or U2361 (N_2361,In_1220,In_735);
or U2362 (N_2362,In_1263,In_768);
or U2363 (N_2363,In_118,In_551);
or U2364 (N_2364,In_332,In_309);
and U2365 (N_2365,In_101,In_480);
and U2366 (N_2366,In_748,In_560);
nand U2367 (N_2367,In_1448,In_1419);
and U2368 (N_2368,In_355,In_1052);
nand U2369 (N_2369,In_1076,In_826);
nor U2370 (N_2370,In_1071,In_494);
and U2371 (N_2371,In_579,In_50);
and U2372 (N_2372,In_409,In_625);
and U2373 (N_2373,In_342,In_595);
nor U2374 (N_2374,In_1205,In_106);
or U2375 (N_2375,In_285,In_199);
and U2376 (N_2376,In_1424,In_159);
nor U2377 (N_2377,In_874,In_309);
and U2378 (N_2378,In_88,In_1193);
nor U2379 (N_2379,In_43,In_1147);
and U2380 (N_2380,In_427,In_133);
nand U2381 (N_2381,In_767,In_1265);
or U2382 (N_2382,In_1467,In_1024);
and U2383 (N_2383,In_1222,In_631);
nor U2384 (N_2384,In_426,In_173);
nor U2385 (N_2385,In_1104,In_617);
or U2386 (N_2386,In_940,In_450);
and U2387 (N_2387,In_525,In_310);
and U2388 (N_2388,In_584,In_468);
and U2389 (N_2389,In_557,In_592);
nand U2390 (N_2390,In_1219,In_530);
and U2391 (N_2391,In_198,In_1251);
or U2392 (N_2392,In_428,In_1252);
nand U2393 (N_2393,In_1216,In_868);
nor U2394 (N_2394,In_168,In_872);
or U2395 (N_2395,In_1477,In_1014);
or U2396 (N_2396,In_434,In_448);
or U2397 (N_2397,In_376,In_1482);
nand U2398 (N_2398,In_721,In_94);
nor U2399 (N_2399,In_717,In_1280);
nand U2400 (N_2400,In_565,In_1351);
and U2401 (N_2401,In_836,In_1476);
nand U2402 (N_2402,In_1447,In_293);
nor U2403 (N_2403,In_558,In_254);
or U2404 (N_2404,In_1175,In_1336);
or U2405 (N_2405,In_762,In_309);
nor U2406 (N_2406,In_1455,In_581);
nand U2407 (N_2407,In_1421,In_1255);
nand U2408 (N_2408,In_1072,In_59);
nand U2409 (N_2409,In_630,In_799);
or U2410 (N_2410,In_231,In_338);
and U2411 (N_2411,In_541,In_1147);
nor U2412 (N_2412,In_1049,In_1154);
or U2413 (N_2413,In_1089,In_975);
or U2414 (N_2414,In_664,In_635);
and U2415 (N_2415,In_838,In_807);
nor U2416 (N_2416,In_262,In_645);
or U2417 (N_2417,In_1147,In_342);
nor U2418 (N_2418,In_255,In_857);
and U2419 (N_2419,In_972,In_653);
nand U2420 (N_2420,In_483,In_696);
or U2421 (N_2421,In_635,In_974);
nand U2422 (N_2422,In_545,In_261);
nand U2423 (N_2423,In_226,In_1313);
nor U2424 (N_2424,In_1275,In_1266);
nand U2425 (N_2425,In_1358,In_1009);
nor U2426 (N_2426,In_962,In_1244);
and U2427 (N_2427,In_529,In_62);
or U2428 (N_2428,In_334,In_1144);
nor U2429 (N_2429,In_457,In_297);
nor U2430 (N_2430,In_146,In_1405);
nand U2431 (N_2431,In_939,In_280);
nand U2432 (N_2432,In_43,In_299);
or U2433 (N_2433,In_196,In_1044);
or U2434 (N_2434,In_167,In_997);
xnor U2435 (N_2435,In_530,In_475);
and U2436 (N_2436,In_467,In_388);
or U2437 (N_2437,In_783,In_462);
or U2438 (N_2438,In_487,In_595);
and U2439 (N_2439,In_948,In_1165);
nor U2440 (N_2440,In_18,In_514);
or U2441 (N_2441,In_215,In_143);
nand U2442 (N_2442,In_237,In_1184);
or U2443 (N_2443,In_672,In_368);
nand U2444 (N_2444,In_125,In_75);
nor U2445 (N_2445,In_653,In_350);
nor U2446 (N_2446,In_869,In_1281);
nor U2447 (N_2447,In_239,In_1422);
or U2448 (N_2448,In_1201,In_53);
nand U2449 (N_2449,In_587,In_201);
nor U2450 (N_2450,In_421,In_302);
or U2451 (N_2451,In_696,In_838);
nand U2452 (N_2452,In_1401,In_588);
and U2453 (N_2453,In_204,In_149);
nand U2454 (N_2454,In_1347,In_1000);
or U2455 (N_2455,In_351,In_415);
or U2456 (N_2456,In_827,In_611);
or U2457 (N_2457,In_1108,In_397);
or U2458 (N_2458,In_524,In_1242);
or U2459 (N_2459,In_672,In_710);
nor U2460 (N_2460,In_1431,In_811);
or U2461 (N_2461,In_1167,In_1274);
xnor U2462 (N_2462,In_327,In_754);
and U2463 (N_2463,In_297,In_305);
and U2464 (N_2464,In_296,In_852);
nor U2465 (N_2465,In_542,In_1265);
nor U2466 (N_2466,In_206,In_1110);
or U2467 (N_2467,In_782,In_1257);
nand U2468 (N_2468,In_470,In_1448);
or U2469 (N_2469,In_368,In_778);
nand U2470 (N_2470,In_1331,In_115);
or U2471 (N_2471,In_243,In_590);
nor U2472 (N_2472,In_1291,In_669);
nor U2473 (N_2473,In_31,In_844);
or U2474 (N_2474,In_360,In_37);
and U2475 (N_2475,In_18,In_705);
nand U2476 (N_2476,In_486,In_461);
and U2477 (N_2477,In_1225,In_1123);
nor U2478 (N_2478,In_344,In_1119);
nor U2479 (N_2479,In_1349,In_632);
or U2480 (N_2480,In_558,In_344);
nor U2481 (N_2481,In_385,In_409);
nor U2482 (N_2482,In_29,In_1309);
nor U2483 (N_2483,In_1164,In_485);
and U2484 (N_2484,In_854,In_713);
nor U2485 (N_2485,In_685,In_957);
and U2486 (N_2486,In_1073,In_1052);
nand U2487 (N_2487,In_1320,In_153);
and U2488 (N_2488,In_1142,In_1152);
and U2489 (N_2489,In_919,In_1033);
or U2490 (N_2490,In_1153,In_1174);
nor U2491 (N_2491,In_236,In_1139);
and U2492 (N_2492,In_349,In_20);
nor U2493 (N_2493,In_89,In_1044);
nor U2494 (N_2494,In_513,In_1106);
nor U2495 (N_2495,In_650,In_862);
or U2496 (N_2496,In_1396,In_999);
and U2497 (N_2497,In_797,In_888);
and U2498 (N_2498,In_1352,In_691);
nand U2499 (N_2499,In_1206,In_883);
nand U2500 (N_2500,In_2,In_1461);
or U2501 (N_2501,In_275,In_162);
or U2502 (N_2502,In_60,In_845);
or U2503 (N_2503,In_488,In_1333);
or U2504 (N_2504,In_1087,In_701);
nor U2505 (N_2505,In_139,In_815);
nor U2506 (N_2506,In_765,In_811);
and U2507 (N_2507,In_1446,In_1118);
nor U2508 (N_2508,In_1321,In_433);
nor U2509 (N_2509,In_1449,In_1030);
nor U2510 (N_2510,In_799,In_1087);
nand U2511 (N_2511,In_217,In_792);
or U2512 (N_2512,In_1180,In_1003);
nor U2513 (N_2513,In_121,In_783);
nand U2514 (N_2514,In_1258,In_1428);
nand U2515 (N_2515,In_1352,In_169);
nor U2516 (N_2516,In_1205,In_1051);
nor U2517 (N_2517,In_581,In_19);
nand U2518 (N_2518,In_100,In_557);
and U2519 (N_2519,In_423,In_1310);
or U2520 (N_2520,In_1430,In_951);
and U2521 (N_2521,In_861,In_90);
and U2522 (N_2522,In_677,In_1221);
or U2523 (N_2523,In_1441,In_675);
or U2524 (N_2524,In_364,In_1194);
nand U2525 (N_2525,In_777,In_246);
or U2526 (N_2526,In_285,In_329);
nor U2527 (N_2527,In_225,In_1309);
nor U2528 (N_2528,In_913,In_223);
or U2529 (N_2529,In_1311,In_654);
and U2530 (N_2530,In_990,In_1269);
nand U2531 (N_2531,In_285,In_605);
nor U2532 (N_2532,In_815,In_320);
and U2533 (N_2533,In_1088,In_17);
nand U2534 (N_2534,In_1133,In_236);
nor U2535 (N_2535,In_306,In_1152);
nor U2536 (N_2536,In_1128,In_1480);
or U2537 (N_2537,In_115,In_660);
or U2538 (N_2538,In_1209,In_662);
nand U2539 (N_2539,In_1385,In_239);
nand U2540 (N_2540,In_1484,In_772);
nor U2541 (N_2541,In_1367,In_925);
or U2542 (N_2542,In_595,In_1491);
and U2543 (N_2543,In_1484,In_295);
nand U2544 (N_2544,In_1084,In_1392);
nor U2545 (N_2545,In_1411,In_1285);
and U2546 (N_2546,In_1454,In_866);
or U2547 (N_2547,In_427,In_813);
or U2548 (N_2548,In_496,In_1208);
nand U2549 (N_2549,In_1000,In_1499);
or U2550 (N_2550,In_410,In_185);
nor U2551 (N_2551,In_1091,In_202);
or U2552 (N_2552,In_122,In_529);
nor U2553 (N_2553,In_461,In_245);
nand U2554 (N_2554,In_658,In_1282);
and U2555 (N_2555,In_112,In_39);
or U2556 (N_2556,In_1349,In_533);
nand U2557 (N_2557,In_869,In_1153);
nand U2558 (N_2558,In_76,In_971);
or U2559 (N_2559,In_868,In_1231);
or U2560 (N_2560,In_983,In_1394);
nand U2561 (N_2561,In_853,In_714);
and U2562 (N_2562,In_1471,In_885);
nor U2563 (N_2563,In_270,In_1203);
nand U2564 (N_2564,In_841,In_1057);
nand U2565 (N_2565,In_116,In_1016);
nor U2566 (N_2566,In_1218,In_261);
nor U2567 (N_2567,In_1123,In_821);
and U2568 (N_2568,In_999,In_694);
nand U2569 (N_2569,In_78,In_813);
or U2570 (N_2570,In_1279,In_996);
or U2571 (N_2571,In_695,In_781);
and U2572 (N_2572,In_637,In_251);
or U2573 (N_2573,In_472,In_998);
or U2574 (N_2574,In_949,In_1185);
nand U2575 (N_2575,In_1446,In_1101);
and U2576 (N_2576,In_45,In_804);
nand U2577 (N_2577,In_204,In_596);
and U2578 (N_2578,In_818,In_27);
and U2579 (N_2579,In_72,In_26);
nor U2580 (N_2580,In_859,In_1444);
or U2581 (N_2581,In_1343,In_210);
nor U2582 (N_2582,In_773,In_940);
and U2583 (N_2583,In_649,In_237);
or U2584 (N_2584,In_408,In_1304);
and U2585 (N_2585,In_740,In_1289);
nand U2586 (N_2586,In_191,In_205);
and U2587 (N_2587,In_1201,In_442);
and U2588 (N_2588,In_1136,In_365);
or U2589 (N_2589,In_1009,In_648);
nand U2590 (N_2590,In_333,In_1129);
or U2591 (N_2591,In_622,In_1413);
nand U2592 (N_2592,In_1067,In_693);
and U2593 (N_2593,In_1051,In_1086);
or U2594 (N_2594,In_847,In_952);
nor U2595 (N_2595,In_1149,In_818);
nand U2596 (N_2596,In_508,In_880);
or U2597 (N_2597,In_1144,In_41);
or U2598 (N_2598,In_1103,In_854);
nor U2599 (N_2599,In_304,In_877);
nand U2600 (N_2600,In_1129,In_587);
nor U2601 (N_2601,In_873,In_626);
nand U2602 (N_2602,In_1020,In_1227);
nor U2603 (N_2603,In_1170,In_687);
nand U2604 (N_2604,In_130,In_360);
nor U2605 (N_2605,In_510,In_195);
nand U2606 (N_2606,In_30,In_976);
nand U2607 (N_2607,In_1419,In_1256);
nor U2608 (N_2608,In_826,In_294);
or U2609 (N_2609,In_789,In_1313);
nand U2610 (N_2610,In_16,In_1495);
and U2611 (N_2611,In_567,In_1161);
nand U2612 (N_2612,In_881,In_112);
and U2613 (N_2613,In_773,In_701);
and U2614 (N_2614,In_608,In_1157);
and U2615 (N_2615,In_790,In_130);
and U2616 (N_2616,In_489,In_349);
nand U2617 (N_2617,In_806,In_1105);
nand U2618 (N_2618,In_1095,In_68);
nand U2619 (N_2619,In_1202,In_216);
and U2620 (N_2620,In_22,In_964);
nand U2621 (N_2621,In_1480,In_343);
nand U2622 (N_2622,In_506,In_1072);
and U2623 (N_2623,In_396,In_729);
or U2624 (N_2624,In_215,In_273);
nor U2625 (N_2625,In_729,In_51);
nand U2626 (N_2626,In_6,In_519);
and U2627 (N_2627,In_1250,In_363);
nand U2628 (N_2628,In_358,In_529);
nand U2629 (N_2629,In_1105,In_381);
nor U2630 (N_2630,In_1130,In_882);
nand U2631 (N_2631,In_1284,In_854);
and U2632 (N_2632,In_1349,In_761);
and U2633 (N_2633,In_148,In_1205);
and U2634 (N_2634,In_1359,In_743);
and U2635 (N_2635,In_498,In_1068);
nor U2636 (N_2636,In_908,In_659);
and U2637 (N_2637,In_454,In_805);
nor U2638 (N_2638,In_56,In_457);
and U2639 (N_2639,In_1395,In_1085);
xor U2640 (N_2640,In_1129,In_138);
or U2641 (N_2641,In_522,In_1175);
nand U2642 (N_2642,In_1375,In_1441);
and U2643 (N_2643,In_940,In_556);
or U2644 (N_2644,In_857,In_792);
or U2645 (N_2645,In_1477,In_932);
and U2646 (N_2646,In_1387,In_1499);
nor U2647 (N_2647,In_60,In_252);
and U2648 (N_2648,In_780,In_881);
nand U2649 (N_2649,In_1377,In_503);
nor U2650 (N_2650,In_462,In_676);
or U2651 (N_2651,In_29,In_1076);
xnor U2652 (N_2652,In_1384,In_261);
and U2653 (N_2653,In_1247,In_1274);
nor U2654 (N_2654,In_1390,In_542);
and U2655 (N_2655,In_84,In_650);
and U2656 (N_2656,In_310,In_263);
nand U2657 (N_2657,In_356,In_858);
nand U2658 (N_2658,In_1321,In_1119);
nand U2659 (N_2659,In_393,In_1312);
and U2660 (N_2660,In_757,In_727);
nor U2661 (N_2661,In_102,In_1352);
nand U2662 (N_2662,In_1079,In_524);
or U2663 (N_2663,In_989,In_1428);
nor U2664 (N_2664,In_1396,In_605);
nor U2665 (N_2665,In_1189,In_1258);
and U2666 (N_2666,In_172,In_837);
or U2667 (N_2667,In_143,In_80);
nor U2668 (N_2668,In_1181,In_275);
or U2669 (N_2669,In_766,In_132);
nor U2670 (N_2670,In_1450,In_758);
nor U2671 (N_2671,In_1124,In_462);
or U2672 (N_2672,In_599,In_233);
nor U2673 (N_2673,In_582,In_684);
or U2674 (N_2674,In_497,In_220);
or U2675 (N_2675,In_734,In_1002);
xnor U2676 (N_2676,In_167,In_1430);
nor U2677 (N_2677,In_185,In_434);
nand U2678 (N_2678,In_1109,In_530);
or U2679 (N_2679,In_1089,In_217);
or U2680 (N_2680,In_58,In_1313);
or U2681 (N_2681,In_192,In_1341);
nor U2682 (N_2682,In_275,In_1114);
nor U2683 (N_2683,In_1129,In_18);
or U2684 (N_2684,In_741,In_436);
or U2685 (N_2685,In_529,In_260);
nand U2686 (N_2686,In_623,In_682);
or U2687 (N_2687,In_899,In_568);
nor U2688 (N_2688,In_908,In_932);
or U2689 (N_2689,In_530,In_1058);
nor U2690 (N_2690,In_601,In_927);
or U2691 (N_2691,In_630,In_26);
and U2692 (N_2692,In_1130,In_62);
or U2693 (N_2693,In_507,In_310);
and U2694 (N_2694,In_1274,In_1071);
or U2695 (N_2695,In_1140,In_1260);
or U2696 (N_2696,In_269,In_570);
and U2697 (N_2697,In_747,In_119);
or U2698 (N_2698,In_0,In_889);
and U2699 (N_2699,In_728,In_1445);
and U2700 (N_2700,In_357,In_1266);
nand U2701 (N_2701,In_466,In_357);
or U2702 (N_2702,In_836,In_639);
nor U2703 (N_2703,In_372,In_106);
and U2704 (N_2704,In_587,In_86);
and U2705 (N_2705,In_401,In_891);
and U2706 (N_2706,In_1169,In_215);
and U2707 (N_2707,In_1342,In_992);
and U2708 (N_2708,In_261,In_132);
nand U2709 (N_2709,In_1135,In_1035);
nand U2710 (N_2710,In_1255,In_1150);
or U2711 (N_2711,In_285,In_10);
nand U2712 (N_2712,In_1195,In_796);
and U2713 (N_2713,In_1419,In_1026);
nand U2714 (N_2714,In_1286,In_61);
or U2715 (N_2715,In_894,In_854);
nor U2716 (N_2716,In_154,In_162);
or U2717 (N_2717,In_652,In_1063);
nor U2718 (N_2718,In_1401,In_71);
nor U2719 (N_2719,In_1458,In_966);
and U2720 (N_2720,In_498,In_553);
nor U2721 (N_2721,In_1281,In_60);
and U2722 (N_2722,In_314,In_577);
nor U2723 (N_2723,In_1117,In_722);
nand U2724 (N_2724,In_824,In_154);
nor U2725 (N_2725,In_818,In_1122);
and U2726 (N_2726,In_741,In_879);
and U2727 (N_2727,In_804,In_226);
nand U2728 (N_2728,In_600,In_175);
nand U2729 (N_2729,In_591,In_669);
or U2730 (N_2730,In_973,In_804);
and U2731 (N_2731,In_1162,In_362);
and U2732 (N_2732,In_603,In_916);
nor U2733 (N_2733,In_335,In_712);
or U2734 (N_2734,In_898,In_528);
nand U2735 (N_2735,In_960,In_748);
or U2736 (N_2736,In_1358,In_1478);
nand U2737 (N_2737,In_1039,In_777);
nor U2738 (N_2738,In_697,In_1343);
or U2739 (N_2739,In_1232,In_1367);
nand U2740 (N_2740,In_945,In_1443);
and U2741 (N_2741,In_1130,In_1109);
nor U2742 (N_2742,In_1309,In_142);
xor U2743 (N_2743,In_859,In_1445);
nor U2744 (N_2744,In_1248,In_487);
or U2745 (N_2745,In_1049,In_131);
and U2746 (N_2746,In_557,In_823);
nand U2747 (N_2747,In_535,In_1215);
nor U2748 (N_2748,In_1198,In_669);
nor U2749 (N_2749,In_462,In_985);
and U2750 (N_2750,In_1145,In_1098);
nor U2751 (N_2751,In_785,In_566);
or U2752 (N_2752,In_362,In_1432);
nand U2753 (N_2753,In_1237,In_1074);
nor U2754 (N_2754,In_692,In_603);
nand U2755 (N_2755,In_1409,In_84);
or U2756 (N_2756,In_732,In_305);
nor U2757 (N_2757,In_216,In_173);
nand U2758 (N_2758,In_421,In_60);
or U2759 (N_2759,In_886,In_334);
nand U2760 (N_2760,In_1410,In_1275);
and U2761 (N_2761,In_852,In_657);
nand U2762 (N_2762,In_1164,In_349);
nor U2763 (N_2763,In_1425,In_1275);
and U2764 (N_2764,In_1375,In_380);
or U2765 (N_2765,In_988,In_862);
or U2766 (N_2766,In_487,In_850);
or U2767 (N_2767,In_204,In_635);
nand U2768 (N_2768,In_269,In_1185);
nand U2769 (N_2769,In_251,In_1152);
nor U2770 (N_2770,In_791,In_481);
nand U2771 (N_2771,In_91,In_1220);
or U2772 (N_2772,In_394,In_1250);
and U2773 (N_2773,In_166,In_1472);
and U2774 (N_2774,In_785,In_43);
nand U2775 (N_2775,In_441,In_1497);
and U2776 (N_2776,In_807,In_1243);
nand U2777 (N_2777,In_159,In_1419);
nand U2778 (N_2778,In_173,In_564);
and U2779 (N_2779,In_907,In_27);
or U2780 (N_2780,In_977,In_351);
or U2781 (N_2781,In_1299,In_731);
or U2782 (N_2782,In_135,In_952);
nor U2783 (N_2783,In_70,In_985);
or U2784 (N_2784,In_493,In_1299);
or U2785 (N_2785,In_277,In_31);
nor U2786 (N_2786,In_1453,In_569);
or U2787 (N_2787,In_1493,In_1456);
and U2788 (N_2788,In_1138,In_890);
nor U2789 (N_2789,In_1419,In_85);
and U2790 (N_2790,In_72,In_1035);
nor U2791 (N_2791,In_1188,In_1233);
nand U2792 (N_2792,In_1426,In_1043);
and U2793 (N_2793,In_71,In_1027);
or U2794 (N_2794,In_773,In_179);
nor U2795 (N_2795,In_1108,In_951);
and U2796 (N_2796,In_1152,In_1326);
nor U2797 (N_2797,In_829,In_470);
and U2798 (N_2798,In_765,In_426);
nor U2799 (N_2799,In_422,In_729);
nand U2800 (N_2800,In_313,In_1088);
nor U2801 (N_2801,In_25,In_1133);
nor U2802 (N_2802,In_680,In_1122);
nand U2803 (N_2803,In_369,In_252);
nand U2804 (N_2804,In_358,In_959);
nor U2805 (N_2805,In_1248,In_1280);
or U2806 (N_2806,In_1075,In_512);
nor U2807 (N_2807,In_1229,In_1080);
nand U2808 (N_2808,In_1211,In_1145);
and U2809 (N_2809,In_31,In_1400);
nor U2810 (N_2810,In_1155,In_353);
nand U2811 (N_2811,In_124,In_638);
nand U2812 (N_2812,In_1442,In_841);
nor U2813 (N_2813,In_1441,In_777);
or U2814 (N_2814,In_962,In_1065);
nor U2815 (N_2815,In_749,In_1436);
or U2816 (N_2816,In_211,In_18);
nand U2817 (N_2817,In_1275,In_1411);
or U2818 (N_2818,In_215,In_213);
and U2819 (N_2819,In_86,In_743);
nand U2820 (N_2820,In_600,In_630);
or U2821 (N_2821,In_1320,In_674);
or U2822 (N_2822,In_843,In_1115);
nand U2823 (N_2823,In_534,In_407);
and U2824 (N_2824,In_1371,In_109);
nand U2825 (N_2825,In_280,In_1214);
nand U2826 (N_2826,In_233,In_74);
or U2827 (N_2827,In_1385,In_768);
nand U2828 (N_2828,In_562,In_712);
nor U2829 (N_2829,In_355,In_1401);
nor U2830 (N_2830,In_46,In_890);
nor U2831 (N_2831,In_0,In_972);
nor U2832 (N_2832,In_456,In_942);
and U2833 (N_2833,In_140,In_408);
nand U2834 (N_2834,In_1198,In_48);
or U2835 (N_2835,In_821,In_457);
and U2836 (N_2836,In_362,In_1209);
or U2837 (N_2837,In_380,In_961);
or U2838 (N_2838,In_1337,In_1235);
nor U2839 (N_2839,In_24,In_228);
nor U2840 (N_2840,In_527,In_357);
nor U2841 (N_2841,In_1043,In_560);
nand U2842 (N_2842,In_331,In_1189);
or U2843 (N_2843,In_681,In_700);
or U2844 (N_2844,In_158,In_417);
nor U2845 (N_2845,In_1264,In_279);
nand U2846 (N_2846,In_3,In_840);
and U2847 (N_2847,In_429,In_682);
nor U2848 (N_2848,In_703,In_919);
or U2849 (N_2849,In_1232,In_447);
nor U2850 (N_2850,In_1493,In_173);
nand U2851 (N_2851,In_1467,In_1072);
nand U2852 (N_2852,In_820,In_870);
nand U2853 (N_2853,In_990,In_855);
and U2854 (N_2854,In_608,In_1203);
nor U2855 (N_2855,In_173,In_1146);
nor U2856 (N_2856,In_240,In_902);
nor U2857 (N_2857,In_1039,In_1433);
or U2858 (N_2858,In_485,In_333);
nand U2859 (N_2859,In_86,In_6);
xor U2860 (N_2860,In_1391,In_660);
nand U2861 (N_2861,In_1342,In_648);
nand U2862 (N_2862,In_660,In_863);
and U2863 (N_2863,In_902,In_1316);
or U2864 (N_2864,In_289,In_831);
nand U2865 (N_2865,In_875,In_9);
nand U2866 (N_2866,In_1489,In_1402);
and U2867 (N_2867,In_981,In_352);
nand U2868 (N_2868,In_745,In_1334);
nor U2869 (N_2869,In_861,In_1041);
nor U2870 (N_2870,In_699,In_1497);
and U2871 (N_2871,In_1355,In_415);
and U2872 (N_2872,In_1236,In_407);
or U2873 (N_2873,In_215,In_128);
or U2874 (N_2874,In_673,In_569);
or U2875 (N_2875,In_317,In_900);
nand U2876 (N_2876,In_767,In_312);
and U2877 (N_2877,In_451,In_1220);
nand U2878 (N_2878,In_562,In_1021);
nand U2879 (N_2879,In_909,In_1363);
and U2880 (N_2880,In_100,In_1066);
or U2881 (N_2881,In_224,In_1406);
or U2882 (N_2882,In_950,In_1491);
and U2883 (N_2883,In_579,In_970);
nand U2884 (N_2884,In_1003,In_408);
and U2885 (N_2885,In_486,In_463);
nand U2886 (N_2886,In_782,In_1009);
and U2887 (N_2887,In_1347,In_595);
or U2888 (N_2888,In_352,In_108);
nand U2889 (N_2889,In_850,In_417);
or U2890 (N_2890,In_350,In_1269);
or U2891 (N_2891,In_481,In_1125);
and U2892 (N_2892,In_631,In_773);
and U2893 (N_2893,In_1344,In_239);
and U2894 (N_2894,In_1377,In_506);
or U2895 (N_2895,In_720,In_23);
or U2896 (N_2896,In_1206,In_830);
and U2897 (N_2897,In_1446,In_1233);
nor U2898 (N_2898,In_1155,In_1035);
nand U2899 (N_2899,In_1051,In_1123);
or U2900 (N_2900,In_995,In_738);
nand U2901 (N_2901,In_313,In_692);
or U2902 (N_2902,In_1084,In_954);
and U2903 (N_2903,In_955,In_625);
nand U2904 (N_2904,In_778,In_1403);
nand U2905 (N_2905,In_1003,In_1366);
and U2906 (N_2906,In_404,In_338);
and U2907 (N_2907,In_479,In_375);
or U2908 (N_2908,In_1397,In_39);
or U2909 (N_2909,In_907,In_45);
nand U2910 (N_2910,In_162,In_627);
nand U2911 (N_2911,In_1258,In_643);
or U2912 (N_2912,In_11,In_633);
nand U2913 (N_2913,In_988,In_1095);
nor U2914 (N_2914,In_895,In_947);
or U2915 (N_2915,In_1101,In_1160);
nor U2916 (N_2916,In_756,In_625);
nor U2917 (N_2917,In_665,In_967);
nand U2918 (N_2918,In_371,In_1334);
or U2919 (N_2919,In_256,In_103);
and U2920 (N_2920,In_208,In_353);
and U2921 (N_2921,In_687,In_1258);
or U2922 (N_2922,In_583,In_671);
nand U2923 (N_2923,In_112,In_16);
nor U2924 (N_2924,In_695,In_1119);
nand U2925 (N_2925,In_486,In_488);
nor U2926 (N_2926,In_645,In_554);
nor U2927 (N_2927,In_314,In_1398);
or U2928 (N_2928,In_1308,In_1437);
nor U2929 (N_2929,In_883,In_1155);
or U2930 (N_2930,In_443,In_545);
nor U2931 (N_2931,In_317,In_10);
nand U2932 (N_2932,In_577,In_315);
and U2933 (N_2933,In_746,In_277);
nand U2934 (N_2934,In_1039,In_138);
nor U2935 (N_2935,In_1246,In_510);
or U2936 (N_2936,In_625,In_1314);
or U2937 (N_2937,In_1197,In_1496);
nand U2938 (N_2938,In_405,In_1104);
nor U2939 (N_2939,In_505,In_211);
and U2940 (N_2940,In_1441,In_1311);
nand U2941 (N_2941,In_408,In_365);
nand U2942 (N_2942,In_624,In_1269);
and U2943 (N_2943,In_1216,In_738);
and U2944 (N_2944,In_1429,In_885);
or U2945 (N_2945,In_1266,In_278);
nand U2946 (N_2946,In_414,In_832);
nand U2947 (N_2947,In_950,In_558);
nor U2948 (N_2948,In_1055,In_1059);
nand U2949 (N_2949,In_937,In_1006);
nor U2950 (N_2950,In_819,In_1086);
and U2951 (N_2951,In_925,In_222);
or U2952 (N_2952,In_1038,In_1490);
and U2953 (N_2953,In_509,In_1089);
or U2954 (N_2954,In_1024,In_1174);
nand U2955 (N_2955,In_984,In_668);
and U2956 (N_2956,In_578,In_1263);
or U2957 (N_2957,In_65,In_648);
nand U2958 (N_2958,In_383,In_864);
nor U2959 (N_2959,In_1061,In_1184);
or U2960 (N_2960,In_28,In_499);
and U2961 (N_2961,In_9,In_115);
nand U2962 (N_2962,In_1268,In_952);
nand U2963 (N_2963,In_615,In_580);
nor U2964 (N_2964,In_1163,In_1018);
and U2965 (N_2965,In_188,In_284);
or U2966 (N_2966,In_360,In_963);
or U2967 (N_2967,In_1153,In_176);
nand U2968 (N_2968,In_94,In_727);
or U2969 (N_2969,In_1132,In_208);
xnor U2970 (N_2970,In_141,In_1156);
or U2971 (N_2971,In_26,In_1185);
and U2972 (N_2972,In_1181,In_1229);
or U2973 (N_2973,In_1379,In_1310);
nor U2974 (N_2974,In_1336,In_1357);
nand U2975 (N_2975,In_1339,In_581);
and U2976 (N_2976,In_1445,In_961);
or U2977 (N_2977,In_1155,In_6);
nor U2978 (N_2978,In_1252,In_795);
and U2979 (N_2979,In_1121,In_1076);
nand U2980 (N_2980,In_746,In_593);
and U2981 (N_2981,In_551,In_1401);
nand U2982 (N_2982,In_534,In_308);
or U2983 (N_2983,In_1161,In_348);
or U2984 (N_2984,In_1296,In_1430);
nor U2985 (N_2985,In_69,In_186);
or U2986 (N_2986,In_1228,In_685);
or U2987 (N_2987,In_1178,In_1071);
and U2988 (N_2988,In_760,In_1178);
nor U2989 (N_2989,In_1455,In_186);
nand U2990 (N_2990,In_1026,In_286);
and U2991 (N_2991,In_371,In_1230);
or U2992 (N_2992,In_971,In_387);
or U2993 (N_2993,In_931,In_1006);
nor U2994 (N_2994,In_442,In_1238);
nor U2995 (N_2995,In_915,In_1152);
nand U2996 (N_2996,In_1208,In_864);
or U2997 (N_2997,In_113,In_1254);
or U2998 (N_2998,In_1143,In_1076);
and U2999 (N_2999,In_752,In_1120);
nand U3000 (N_3000,In_795,In_1116);
nor U3001 (N_3001,In_1186,In_638);
or U3002 (N_3002,In_707,In_1163);
and U3003 (N_3003,In_1103,In_1297);
and U3004 (N_3004,In_384,In_1447);
or U3005 (N_3005,In_1113,In_1131);
nand U3006 (N_3006,In_1190,In_665);
nand U3007 (N_3007,In_277,In_602);
or U3008 (N_3008,In_1159,In_307);
or U3009 (N_3009,In_1280,In_388);
or U3010 (N_3010,In_124,In_715);
nand U3011 (N_3011,In_619,In_1030);
or U3012 (N_3012,In_312,In_776);
and U3013 (N_3013,In_974,In_900);
and U3014 (N_3014,In_1050,In_333);
and U3015 (N_3015,In_1117,In_43);
and U3016 (N_3016,In_362,In_1324);
and U3017 (N_3017,In_633,In_83);
or U3018 (N_3018,In_1362,In_143);
and U3019 (N_3019,In_797,In_89);
nor U3020 (N_3020,In_420,In_124);
or U3021 (N_3021,In_1306,In_425);
and U3022 (N_3022,In_1404,In_1411);
and U3023 (N_3023,In_1243,In_719);
nor U3024 (N_3024,In_38,In_1112);
or U3025 (N_3025,In_1206,In_718);
or U3026 (N_3026,In_1138,In_618);
or U3027 (N_3027,In_18,In_170);
or U3028 (N_3028,In_1227,In_415);
nor U3029 (N_3029,In_701,In_45);
and U3030 (N_3030,In_251,In_853);
nand U3031 (N_3031,In_773,In_243);
and U3032 (N_3032,In_1165,In_123);
and U3033 (N_3033,In_163,In_344);
nor U3034 (N_3034,In_1142,In_888);
and U3035 (N_3035,In_962,In_1142);
or U3036 (N_3036,In_1345,In_248);
nand U3037 (N_3037,In_894,In_729);
nand U3038 (N_3038,In_750,In_476);
and U3039 (N_3039,In_792,In_1376);
or U3040 (N_3040,In_1261,In_652);
or U3041 (N_3041,In_498,In_1306);
nand U3042 (N_3042,In_372,In_507);
nor U3043 (N_3043,In_998,In_878);
nand U3044 (N_3044,In_217,In_840);
and U3045 (N_3045,In_749,In_800);
or U3046 (N_3046,In_228,In_86);
and U3047 (N_3047,In_619,In_796);
or U3048 (N_3048,In_970,In_585);
xnor U3049 (N_3049,In_1190,In_709);
nand U3050 (N_3050,In_698,In_444);
or U3051 (N_3051,In_1386,In_141);
and U3052 (N_3052,In_887,In_142);
or U3053 (N_3053,In_1074,In_911);
and U3054 (N_3054,In_131,In_1018);
or U3055 (N_3055,In_1085,In_1448);
nor U3056 (N_3056,In_37,In_1440);
nor U3057 (N_3057,In_129,In_762);
nand U3058 (N_3058,In_1345,In_1223);
and U3059 (N_3059,In_718,In_1208);
and U3060 (N_3060,In_670,In_1297);
and U3061 (N_3061,In_271,In_901);
or U3062 (N_3062,In_408,In_1265);
nand U3063 (N_3063,In_549,In_226);
and U3064 (N_3064,In_647,In_662);
nand U3065 (N_3065,In_1182,In_1372);
nor U3066 (N_3066,In_1427,In_1476);
or U3067 (N_3067,In_444,In_918);
or U3068 (N_3068,In_262,In_163);
or U3069 (N_3069,In_1489,In_1443);
or U3070 (N_3070,In_557,In_1015);
nor U3071 (N_3071,In_751,In_632);
nand U3072 (N_3072,In_62,In_564);
or U3073 (N_3073,In_503,In_1084);
or U3074 (N_3074,In_736,In_1118);
nand U3075 (N_3075,In_1492,In_798);
nand U3076 (N_3076,In_1157,In_159);
and U3077 (N_3077,In_793,In_267);
or U3078 (N_3078,In_1267,In_1040);
nor U3079 (N_3079,In_233,In_1470);
or U3080 (N_3080,In_786,In_1338);
nand U3081 (N_3081,In_106,In_454);
nand U3082 (N_3082,In_729,In_89);
nand U3083 (N_3083,In_840,In_20);
nand U3084 (N_3084,In_1402,In_391);
nor U3085 (N_3085,In_606,In_1432);
and U3086 (N_3086,In_782,In_1038);
nor U3087 (N_3087,In_643,In_963);
and U3088 (N_3088,In_26,In_633);
and U3089 (N_3089,In_244,In_423);
and U3090 (N_3090,In_783,In_1352);
and U3091 (N_3091,In_385,In_1066);
nor U3092 (N_3092,In_578,In_885);
nand U3093 (N_3093,In_160,In_322);
nor U3094 (N_3094,In_681,In_740);
nor U3095 (N_3095,In_414,In_737);
and U3096 (N_3096,In_670,In_1155);
and U3097 (N_3097,In_745,In_60);
nand U3098 (N_3098,In_889,In_1255);
or U3099 (N_3099,In_1144,In_203);
nor U3100 (N_3100,In_1043,In_378);
or U3101 (N_3101,In_1315,In_685);
and U3102 (N_3102,In_1469,In_758);
nor U3103 (N_3103,In_804,In_466);
xnor U3104 (N_3104,In_297,In_1047);
nand U3105 (N_3105,In_1125,In_594);
and U3106 (N_3106,In_834,In_394);
xnor U3107 (N_3107,In_1135,In_1193);
nand U3108 (N_3108,In_281,In_844);
nand U3109 (N_3109,In_811,In_647);
or U3110 (N_3110,In_891,In_951);
or U3111 (N_3111,In_1151,In_732);
nand U3112 (N_3112,In_365,In_545);
nand U3113 (N_3113,In_955,In_23);
nor U3114 (N_3114,In_916,In_677);
nor U3115 (N_3115,In_125,In_710);
nand U3116 (N_3116,In_980,In_47);
nand U3117 (N_3117,In_1314,In_1226);
and U3118 (N_3118,In_77,In_519);
nand U3119 (N_3119,In_518,In_504);
and U3120 (N_3120,In_779,In_824);
or U3121 (N_3121,In_840,In_184);
or U3122 (N_3122,In_1305,In_872);
nand U3123 (N_3123,In_1145,In_528);
and U3124 (N_3124,In_5,In_564);
nand U3125 (N_3125,In_617,In_1261);
nor U3126 (N_3126,In_510,In_1487);
and U3127 (N_3127,In_400,In_617);
nor U3128 (N_3128,In_159,In_1394);
nand U3129 (N_3129,In_1487,In_612);
or U3130 (N_3130,In_638,In_1118);
nand U3131 (N_3131,In_741,In_502);
and U3132 (N_3132,In_1292,In_758);
and U3133 (N_3133,In_1044,In_924);
or U3134 (N_3134,In_593,In_1197);
or U3135 (N_3135,In_63,In_624);
nor U3136 (N_3136,In_1045,In_210);
and U3137 (N_3137,In_960,In_1248);
nor U3138 (N_3138,In_1153,In_718);
and U3139 (N_3139,In_1329,In_699);
and U3140 (N_3140,In_658,In_938);
nand U3141 (N_3141,In_431,In_1066);
nor U3142 (N_3142,In_671,In_32);
or U3143 (N_3143,In_1392,In_170);
and U3144 (N_3144,In_623,In_1370);
and U3145 (N_3145,In_363,In_443);
or U3146 (N_3146,In_897,In_406);
or U3147 (N_3147,In_500,In_798);
or U3148 (N_3148,In_1432,In_828);
nor U3149 (N_3149,In_1322,In_580);
and U3150 (N_3150,In_959,In_1314);
nor U3151 (N_3151,In_1255,In_51);
or U3152 (N_3152,In_1425,In_970);
or U3153 (N_3153,In_351,In_1226);
and U3154 (N_3154,In_732,In_1263);
nand U3155 (N_3155,In_272,In_201);
xor U3156 (N_3156,In_15,In_989);
nor U3157 (N_3157,In_608,In_1355);
nand U3158 (N_3158,In_528,In_350);
nor U3159 (N_3159,In_1180,In_476);
and U3160 (N_3160,In_1185,In_334);
or U3161 (N_3161,In_1386,In_875);
or U3162 (N_3162,In_517,In_222);
and U3163 (N_3163,In_53,In_178);
or U3164 (N_3164,In_1137,In_779);
and U3165 (N_3165,In_164,In_742);
nand U3166 (N_3166,In_985,In_690);
nor U3167 (N_3167,In_1208,In_742);
and U3168 (N_3168,In_1094,In_1463);
or U3169 (N_3169,In_565,In_808);
and U3170 (N_3170,In_162,In_1226);
nand U3171 (N_3171,In_519,In_88);
nor U3172 (N_3172,In_912,In_125);
nor U3173 (N_3173,In_75,In_800);
nand U3174 (N_3174,In_860,In_1360);
nand U3175 (N_3175,In_1186,In_546);
nor U3176 (N_3176,In_934,In_636);
nand U3177 (N_3177,In_540,In_866);
or U3178 (N_3178,In_179,In_1371);
nand U3179 (N_3179,In_363,In_105);
nor U3180 (N_3180,In_739,In_1289);
nor U3181 (N_3181,In_1294,In_190);
nand U3182 (N_3182,In_1252,In_1010);
nand U3183 (N_3183,In_979,In_316);
or U3184 (N_3184,In_1334,In_292);
nor U3185 (N_3185,In_352,In_275);
and U3186 (N_3186,In_1399,In_65);
nor U3187 (N_3187,In_494,In_1114);
nor U3188 (N_3188,In_510,In_1200);
and U3189 (N_3189,In_102,In_340);
nand U3190 (N_3190,In_256,In_860);
and U3191 (N_3191,In_390,In_1296);
nand U3192 (N_3192,In_932,In_1121);
and U3193 (N_3193,In_559,In_1480);
or U3194 (N_3194,In_1358,In_1455);
and U3195 (N_3195,In_525,In_1186);
or U3196 (N_3196,In_1075,In_237);
nor U3197 (N_3197,In_698,In_446);
and U3198 (N_3198,In_268,In_244);
nand U3199 (N_3199,In_522,In_612);
and U3200 (N_3200,In_1114,In_1270);
nand U3201 (N_3201,In_561,In_311);
nand U3202 (N_3202,In_94,In_1051);
nand U3203 (N_3203,In_1381,In_395);
nor U3204 (N_3204,In_746,In_577);
and U3205 (N_3205,In_846,In_1456);
nor U3206 (N_3206,In_715,In_450);
nand U3207 (N_3207,In_969,In_898);
and U3208 (N_3208,In_1459,In_254);
xor U3209 (N_3209,In_1456,In_1419);
nor U3210 (N_3210,In_820,In_1167);
nor U3211 (N_3211,In_281,In_714);
or U3212 (N_3212,In_639,In_1096);
and U3213 (N_3213,In_1208,In_682);
and U3214 (N_3214,In_320,In_1474);
and U3215 (N_3215,In_281,In_128);
or U3216 (N_3216,In_142,In_401);
and U3217 (N_3217,In_586,In_490);
nor U3218 (N_3218,In_290,In_518);
nor U3219 (N_3219,In_210,In_107);
or U3220 (N_3220,In_1260,In_426);
nor U3221 (N_3221,In_365,In_1121);
nor U3222 (N_3222,In_862,In_772);
and U3223 (N_3223,In_289,In_633);
nand U3224 (N_3224,In_451,In_479);
nand U3225 (N_3225,In_817,In_0);
or U3226 (N_3226,In_1172,In_563);
or U3227 (N_3227,In_954,In_20);
nor U3228 (N_3228,In_834,In_1019);
nor U3229 (N_3229,In_1313,In_326);
nand U3230 (N_3230,In_1112,In_832);
or U3231 (N_3231,In_421,In_993);
nand U3232 (N_3232,In_648,In_1226);
nand U3233 (N_3233,In_1447,In_419);
nor U3234 (N_3234,In_1260,In_457);
or U3235 (N_3235,In_361,In_1359);
nand U3236 (N_3236,In_1292,In_856);
or U3237 (N_3237,In_311,In_565);
or U3238 (N_3238,In_810,In_593);
nand U3239 (N_3239,In_269,In_387);
nor U3240 (N_3240,In_1413,In_260);
nor U3241 (N_3241,In_1326,In_1281);
or U3242 (N_3242,In_617,In_89);
or U3243 (N_3243,In_17,In_180);
nand U3244 (N_3244,In_798,In_1408);
or U3245 (N_3245,In_1321,In_942);
nor U3246 (N_3246,In_959,In_292);
and U3247 (N_3247,In_159,In_94);
nand U3248 (N_3248,In_1013,In_842);
nor U3249 (N_3249,In_749,In_30);
nand U3250 (N_3250,In_1288,In_1453);
or U3251 (N_3251,In_1263,In_1132);
nand U3252 (N_3252,In_706,In_356);
nor U3253 (N_3253,In_1041,In_190);
and U3254 (N_3254,In_776,In_1396);
or U3255 (N_3255,In_1083,In_524);
nand U3256 (N_3256,In_431,In_323);
and U3257 (N_3257,In_1437,In_1113);
or U3258 (N_3258,In_1125,In_825);
nor U3259 (N_3259,In_740,In_176);
and U3260 (N_3260,In_372,In_1356);
nor U3261 (N_3261,In_1260,In_963);
nor U3262 (N_3262,In_1409,In_1075);
and U3263 (N_3263,In_1136,In_1413);
or U3264 (N_3264,In_1187,In_480);
nor U3265 (N_3265,In_655,In_1337);
nand U3266 (N_3266,In_376,In_918);
and U3267 (N_3267,In_1099,In_901);
and U3268 (N_3268,In_578,In_1398);
nor U3269 (N_3269,In_1359,In_228);
nor U3270 (N_3270,In_1110,In_156);
nand U3271 (N_3271,In_794,In_1280);
nor U3272 (N_3272,In_779,In_482);
and U3273 (N_3273,In_900,In_397);
or U3274 (N_3274,In_1264,In_706);
nor U3275 (N_3275,In_1450,In_781);
or U3276 (N_3276,In_1063,In_839);
or U3277 (N_3277,In_951,In_1300);
and U3278 (N_3278,In_302,In_777);
and U3279 (N_3279,In_665,In_28);
and U3280 (N_3280,In_1039,In_1163);
nand U3281 (N_3281,In_183,In_350);
nor U3282 (N_3282,In_1263,In_747);
and U3283 (N_3283,In_628,In_1289);
and U3284 (N_3284,In_1117,In_681);
and U3285 (N_3285,In_984,In_385);
nor U3286 (N_3286,In_995,In_956);
or U3287 (N_3287,In_343,In_1496);
or U3288 (N_3288,In_371,In_887);
and U3289 (N_3289,In_1460,In_328);
nand U3290 (N_3290,In_662,In_712);
and U3291 (N_3291,In_265,In_1313);
or U3292 (N_3292,In_508,In_66);
nand U3293 (N_3293,In_368,In_421);
nand U3294 (N_3294,In_616,In_761);
or U3295 (N_3295,In_840,In_1498);
or U3296 (N_3296,In_1344,In_1170);
or U3297 (N_3297,In_331,In_570);
or U3298 (N_3298,In_285,In_700);
nor U3299 (N_3299,In_895,In_927);
or U3300 (N_3300,In_518,In_623);
nor U3301 (N_3301,In_773,In_1042);
nand U3302 (N_3302,In_805,In_54);
nor U3303 (N_3303,In_245,In_38);
or U3304 (N_3304,In_1156,In_1435);
and U3305 (N_3305,In_750,In_1475);
or U3306 (N_3306,In_43,In_650);
and U3307 (N_3307,In_250,In_77);
and U3308 (N_3308,In_714,In_721);
nand U3309 (N_3309,In_494,In_334);
or U3310 (N_3310,In_1233,In_932);
and U3311 (N_3311,In_207,In_852);
and U3312 (N_3312,In_1342,In_816);
and U3313 (N_3313,In_864,In_416);
and U3314 (N_3314,In_804,In_306);
and U3315 (N_3315,In_136,In_358);
nand U3316 (N_3316,In_817,In_316);
nor U3317 (N_3317,In_194,In_1205);
and U3318 (N_3318,In_733,In_920);
and U3319 (N_3319,In_1441,In_711);
and U3320 (N_3320,In_1482,In_227);
nor U3321 (N_3321,In_1310,In_1001);
nand U3322 (N_3322,In_959,In_1169);
and U3323 (N_3323,In_1324,In_958);
nand U3324 (N_3324,In_661,In_1202);
nand U3325 (N_3325,In_364,In_854);
and U3326 (N_3326,In_360,In_1464);
nor U3327 (N_3327,In_1471,In_197);
nand U3328 (N_3328,In_1207,In_240);
or U3329 (N_3329,In_1055,In_1217);
or U3330 (N_3330,In_601,In_1154);
nor U3331 (N_3331,In_1475,In_364);
nor U3332 (N_3332,In_644,In_1171);
nor U3333 (N_3333,In_1498,In_1312);
nand U3334 (N_3334,In_652,In_1106);
nand U3335 (N_3335,In_403,In_1269);
and U3336 (N_3336,In_1440,In_1115);
or U3337 (N_3337,In_719,In_247);
or U3338 (N_3338,In_1050,In_1348);
or U3339 (N_3339,In_1435,In_1006);
nor U3340 (N_3340,In_433,In_222);
or U3341 (N_3341,In_386,In_650);
nor U3342 (N_3342,In_714,In_667);
nand U3343 (N_3343,In_942,In_795);
nand U3344 (N_3344,In_1148,In_869);
and U3345 (N_3345,In_860,In_721);
and U3346 (N_3346,In_1383,In_1234);
nand U3347 (N_3347,In_782,In_140);
nor U3348 (N_3348,In_983,In_597);
and U3349 (N_3349,In_1277,In_1016);
or U3350 (N_3350,In_279,In_1222);
nand U3351 (N_3351,In_1485,In_1164);
or U3352 (N_3352,In_1371,In_223);
nand U3353 (N_3353,In_411,In_303);
nor U3354 (N_3354,In_214,In_195);
and U3355 (N_3355,In_338,In_114);
nand U3356 (N_3356,In_48,In_687);
nand U3357 (N_3357,In_84,In_129);
and U3358 (N_3358,In_1265,In_359);
nor U3359 (N_3359,In_4,In_717);
nor U3360 (N_3360,In_1259,In_512);
nand U3361 (N_3361,In_808,In_900);
nor U3362 (N_3362,In_1002,In_888);
nand U3363 (N_3363,In_9,In_799);
and U3364 (N_3364,In_337,In_1357);
or U3365 (N_3365,In_1211,In_316);
nand U3366 (N_3366,In_1343,In_504);
nand U3367 (N_3367,In_860,In_466);
nand U3368 (N_3368,In_55,In_830);
nor U3369 (N_3369,In_305,In_206);
and U3370 (N_3370,In_912,In_1166);
nand U3371 (N_3371,In_1416,In_519);
or U3372 (N_3372,In_28,In_534);
and U3373 (N_3373,In_214,In_1062);
nand U3374 (N_3374,In_1284,In_520);
or U3375 (N_3375,In_1113,In_1041);
nand U3376 (N_3376,In_876,In_1104);
nand U3377 (N_3377,In_155,In_848);
and U3378 (N_3378,In_816,In_35);
and U3379 (N_3379,In_1042,In_323);
nor U3380 (N_3380,In_593,In_666);
nor U3381 (N_3381,In_1152,In_631);
nand U3382 (N_3382,In_358,In_572);
nor U3383 (N_3383,In_1377,In_1217);
nand U3384 (N_3384,In_1283,In_1478);
nand U3385 (N_3385,In_768,In_1031);
or U3386 (N_3386,In_153,In_1274);
and U3387 (N_3387,In_1146,In_595);
or U3388 (N_3388,In_863,In_696);
nor U3389 (N_3389,In_1241,In_249);
nor U3390 (N_3390,In_344,In_971);
nand U3391 (N_3391,In_643,In_1302);
nand U3392 (N_3392,In_339,In_1360);
and U3393 (N_3393,In_968,In_1027);
or U3394 (N_3394,In_1494,In_670);
nor U3395 (N_3395,In_1223,In_1393);
nand U3396 (N_3396,In_4,In_1166);
nand U3397 (N_3397,In_1254,In_358);
and U3398 (N_3398,In_1400,In_507);
or U3399 (N_3399,In_906,In_58);
and U3400 (N_3400,In_778,In_1226);
and U3401 (N_3401,In_109,In_604);
nor U3402 (N_3402,In_513,In_504);
and U3403 (N_3403,In_1049,In_822);
and U3404 (N_3404,In_357,In_92);
nor U3405 (N_3405,In_1121,In_96);
or U3406 (N_3406,In_765,In_865);
nor U3407 (N_3407,In_954,In_1059);
and U3408 (N_3408,In_961,In_1332);
and U3409 (N_3409,In_874,In_355);
and U3410 (N_3410,In_481,In_1197);
and U3411 (N_3411,In_1128,In_1014);
and U3412 (N_3412,In_1235,In_769);
and U3413 (N_3413,In_1364,In_1472);
or U3414 (N_3414,In_1147,In_59);
or U3415 (N_3415,In_700,In_552);
nor U3416 (N_3416,In_654,In_1170);
and U3417 (N_3417,In_148,In_421);
nand U3418 (N_3418,In_331,In_1207);
nand U3419 (N_3419,In_1050,In_205);
or U3420 (N_3420,In_638,In_1496);
or U3421 (N_3421,In_933,In_78);
or U3422 (N_3422,In_854,In_428);
xor U3423 (N_3423,In_956,In_942);
nand U3424 (N_3424,In_372,In_1432);
nor U3425 (N_3425,In_1349,In_767);
or U3426 (N_3426,In_737,In_1152);
nor U3427 (N_3427,In_748,In_1244);
nand U3428 (N_3428,In_721,In_1245);
or U3429 (N_3429,In_986,In_149);
or U3430 (N_3430,In_722,In_746);
nand U3431 (N_3431,In_1366,In_248);
nand U3432 (N_3432,In_655,In_952);
and U3433 (N_3433,In_275,In_875);
and U3434 (N_3434,In_1283,In_836);
and U3435 (N_3435,In_66,In_1397);
or U3436 (N_3436,In_517,In_698);
or U3437 (N_3437,In_958,In_869);
nor U3438 (N_3438,In_1070,In_1005);
or U3439 (N_3439,In_528,In_395);
nand U3440 (N_3440,In_484,In_328);
nor U3441 (N_3441,In_1301,In_1339);
or U3442 (N_3442,In_396,In_1295);
nor U3443 (N_3443,In_1224,In_55);
and U3444 (N_3444,In_1338,In_667);
nand U3445 (N_3445,In_658,In_1436);
nor U3446 (N_3446,In_1066,In_3);
and U3447 (N_3447,In_499,In_80);
or U3448 (N_3448,In_1256,In_484);
nor U3449 (N_3449,In_1124,In_345);
nand U3450 (N_3450,In_365,In_317);
and U3451 (N_3451,In_478,In_416);
nor U3452 (N_3452,In_957,In_829);
and U3453 (N_3453,In_390,In_1002);
or U3454 (N_3454,In_1479,In_1248);
nor U3455 (N_3455,In_615,In_465);
and U3456 (N_3456,In_1111,In_1172);
nor U3457 (N_3457,In_547,In_798);
and U3458 (N_3458,In_942,In_199);
or U3459 (N_3459,In_691,In_257);
and U3460 (N_3460,In_980,In_158);
nand U3461 (N_3461,In_935,In_1093);
nand U3462 (N_3462,In_488,In_120);
or U3463 (N_3463,In_1406,In_99);
and U3464 (N_3464,In_1330,In_1120);
and U3465 (N_3465,In_1251,In_431);
and U3466 (N_3466,In_1052,In_426);
and U3467 (N_3467,In_58,In_1489);
nor U3468 (N_3468,In_256,In_725);
nor U3469 (N_3469,In_1448,In_207);
nand U3470 (N_3470,In_342,In_332);
or U3471 (N_3471,In_1095,In_104);
or U3472 (N_3472,In_1232,In_1192);
nor U3473 (N_3473,In_545,In_716);
nor U3474 (N_3474,In_1321,In_444);
and U3475 (N_3475,In_1269,In_1261);
or U3476 (N_3476,In_1467,In_903);
and U3477 (N_3477,In_515,In_1385);
nand U3478 (N_3478,In_1245,In_5);
and U3479 (N_3479,In_102,In_934);
and U3480 (N_3480,In_705,In_686);
nand U3481 (N_3481,In_129,In_256);
nand U3482 (N_3482,In_1226,In_793);
nor U3483 (N_3483,In_242,In_163);
nand U3484 (N_3484,In_701,In_1225);
nand U3485 (N_3485,In_1107,In_1030);
or U3486 (N_3486,In_1017,In_1229);
and U3487 (N_3487,In_801,In_1009);
and U3488 (N_3488,In_674,In_1488);
nor U3489 (N_3489,In_1377,In_779);
or U3490 (N_3490,In_1084,In_897);
nor U3491 (N_3491,In_907,In_1471);
nand U3492 (N_3492,In_879,In_598);
nor U3493 (N_3493,In_126,In_1201);
nand U3494 (N_3494,In_807,In_328);
nor U3495 (N_3495,In_327,In_1066);
nand U3496 (N_3496,In_53,In_857);
nand U3497 (N_3497,In_114,In_321);
and U3498 (N_3498,In_120,In_1099);
and U3499 (N_3499,In_1150,In_207);
nand U3500 (N_3500,In_1119,In_558);
and U3501 (N_3501,In_120,In_96);
or U3502 (N_3502,In_930,In_1173);
or U3503 (N_3503,In_1174,In_632);
nor U3504 (N_3504,In_1305,In_610);
nand U3505 (N_3505,In_952,In_1313);
or U3506 (N_3506,In_1155,In_543);
nor U3507 (N_3507,In_1407,In_336);
or U3508 (N_3508,In_381,In_661);
nor U3509 (N_3509,In_1021,In_107);
or U3510 (N_3510,In_359,In_1147);
nand U3511 (N_3511,In_441,In_814);
and U3512 (N_3512,In_1139,In_1400);
and U3513 (N_3513,In_463,In_223);
and U3514 (N_3514,In_104,In_31);
or U3515 (N_3515,In_586,In_1322);
and U3516 (N_3516,In_78,In_1131);
and U3517 (N_3517,In_1257,In_362);
nand U3518 (N_3518,In_87,In_493);
nor U3519 (N_3519,In_987,In_1224);
or U3520 (N_3520,In_1167,In_211);
nor U3521 (N_3521,In_1134,In_951);
nor U3522 (N_3522,In_879,In_1433);
and U3523 (N_3523,In_823,In_1354);
and U3524 (N_3524,In_650,In_76);
nand U3525 (N_3525,In_1172,In_108);
or U3526 (N_3526,In_687,In_1279);
nand U3527 (N_3527,In_76,In_20);
or U3528 (N_3528,In_787,In_215);
or U3529 (N_3529,In_93,In_617);
and U3530 (N_3530,In_245,In_1129);
and U3531 (N_3531,In_643,In_21);
nand U3532 (N_3532,In_601,In_1450);
nand U3533 (N_3533,In_421,In_1338);
or U3534 (N_3534,In_817,In_714);
or U3535 (N_3535,In_198,In_241);
or U3536 (N_3536,In_472,In_362);
nor U3537 (N_3537,In_1458,In_809);
nand U3538 (N_3538,In_1390,In_1250);
or U3539 (N_3539,In_1491,In_775);
nor U3540 (N_3540,In_266,In_302);
nand U3541 (N_3541,In_954,In_848);
and U3542 (N_3542,In_1112,In_525);
nor U3543 (N_3543,In_43,In_1494);
nand U3544 (N_3544,In_920,In_1097);
and U3545 (N_3545,In_960,In_421);
or U3546 (N_3546,In_699,In_726);
nor U3547 (N_3547,In_1077,In_1426);
or U3548 (N_3548,In_166,In_911);
or U3549 (N_3549,In_300,In_122);
and U3550 (N_3550,In_840,In_222);
nand U3551 (N_3551,In_406,In_454);
and U3552 (N_3552,In_240,In_1223);
and U3553 (N_3553,In_442,In_781);
nor U3554 (N_3554,In_845,In_701);
nor U3555 (N_3555,In_151,In_165);
nand U3556 (N_3556,In_447,In_535);
or U3557 (N_3557,In_1261,In_1309);
nor U3558 (N_3558,In_217,In_356);
or U3559 (N_3559,In_877,In_1382);
nand U3560 (N_3560,In_940,In_587);
and U3561 (N_3561,In_356,In_960);
nand U3562 (N_3562,In_235,In_56);
nor U3563 (N_3563,In_1204,In_694);
and U3564 (N_3564,In_593,In_1148);
or U3565 (N_3565,In_842,In_847);
and U3566 (N_3566,In_547,In_223);
nand U3567 (N_3567,In_419,In_18);
and U3568 (N_3568,In_821,In_315);
or U3569 (N_3569,In_1211,In_398);
or U3570 (N_3570,In_1349,In_1158);
nand U3571 (N_3571,In_394,In_1455);
nand U3572 (N_3572,In_12,In_65);
nand U3573 (N_3573,In_912,In_697);
nand U3574 (N_3574,In_1190,In_624);
and U3575 (N_3575,In_1270,In_33);
nand U3576 (N_3576,In_632,In_817);
or U3577 (N_3577,In_1075,In_298);
nand U3578 (N_3578,In_1331,In_327);
and U3579 (N_3579,In_967,In_1131);
nand U3580 (N_3580,In_1065,In_899);
nor U3581 (N_3581,In_615,In_1379);
nor U3582 (N_3582,In_1446,In_47);
and U3583 (N_3583,In_79,In_356);
and U3584 (N_3584,In_125,In_1318);
nand U3585 (N_3585,In_427,In_128);
nand U3586 (N_3586,In_0,In_1386);
nand U3587 (N_3587,In_455,In_1435);
and U3588 (N_3588,In_687,In_108);
nand U3589 (N_3589,In_1191,In_1142);
and U3590 (N_3590,In_107,In_626);
or U3591 (N_3591,In_1257,In_1135);
nand U3592 (N_3592,In_812,In_1398);
or U3593 (N_3593,In_592,In_676);
and U3594 (N_3594,In_1095,In_476);
nand U3595 (N_3595,In_439,In_84);
nand U3596 (N_3596,In_609,In_81);
nor U3597 (N_3597,In_541,In_831);
and U3598 (N_3598,In_36,In_1373);
nand U3599 (N_3599,In_250,In_936);
and U3600 (N_3600,In_123,In_135);
nand U3601 (N_3601,In_217,In_1269);
and U3602 (N_3602,In_297,In_1323);
nand U3603 (N_3603,In_734,In_1153);
and U3604 (N_3604,In_163,In_1198);
and U3605 (N_3605,In_68,In_422);
or U3606 (N_3606,In_545,In_240);
nor U3607 (N_3607,In_1304,In_694);
or U3608 (N_3608,In_824,In_1449);
or U3609 (N_3609,In_186,In_183);
or U3610 (N_3610,In_534,In_803);
nor U3611 (N_3611,In_1073,In_105);
and U3612 (N_3612,In_1327,In_903);
nand U3613 (N_3613,In_1256,In_955);
and U3614 (N_3614,In_713,In_925);
and U3615 (N_3615,In_389,In_870);
nand U3616 (N_3616,In_172,In_1392);
nor U3617 (N_3617,In_115,In_401);
nand U3618 (N_3618,In_219,In_223);
nand U3619 (N_3619,In_1030,In_624);
or U3620 (N_3620,In_1254,In_724);
or U3621 (N_3621,In_1270,In_854);
or U3622 (N_3622,In_20,In_1448);
or U3623 (N_3623,In_761,In_756);
nor U3624 (N_3624,In_1009,In_415);
nand U3625 (N_3625,In_803,In_1423);
nor U3626 (N_3626,In_1433,In_456);
or U3627 (N_3627,In_166,In_988);
nor U3628 (N_3628,In_445,In_358);
nor U3629 (N_3629,In_530,In_369);
and U3630 (N_3630,In_1146,In_51);
nor U3631 (N_3631,In_1045,In_894);
and U3632 (N_3632,In_1497,In_1451);
or U3633 (N_3633,In_1046,In_202);
or U3634 (N_3634,In_974,In_788);
or U3635 (N_3635,In_245,In_971);
nand U3636 (N_3636,In_1094,In_805);
nor U3637 (N_3637,In_1496,In_397);
or U3638 (N_3638,In_1387,In_159);
nand U3639 (N_3639,In_594,In_914);
nand U3640 (N_3640,In_571,In_747);
or U3641 (N_3641,In_476,In_32);
or U3642 (N_3642,In_755,In_1465);
nand U3643 (N_3643,In_1116,In_90);
nand U3644 (N_3644,In_958,In_210);
or U3645 (N_3645,In_538,In_74);
and U3646 (N_3646,In_1036,In_211);
or U3647 (N_3647,In_56,In_1180);
and U3648 (N_3648,In_26,In_1356);
nor U3649 (N_3649,In_462,In_330);
or U3650 (N_3650,In_1202,In_1219);
or U3651 (N_3651,In_1203,In_338);
nor U3652 (N_3652,In_856,In_1049);
or U3653 (N_3653,In_422,In_14);
and U3654 (N_3654,In_1250,In_470);
or U3655 (N_3655,In_499,In_711);
and U3656 (N_3656,In_1301,In_1026);
and U3657 (N_3657,In_153,In_1158);
nor U3658 (N_3658,In_1271,In_930);
and U3659 (N_3659,In_290,In_198);
or U3660 (N_3660,In_1354,In_534);
or U3661 (N_3661,In_1361,In_1092);
or U3662 (N_3662,In_912,In_1345);
and U3663 (N_3663,In_1231,In_331);
nor U3664 (N_3664,In_615,In_343);
or U3665 (N_3665,In_386,In_173);
and U3666 (N_3666,In_527,In_1111);
nand U3667 (N_3667,In_52,In_499);
or U3668 (N_3668,In_9,In_496);
or U3669 (N_3669,In_65,In_681);
or U3670 (N_3670,In_1006,In_154);
nor U3671 (N_3671,In_1358,In_1263);
nor U3672 (N_3672,In_568,In_1427);
xor U3673 (N_3673,In_1280,In_760);
and U3674 (N_3674,In_330,In_1349);
nor U3675 (N_3675,In_651,In_158);
nor U3676 (N_3676,In_1279,In_1356);
nand U3677 (N_3677,In_658,In_1038);
nand U3678 (N_3678,In_995,In_1422);
and U3679 (N_3679,In_120,In_702);
or U3680 (N_3680,In_566,In_276);
nand U3681 (N_3681,In_1126,In_558);
and U3682 (N_3682,In_941,In_732);
nor U3683 (N_3683,In_798,In_313);
nor U3684 (N_3684,In_207,In_393);
and U3685 (N_3685,In_1027,In_366);
or U3686 (N_3686,In_207,In_1261);
and U3687 (N_3687,In_1193,In_1439);
or U3688 (N_3688,In_1276,In_559);
nand U3689 (N_3689,In_1073,In_1372);
nor U3690 (N_3690,In_446,In_546);
or U3691 (N_3691,In_564,In_1283);
or U3692 (N_3692,In_187,In_1122);
and U3693 (N_3693,In_1230,In_935);
or U3694 (N_3694,In_785,In_375);
nor U3695 (N_3695,In_214,In_623);
nor U3696 (N_3696,In_1438,In_818);
or U3697 (N_3697,In_906,In_365);
nand U3698 (N_3698,In_642,In_321);
and U3699 (N_3699,In_768,In_534);
or U3700 (N_3700,In_1426,In_1256);
and U3701 (N_3701,In_1253,In_824);
nand U3702 (N_3702,In_961,In_726);
nor U3703 (N_3703,In_1102,In_413);
nand U3704 (N_3704,In_745,In_280);
nor U3705 (N_3705,In_10,In_1193);
and U3706 (N_3706,In_1383,In_4);
nor U3707 (N_3707,In_430,In_664);
and U3708 (N_3708,In_372,In_702);
and U3709 (N_3709,In_292,In_635);
nor U3710 (N_3710,In_1166,In_881);
and U3711 (N_3711,In_1349,In_759);
nand U3712 (N_3712,In_72,In_1274);
and U3713 (N_3713,In_353,In_574);
nor U3714 (N_3714,In_1216,In_36);
and U3715 (N_3715,In_683,In_429);
nand U3716 (N_3716,In_860,In_338);
and U3717 (N_3717,In_594,In_995);
nand U3718 (N_3718,In_792,In_132);
and U3719 (N_3719,In_550,In_556);
or U3720 (N_3720,In_456,In_1377);
nand U3721 (N_3721,In_146,In_90);
or U3722 (N_3722,In_1105,In_154);
or U3723 (N_3723,In_518,In_302);
nand U3724 (N_3724,In_1368,In_464);
and U3725 (N_3725,In_749,In_74);
and U3726 (N_3726,In_1441,In_864);
nor U3727 (N_3727,In_107,In_247);
or U3728 (N_3728,In_432,In_325);
or U3729 (N_3729,In_1179,In_1226);
nand U3730 (N_3730,In_870,In_254);
or U3731 (N_3731,In_1487,In_735);
and U3732 (N_3732,In_664,In_1222);
nand U3733 (N_3733,In_505,In_636);
and U3734 (N_3734,In_942,In_1227);
nor U3735 (N_3735,In_368,In_246);
and U3736 (N_3736,In_993,In_741);
nor U3737 (N_3737,In_851,In_12);
and U3738 (N_3738,In_355,In_6);
nand U3739 (N_3739,In_892,In_1117);
nor U3740 (N_3740,In_843,In_701);
nand U3741 (N_3741,In_773,In_1044);
nor U3742 (N_3742,In_1088,In_1377);
and U3743 (N_3743,In_1375,In_754);
nor U3744 (N_3744,In_815,In_146);
nor U3745 (N_3745,In_1179,In_1467);
and U3746 (N_3746,In_1423,In_125);
nor U3747 (N_3747,In_1167,In_234);
or U3748 (N_3748,In_1264,In_719);
nor U3749 (N_3749,In_1153,In_1237);
or U3750 (N_3750,In_6,In_1136);
nand U3751 (N_3751,In_55,In_1253);
nor U3752 (N_3752,In_1078,In_1168);
or U3753 (N_3753,In_442,In_1339);
and U3754 (N_3754,In_853,In_484);
nand U3755 (N_3755,In_910,In_1447);
nand U3756 (N_3756,In_69,In_1287);
nand U3757 (N_3757,In_850,In_1344);
and U3758 (N_3758,In_162,In_927);
and U3759 (N_3759,In_707,In_536);
or U3760 (N_3760,In_487,In_1364);
nor U3761 (N_3761,In_470,In_1367);
nor U3762 (N_3762,In_1078,In_1421);
nor U3763 (N_3763,In_437,In_1038);
or U3764 (N_3764,In_410,In_588);
nand U3765 (N_3765,In_861,In_1388);
nand U3766 (N_3766,In_46,In_1198);
nor U3767 (N_3767,In_337,In_1389);
nand U3768 (N_3768,In_390,In_584);
nand U3769 (N_3769,In_235,In_607);
and U3770 (N_3770,In_1496,In_172);
or U3771 (N_3771,In_870,In_1112);
and U3772 (N_3772,In_228,In_745);
nor U3773 (N_3773,In_395,In_1183);
nand U3774 (N_3774,In_1315,In_1051);
nor U3775 (N_3775,In_464,In_687);
nand U3776 (N_3776,In_1054,In_1024);
nand U3777 (N_3777,In_69,In_662);
and U3778 (N_3778,In_87,In_134);
and U3779 (N_3779,In_723,In_1307);
nand U3780 (N_3780,In_869,In_64);
nand U3781 (N_3781,In_90,In_826);
and U3782 (N_3782,In_1345,In_1340);
or U3783 (N_3783,In_306,In_50);
nor U3784 (N_3784,In_220,In_1386);
nand U3785 (N_3785,In_1498,In_831);
nand U3786 (N_3786,In_1408,In_1326);
or U3787 (N_3787,In_1453,In_522);
or U3788 (N_3788,In_1391,In_230);
and U3789 (N_3789,In_942,In_392);
or U3790 (N_3790,In_750,In_218);
or U3791 (N_3791,In_1219,In_718);
or U3792 (N_3792,In_915,In_1066);
and U3793 (N_3793,In_915,In_716);
nor U3794 (N_3794,In_1457,In_558);
xor U3795 (N_3795,In_1307,In_573);
or U3796 (N_3796,In_491,In_835);
and U3797 (N_3797,In_1153,In_529);
nor U3798 (N_3798,In_414,In_162);
nand U3799 (N_3799,In_1476,In_783);
and U3800 (N_3800,In_842,In_210);
and U3801 (N_3801,In_934,In_467);
nand U3802 (N_3802,In_815,In_423);
and U3803 (N_3803,In_9,In_862);
nor U3804 (N_3804,In_849,In_382);
and U3805 (N_3805,In_891,In_503);
or U3806 (N_3806,In_710,In_1132);
or U3807 (N_3807,In_1466,In_283);
nor U3808 (N_3808,In_362,In_1418);
nand U3809 (N_3809,In_427,In_686);
and U3810 (N_3810,In_266,In_695);
nor U3811 (N_3811,In_106,In_470);
and U3812 (N_3812,In_1436,In_787);
and U3813 (N_3813,In_713,In_1482);
nor U3814 (N_3814,In_1214,In_449);
nand U3815 (N_3815,In_56,In_1090);
or U3816 (N_3816,In_397,In_257);
nor U3817 (N_3817,In_605,In_234);
nand U3818 (N_3818,In_1117,In_470);
nand U3819 (N_3819,In_1476,In_133);
and U3820 (N_3820,In_1237,In_445);
nand U3821 (N_3821,In_131,In_1426);
or U3822 (N_3822,In_957,In_936);
nand U3823 (N_3823,In_455,In_20);
or U3824 (N_3824,In_967,In_461);
nor U3825 (N_3825,In_4,In_1340);
nor U3826 (N_3826,In_983,In_1181);
nor U3827 (N_3827,In_532,In_342);
and U3828 (N_3828,In_107,In_823);
nand U3829 (N_3829,In_192,In_30);
xnor U3830 (N_3830,In_795,In_740);
and U3831 (N_3831,In_447,In_1193);
and U3832 (N_3832,In_1333,In_521);
and U3833 (N_3833,In_1352,In_12);
or U3834 (N_3834,In_428,In_557);
nand U3835 (N_3835,In_285,In_1020);
and U3836 (N_3836,In_1499,In_1406);
or U3837 (N_3837,In_33,In_233);
and U3838 (N_3838,In_1317,In_613);
and U3839 (N_3839,In_1267,In_1303);
or U3840 (N_3840,In_204,In_745);
and U3841 (N_3841,In_1003,In_707);
or U3842 (N_3842,In_281,In_191);
nand U3843 (N_3843,In_922,In_498);
nand U3844 (N_3844,In_807,In_81);
nor U3845 (N_3845,In_313,In_280);
and U3846 (N_3846,In_244,In_1186);
nor U3847 (N_3847,In_226,In_501);
or U3848 (N_3848,In_699,In_115);
nand U3849 (N_3849,In_321,In_644);
and U3850 (N_3850,In_604,In_529);
nor U3851 (N_3851,In_452,In_474);
nor U3852 (N_3852,In_347,In_1269);
nand U3853 (N_3853,In_751,In_1333);
nand U3854 (N_3854,In_1316,In_854);
nand U3855 (N_3855,In_905,In_89);
and U3856 (N_3856,In_238,In_138);
nor U3857 (N_3857,In_312,In_994);
nand U3858 (N_3858,In_88,In_762);
nor U3859 (N_3859,In_832,In_507);
nor U3860 (N_3860,In_775,In_1307);
and U3861 (N_3861,In_430,In_242);
nor U3862 (N_3862,In_452,In_509);
and U3863 (N_3863,In_1047,In_843);
nor U3864 (N_3864,In_1158,In_1489);
nor U3865 (N_3865,In_107,In_739);
nand U3866 (N_3866,In_488,In_738);
nor U3867 (N_3867,In_650,In_571);
nand U3868 (N_3868,In_284,In_1190);
nand U3869 (N_3869,In_229,In_672);
or U3870 (N_3870,In_689,In_568);
xor U3871 (N_3871,In_369,In_1036);
or U3872 (N_3872,In_918,In_533);
nor U3873 (N_3873,In_1322,In_1082);
nand U3874 (N_3874,In_465,In_419);
nor U3875 (N_3875,In_134,In_1446);
nand U3876 (N_3876,In_1255,In_184);
nand U3877 (N_3877,In_1041,In_632);
and U3878 (N_3878,In_847,In_170);
nand U3879 (N_3879,In_152,In_1446);
nor U3880 (N_3880,In_114,In_761);
or U3881 (N_3881,In_445,In_252);
or U3882 (N_3882,In_88,In_287);
nand U3883 (N_3883,In_260,In_632);
and U3884 (N_3884,In_223,In_1321);
and U3885 (N_3885,In_659,In_1158);
and U3886 (N_3886,In_400,In_664);
nand U3887 (N_3887,In_1097,In_222);
nand U3888 (N_3888,In_1097,In_1168);
and U3889 (N_3889,In_920,In_19);
or U3890 (N_3890,In_171,In_289);
nand U3891 (N_3891,In_1092,In_435);
nand U3892 (N_3892,In_1090,In_517);
nor U3893 (N_3893,In_533,In_814);
and U3894 (N_3894,In_702,In_171);
nor U3895 (N_3895,In_549,In_1319);
nor U3896 (N_3896,In_41,In_951);
nor U3897 (N_3897,In_354,In_1375);
nand U3898 (N_3898,In_1310,In_10);
nor U3899 (N_3899,In_494,In_488);
nand U3900 (N_3900,In_215,In_1065);
nand U3901 (N_3901,In_611,In_705);
and U3902 (N_3902,In_75,In_359);
nand U3903 (N_3903,In_457,In_777);
nand U3904 (N_3904,In_706,In_1184);
or U3905 (N_3905,In_1212,In_15);
or U3906 (N_3906,In_69,In_804);
or U3907 (N_3907,In_1056,In_1011);
and U3908 (N_3908,In_8,In_446);
nor U3909 (N_3909,In_362,In_1229);
nor U3910 (N_3910,In_1300,In_263);
or U3911 (N_3911,In_1206,In_418);
nor U3912 (N_3912,In_1109,In_731);
or U3913 (N_3913,In_961,In_1322);
and U3914 (N_3914,In_1497,In_797);
nand U3915 (N_3915,In_357,In_975);
or U3916 (N_3916,In_842,In_548);
xnor U3917 (N_3917,In_90,In_1003);
nor U3918 (N_3918,In_1404,In_395);
or U3919 (N_3919,In_804,In_1432);
nor U3920 (N_3920,In_1102,In_200);
nand U3921 (N_3921,In_552,In_207);
or U3922 (N_3922,In_446,In_425);
and U3923 (N_3923,In_1403,In_1315);
nand U3924 (N_3924,In_386,In_709);
or U3925 (N_3925,In_97,In_671);
or U3926 (N_3926,In_1338,In_1242);
and U3927 (N_3927,In_1414,In_946);
nor U3928 (N_3928,In_801,In_863);
or U3929 (N_3929,In_192,In_128);
nor U3930 (N_3930,In_955,In_475);
nand U3931 (N_3931,In_870,In_950);
and U3932 (N_3932,In_1102,In_1058);
nand U3933 (N_3933,In_880,In_631);
nand U3934 (N_3934,In_978,In_796);
or U3935 (N_3935,In_1283,In_521);
and U3936 (N_3936,In_638,In_281);
nor U3937 (N_3937,In_346,In_258);
and U3938 (N_3938,In_643,In_521);
and U3939 (N_3939,In_1058,In_234);
or U3940 (N_3940,In_672,In_135);
and U3941 (N_3941,In_1072,In_1058);
and U3942 (N_3942,In_1114,In_1079);
nand U3943 (N_3943,In_500,In_680);
or U3944 (N_3944,In_833,In_957);
nor U3945 (N_3945,In_1324,In_1425);
nand U3946 (N_3946,In_658,In_1300);
and U3947 (N_3947,In_1354,In_959);
nand U3948 (N_3948,In_1421,In_963);
nand U3949 (N_3949,In_51,In_898);
and U3950 (N_3950,In_773,In_540);
or U3951 (N_3951,In_1310,In_1222);
nor U3952 (N_3952,In_1136,In_61);
or U3953 (N_3953,In_809,In_274);
nand U3954 (N_3954,In_9,In_15);
nor U3955 (N_3955,In_64,In_573);
nand U3956 (N_3956,In_1051,In_645);
and U3957 (N_3957,In_441,In_1331);
and U3958 (N_3958,In_327,In_128);
nor U3959 (N_3959,In_808,In_254);
and U3960 (N_3960,In_275,In_513);
or U3961 (N_3961,In_1338,In_346);
nor U3962 (N_3962,In_1270,In_1101);
nor U3963 (N_3963,In_1428,In_885);
nor U3964 (N_3964,In_204,In_1215);
nor U3965 (N_3965,In_676,In_1175);
nor U3966 (N_3966,In_773,In_320);
nor U3967 (N_3967,In_1157,In_812);
nor U3968 (N_3968,In_651,In_494);
nor U3969 (N_3969,In_419,In_219);
nand U3970 (N_3970,In_993,In_967);
nor U3971 (N_3971,In_1312,In_1303);
and U3972 (N_3972,In_1074,In_518);
nand U3973 (N_3973,In_200,In_1490);
nand U3974 (N_3974,In_1267,In_1389);
and U3975 (N_3975,In_863,In_1231);
nand U3976 (N_3976,In_1071,In_763);
nor U3977 (N_3977,In_819,In_303);
or U3978 (N_3978,In_572,In_1354);
or U3979 (N_3979,In_817,In_1399);
or U3980 (N_3980,In_487,In_402);
nand U3981 (N_3981,In_542,In_1141);
and U3982 (N_3982,In_1069,In_234);
and U3983 (N_3983,In_1266,In_1291);
nand U3984 (N_3984,In_1229,In_682);
nand U3985 (N_3985,In_1323,In_661);
nor U3986 (N_3986,In_701,In_22);
nand U3987 (N_3987,In_1036,In_1091);
or U3988 (N_3988,In_1102,In_1374);
nor U3989 (N_3989,In_152,In_191);
or U3990 (N_3990,In_249,In_331);
nor U3991 (N_3991,In_875,In_662);
or U3992 (N_3992,In_1050,In_160);
nor U3993 (N_3993,In_1485,In_784);
and U3994 (N_3994,In_929,In_1119);
and U3995 (N_3995,In_1395,In_628);
nand U3996 (N_3996,In_1278,In_82);
nor U3997 (N_3997,In_396,In_69);
nor U3998 (N_3998,In_447,In_400);
and U3999 (N_3999,In_792,In_168);
and U4000 (N_4000,In_941,In_1220);
nor U4001 (N_4001,In_698,In_301);
nand U4002 (N_4002,In_197,In_1247);
and U4003 (N_4003,In_16,In_1432);
nor U4004 (N_4004,In_895,In_675);
nand U4005 (N_4005,In_879,In_570);
and U4006 (N_4006,In_722,In_527);
nand U4007 (N_4007,In_403,In_385);
nor U4008 (N_4008,In_879,In_198);
and U4009 (N_4009,In_1162,In_1452);
and U4010 (N_4010,In_639,In_473);
and U4011 (N_4011,In_1128,In_876);
and U4012 (N_4012,In_395,In_986);
nor U4013 (N_4013,In_1073,In_506);
nor U4014 (N_4014,In_84,In_1199);
and U4015 (N_4015,In_1464,In_479);
or U4016 (N_4016,In_995,In_985);
nor U4017 (N_4017,In_661,In_780);
nand U4018 (N_4018,In_620,In_1311);
nor U4019 (N_4019,In_459,In_324);
nor U4020 (N_4020,In_1000,In_268);
and U4021 (N_4021,In_896,In_1316);
or U4022 (N_4022,In_671,In_679);
and U4023 (N_4023,In_254,In_1159);
and U4024 (N_4024,In_122,In_804);
nand U4025 (N_4025,In_1413,In_151);
or U4026 (N_4026,In_1080,In_520);
and U4027 (N_4027,In_1078,In_603);
and U4028 (N_4028,In_1301,In_817);
nor U4029 (N_4029,In_1478,In_446);
nor U4030 (N_4030,In_484,In_965);
and U4031 (N_4031,In_845,In_938);
nor U4032 (N_4032,In_751,In_626);
nand U4033 (N_4033,In_1167,In_923);
nand U4034 (N_4034,In_16,In_262);
or U4035 (N_4035,In_1296,In_558);
nand U4036 (N_4036,In_1320,In_804);
nor U4037 (N_4037,In_277,In_145);
or U4038 (N_4038,In_1493,In_799);
or U4039 (N_4039,In_349,In_595);
or U4040 (N_4040,In_1315,In_488);
and U4041 (N_4041,In_91,In_1422);
or U4042 (N_4042,In_1061,In_140);
nand U4043 (N_4043,In_204,In_979);
and U4044 (N_4044,In_944,In_61);
nor U4045 (N_4045,In_36,In_107);
nand U4046 (N_4046,In_97,In_261);
and U4047 (N_4047,In_324,In_958);
nand U4048 (N_4048,In_880,In_928);
nand U4049 (N_4049,In_504,In_1342);
and U4050 (N_4050,In_508,In_1064);
or U4051 (N_4051,In_1003,In_886);
nor U4052 (N_4052,In_391,In_1196);
and U4053 (N_4053,In_1085,In_164);
or U4054 (N_4054,In_1311,In_659);
or U4055 (N_4055,In_1252,In_1003);
nor U4056 (N_4056,In_570,In_328);
nand U4057 (N_4057,In_304,In_1223);
or U4058 (N_4058,In_988,In_618);
nor U4059 (N_4059,In_457,In_89);
or U4060 (N_4060,In_1153,In_1171);
nor U4061 (N_4061,In_1488,In_1067);
nor U4062 (N_4062,In_327,In_1127);
or U4063 (N_4063,In_811,In_518);
or U4064 (N_4064,In_354,In_502);
nand U4065 (N_4065,In_1275,In_503);
nor U4066 (N_4066,In_1490,In_738);
or U4067 (N_4067,In_62,In_271);
or U4068 (N_4068,In_1191,In_910);
or U4069 (N_4069,In_663,In_387);
or U4070 (N_4070,In_438,In_112);
and U4071 (N_4071,In_1009,In_331);
or U4072 (N_4072,In_1443,In_242);
or U4073 (N_4073,In_121,In_985);
or U4074 (N_4074,In_331,In_413);
nand U4075 (N_4075,In_1116,In_161);
xor U4076 (N_4076,In_1436,In_536);
nor U4077 (N_4077,In_344,In_748);
nand U4078 (N_4078,In_483,In_163);
and U4079 (N_4079,In_233,In_731);
or U4080 (N_4080,In_96,In_241);
and U4081 (N_4081,In_611,In_485);
and U4082 (N_4082,In_839,In_1108);
and U4083 (N_4083,In_630,In_801);
and U4084 (N_4084,In_131,In_893);
or U4085 (N_4085,In_1219,In_1390);
and U4086 (N_4086,In_1278,In_954);
nand U4087 (N_4087,In_20,In_821);
nand U4088 (N_4088,In_1046,In_491);
nor U4089 (N_4089,In_1058,In_1089);
nor U4090 (N_4090,In_581,In_994);
or U4091 (N_4091,In_1410,In_612);
nor U4092 (N_4092,In_1017,In_472);
and U4093 (N_4093,In_92,In_1463);
and U4094 (N_4094,In_1417,In_691);
nand U4095 (N_4095,In_528,In_388);
or U4096 (N_4096,In_654,In_1079);
nor U4097 (N_4097,In_75,In_1142);
nor U4098 (N_4098,In_189,In_383);
or U4099 (N_4099,In_565,In_349);
and U4100 (N_4100,In_964,In_526);
nor U4101 (N_4101,In_95,In_935);
nand U4102 (N_4102,In_169,In_1078);
nand U4103 (N_4103,In_1218,In_796);
or U4104 (N_4104,In_428,In_317);
nor U4105 (N_4105,In_1009,In_1372);
nor U4106 (N_4106,In_793,In_1051);
nand U4107 (N_4107,In_132,In_1051);
and U4108 (N_4108,In_937,In_413);
and U4109 (N_4109,In_750,In_509);
and U4110 (N_4110,In_79,In_1199);
and U4111 (N_4111,In_1319,In_956);
or U4112 (N_4112,In_1435,In_726);
nand U4113 (N_4113,In_1483,In_373);
and U4114 (N_4114,In_1049,In_979);
nor U4115 (N_4115,In_525,In_219);
nor U4116 (N_4116,In_363,In_652);
or U4117 (N_4117,In_189,In_1223);
nor U4118 (N_4118,In_115,In_219);
and U4119 (N_4119,In_1049,In_197);
nand U4120 (N_4120,In_1008,In_711);
nor U4121 (N_4121,In_1497,In_940);
and U4122 (N_4122,In_67,In_1083);
and U4123 (N_4123,In_1341,In_882);
and U4124 (N_4124,In_746,In_859);
and U4125 (N_4125,In_695,In_568);
and U4126 (N_4126,In_681,In_314);
nor U4127 (N_4127,In_729,In_49);
nor U4128 (N_4128,In_741,In_470);
or U4129 (N_4129,In_1321,In_410);
and U4130 (N_4130,In_74,In_920);
nand U4131 (N_4131,In_520,In_1495);
nor U4132 (N_4132,In_1255,In_329);
and U4133 (N_4133,In_411,In_910);
nand U4134 (N_4134,In_541,In_623);
nor U4135 (N_4135,In_745,In_1228);
or U4136 (N_4136,In_78,In_916);
and U4137 (N_4137,In_726,In_14);
nor U4138 (N_4138,In_138,In_659);
or U4139 (N_4139,In_1338,In_492);
nor U4140 (N_4140,In_519,In_1398);
and U4141 (N_4141,In_811,In_1494);
or U4142 (N_4142,In_1313,In_649);
nor U4143 (N_4143,In_93,In_224);
or U4144 (N_4144,In_1482,In_434);
and U4145 (N_4145,In_27,In_1024);
nor U4146 (N_4146,In_1123,In_1088);
nor U4147 (N_4147,In_786,In_206);
and U4148 (N_4148,In_1404,In_806);
nand U4149 (N_4149,In_1352,In_305);
or U4150 (N_4150,In_364,In_938);
nor U4151 (N_4151,In_237,In_457);
or U4152 (N_4152,In_1355,In_771);
nand U4153 (N_4153,In_764,In_981);
or U4154 (N_4154,In_1413,In_638);
nand U4155 (N_4155,In_1146,In_1414);
or U4156 (N_4156,In_1420,In_1157);
and U4157 (N_4157,In_314,In_1480);
nand U4158 (N_4158,In_1395,In_1367);
or U4159 (N_4159,In_781,In_232);
and U4160 (N_4160,In_325,In_873);
and U4161 (N_4161,In_1211,In_289);
and U4162 (N_4162,In_144,In_171);
nor U4163 (N_4163,In_607,In_732);
and U4164 (N_4164,In_795,In_727);
and U4165 (N_4165,In_993,In_159);
or U4166 (N_4166,In_686,In_230);
and U4167 (N_4167,In_1218,In_845);
or U4168 (N_4168,In_588,In_675);
nand U4169 (N_4169,In_1332,In_1019);
and U4170 (N_4170,In_1123,In_163);
nor U4171 (N_4171,In_1102,In_1479);
and U4172 (N_4172,In_281,In_114);
and U4173 (N_4173,In_46,In_586);
nand U4174 (N_4174,In_1453,In_1167);
or U4175 (N_4175,In_1475,In_831);
nor U4176 (N_4176,In_942,In_1216);
and U4177 (N_4177,In_828,In_292);
nand U4178 (N_4178,In_1315,In_31);
and U4179 (N_4179,In_1405,In_759);
or U4180 (N_4180,In_660,In_1497);
nand U4181 (N_4181,In_1372,In_621);
or U4182 (N_4182,In_233,In_401);
nor U4183 (N_4183,In_647,In_705);
and U4184 (N_4184,In_330,In_22);
and U4185 (N_4185,In_290,In_1087);
nor U4186 (N_4186,In_1292,In_63);
xnor U4187 (N_4187,In_1181,In_242);
nor U4188 (N_4188,In_875,In_777);
nor U4189 (N_4189,In_547,In_420);
and U4190 (N_4190,In_68,In_1430);
and U4191 (N_4191,In_425,In_691);
nor U4192 (N_4192,In_606,In_744);
and U4193 (N_4193,In_1007,In_488);
and U4194 (N_4194,In_589,In_396);
and U4195 (N_4195,In_522,In_424);
nor U4196 (N_4196,In_449,In_1265);
and U4197 (N_4197,In_771,In_473);
nor U4198 (N_4198,In_1167,In_1112);
or U4199 (N_4199,In_1439,In_60);
nand U4200 (N_4200,In_1067,In_1367);
nand U4201 (N_4201,In_832,In_742);
and U4202 (N_4202,In_1284,In_631);
and U4203 (N_4203,In_1436,In_1408);
nand U4204 (N_4204,In_1417,In_752);
or U4205 (N_4205,In_597,In_120);
nand U4206 (N_4206,In_640,In_988);
nand U4207 (N_4207,In_1256,In_1339);
or U4208 (N_4208,In_884,In_336);
or U4209 (N_4209,In_1226,In_602);
or U4210 (N_4210,In_1284,In_709);
xnor U4211 (N_4211,In_452,In_1118);
or U4212 (N_4212,In_627,In_921);
or U4213 (N_4213,In_15,In_821);
nand U4214 (N_4214,In_1343,In_1026);
nor U4215 (N_4215,In_195,In_88);
and U4216 (N_4216,In_853,In_70);
nand U4217 (N_4217,In_855,In_1460);
nand U4218 (N_4218,In_196,In_1206);
nor U4219 (N_4219,In_1118,In_5);
nor U4220 (N_4220,In_945,In_1444);
nor U4221 (N_4221,In_382,In_54);
nand U4222 (N_4222,In_54,In_185);
and U4223 (N_4223,In_922,In_100);
xnor U4224 (N_4224,In_632,In_292);
and U4225 (N_4225,In_725,In_528);
and U4226 (N_4226,In_1343,In_620);
or U4227 (N_4227,In_1066,In_446);
nand U4228 (N_4228,In_513,In_1479);
or U4229 (N_4229,In_747,In_1270);
nor U4230 (N_4230,In_1344,In_802);
or U4231 (N_4231,In_612,In_1032);
nor U4232 (N_4232,In_1110,In_16);
or U4233 (N_4233,In_979,In_1190);
and U4234 (N_4234,In_27,In_1403);
nand U4235 (N_4235,In_454,In_1423);
and U4236 (N_4236,In_9,In_1111);
and U4237 (N_4237,In_402,In_326);
nor U4238 (N_4238,In_1281,In_951);
nor U4239 (N_4239,In_1058,In_1356);
nor U4240 (N_4240,In_737,In_1175);
or U4241 (N_4241,In_1,In_666);
nor U4242 (N_4242,In_834,In_824);
nand U4243 (N_4243,In_606,In_966);
nand U4244 (N_4244,In_327,In_393);
and U4245 (N_4245,In_653,In_25);
or U4246 (N_4246,In_975,In_1338);
and U4247 (N_4247,In_1449,In_1117);
nand U4248 (N_4248,In_127,In_605);
nand U4249 (N_4249,In_1202,In_1334);
or U4250 (N_4250,In_64,In_1295);
nor U4251 (N_4251,In_1009,In_539);
and U4252 (N_4252,In_1077,In_1091);
nand U4253 (N_4253,In_1081,In_670);
or U4254 (N_4254,In_1491,In_485);
nand U4255 (N_4255,In_1491,In_138);
nor U4256 (N_4256,In_1333,In_1222);
or U4257 (N_4257,In_821,In_517);
and U4258 (N_4258,In_55,In_1073);
nor U4259 (N_4259,In_940,In_1201);
and U4260 (N_4260,In_1240,In_355);
nand U4261 (N_4261,In_194,In_388);
and U4262 (N_4262,In_761,In_1170);
xor U4263 (N_4263,In_1108,In_614);
nor U4264 (N_4264,In_964,In_1211);
and U4265 (N_4265,In_1100,In_257);
or U4266 (N_4266,In_1188,In_406);
or U4267 (N_4267,In_274,In_1277);
nor U4268 (N_4268,In_502,In_1431);
and U4269 (N_4269,In_1301,In_628);
nand U4270 (N_4270,In_258,In_1102);
or U4271 (N_4271,In_241,In_745);
or U4272 (N_4272,In_1219,In_143);
nor U4273 (N_4273,In_8,In_181);
or U4274 (N_4274,In_436,In_1465);
nand U4275 (N_4275,In_956,In_630);
or U4276 (N_4276,In_669,In_893);
nor U4277 (N_4277,In_360,In_1495);
nor U4278 (N_4278,In_374,In_265);
or U4279 (N_4279,In_803,In_796);
nor U4280 (N_4280,In_1153,In_36);
or U4281 (N_4281,In_316,In_479);
and U4282 (N_4282,In_454,In_1026);
and U4283 (N_4283,In_1231,In_506);
or U4284 (N_4284,In_324,In_1311);
or U4285 (N_4285,In_1213,In_848);
or U4286 (N_4286,In_931,In_1155);
or U4287 (N_4287,In_1028,In_947);
or U4288 (N_4288,In_270,In_830);
nand U4289 (N_4289,In_458,In_1376);
nor U4290 (N_4290,In_250,In_136);
or U4291 (N_4291,In_57,In_76);
nand U4292 (N_4292,In_305,In_1169);
or U4293 (N_4293,In_1429,In_1165);
nand U4294 (N_4294,In_711,In_1241);
or U4295 (N_4295,In_1210,In_1009);
or U4296 (N_4296,In_1391,In_1100);
nor U4297 (N_4297,In_1271,In_981);
xor U4298 (N_4298,In_579,In_1251);
nor U4299 (N_4299,In_537,In_581);
nand U4300 (N_4300,In_940,In_1435);
nand U4301 (N_4301,In_1050,In_1480);
and U4302 (N_4302,In_736,In_1366);
nor U4303 (N_4303,In_1382,In_1467);
nor U4304 (N_4304,In_1136,In_289);
or U4305 (N_4305,In_554,In_301);
and U4306 (N_4306,In_525,In_1366);
or U4307 (N_4307,In_1352,In_257);
or U4308 (N_4308,In_1189,In_865);
or U4309 (N_4309,In_514,In_630);
and U4310 (N_4310,In_1125,In_615);
or U4311 (N_4311,In_587,In_245);
nand U4312 (N_4312,In_720,In_584);
nor U4313 (N_4313,In_663,In_304);
and U4314 (N_4314,In_431,In_570);
nor U4315 (N_4315,In_93,In_493);
or U4316 (N_4316,In_1368,In_857);
nand U4317 (N_4317,In_1448,In_413);
nor U4318 (N_4318,In_1049,In_1184);
and U4319 (N_4319,In_1299,In_631);
nor U4320 (N_4320,In_835,In_276);
and U4321 (N_4321,In_15,In_388);
nor U4322 (N_4322,In_10,In_93);
or U4323 (N_4323,In_1037,In_778);
nand U4324 (N_4324,In_172,In_1038);
nand U4325 (N_4325,In_483,In_351);
or U4326 (N_4326,In_98,In_1017);
nand U4327 (N_4327,In_42,In_1196);
or U4328 (N_4328,In_935,In_319);
or U4329 (N_4329,In_723,In_375);
nor U4330 (N_4330,In_100,In_1373);
and U4331 (N_4331,In_1037,In_1335);
nor U4332 (N_4332,In_1440,In_434);
nand U4333 (N_4333,In_1151,In_1258);
or U4334 (N_4334,In_95,In_1308);
nand U4335 (N_4335,In_506,In_139);
nand U4336 (N_4336,In_364,In_128);
nand U4337 (N_4337,In_90,In_1129);
and U4338 (N_4338,In_1318,In_151);
nor U4339 (N_4339,In_473,In_490);
and U4340 (N_4340,In_888,In_403);
nor U4341 (N_4341,In_1127,In_1282);
nor U4342 (N_4342,In_456,In_1211);
or U4343 (N_4343,In_59,In_1053);
or U4344 (N_4344,In_472,In_707);
and U4345 (N_4345,In_1337,In_1319);
nand U4346 (N_4346,In_458,In_76);
and U4347 (N_4347,In_815,In_873);
and U4348 (N_4348,In_569,In_19);
or U4349 (N_4349,In_1061,In_561);
nor U4350 (N_4350,In_137,In_307);
and U4351 (N_4351,In_438,In_576);
and U4352 (N_4352,In_991,In_164);
or U4353 (N_4353,In_868,In_968);
or U4354 (N_4354,In_499,In_1405);
nor U4355 (N_4355,In_817,In_1409);
and U4356 (N_4356,In_905,In_23);
or U4357 (N_4357,In_957,In_1158);
or U4358 (N_4358,In_488,In_927);
and U4359 (N_4359,In_1117,In_922);
and U4360 (N_4360,In_155,In_356);
nor U4361 (N_4361,In_400,In_557);
nand U4362 (N_4362,In_1114,In_731);
nor U4363 (N_4363,In_194,In_1166);
nor U4364 (N_4364,In_636,In_427);
nor U4365 (N_4365,In_810,In_1430);
or U4366 (N_4366,In_1224,In_1371);
nor U4367 (N_4367,In_940,In_1366);
or U4368 (N_4368,In_1427,In_498);
and U4369 (N_4369,In_1150,In_1287);
nand U4370 (N_4370,In_390,In_292);
nand U4371 (N_4371,In_237,In_314);
and U4372 (N_4372,In_314,In_1060);
nand U4373 (N_4373,In_1337,In_669);
or U4374 (N_4374,In_991,In_265);
nand U4375 (N_4375,In_706,In_1283);
or U4376 (N_4376,In_173,In_174);
nor U4377 (N_4377,In_1282,In_1042);
and U4378 (N_4378,In_582,In_186);
and U4379 (N_4379,In_323,In_1225);
or U4380 (N_4380,In_1102,In_12);
or U4381 (N_4381,In_1109,In_1127);
and U4382 (N_4382,In_153,In_1050);
or U4383 (N_4383,In_264,In_356);
or U4384 (N_4384,In_379,In_1161);
nor U4385 (N_4385,In_368,In_1460);
nand U4386 (N_4386,In_225,In_157);
nand U4387 (N_4387,In_367,In_822);
nor U4388 (N_4388,In_51,In_510);
nor U4389 (N_4389,In_1238,In_634);
nor U4390 (N_4390,In_1053,In_1199);
or U4391 (N_4391,In_49,In_575);
nor U4392 (N_4392,In_337,In_401);
xor U4393 (N_4393,In_8,In_1288);
nand U4394 (N_4394,In_1496,In_1114);
nor U4395 (N_4395,In_151,In_1007);
nand U4396 (N_4396,In_518,In_115);
nor U4397 (N_4397,In_1140,In_1089);
or U4398 (N_4398,In_294,In_1250);
or U4399 (N_4399,In_261,In_1199);
or U4400 (N_4400,In_1205,In_1050);
nor U4401 (N_4401,In_1072,In_1217);
nor U4402 (N_4402,In_1058,In_155);
or U4403 (N_4403,In_341,In_868);
nor U4404 (N_4404,In_837,In_415);
and U4405 (N_4405,In_175,In_856);
nor U4406 (N_4406,In_954,In_1095);
nor U4407 (N_4407,In_18,In_543);
and U4408 (N_4408,In_1432,In_423);
nor U4409 (N_4409,In_804,In_1431);
nor U4410 (N_4410,In_341,In_982);
nand U4411 (N_4411,In_1279,In_641);
and U4412 (N_4412,In_1148,In_356);
nor U4413 (N_4413,In_1007,In_1438);
or U4414 (N_4414,In_174,In_493);
and U4415 (N_4415,In_735,In_704);
and U4416 (N_4416,In_647,In_1241);
or U4417 (N_4417,In_1328,In_305);
and U4418 (N_4418,In_1,In_1258);
nand U4419 (N_4419,In_265,In_1141);
or U4420 (N_4420,In_657,In_93);
nand U4421 (N_4421,In_358,In_365);
and U4422 (N_4422,In_753,In_60);
nand U4423 (N_4423,In_1144,In_1028);
or U4424 (N_4424,In_192,In_223);
nor U4425 (N_4425,In_1351,In_134);
or U4426 (N_4426,In_22,In_241);
or U4427 (N_4427,In_738,In_485);
nand U4428 (N_4428,In_410,In_433);
nand U4429 (N_4429,In_851,In_1298);
or U4430 (N_4430,In_766,In_1035);
or U4431 (N_4431,In_1393,In_291);
nor U4432 (N_4432,In_1232,In_903);
nand U4433 (N_4433,In_398,In_430);
or U4434 (N_4434,In_702,In_833);
nor U4435 (N_4435,In_633,In_734);
and U4436 (N_4436,In_579,In_860);
nand U4437 (N_4437,In_322,In_152);
nand U4438 (N_4438,In_163,In_657);
nand U4439 (N_4439,In_67,In_882);
and U4440 (N_4440,In_793,In_1206);
nand U4441 (N_4441,In_309,In_111);
nand U4442 (N_4442,In_190,In_253);
or U4443 (N_4443,In_1202,In_890);
nand U4444 (N_4444,In_1258,In_50);
nor U4445 (N_4445,In_149,In_185);
or U4446 (N_4446,In_705,In_453);
or U4447 (N_4447,In_525,In_577);
nor U4448 (N_4448,In_219,In_1135);
and U4449 (N_4449,In_362,In_750);
and U4450 (N_4450,In_512,In_501);
nor U4451 (N_4451,In_487,In_1047);
or U4452 (N_4452,In_553,In_478);
or U4453 (N_4453,In_1392,In_611);
nor U4454 (N_4454,In_33,In_428);
nand U4455 (N_4455,In_365,In_51);
or U4456 (N_4456,In_613,In_625);
nand U4457 (N_4457,In_1136,In_825);
nand U4458 (N_4458,In_953,In_942);
and U4459 (N_4459,In_1048,In_333);
or U4460 (N_4460,In_1005,In_960);
or U4461 (N_4461,In_691,In_1086);
xor U4462 (N_4462,In_617,In_297);
or U4463 (N_4463,In_511,In_558);
or U4464 (N_4464,In_600,In_945);
nand U4465 (N_4465,In_300,In_1205);
and U4466 (N_4466,In_982,In_277);
nor U4467 (N_4467,In_1286,In_581);
or U4468 (N_4468,In_784,In_417);
or U4469 (N_4469,In_921,In_886);
and U4470 (N_4470,In_837,In_514);
nor U4471 (N_4471,In_1300,In_1025);
nand U4472 (N_4472,In_1188,In_1377);
nand U4473 (N_4473,In_238,In_1458);
nand U4474 (N_4474,In_965,In_156);
or U4475 (N_4475,In_1406,In_227);
and U4476 (N_4476,In_406,In_474);
and U4477 (N_4477,In_59,In_389);
nor U4478 (N_4478,In_239,In_555);
and U4479 (N_4479,In_1006,In_1135);
and U4480 (N_4480,In_1054,In_851);
and U4481 (N_4481,In_1331,In_1137);
and U4482 (N_4482,In_797,In_477);
nand U4483 (N_4483,In_1104,In_639);
or U4484 (N_4484,In_1250,In_1305);
and U4485 (N_4485,In_896,In_723);
nor U4486 (N_4486,In_1279,In_1482);
and U4487 (N_4487,In_404,In_700);
nand U4488 (N_4488,In_832,In_63);
nand U4489 (N_4489,In_12,In_1475);
and U4490 (N_4490,In_229,In_317);
nand U4491 (N_4491,In_842,In_239);
and U4492 (N_4492,In_994,In_562);
nor U4493 (N_4493,In_367,In_1306);
nor U4494 (N_4494,In_1284,In_1274);
and U4495 (N_4495,In_1468,In_86);
and U4496 (N_4496,In_1228,In_929);
nand U4497 (N_4497,In_324,In_1177);
nand U4498 (N_4498,In_269,In_215);
xor U4499 (N_4499,In_830,In_439);
or U4500 (N_4500,In_538,In_375);
or U4501 (N_4501,In_901,In_1241);
nor U4502 (N_4502,In_951,In_443);
nor U4503 (N_4503,In_673,In_1056);
and U4504 (N_4504,In_1203,In_1152);
and U4505 (N_4505,In_1021,In_1346);
nor U4506 (N_4506,In_399,In_463);
nor U4507 (N_4507,In_311,In_793);
nor U4508 (N_4508,In_325,In_634);
and U4509 (N_4509,In_679,In_760);
nand U4510 (N_4510,In_941,In_1157);
or U4511 (N_4511,In_705,In_783);
nor U4512 (N_4512,In_11,In_1295);
or U4513 (N_4513,In_539,In_401);
nand U4514 (N_4514,In_477,In_509);
nand U4515 (N_4515,In_1327,In_255);
nand U4516 (N_4516,In_870,In_1292);
nand U4517 (N_4517,In_945,In_994);
nor U4518 (N_4518,In_703,In_48);
and U4519 (N_4519,In_972,In_584);
nor U4520 (N_4520,In_1040,In_664);
or U4521 (N_4521,In_1083,In_988);
nand U4522 (N_4522,In_78,In_637);
and U4523 (N_4523,In_1171,In_26);
and U4524 (N_4524,In_1314,In_1359);
or U4525 (N_4525,In_1300,In_1469);
and U4526 (N_4526,In_4,In_89);
nor U4527 (N_4527,In_1422,In_967);
nor U4528 (N_4528,In_461,In_677);
and U4529 (N_4529,In_166,In_1381);
and U4530 (N_4530,In_362,In_291);
or U4531 (N_4531,In_1130,In_713);
and U4532 (N_4532,In_76,In_149);
nand U4533 (N_4533,In_790,In_1284);
nand U4534 (N_4534,In_878,In_917);
nor U4535 (N_4535,In_282,In_224);
nor U4536 (N_4536,In_1269,In_183);
nand U4537 (N_4537,In_66,In_972);
and U4538 (N_4538,In_483,In_1463);
or U4539 (N_4539,In_530,In_190);
nor U4540 (N_4540,In_13,In_1228);
and U4541 (N_4541,In_1198,In_1272);
nor U4542 (N_4542,In_1100,In_634);
nor U4543 (N_4543,In_619,In_1291);
nand U4544 (N_4544,In_768,In_1452);
or U4545 (N_4545,In_173,In_612);
nor U4546 (N_4546,In_760,In_1005);
or U4547 (N_4547,In_889,In_1412);
and U4548 (N_4548,In_1269,In_1447);
nor U4549 (N_4549,In_494,In_296);
and U4550 (N_4550,In_881,In_1041);
nor U4551 (N_4551,In_116,In_553);
and U4552 (N_4552,In_485,In_1320);
nand U4553 (N_4553,In_193,In_1419);
nand U4554 (N_4554,In_560,In_74);
nand U4555 (N_4555,In_1450,In_515);
nand U4556 (N_4556,In_136,In_691);
nand U4557 (N_4557,In_629,In_289);
nor U4558 (N_4558,In_190,In_930);
nor U4559 (N_4559,In_759,In_881);
and U4560 (N_4560,In_1415,In_1368);
nand U4561 (N_4561,In_9,In_765);
and U4562 (N_4562,In_487,In_618);
and U4563 (N_4563,In_1054,In_1390);
and U4564 (N_4564,In_478,In_343);
nor U4565 (N_4565,In_1130,In_487);
nand U4566 (N_4566,In_694,In_1224);
and U4567 (N_4567,In_1119,In_921);
nor U4568 (N_4568,In_1303,In_598);
or U4569 (N_4569,In_885,In_1451);
nor U4570 (N_4570,In_140,In_874);
or U4571 (N_4571,In_1036,In_107);
and U4572 (N_4572,In_1384,In_500);
nand U4573 (N_4573,In_920,In_1296);
or U4574 (N_4574,In_983,In_1399);
nor U4575 (N_4575,In_269,In_1106);
or U4576 (N_4576,In_904,In_1263);
nor U4577 (N_4577,In_803,In_1052);
nor U4578 (N_4578,In_730,In_1187);
nand U4579 (N_4579,In_476,In_695);
and U4580 (N_4580,In_296,In_174);
nor U4581 (N_4581,In_176,In_1461);
or U4582 (N_4582,In_704,In_1356);
and U4583 (N_4583,In_40,In_1239);
or U4584 (N_4584,In_344,In_28);
nor U4585 (N_4585,In_1256,In_1075);
and U4586 (N_4586,In_976,In_71);
nand U4587 (N_4587,In_881,In_955);
nand U4588 (N_4588,In_1139,In_274);
nand U4589 (N_4589,In_194,In_1126);
nor U4590 (N_4590,In_621,In_1333);
nand U4591 (N_4591,In_746,In_299);
and U4592 (N_4592,In_1445,In_1325);
nand U4593 (N_4593,In_426,In_592);
or U4594 (N_4594,In_321,In_524);
or U4595 (N_4595,In_651,In_611);
xnor U4596 (N_4596,In_1452,In_1094);
and U4597 (N_4597,In_1306,In_353);
or U4598 (N_4598,In_700,In_497);
or U4599 (N_4599,In_755,In_1235);
nand U4600 (N_4600,In_649,In_1422);
and U4601 (N_4601,In_369,In_704);
and U4602 (N_4602,In_132,In_735);
nand U4603 (N_4603,In_531,In_917);
or U4604 (N_4604,In_1209,In_160);
nand U4605 (N_4605,In_291,In_336);
nor U4606 (N_4606,In_361,In_295);
and U4607 (N_4607,In_1429,In_879);
or U4608 (N_4608,In_940,In_7);
nand U4609 (N_4609,In_273,In_263);
nand U4610 (N_4610,In_594,In_358);
nor U4611 (N_4611,In_850,In_1205);
nor U4612 (N_4612,In_4,In_1480);
and U4613 (N_4613,In_52,In_1063);
nor U4614 (N_4614,In_363,In_1484);
nand U4615 (N_4615,In_1189,In_653);
nor U4616 (N_4616,In_1462,In_573);
xor U4617 (N_4617,In_527,In_234);
or U4618 (N_4618,In_244,In_1397);
nand U4619 (N_4619,In_190,In_13);
nand U4620 (N_4620,In_458,In_44);
and U4621 (N_4621,In_441,In_1241);
and U4622 (N_4622,In_43,In_993);
and U4623 (N_4623,In_603,In_140);
and U4624 (N_4624,In_1238,In_1035);
and U4625 (N_4625,In_544,In_671);
xnor U4626 (N_4626,In_637,In_1326);
or U4627 (N_4627,In_700,In_435);
nand U4628 (N_4628,In_90,In_832);
or U4629 (N_4629,In_1049,In_791);
nor U4630 (N_4630,In_949,In_428);
nand U4631 (N_4631,In_599,In_444);
nand U4632 (N_4632,In_538,In_1003);
and U4633 (N_4633,In_847,In_388);
or U4634 (N_4634,In_322,In_1280);
nand U4635 (N_4635,In_255,In_1082);
nand U4636 (N_4636,In_950,In_280);
nor U4637 (N_4637,In_495,In_772);
nand U4638 (N_4638,In_1024,In_759);
nor U4639 (N_4639,In_26,In_114);
nand U4640 (N_4640,In_243,In_1223);
or U4641 (N_4641,In_508,In_734);
or U4642 (N_4642,In_233,In_1192);
nand U4643 (N_4643,In_910,In_924);
and U4644 (N_4644,In_465,In_1017);
nor U4645 (N_4645,In_373,In_1298);
nand U4646 (N_4646,In_314,In_986);
nand U4647 (N_4647,In_706,In_778);
or U4648 (N_4648,In_318,In_838);
nand U4649 (N_4649,In_675,In_1483);
and U4650 (N_4650,In_40,In_1247);
and U4651 (N_4651,In_507,In_1141);
and U4652 (N_4652,In_507,In_1176);
nand U4653 (N_4653,In_805,In_1358);
or U4654 (N_4654,In_1175,In_795);
or U4655 (N_4655,In_576,In_746);
or U4656 (N_4656,In_606,In_1109);
or U4657 (N_4657,In_1247,In_868);
nor U4658 (N_4658,In_778,In_342);
nor U4659 (N_4659,In_1290,In_1424);
and U4660 (N_4660,In_1371,In_923);
nand U4661 (N_4661,In_370,In_31);
nor U4662 (N_4662,In_875,In_312);
nor U4663 (N_4663,In_500,In_306);
nor U4664 (N_4664,In_1327,In_283);
nor U4665 (N_4665,In_200,In_740);
nor U4666 (N_4666,In_805,In_968);
or U4667 (N_4667,In_971,In_399);
or U4668 (N_4668,In_167,In_378);
or U4669 (N_4669,In_1325,In_696);
and U4670 (N_4670,In_338,In_1432);
nand U4671 (N_4671,In_1421,In_1203);
nor U4672 (N_4672,In_1336,In_395);
nor U4673 (N_4673,In_1133,In_1230);
and U4674 (N_4674,In_481,In_1204);
and U4675 (N_4675,In_487,In_1201);
nor U4676 (N_4676,In_337,In_920);
nor U4677 (N_4677,In_1255,In_978);
or U4678 (N_4678,In_510,In_1075);
nand U4679 (N_4679,In_404,In_1173);
and U4680 (N_4680,In_615,In_903);
or U4681 (N_4681,In_256,In_1056);
and U4682 (N_4682,In_443,In_484);
and U4683 (N_4683,In_1382,In_1142);
or U4684 (N_4684,In_1446,In_1167);
and U4685 (N_4685,In_619,In_1146);
nor U4686 (N_4686,In_1163,In_1285);
or U4687 (N_4687,In_862,In_486);
and U4688 (N_4688,In_888,In_416);
nor U4689 (N_4689,In_465,In_832);
or U4690 (N_4690,In_747,In_573);
or U4691 (N_4691,In_1189,In_193);
and U4692 (N_4692,In_962,In_754);
nor U4693 (N_4693,In_1388,In_653);
nor U4694 (N_4694,In_251,In_187);
or U4695 (N_4695,In_144,In_456);
or U4696 (N_4696,In_1129,In_807);
nand U4697 (N_4697,In_369,In_627);
or U4698 (N_4698,In_140,In_897);
or U4699 (N_4699,In_884,In_581);
and U4700 (N_4700,In_43,In_1414);
nor U4701 (N_4701,In_1406,In_1296);
or U4702 (N_4702,In_436,In_160);
nor U4703 (N_4703,In_964,In_319);
nand U4704 (N_4704,In_139,In_456);
nor U4705 (N_4705,In_1020,In_1375);
and U4706 (N_4706,In_61,In_763);
or U4707 (N_4707,In_160,In_69);
or U4708 (N_4708,In_658,In_342);
nand U4709 (N_4709,In_215,In_1208);
or U4710 (N_4710,In_158,In_418);
nand U4711 (N_4711,In_1468,In_636);
or U4712 (N_4712,In_1314,In_275);
nor U4713 (N_4713,In_814,In_1137);
and U4714 (N_4714,In_190,In_702);
nor U4715 (N_4715,In_707,In_933);
nand U4716 (N_4716,In_565,In_1126);
and U4717 (N_4717,In_192,In_138);
and U4718 (N_4718,In_734,In_1423);
or U4719 (N_4719,In_884,In_478);
or U4720 (N_4720,In_756,In_909);
or U4721 (N_4721,In_1161,In_196);
nor U4722 (N_4722,In_1499,In_958);
and U4723 (N_4723,In_237,In_506);
and U4724 (N_4724,In_1308,In_352);
nor U4725 (N_4725,In_1266,In_1180);
nor U4726 (N_4726,In_27,In_345);
nand U4727 (N_4727,In_138,In_1006);
or U4728 (N_4728,In_318,In_1487);
nor U4729 (N_4729,In_1046,In_1256);
nor U4730 (N_4730,In_537,In_1096);
nor U4731 (N_4731,In_1103,In_1225);
nor U4732 (N_4732,In_683,In_462);
nor U4733 (N_4733,In_864,In_1033);
nand U4734 (N_4734,In_909,In_772);
nand U4735 (N_4735,In_1305,In_1229);
nand U4736 (N_4736,In_566,In_166);
and U4737 (N_4737,In_1367,In_1208);
and U4738 (N_4738,In_999,In_1439);
and U4739 (N_4739,In_618,In_1170);
or U4740 (N_4740,In_1065,In_382);
or U4741 (N_4741,In_1091,In_1303);
nor U4742 (N_4742,In_208,In_823);
nand U4743 (N_4743,In_1087,In_1217);
nand U4744 (N_4744,In_1294,In_724);
and U4745 (N_4745,In_1082,In_643);
nor U4746 (N_4746,In_340,In_354);
nand U4747 (N_4747,In_521,In_727);
and U4748 (N_4748,In_906,In_57);
nor U4749 (N_4749,In_889,In_428);
nor U4750 (N_4750,In_89,In_21);
xor U4751 (N_4751,In_831,In_1350);
nor U4752 (N_4752,In_351,In_596);
nand U4753 (N_4753,In_92,In_949);
nor U4754 (N_4754,In_1297,In_770);
nand U4755 (N_4755,In_947,In_200);
or U4756 (N_4756,In_457,In_1165);
nor U4757 (N_4757,In_1233,In_66);
or U4758 (N_4758,In_1017,In_1480);
nor U4759 (N_4759,In_1433,In_566);
and U4760 (N_4760,In_1293,In_537);
nand U4761 (N_4761,In_909,In_1062);
nand U4762 (N_4762,In_741,In_72);
nand U4763 (N_4763,In_912,In_797);
nand U4764 (N_4764,In_431,In_1016);
xor U4765 (N_4765,In_842,In_420);
nor U4766 (N_4766,In_407,In_199);
and U4767 (N_4767,In_1029,In_1056);
nor U4768 (N_4768,In_267,In_771);
nand U4769 (N_4769,In_406,In_163);
and U4770 (N_4770,In_691,In_261);
and U4771 (N_4771,In_197,In_306);
and U4772 (N_4772,In_889,In_957);
or U4773 (N_4773,In_193,In_882);
nor U4774 (N_4774,In_1037,In_1438);
or U4775 (N_4775,In_933,In_924);
xor U4776 (N_4776,In_1219,In_1423);
and U4777 (N_4777,In_666,In_714);
or U4778 (N_4778,In_713,In_83);
nor U4779 (N_4779,In_518,In_407);
xnor U4780 (N_4780,In_1139,In_1132);
and U4781 (N_4781,In_1178,In_1247);
nand U4782 (N_4782,In_1170,In_1385);
xnor U4783 (N_4783,In_546,In_258);
nand U4784 (N_4784,In_858,In_779);
and U4785 (N_4785,In_1236,In_1451);
or U4786 (N_4786,In_488,In_1087);
nand U4787 (N_4787,In_1355,In_930);
nand U4788 (N_4788,In_229,In_742);
nor U4789 (N_4789,In_231,In_1079);
nor U4790 (N_4790,In_1319,In_1052);
nand U4791 (N_4791,In_1425,In_662);
and U4792 (N_4792,In_914,In_1049);
and U4793 (N_4793,In_980,In_1210);
nand U4794 (N_4794,In_510,In_799);
nand U4795 (N_4795,In_169,In_10);
or U4796 (N_4796,In_89,In_476);
or U4797 (N_4797,In_691,In_802);
or U4798 (N_4798,In_876,In_328);
and U4799 (N_4799,In_1321,In_1294);
xnor U4800 (N_4800,In_1225,In_1448);
nand U4801 (N_4801,In_974,In_624);
or U4802 (N_4802,In_783,In_698);
nor U4803 (N_4803,In_127,In_296);
nand U4804 (N_4804,In_386,In_305);
nand U4805 (N_4805,In_601,In_243);
or U4806 (N_4806,In_1369,In_1063);
or U4807 (N_4807,In_141,In_223);
and U4808 (N_4808,In_920,In_866);
and U4809 (N_4809,In_1271,In_129);
nor U4810 (N_4810,In_986,In_56);
nor U4811 (N_4811,In_1371,In_270);
nand U4812 (N_4812,In_508,In_1364);
and U4813 (N_4813,In_1265,In_688);
or U4814 (N_4814,In_183,In_45);
and U4815 (N_4815,In_1086,In_1471);
or U4816 (N_4816,In_540,In_509);
nand U4817 (N_4817,In_287,In_309);
nand U4818 (N_4818,In_1245,In_855);
nand U4819 (N_4819,In_962,In_581);
nand U4820 (N_4820,In_599,In_25);
or U4821 (N_4821,In_49,In_1464);
nor U4822 (N_4822,In_1483,In_708);
or U4823 (N_4823,In_698,In_1013);
or U4824 (N_4824,In_231,In_750);
nor U4825 (N_4825,In_583,In_1071);
nand U4826 (N_4826,In_1048,In_472);
or U4827 (N_4827,In_696,In_327);
nand U4828 (N_4828,In_1132,In_534);
nand U4829 (N_4829,In_1395,In_1210);
nor U4830 (N_4830,In_634,In_1207);
nor U4831 (N_4831,In_1071,In_437);
and U4832 (N_4832,In_1113,In_70);
or U4833 (N_4833,In_1421,In_680);
nand U4834 (N_4834,In_624,In_1405);
and U4835 (N_4835,In_595,In_995);
and U4836 (N_4836,In_1095,In_593);
or U4837 (N_4837,In_332,In_1258);
nand U4838 (N_4838,In_561,In_697);
or U4839 (N_4839,In_239,In_1347);
or U4840 (N_4840,In_993,In_772);
and U4841 (N_4841,In_1456,In_664);
nor U4842 (N_4842,In_100,In_774);
nand U4843 (N_4843,In_305,In_934);
nand U4844 (N_4844,In_805,In_1019);
nand U4845 (N_4845,In_143,In_41);
or U4846 (N_4846,In_1407,In_595);
nor U4847 (N_4847,In_1321,In_21);
or U4848 (N_4848,In_1160,In_43);
nand U4849 (N_4849,In_1088,In_674);
nand U4850 (N_4850,In_665,In_187);
nand U4851 (N_4851,In_766,In_1020);
nor U4852 (N_4852,In_242,In_645);
nand U4853 (N_4853,In_1401,In_422);
or U4854 (N_4854,In_1305,In_68);
and U4855 (N_4855,In_235,In_1491);
or U4856 (N_4856,In_406,In_777);
or U4857 (N_4857,In_994,In_153);
or U4858 (N_4858,In_571,In_582);
xor U4859 (N_4859,In_848,In_129);
and U4860 (N_4860,In_230,In_497);
or U4861 (N_4861,In_487,In_181);
and U4862 (N_4862,In_1042,In_287);
nor U4863 (N_4863,In_799,In_1);
or U4864 (N_4864,In_1208,In_1236);
nor U4865 (N_4865,In_1029,In_1340);
or U4866 (N_4866,In_1461,In_516);
or U4867 (N_4867,In_367,In_522);
nand U4868 (N_4868,In_1255,In_1029);
or U4869 (N_4869,In_154,In_659);
nor U4870 (N_4870,In_702,In_962);
or U4871 (N_4871,In_1229,In_1368);
nor U4872 (N_4872,In_1301,In_349);
and U4873 (N_4873,In_544,In_686);
and U4874 (N_4874,In_427,In_363);
nand U4875 (N_4875,In_1464,In_801);
nor U4876 (N_4876,In_1046,In_564);
or U4877 (N_4877,In_1016,In_1083);
nor U4878 (N_4878,In_1328,In_649);
nor U4879 (N_4879,In_1035,In_835);
nand U4880 (N_4880,In_417,In_410);
nand U4881 (N_4881,In_693,In_1018);
and U4882 (N_4882,In_80,In_53);
nor U4883 (N_4883,In_166,In_33);
and U4884 (N_4884,In_713,In_824);
or U4885 (N_4885,In_640,In_974);
nand U4886 (N_4886,In_1004,In_836);
nand U4887 (N_4887,In_1261,In_95);
nor U4888 (N_4888,In_1209,In_256);
nor U4889 (N_4889,In_443,In_993);
and U4890 (N_4890,In_760,In_313);
nand U4891 (N_4891,In_186,In_72);
and U4892 (N_4892,In_956,In_316);
nor U4893 (N_4893,In_497,In_41);
nor U4894 (N_4894,In_136,In_69);
nor U4895 (N_4895,In_241,In_1174);
nand U4896 (N_4896,In_400,In_573);
and U4897 (N_4897,In_175,In_1180);
and U4898 (N_4898,In_1103,In_427);
nand U4899 (N_4899,In_866,In_393);
nor U4900 (N_4900,In_1053,In_19);
nor U4901 (N_4901,In_809,In_968);
nand U4902 (N_4902,In_326,In_1048);
or U4903 (N_4903,In_1214,In_1396);
and U4904 (N_4904,In_932,In_1304);
nor U4905 (N_4905,In_1499,In_1293);
nor U4906 (N_4906,In_918,In_83);
and U4907 (N_4907,In_1151,In_319);
or U4908 (N_4908,In_542,In_977);
or U4909 (N_4909,In_69,In_1343);
nor U4910 (N_4910,In_1312,In_742);
nor U4911 (N_4911,In_82,In_120);
nor U4912 (N_4912,In_1099,In_727);
or U4913 (N_4913,In_839,In_1451);
and U4914 (N_4914,In_297,In_1317);
xnor U4915 (N_4915,In_883,In_439);
nand U4916 (N_4916,In_322,In_379);
or U4917 (N_4917,In_712,In_1112);
nand U4918 (N_4918,In_1417,In_562);
or U4919 (N_4919,In_1333,In_393);
nand U4920 (N_4920,In_1427,In_25);
nand U4921 (N_4921,In_369,In_740);
nor U4922 (N_4922,In_495,In_247);
nand U4923 (N_4923,In_581,In_1435);
and U4924 (N_4924,In_503,In_23);
nand U4925 (N_4925,In_711,In_440);
nand U4926 (N_4926,In_398,In_1413);
or U4927 (N_4927,In_556,In_1038);
nor U4928 (N_4928,In_1026,In_627);
xor U4929 (N_4929,In_1066,In_262);
nor U4930 (N_4930,In_696,In_1076);
nor U4931 (N_4931,In_845,In_277);
and U4932 (N_4932,In_1146,In_803);
nor U4933 (N_4933,In_1228,In_361);
nor U4934 (N_4934,In_88,In_548);
nor U4935 (N_4935,In_620,In_74);
nand U4936 (N_4936,In_605,In_606);
nand U4937 (N_4937,In_784,In_1394);
nand U4938 (N_4938,In_173,In_855);
nand U4939 (N_4939,In_1146,In_1152);
or U4940 (N_4940,In_368,In_807);
and U4941 (N_4941,In_1369,In_93);
nand U4942 (N_4942,In_67,In_1148);
nor U4943 (N_4943,In_780,In_465);
or U4944 (N_4944,In_377,In_566);
or U4945 (N_4945,In_650,In_855);
and U4946 (N_4946,In_1481,In_1325);
nand U4947 (N_4947,In_1306,In_127);
or U4948 (N_4948,In_1394,In_939);
nand U4949 (N_4949,In_954,In_813);
and U4950 (N_4950,In_318,In_1113);
and U4951 (N_4951,In_704,In_693);
and U4952 (N_4952,In_897,In_391);
and U4953 (N_4953,In_153,In_1235);
or U4954 (N_4954,In_144,In_714);
nor U4955 (N_4955,In_96,In_581);
nand U4956 (N_4956,In_773,In_250);
nor U4957 (N_4957,In_1020,In_730);
or U4958 (N_4958,In_219,In_1247);
nor U4959 (N_4959,In_1206,In_1416);
nor U4960 (N_4960,In_742,In_405);
xnor U4961 (N_4961,In_177,In_566);
nor U4962 (N_4962,In_259,In_1468);
nand U4963 (N_4963,In_450,In_1063);
nor U4964 (N_4964,In_1212,In_1091);
and U4965 (N_4965,In_11,In_87);
and U4966 (N_4966,In_1268,In_1207);
nand U4967 (N_4967,In_39,In_1323);
nand U4968 (N_4968,In_1039,In_1094);
and U4969 (N_4969,In_930,In_1);
nor U4970 (N_4970,In_620,In_950);
nor U4971 (N_4971,In_782,In_176);
or U4972 (N_4972,In_51,In_373);
nand U4973 (N_4973,In_84,In_584);
or U4974 (N_4974,In_909,In_1404);
nand U4975 (N_4975,In_152,In_1369);
or U4976 (N_4976,In_1399,In_1160);
and U4977 (N_4977,In_63,In_222);
and U4978 (N_4978,In_1389,In_1025);
or U4979 (N_4979,In_816,In_858);
and U4980 (N_4980,In_1372,In_395);
nor U4981 (N_4981,In_435,In_1234);
or U4982 (N_4982,In_1425,In_361);
nor U4983 (N_4983,In_131,In_789);
and U4984 (N_4984,In_26,In_809);
nor U4985 (N_4985,In_419,In_104);
nand U4986 (N_4986,In_381,In_192);
nand U4987 (N_4987,In_1418,In_1495);
nor U4988 (N_4988,In_526,In_305);
or U4989 (N_4989,In_642,In_705);
nand U4990 (N_4990,In_57,In_554);
nor U4991 (N_4991,In_47,In_400);
nand U4992 (N_4992,In_811,In_707);
nor U4993 (N_4993,In_525,In_727);
and U4994 (N_4994,In_981,In_1146);
nor U4995 (N_4995,In_918,In_1241);
and U4996 (N_4996,In_63,In_380);
and U4997 (N_4997,In_1155,In_282);
and U4998 (N_4998,In_660,In_498);
nor U4999 (N_4999,In_763,In_1383);
nor U5000 (N_5000,N_1385,N_2499);
nand U5001 (N_5001,N_3483,N_1995);
or U5002 (N_5002,N_4126,N_841);
and U5003 (N_5003,N_3563,N_1042);
nand U5004 (N_5004,N_4585,N_1347);
nand U5005 (N_5005,N_2628,N_3816);
and U5006 (N_5006,N_2920,N_1990);
or U5007 (N_5007,N_863,N_4952);
nor U5008 (N_5008,N_1678,N_385);
nand U5009 (N_5009,N_2571,N_3450);
nor U5010 (N_5010,N_4383,N_3278);
nor U5011 (N_5011,N_3996,N_3260);
or U5012 (N_5012,N_3489,N_3494);
and U5013 (N_5013,N_1548,N_3345);
nor U5014 (N_5014,N_1834,N_4964);
and U5015 (N_5015,N_2901,N_536);
xnor U5016 (N_5016,N_1756,N_3791);
and U5017 (N_5017,N_151,N_1026);
nand U5018 (N_5018,N_1901,N_839);
and U5019 (N_5019,N_3919,N_2925);
nor U5020 (N_5020,N_3043,N_3600);
or U5021 (N_5021,N_3928,N_3209);
nor U5022 (N_5022,N_4543,N_3535);
and U5023 (N_5023,N_1640,N_4444);
nand U5024 (N_5024,N_4826,N_3534);
or U5025 (N_5025,N_4834,N_816);
or U5026 (N_5026,N_758,N_4201);
and U5027 (N_5027,N_1169,N_4986);
or U5028 (N_5028,N_4002,N_2587);
and U5029 (N_5029,N_2205,N_4266);
nand U5030 (N_5030,N_1673,N_1080);
or U5031 (N_5031,N_836,N_4994);
and U5032 (N_5032,N_4216,N_2932);
nand U5033 (N_5033,N_3789,N_2055);
or U5034 (N_5034,N_1582,N_2573);
nor U5035 (N_5035,N_3096,N_2032);
and U5036 (N_5036,N_3861,N_2503);
nand U5037 (N_5037,N_895,N_2715);
nor U5038 (N_5038,N_501,N_1105);
nand U5039 (N_5039,N_4354,N_556);
nand U5040 (N_5040,N_4907,N_4479);
nand U5041 (N_5041,N_1575,N_1109);
or U5042 (N_5042,N_1341,N_2871);
and U5043 (N_5043,N_4388,N_3267);
nand U5044 (N_5044,N_1101,N_100);
or U5045 (N_5045,N_4022,N_3007);
nor U5046 (N_5046,N_2583,N_2462);
and U5047 (N_5047,N_3117,N_709);
or U5048 (N_5048,N_2885,N_886);
nor U5049 (N_5049,N_4655,N_4620);
and U5050 (N_5050,N_3449,N_996);
nor U5051 (N_5051,N_1938,N_3812);
or U5052 (N_5052,N_1794,N_2726);
nand U5053 (N_5053,N_3960,N_1389);
or U5054 (N_5054,N_2412,N_3726);
or U5055 (N_5055,N_4694,N_2127);
and U5056 (N_5056,N_4249,N_1456);
nor U5057 (N_5057,N_1701,N_2098);
nand U5058 (N_5058,N_3474,N_4823);
nor U5059 (N_5059,N_3686,N_2816);
nand U5060 (N_5060,N_1129,N_506);
nor U5061 (N_5061,N_2543,N_1257);
and U5062 (N_5062,N_2480,N_2263);
nand U5063 (N_5063,N_3508,N_4146);
nand U5064 (N_5064,N_3648,N_358);
nor U5065 (N_5065,N_4765,N_3392);
and U5066 (N_5066,N_1335,N_305);
and U5067 (N_5067,N_2709,N_2364);
or U5068 (N_5068,N_3492,N_4874);
nand U5069 (N_5069,N_3778,N_2598);
nor U5070 (N_5070,N_1366,N_3281);
nand U5071 (N_5071,N_2842,N_4211);
xnor U5072 (N_5072,N_384,N_3417);
nand U5073 (N_5073,N_2525,N_2478);
xor U5074 (N_5074,N_4853,N_4919);
or U5075 (N_5075,N_3635,N_163);
xnor U5076 (N_5076,N_3703,N_350);
or U5077 (N_5077,N_3292,N_4367);
and U5078 (N_5078,N_167,N_630);
nand U5079 (N_5079,N_1510,N_2892);
and U5080 (N_5080,N_1626,N_2231);
and U5081 (N_5081,N_3228,N_926);
and U5082 (N_5082,N_1528,N_2728);
nand U5083 (N_5083,N_1061,N_3324);
and U5084 (N_5084,N_2563,N_3039);
nand U5085 (N_5085,N_4536,N_2176);
or U5086 (N_5086,N_1744,N_2374);
nand U5087 (N_5087,N_1937,N_2481);
and U5088 (N_5088,N_3465,N_2859);
or U5089 (N_5089,N_3030,N_3800);
nand U5090 (N_5090,N_168,N_3408);
nor U5091 (N_5091,N_1559,N_3750);
or U5092 (N_5092,N_583,N_4974);
and U5093 (N_5093,N_3943,N_3058);
or U5094 (N_5094,N_161,N_1816);
nor U5095 (N_5095,N_3366,N_2274);
and U5096 (N_5096,N_4712,N_3978);
or U5097 (N_5097,N_2259,N_1910);
or U5098 (N_5098,N_4631,N_998);
or U5099 (N_5099,N_4251,N_4077);
nand U5100 (N_5100,N_2547,N_4263);
nor U5101 (N_5101,N_65,N_451);
or U5102 (N_5102,N_4340,N_2665);
or U5103 (N_5103,N_37,N_3140);
and U5104 (N_5104,N_3380,N_27);
nand U5105 (N_5105,N_1542,N_2948);
or U5106 (N_5106,N_2201,N_2146);
or U5107 (N_5107,N_3578,N_4095);
and U5108 (N_5108,N_4108,N_4026);
nor U5109 (N_5109,N_3241,N_2003);
nand U5110 (N_5110,N_3777,N_1261);
nor U5111 (N_5111,N_4616,N_3185);
and U5112 (N_5112,N_2782,N_2985);
or U5113 (N_5113,N_4877,N_2366);
and U5114 (N_5114,N_3732,N_4165);
nor U5115 (N_5115,N_1961,N_3549);
or U5116 (N_5116,N_2335,N_4054);
nor U5117 (N_5117,N_1209,N_1228);
nand U5118 (N_5118,N_838,N_2379);
or U5119 (N_5119,N_2221,N_21);
or U5120 (N_5120,N_4041,N_2195);
nor U5121 (N_5121,N_380,N_3136);
and U5122 (N_5122,N_920,N_1386);
nand U5123 (N_5123,N_4474,N_1399);
or U5124 (N_5124,N_4295,N_2037);
nand U5125 (N_5125,N_2053,N_4961);
and U5126 (N_5126,N_1522,N_4695);
nand U5127 (N_5127,N_891,N_3505);
nor U5128 (N_5128,N_733,N_1409);
nor U5129 (N_5129,N_143,N_773);
and U5130 (N_5130,N_2220,N_2243);
nor U5131 (N_5131,N_3655,N_837);
nand U5132 (N_5132,N_4061,N_3356);
and U5133 (N_5133,N_3968,N_0);
and U5134 (N_5134,N_4330,N_2044);
nor U5135 (N_5135,N_3832,N_4649);
nor U5136 (N_5136,N_4158,N_3592);
nor U5137 (N_5137,N_1793,N_589);
nor U5138 (N_5138,N_3717,N_1507);
nor U5139 (N_5139,N_1665,N_3132);
or U5140 (N_5140,N_2271,N_3471);
and U5141 (N_5141,N_2238,N_3807);
nor U5142 (N_5142,N_4102,N_3336);
nor U5143 (N_5143,N_2991,N_4861);
nand U5144 (N_5144,N_4801,N_1384);
nor U5145 (N_5145,N_2246,N_3937);
nor U5146 (N_5146,N_1010,N_205);
or U5147 (N_5147,N_3873,N_2631);
nand U5148 (N_5148,N_748,N_3802);
xor U5149 (N_5149,N_3151,N_4074);
nor U5150 (N_5150,N_138,N_884);
and U5151 (N_5151,N_3944,N_1193);
nand U5152 (N_5152,N_1764,N_4334);
nand U5153 (N_5153,N_4854,N_3216);
and U5154 (N_5154,N_1614,N_3837);
and U5155 (N_5155,N_2818,N_4575);
or U5156 (N_5156,N_3880,N_1022);
or U5157 (N_5157,N_4972,N_4403);
and U5158 (N_5158,N_4900,N_2616);
or U5159 (N_5159,N_2953,N_749);
nand U5160 (N_5160,N_2415,N_2439);
nand U5161 (N_5161,N_2687,N_735);
nor U5162 (N_5162,N_1119,N_1600);
or U5163 (N_5163,N_2720,N_4315);
or U5164 (N_5164,N_4773,N_3990);
or U5165 (N_5165,N_762,N_1723);
nor U5166 (N_5166,N_1066,N_4879);
nand U5167 (N_5167,N_171,N_1999);
or U5168 (N_5168,N_4082,N_1486);
or U5169 (N_5169,N_1375,N_3657);
or U5170 (N_5170,N_3728,N_2472);
nand U5171 (N_5171,N_3306,N_3052);
nor U5172 (N_5172,N_4031,N_1235);
nand U5173 (N_5173,N_1234,N_4419);
or U5174 (N_5174,N_439,N_2319);
or U5175 (N_5175,N_1871,N_969);
nand U5176 (N_5176,N_905,N_2442);
and U5177 (N_5177,N_3285,N_3986);
or U5178 (N_5178,N_3116,N_1952);
and U5179 (N_5179,N_4398,N_372);
nor U5180 (N_5180,N_2361,N_474);
and U5181 (N_5181,N_1333,N_1822);
nor U5182 (N_5182,N_3537,N_775);
nor U5183 (N_5183,N_3857,N_726);
nand U5184 (N_5184,N_4921,N_19);
or U5185 (N_5185,N_2664,N_1063);
nor U5186 (N_5186,N_410,N_3053);
and U5187 (N_5187,N_1000,N_538);
nand U5188 (N_5188,N_1949,N_3407);
or U5189 (N_5189,N_4098,N_1623);
and U5190 (N_5190,N_4206,N_4154);
nand U5191 (N_5191,N_3390,N_4100);
or U5192 (N_5192,N_1391,N_10);
nand U5193 (N_5193,N_835,N_1684);
nand U5194 (N_5194,N_2018,N_2548);
or U5195 (N_5195,N_431,N_4272);
nor U5196 (N_5196,N_4566,N_1955);
or U5197 (N_5197,N_1588,N_2986);
nand U5198 (N_5198,N_3419,N_1849);
and U5199 (N_5199,N_3027,N_1459);
or U5200 (N_5200,N_3862,N_4264);
or U5201 (N_5201,N_3518,N_4567);
or U5202 (N_5202,N_1545,N_4179);
and U5203 (N_5203,N_3615,N_4762);
and U5204 (N_5204,N_1812,N_3014);
nor U5205 (N_5205,N_1305,N_2309);
and U5206 (N_5206,N_3059,N_4958);
nor U5207 (N_5207,N_4604,N_2546);
and U5208 (N_5208,N_2742,N_2040);
nand U5209 (N_5209,N_3341,N_738);
nor U5210 (N_5210,N_333,N_4938);
nor U5211 (N_5211,N_2869,N_2967);
nor U5212 (N_5212,N_1357,N_162);
nand U5213 (N_5213,N_4718,N_4020);
and U5214 (N_5214,N_1570,N_3212);
nand U5215 (N_5215,N_1795,N_3868);
nand U5216 (N_5216,N_2740,N_4906);
or U5217 (N_5217,N_4745,N_2817);
and U5218 (N_5218,N_4759,N_3332);
nand U5219 (N_5219,N_1466,N_3065);
nand U5220 (N_5220,N_1926,N_1683);
nand U5221 (N_5221,N_4121,N_2502);
nand U5222 (N_5222,N_1024,N_377);
nor U5223 (N_5223,N_4609,N_2595);
nor U5224 (N_5224,N_3593,N_1874);
or U5225 (N_5225,N_252,N_2203);
nor U5226 (N_5226,N_1358,N_1819);
or U5227 (N_5227,N_293,N_1579);
nor U5228 (N_5228,N_1254,N_1846);
or U5229 (N_5229,N_4503,N_2209);
and U5230 (N_5230,N_3439,N_2891);
nor U5231 (N_5231,N_2156,N_802);
or U5232 (N_5232,N_4587,N_2693);
or U5233 (N_5233,N_4352,N_2091);
nand U5234 (N_5234,N_1072,N_2448);
nor U5235 (N_5235,N_3491,N_2744);
nand U5236 (N_5236,N_4318,N_718);
or U5237 (N_5237,N_1173,N_2717);
or U5238 (N_5238,N_755,N_668);
or U5239 (N_5239,N_3273,N_228);
nand U5240 (N_5240,N_1093,N_676);
nor U5241 (N_5241,N_4129,N_4520);
nand U5242 (N_5242,N_867,N_4382);
nand U5243 (N_5243,N_4560,N_363);
nor U5244 (N_5244,N_3740,N_812);
and U5245 (N_5245,N_4622,N_3519);
and U5246 (N_5246,N_2192,N_1495);
and U5247 (N_5247,N_3542,N_1974);
nor U5248 (N_5248,N_3509,N_159);
and U5249 (N_5249,N_3298,N_3378);
or U5250 (N_5250,N_4528,N_4173);
or U5251 (N_5251,N_4110,N_3016);
and U5252 (N_5252,N_4013,N_2000);
or U5253 (N_5253,N_4291,N_3500);
nor U5254 (N_5254,N_1670,N_4953);
and U5255 (N_5255,N_4120,N_4664);
nand U5256 (N_5256,N_278,N_1869);
or U5257 (N_5257,N_191,N_154);
nand U5258 (N_5258,N_4410,N_3538);
nor U5259 (N_5259,N_3568,N_1798);
nand U5260 (N_5260,N_465,N_610);
and U5261 (N_5261,N_4092,N_4314);
or U5262 (N_5262,N_2660,N_2642);
nand U5263 (N_5263,N_1062,N_4946);
and U5264 (N_5264,N_3819,N_1963);
nand U5265 (N_5265,N_4579,N_1197);
and U5266 (N_5266,N_517,N_1411);
nand U5267 (N_5267,N_725,N_3259);
and U5268 (N_5268,N_1083,N_1100);
and U5269 (N_5269,N_3875,N_4621);
nor U5270 (N_5270,N_2071,N_1612);
nand U5271 (N_5271,N_3609,N_1767);
or U5272 (N_5272,N_240,N_4227);
nor U5273 (N_5273,N_3300,N_1082);
nand U5274 (N_5274,N_4784,N_3409);
and U5275 (N_5275,N_2486,N_4524);
or U5276 (N_5276,N_3435,N_2099);
or U5277 (N_5277,N_447,N_1900);
nor U5278 (N_5278,N_4839,N_4331);
and U5279 (N_5279,N_4989,N_4565);
or U5280 (N_5280,N_4637,N_4239);
and U5281 (N_5281,N_3191,N_3467);
or U5282 (N_5282,N_1480,N_761);
and U5283 (N_5283,N_33,N_395);
or U5284 (N_5284,N_1658,N_4260);
or U5285 (N_5285,N_1635,N_3351);
and U5286 (N_5286,N_1520,N_1923);
nand U5287 (N_5287,N_1643,N_3057);
or U5288 (N_5288,N_2250,N_3204);
or U5289 (N_5289,N_4420,N_1236);
or U5290 (N_5290,N_4584,N_4015);
or U5291 (N_5291,N_4626,N_489);
nand U5292 (N_5292,N_834,N_4289);
and U5293 (N_5293,N_548,N_2678);
nor U5294 (N_5294,N_2959,N_4235);
nor U5295 (N_5295,N_3301,N_1351);
or U5296 (N_5296,N_3527,N_1526);
nor U5297 (N_5297,N_2402,N_730);
and U5298 (N_5298,N_1132,N_2611);
nor U5299 (N_5299,N_1426,N_553);
nor U5300 (N_5300,N_2919,N_3804);
nor U5301 (N_5301,N_4598,N_1738);
nor U5302 (N_5302,N_4661,N_3675);
nor U5303 (N_5303,N_1425,N_4997);
or U5304 (N_5304,N_3822,N_4039);
nor U5305 (N_5305,N_915,N_2315);
nand U5306 (N_5306,N_4445,N_4673);
and U5307 (N_5307,N_2437,N_4648);
nand U5308 (N_5308,N_3774,N_2421);
xnor U5309 (N_5309,N_4732,N_2897);
and U5310 (N_5310,N_204,N_15);
nand U5311 (N_5311,N_3654,N_3397);
nand U5312 (N_5312,N_3785,N_783);
and U5313 (N_5313,N_2676,N_195);
nor U5314 (N_5314,N_304,N_4650);
or U5315 (N_5315,N_892,N_1933);
nand U5316 (N_5316,N_4777,N_4461);
or U5317 (N_5317,N_1380,N_3236);
nand U5318 (N_5318,N_3369,N_189);
nor U5319 (N_5319,N_3656,N_855);
or U5320 (N_5320,N_1291,N_1714);
or U5321 (N_5321,N_2970,N_2081);
nor U5322 (N_5322,N_4888,N_3025);
and U5323 (N_5323,N_3756,N_2941);
and U5324 (N_5324,N_4709,N_3452);
nor U5325 (N_5325,N_2574,N_4430);
nor U5326 (N_5326,N_2849,N_2917);
or U5327 (N_5327,N_2681,N_472);
and U5328 (N_5328,N_4654,N_873);
nand U5329 (N_5329,N_4666,N_2894);
or U5330 (N_5330,N_3589,N_3088);
nand U5331 (N_5331,N_2599,N_4488);
nor U5332 (N_5332,N_1262,N_1557);
and U5333 (N_5333,N_1041,N_2360);
nor U5334 (N_5334,N_639,N_655);
nand U5335 (N_5335,N_2289,N_4433);
nand U5336 (N_5336,N_185,N_4707);
and U5337 (N_5337,N_1455,N_4908);
nand U5338 (N_5338,N_2172,N_2166);
and U5339 (N_5339,N_379,N_1404);
nor U5340 (N_5340,N_1152,N_170);
or U5341 (N_5341,N_4435,N_57);
and U5342 (N_5342,N_2164,N_3823);
and U5343 (N_5343,N_1070,N_3214);
nand U5344 (N_5344,N_770,N_364);
or U5345 (N_5345,N_931,N_3904);
nand U5346 (N_5346,N_2339,N_3359);
and U5347 (N_5347,N_1571,N_4177);
or U5348 (N_5348,N_1732,N_97);
and U5349 (N_5349,N_2695,N_4164);
nor U5350 (N_5350,N_4929,N_3074);
and U5351 (N_5351,N_1472,N_1047);
nor U5352 (N_5352,N_3671,N_2990);
nor U5353 (N_5353,N_981,N_2295);
and U5354 (N_5354,N_496,N_3882);
nor U5355 (N_5355,N_2162,N_2513);
nand U5356 (N_5356,N_4651,N_4639);
nor U5357 (N_5357,N_3035,N_3068);
nor U5358 (N_5358,N_4192,N_4522);
nor U5359 (N_5359,N_1598,N_3091);
nand U5360 (N_5360,N_264,N_3806);
nor U5361 (N_5361,N_2035,N_4099);
nand U5362 (N_5362,N_3248,N_2969);
or U5363 (N_5363,N_1563,N_513);
and U5364 (N_5364,N_1986,N_3627);
nor U5365 (N_5365,N_3142,N_499);
or U5366 (N_5366,N_1506,N_4030);
nand U5367 (N_5367,N_2378,N_2786);
nand U5368 (N_5368,N_4628,N_928);
nand U5369 (N_5369,N_2692,N_3621);
and U5370 (N_5370,N_1318,N_2080);
nand U5371 (N_5371,N_2857,N_4456);
or U5372 (N_5372,N_2070,N_2479);
nand U5373 (N_5373,N_4603,N_3524);
nor U5374 (N_5374,N_699,N_2700);
nor U5375 (N_5375,N_752,N_4810);
nand U5376 (N_5376,N_1020,N_4730);
or U5377 (N_5377,N_3,N_2988);
nor U5378 (N_5378,N_2934,N_433);
nor U5379 (N_5379,N_2373,N_404);
or U5380 (N_5380,N_3961,N_590);
xnor U5381 (N_5381,N_1650,N_365);
or U5382 (N_5382,N_4999,N_3163);
and U5383 (N_5383,N_3888,N_4889);
or U5384 (N_5384,N_99,N_1709);
nor U5385 (N_5385,N_4830,N_1525);
and U5386 (N_5386,N_3174,N_2432);
or U5387 (N_5387,N_907,N_4789);
nor U5388 (N_5388,N_4337,N_3530);
or U5389 (N_5389,N_2022,N_702);
or U5390 (N_5390,N_435,N_1224);
or U5391 (N_5391,N_1975,N_4531);
and U5392 (N_5392,N_2625,N_557);
nand U5393 (N_5393,N_3282,N_2073);
and U5394 (N_5394,N_4969,N_1602);
nand U5395 (N_5395,N_2677,N_1699);
nand U5396 (N_5396,N_2034,N_2331);
nor U5397 (N_5397,N_994,N_4866);
and U5398 (N_5398,N_3689,N_1126);
nor U5399 (N_5399,N_3669,N_2673);
and U5400 (N_5400,N_2626,N_289);
nand U5401 (N_5401,N_2408,N_1097);
or U5402 (N_5402,N_66,N_2386);
or U5403 (N_5403,N_2100,N_4595);
and U5404 (N_5404,N_1927,N_3539);
and U5405 (N_5405,N_2511,N_1148);
or U5406 (N_5406,N_2468,N_2950);
and U5407 (N_5407,N_2647,N_2355);
nor U5408 (N_5408,N_479,N_3370);
or U5409 (N_5409,N_174,N_3644);
nor U5410 (N_5410,N_349,N_4629);
nand U5411 (N_5411,N_3545,N_1644);
or U5412 (N_5412,N_3735,N_468);
and U5413 (N_5413,N_2072,N_2157);
or U5414 (N_5414,N_3818,N_1988);
or U5415 (N_5415,N_4781,N_1809);
nor U5416 (N_5416,N_3325,N_505);
nor U5417 (N_5417,N_3314,N_924);
nor U5418 (N_5418,N_3275,N_3115);
nor U5419 (N_5419,N_859,N_4904);
nand U5420 (N_5420,N_1698,N_896);
nand U5421 (N_5421,N_750,N_3427);
nor U5422 (N_5422,N_44,N_1204);
nand U5423 (N_5423,N_255,N_2292);
nand U5424 (N_5424,N_3291,N_124);
nand U5425 (N_5425,N_1292,N_4296);
nor U5426 (N_5426,N_4814,N_3456);
xnor U5427 (N_5427,N_2169,N_1099);
nand U5428 (N_5428,N_525,N_2646);
nand U5429 (N_5429,N_700,N_153);
nand U5430 (N_5430,N_4829,N_196);
and U5431 (N_5431,N_3123,N_421);
nor U5432 (N_5432,N_3895,N_1958);
or U5433 (N_5433,N_1239,N_2377);
or U5434 (N_5434,N_4018,N_3160);
nand U5435 (N_5435,N_2512,N_3041);
nand U5436 (N_5436,N_587,N_1181);
and U5437 (N_5437,N_1011,N_1915);
nand U5438 (N_5438,N_211,N_3404);
nand U5439 (N_5439,N_820,N_4396);
nand U5440 (N_5440,N_272,N_2890);
nand U5441 (N_5441,N_1719,N_1511);
or U5442 (N_5442,N_4424,N_3148);
and U5443 (N_5443,N_337,N_1713);
or U5444 (N_5444,N_845,N_4691);
nand U5445 (N_5445,N_3570,N_4415);
nor U5446 (N_5446,N_4477,N_1429);
and U5447 (N_5447,N_2333,N_3649);
and U5448 (N_5448,N_4590,N_4175);
and U5449 (N_5449,N_110,N_3936);
nor U5450 (N_5450,N_4828,N_106);
nand U5451 (N_5451,N_2608,N_2452);
and U5452 (N_5452,N_4483,N_150);
nor U5453 (N_5453,N_1387,N_1448);
nor U5454 (N_5454,N_2734,N_3418);
nand U5455 (N_5455,N_1837,N_2500);
xnor U5456 (N_5456,N_1156,N_3008);
and U5457 (N_5457,N_2637,N_623);
nor U5458 (N_5458,N_3352,N_1815);
or U5459 (N_5459,N_1012,N_4321);
nand U5460 (N_5460,N_3497,N_4710);
and U5461 (N_5461,N_3573,N_1482);
nand U5462 (N_5462,N_3942,N_2337);
or U5463 (N_5463,N_4033,N_182);
nor U5464 (N_5464,N_2281,N_466);
nand U5465 (N_5465,N_3410,N_178);
or U5466 (N_5466,N_1434,N_2257);
xor U5467 (N_5467,N_3725,N_1218);
nand U5468 (N_5468,N_4172,N_2954);
xnor U5469 (N_5469,N_3313,N_3349);
and U5470 (N_5470,N_2588,N_369);
nand U5471 (N_5471,N_4343,N_1948);
and U5472 (N_5472,N_3881,N_1465);
nand U5473 (N_5473,N_1069,N_446);
and U5474 (N_5474,N_4914,N_2325);
nand U5475 (N_5475,N_3402,N_1221);
nand U5476 (N_5476,N_469,N_3820);
or U5477 (N_5477,N_2719,N_4942);
nand U5478 (N_5478,N_663,N_4449);
nand U5479 (N_5479,N_130,N_2751);
and U5480 (N_5480,N_246,N_2407);
nor U5481 (N_5481,N_2848,N_2644);
nor U5482 (N_5482,N_3926,N_3386);
and U5483 (N_5483,N_781,N_823);
or U5484 (N_5484,N_4047,N_4482);
xor U5485 (N_5485,N_3536,N_4821);
and U5486 (N_5486,N_3585,N_4669);
or U5487 (N_5487,N_3131,N_213);
nor U5488 (N_5488,N_244,N_4446);
and U5489 (N_5489,N_646,N_2980);
nor U5490 (N_5490,N_4288,N_3211);
nor U5491 (N_5491,N_4723,N_1922);
or U5492 (N_5492,N_1867,N_1946);
nand U5493 (N_5493,N_216,N_3168);
nor U5494 (N_5494,N_1604,N_3983);
and U5495 (N_5495,N_2342,N_425);
nand U5496 (N_5496,N_2519,N_416);
nor U5497 (N_5497,N_1414,N_856);
nand U5498 (N_5498,N_1483,N_4960);
nor U5499 (N_5499,N_3289,N_4364);
and U5500 (N_5500,N_2310,N_4066);
or U5501 (N_5501,N_3901,N_4996);
nand U5502 (N_5502,N_4686,N_1142);
nand U5503 (N_5503,N_28,N_3133);
or U5504 (N_5504,N_2232,N_3821);
and U5505 (N_5505,N_3765,N_378);
nand U5506 (N_5506,N_370,N_1907);
nor U5507 (N_5507,N_2194,N_2495);
and U5508 (N_5508,N_1947,N_1692);
nand U5509 (N_5509,N_1763,N_1704);
or U5510 (N_5510,N_1691,N_3327);
or U5511 (N_5511,N_847,N_3192);
and U5512 (N_5512,N_2193,N_1092);
xnor U5513 (N_5513,N_1303,N_1345);
or U5514 (N_5514,N_1799,N_3238);
nor U5515 (N_5515,N_2661,N_3257);
nand U5516 (N_5516,N_1865,N_4918);
nand U5517 (N_5517,N_2864,N_2230);
nand U5518 (N_5518,N_4842,N_1240);
nand U5519 (N_5519,N_4212,N_486);
and U5520 (N_5520,N_1605,N_2027);
and U5521 (N_5521,N_1883,N_3680);
nand U5522 (N_5522,N_736,N_1740);
nor U5523 (N_5523,N_2643,N_2888);
nand U5524 (N_5524,N_4271,N_4899);
or U5525 (N_5525,N_1583,N_1680);
and U5526 (N_5526,N_3100,N_2508);
nand U5527 (N_5527,N_1504,N_3230);
nand U5528 (N_5528,N_4797,N_3321);
nor U5529 (N_5529,N_2320,N_1788);
nor U5530 (N_5530,N_179,N_4513);
nor U5531 (N_5531,N_719,N_3139);
and U5532 (N_5532,N_2436,N_1469);
nand U5533 (N_5533,N_1308,N_1726);
and U5534 (N_5534,N_3437,N_3358);
nand U5535 (N_5535,N_2995,N_1107);
and U5536 (N_5536,N_670,N_3826);
nand U5537 (N_5537,N_1231,N_3997);
or U5538 (N_5538,N_4375,N_885);
nand U5539 (N_5539,N_3958,N_1786);
and U5540 (N_5540,N_2385,N_4376);
nor U5541 (N_5541,N_2593,N_1123);
nor U5542 (N_5542,N_4662,N_1728);
nand U5543 (N_5543,N_2084,N_299);
or U5544 (N_5544,N_4702,N_3502);
or U5545 (N_5545,N_4426,N_4511);
nand U5546 (N_5546,N_1572,N_889);
or U5547 (N_5547,N_2639,N_591);
nand U5548 (N_5548,N_2620,N_4127);
and U5549 (N_5549,N_4688,N_101);
nand U5550 (N_5550,N_1880,N_3878);
nor U5551 (N_5551,N_2494,N_1230);
nand U5552 (N_5552,N_2581,N_2460);
or U5553 (N_5553,N_41,N_4298);
or U5554 (N_5554,N_4555,N_1771);
nand U5555 (N_5555,N_4007,N_478);
and U5556 (N_5556,N_180,N_1589);
nand U5557 (N_5557,N_964,N_2210);
nand U5558 (N_5558,N_956,N_258);
or U5559 (N_5559,N_3697,N_2884);
or U5560 (N_5560,N_888,N_4804);
or U5561 (N_5561,N_4684,N_4062);
nor U5562 (N_5562,N_3165,N_1773);
and U5563 (N_5563,N_3233,N_2306);
or U5564 (N_5564,N_772,N_2819);
or U5565 (N_5565,N_2861,N_361);
or U5566 (N_5566,N_2947,N_3019);
nand U5567 (N_5567,N_4353,N_4351);
or U5568 (N_5568,N_4977,N_4094);
nor U5569 (N_5569,N_2509,N_3967);
nor U5570 (N_5570,N_2493,N_4068);
nor U5571 (N_5571,N_523,N_763);
and U5572 (N_5572,N_2304,N_1214);
nor U5573 (N_5573,N_1942,N_4577);
nor U5574 (N_5574,N_4970,N_2347);
nand U5575 (N_5575,N_4903,N_1935);
nand U5576 (N_5576,N_4507,N_1436);
nand U5577 (N_5577,N_208,N_1420);
and U5578 (N_5578,N_4740,N_1360);
nor U5579 (N_5579,N_4465,N_286);
nor U5580 (N_5580,N_1237,N_2160);
or U5581 (N_5581,N_4051,N_4612);
nor U5582 (N_5582,N_4862,N_4736);
nand U5583 (N_5583,N_1280,N_584);
nand U5584 (N_5584,N_2982,N_581);
nand U5585 (N_5585,N_4987,N_765);
nor U5586 (N_5586,N_1167,N_229);
and U5587 (N_5587,N_2128,N_4581);
nor U5588 (N_5588,N_462,N_1803);
nor U5589 (N_5589,N_2569,N_967);
or U5590 (N_5590,N_3532,N_4838);
or U5591 (N_5591,N_1941,N_2178);
and U5592 (N_5592,N_4156,N_939);
nand U5593 (N_5593,N_2125,N_934);
and U5594 (N_5594,N_51,N_3367);
and U5595 (N_5595,N_2404,N_4835);
or U5596 (N_5596,N_2933,N_4200);
nor U5597 (N_5597,N_1730,N_3095);
and U5598 (N_5598,N_1906,N_320);
nand U5599 (N_5599,N_89,N_4105);
or U5600 (N_5600,N_4226,N_1885);
or U5601 (N_5601,N_2951,N_3751);
xnor U5602 (N_5602,N_3244,N_3433);
nand U5603 (N_5603,N_2668,N_2667);
or U5604 (N_5604,N_310,N_1210);
nand U5605 (N_5605,N_4549,N_4574);
or U5606 (N_5606,N_3957,N_3460);
nand U5607 (N_5607,N_3769,N_4176);
or U5608 (N_5608,N_222,N_4317);
or U5609 (N_5609,N_2708,N_2679);
and U5610 (N_5610,N_49,N_4389);
and U5611 (N_5611,N_791,N_1558);
nor U5612 (N_5612,N_786,N_3135);
nor U5613 (N_5613,N_3242,N_2518);
and U5614 (N_5614,N_2797,N_2471);
nor U5615 (N_5615,N_132,N_4901);
nand U5616 (N_5616,N_4816,N_360);
nor U5617 (N_5617,N_1182,N_493);
nand U5618 (N_5618,N_340,N_3708);
nor U5619 (N_5619,N_3528,N_3394);
nor U5620 (N_5620,N_4390,N_2154);
or U5621 (N_5621,N_4749,N_806);
nand U5622 (N_5622,N_3032,N_1766);
or U5623 (N_5623,N_4252,N_1841);
and U5624 (N_5624,N_2622,N_1518);
nor U5625 (N_5625,N_2014,N_4016);
or U5626 (N_5626,N_503,N_3984);
and U5627 (N_5627,N_3342,N_3219);
and U5628 (N_5628,N_911,N_1121);
and U5629 (N_5629,N_1154,N_944);
or U5630 (N_5630,N_1004,N_4800);
nor U5631 (N_5631,N_588,N_3801);
nand U5632 (N_5632,N_2795,N_2900);
and U5633 (N_5633,N_1718,N_3328);
nor U5634 (N_5634,N_637,N_3286);
or U5635 (N_5635,N_516,N_1117);
or U5636 (N_5636,N_3190,N_672);
nor U5637 (N_5637,N_1125,N_1338);
or U5638 (N_5638,N_667,N_1932);
nor U5639 (N_5639,N_3613,N_807);
or U5640 (N_5640,N_599,N_2005);
nor U5641 (N_5641,N_869,N_2324);
nor U5642 (N_5642,N_2614,N_3931);
or U5643 (N_5643,N_3443,N_2489);
or U5644 (N_5644,N_1348,N_2641);
nor U5645 (N_5645,N_4072,N_3595);
nand U5646 (N_5646,N_1120,N_2228);
and U5647 (N_5647,N_1615,N_61);
and U5648 (N_5648,N_2653,N_2821);
or U5649 (N_5649,N_4378,N_3112);
and U5650 (N_5650,N_292,N_3158);
nor U5651 (N_5651,N_1594,N_2580);
or U5652 (N_5652,N_779,N_3220);
or U5653 (N_5653,N_2496,N_2039);
or U5654 (N_5654,N_26,N_3599);
or U5655 (N_5655,N_20,N_4634);
nor U5656 (N_5656,N_619,N_804);
nand U5657 (N_5657,N_3103,N_1634);
or U5658 (N_5658,N_916,N_2741);
nor U5659 (N_5659,N_3667,N_232);
nor U5660 (N_5660,N_4122,N_1002);
and U5661 (N_5661,N_4625,N_4219);
or U5662 (N_5662,N_3827,N_4870);
or U5663 (N_5663,N_393,N_3063);
nor U5664 (N_5664,N_1706,N_1336);
and U5665 (N_5665,N_1213,N_4728);
nor U5666 (N_5666,N_4135,N_2710);
nor U5667 (N_5667,N_2394,N_60);
nor U5668 (N_5668,N_1750,N_1279);
nand U5669 (N_5669,N_3579,N_1888);
nor U5670 (N_5670,N_1439,N_1928);
and U5671 (N_5671,N_1821,N_2612);
and U5672 (N_5672,N_1857,N_87);
nand U5673 (N_5673,N_4897,N_187);
and U5674 (N_5674,N_782,N_764);
nand U5675 (N_5675,N_1553,N_3196);
nand U5676 (N_5676,N_4515,N_3363);
and U5677 (N_5677,N_2383,N_2444);
nor U5678 (N_5678,N_2485,N_3205);
and U5679 (N_5679,N_3582,N_757);
nor U5680 (N_5680,N_4545,N_4161);
and U5681 (N_5681,N_4010,N_3377);
and U5682 (N_5682,N_401,N_1096);
nand U5683 (N_5683,N_118,N_4478);
nor U5684 (N_5684,N_3533,N_4852);
or U5685 (N_5685,N_2886,N_2896);
or U5686 (N_5686,N_4231,N_1285);
nor U5687 (N_5687,N_1065,N_3182);
and U5688 (N_5688,N_3659,N_294);
nor U5689 (N_5689,N_3766,N_4090);
and U5690 (N_5690,N_3485,N_4148);
or U5691 (N_5691,N_1219,N_3329);
nand U5692 (N_5692,N_4486,N_1325);
or U5693 (N_5693,N_4949,N_3704);
and U5694 (N_5694,N_4056,N_2414);
nor U5695 (N_5695,N_4402,N_4771);
or U5696 (N_5696,N_4787,N_3266);
nor U5697 (N_5697,N_2689,N_691);
nor U5698 (N_5698,N_1945,N_1653);
nand U5699 (N_5699,N_1017,N_638);
nand U5700 (N_5700,N_1300,N_4665);
or U5701 (N_5701,N_3650,N_3475);
or U5702 (N_5702,N_3181,N_4775);
and U5703 (N_5703,N_2457,N_427);
nor U5704 (N_5704,N_2020,N_3179);
nor U5705 (N_5705,N_842,N_810);
nand U5706 (N_5706,N_4348,N_711);
or U5707 (N_5707,N_2121,N_4532);
nor U5708 (N_5708,N_1994,N_978);
and U5709 (N_5709,N_4308,N_2732);
nand U5710 (N_5710,N_2584,N_355);
or U5711 (N_5711,N_3694,N_1627);
nor U5712 (N_5712,N_2026,N_3577);
nor U5713 (N_5713,N_3716,N_1059);
nand U5714 (N_5714,N_3153,N_2929);
and U5715 (N_5715,N_4310,N_4497);
and U5716 (N_5716,N_3836,N_1267);
nor U5717 (N_5717,N_1532,N_2240);
nand U5718 (N_5718,N_2475,N_4040);
and U5719 (N_5719,N_3770,N_4244);
or U5720 (N_5720,N_933,N_243);
nor U5721 (N_5721,N_3186,N_1610);
and U5722 (N_5722,N_2330,N_2912);
and U5723 (N_5723,N_2367,N_2787);
nand U5724 (N_5724,N_1752,N_3146);
nor U5725 (N_5725,N_383,N_722);
nor U5726 (N_5726,N_1301,N_227);
or U5727 (N_5727,N_2697,N_4405);
nor U5728 (N_5728,N_3885,N_1783);
or U5729 (N_5729,N_4300,N_311);
nor U5730 (N_5730,N_2317,N_4915);
or U5731 (N_5731,N_2570,N_1866);
or U5732 (N_5732,N_4819,N_4955);
and U5733 (N_5733,N_852,N_3900);
nor U5734 (N_5734,N_2036,N_2430);
and U5735 (N_5735,N_42,N_356);
and U5736 (N_5736,N_1215,N_2057);
nor U5737 (N_5737,N_3101,N_4825);
nor U5738 (N_5738,N_776,N_1823);
or U5739 (N_5739,N_4186,N_1071);
nand U5740 (N_5740,N_1886,N_3884);
or U5741 (N_5741,N_3548,N_4453);
and U5742 (N_5742,N_3724,N_1685);
nand U5743 (N_5743,N_1792,N_2820);
and U5744 (N_5744,N_4674,N_923);
nand U5745 (N_5745,N_4692,N_73);
nand U5746 (N_5746,N_3564,N_4408);
nor U5747 (N_5747,N_2536,N_2976);
or U5748 (N_5748,N_4573,N_3365);
or U5749 (N_5749,N_4586,N_4931);
nor U5750 (N_5750,N_277,N_3779);
and U5751 (N_5751,N_3304,N_1086);
nor U5752 (N_5752,N_1877,N_3811);
nand U5753 (N_5753,N_1960,N_1970);
or U5754 (N_5754,N_2841,N_3541);
or U5755 (N_5755,N_4758,N_1541);
and U5756 (N_5756,N_3256,N_2380);
and U5757 (N_5757,N_3482,N_1211);
nor U5758 (N_5758,N_4046,N_1687);
and U5759 (N_5759,N_3626,N_560);
nor U5760 (N_5760,N_3540,N_3664);
nor U5761 (N_5761,N_3362,N_4134);
nand U5762 (N_5762,N_695,N_335);
and U5763 (N_5763,N_4633,N_3287);
and U5764 (N_5764,N_2123,N_3490);
nand U5765 (N_5765,N_3155,N_242);
nand U5766 (N_5766,N_592,N_4769);
nand U5767 (N_5767,N_833,N_1031);
nor U5768 (N_5768,N_1238,N_1272);
and U5769 (N_5769,N_4860,N_3620);
or U5770 (N_5770,N_4582,N_3247);
nor U5771 (N_5771,N_1151,N_3556);
and U5772 (N_5772,N_2694,N_4190);
or U5773 (N_5773,N_2305,N_1882);
or U5774 (N_5774,N_2839,N_2108);
xor U5775 (N_5775,N_248,N_626);
and U5776 (N_5776,N_1367,N_283);
or U5777 (N_5777,N_2657,N_2730);
nor U5778 (N_5778,N_8,N_1920);
and U5779 (N_5779,N_3744,N_4882);
and U5780 (N_5780,N_492,N_3784);
or U5781 (N_5781,N_1198,N_3302);
nor U5782 (N_5782,N_1478,N_4163);
and U5783 (N_5783,N_2273,N_1484);
nor U5784 (N_5784,N_4841,N_2217);
nor U5785 (N_5785,N_4205,N_848);
nor U5786 (N_5786,N_1140,N_4253);
nand U5787 (N_5787,N_2952,N_3742);
xnor U5788 (N_5788,N_2069,N_4021);
nor U5789 (N_5789,N_4706,N_4391);
or U5790 (N_5790,N_464,N_3470);
or U5791 (N_5791,N_2576,N_1074);
nor U5792 (N_5792,N_3299,N_3623);
nor U5793 (N_5793,N_526,N_1524);
or U5794 (N_5794,N_3330,N_918);
nor U5795 (N_5795,N_937,N_3020);
nand U5796 (N_5796,N_2208,N_3188);
or U5797 (N_5797,N_4911,N_2945);
nand U5798 (N_5798,N_617,N_2356);
or U5799 (N_5799,N_1645,N_813);
and U5800 (N_5800,N_606,N_2898);
and U5801 (N_5801,N_504,N_4910);
xnor U5802 (N_5802,N_144,N_1695);
nor U5803 (N_5803,N_3619,N_4459);
or U5804 (N_5804,N_514,N_4541);
and U5805 (N_5805,N_2895,N_2556);
or U5806 (N_5806,N_1659,N_4847);
or U5807 (N_5807,N_25,N_1006);
nand U5808 (N_5808,N_2759,N_1925);
nor U5809 (N_5809,N_357,N_4323);
nor U5810 (N_5810,N_212,N_771);
nand U5811 (N_5811,N_4362,N_4538);
or U5812 (N_5812,N_3023,N_4407);
nand U5813 (N_5813,N_3975,N_113);
and U5814 (N_5814,N_428,N_3754);
and U5815 (N_5815,N_1094,N_2926);
nor U5816 (N_5816,N_1836,N_2046);
or U5817 (N_5817,N_3894,N_4069);
nor U5818 (N_5818,N_4413,N_551);
and U5819 (N_5819,N_3580,N_2618);
nor U5820 (N_5820,N_2640,N_4181);
nor U5821 (N_5821,N_3495,N_671);
and U5822 (N_5822,N_2190,N_3892);
or U5823 (N_5823,N_9,N_2398);
and U5824 (N_5824,N_268,N_64);
and U5825 (N_5825,N_2224,N_2351);
or U5826 (N_5826,N_3213,N_2158);
nand U5827 (N_5827,N_795,N_4466);
xnor U5828 (N_5828,N_1533,N_2538);
or U5829 (N_5829,N_2346,N_4374);
nand U5830 (N_5830,N_4360,N_307);
and U5831 (N_5831,N_3372,N_4822);
nor U5832 (N_5832,N_2780,N_145);
and U5833 (N_5833,N_1346,N_4599);
and U5834 (N_5834,N_1811,N_152);
nand U5835 (N_5835,N_2783,N_2218);
nor U5836 (N_5836,N_3929,N_3406);
nor U5837 (N_5837,N_3145,N_2300);
or U5838 (N_5838,N_3164,N_4529);
or U5839 (N_5839,N_1371,N_598);
nor U5840 (N_5840,N_4499,N_1777);
and U5841 (N_5841,N_1765,N_131);
or U5842 (N_5842,N_2532,N_1531);
nand U5843 (N_5843,N_1838,N_220);
and U5844 (N_5844,N_3572,N_1761);
or U5845 (N_5845,N_4966,N_3786);
nor U5846 (N_5846,N_1450,N_1273);
nor U5847 (N_5847,N_2434,N_3442);
nor U5848 (N_5848,N_1276,N_403);
and U5849 (N_5849,N_1617,N_3513);
nor U5850 (N_5850,N_975,N_4349);
nor U5851 (N_5851,N_4552,N_3055);
or U5852 (N_5852,N_729,N_615);
nor U5853 (N_5853,N_2585,N_430);
nand U5854 (N_5854,N_1200,N_482);
nor U5855 (N_5855,N_4793,N_3463);
nand U5856 (N_5856,N_215,N_4656);
and U5857 (N_5857,N_3271,N_3134);
or U5858 (N_5858,N_727,N_1118);
nor U5859 (N_5859,N_4409,N_530);
nor U5860 (N_5860,N_4988,N_1527);
nor U5861 (N_5861,N_1893,N_4436);
or U5862 (N_5862,N_2696,N_2298);
nor U5863 (N_5863,N_2399,N_1818);
and U5864 (N_5864,N_2757,N_4267);
and U5865 (N_5865,N_4277,N_4157);
nand U5866 (N_5866,N_3371,N_4393);
nor U5867 (N_5867,N_1843,N_4043);
or U5868 (N_5868,N_1980,N_1260);
nor U5869 (N_5869,N_3687,N_3234);
and U5870 (N_5870,N_2147,N_1712);
nor U5871 (N_5871,N_3631,N_1021);
or U5872 (N_5872,N_1584,N_3838);
and U5873 (N_5873,N_3288,N_814);
nor U5874 (N_5874,N_3863,N_3798);
and U5875 (N_5875,N_2138,N_1134);
nor U5876 (N_5876,N_3560,N_614);
nor U5877 (N_5877,N_3641,N_3783);
and U5878 (N_5878,N_2750,N_3172);
nand U5879 (N_5879,N_1269,N_4241);
nand U5880 (N_5880,N_3601,N_4887);
nand U5881 (N_5881,N_2019,N_3064);
nor U5882 (N_5882,N_529,N_1014);
nand U5883 (N_5883,N_454,N_4432);
and U5884 (N_5884,N_4329,N_3102);
and U5885 (N_5885,N_4856,N_3974);
and U5886 (N_5886,N_2149,N_893);
or U5887 (N_5887,N_4752,N_3520);
nor U5888 (N_5888,N_3554,N_1166);
or U5889 (N_5889,N_1641,N_1067);
nand U5890 (N_5890,N_4000,N_946);
nand U5891 (N_5891,N_2735,N_1861);
nand U5892 (N_5892,N_1611,N_2997);
or U5893 (N_5893,N_4905,N_4926);
and U5894 (N_5894,N_3221,N_175);
nor U5895 (N_5895,N_3834,N_1757);
nand U5896 (N_5896,N_4619,N_2516);
nand U5897 (N_5897,N_4290,N_3468);
nor U5898 (N_5898,N_4589,N_2812);
nand U5899 (N_5899,N_50,N_4036);
or U5900 (N_5900,N_3890,N_2277);
and U5901 (N_5901,N_1076,N_2140);
nor U5902 (N_5902,N_3312,N_2459);
nor U5903 (N_5903,N_543,N_3350);
or U5904 (N_5904,N_4194,N_225);
nand U5905 (N_5905,N_1251,N_4070);
and U5906 (N_5906,N_4554,N_1898);
and U5907 (N_5907,N_657,N_2303);
xor U5908 (N_5908,N_4139,N_3217);
and U5909 (N_5909,N_4370,N_239);
or U5910 (N_5910,N_3337,N_4320);
nand U5911 (N_5911,N_3739,N_2702);
or U5912 (N_5912,N_3683,N_2297);
and U5913 (N_5913,N_4191,N_940);
nand U5914 (N_5914,N_1930,N_3898);
or U5915 (N_5915,N_1468,N_2866);
or U5916 (N_5916,N_4434,N_2136);
nand U5917 (N_5917,N_4233,N_4471);
nand U5918 (N_5918,N_4485,N_950);
nor U5919 (N_5919,N_3718,N_4115);
nor U5920 (N_5920,N_2977,N_2586);
or U5921 (N_5921,N_2168,N_3226);
and U5922 (N_5922,N_2843,N_3169);
nor U5923 (N_5923,N_4876,N_792);
and U5924 (N_5924,N_3856,N_4417);
nor U5925 (N_5925,N_4437,N_2749);
or U5926 (N_5926,N_1929,N_230);
nor U5927 (N_5927,N_3993,N_3081);
and U5928 (N_5928,N_705,N_397);
nor U5929 (N_5929,N_488,N_4848);
nand U5930 (N_5930,N_2348,N_1403);
and U5931 (N_5931,N_1274,N_2011);
and U5932 (N_5932,N_1500,N_3381);
nor U5933 (N_5933,N_2180,N_2778);
and U5934 (N_5934,N_3938,N_3633);
nor U5935 (N_5935,N_580,N_4725);
nand U5936 (N_5936,N_1973,N_3775);
and U5937 (N_5937,N_2179,N_2200);
and U5938 (N_5938,N_1157,N_1390);
and U5939 (N_5939,N_547,N_4954);
nor U5940 (N_5940,N_984,N_4761);
nand U5941 (N_5941,N_279,N_528);
or U5942 (N_5942,N_4073,N_3969);
nand U5943 (N_5943,N_734,N_1033);
nand U5944 (N_5944,N_3061,N_4670);
and U5945 (N_5945,N_109,N_4505);
nand U5946 (N_5946,N_1807,N_2999);
or U5947 (N_5947,N_4788,N_2328);
and U5948 (N_5948,N_203,N_342);
and U5949 (N_5949,N_4681,N_4473);
and U5950 (N_5950,N_3396,N_4058);
nor U5951 (N_5951,N_3653,N_3889);
or U5952 (N_5952,N_4255,N_1477);
nand U5953 (N_5953,N_4293,N_233);
nand U5954 (N_5954,N_2527,N_4232);
and U5955 (N_5955,N_3591,N_1774);
or U5956 (N_5956,N_2077,N_2323);
nand U5957 (N_5957,N_3232,N_3691);
and U5958 (N_5958,N_2853,N_4299);
or U5959 (N_5959,N_231,N_36);
or U5960 (N_5960,N_3021,N_4057);
and U5961 (N_5961,N_2860,N_4183);
or U5962 (N_5962,N_1647,N_527);
nand U5963 (N_5963,N_192,N_3464);
or U5964 (N_5964,N_1720,N_2863);
or U5965 (N_5965,N_686,N_4799);
nand U5966 (N_5966,N_4307,N_3089);
nor U5967 (N_5967,N_879,N_4611);
nand U5968 (N_5968,N_4635,N_2921);
and U5969 (N_5969,N_4228,N_221);
or U5970 (N_5970,N_563,N_3598);
nand U5971 (N_5971,N_2248,N_434);
and U5972 (N_5972,N_1161,N_4884);
and U5973 (N_5973,N_3322,N_2141);
nand U5974 (N_5974,N_4583,N_325);
nand U5975 (N_5975,N_3009,N_2187);
nor U5976 (N_5976,N_3147,N_3038);
or U5977 (N_5977,N_2237,N_4377);
and U5978 (N_5978,N_509,N_1832);
nor U5979 (N_5979,N_3012,N_4717);
nor U5980 (N_5980,N_3905,N_1593);
and U5981 (N_5981,N_4731,N_930);
nor U5982 (N_5982,N_1535,N_794);
nand U5983 (N_5983,N_2979,N_2773);
or U5984 (N_5984,N_3031,N_613);
and U5985 (N_5985,N_183,N_4050);
and U5986 (N_5986,N_652,N_2350);
nand U5987 (N_5987,N_1789,N_1697);
or U5988 (N_5988,N_1707,N_3079);
nor U5989 (N_5989,N_199,N_2723);
and U5990 (N_5990,N_2183,N_1188);
nor U5991 (N_5991,N_344,N_4411);
nand U5992 (N_5992,N_4333,N_470);
nor U5993 (N_5993,N_643,N_3000);
or U5994 (N_5994,N_1830,N_1689);
or U5995 (N_5995,N_850,N_3507);
and U5996 (N_5996,N_4336,N_1220);
and U5997 (N_5997,N_381,N_965);
or U5998 (N_5998,N_1555,N_2680);
and U5999 (N_5999,N_4737,N_3712);
or U6000 (N_6000,N_3952,N_3886);
nor U6001 (N_6001,N_2804,N_3590);
nand U6002 (N_6002,N_2753,N_1636);
nor U6003 (N_6003,N_1191,N_3246);
or U6004 (N_6004,N_1258,N_4246);
and U6005 (N_6005,N_3877,N_1015);
or U6006 (N_6006,N_4103,N_2186);
or U6007 (N_6007,N_1199,N_120);
nand U6008 (N_6008,N_1564,N_4509);
and U6009 (N_6009,N_4849,N_3698);
nand U6010 (N_6010,N_45,N_621);
nand U6011 (N_6011,N_4372,N_3412);
nor U6012 (N_6012,N_2048,N_103);
nand U6013 (N_6013,N_4152,N_3566);
or U6014 (N_6014,N_1581,N_1413);
and U6015 (N_6015,N_1060,N_122);
or U6016 (N_6016,N_46,N_2572);
or U6017 (N_6017,N_194,N_4475);
nand U6018 (N_6018,N_3663,N_4936);
nand U6019 (N_6019,N_4229,N_4658);
nand U6020 (N_6020,N_2001,N_1038);
nor U6021 (N_6021,N_4806,N_3416);
nand U6022 (N_6022,N_2061,N_3274);
and U6023 (N_6023,N_3105,N_4138);
nor U6024 (N_6024,N_2204,N_4355);
and U6025 (N_6025,N_3829,N_4481);
nor U6026 (N_6026,N_12,N_4783);
nand U6027 (N_6027,N_1470,N_1521);
nor U6028 (N_6028,N_3632,N_843);
nand U6029 (N_6029,N_4425,N_568);
nor U6030 (N_6030,N_4431,N_4803);
nand U6031 (N_6031,N_2251,N_2962);
and U6032 (N_6032,N_1551,N_4846);
nor U6033 (N_6033,N_1562,N_1772);
and U6034 (N_6034,N_1863,N_4223);
or U6035 (N_6035,N_1519,N_4504);
nand U6036 (N_6036,N_1590,N_3897);
nand U6037 (N_6037,N_3504,N_417);
nand U6038 (N_6038,N_708,N_2731);
or U6039 (N_6039,N_4753,N_105);
nor U6040 (N_6040,N_1538,N_39);
nand U6041 (N_6041,N_4517,N_4594);
and U6042 (N_6042,N_1331,N_4894);
nand U6043 (N_6043,N_3989,N_1782);
nor U6044 (N_6044,N_3876,N_1233);
or U6045 (N_6045,N_4371,N_3383);
and U6046 (N_6046,N_3389,N_3730);
nand U6047 (N_6047,N_3166,N_3488);
and U6048 (N_6048,N_4469,N_3307);
nor U6049 (N_6049,N_3584,N_1055);
nand U6050 (N_6050,N_4489,N_415);
nor U6051 (N_6051,N_4395,N_3254);
xnor U6052 (N_6052,N_83,N_4067);
nor U6053 (N_6053,N_1796,N_4282);
and U6054 (N_6054,N_575,N_744);
nand U6055 (N_6055,N_1441,N_339);
or U6056 (N_6056,N_904,N_329);
and U6057 (N_6057,N_919,N_2307);
and U6058 (N_6058,N_3646,N_3250);
and U6059 (N_6059,N_210,N_4309);
and U6060 (N_6060,N_4680,N_407);
and U6061 (N_6061,N_4676,N_2601);
nand U6062 (N_6062,N_2845,N_259);
xor U6063 (N_6063,N_2426,N_1686);
nor U6064 (N_6064,N_2344,N_3373);
and U6065 (N_6065,N_2701,N_367);
nand U6066 (N_6066,N_941,N_586);
nand U6067 (N_6067,N_1851,N_717);
or U6068 (N_6068,N_4945,N_2906);
nor U6069 (N_6069,N_4247,N_6);
and U6070 (N_6070,N_1207,N_4556);
nand U6071 (N_6071,N_851,N_3245);
or U6072 (N_6072,N_4935,N_868);
or U6073 (N_6073,N_4898,N_1302);
nor U6074 (N_6074,N_2770,N_4167);
or U6075 (N_6075,N_4813,N_3771);
nand U6076 (N_6076,N_1225,N_1735);
or U6077 (N_6077,N_2139,N_2766);
nor U6078 (N_6078,N_4230,N_4303);
nand U6079 (N_6079,N_2287,N_4498);
nand U6080 (N_6080,N_3127,N_3098);
nor U6081 (N_6081,N_4940,N_7);
nor U6082 (N_6082,N_3431,N_487);
nand U6083 (N_6083,N_4422,N_3973);
or U6084 (N_6084,N_554,N_3747);
nand U6085 (N_6085,N_2984,N_3364);
and U6086 (N_6086,N_373,N_4492);
xnor U6087 (N_6087,N_3277,N_81);
nand U6088 (N_6088,N_3210,N_2206);
nand U6089 (N_6089,N_4064,N_1394);
xnor U6090 (N_6090,N_408,N_2089);
nor U6091 (N_6091,N_3603,N_1284);
nand U6092 (N_6092,N_2805,N_2362);
nand U6093 (N_6093,N_3970,N_2245);
nand U6094 (N_6094,N_3316,N_1315);
nand U6095 (N_6095,N_1058,N_3760);
or U6096 (N_6096,N_1128,N_2409);
or U6097 (N_6097,N_2603,N_4166);
or U6098 (N_6098,N_3072,N_3514);
and U6099 (N_6099,N_1784,N_366);
nor U6100 (N_6100,N_2110,N_4236);
and U6101 (N_6101,N_3354,N_871);
nor U6102 (N_6102,N_2975,N_552);
nor U6103 (N_6103,N_1137,N_1595);
and U6104 (N_6104,N_4399,N_1515);
and U6105 (N_6105,N_3085,N_1657);
and U6106 (N_6106,N_3643,N_2792);
and U6107 (N_6107,N_480,N_2332);
or U6108 (N_6108,N_2784,N_3741);
and U6109 (N_6109,N_4867,N_2776);
nor U6110 (N_6110,N_2148,N_3637);
or U6111 (N_6111,N_4886,N_2942);
nand U6112 (N_6112,N_4869,N_62);
and U6113 (N_6113,N_3831,N_2936);
nand U6114 (N_6114,N_4927,N_3954);
nor U6115 (N_6115,N_669,N_3666);
nor U6116 (N_6116,N_3318,N_4312);
nand U6117 (N_6117,N_1122,N_1677);
nor U6118 (N_6118,N_149,N_4948);
nor U6119 (N_6119,N_4356,N_540);
or U6120 (N_6120,N_2791,N_3920);
and U6121 (N_6121,N_788,N_1189);
and U6122 (N_6122,N_3355,N_2008);
and U6123 (N_6123,N_1804,N_688);
nand U6124 (N_6124,N_471,N_1586);
or U6125 (N_6125,N_914,N_1113);
nor U6126 (N_6126,N_3713,N_3682);
nand U6127 (N_6127,N_3896,N_3731);
nand U6128 (N_6128,N_4512,N_3374);
or U6129 (N_6129,N_2109,N_405);
nor U6130 (N_6130,N_3152,N_2117);
and U6131 (N_6131,N_3734,N_3202);
and U6132 (N_6132,N_200,N_442);
nor U6133 (N_6133,N_172,N_3612);
xnor U6134 (N_6134,N_4811,N_3013);
and U6135 (N_6135,N_2649,N_3700);
and U6136 (N_6136,N_346,N_945);
nor U6137 (N_6137,N_3264,N_1565);
nand U6138 (N_6138,N_3634,N_56);
nor U6139 (N_6139,N_4168,N_774);
nand U6140 (N_6140,N_625,N_3093);
nor U6141 (N_6141,N_4171,N_1362);
and U6142 (N_6142,N_3845,N_4028);
xnor U6143 (N_6143,N_4690,N_800);
nand U6144 (N_6144,N_741,N_1155);
or U6145 (N_6145,N_991,N_308);
nand U6146 (N_6146,N_43,N_125);
nor U6147 (N_6147,N_1388,N_808);
and U6148 (N_6148,N_426,N_1943);
nand U6149 (N_6149,N_4151,N_3249);
nand U6150 (N_6150,N_4824,N_983);
or U6151 (N_6151,N_585,N_986);
nand U6152 (N_6152,N_1810,N_1244);
or U6153 (N_6153,N_1913,N_849);
nor U6154 (N_6154,N_1902,N_2654);
or U6155 (N_6155,N_579,N_4741);
nor U6156 (N_6156,N_2137,N_2382);
nand U6157 (N_6157,N_3276,N_1194);
or U6158 (N_6158,N_441,N_133);
nand U6159 (N_6159,N_2425,N_1298);
or U6160 (N_6160,N_1030,N_1044);
or U6161 (N_6161,N_2249,N_1668);
xor U6162 (N_6162,N_3587,N_2107);
and U6163 (N_6163,N_1028,N_4);
nor U6164 (N_6164,N_4733,N_2579);
nor U6165 (N_6165,N_3073,N_687);
and U6166 (N_6166,N_3860,N_1656);
or U6167 (N_6167,N_2092,N_2767);
nor U6168 (N_6168,N_173,N_2131);
or U6169 (N_6169,N_977,N_1596);
and U6170 (N_6170,N_3709,N_4893);
or U6171 (N_6171,N_3796,N_1401);
or U6172 (N_6172,N_3565,N_1530);
or U6173 (N_6173,N_651,N_681);
nand U6174 (N_6174,N_4843,N_424);
and U6175 (N_6175,N_351,N_2021);
nand U6176 (N_6176,N_1025,N_4965);
nand U6177 (N_6177,N_1475,N_4418);
nand U6178 (N_6178,N_4495,N_3814);
and U6179 (N_6179,N_2010,N_3121);
nor U6180 (N_6180,N_644,N_2417);
or U6181 (N_6181,N_2703,N_302);
nand U6182 (N_6182,N_515,N_2650);
nand U6183 (N_6183,N_3237,N_4093);
or U6184 (N_6184,N_860,N_3479);
nand U6185 (N_6185,N_2597,N_1035);
and U6186 (N_6186,N_3458,N_2714);
or U6187 (N_6187,N_549,N_3379);
xnor U6188 (N_6188,N_1824,N_2909);
nor U6189 (N_6189,N_714,N_947);
nand U6190 (N_6190,N_1311,N_3658);
and U6191 (N_6191,N_1502,N_1508);
or U6192 (N_6192,N_4081,N_4208);
or U6193 (N_6193,N_2222,N_4932);
nand U6194 (N_6194,N_1485,N_4130);
nand U6195 (N_6195,N_3618,N_2858);
nand U6196 (N_6196,N_4001,N_4442);
nor U6197 (N_6197,N_4204,N_3391);
or U6198 (N_6198,N_1835,N_942);
and U6199 (N_6199,N_756,N_787);
nor U6200 (N_6200,N_4934,N_332);
and U6201 (N_6201,N_1246,N_4197);
nand U6202 (N_6202,N_1802,N_2867);
nand U6203 (N_6203,N_2461,N_1314);
nand U6204 (N_6204,N_1546,N_825);
and U6205 (N_6205,N_3795,N_1864);
nand U6206 (N_6206,N_1639,N_1694);
and U6207 (N_6207,N_331,N_1591);
or U6208 (N_6208,N_3525,N_4005);
nor U6209 (N_6209,N_3149,N_2278);
or U6210 (N_6210,N_2550,N_1232);
and U6211 (N_6211,N_1433,N_742);
nor U6212 (N_6212,N_2120,N_4902);
nor U6213 (N_6213,N_936,N_4701);
or U6214 (N_6214,N_4273,N_4464);
nand U6215 (N_6215,N_4302,N_4976);
nor U6216 (N_6216,N_1609,N_4802);
nand U6217 (N_6217,N_3864,N_3347);
nand U6218 (N_6218,N_2431,N_4748);
nor U6219 (N_6219,N_2725,N_198);
and U6220 (N_6220,N_1467,N_2214);
nand U6221 (N_6221,N_266,N_2393);
or U6222 (N_6222,N_330,N_2318);
nor U6223 (N_6223,N_1587,N_4049);
and U6224 (N_6224,N_3137,N_280);
nor U6225 (N_6225,N_306,N_2283);
nor U6226 (N_6226,N_2809,N_4279);
nand U6227 (N_6227,N_2549,N_116);
and U6228 (N_6228,N_4140,N_241);
nand U6229 (N_6229,N_1277,N_2779);
or U6230 (N_6230,N_4913,N_1372);
nor U6231 (N_6231,N_1460,N_2291);
and U6232 (N_6232,N_1009,N_2043);
and U6233 (N_6233,N_1075,N_476);
or U6234 (N_6234,N_362,N_532);
nor U6235 (N_6235,N_3029,N_4865);
nand U6236 (N_6236,N_3476,N_4210);
nor U6237 (N_6237,N_4627,N_3076);
and U6238 (N_6238,N_2116,N_3711);
nor U6239 (N_6239,N_3054,N_1422);
and U6240 (N_6240,N_2052,N_1179);
or U6241 (N_6241,N_224,N_2047);
nand U6242 (N_6242,N_1354,N_2528);
nor U6243 (N_6243,N_1646,N_3569);
nand U6244 (N_6244,N_4817,N_24);
nand U6245 (N_6245,N_1785,N_4719);
nor U6246 (N_6246,N_3050,N_4959);
nor U6247 (N_6247,N_376,N_4896);
nand U6248 (N_6248,N_4294,N_4596);
nand U6249 (N_6249,N_88,N_1870);
and U6250 (N_6250,N_4880,N_3923);
nor U6251 (N_6251,N_4978,N_728);
and U6252 (N_6252,N_3842,N_831);
nand U6253 (N_6253,N_3189,N_3451);
or U6254 (N_6254,N_675,N_4357);
nand U6255 (N_6255,N_3678,N_4672);
nor U6256 (N_6256,N_4542,N_2904);
or U6257 (N_6257,N_1800,N_3184);
and U6258 (N_6258,N_2106,N_3543);
or U6259 (N_6259,N_3049,N_2840);
and U6260 (N_6260,N_1365,N_309);
or U6261 (N_6261,N_4782,N_846);
nor U6262 (N_6262,N_4951,N_1417);
and U6263 (N_6263,N_2798,N_3696);
or U6264 (N_6264,N_423,N_3776);
nand U6265 (N_6265,N_3672,N_2066);
or U6266 (N_6266,N_3413,N_4470);
nand U6267 (N_6267,N_4791,N_2419);
nor U6268 (N_6268,N_453,N_2012);
nand U6269 (N_6269,N_2799,N_1294);
or U6270 (N_6270,N_3586,N_4301);
and U6271 (N_6271,N_4222,N_534);
and U6272 (N_6272,N_4990,N_3086);
nand U6273 (N_6273,N_4404,N_4613);
or U6274 (N_6274,N_4150,N_1711);
nor U6275 (N_6275,N_2923,N_4716);
nand U6276 (N_6276,N_3297,N_2545);
nor U6277 (N_6277,N_1696,N_4225);
or U6278 (N_6278,N_2875,N_666);
and U6279 (N_6279,N_2113,N_3559);
and U6280 (N_6280,N_1136,N_262);
or U6281 (N_6281,N_1853,N_2197);
xnor U6282 (N_6282,N_3200,N_1517);
and U6283 (N_6283,N_3887,N_317);
nand U6284 (N_6284,N_3824,N_2134);
nor U6285 (N_6285,N_184,N_2617);
or U6286 (N_6286,N_1578,N_1150);
and U6287 (N_6287,N_2882,N_4858);
nor U6288 (N_6288,N_903,N_4742);
and U6289 (N_6289,N_3748,N_1939);
nand U6290 (N_6290,N_4097,N_3930);
or U6291 (N_6291,N_4160,N_2363);
and U6292 (N_6292,N_4644,N_3839);
nand U6293 (N_6293,N_4571,N_4133);
nand U6294 (N_6294,N_3486,N_2727);
nand U6295 (N_6295,N_1255,N_4017);
or U6296 (N_6296,N_3308,N_2633);
or U6297 (N_6297,N_2338,N_3951);
nor U6298 (N_6298,N_2049,N_4327);
or U6299 (N_6299,N_1632,N_3915);
and U6300 (N_6300,N_5,N_594);
or U6301 (N_6301,N_4141,N_1911);
or U6302 (N_6302,N_2946,N_3454);
nand U6303 (N_6303,N_2604,N_664);
and U6304 (N_6304,N_2226,N_412);
nand U6305 (N_6305,N_2235,N_1875);
and U6306 (N_6306,N_2865,N_3780);
nor U6307 (N_6307,N_4614,N_4346);
or U6308 (N_6308,N_4116,N_4045);
and U6309 (N_6309,N_2989,N_1839);
or U6310 (N_6310,N_117,N_938);
nand U6311 (N_6311,N_511,N_1852);
or U6312 (N_6312,N_3150,N_1747);
nand U6313 (N_6313,N_1881,N_811);
and U6314 (N_6314,N_34,N_281);
or U6315 (N_6315,N_1135,N_3866);
nand U6316 (N_6316,N_3628,N_2748);
nor U6317 (N_6317,N_2655,N_4257);
and U6318 (N_6318,N_2241,N_2793);
or U6319 (N_6319,N_2589,N_4698);
nand U6320 (N_6320,N_119,N_1081);
and U6321 (N_6321,N_2159,N_1158);
nand U6322 (N_6322,N_160,N_4075);
and U6323 (N_6323,N_3772,N_390);
and U6324 (N_6324,N_2862,N_2463);
nor U6325 (N_6325,N_878,N_3959);
and U6326 (N_6326,N_4677,N_3581);
and U6327 (N_6327,N_604,N_3625);
or U6328 (N_6328,N_2207,N_2596);
nor U6329 (N_6329,N_1098,N_53);
or U6330 (N_6330,N_2410,N_2009);
or U6331 (N_6331,N_4630,N_992);
nand U6332 (N_6332,N_135,N_2267);
nand U6333 (N_6333,N_2627,N_1164);
and U6334 (N_6334,N_3911,N_629);
and U6335 (N_6335,N_4209,N_2652);
nor U6336 (N_6336,N_52,N_2520);
or U6337 (N_6337,N_3075,N_4142);
or U6338 (N_6338,N_2067,N_4798);
or U6339 (N_6339,N_1287,N_1592);
nor U6340 (N_6340,N_2474,N_4746);
and U6341 (N_6341,N_2229,N_1440);
nor U6342 (N_6342,N_3561,N_784);
nand U6343 (N_6343,N_2577,N_3526);
or U6344 (N_6344,N_3604,N_314);
nor U6345 (N_6345,N_2096,N_2931);
and U6346 (N_6346,N_4550,N_3719);
or U6347 (N_6347,N_206,N_607);
nor U6348 (N_6348,N_1956,N_3516);
nand U6349 (N_6349,N_3126,N_1023);
or U6350 (N_6350,N_3893,N_176);
nor U6351 (N_6351,N_267,N_2181);
nor U6352 (N_6352,N_3067,N_4984);
nand U6353 (N_6353,N_3714,N_3319);
nand U6354 (N_6354,N_1702,N_1087);
nor U6355 (N_6355,N_1392,N_4917);
and U6356 (N_6356,N_3833,N_2998);
nand U6357 (N_6357,N_642,N_3562);
nand U6358 (N_6358,N_3434,N_1127);
nand U6359 (N_6359,N_2555,N_3255);
or U6360 (N_6360,N_768,N_1299);
or U6361 (N_6361,N_4660,N_680);
xnor U6362 (N_6362,N_3858,N_743);
and U6363 (N_6363,N_3909,N_1717);
or U6364 (N_6364,N_4198,N_2956);
nand U6365 (N_6365,N_3673,N_1724);
nand U6366 (N_6366,N_649,N_4452);
nand U6367 (N_6367,N_291,N_1981);
and U6368 (N_6368,N_2171,N_1755);
nand U6369 (N_6369,N_3156,N_1084);
nor U6370 (N_6370,N_987,N_2030);
nor U6371 (N_6371,N_3692,N_2949);
or U6372 (N_6372,N_4667,N_3120);
nor U6373 (N_6373,N_94,N_1991);
nor U6374 (N_6374,N_4659,N_2705);
or U6375 (N_6375,N_1293,N_1170);
and U6376 (N_6376,N_4240,N_1271);
and U6377 (N_6377,N_660,N_4591);
nor U6378 (N_6378,N_1496,N_976);
or U6379 (N_6379,N_2253,N_1638);
nor U6380 (N_6380,N_2392,N_3106);
and U6381 (N_6381,N_3668,N_2754);
xor U6382 (N_6382,N_2458,N_30);
nor U6383 (N_6383,N_953,N_628);
nor U6384 (N_6384,N_2592,N_4366);
or U6385 (N_6385,N_3966,N_4079);
or U6386 (N_6386,N_2395,N_4930);
or U6387 (N_6387,N_2054,N_4044);
and U6388 (N_6388,N_2400,N_297);
or U6389 (N_6389,N_4533,N_4607);
or U6390 (N_6390,N_490,N_3729);
nor U6391 (N_6391,N_80,N_3722);
nand U6392 (N_6392,N_518,N_4850);
nor U6393 (N_6393,N_2544,N_2491);
nand U6394 (N_6394,N_319,N_2082);
or U6395 (N_6395,N_4729,N_445);
or U6396 (N_6396,N_2827,N_2288);
nand U6397 (N_6397,N_2807,N_4941);
nor U6398 (N_6398,N_3640,N_2764);
or U6399 (N_6399,N_853,N_2965);
nor U6400 (N_6400,N_1342,N_1778);
nand U6401 (N_6401,N_2674,N_3972);
and U6402 (N_6402,N_1606,N_3208);
xor U6403 (N_6403,N_3998,N_1652);
nand U6404 (N_6404,N_2971,N_1003);
or U6405 (N_6405,N_2698,N_4820);
nand U6406 (N_6406,N_2236,N_1895);
and U6407 (N_6407,N_261,N_4646);
nor U6408 (N_6408,N_4350,N_4071);
nand U6409 (N_6409,N_3154,N_298);
nand U6410 (N_6410,N_524,N_4693);
nand U6411 (N_6411,N_1498,N_2635);
or U6412 (N_6412,N_1934,N_988);
nand U6413 (N_6413,N_620,N_4202);
and U6414 (N_6414,N_4467,N_2889);
nor U6415 (N_6415,N_1918,N_1437);
and U6416 (N_6416,N_455,N_1250);
and U6417 (N_6417,N_3340,N_2182);
nand U6418 (N_6418,N_3187,N_2524);
or U6419 (N_6419,N_4258,N_4760);
and U6420 (N_6420,N_2691,N_4547);
or U6421 (N_6421,N_634,N_2114);
or U6422 (N_6422,N_2844,N_1534);
or U6423 (N_6423,N_2568,N_2170);
and U6424 (N_6424,N_3426,N_951);
nand U6425 (N_6425,N_3040,N_1398);
nor U6426 (N_6426,N_4909,N_202);
nor U6427 (N_6427,N_4786,N_4184);
and U6428 (N_6428,N_402,N_4450);
nor U6429 (N_6429,N_4387,N_2666);
and U6430 (N_6430,N_4540,N_2762);
nor U6431 (N_6431,N_2258,N_4118);
nand U6432 (N_6432,N_2063,N_2847);
or U6433 (N_6433,N_4414,N_3401);
or U6434 (N_6434,N_3071,N_1628);
nand U6435 (N_6435,N_2806,N_4034);
xnor U6436 (N_6436,N_2023,N_1451);
or U6437 (N_6437,N_1264,N_1854);
nor U6438 (N_6438,N_4578,N_1177);
and U6439 (N_6439,N_440,N_2938);
xor U6440 (N_6440,N_1501,N_32);
or U6441 (N_6441,N_3947,N_3523);
xor U6442 (N_6442,N_4734,N_1453);
and U6443 (N_6443,N_4306,N_2247);
or U6444 (N_6444,N_4107,N_4128);
xnor U6445 (N_6445,N_4416,N_2007);
nand U6446 (N_6446,N_3080,N_3515);
and U6447 (N_6447,N_1330,N_4569);
and U6448 (N_6448,N_3607,N_1185);
or U6449 (N_6449,N_2957,N_3268);
nor U6450 (N_6450,N_1654,N_2899);
or U6451 (N_6451,N_3925,N_1873);
nand U6452 (N_6452,N_1556,N_3953);
or U6453 (N_6453,N_4123,N_1406);
nand U6454 (N_6454,N_550,N_3171);
nor U6455 (N_6455,N_962,N_4180);
nand U6456 (N_6456,N_3854,N_822);
nand U6457 (N_6457,N_4640,N_1967);
nand U6458 (N_6458,N_4527,N_704);
and U6459 (N_6459,N_4605,N_406);
nand U6460 (N_6460,N_4992,N_3384);
and U6461 (N_6461,N_4215,N_4890);
nand U6462 (N_6462,N_3066,N_1664);
nand U6463 (N_6463,N_2358,N_47);
nor U6464 (N_6464,N_3444,N_898);
or U6465 (N_6465,N_1977,N_2944);
and U6466 (N_6466,N_3964,N_3602);
nor U6467 (N_6467,N_2837,N_3090);
or U6468 (N_6468,N_578,N_1243);
or U6469 (N_6469,N_256,N_3173);
nor U6470 (N_6470,N_759,N_4401);
and U6471 (N_6471,N_2830,N_3622);
nand U6472 (N_6472,N_2813,N_1737);
nand U6473 (N_6473,N_3846,N_3982);
nand U6474 (N_6474,N_2704,N_4980);
or U6475 (N_6475,N_2789,N_169);
and U6476 (N_6476,N_1222,N_1894);
nor U6477 (N_6477,N_840,N_1523);
nor U6478 (N_6478,N_4679,N_3034);
and U6479 (N_6479,N_4397,N_3425);
nand U6480 (N_6480,N_3141,N_96);
and U6481 (N_6481,N_1032,N_922);
nor U6482 (N_6482,N_2284,N_2006);
and U6483 (N_6483,N_1566,N_2711);
xor U6484 (N_6484,N_3124,N_3143);
nor U6485 (N_6485,N_1681,N_1987);
or U6486 (N_6486,N_1310,N_2716);
or U6487 (N_6487,N_1168,N_880);
nor U6488 (N_6488,N_2557,N_4933);
and U6489 (N_6489,N_1716,N_2987);
or U6490 (N_6490,N_59,N_1089);
nand U6491 (N_6491,N_897,N_3044);
and U6492 (N_6492,N_1962,N_3908);
and U6493 (N_6493,N_4458,N_4562);
and U6494 (N_6494,N_3077,N_971);
nor U6495 (N_6495,N_648,N_3991);
nor U6496 (N_6496,N_754,N_3917);
and U6497 (N_6497,N_494,N_2765);
or U6498 (N_6498,N_2874,N_2119);
nor U6499 (N_6499,N_2418,N_4872);
or U6500 (N_6500,N_1577,N_2768);
nand U6501 (N_6501,N_683,N_2854);
nand U6502 (N_6502,N_4523,N_3472);
and U6503 (N_6503,N_3999,N_1103);
and U6504 (N_6504,N_1779,N_1073);
and U6505 (N_6505,N_484,N_4968);
nor U6506 (N_6506,N_4832,N_3522);
or U6507 (N_6507,N_1831,N_2808);
or U6508 (N_6508,N_731,N_1007);
and U6509 (N_6509,N_3036,N_2825);
and U6510 (N_6510,N_1703,N_3197);
or U6511 (N_6511,N_2619,N_4895);
and U6512 (N_6512,N_2523,N_3343);
and U6513 (N_6513,N_828,N_654);
nor U6514 (N_6514,N_3987,N_3006);
or U6515 (N_6515,N_1917,N_2466);
or U6516 (N_6516,N_737,N_1931);
or U6517 (N_6517,N_3701,N_2836);
nor U6518 (N_6518,N_2216,N_29);
nand U6519 (N_6519,N_2567,N_303);
and U6520 (N_6520,N_4892,N_4155);
nand U6521 (N_6521,N_92,N_862);
nand U6522 (N_6522,N_2152,N_2296);
or U6523 (N_6523,N_3963,N_658);
and U6524 (N_6524,N_1769,N_4525);
nor U6525 (N_6525,N_4136,N_3395);
or U6526 (N_6526,N_18,N_2755);
and U6527 (N_6527,N_1710,N_3547);
and U6528 (N_6528,N_201,N_1982);
nor U6529 (N_6529,N_4384,N_3844);
and U6530 (N_6530,N_2135,N_3118);
or U6531 (N_6531,N_1045,N_2470);
and U6532 (N_6532,N_3720,N_1876);
nand U6533 (N_6533,N_63,N_4332);
nand U6534 (N_6534,N_3849,N_2602);
nand U6535 (N_6535,N_4006,N_1162);
nor U6536 (N_6536,N_809,N_2684);
nand U6537 (N_6537,N_3670,N_2438);
and U6538 (N_6538,N_2542,N_1307);
or U6539 (N_6539,N_1400,N_4037);
nor U6540 (N_6540,N_295,N_3531);
nand U6541 (N_6541,N_4514,N_399);
or U6542 (N_6542,N_3977,N_2);
nand U6543 (N_6543,N_1085,N_1859);
nand U6544 (N_6544,N_4052,N_2561);
nor U6545 (N_6545,N_875,N_429);
and U6546 (N_6546,N_2058,N_2334);
or U6547 (N_6547,N_4632,N_864);
or U6548 (N_6548,N_2144,N_388);
or U6549 (N_6549,N_4510,N_4193);
or U6550 (N_6550,N_4214,N_1481);
or U6551 (N_6551,N_93,N_1454);
or U6552 (N_6552,N_3512,N_2846);
and U6553 (N_6553,N_82,N_1856);
nand U6554 (N_6554,N_359,N_3630);
nor U6555 (N_6555,N_2487,N_3484);
nand U6556 (N_6556,N_801,N_4113);
or U6557 (N_6557,N_4224,N_4967);
and U6558 (N_6558,N_1474,N_1505);
or U6559 (N_6559,N_1878,N_4174);
or U6560 (N_6560,N_3610,N_1435);
and U6561 (N_6561,N_3466,N_2103);
nand U6562 (N_6562,N_4713,N_3557);
nand U6563 (N_6563,N_894,N_2262);
nor U6564 (N_6564,N_3955,N_3851);
nand U6565 (N_6565,N_2636,N_2712);
and U6566 (N_6566,N_2381,N_218);
or U6567 (N_6567,N_4568,N_1005);
nand U6568 (N_6568,N_1370,N_2371);
nor U6569 (N_6569,N_724,N_1842);
nor U6570 (N_6570,N_146,N_3761);
nor U6571 (N_6571,N_3922,N_1550);
and U6572 (N_6572,N_2428,N_2775);
nand U6573 (N_6573,N_572,N_126);
nand U6574 (N_6574,N_874,N_2051);
and U6575 (N_6575,N_4250,N_2881);
nor U6576 (N_6576,N_785,N_641);
nand U6577 (N_6577,N_2834,N_1447);
nor U6578 (N_6578,N_973,N_3348);
nor U6579 (N_6579,N_3252,N_982);
and U6580 (N_6580,N_1130,N_4125);
nand U6581 (N_6581,N_1334,N_121);
and U6582 (N_6582,N_491,N_2973);
or U6583 (N_6583,N_1078,N_4636);
or U6584 (N_6584,N_1746,N_1560);
or U6585 (N_6585,N_2497,N_495);
nand U6586 (N_6586,N_1736,N_1944);
and U6587 (N_6587,N_4572,N_3870);
and U6588 (N_6588,N_1607,N_4106);
and U6589 (N_6589,N_3428,N_4487);
nand U6590 (N_6590,N_4638,N_565);
nor U6591 (N_6591,N_899,N_4878);
nand U6592 (N_6592,N_2074,N_1544);
nor U6593 (N_6593,N_1091,N_3867);
xnor U6594 (N_6594,N_4682,N_4278);
nor U6595 (N_6595,N_1393,N_3263);
and U6596 (N_6596,N_1499,N_2260);
and U6597 (N_6597,N_4993,N_1457);
nand U6598 (N_6598,N_4570,N_1826);
and U6599 (N_6599,N_963,N_1806);
nor U6600 (N_6600,N_1266,N_2405);
or U6601 (N_6601,N_4111,N_4269);
or U6602 (N_6602,N_2690,N_3487);
nand U6603 (N_6603,N_1576,N_4652);
nor U6604 (N_6604,N_4982,N_2056);
or U6605 (N_6605,N_1682,N_2907);
nor U6606 (N_6606,N_3099,N_386);
nor U6607 (N_6607,N_2388,N_71);
and U6608 (N_6608,N_3976,N_1879);
nand U6609 (N_6609,N_2707,N_3684);
nor U6610 (N_6610,N_345,N_2042);
nand U6611 (N_6611,N_4406,N_2670);
nand U6612 (N_6612,N_457,N_1787);
and U6613 (N_6613,N_1547,N_2341);
or U6614 (N_6614,N_4502,N_753);
nand U6615 (N_6615,N_4551,N_4379);
nor U6616 (N_6616,N_3104,N_2211);
and U6617 (N_6617,N_270,N_4268);
nor U6618 (N_6618,N_1253,N_3045);
nor U6619 (N_6619,N_4083,N_901);
nor U6620 (N_6620,N_4602,N_4500);
nand U6621 (N_6621,N_2613,N_980);
or U6622 (N_6622,N_3985,N_640);
nor U6623 (N_6623,N_887,N_1540);
nand U6624 (N_6624,N_4851,N_1891);
nor U6625 (N_6625,N_69,N_4610);
nor U6626 (N_6626,N_2340,N_414);
or U6627 (N_6627,N_1715,N_2345);
nand U6628 (N_6628,N_3809,N_4496);
and U6629 (N_6629,N_1039,N_832);
or U6630 (N_6630,N_1805,N_3457);
and U6631 (N_6631,N_1405,N_1631);
nand U6632 (N_6632,N_4995,N_2076);
and U6633 (N_6633,N_1491,N_1452);
and U6634 (N_6634,N_3706,N_4207);
and U6635 (N_6635,N_1733,N_3521);
or U6636 (N_6636,N_108,N_1781);
and U6637 (N_6637,N_3753,N_2883);
nor U6638 (N_6638,N_1829,N_2422);
and U6639 (N_6639,N_4494,N_3398);
and U6640 (N_6640,N_3707,N_1057);
or U6641 (N_6641,N_2290,N_4928);
nor U6642 (N_6642,N_4576,N_3571);
nand U6643 (N_6643,N_1149,N_463);
or U6644 (N_6644,N_3339,N_3046);
or U6645 (N_6645,N_2534,N_3550);
or U6646 (N_6646,N_1229,N_2566);
nor U6647 (N_6647,N_4086,N_2033);
or U6648 (N_6648,N_2656,N_1282);
nand U6649 (N_6649,N_2256,N_4561);
and U6650 (N_6650,N_140,N_84);
nand U6651 (N_6651,N_1361,N_861);
nand U6652 (N_6652,N_347,N_1184);
nand U6653 (N_6653,N_2453,N_4606);
and U6654 (N_6654,N_1813,N_1554);
nand U6655 (N_6655,N_4096,N_4881);
and U6656 (N_6656,N_2353,N_3070);
nor U6657 (N_6657,N_4462,N_1013);
or U6658 (N_6658,N_3360,N_3436);
nor U6659 (N_6659,N_2423,N_1165);
nor U6660 (N_6660,N_3695,N_2387);
or U6661 (N_6661,N_4519,N_2777);
nor U6662 (N_6662,N_611,N_443);
or U6663 (N_6663,N_2833,N_650);
or U6664 (N_6664,N_1328,N_521);
and U6665 (N_6665,N_3477,N_4328);
or U6666 (N_6666,N_448,N_502);
and U6667 (N_6667,N_2838,N_3794);
or U6668 (N_6668,N_2372,N_1667);
nand U6669 (N_6669,N_3743,N_2747);
nand U6670 (N_6670,N_2814,N_3290);
nand U6671 (N_6671,N_4703,N_86);
or U6672 (N_6672,N_3859,N_3293);
nand U6673 (N_6673,N_2269,N_3480);
nor U6674 (N_6674,N_1064,N_1048);
nor U6675 (N_6675,N_4019,N_2565);
nor U6676 (N_6676,N_3906,N_2645);
nand U6677 (N_6677,N_3555,N_2629);
nand U6678 (N_6678,N_2173,N_2467);
nand U6679 (N_6679,N_685,N_3924);
or U6680 (N_6680,N_818,N_4101);
nor U6681 (N_6681,N_3891,N_596);
and U6682 (N_6682,N_943,N_290);
or U6683 (N_6683,N_2850,N_2403);
and U6684 (N_6684,N_3752,N_4751);
nand U6685 (N_6685,N_1397,N_247);
nand U6686 (N_6686,N_1143,N_3933);
nor U6687 (N_6687,N_3617,N_1721);
nor U6688 (N_6688,N_2908,N_4011);
or U6689 (N_6689,N_1205,N_4833);
or U6690 (N_6690,N_2492,N_4827);
nor U6691 (N_6691,N_3949,N_3597);
and U6692 (N_6692,N_2265,N_4875);
or U6693 (N_6693,N_1868,N_4048);
nor U6694 (N_6694,N_2411,N_1313);
and U6695 (N_6695,N_559,N_2826);
and U6696 (N_6696,N_830,N_4004);
or U6697 (N_6697,N_2937,N_1421);
nor U6698 (N_6698,N_1490,N_1160);
or U6699 (N_6699,N_2155,N_1827);
or U6700 (N_6700,N_3865,N_1473);
or U6701 (N_6701,N_4790,N_1252);
or U6702 (N_6702,N_3331,N_1914);
and U6703 (N_6703,N_1820,N_510);
or U6704 (N_6704,N_673,N_2266);
nor U6705 (N_6705,N_689,N_601);
or U6706 (N_6706,N_1053,N_2610);
and U6707 (N_6707,N_1768,N_546);
nand U6708 (N_6708,N_4506,N_1195);
nor U6709 (N_6709,N_2390,N_4675);
nand U6710 (N_6710,N_3421,N_3869);
and U6711 (N_6711,N_477,N_4592);
nor U6712 (N_6712,N_2456,N_4144);
nand U6713 (N_6713,N_1147,N_739);
nand U6714 (N_6714,N_450,N_3498);
and U6715 (N_6715,N_3768,N_1860);
nor U6716 (N_6716,N_1355,N_4754);
nor U6717 (N_6717,N_1376,N_1951);
nor U6718 (N_6718,N_3315,N_3459);
or U6719 (N_6719,N_271,N_2429);
nor U6720 (N_6720,N_3914,N_1479);
and U6721 (N_6721,N_2878,N_4185);
nand U6722 (N_6722,N_2966,N_197);
nand U6723 (N_6723,N_531,N_4009);
and U6724 (N_6724,N_4063,N_3847);
nor U6725 (N_6725,N_3705,N_3222);
nand U6726 (N_6726,N_4785,N_4386);
nor U6727 (N_6727,N_115,N_2913);
and U6728 (N_6728,N_1618,N_4537);
nand U6729 (N_6729,N_958,N_3231);
or U6730 (N_6730,N_1183,N_396);
nand U6731 (N_6731,N_2122,N_3994);
and U6732 (N_6732,N_2268,N_22);
nor U6733 (N_6733,N_1924,N_3129);
nand U6734 (N_6734,N_348,N_3411);
or U6735 (N_6735,N_4484,N_698);
nand U6736 (N_6736,N_2648,N_2551);
or U6737 (N_6737,N_4147,N_3481);
nand U6738 (N_6738,N_3334,N_4971);
and U6739 (N_6739,N_2752,N_935);
and U6740 (N_6740,N_1552,N_3746);
or U6741 (N_6741,N_2609,N_2199);
and U6742 (N_6742,N_3813,N_2198);
and U6743 (N_6743,N_2354,N_3125);
nor U6744 (N_6744,N_2294,N_2914);
nand U6745 (N_6745,N_3608,N_2185);
nand U6746 (N_6746,N_1382,N_2104);
nand U6747 (N_6747,N_966,N_2803);
and U6748 (N_6748,N_4159,N_1629);
and U6749 (N_6749,N_2329,N_2915);
or U6750 (N_6750,N_1537,N_1637);
or U6751 (N_6751,N_3399,N_2029);
or U6752 (N_6752,N_4985,N_190);
and U6753 (N_6753,N_4837,N_2454);
and U6754 (N_6754,N_4696,N_3159);
or U6755 (N_6755,N_3109,N_2721);
or U6756 (N_6756,N_400,N_139);
and U6757 (N_6757,N_260,N_3424);
nand U6758 (N_6758,N_3927,N_4744);
nor U6759 (N_6759,N_2312,N_2560);
nor U6760 (N_6760,N_3850,N_1725);
nor U6761 (N_6761,N_4683,N_1953);
or U6762 (N_6762,N_2659,N_1106);
nand U6763 (N_6763,N_3567,N_4726);
and U6764 (N_6764,N_3092,N_4615);
or U6765 (N_6765,N_1202,N_2369);
and U6766 (N_6766,N_104,N_4400);
and U6767 (N_6767,N_312,N_3157);
and U6768 (N_6768,N_2893,N_4491);
or U6769 (N_6769,N_432,N_778);
nor U6770 (N_6770,N_4254,N_4947);
nand U6771 (N_6771,N_2349,N_1753);
or U6772 (N_6772,N_2254,N_954);
nand U6773 (N_6773,N_1296,N_186);
nor U6774 (N_6774,N_1163,N_1674);
nand U6775 (N_6775,N_2539,N_1909);
nor U6776 (N_6776,N_4943,N_2016);
nor U6777 (N_6777,N_418,N_249);
nor U6778 (N_6778,N_3461,N_1996);
or U6779 (N_6779,N_3193,N_4280);
and U6780 (N_6780,N_285,N_2424);
nand U6781 (N_6781,N_3110,N_1329);
or U6782 (N_6782,N_2594,N_1051);
nand U6783 (N_6783,N_54,N_4657);
nor U6784 (N_6784,N_1245,N_1954);
nand U6785 (N_6785,N_3932,N_3636);
nand U6786 (N_6786,N_605,N_3114);
and U6787 (N_6787,N_4871,N_3797);
nand U6788 (N_6788,N_2994,N_1418);
nor U6789 (N_6789,N_1817,N_3871);
or U6790 (N_6790,N_1622,N_1110);
or U6791 (N_6791,N_4338,N_1993);
nand U6792 (N_6792,N_2252,N_4700);
or U6793 (N_6793,N_2810,N_512);
nand U6794 (N_6794,N_67,N_2802);
and U6795 (N_6795,N_263,N_3176);
and U6796 (N_6796,N_1461,N_2469);
or U6797 (N_6797,N_1187,N_4857);
or U6798 (N_6798,N_1529,N_1971);
or U6799 (N_6799,N_3793,N_1959);
nor U6800 (N_6800,N_254,N_3934);
or U6801 (N_6801,N_4259,N_112);
nor U6802 (N_6802,N_927,N_3017);
nor U6803 (N_6803,N_1190,N_3576);
or U6804 (N_6804,N_1896,N_3517);
and U6805 (N_6805,N_3499,N_2600);
nor U6806 (N_6806,N_2050,N_2564);
nand U6807 (N_6807,N_1741,N_1722);
nand U6808 (N_6808,N_1368,N_2314);
nor U6809 (N_6809,N_3224,N_1858);
nor U6810 (N_6810,N_2079,N_1111);
and U6811 (N_6811,N_912,N_1036);
or U6812 (N_6812,N_2958,N_1442);
nand U6813 (N_6813,N_1464,N_2443);
or U6814 (N_6814,N_4708,N_3594);
or U6815 (N_6815,N_4472,N_1217);
nor U6816 (N_6816,N_2852,N_3062);
or U6817 (N_6817,N_1908,N_1762);
or U6818 (N_6818,N_1144,N_2086);
or U6819 (N_6819,N_2308,N_4776);
or U6820 (N_6820,N_3962,N_4285);
and U6821 (N_6821,N_2124,N_158);
and U6822 (N_6822,N_77,N_760);
xor U6823 (N_6823,N_2167,N_4796);
nand U6824 (N_6824,N_3745,N_238);
and U6825 (N_6825,N_769,N_2993);
nand U6826 (N_6826,N_3757,N_2413);
nor U6827 (N_6827,N_1992,N_2974);
or U6828 (N_6828,N_2272,N_2446);
or U6829 (N_6829,N_4365,N_790);
or U6830 (N_6830,N_1145,N_166);
and U6831 (N_6831,N_2115,N_1642);
and U6832 (N_6832,N_2242,N_1428);
nor U6833 (N_6833,N_2658,N_164);
nand U6834 (N_6834,N_3913,N_316);
and U6835 (N_6835,N_2504,N_631);
nand U6836 (N_6836,N_2872,N_4772);
and U6837 (N_6837,N_3357,N_1936);
or U6838 (N_6838,N_1957,N_2175);
and U6839 (N_6839,N_1008,N_1186);
nand U6840 (N_6840,N_3737,N_4025);
nand U6841 (N_6841,N_1309,N_4080);
nor U6842 (N_6842,N_3946,N_23);
nor U6843 (N_6843,N_4678,N_574);
and U6844 (N_6844,N_925,N_2142);
or U6845 (N_6845,N_4394,N_877);
nand U6846 (N_6846,N_223,N_3652);
and U6847 (N_6847,N_1319,N_1916);
and U6848 (N_6848,N_2041,N_4831);
or U6849 (N_6849,N_1489,N_2763);
or U6850 (N_6850,N_3638,N_1138);
nand U6851 (N_6851,N_2126,N_2352);
and U6852 (N_6852,N_1249,N_2713);
and U6853 (N_6853,N_2992,N_2391);
or U6854 (N_6854,N_4962,N_3047);
and U6855 (N_6855,N_2831,N_3258);
nand U6856 (N_6856,N_3645,N_3048);
nor U6857 (N_6857,N_4220,N_2311);
nor U6858 (N_6858,N_2758,N_3323);
nor U6859 (N_6859,N_1216,N_31);
and U6860 (N_6860,N_1029,N_177);
nand U6861 (N_6861,N_1206,N_3553);
or U6862 (N_6862,N_1095,N_2177);
nand U6863 (N_6863,N_707,N_2264);
nor U6864 (N_6864,N_2234,N_803);
and U6865 (N_6865,N_2718,N_1259);
nor U6866 (N_6866,N_3715,N_4304);
or U6867 (N_6867,N_4218,N_2815);
nand U6868 (N_6868,N_603,N_1381);
nor U6869 (N_6869,N_2447,N_456);
and U6870 (N_6870,N_3762,N_1043);
and U6871 (N_6871,N_98,N_4153);
and U6872 (N_6872,N_4275,N_4836);
nand U6873 (N_6873,N_1352,N_2940);
or U6874 (N_6874,N_2397,N_1049);
and U6875 (N_6875,N_3710,N_4618);
nand U6876 (N_6876,N_571,N_3916);
nand U6877 (N_6877,N_653,N_2855);
nand U6878 (N_6878,N_2015,N_1159);
nor U6879 (N_6879,N_1248,N_1353);
nor U6880 (N_6880,N_566,N_3162);
and U6881 (N_6881,N_1016,N_2683);
or U6882 (N_6882,N_2233,N_1349);
and U6883 (N_6883,N_438,N_819);
nor U6884 (N_6884,N_3679,N_2774);
nand U6885 (N_6885,N_3501,N_3144);
or U6886 (N_6886,N_1019,N_4104);
or U6887 (N_6887,N_2163,N_55);
or U6888 (N_6888,N_2130,N_4641);
nand U6889 (N_6889,N_4553,N_4844);
nor U6890 (N_6890,N_2449,N_2359);
and U6891 (N_6891,N_2326,N_902);
and U6892 (N_6892,N_2722,N_4735);
nand U6893 (N_6893,N_3223,N_1494);
or U6894 (N_6894,N_2188,N_857);
and U6895 (N_6895,N_301,N_865);
or U6896 (N_6896,N_1288,N_3128);
xor U6897 (N_6897,N_2133,N_2515);
nor U6898 (N_6898,N_157,N_2510);
nand U6899 (N_6899,N_4335,N_3320);
and U6900 (N_6900,N_519,N_1174);
or U6901 (N_6901,N_1905,N_1972);
or U6902 (N_6902,N_4137,N_2420);
and U6903 (N_6903,N_368,N_4441);
nor U6904 (N_6904,N_1412,N_76);
nand U6905 (N_6905,N_4325,N_4624);
nor U6906 (N_6906,N_970,N_4563);
nor U6907 (N_6907,N_2632,N_535);
and U6908 (N_6908,N_4863,N_4855);
or U6909 (N_6909,N_237,N_72);
and U6910 (N_6910,N_957,N_16);
and U6911 (N_6911,N_1379,N_799);
nand U6912 (N_6912,N_1903,N_4221);
nor U6913 (N_6913,N_3629,N_1775);
nand U6914 (N_6914,N_2196,N_1306);
nor U6915 (N_6915,N_2961,N_3195);
or U6916 (N_6916,N_777,N_123);
or U6917 (N_6917,N_2416,N_2729);
or U6918 (N_6918,N_2261,N_4774);
or U6919 (N_6919,N_2031,N_354);
nor U6920 (N_6920,N_682,N_147);
or U6921 (N_6921,N_1690,N_3749);
nand U6922 (N_6922,N_692,N_3207);
nor U6923 (N_6923,N_2688,N_2552);
and U6924 (N_6924,N_4764,N_95);
or U6925 (N_6925,N_3874,N_2983);
nor U6926 (N_6926,N_3361,N_3375);
nor U6927 (N_6927,N_4248,N_2769);
nor U6928 (N_6928,N_4326,N_2477);
nor U6929 (N_6929,N_1780,N_1415);
nand U6930 (N_6930,N_1567,N_4864);
nor U6931 (N_6931,N_485,N_4739);
nand U6932 (N_6932,N_452,N_2161);
xnor U6933 (N_6933,N_4261,N_1133);
nand U6934 (N_6934,N_4029,N_2605);
nand U6935 (N_6935,N_4920,N_315);
nand U6936 (N_6936,N_997,N_3677);
nand U6937 (N_6937,N_1897,N_4412);
nand U6938 (N_6938,N_701,N_677);
or U6939 (N_6939,N_1950,N_1825);
nand U6940 (N_6940,N_2675,N_1408);
nand U6941 (N_6941,N_2427,N_1613);
or U6942 (N_6942,N_3941,N_3382);
and U6943 (N_6943,N_3387,N_3662);
or U6944 (N_6944,N_4963,N_883);
nor U6945 (N_6945,N_3681,N_3511);
and U6946 (N_6946,N_1808,N_3852);
nor U6947 (N_6947,N_3574,N_4170);
or U6948 (N_6948,N_3119,N_1373);
and U6949 (N_6949,N_2800,N_1471);
nor U6950 (N_6950,N_2737,N_3283);
or U6951 (N_6951,N_4023,N_2922);
or U6952 (N_6952,N_2095,N_1889);
nand U6953 (N_6953,N_3130,N_1619);
nor U6954 (N_6954,N_1052,N_2013);
or U6955 (N_6955,N_829,N_1077);
nor U6956 (N_6956,N_3616,N_2505);
and U6957 (N_6957,N_4359,N_1289);
nand U6958 (N_6958,N_1343,N_636);
nand U6959 (N_6959,N_2153,N_1312);
nand U6960 (N_6960,N_4084,N_1172);
or U6961 (N_6961,N_3660,N_300);
nand U6962 (N_6962,N_1585,N_2856);
nor U6963 (N_6963,N_3309,N_1);
or U6964 (N_6964,N_188,N_3503);
nor U6965 (N_6965,N_1979,N_3198);
nand U6966 (N_6966,N_3400,N_2963);
and U6967 (N_6967,N_4003,N_422);
or U6968 (N_6968,N_1027,N_789);
nand U6969 (N_6969,N_3883,N_4345);
nand U6970 (N_6970,N_1630,N_4979);
nor U6971 (N_6971,N_2851,N_3215);
and U6972 (N_6972,N_507,N_3736);
and U6973 (N_6973,N_2464,N_411);
nand U6974 (N_6974,N_2623,N_2064);
and U6975 (N_6975,N_274,N_4286);
or U6976 (N_6976,N_3980,N_3551);
nand U6977 (N_6977,N_703,N_2672);
nand U6978 (N_6978,N_1175,N_3024);
and U6979 (N_6979,N_4245,N_1374);
nand U6980 (N_6980,N_2498,N_3755);
and U6981 (N_6981,N_1845,N_1968);
or U6982 (N_6982,N_3506,N_4738);
nor U6983 (N_6983,N_4859,N_1438);
or U6984 (N_6984,N_2916,N_4392);
nor U6985 (N_6985,N_1034,N_4593);
or U6986 (N_6986,N_2943,N_989);
nand U6987 (N_6987,N_1742,N_444);
or U6988 (N_6988,N_713,N_537);
nor U6989 (N_6989,N_3326,N_3788);
and U6990 (N_6990,N_2964,N_3447);
or U6991 (N_6991,N_287,N_1976);
and U6992 (N_6992,N_322,N_4145);
and U6993 (N_6993,N_4808,N_1648);
nand U6994 (N_6994,N_3853,N_3702);
or U6995 (N_6995,N_1320,N_1223);
and U6996 (N_6996,N_2313,N_2118);
nor U6997 (N_6997,N_2433,N_3790);
nand U6998 (N_6998,N_2739,N_1791);
and U6999 (N_6999,N_4076,N_4493);
nor U7000 (N_7000,N_40,N_1488);
nand U7001 (N_7001,N_284,N_4342);
nor U7002 (N_7002,N_1904,N_1141);
and U7003 (N_7003,N_1597,N_4534);
nor U7004 (N_7004,N_2028,N_3462);
and U7005 (N_7005,N_2760,N_181);
nor U7006 (N_7006,N_1568,N_4912);
or U7007 (N_7007,N_2972,N_4975);
nand U7008 (N_7008,N_2724,N_2873);
nor U7009 (N_7009,N_4265,N_3773);
or U7010 (N_7010,N_4763,N_2105);
and U7011 (N_7011,N_2024,N_4238);
and U7012 (N_7012,N_1671,N_908);
and U7013 (N_7013,N_4608,N_1751);
nand U7014 (N_7014,N_1509,N_4143);
and U7015 (N_7015,N_3225,N_3453);
nor U7016 (N_7016,N_1350,N_1965);
and U7017 (N_7017,N_4195,N_582);
nor U7018 (N_7018,N_459,N_475);
and U7019 (N_7019,N_609,N_226);
or U7020 (N_7020,N_1844,N_573);
nor U7021 (N_7021,N_1708,N_3388);
or U7022 (N_7022,N_4199,N_3992);
or U7023 (N_7023,N_1263,N_3988);
nand U7024 (N_7024,N_4324,N_4750);
nor U7025 (N_7025,N_817,N_2276);
nand U7026 (N_7026,N_1037,N_2280);
and U7027 (N_7027,N_715,N_2829);
or U7028 (N_7028,N_2286,N_4885);
nand U7029 (N_7029,N_2085,N_1268);
nor U7030 (N_7030,N_4276,N_1383);
and U7031 (N_7031,N_3690,N_4281);
nand U7032 (N_7032,N_3910,N_3624);
and U7033 (N_7033,N_720,N_1327);
and U7034 (N_7034,N_4805,N_4187);
nand U7035 (N_7035,N_2870,N_3376);
or U7036 (N_7036,N_1662,N_3294);
or U7037 (N_7037,N_4546,N_990);
nand U7038 (N_7038,N_2075,N_2903);
nand U7039 (N_7039,N_3113,N_1731);
or U7040 (N_7040,N_2087,N_881);
nor U7041 (N_7041,N_1985,N_3799);
or U7042 (N_7042,N_2093,N_4724);
and U7043 (N_7043,N_3872,N_1580);
and U7044 (N_7044,N_622,N_2671);
xor U7045 (N_7045,N_569,N_1424);
nand U7046 (N_7046,N_4380,N_35);
nand U7047 (N_7047,N_1378,N_624);
and U7048 (N_7048,N_313,N_961);
nand U7049 (N_7049,N_555,N_522);
nor U7050 (N_7050,N_2880,N_235);
and U7051 (N_7051,N_3203,N_1770);
and U7052 (N_7052,N_796,N_4124);
nand U7053 (N_7053,N_2738,N_4287);
xor U7054 (N_7054,N_2215,N_4642);
and U7055 (N_7055,N_2811,N_3956);
nor U7056 (N_7056,N_4767,N_296);
nor U7057 (N_7057,N_2743,N_1790);
or U7058 (N_7058,N_4998,N_2357);
nor U7059 (N_7059,N_1090,N_4780);
and U7060 (N_7060,N_273,N_2507);
and U7061 (N_7061,N_1940,N_1599);
and U7062 (N_7062,N_4645,N_1989);
nor U7063 (N_7063,N_4476,N_498);
or U7064 (N_7064,N_2090,N_3948);
nor U7065 (N_7065,N_1445,N_4687);
nand U7066 (N_7066,N_2699,N_2088);
or U7067 (N_7067,N_353,N_1407);
or U7068 (N_7068,N_2706,N_4647);
nor U7069 (N_7069,N_2559,N_1919);
nand U7070 (N_7070,N_544,N_1283);
or U7071 (N_7071,N_2517,N_4617);
or U7072 (N_7072,N_4341,N_282);
nor U7073 (N_7073,N_3808,N_2165);
nor U7074 (N_7074,N_866,N_1661);
nand U7075 (N_7075,N_375,N_3493);
or U7076 (N_7076,N_2996,N_265);
nor U7077 (N_7077,N_371,N_4580);
and U7078 (N_7078,N_4792,N_633);
nand U7079 (N_7079,N_1539,N_3368);
or U7080 (N_7080,N_343,N_2978);
nor U7081 (N_7081,N_288,N_3614);
and U7082 (N_7082,N_635,N_141);
or U7083 (N_7083,N_3177,N_4131);
nor U7084 (N_7084,N_4344,N_275);
nor U7085 (N_7085,N_2450,N_1180);
nand U7086 (N_7086,N_858,N_3022);
or U7087 (N_7087,N_4937,N_1068);
and U7088 (N_7088,N_2202,N_2322);
or U7089 (N_7089,N_561,N_4756);
or U7090 (N_7090,N_3787,N_1431);
nor U7091 (N_7091,N_3279,N_3935);
and U7092 (N_7092,N_3981,N_3251);
nor U7093 (N_7093,N_1887,N_58);
and U7094 (N_7094,N_3552,N_2065);
nand U7095 (N_7095,N_972,N_2745);
and U7096 (N_7096,N_949,N_1543);
nand U7097 (N_7097,N_1364,N_1241);
or U7098 (N_7098,N_1443,N_3764);
or U7099 (N_7099,N_4807,N_1758);
nand U7100 (N_7100,N_2327,N_4038);
nor U7101 (N_7101,N_2506,N_2455);
nor U7102 (N_7102,N_4840,N_3042);
nand U7103 (N_7103,N_155,N_3083);
or U7104 (N_7104,N_17,N_558);
and U7105 (N_7105,N_4213,N_1514);
and U7106 (N_7106,N_1449,N_2370);
and U7107 (N_7107,N_1884,N_2145);
nor U7108 (N_7108,N_890,N_4024);
nor U7109 (N_7109,N_3108,N_3005);
nand U7110 (N_7110,N_4747,N_2531);
and U7111 (N_7111,N_4778,N_1316);
nand U7112 (N_7112,N_4234,N_4564);
and U7113 (N_7113,N_1760,N_142);
nand U7114 (N_7114,N_805,N_458);
and U7115 (N_7115,N_78,N_4643);
or U7116 (N_7116,N_541,N_798);
nor U7117 (N_7117,N_2255,N_2279);
nand U7118 (N_7118,N_3004,N_128);
and U7119 (N_7119,N_4132,N_2606);
or U7120 (N_7120,N_3448,N_1124);
nor U7121 (N_7121,N_3180,N_4957);
nand U7122 (N_7122,N_678,N_1729);
and U7123 (N_7123,N_1574,N_1693);
nor U7124 (N_7124,N_3469,N_1669);
nor U7125 (N_7125,N_1018,N_4217);
or U7126 (N_7126,N_721,N_2004);
nor U7127 (N_7127,N_3767,N_1493);
nand U7128 (N_7128,N_3199,N_391);
nor U7129 (N_7129,N_1040,N_4721);
or U7130 (N_7130,N_4704,N_336);
or U7131 (N_7131,N_2435,N_1363);
or U7132 (N_7132,N_2968,N_1332);
nor U7133 (N_7133,N_1679,N_3284);
nand U7134 (N_7134,N_217,N_253);
or U7135 (N_7135,N_4883,N_38);
or U7136 (N_7136,N_3338,N_797);
and U7137 (N_7137,N_1432,N_3122);
or U7138 (N_7138,N_2097,N_3763);
and U7139 (N_7139,N_2336,N_4770);
and U7140 (N_7140,N_909,N_107);
nand U7141 (N_7141,N_2801,N_3921);
and U7142 (N_7142,N_2591,N_4557);
nor U7143 (N_7143,N_2484,N_2535);
nand U7144 (N_7144,N_1776,N_1633);
and U7145 (N_7145,N_1295,N_2094);
or U7146 (N_7146,N_1675,N_2213);
nor U7147 (N_7147,N_948,N_2662);
nand U7148 (N_7148,N_102,N_4653);
or U7149 (N_7149,N_3403,N_766);
nor U7150 (N_7150,N_3261,N_2530);
nor U7151 (N_7151,N_3415,N_4347);
nand U7152 (N_7152,N_3087,N_3529);
or U7153 (N_7153,N_2227,N_4012);
nor U7154 (N_7154,N_3965,N_1192);
or U7155 (N_7155,N_4182,N_4053);
nor U7156 (N_7156,N_1247,N_352);
and U7157 (N_7157,N_3311,N_2634);
and U7158 (N_7158,N_1208,N_1978);
or U7159 (N_7159,N_70,N_1359);
nor U7160 (N_7160,N_3335,N_1290);
or U7161 (N_7161,N_1444,N_2736);
or U7162 (N_7162,N_2129,N_1621);
or U7163 (N_7163,N_960,N_3971);
nand U7164 (N_7164,N_3699,N_3446);
nor U7165 (N_7165,N_4809,N_4711);
nand U7166 (N_7166,N_127,N_2316);
or U7167 (N_7167,N_4516,N_1104);
and U7168 (N_7168,N_4369,N_4008);
and U7169 (N_7169,N_1212,N_1921);
or U7170 (N_7170,N_219,N_4922);
nor U7171 (N_7171,N_2924,N_740);
nand U7172 (N_7172,N_3546,N_632);
nand U7173 (N_7173,N_952,N_4526);
or U7174 (N_7174,N_3674,N_2554);
nor U7175 (N_7175,N_793,N_4319);
nor U7176 (N_7176,N_321,N_732);
nor U7177 (N_7177,N_2045,N_4597);
nor U7178 (N_7178,N_4112,N_993);
and U7179 (N_7179,N_564,N_612);
and U7180 (N_7180,N_3782,N_1828);
nand U7181 (N_7181,N_4274,N_4311);
nor U7182 (N_7182,N_85,N_4697);
and U7183 (N_7183,N_2025,N_3423);
xnor U7184 (N_7184,N_712,N_4455);
nor U7185 (N_7185,N_4448,N_1833);
nand U7186 (N_7186,N_2219,N_3262);
nor U7187 (N_7187,N_4429,N_1046);
or U7188 (N_7188,N_2835,N_2638);
nand U7189 (N_7189,N_409,N_4623);
nand U7190 (N_7190,N_68,N_4544);
nand U7191 (N_7191,N_3841,N_148);
nor U7192 (N_7192,N_1487,N_844);
nand U7193 (N_7193,N_4262,N_4868);
or U7194 (N_7194,N_985,N_3803);
or U7195 (N_7195,N_3606,N_1281);
and U7196 (N_7196,N_4457,N_3206);
nand U7197 (N_7197,N_684,N_3478);
nand U7198 (N_7198,N_4270,N_2368);
or U7199 (N_7199,N_13,N_389);
nand U7200 (N_7200,N_1323,N_3950);
nand U7201 (N_7201,N_2935,N_1672);
or U7202 (N_7202,N_382,N_4671);
and U7203 (N_7203,N_1171,N_2615);
nor U7204 (N_7204,N_4663,N_3272);
or U7205 (N_7205,N_4795,N_3685);
or U7206 (N_7206,N_2002,N_4109);
nor U7207 (N_7207,N_129,N_679);
or U7208 (N_7208,N_4117,N_4727);
or U7209 (N_7209,N_3879,N_3758);
nand U7210 (N_7210,N_900,N_1969);
xnor U7211 (N_7211,N_2772,N_4973);
and U7212 (N_7212,N_1340,N_665);
nand U7213 (N_7213,N_2537,N_1056);
nor U7214 (N_7214,N_3405,N_1322);
nand U7215 (N_7215,N_1326,N_500);
nand U7216 (N_7216,N_2150,N_3227);
nor U7217 (N_7217,N_2239,N_4950);
nor U7218 (N_7218,N_2501,N_3018);
and U7219 (N_7219,N_3438,N_1396);
and U7220 (N_7220,N_4845,N_1700);
and U7221 (N_7221,N_1419,N_3011);
nor U7222 (N_7222,N_1054,N_4428);
nand U7223 (N_7223,N_4983,N_723);
and U7224 (N_7224,N_3253,N_1964);
and U7225 (N_7225,N_3270,N_1655);
nand U7226 (N_7226,N_1377,N_328);
and U7227 (N_7227,N_2930,N_136);
nand U7228 (N_7228,N_3828,N_1666);
and U7229 (N_7229,N_4439,N_3107);
or U7230 (N_7230,N_3792,N_627);
nor U7231 (N_7231,N_3611,N_647);
nor U7232 (N_7232,N_597,N_2375);
and U7233 (N_7233,N_79,N_1153);
and U7234 (N_7234,N_2059,N_2225);
nand U7235 (N_7235,N_3939,N_4705);
or U7236 (N_7236,N_1427,N_234);
nand U7237 (N_7237,N_1998,N_1050);
nand U7238 (N_7238,N_413,N_4812);
nor U7239 (N_7239,N_815,N_193);
nor U7240 (N_7240,N_4322,N_4316);
nand U7241 (N_7241,N_872,N_4685);
or U7242 (N_7242,N_2529,N_2396);
nor U7243 (N_7243,N_3912,N_1608);
nand U7244 (N_7244,N_1624,N_236);
or U7245 (N_7245,N_4423,N_4815);
xor U7246 (N_7246,N_1601,N_4283);
and U7247 (N_7247,N_461,N_3835);
nor U7248 (N_7248,N_1462,N_3333);
nor U7249 (N_7249,N_1112,N_1966);
nor U7250 (N_7250,N_929,N_1983);
or U7251 (N_7251,N_4313,N_2174);
or U7252 (N_7252,N_2824,N_473);
nor U7253 (N_7253,N_913,N_2384);
nand U7254 (N_7254,N_4451,N_2876);
nand U7255 (N_7255,N_1423,N_1625);
nor U7256 (N_7256,N_3688,N_4722);
and U7257 (N_7257,N_2887,N_4089);
nand U7258 (N_7258,N_693,N_2939);
and U7259 (N_7259,N_2630,N_4059);
or U7260 (N_7260,N_318,N_4521);
and U7261 (N_7261,N_2781,N_1203);
nand U7262 (N_7262,N_4440,N_3805);
nor U7263 (N_7263,N_3265,N_114);
and U7264 (N_7264,N_4518,N_1369);
or U7265 (N_7265,N_4361,N_1850);
nand U7266 (N_7266,N_4755,N_2832);
nand U7267 (N_7267,N_3015,N_3723);
nand U7268 (N_7268,N_3094,N_3239);
nand U7269 (N_7269,N_436,N_2514);
nor U7270 (N_7270,N_2796,N_539);
nor U7271 (N_7271,N_2558,N_269);
or U7272 (N_7272,N_394,N_3441);
nand U7273 (N_7273,N_4501,N_2794);
or U7274 (N_7274,N_2293,N_2756);
nand U7275 (N_7275,N_4443,N_4203);
or U7276 (N_7276,N_1603,N_1743);
and U7277 (N_7277,N_4169,N_323);
nor U7278 (N_7278,N_4284,N_1108);
nor U7279 (N_7279,N_4381,N_1227);
nor U7280 (N_7280,N_3642,N_214);
and U7281 (N_7281,N_1446,N_3440);
and U7282 (N_7282,N_4480,N_645);
nand U7283 (N_7283,N_2490,N_2686);
nor U7284 (N_7284,N_2068,N_156);
or U7285 (N_7285,N_821,N_2621);
nor U7286 (N_7286,N_3310,N_600);
nor U7287 (N_7287,N_3575,N_3945);
or U7288 (N_7288,N_4162,N_2910);
and U7289 (N_7289,N_338,N_3830);
or U7290 (N_7290,N_4588,N_3346);
nor U7291 (N_7291,N_4242,N_1759);
nor U7292 (N_7292,N_2270,N_751);
and U7293 (N_7293,N_2553,N_2321);
or U7294 (N_7294,N_4924,N_1278);
or U7295 (N_7295,N_2960,N_746);
or U7296 (N_7296,N_3496,N_1321);
or U7297 (N_7297,N_3510,N_4363);
nor U7298 (N_7298,N_1848,N_3280);
or U7299 (N_7299,N_1201,N_2651);
or U7300 (N_7300,N_4014,N_3069);
nand U7301 (N_7301,N_3240,N_4939);
nand U7302 (N_7302,N_2771,N_419);
nor U7303 (N_7303,N_3414,N_1862);
nor U7304 (N_7304,N_3344,N_780);
and U7305 (N_7305,N_595,N_690);
or U7306 (N_7306,N_74,N_542);
and U7307 (N_7307,N_3817,N_2562);
or U7308 (N_7308,N_1997,N_1649);
or U7309 (N_7309,N_2669,N_3051);
or U7310 (N_7310,N_4490,N_968);
nand U7311 (N_7311,N_910,N_3738);
nand U7312 (N_7312,N_1463,N_2682);
and U7313 (N_7313,N_1814,N_3010);
xnor U7314 (N_7314,N_3194,N_979);
nor U7315 (N_7315,N_3138,N_3161);
nor U7316 (N_7316,N_2526,N_420);
and U7317 (N_7317,N_3855,N_4601);
nand U7318 (N_7318,N_1569,N_3651);
and U7319 (N_7319,N_4916,N_2282);
and U7320 (N_7320,N_497,N_4468);
nor U7321 (N_7321,N_1324,N_387);
nand U7322 (N_7322,N_2017,N_1114);
nor U7323 (N_7323,N_2060,N_398);
and U7324 (N_7324,N_827,N_4720);
and U7325 (N_7325,N_1356,N_4178);
and U7326 (N_7326,N_4088,N_1516);
nor U7327 (N_7327,N_2521,N_616);
or U7328 (N_7328,N_90,N_4297);
or U7329 (N_7329,N_4438,N_1131);
nand U7330 (N_7330,N_562,N_4087);
nand U7331 (N_7331,N_449,N_1339);
nand U7332 (N_7332,N_4427,N_2184);
and U7333 (N_7333,N_1304,N_662);
nor U7334 (N_7334,N_1297,N_111);
nor U7335 (N_7335,N_4078,N_3037);
nor U7336 (N_7336,N_2299,N_1196);
nor U7337 (N_7337,N_4373,N_4027);
nor U7338 (N_7338,N_4256,N_1337);
nand U7339 (N_7339,N_3269,N_2905);
and U7340 (N_7340,N_1847,N_1855);
nand U7341 (N_7341,N_1270,N_4447);
or U7342 (N_7342,N_2062,N_999);
nor U7343 (N_7343,N_4243,N_2575);
and U7344 (N_7344,N_4149,N_4508);
or U7345 (N_7345,N_656,N_1739);
and U7346 (N_7346,N_4065,N_3001);
nand U7347 (N_7347,N_3825,N_1256);
and U7348 (N_7348,N_1410,N_2823);
nand U7349 (N_7349,N_4699,N_334);
nor U7350 (N_7350,N_694,N_3918);
and U7351 (N_7351,N_3596,N_2902);
nand U7352 (N_7352,N_1265,N_767);
or U7353 (N_7353,N_1115,N_4237);
nor U7354 (N_7354,N_4757,N_1727);
or U7355 (N_7355,N_2785,N_4189);
nand U7356 (N_7356,N_2285,N_392);
and U7357 (N_7357,N_3815,N_4766);
nand U7358 (N_7358,N_1651,N_1705);
or U7359 (N_7359,N_3097,N_602);
and U7360 (N_7360,N_2302,N_959);
and U7361 (N_7361,N_2761,N_2143);
and U7362 (N_7362,N_1088,N_4925);
nand U7363 (N_7363,N_4114,N_3588);
nor U7364 (N_7364,N_2981,N_134);
and U7365 (N_7365,N_921,N_4981);
or U7366 (N_7366,N_2189,N_2083);
and U7367 (N_7367,N_3033,N_1620);
nand U7368 (N_7368,N_659,N_4305);
nand U7369 (N_7369,N_2685,N_3243);
or U7370 (N_7370,N_91,N_1745);
and U7371 (N_7371,N_2102,N_4873);
nand U7372 (N_7372,N_11,N_2401);
and U7373 (N_7373,N_2151,N_995);
or U7374 (N_7374,N_3605,N_1561);
nor U7375 (N_7375,N_4559,N_3078);
nor U7376 (N_7376,N_876,N_3385);
and U7377 (N_7377,N_3843,N_710);
xnor U7378 (N_7378,N_3183,N_2522);
and U7379 (N_7379,N_1748,N_1102);
nand U7380 (N_7380,N_1001,N_3445);
and U7381 (N_7381,N_3583,N_1416);
nor U7382 (N_7382,N_706,N_4035);
nor U7383 (N_7383,N_3082,N_674);
nand U7384 (N_7384,N_2191,N_3676);
or U7385 (N_7385,N_4991,N_2445);
or U7386 (N_7386,N_1616,N_2911);
nor U7387 (N_7387,N_2038,N_2376);
and U7388 (N_7388,N_1797,N_2533);
nor U7389 (N_7389,N_3393,N_3781);
nand U7390 (N_7390,N_1663,N_2389);
or U7391 (N_7391,N_4454,N_520);
and U7392 (N_7392,N_570,N_250);
or U7393 (N_7393,N_1503,N_567);
nand U7394 (N_7394,N_3810,N_1660);
nand U7395 (N_7395,N_137,N_3028);
and U7396 (N_7396,N_2541,N_3899);
nor U7397 (N_7397,N_3903,N_1513);
or U7398 (N_7398,N_3235,N_2212);
nand U7399 (N_7399,N_3420,N_932);
and U7400 (N_7400,N_577,N_917);
nand U7401 (N_7401,N_3693,N_4292);
nand U7402 (N_7402,N_1912,N_4956);
nand U7403 (N_7403,N_696,N_1536);
nor U7404 (N_7404,N_4539,N_3995);
or U7405 (N_7405,N_3733,N_4779);
nor U7406 (N_7406,N_4891,N_906);
and U7407 (N_7407,N_1573,N_1430);
or U7408 (N_7408,N_341,N_1872);
nor U7409 (N_7409,N_1402,N_4188);
nand U7410 (N_7410,N_2928,N_2607);
nor U7411 (N_7411,N_545,N_3303);
nor U7412 (N_7412,N_4091,N_1116);
and U7413 (N_7413,N_3430,N_2582);
nor U7414 (N_7414,N_4196,N_2482);
nor U7415 (N_7415,N_3175,N_326);
nand U7416 (N_7416,N_3353,N_3317);
and U7417 (N_7417,N_618,N_661);
nand U7418 (N_7418,N_1395,N_1749);
and U7419 (N_7419,N_257,N_533);
and U7420 (N_7420,N_3544,N_1984);
or U7421 (N_7421,N_483,N_745);
or U7422 (N_7422,N_1512,N_1492);
nand U7423 (N_7423,N_2788,N_4743);
nor U7424 (N_7424,N_3167,N_324);
nor U7425 (N_7425,N_854,N_2746);
nand U7426 (N_7426,N_2473,N_697);
or U7427 (N_7427,N_3229,N_1139);
and U7428 (N_7428,N_4385,N_4358);
or U7429 (N_7429,N_3201,N_75);
or U7430 (N_7430,N_481,N_2578);
or U7431 (N_7431,N_3429,N_1146);
or U7432 (N_7432,N_1801,N_3002);
nor U7433 (N_7433,N_1688,N_327);
or U7434 (N_7434,N_4548,N_2112);
or U7435 (N_7435,N_2301,N_1476);
and U7436 (N_7436,N_882,N_2663);
nand U7437 (N_7437,N_207,N_3665);
and U7438 (N_7438,N_2877,N_3111);
and U7439 (N_7439,N_1892,N_460);
or U7440 (N_7440,N_2733,N_4368);
or U7441 (N_7441,N_3907,N_3759);
nand U7442 (N_7442,N_824,N_593);
and U7443 (N_7443,N_3026,N_467);
or U7444 (N_7444,N_2441,N_4768);
nor U7445 (N_7445,N_4055,N_747);
nand U7446 (N_7446,N_3084,N_3170);
and U7447 (N_7447,N_576,N_1176);
nor U7448 (N_7448,N_2624,N_4944);
and U7449 (N_7449,N_374,N_4085);
or U7450 (N_7450,N_4042,N_1178);
nand U7451 (N_7451,N_1079,N_4060);
or U7452 (N_7452,N_716,N_4460);
or U7453 (N_7453,N_1275,N_4715);
or U7454 (N_7454,N_3295,N_2879);
or U7455 (N_7455,N_4558,N_1286);
nand U7456 (N_7456,N_3979,N_3422);
and U7457 (N_7457,N_2540,N_2111);
nor U7458 (N_7458,N_4818,N_3455);
nor U7459 (N_7459,N_4339,N_3727);
or U7460 (N_7460,N_1317,N_3902);
and U7461 (N_7461,N_1344,N_2927);
and U7462 (N_7462,N_276,N_1242);
nand U7463 (N_7463,N_245,N_251);
nand U7464 (N_7464,N_1754,N_2406);
nor U7465 (N_7465,N_4923,N_209);
xnor U7466 (N_7466,N_4600,N_4421);
nor U7467 (N_7467,N_4119,N_3558);
and U7468 (N_7468,N_4535,N_437);
and U7469 (N_7469,N_870,N_4689);
nor U7470 (N_7470,N_2828,N_3639);
nand U7471 (N_7471,N_1226,N_3432);
and U7472 (N_7472,N_3721,N_3296);
and U7473 (N_7473,N_2451,N_1549);
nor U7474 (N_7474,N_2868,N_2365);
nand U7475 (N_7475,N_4463,N_2343);
and U7476 (N_7476,N_2822,N_826);
or U7477 (N_7477,N_2223,N_2244);
xnor U7478 (N_7478,N_3056,N_4530);
nand U7479 (N_7479,N_3305,N_3218);
nand U7480 (N_7480,N_4668,N_48);
and U7481 (N_7481,N_955,N_2488);
or U7482 (N_7482,N_3473,N_2918);
or U7483 (N_7483,N_2790,N_2955);
and U7484 (N_7484,N_4714,N_974);
or U7485 (N_7485,N_3661,N_2132);
and U7486 (N_7486,N_1458,N_3848);
and U7487 (N_7487,N_165,N_3647);
or U7488 (N_7488,N_14,N_1676);
xnor U7489 (N_7489,N_3840,N_3003);
nor U7490 (N_7490,N_3940,N_1497);
and U7491 (N_7491,N_2275,N_4794);
or U7492 (N_7492,N_2078,N_2101);
and U7493 (N_7493,N_508,N_2465);
or U7494 (N_7494,N_2590,N_1734);
and U7495 (N_7495,N_1890,N_3178);
and U7496 (N_7496,N_2483,N_3060);
and U7497 (N_7497,N_2476,N_2440);
and U7498 (N_7498,N_4032,N_1840);
and U7499 (N_7499,N_608,N_1899);
and U7500 (N_7500,N_2685,N_1632);
or U7501 (N_7501,N_253,N_4489);
nor U7502 (N_7502,N_1484,N_3053);
nand U7503 (N_7503,N_3112,N_1992);
and U7504 (N_7504,N_477,N_2507);
or U7505 (N_7505,N_4009,N_20);
nand U7506 (N_7506,N_4569,N_3407);
nand U7507 (N_7507,N_48,N_2650);
or U7508 (N_7508,N_495,N_4331);
and U7509 (N_7509,N_4859,N_1072);
or U7510 (N_7510,N_853,N_3910);
and U7511 (N_7511,N_2961,N_2463);
nor U7512 (N_7512,N_4525,N_4199);
nor U7513 (N_7513,N_3354,N_4645);
or U7514 (N_7514,N_2538,N_1056);
or U7515 (N_7515,N_1261,N_4009);
or U7516 (N_7516,N_3996,N_2278);
xor U7517 (N_7517,N_3826,N_232);
nor U7518 (N_7518,N_841,N_2937);
and U7519 (N_7519,N_2008,N_219);
and U7520 (N_7520,N_1967,N_2072);
and U7521 (N_7521,N_2071,N_2933);
and U7522 (N_7522,N_50,N_2005);
nor U7523 (N_7523,N_2898,N_1059);
nand U7524 (N_7524,N_716,N_972);
and U7525 (N_7525,N_747,N_2942);
and U7526 (N_7526,N_4648,N_4149);
nand U7527 (N_7527,N_4016,N_3218);
nand U7528 (N_7528,N_751,N_3559);
or U7529 (N_7529,N_929,N_1980);
and U7530 (N_7530,N_792,N_588);
and U7531 (N_7531,N_3834,N_640);
or U7532 (N_7532,N_4073,N_1073);
or U7533 (N_7533,N_1892,N_4307);
nor U7534 (N_7534,N_3402,N_951);
nor U7535 (N_7535,N_4049,N_2302);
nor U7536 (N_7536,N_3898,N_850);
nor U7537 (N_7537,N_3197,N_605);
nor U7538 (N_7538,N_1550,N_4071);
nand U7539 (N_7539,N_909,N_3388);
and U7540 (N_7540,N_3053,N_3054);
nor U7541 (N_7541,N_2061,N_4886);
nor U7542 (N_7542,N_4970,N_1308);
and U7543 (N_7543,N_2753,N_3883);
and U7544 (N_7544,N_3587,N_1765);
nor U7545 (N_7545,N_4025,N_121);
or U7546 (N_7546,N_4645,N_1098);
or U7547 (N_7547,N_2212,N_4020);
or U7548 (N_7548,N_4769,N_4890);
nor U7549 (N_7549,N_2960,N_1124);
or U7550 (N_7550,N_3840,N_4889);
and U7551 (N_7551,N_2123,N_305);
or U7552 (N_7552,N_3053,N_2054);
nor U7553 (N_7553,N_704,N_2830);
or U7554 (N_7554,N_2277,N_4787);
nand U7555 (N_7555,N_527,N_1403);
and U7556 (N_7556,N_4940,N_2291);
and U7557 (N_7557,N_2120,N_1815);
nand U7558 (N_7558,N_4160,N_424);
nor U7559 (N_7559,N_4275,N_2094);
nand U7560 (N_7560,N_350,N_45);
and U7561 (N_7561,N_4223,N_2171);
or U7562 (N_7562,N_651,N_391);
nand U7563 (N_7563,N_283,N_2034);
nand U7564 (N_7564,N_2487,N_275);
or U7565 (N_7565,N_1055,N_2401);
and U7566 (N_7566,N_745,N_3747);
or U7567 (N_7567,N_1962,N_934);
nand U7568 (N_7568,N_1543,N_3802);
nor U7569 (N_7569,N_426,N_3770);
nand U7570 (N_7570,N_617,N_2670);
and U7571 (N_7571,N_168,N_1496);
and U7572 (N_7572,N_2604,N_1053);
and U7573 (N_7573,N_2766,N_3223);
nor U7574 (N_7574,N_2007,N_124);
or U7575 (N_7575,N_83,N_523);
nor U7576 (N_7576,N_734,N_1264);
nor U7577 (N_7577,N_4961,N_2983);
or U7578 (N_7578,N_1390,N_2943);
nand U7579 (N_7579,N_365,N_1080);
nand U7580 (N_7580,N_2195,N_2068);
nand U7581 (N_7581,N_491,N_1537);
nand U7582 (N_7582,N_2703,N_1261);
nor U7583 (N_7583,N_4157,N_4112);
nor U7584 (N_7584,N_3916,N_920);
and U7585 (N_7585,N_4670,N_60);
and U7586 (N_7586,N_1434,N_2589);
nor U7587 (N_7587,N_2439,N_2307);
and U7588 (N_7588,N_4234,N_663);
or U7589 (N_7589,N_2967,N_2168);
or U7590 (N_7590,N_1425,N_966);
or U7591 (N_7591,N_4841,N_4401);
or U7592 (N_7592,N_3616,N_1473);
nor U7593 (N_7593,N_139,N_3656);
xnor U7594 (N_7594,N_3257,N_4703);
or U7595 (N_7595,N_2645,N_631);
or U7596 (N_7596,N_925,N_1133);
or U7597 (N_7597,N_1362,N_1634);
nand U7598 (N_7598,N_3425,N_3827);
nand U7599 (N_7599,N_2581,N_2979);
and U7600 (N_7600,N_2920,N_1694);
nand U7601 (N_7601,N_2499,N_4638);
xor U7602 (N_7602,N_1122,N_1845);
nor U7603 (N_7603,N_2007,N_2628);
nand U7604 (N_7604,N_46,N_3946);
nor U7605 (N_7605,N_1467,N_275);
and U7606 (N_7606,N_3235,N_3782);
nor U7607 (N_7607,N_2295,N_642);
and U7608 (N_7608,N_2624,N_129);
nand U7609 (N_7609,N_2314,N_4077);
nor U7610 (N_7610,N_1734,N_270);
nor U7611 (N_7611,N_363,N_4050);
or U7612 (N_7612,N_2314,N_2590);
or U7613 (N_7613,N_3303,N_1349);
nand U7614 (N_7614,N_988,N_2423);
or U7615 (N_7615,N_4080,N_2094);
or U7616 (N_7616,N_2196,N_3484);
nand U7617 (N_7617,N_3048,N_2194);
and U7618 (N_7618,N_1178,N_766);
nor U7619 (N_7619,N_4294,N_2108);
nor U7620 (N_7620,N_2153,N_1662);
nand U7621 (N_7621,N_1473,N_812);
and U7622 (N_7622,N_3147,N_4390);
nand U7623 (N_7623,N_1524,N_4830);
nand U7624 (N_7624,N_2839,N_2095);
nand U7625 (N_7625,N_3219,N_1217);
nor U7626 (N_7626,N_4752,N_908);
nor U7627 (N_7627,N_2061,N_292);
or U7628 (N_7628,N_4238,N_1991);
nand U7629 (N_7629,N_1521,N_292);
nand U7630 (N_7630,N_1366,N_462);
and U7631 (N_7631,N_4766,N_1009);
and U7632 (N_7632,N_3489,N_3849);
nor U7633 (N_7633,N_87,N_3989);
nand U7634 (N_7634,N_4189,N_1235);
and U7635 (N_7635,N_2336,N_3547);
nand U7636 (N_7636,N_1187,N_658);
and U7637 (N_7637,N_511,N_3538);
nand U7638 (N_7638,N_3390,N_1270);
or U7639 (N_7639,N_3213,N_370);
and U7640 (N_7640,N_2967,N_1109);
and U7641 (N_7641,N_2245,N_1181);
xnor U7642 (N_7642,N_2502,N_4926);
or U7643 (N_7643,N_4884,N_2502);
and U7644 (N_7644,N_2431,N_4268);
nand U7645 (N_7645,N_440,N_17);
or U7646 (N_7646,N_1282,N_261);
and U7647 (N_7647,N_4952,N_1075);
and U7648 (N_7648,N_4884,N_4408);
and U7649 (N_7649,N_220,N_726);
nand U7650 (N_7650,N_3602,N_2879);
nor U7651 (N_7651,N_578,N_2277);
nor U7652 (N_7652,N_3159,N_1229);
and U7653 (N_7653,N_3427,N_1629);
and U7654 (N_7654,N_4210,N_2683);
and U7655 (N_7655,N_741,N_4469);
nor U7656 (N_7656,N_1579,N_1091);
nand U7657 (N_7657,N_2344,N_3782);
and U7658 (N_7658,N_3034,N_754);
and U7659 (N_7659,N_4365,N_4499);
or U7660 (N_7660,N_2235,N_547);
and U7661 (N_7661,N_2657,N_989);
and U7662 (N_7662,N_3147,N_3675);
and U7663 (N_7663,N_1618,N_1694);
or U7664 (N_7664,N_4991,N_2661);
and U7665 (N_7665,N_4737,N_256);
or U7666 (N_7666,N_681,N_1226);
nand U7667 (N_7667,N_3838,N_1789);
and U7668 (N_7668,N_976,N_4701);
nand U7669 (N_7669,N_4382,N_4765);
and U7670 (N_7670,N_1579,N_2199);
nor U7671 (N_7671,N_4516,N_2343);
and U7672 (N_7672,N_4182,N_2297);
nor U7673 (N_7673,N_767,N_4709);
and U7674 (N_7674,N_3245,N_1320);
nand U7675 (N_7675,N_2997,N_2272);
or U7676 (N_7676,N_4372,N_2613);
nor U7677 (N_7677,N_112,N_1988);
or U7678 (N_7678,N_241,N_1433);
nor U7679 (N_7679,N_3416,N_3621);
nor U7680 (N_7680,N_3341,N_2947);
nand U7681 (N_7681,N_1770,N_2877);
nand U7682 (N_7682,N_4682,N_3071);
or U7683 (N_7683,N_4858,N_4621);
and U7684 (N_7684,N_829,N_2171);
nor U7685 (N_7685,N_2512,N_608);
nand U7686 (N_7686,N_2717,N_1321);
nor U7687 (N_7687,N_1134,N_1797);
or U7688 (N_7688,N_320,N_2708);
or U7689 (N_7689,N_3076,N_1070);
and U7690 (N_7690,N_2389,N_983);
nor U7691 (N_7691,N_100,N_4646);
or U7692 (N_7692,N_605,N_366);
nand U7693 (N_7693,N_3904,N_583);
and U7694 (N_7694,N_3500,N_360);
and U7695 (N_7695,N_2878,N_3870);
or U7696 (N_7696,N_573,N_906);
and U7697 (N_7697,N_847,N_1498);
and U7698 (N_7698,N_4662,N_2925);
or U7699 (N_7699,N_1339,N_3945);
nor U7700 (N_7700,N_3796,N_2752);
or U7701 (N_7701,N_3487,N_1077);
and U7702 (N_7702,N_1203,N_4726);
nand U7703 (N_7703,N_4508,N_2078);
nor U7704 (N_7704,N_2260,N_4447);
and U7705 (N_7705,N_4796,N_352);
or U7706 (N_7706,N_4567,N_1370);
and U7707 (N_7707,N_109,N_3320);
or U7708 (N_7708,N_2775,N_2057);
or U7709 (N_7709,N_4365,N_2235);
nor U7710 (N_7710,N_2290,N_4927);
and U7711 (N_7711,N_4797,N_4548);
and U7712 (N_7712,N_1003,N_2167);
nand U7713 (N_7713,N_4523,N_909);
nand U7714 (N_7714,N_1140,N_3693);
nor U7715 (N_7715,N_2604,N_1580);
nor U7716 (N_7716,N_3081,N_194);
or U7717 (N_7717,N_1315,N_1745);
or U7718 (N_7718,N_1094,N_3702);
nor U7719 (N_7719,N_4142,N_2699);
and U7720 (N_7720,N_1651,N_3189);
or U7721 (N_7721,N_3076,N_1183);
or U7722 (N_7722,N_4949,N_3936);
nor U7723 (N_7723,N_1533,N_2064);
nor U7724 (N_7724,N_3873,N_4602);
nand U7725 (N_7725,N_100,N_535);
or U7726 (N_7726,N_2950,N_2153);
nand U7727 (N_7727,N_3377,N_1453);
and U7728 (N_7728,N_1305,N_1508);
or U7729 (N_7729,N_2651,N_3437);
nor U7730 (N_7730,N_4327,N_4640);
and U7731 (N_7731,N_3456,N_4061);
nand U7732 (N_7732,N_1873,N_1097);
or U7733 (N_7733,N_4224,N_4367);
nand U7734 (N_7734,N_2559,N_104);
nor U7735 (N_7735,N_4562,N_806);
nand U7736 (N_7736,N_976,N_2406);
or U7737 (N_7737,N_233,N_3926);
nor U7738 (N_7738,N_4711,N_2240);
nand U7739 (N_7739,N_1856,N_1431);
or U7740 (N_7740,N_4598,N_1918);
and U7741 (N_7741,N_3498,N_4417);
or U7742 (N_7742,N_1310,N_4033);
and U7743 (N_7743,N_1043,N_1001);
nand U7744 (N_7744,N_4927,N_4074);
and U7745 (N_7745,N_484,N_4832);
xnor U7746 (N_7746,N_3000,N_529);
and U7747 (N_7747,N_262,N_330);
nand U7748 (N_7748,N_1546,N_2123);
and U7749 (N_7749,N_3234,N_1124);
and U7750 (N_7750,N_4424,N_2116);
and U7751 (N_7751,N_2171,N_1972);
and U7752 (N_7752,N_3244,N_2706);
nand U7753 (N_7753,N_3930,N_1125);
and U7754 (N_7754,N_4538,N_2548);
nand U7755 (N_7755,N_1700,N_2862);
nor U7756 (N_7756,N_1316,N_3616);
nor U7757 (N_7757,N_1048,N_3637);
and U7758 (N_7758,N_4613,N_2638);
or U7759 (N_7759,N_4991,N_2438);
nand U7760 (N_7760,N_3865,N_3570);
nor U7761 (N_7761,N_2073,N_690);
and U7762 (N_7762,N_3057,N_192);
nor U7763 (N_7763,N_1628,N_535);
nand U7764 (N_7764,N_1235,N_126);
or U7765 (N_7765,N_2290,N_4801);
nand U7766 (N_7766,N_172,N_4851);
or U7767 (N_7767,N_4923,N_1934);
and U7768 (N_7768,N_317,N_817);
or U7769 (N_7769,N_2048,N_4526);
nand U7770 (N_7770,N_1264,N_2627);
nand U7771 (N_7771,N_4449,N_1132);
and U7772 (N_7772,N_3547,N_2293);
or U7773 (N_7773,N_2370,N_4365);
and U7774 (N_7774,N_4896,N_238);
nand U7775 (N_7775,N_2649,N_4340);
nor U7776 (N_7776,N_4695,N_2645);
and U7777 (N_7777,N_4521,N_4404);
nand U7778 (N_7778,N_900,N_2523);
or U7779 (N_7779,N_634,N_1337);
and U7780 (N_7780,N_430,N_365);
nand U7781 (N_7781,N_3146,N_1743);
nor U7782 (N_7782,N_1890,N_3518);
and U7783 (N_7783,N_3161,N_4850);
and U7784 (N_7784,N_4607,N_1381);
nand U7785 (N_7785,N_1941,N_1497);
nand U7786 (N_7786,N_545,N_2977);
nand U7787 (N_7787,N_4948,N_1347);
nor U7788 (N_7788,N_4491,N_1933);
nand U7789 (N_7789,N_2362,N_2075);
nand U7790 (N_7790,N_559,N_4677);
and U7791 (N_7791,N_561,N_2972);
or U7792 (N_7792,N_1660,N_4727);
or U7793 (N_7793,N_4946,N_3918);
nor U7794 (N_7794,N_3400,N_3954);
and U7795 (N_7795,N_2152,N_358);
nor U7796 (N_7796,N_1548,N_2450);
and U7797 (N_7797,N_2614,N_1275);
nor U7798 (N_7798,N_2932,N_2241);
and U7799 (N_7799,N_2872,N_629);
or U7800 (N_7800,N_1235,N_2318);
nand U7801 (N_7801,N_1981,N_940);
nand U7802 (N_7802,N_471,N_239);
and U7803 (N_7803,N_351,N_2480);
and U7804 (N_7804,N_4033,N_3948);
nand U7805 (N_7805,N_4115,N_3771);
and U7806 (N_7806,N_3030,N_1253);
and U7807 (N_7807,N_278,N_2302);
nor U7808 (N_7808,N_2044,N_1684);
nor U7809 (N_7809,N_1736,N_3206);
nor U7810 (N_7810,N_4815,N_2315);
and U7811 (N_7811,N_4747,N_517);
and U7812 (N_7812,N_2542,N_162);
or U7813 (N_7813,N_2497,N_934);
or U7814 (N_7814,N_2228,N_2493);
or U7815 (N_7815,N_3917,N_158);
nand U7816 (N_7816,N_1473,N_3126);
and U7817 (N_7817,N_4828,N_2479);
and U7818 (N_7818,N_1766,N_433);
and U7819 (N_7819,N_129,N_3676);
and U7820 (N_7820,N_4742,N_1370);
and U7821 (N_7821,N_3292,N_2096);
or U7822 (N_7822,N_2382,N_3055);
or U7823 (N_7823,N_3102,N_766);
or U7824 (N_7824,N_311,N_2020);
or U7825 (N_7825,N_676,N_500);
or U7826 (N_7826,N_102,N_2374);
and U7827 (N_7827,N_1030,N_2720);
nor U7828 (N_7828,N_2652,N_2232);
or U7829 (N_7829,N_1565,N_3502);
and U7830 (N_7830,N_3966,N_4885);
nand U7831 (N_7831,N_255,N_3204);
or U7832 (N_7832,N_1644,N_4212);
nor U7833 (N_7833,N_2062,N_3899);
nand U7834 (N_7834,N_1342,N_3938);
nor U7835 (N_7835,N_2705,N_2952);
nand U7836 (N_7836,N_3164,N_1784);
or U7837 (N_7837,N_4523,N_3526);
nand U7838 (N_7838,N_4942,N_3363);
nand U7839 (N_7839,N_3425,N_4709);
nor U7840 (N_7840,N_3612,N_1955);
nand U7841 (N_7841,N_4046,N_3814);
nor U7842 (N_7842,N_480,N_4092);
nand U7843 (N_7843,N_2994,N_2175);
nor U7844 (N_7844,N_4489,N_807);
nand U7845 (N_7845,N_3812,N_3879);
or U7846 (N_7846,N_3907,N_2768);
nor U7847 (N_7847,N_1923,N_1025);
and U7848 (N_7848,N_2462,N_4418);
nor U7849 (N_7849,N_3609,N_1949);
nand U7850 (N_7850,N_3279,N_583);
nand U7851 (N_7851,N_3806,N_396);
or U7852 (N_7852,N_4406,N_4068);
or U7853 (N_7853,N_4521,N_4323);
or U7854 (N_7854,N_958,N_1050);
nor U7855 (N_7855,N_4356,N_581);
and U7856 (N_7856,N_426,N_4407);
nor U7857 (N_7857,N_4375,N_3017);
and U7858 (N_7858,N_367,N_3358);
or U7859 (N_7859,N_4381,N_3165);
nor U7860 (N_7860,N_1569,N_4023);
and U7861 (N_7861,N_1516,N_1119);
and U7862 (N_7862,N_293,N_2896);
nor U7863 (N_7863,N_752,N_4802);
nand U7864 (N_7864,N_1172,N_300);
nand U7865 (N_7865,N_3680,N_89);
and U7866 (N_7866,N_2989,N_1328);
nand U7867 (N_7867,N_3289,N_2429);
nor U7868 (N_7868,N_537,N_19);
nor U7869 (N_7869,N_3000,N_3304);
or U7870 (N_7870,N_3244,N_1775);
and U7871 (N_7871,N_4846,N_1237);
or U7872 (N_7872,N_4661,N_3563);
nor U7873 (N_7873,N_2003,N_3234);
or U7874 (N_7874,N_1658,N_1656);
nand U7875 (N_7875,N_4605,N_108);
nand U7876 (N_7876,N_1413,N_3652);
or U7877 (N_7877,N_4903,N_539);
or U7878 (N_7878,N_3177,N_4870);
and U7879 (N_7879,N_3762,N_273);
xor U7880 (N_7880,N_4176,N_4926);
nor U7881 (N_7881,N_1165,N_4208);
nor U7882 (N_7882,N_3804,N_264);
nor U7883 (N_7883,N_1532,N_596);
nor U7884 (N_7884,N_3863,N_3456);
and U7885 (N_7885,N_4565,N_1473);
nor U7886 (N_7886,N_1114,N_3836);
and U7887 (N_7887,N_176,N_787);
nor U7888 (N_7888,N_3407,N_4733);
or U7889 (N_7889,N_1589,N_258);
or U7890 (N_7890,N_2073,N_1507);
nor U7891 (N_7891,N_1251,N_433);
or U7892 (N_7892,N_1040,N_753);
nand U7893 (N_7893,N_4152,N_4114);
xor U7894 (N_7894,N_298,N_1861);
nor U7895 (N_7895,N_2856,N_4395);
nor U7896 (N_7896,N_980,N_2195);
and U7897 (N_7897,N_4266,N_2163);
nor U7898 (N_7898,N_421,N_3020);
nor U7899 (N_7899,N_2601,N_310);
or U7900 (N_7900,N_3663,N_373);
or U7901 (N_7901,N_4004,N_3475);
nor U7902 (N_7902,N_3385,N_978);
and U7903 (N_7903,N_4204,N_3350);
or U7904 (N_7904,N_2556,N_4212);
or U7905 (N_7905,N_3014,N_4583);
and U7906 (N_7906,N_3646,N_1083);
or U7907 (N_7907,N_249,N_1681);
nand U7908 (N_7908,N_58,N_1467);
or U7909 (N_7909,N_1628,N_4793);
nor U7910 (N_7910,N_4223,N_3187);
nand U7911 (N_7911,N_4211,N_2536);
or U7912 (N_7912,N_2077,N_2181);
nand U7913 (N_7913,N_3598,N_166);
nor U7914 (N_7914,N_4173,N_2300);
nand U7915 (N_7915,N_4073,N_2996);
or U7916 (N_7916,N_3704,N_3801);
and U7917 (N_7917,N_1396,N_2387);
or U7918 (N_7918,N_1952,N_4146);
nand U7919 (N_7919,N_3714,N_1625);
or U7920 (N_7920,N_411,N_315);
or U7921 (N_7921,N_4757,N_2710);
nand U7922 (N_7922,N_4965,N_847);
nand U7923 (N_7923,N_231,N_2087);
nand U7924 (N_7924,N_4462,N_2496);
nand U7925 (N_7925,N_1260,N_3224);
or U7926 (N_7926,N_3043,N_1224);
nand U7927 (N_7927,N_1831,N_1809);
nor U7928 (N_7928,N_30,N_2311);
nand U7929 (N_7929,N_3034,N_3148);
nand U7930 (N_7930,N_3845,N_1194);
nand U7931 (N_7931,N_3800,N_2051);
nand U7932 (N_7932,N_1049,N_4499);
nand U7933 (N_7933,N_4680,N_799);
nand U7934 (N_7934,N_927,N_262);
or U7935 (N_7935,N_3709,N_1002);
nor U7936 (N_7936,N_1573,N_4430);
nor U7937 (N_7937,N_233,N_1050);
and U7938 (N_7938,N_3624,N_3642);
nor U7939 (N_7939,N_4927,N_1595);
xor U7940 (N_7940,N_4316,N_369);
or U7941 (N_7941,N_4533,N_4381);
or U7942 (N_7942,N_4686,N_4797);
nor U7943 (N_7943,N_3526,N_4917);
or U7944 (N_7944,N_4863,N_3696);
or U7945 (N_7945,N_2339,N_3725);
nor U7946 (N_7946,N_2826,N_2604);
nor U7947 (N_7947,N_2169,N_1692);
and U7948 (N_7948,N_890,N_1472);
or U7949 (N_7949,N_4665,N_11);
nor U7950 (N_7950,N_4981,N_4837);
or U7951 (N_7951,N_3998,N_2663);
nand U7952 (N_7952,N_3742,N_187);
nand U7953 (N_7953,N_1565,N_3615);
and U7954 (N_7954,N_753,N_618);
or U7955 (N_7955,N_3579,N_4472);
and U7956 (N_7956,N_3826,N_1839);
nand U7957 (N_7957,N_4794,N_2196);
and U7958 (N_7958,N_1592,N_1364);
or U7959 (N_7959,N_2112,N_1435);
nor U7960 (N_7960,N_352,N_2823);
and U7961 (N_7961,N_2863,N_3888);
or U7962 (N_7962,N_3331,N_3222);
nor U7963 (N_7963,N_4124,N_1271);
and U7964 (N_7964,N_337,N_145);
or U7965 (N_7965,N_2060,N_3689);
nor U7966 (N_7966,N_4328,N_343);
nor U7967 (N_7967,N_3305,N_4395);
nor U7968 (N_7968,N_2383,N_4975);
and U7969 (N_7969,N_4946,N_4895);
nand U7970 (N_7970,N_1863,N_1992);
and U7971 (N_7971,N_3431,N_1916);
or U7972 (N_7972,N_1878,N_4287);
nand U7973 (N_7973,N_1816,N_1656);
nor U7974 (N_7974,N_2859,N_3047);
or U7975 (N_7975,N_255,N_2138);
nand U7976 (N_7976,N_2952,N_2939);
xnor U7977 (N_7977,N_3823,N_1318);
nor U7978 (N_7978,N_890,N_1959);
nor U7979 (N_7979,N_4171,N_4751);
or U7980 (N_7980,N_896,N_998);
nor U7981 (N_7981,N_4106,N_1128);
and U7982 (N_7982,N_3751,N_2367);
nor U7983 (N_7983,N_3303,N_2238);
nor U7984 (N_7984,N_2699,N_2761);
nand U7985 (N_7985,N_4297,N_3604);
and U7986 (N_7986,N_3099,N_2119);
or U7987 (N_7987,N_4734,N_430);
nor U7988 (N_7988,N_3939,N_2714);
or U7989 (N_7989,N_3289,N_1769);
and U7990 (N_7990,N_463,N_3631);
nor U7991 (N_7991,N_4019,N_1677);
and U7992 (N_7992,N_2808,N_3576);
or U7993 (N_7993,N_2811,N_750);
or U7994 (N_7994,N_3678,N_381);
nor U7995 (N_7995,N_1911,N_685);
and U7996 (N_7996,N_1941,N_3181);
nor U7997 (N_7997,N_596,N_3495);
nand U7998 (N_7998,N_1733,N_1411);
xor U7999 (N_7999,N_2962,N_199);
or U8000 (N_8000,N_1923,N_3652);
xnor U8001 (N_8001,N_745,N_920);
and U8002 (N_8002,N_2045,N_563);
nand U8003 (N_8003,N_2417,N_2122);
xnor U8004 (N_8004,N_1871,N_4246);
or U8005 (N_8005,N_648,N_1718);
nor U8006 (N_8006,N_2679,N_4409);
or U8007 (N_8007,N_2055,N_2028);
or U8008 (N_8008,N_4836,N_3817);
and U8009 (N_8009,N_1887,N_213);
nand U8010 (N_8010,N_846,N_59);
nand U8011 (N_8011,N_3980,N_4101);
nor U8012 (N_8012,N_4925,N_1296);
nor U8013 (N_8013,N_485,N_4468);
nor U8014 (N_8014,N_4117,N_1862);
or U8015 (N_8015,N_974,N_716);
or U8016 (N_8016,N_1500,N_2962);
and U8017 (N_8017,N_2382,N_869);
or U8018 (N_8018,N_2888,N_2898);
or U8019 (N_8019,N_1021,N_2207);
and U8020 (N_8020,N_3808,N_9);
or U8021 (N_8021,N_511,N_3632);
or U8022 (N_8022,N_67,N_4521);
or U8023 (N_8023,N_4622,N_3458);
or U8024 (N_8024,N_1227,N_831);
nand U8025 (N_8025,N_3433,N_1545);
and U8026 (N_8026,N_1884,N_3823);
or U8027 (N_8027,N_3738,N_2211);
or U8028 (N_8028,N_4192,N_2426);
nor U8029 (N_8029,N_2756,N_2280);
nand U8030 (N_8030,N_2605,N_850);
nor U8031 (N_8031,N_206,N_441);
and U8032 (N_8032,N_3637,N_349);
nor U8033 (N_8033,N_1282,N_616);
and U8034 (N_8034,N_2155,N_1225);
or U8035 (N_8035,N_3634,N_2028);
or U8036 (N_8036,N_3337,N_4839);
nor U8037 (N_8037,N_2878,N_3309);
nor U8038 (N_8038,N_2335,N_326);
and U8039 (N_8039,N_4838,N_309);
nor U8040 (N_8040,N_101,N_2199);
xnor U8041 (N_8041,N_1163,N_149);
nor U8042 (N_8042,N_909,N_151);
or U8043 (N_8043,N_1603,N_1821);
or U8044 (N_8044,N_3654,N_596);
or U8045 (N_8045,N_842,N_1445);
or U8046 (N_8046,N_3787,N_3872);
nor U8047 (N_8047,N_2332,N_2997);
or U8048 (N_8048,N_1947,N_1467);
nor U8049 (N_8049,N_137,N_4951);
and U8050 (N_8050,N_4385,N_3562);
nor U8051 (N_8051,N_1862,N_3576);
or U8052 (N_8052,N_3353,N_2957);
and U8053 (N_8053,N_1898,N_4134);
or U8054 (N_8054,N_3484,N_4783);
and U8055 (N_8055,N_2428,N_5);
or U8056 (N_8056,N_4,N_2934);
nand U8057 (N_8057,N_4802,N_4027);
or U8058 (N_8058,N_3579,N_4146);
and U8059 (N_8059,N_324,N_1044);
or U8060 (N_8060,N_4650,N_921);
nor U8061 (N_8061,N_971,N_1777);
nor U8062 (N_8062,N_4225,N_812);
nand U8063 (N_8063,N_2647,N_3970);
or U8064 (N_8064,N_1636,N_258);
and U8065 (N_8065,N_840,N_4375);
nor U8066 (N_8066,N_4734,N_2847);
nor U8067 (N_8067,N_4576,N_4297);
nor U8068 (N_8068,N_509,N_2880);
and U8069 (N_8069,N_3005,N_4704);
and U8070 (N_8070,N_1344,N_524);
or U8071 (N_8071,N_354,N_2868);
nand U8072 (N_8072,N_165,N_2558);
nor U8073 (N_8073,N_1883,N_3048);
nor U8074 (N_8074,N_4597,N_3989);
nand U8075 (N_8075,N_2180,N_1677);
nand U8076 (N_8076,N_2795,N_1894);
nand U8077 (N_8077,N_1646,N_1928);
or U8078 (N_8078,N_4616,N_3511);
nand U8079 (N_8079,N_4351,N_1244);
nor U8080 (N_8080,N_2908,N_577);
or U8081 (N_8081,N_3760,N_530);
nand U8082 (N_8082,N_4853,N_4174);
and U8083 (N_8083,N_1429,N_4850);
or U8084 (N_8084,N_1104,N_274);
nor U8085 (N_8085,N_3630,N_90);
nor U8086 (N_8086,N_4403,N_3801);
and U8087 (N_8087,N_3302,N_3416);
or U8088 (N_8088,N_2589,N_2088);
and U8089 (N_8089,N_2790,N_980);
nor U8090 (N_8090,N_4914,N_3284);
or U8091 (N_8091,N_312,N_2101);
or U8092 (N_8092,N_1844,N_2239);
nand U8093 (N_8093,N_3312,N_3881);
and U8094 (N_8094,N_1791,N_2342);
nor U8095 (N_8095,N_120,N_2143);
or U8096 (N_8096,N_4793,N_4877);
or U8097 (N_8097,N_3144,N_345);
nand U8098 (N_8098,N_3659,N_211);
nor U8099 (N_8099,N_2096,N_4673);
and U8100 (N_8100,N_4455,N_849);
or U8101 (N_8101,N_588,N_3109);
nand U8102 (N_8102,N_4241,N_4248);
or U8103 (N_8103,N_4497,N_1015);
nand U8104 (N_8104,N_3470,N_4864);
xor U8105 (N_8105,N_3485,N_4252);
nand U8106 (N_8106,N_2031,N_2534);
nand U8107 (N_8107,N_1546,N_4211);
nor U8108 (N_8108,N_546,N_3309);
or U8109 (N_8109,N_4348,N_947);
or U8110 (N_8110,N_2337,N_2004);
nor U8111 (N_8111,N_1678,N_2859);
or U8112 (N_8112,N_3989,N_4103);
nor U8113 (N_8113,N_467,N_1810);
nand U8114 (N_8114,N_3945,N_4475);
nand U8115 (N_8115,N_3695,N_541);
or U8116 (N_8116,N_1232,N_2562);
and U8117 (N_8117,N_2516,N_3753);
or U8118 (N_8118,N_4708,N_2400);
and U8119 (N_8119,N_2822,N_4731);
or U8120 (N_8120,N_4789,N_3845);
and U8121 (N_8121,N_2949,N_1906);
or U8122 (N_8122,N_2540,N_3217);
and U8123 (N_8123,N_1813,N_1801);
nor U8124 (N_8124,N_1633,N_4801);
and U8125 (N_8125,N_3922,N_2496);
or U8126 (N_8126,N_4954,N_723);
and U8127 (N_8127,N_624,N_820);
or U8128 (N_8128,N_3573,N_3038);
and U8129 (N_8129,N_1904,N_3353);
and U8130 (N_8130,N_241,N_2341);
nand U8131 (N_8131,N_4795,N_2132);
nand U8132 (N_8132,N_359,N_1116);
nand U8133 (N_8133,N_2780,N_1955);
nand U8134 (N_8134,N_4681,N_2672);
nor U8135 (N_8135,N_2198,N_368);
and U8136 (N_8136,N_397,N_1830);
nand U8137 (N_8137,N_1615,N_1806);
and U8138 (N_8138,N_4149,N_1833);
and U8139 (N_8139,N_417,N_4046);
nand U8140 (N_8140,N_3810,N_373);
or U8141 (N_8141,N_4850,N_1257);
and U8142 (N_8142,N_2668,N_3916);
or U8143 (N_8143,N_1123,N_2471);
nand U8144 (N_8144,N_713,N_155);
nand U8145 (N_8145,N_2870,N_3286);
nand U8146 (N_8146,N_3902,N_4889);
and U8147 (N_8147,N_4453,N_818);
and U8148 (N_8148,N_2119,N_4088);
nor U8149 (N_8149,N_3202,N_518);
or U8150 (N_8150,N_1061,N_1227);
nand U8151 (N_8151,N_2379,N_2629);
nor U8152 (N_8152,N_570,N_4896);
xnor U8153 (N_8153,N_1968,N_1112);
and U8154 (N_8154,N_2676,N_3995);
and U8155 (N_8155,N_3543,N_1424);
nand U8156 (N_8156,N_1101,N_2301);
and U8157 (N_8157,N_635,N_4332);
or U8158 (N_8158,N_2044,N_1892);
or U8159 (N_8159,N_2037,N_4526);
nand U8160 (N_8160,N_926,N_4758);
nor U8161 (N_8161,N_2652,N_1963);
nor U8162 (N_8162,N_3908,N_563);
xnor U8163 (N_8163,N_131,N_3689);
nand U8164 (N_8164,N_118,N_2655);
and U8165 (N_8165,N_685,N_1280);
nor U8166 (N_8166,N_1403,N_413);
and U8167 (N_8167,N_3264,N_3949);
nor U8168 (N_8168,N_1573,N_1014);
nor U8169 (N_8169,N_1643,N_3074);
and U8170 (N_8170,N_2759,N_1202);
nand U8171 (N_8171,N_4336,N_1350);
nand U8172 (N_8172,N_1244,N_1068);
and U8173 (N_8173,N_4574,N_2690);
xnor U8174 (N_8174,N_2162,N_1268);
nand U8175 (N_8175,N_2500,N_4656);
nor U8176 (N_8176,N_3380,N_2684);
nand U8177 (N_8177,N_351,N_2591);
and U8178 (N_8178,N_919,N_1515);
or U8179 (N_8179,N_2904,N_25);
nand U8180 (N_8180,N_4143,N_1667);
and U8181 (N_8181,N_1387,N_908);
or U8182 (N_8182,N_3108,N_2402);
and U8183 (N_8183,N_1166,N_2442);
or U8184 (N_8184,N_1026,N_1402);
nand U8185 (N_8185,N_2456,N_1983);
nor U8186 (N_8186,N_3388,N_2833);
nand U8187 (N_8187,N_4010,N_4634);
or U8188 (N_8188,N_2891,N_1978);
or U8189 (N_8189,N_4582,N_543);
or U8190 (N_8190,N_3284,N_340);
nand U8191 (N_8191,N_4847,N_245);
and U8192 (N_8192,N_3270,N_3188);
nor U8193 (N_8193,N_2442,N_3389);
or U8194 (N_8194,N_3941,N_2842);
or U8195 (N_8195,N_2703,N_4125);
nand U8196 (N_8196,N_1404,N_4704);
or U8197 (N_8197,N_2256,N_4822);
nor U8198 (N_8198,N_3712,N_667);
nor U8199 (N_8199,N_1518,N_573);
and U8200 (N_8200,N_4752,N_1750);
and U8201 (N_8201,N_668,N_2170);
nand U8202 (N_8202,N_3800,N_3658);
and U8203 (N_8203,N_2722,N_2120);
or U8204 (N_8204,N_3968,N_4582);
or U8205 (N_8205,N_679,N_1061);
or U8206 (N_8206,N_1042,N_4695);
nand U8207 (N_8207,N_1393,N_3952);
and U8208 (N_8208,N_2327,N_4247);
nand U8209 (N_8209,N_1708,N_624);
nor U8210 (N_8210,N_313,N_3159);
nand U8211 (N_8211,N_2529,N_3997);
nor U8212 (N_8212,N_4664,N_3469);
nor U8213 (N_8213,N_807,N_2338);
nand U8214 (N_8214,N_2143,N_3822);
or U8215 (N_8215,N_1497,N_3965);
nand U8216 (N_8216,N_1479,N_2207);
and U8217 (N_8217,N_1020,N_2392);
or U8218 (N_8218,N_3945,N_87);
and U8219 (N_8219,N_4609,N_3435);
and U8220 (N_8220,N_1795,N_3160);
nand U8221 (N_8221,N_1276,N_1273);
and U8222 (N_8222,N_550,N_1548);
or U8223 (N_8223,N_1917,N_2322);
nor U8224 (N_8224,N_1680,N_212);
or U8225 (N_8225,N_1196,N_3196);
nor U8226 (N_8226,N_3843,N_789);
or U8227 (N_8227,N_1401,N_4184);
or U8228 (N_8228,N_878,N_779);
nand U8229 (N_8229,N_2824,N_3857);
nand U8230 (N_8230,N_2907,N_3235);
or U8231 (N_8231,N_2589,N_1991);
nand U8232 (N_8232,N_3316,N_4976);
and U8233 (N_8233,N_71,N_101);
nor U8234 (N_8234,N_4595,N_3029);
and U8235 (N_8235,N_297,N_4912);
xor U8236 (N_8236,N_4359,N_199);
nand U8237 (N_8237,N_6,N_698);
and U8238 (N_8238,N_419,N_247);
nor U8239 (N_8239,N_70,N_3315);
nor U8240 (N_8240,N_4452,N_4148);
nor U8241 (N_8241,N_3188,N_3724);
nor U8242 (N_8242,N_30,N_4416);
or U8243 (N_8243,N_4665,N_4909);
nand U8244 (N_8244,N_1003,N_2860);
and U8245 (N_8245,N_3521,N_525);
or U8246 (N_8246,N_3253,N_1417);
or U8247 (N_8247,N_4648,N_1932);
and U8248 (N_8248,N_305,N_3679);
nor U8249 (N_8249,N_3213,N_462);
nor U8250 (N_8250,N_4191,N_2447);
and U8251 (N_8251,N_4579,N_578);
nand U8252 (N_8252,N_2672,N_92);
and U8253 (N_8253,N_2159,N_2009);
or U8254 (N_8254,N_1631,N_1996);
and U8255 (N_8255,N_3335,N_919);
nor U8256 (N_8256,N_1159,N_3109);
and U8257 (N_8257,N_4511,N_1917);
and U8258 (N_8258,N_431,N_4557);
and U8259 (N_8259,N_2415,N_1322);
nand U8260 (N_8260,N_1390,N_1585);
or U8261 (N_8261,N_2233,N_130);
nand U8262 (N_8262,N_3320,N_4646);
nor U8263 (N_8263,N_383,N_3544);
and U8264 (N_8264,N_1200,N_2138);
or U8265 (N_8265,N_1133,N_1375);
nand U8266 (N_8266,N_2766,N_2371);
or U8267 (N_8267,N_1671,N_3106);
or U8268 (N_8268,N_1545,N_1352);
or U8269 (N_8269,N_1769,N_1153);
and U8270 (N_8270,N_40,N_3630);
and U8271 (N_8271,N_3902,N_634);
nand U8272 (N_8272,N_1006,N_544);
nor U8273 (N_8273,N_4666,N_611);
nor U8274 (N_8274,N_2884,N_1206);
and U8275 (N_8275,N_3627,N_1027);
nor U8276 (N_8276,N_1313,N_4742);
nor U8277 (N_8277,N_1025,N_4760);
nand U8278 (N_8278,N_1307,N_2384);
or U8279 (N_8279,N_3492,N_3792);
nand U8280 (N_8280,N_3260,N_3928);
nor U8281 (N_8281,N_2720,N_673);
nand U8282 (N_8282,N_792,N_2171);
nand U8283 (N_8283,N_3293,N_95);
or U8284 (N_8284,N_3599,N_678);
nor U8285 (N_8285,N_3380,N_2140);
nand U8286 (N_8286,N_2214,N_4112);
nand U8287 (N_8287,N_239,N_3009);
xnor U8288 (N_8288,N_2050,N_1387);
and U8289 (N_8289,N_4472,N_2521);
and U8290 (N_8290,N_1019,N_4622);
nor U8291 (N_8291,N_2340,N_2686);
nand U8292 (N_8292,N_145,N_4046);
nor U8293 (N_8293,N_2304,N_3528);
or U8294 (N_8294,N_20,N_1406);
or U8295 (N_8295,N_549,N_4174);
and U8296 (N_8296,N_3303,N_3498);
or U8297 (N_8297,N_3441,N_2695);
nor U8298 (N_8298,N_4589,N_4087);
and U8299 (N_8299,N_2546,N_3061);
and U8300 (N_8300,N_1007,N_1739);
nor U8301 (N_8301,N_4241,N_1643);
nand U8302 (N_8302,N_2306,N_4362);
nand U8303 (N_8303,N_220,N_3288);
and U8304 (N_8304,N_1463,N_831);
nor U8305 (N_8305,N_356,N_3845);
nand U8306 (N_8306,N_2521,N_535);
and U8307 (N_8307,N_2422,N_1401);
nor U8308 (N_8308,N_2368,N_4229);
nand U8309 (N_8309,N_3949,N_354);
and U8310 (N_8310,N_4824,N_2479);
nor U8311 (N_8311,N_3162,N_3400);
nor U8312 (N_8312,N_3466,N_605);
nor U8313 (N_8313,N_210,N_4376);
or U8314 (N_8314,N_807,N_145);
and U8315 (N_8315,N_146,N_2342);
nor U8316 (N_8316,N_1964,N_2856);
or U8317 (N_8317,N_3727,N_2515);
or U8318 (N_8318,N_4632,N_1014);
and U8319 (N_8319,N_3114,N_2060);
nor U8320 (N_8320,N_2689,N_4841);
nor U8321 (N_8321,N_1967,N_1324);
nand U8322 (N_8322,N_1079,N_2039);
xnor U8323 (N_8323,N_2433,N_3456);
or U8324 (N_8324,N_3220,N_4246);
and U8325 (N_8325,N_2350,N_3794);
and U8326 (N_8326,N_2542,N_3288);
nand U8327 (N_8327,N_2639,N_344);
or U8328 (N_8328,N_1635,N_2553);
or U8329 (N_8329,N_3083,N_4745);
nor U8330 (N_8330,N_640,N_385);
and U8331 (N_8331,N_3236,N_1657);
nand U8332 (N_8332,N_4831,N_538);
nand U8333 (N_8333,N_1190,N_4449);
nand U8334 (N_8334,N_4826,N_2455);
or U8335 (N_8335,N_2416,N_129);
or U8336 (N_8336,N_2837,N_365);
and U8337 (N_8337,N_3271,N_2373);
or U8338 (N_8338,N_4288,N_1485);
nand U8339 (N_8339,N_40,N_3365);
or U8340 (N_8340,N_3625,N_3502);
nor U8341 (N_8341,N_928,N_1466);
or U8342 (N_8342,N_4381,N_4072);
or U8343 (N_8343,N_547,N_3097);
nand U8344 (N_8344,N_3407,N_4016);
nand U8345 (N_8345,N_1584,N_2515);
and U8346 (N_8346,N_4068,N_1785);
nor U8347 (N_8347,N_2689,N_2889);
or U8348 (N_8348,N_4794,N_160);
nand U8349 (N_8349,N_4557,N_3603);
nor U8350 (N_8350,N_1621,N_2733);
and U8351 (N_8351,N_2132,N_2265);
and U8352 (N_8352,N_2447,N_1659);
and U8353 (N_8353,N_1952,N_3831);
nor U8354 (N_8354,N_4562,N_4591);
or U8355 (N_8355,N_4118,N_1436);
and U8356 (N_8356,N_3872,N_4766);
and U8357 (N_8357,N_2499,N_2232);
and U8358 (N_8358,N_3427,N_218);
and U8359 (N_8359,N_1967,N_2992);
nor U8360 (N_8360,N_3620,N_2229);
or U8361 (N_8361,N_1220,N_219);
nor U8362 (N_8362,N_4884,N_4596);
nand U8363 (N_8363,N_2058,N_3356);
nand U8364 (N_8364,N_3404,N_3955);
and U8365 (N_8365,N_998,N_360);
nor U8366 (N_8366,N_4217,N_1829);
nand U8367 (N_8367,N_280,N_3477);
and U8368 (N_8368,N_4336,N_2217);
xor U8369 (N_8369,N_3107,N_4401);
nor U8370 (N_8370,N_937,N_3441);
or U8371 (N_8371,N_4384,N_4003);
nor U8372 (N_8372,N_2380,N_3162);
and U8373 (N_8373,N_721,N_777);
and U8374 (N_8374,N_2985,N_1807);
nand U8375 (N_8375,N_3162,N_2576);
and U8376 (N_8376,N_455,N_7);
and U8377 (N_8377,N_3359,N_1368);
nor U8378 (N_8378,N_4436,N_4050);
and U8379 (N_8379,N_4381,N_1218);
and U8380 (N_8380,N_4206,N_1201);
and U8381 (N_8381,N_2581,N_1837);
nand U8382 (N_8382,N_1387,N_792);
or U8383 (N_8383,N_2756,N_1848);
and U8384 (N_8384,N_569,N_2241);
nand U8385 (N_8385,N_1201,N_3379);
nand U8386 (N_8386,N_3292,N_1157);
and U8387 (N_8387,N_2217,N_1720);
and U8388 (N_8388,N_1343,N_4459);
or U8389 (N_8389,N_548,N_4592);
or U8390 (N_8390,N_3726,N_2531);
nand U8391 (N_8391,N_3459,N_232);
nor U8392 (N_8392,N_3387,N_2193);
nor U8393 (N_8393,N_826,N_81);
nor U8394 (N_8394,N_3868,N_3837);
or U8395 (N_8395,N_933,N_3575);
and U8396 (N_8396,N_1970,N_3947);
and U8397 (N_8397,N_4157,N_320);
and U8398 (N_8398,N_2306,N_3563);
and U8399 (N_8399,N_4681,N_3728);
nor U8400 (N_8400,N_1150,N_2733);
or U8401 (N_8401,N_594,N_4789);
nor U8402 (N_8402,N_1884,N_1866);
and U8403 (N_8403,N_3757,N_4000);
nand U8404 (N_8404,N_1447,N_551);
nor U8405 (N_8405,N_2146,N_2354);
nand U8406 (N_8406,N_1641,N_1381);
or U8407 (N_8407,N_393,N_3437);
xnor U8408 (N_8408,N_4410,N_2262);
and U8409 (N_8409,N_760,N_556);
nand U8410 (N_8410,N_4177,N_3587);
nor U8411 (N_8411,N_678,N_3282);
nand U8412 (N_8412,N_2198,N_1522);
xor U8413 (N_8413,N_4835,N_1376);
nand U8414 (N_8414,N_389,N_1442);
or U8415 (N_8415,N_2259,N_4559);
nand U8416 (N_8416,N_335,N_3353);
nor U8417 (N_8417,N_2713,N_3528);
or U8418 (N_8418,N_4059,N_3980);
and U8419 (N_8419,N_4062,N_2875);
and U8420 (N_8420,N_4697,N_2483);
or U8421 (N_8421,N_2398,N_3124);
or U8422 (N_8422,N_2802,N_1423);
and U8423 (N_8423,N_1747,N_2427);
and U8424 (N_8424,N_2229,N_600);
or U8425 (N_8425,N_835,N_823);
nor U8426 (N_8426,N_2975,N_1454);
and U8427 (N_8427,N_2749,N_3478);
and U8428 (N_8428,N_4049,N_3514);
and U8429 (N_8429,N_3766,N_1577);
nand U8430 (N_8430,N_852,N_3111);
nor U8431 (N_8431,N_2991,N_1716);
nand U8432 (N_8432,N_2495,N_1837);
or U8433 (N_8433,N_3174,N_4345);
and U8434 (N_8434,N_4368,N_3539);
or U8435 (N_8435,N_4978,N_4571);
or U8436 (N_8436,N_1577,N_4892);
nor U8437 (N_8437,N_2384,N_1900);
xor U8438 (N_8438,N_3630,N_3467);
nand U8439 (N_8439,N_2938,N_1247);
or U8440 (N_8440,N_963,N_2766);
and U8441 (N_8441,N_838,N_1317);
nor U8442 (N_8442,N_1046,N_2633);
or U8443 (N_8443,N_154,N_1635);
or U8444 (N_8444,N_1892,N_821);
or U8445 (N_8445,N_3702,N_3760);
nor U8446 (N_8446,N_351,N_2572);
nor U8447 (N_8447,N_4111,N_1346);
nand U8448 (N_8448,N_4352,N_4092);
and U8449 (N_8449,N_2251,N_137);
nor U8450 (N_8450,N_1380,N_2501);
and U8451 (N_8451,N_3519,N_1313);
nor U8452 (N_8452,N_421,N_2937);
or U8453 (N_8453,N_3647,N_3105);
nand U8454 (N_8454,N_2137,N_3850);
nand U8455 (N_8455,N_1783,N_1675);
nand U8456 (N_8456,N_2122,N_1898);
nand U8457 (N_8457,N_2026,N_1793);
and U8458 (N_8458,N_1872,N_4233);
or U8459 (N_8459,N_656,N_4787);
nand U8460 (N_8460,N_2163,N_3085);
or U8461 (N_8461,N_2004,N_3952);
nor U8462 (N_8462,N_3086,N_1038);
or U8463 (N_8463,N_3898,N_2625);
nor U8464 (N_8464,N_356,N_551);
or U8465 (N_8465,N_2465,N_4558);
or U8466 (N_8466,N_3379,N_1520);
and U8467 (N_8467,N_1219,N_743);
and U8468 (N_8468,N_3938,N_1222);
nand U8469 (N_8469,N_3786,N_1826);
or U8470 (N_8470,N_446,N_623);
and U8471 (N_8471,N_1139,N_1192);
or U8472 (N_8472,N_4286,N_3151);
nand U8473 (N_8473,N_1753,N_3767);
and U8474 (N_8474,N_17,N_95);
nor U8475 (N_8475,N_3037,N_3222);
nor U8476 (N_8476,N_2423,N_3908);
and U8477 (N_8477,N_3939,N_1107);
or U8478 (N_8478,N_4311,N_3626);
and U8479 (N_8479,N_2486,N_1463);
and U8480 (N_8480,N_1171,N_2751);
and U8481 (N_8481,N_2241,N_4430);
xnor U8482 (N_8482,N_252,N_260);
nand U8483 (N_8483,N_4755,N_2342);
or U8484 (N_8484,N_3127,N_4245);
and U8485 (N_8485,N_3119,N_3619);
nor U8486 (N_8486,N_4857,N_3016);
nor U8487 (N_8487,N_2803,N_1479);
or U8488 (N_8488,N_4108,N_4610);
and U8489 (N_8489,N_4182,N_4197);
xor U8490 (N_8490,N_2467,N_351);
nand U8491 (N_8491,N_2725,N_149);
and U8492 (N_8492,N_993,N_1317);
and U8493 (N_8493,N_2463,N_2125);
nor U8494 (N_8494,N_1768,N_1729);
nand U8495 (N_8495,N_2902,N_4699);
nand U8496 (N_8496,N_299,N_3821);
nand U8497 (N_8497,N_95,N_2540);
and U8498 (N_8498,N_2008,N_2349);
and U8499 (N_8499,N_1722,N_2133);
nand U8500 (N_8500,N_697,N_4314);
or U8501 (N_8501,N_831,N_1785);
or U8502 (N_8502,N_4419,N_4907);
nand U8503 (N_8503,N_3982,N_3203);
or U8504 (N_8504,N_1637,N_475);
nor U8505 (N_8505,N_504,N_748);
or U8506 (N_8506,N_652,N_419);
nor U8507 (N_8507,N_4953,N_4203);
nand U8508 (N_8508,N_2876,N_207);
and U8509 (N_8509,N_3162,N_239);
or U8510 (N_8510,N_4387,N_127);
or U8511 (N_8511,N_2205,N_1609);
nor U8512 (N_8512,N_3740,N_4065);
nand U8513 (N_8513,N_2499,N_976);
or U8514 (N_8514,N_1626,N_321);
or U8515 (N_8515,N_2140,N_40);
nand U8516 (N_8516,N_3424,N_3214);
or U8517 (N_8517,N_501,N_458);
and U8518 (N_8518,N_116,N_1411);
or U8519 (N_8519,N_603,N_687);
nand U8520 (N_8520,N_3005,N_3653);
nand U8521 (N_8521,N_430,N_2527);
nand U8522 (N_8522,N_3376,N_1780);
or U8523 (N_8523,N_634,N_3763);
or U8524 (N_8524,N_3071,N_2706);
and U8525 (N_8525,N_1754,N_587);
nand U8526 (N_8526,N_3218,N_4437);
nor U8527 (N_8527,N_1656,N_1467);
nand U8528 (N_8528,N_2398,N_1992);
and U8529 (N_8529,N_1719,N_239);
and U8530 (N_8530,N_3560,N_266);
or U8531 (N_8531,N_3554,N_3656);
and U8532 (N_8532,N_2096,N_1549);
and U8533 (N_8533,N_719,N_2539);
or U8534 (N_8534,N_1993,N_3555);
and U8535 (N_8535,N_638,N_2768);
or U8536 (N_8536,N_2205,N_1342);
or U8537 (N_8537,N_3714,N_2765);
or U8538 (N_8538,N_410,N_3144);
and U8539 (N_8539,N_3263,N_3296);
and U8540 (N_8540,N_832,N_4563);
nand U8541 (N_8541,N_2277,N_1241);
nor U8542 (N_8542,N_2618,N_4400);
and U8543 (N_8543,N_3984,N_499);
nand U8544 (N_8544,N_1114,N_4698);
nor U8545 (N_8545,N_4349,N_4222);
nor U8546 (N_8546,N_3617,N_2895);
xnor U8547 (N_8547,N_2666,N_3190);
or U8548 (N_8548,N_2720,N_2444);
and U8549 (N_8549,N_2181,N_1074);
nor U8550 (N_8550,N_4005,N_4419);
nand U8551 (N_8551,N_1450,N_4615);
or U8552 (N_8552,N_1737,N_4657);
nand U8553 (N_8553,N_959,N_3546);
nand U8554 (N_8554,N_229,N_144);
or U8555 (N_8555,N_220,N_778);
nor U8556 (N_8556,N_4609,N_1656);
and U8557 (N_8557,N_2401,N_4665);
or U8558 (N_8558,N_100,N_3447);
and U8559 (N_8559,N_2858,N_1705);
and U8560 (N_8560,N_4923,N_1665);
and U8561 (N_8561,N_4825,N_373);
nor U8562 (N_8562,N_2022,N_1802);
or U8563 (N_8563,N_740,N_2376);
or U8564 (N_8564,N_4471,N_4545);
or U8565 (N_8565,N_154,N_458);
nor U8566 (N_8566,N_2388,N_1519);
or U8567 (N_8567,N_1999,N_3459);
nand U8568 (N_8568,N_1883,N_604);
nor U8569 (N_8569,N_443,N_1223);
nand U8570 (N_8570,N_477,N_100);
and U8571 (N_8571,N_29,N_3739);
and U8572 (N_8572,N_1272,N_65);
nor U8573 (N_8573,N_3398,N_2694);
nor U8574 (N_8574,N_3123,N_3889);
nand U8575 (N_8575,N_1130,N_1168);
or U8576 (N_8576,N_2507,N_3552);
and U8577 (N_8577,N_4352,N_3226);
nor U8578 (N_8578,N_558,N_4061);
and U8579 (N_8579,N_4516,N_1849);
or U8580 (N_8580,N_3803,N_3269);
or U8581 (N_8581,N_4042,N_2759);
nand U8582 (N_8582,N_4563,N_1693);
nand U8583 (N_8583,N_3703,N_3404);
or U8584 (N_8584,N_91,N_89);
or U8585 (N_8585,N_2096,N_1899);
or U8586 (N_8586,N_478,N_397);
or U8587 (N_8587,N_598,N_2615);
and U8588 (N_8588,N_3427,N_1985);
and U8589 (N_8589,N_4828,N_959);
nand U8590 (N_8590,N_661,N_4093);
and U8591 (N_8591,N_1119,N_4052);
or U8592 (N_8592,N_657,N_2762);
nor U8593 (N_8593,N_1928,N_3231);
or U8594 (N_8594,N_479,N_130);
or U8595 (N_8595,N_471,N_3759);
xor U8596 (N_8596,N_4543,N_1129);
nor U8597 (N_8597,N_3757,N_3204);
and U8598 (N_8598,N_1779,N_578);
nor U8599 (N_8599,N_2603,N_4338);
or U8600 (N_8600,N_4891,N_1803);
nor U8601 (N_8601,N_3372,N_3499);
nand U8602 (N_8602,N_4566,N_291);
nand U8603 (N_8603,N_4202,N_328);
and U8604 (N_8604,N_567,N_1653);
nor U8605 (N_8605,N_4518,N_1707);
nor U8606 (N_8606,N_2267,N_1869);
or U8607 (N_8607,N_2417,N_3851);
or U8608 (N_8608,N_2345,N_4534);
or U8609 (N_8609,N_3023,N_3073);
and U8610 (N_8610,N_4299,N_4320);
nand U8611 (N_8611,N_578,N_720);
nor U8612 (N_8612,N_2027,N_1213);
or U8613 (N_8613,N_4562,N_4227);
or U8614 (N_8614,N_4452,N_2350);
and U8615 (N_8615,N_3164,N_2152);
and U8616 (N_8616,N_4443,N_4786);
nor U8617 (N_8617,N_3639,N_34);
and U8618 (N_8618,N_1285,N_4408);
nand U8619 (N_8619,N_972,N_4186);
or U8620 (N_8620,N_1125,N_4497);
or U8621 (N_8621,N_3539,N_2652);
nor U8622 (N_8622,N_3336,N_2382);
nor U8623 (N_8623,N_3839,N_3609);
or U8624 (N_8624,N_3124,N_2529);
nand U8625 (N_8625,N_4731,N_524);
or U8626 (N_8626,N_363,N_2505);
or U8627 (N_8627,N_2869,N_2941);
nor U8628 (N_8628,N_1308,N_906);
xor U8629 (N_8629,N_1208,N_4243);
nand U8630 (N_8630,N_3061,N_3008);
nand U8631 (N_8631,N_4148,N_932);
or U8632 (N_8632,N_762,N_2571);
and U8633 (N_8633,N_2259,N_2399);
nand U8634 (N_8634,N_1544,N_1646);
nor U8635 (N_8635,N_3047,N_4809);
or U8636 (N_8636,N_3793,N_4026);
and U8637 (N_8637,N_1935,N_2333);
or U8638 (N_8638,N_2200,N_1619);
and U8639 (N_8639,N_1732,N_1892);
nand U8640 (N_8640,N_260,N_727);
and U8641 (N_8641,N_388,N_539);
and U8642 (N_8642,N_1590,N_4751);
and U8643 (N_8643,N_4203,N_2814);
nor U8644 (N_8644,N_4836,N_3897);
nor U8645 (N_8645,N_634,N_1402);
or U8646 (N_8646,N_2712,N_3586);
and U8647 (N_8647,N_4224,N_4865);
nand U8648 (N_8648,N_3235,N_3789);
or U8649 (N_8649,N_303,N_4404);
and U8650 (N_8650,N_901,N_2874);
nor U8651 (N_8651,N_4912,N_2425);
or U8652 (N_8652,N_4330,N_893);
or U8653 (N_8653,N_2141,N_4456);
nand U8654 (N_8654,N_2729,N_3854);
and U8655 (N_8655,N_2308,N_3123);
nand U8656 (N_8656,N_2200,N_3556);
nand U8657 (N_8657,N_1508,N_4307);
nand U8658 (N_8658,N_3126,N_3012);
and U8659 (N_8659,N_648,N_3618);
or U8660 (N_8660,N_3516,N_56);
nor U8661 (N_8661,N_139,N_3100);
or U8662 (N_8662,N_3873,N_2665);
nand U8663 (N_8663,N_4856,N_731);
nand U8664 (N_8664,N_3484,N_1478);
nand U8665 (N_8665,N_275,N_3738);
nor U8666 (N_8666,N_3280,N_413);
nor U8667 (N_8667,N_2098,N_2500);
and U8668 (N_8668,N_589,N_2907);
or U8669 (N_8669,N_2046,N_4575);
nor U8670 (N_8670,N_2220,N_3994);
nand U8671 (N_8671,N_3301,N_65);
nor U8672 (N_8672,N_1196,N_1540);
or U8673 (N_8673,N_3370,N_1317);
nand U8674 (N_8674,N_4299,N_3361);
or U8675 (N_8675,N_3485,N_3641);
nand U8676 (N_8676,N_3325,N_3723);
nand U8677 (N_8677,N_4363,N_4097);
or U8678 (N_8678,N_3576,N_3836);
and U8679 (N_8679,N_3868,N_2858);
and U8680 (N_8680,N_3144,N_1962);
nand U8681 (N_8681,N_4236,N_2703);
or U8682 (N_8682,N_3086,N_3009);
nor U8683 (N_8683,N_3887,N_4365);
nor U8684 (N_8684,N_101,N_648);
and U8685 (N_8685,N_1782,N_931);
nor U8686 (N_8686,N_894,N_4628);
and U8687 (N_8687,N_3579,N_2739);
nand U8688 (N_8688,N_1584,N_2474);
and U8689 (N_8689,N_1704,N_1480);
nor U8690 (N_8690,N_509,N_2306);
and U8691 (N_8691,N_1951,N_3809);
nand U8692 (N_8692,N_1369,N_515);
and U8693 (N_8693,N_380,N_4940);
nand U8694 (N_8694,N_2617,N_122);
xor U8695 (N_8695,N_2154,N_2577);
or U8696 (N_8696,N_660,N_4931);
nor U8697 (N_8697,N_1940,N_681);
and U8698 (N_8698,N_4332,N_632);
nand U8699 (N_8699,N_4574,N_1050);
nand U8700 (N_8700,N_2989,N_3136);
and U8701 (N_8701,N_4307,N_2433);
or U8702 (N_8702,N_4980,N_168);
and U8703 (N_8703,N_2089,N_1611);
nand U8704 (N_8704,N_32,N_1039);
nand U8705 (N_8705,N_4526,N_2665);
and U8706 (N_8706,N_981,N_3760);
nand U8707 (N_8707,N_4582,N_1721);
nand U8708 (N_8708,N_1560,N_4890);
and U8709 (N_8709,N_3885,N_4852);
nor U8710 (N_8710,N_169,N_2524);
nand U8711 (N_8711,N_4552,N_2626);
or U8712 (N_8712,N_4545,N_292);
nor U8713 (N_8713,N_994,N_1547);
and U8714 (N_8714,N_1454,N_4071);
nand U8715 (N_8715,N_3610,N_1073);
or U8716 (N_8716,N_368,N_4252);
nand U8717 (N_8717,N_3568,N_3711);
nand U8718 (N_8718,N_3169,N_3512);
and U8719 (N_8719,N_1745,N_1312);
nand U8720 (N_8720,N_1133,N_3014);
nor U8721 (N_8721,N_215,N_3053);
nor U8722 (N_8722,N_1475,N_4008);
nor U8723 (N_8723,N_2969,N_3699);
nor U8724 (N_8724,N_2995,N_4883);
nand U8725 (N_8725,N_3329,N_1923);
or U8726 (N_8726,N_3516,N_780);
and U8727 (N_8727,N_491,N_2719);
or U8728 (N_8728,N_596,N_3862);
or U8729 (N_8729,N_1066,N_3247);
nor U8730 (N_8730,N_3393,N_927);
and U8731 (N_8731,N_789,N_197);
nand U8732 (N_8732,N_4431,N_4179);
nand U8733 (N_8733,N_685,N_81);
nor U8734 (N_8734,N_1294,N_2111);
and U8735 (N_8735,N_3227,N_1849);
and U8736 (N_8736,N_3037,N_4254);
xnor U8737 (N_8737,N_4599,N_1500);
nand U8738 (N_8738,N_2612,N_4653);
and U8739 (N_8739,N_501,N_1379);
nand U8740 (N_8740,N_510,N_2940);
and U8741 (N_8741,N_2754,N_2832);
nor U8742 (N_8742,N_4474,N_2668);
nor U8743 (N_8743,N_3849,N_31);
nand U8744 (N_8744,N_4300,N_4801);
nor U8745 (N_8745,N_2821,N_1241);
nand U8746 (N_8746,N_3439,N_3285);
and U8747 (N_8747,N_2038,N_812);
nand U8748 (N_8748,N_2522,N_3254);
nor U8749 (N_8749,N_4366,N_3713);
nand U8750 (N_8750,N_954,N_2511);
and U8751 (N_8751,N_2797,N_2024);
nor U8752 (N_8752,N_3213,N_2206);
nor U8753 (N_8753,N_2612,N_1484);
nand U8754 (N_8754,N_3988,N_3959);
nor U8755 (N_8755,N_1561,N_3042);
or U8756 (N_8756,N_1150,N_2750);
or U8757 (N_8757,N_2478,N_2351);
nor U8758 (N_8758,N_4943,N_4135);
and U8759 (N_8759,N_4254,N_4444);
nand U8760 (N_8760,N_476,N_1787);
or U8761 (N_8761,N_350,N_2339);
and U8762 (N_8762,N_2120,N_3765);
and U8763 (N_8763,N_2689,N_2049);
nor U8764 (N_8764,N_4105,N_3309);
or U8765 (N_8765,N_4796,N_254);
and U8766 (N_8766,N_2774,N_1383);
nand U8767 (N_8767,N_1334,N_275);
nand U8768 (N_8768,N_223,N_3788);
or U8769 (N_8769,N_4777,N_1155);
nand U8770 (N_8770,N_4772,N_4011);
xnor U8771 (N_8771,N_405,N_2308);
and U8772 (N_8772,N_2066,N_4437);
nor U8773 (N_8773,N_2701,N_3162);
nand U8774 (N_8774,N_1042,N_2627);
and U8775 (N_8775,N_894,N_611);
nand U8776 (N_8776,N_134,N_1258);
or U8777 (N_8777,N_3988,N_331);
and U8778 (N_8778,N_105,N_837);
and U8779 (N_8779,N_4674,N_4068);
nor U8780 (N_8780,N_1731,N_1460);
nor U8781 (N_8781,N_2244,N_820);
xor U8782 (N_8782,N_4636,N_4652);
nand U8783 (N_8783,N_3502,N_3960);
and U8784 (N_8784,N_1716,N_473);
nor U8785 (N_8785,N_4396,N_2813);
nand U8786 (N_8786,N_2042,N_2687);
or U8787 (N_8787,N_945,N_819);
and U8788 (N_8788,N_4908,N_2331);
nand U8789 (N_8789,N_334,N_988);
nor U8790 (N_8790,N_1968,N_2055);
nor U8791 (N_8791,N_4375,N_823);
nor U8792 (N_8792,N_920,N_4401);
and U8793 (N_8793,N_2358,N_4114);
xnor U8794 (N_8794,N_3606,N_4307);
nand U8795 (N_8795,N_1508,N_3124);
and U8796 (N_8796,N_2480,N_2944);
or U8797 (N_8797,N_2384,N_3208);
nor U8798 (N_8798,N_4495,N_201);
xor U8799 (N_8799,N_1267,N_4761);
nand U8800 (N_8800,N_2624,N_3321);
or U8801 (N_8801,N_402,N_1058);
and U8802 (N_8802,N_3105,N_3545);
and U8803 (N_8803,N_2938,N_4624);
or U8804 (N_8804,N_2141,N_2378);
and U8805 (N_8805,N_1351,N_4019);
or U8806 (N_8806,N_3013,N_3805);
or U8807 (N_8807,N_2979,N_1106);
nor U8808 (N_8808,N_3531,N_4675);
and U8809 (N_8809,N_1696,N_2742);
and U8810 (N_8810,N_1506,N_4026);
nor U8811 (N_8811,N_278,N_2220);
nor U8812 (N_8812,N_1848,N_4983);
or U8813 (N_8813,N_3782,N_945);
and U8814 (N_8814,N_1845,N_1920);
nor U8815 (N_8815,N_939,N_2017);
nand U8816 (N_8816,N_1605,N_366);
and U8817 (N_8817,N_286,N_458);
nor U8818 (N_8818,N_1903,N_33);
or U8819 (N_8819,N_2738,N_3158);
or U8820 (N_8820,N_4717,N_3807);
nand U8821 (N_8821,N_3159,N_3186);
or U8822 (N_8822,N_3650,N_24);
nand U8823 (N_8823,N_4402,N_4436);
nand U8824 (N_8824,N_67,N_4558);
nor U8825 (N_8825,N_4813,N_4761);
and U8826 (N_8826,N_1927,N_4373);
nor U8827 (N_8827,N_4862,N_3456);
or U8828 (N_8828,N_1292,N_4298);
and U8829 (N_8829,N_770,N_474);
or U8830 (N_8830,N_1270,N_1850);
and U8831 (N_8831,N_4514,N_1129);
and U8832 (N_8832,N_1739,N_2914);
or U8833 (N_8833,N_4572,N_3785);
and U8834 (N_8834,N_710,N_628);
nand U8835 (N_8835,N_497,N_2221);
nand U8836 (N_8836,N_1369,N_2687);
or U8837 (N_8837,N_3872,N_2835);
or U8838 (N_8838,N_3775,N_372);
nand U8839 (N_8839,N_671,N_4026);
nand U8840 (N_8840,N_3267,N_1863);
nand U8841 (N_8841,N_370,N_4847);
or U8842 (N_8842,N_4112,N_1136);
nand U8843 (N_8843,N_3406,N_2399);
or U8844 (N_8844,N_1341,N_3103);
or U8845 (N_8845,N_1269,N_2781);
or U8846 (N_8846,N_2133,N_3784);
nor U8847 (N_8847,N_3223,N_1101);
nor U8848 (N_8848,N_911,N_1010);
nor U8849 (N_8849,N_1305,N_2343);
nand U8850 (N_8850,N_60,N_2088);
nor U8851 (N_8851,N_3594,N_305);
nand U8852 (N_8852,N_3644,N_2106);
nand U8853 (N_8853,N_3313,N_279);
nor U8854 (N_8854,N_3394,N_164);
nand U8855 (N_8855,N_3918,N_2932);
and U8856 (N_8856,N_4535,N_1332);
and U8857 (N_8857,N_133,N_4700);
or U8858 (N_8858,N_3413,N_2311);
and U8859 (N_8859,N_975,N_3955);
and U8860 (N_8860,N_2757,N_4390);
nand U8861 (N_8861,N_4706,N_4372);
nand U8862 (N_8862,N_1895,N_519);
or U8863 (N_8863,N_4487,N_3624);
nand U8864 (N_8864,N_4259,N_2737);
and U8865 (N_8865,N_3738,N_3051);
or U8866 (N_8866,N_3071,N_197);
and U8867 (N_8867,N_511,N_1227);
nor U8868 (N_8868,N_2507,N_1378);
or U8869 (N_8869,N_1645,N_850);
nand U8870 (N_8870,N_3759,N_4011);
nor U8871 (N_8871,N_3185,N_3158);
or U8872 (N_8872,N_3963,N_4106);
nor U8873 (N_8873,N_4469,N_3168);
nor U8874 (N_8874,N_869,N_4182);
or U8875 (N_8875,N_4101,N_951);
and U8876 (N_8876,N_3032,N_390);
nand U8877 (N_8877,N_3948,N_1758);
and U8878 (N_8878,N_2341,N_2580);
or U8879 (N_8879,N_149,N_4770);
nor U8880 (N_8880,N_4246,N_2852);
and U8881 (N_8881,N_3441,N_439);
and U8882 (N_8882,N_4186,N_2865);
or U8883 (N_8883,N_2477,N_3687);
and U8884 (N_8884,N_4477,N_1718);
nand U8885 (N_8885,N_1196,N_1554);
and U8886 (N_8886,N_4406,N_2264);
nor U8887 (N_8887,N_297,N_197);
and U8888 (N_8888,N_3637,N_955);
or U8889 (N_8889,N_3719,N_4192);
and U8890 (N_8890,N_632,N_2568);
nor U8891 (N_8891,N_1516,N_2357);
or U8892 (N_8892,N_2440,N_3669);
and U8893 (N_8893,N_992,N_3457);
and U8894 (N_8894,N_843,N_4221);
and U8895 (N_8895,N_3244,N_4110);
nor U8896 (N_8896,N_241,N_706);
xor U8897 (N_8897,N_4874,N_1030);
and U8898 (N_8898,N_4031,N_2754);
nand U8899 (N_8899,N_3799,N_3696);
nand U8900 (N_8900,N_3406,N_375);
nor U8901 (N_8901,N_2208,N_1494);
and U8902 (N_8902,N_3800,N_3355);
or U8903 (N_8903,N_261,N_2188);
nor U8904 (N_8904,N_248,N_2635);
and U8905 (N_8905,N_235,N_4087);
or U8906 (N_8906,N_2761,N_2077);
and U8907 (N_8907,N_4867,N_1358);
nor U8908 (N_8908,N_3938,N_5);
and U8909 (N_8909,N_3161,N_2104);
or U8910 (N_8910,N_801,N_3167);
nand U8911 (N_8911,N_954,N_4313);
nor U8912 (N_8912,N_3160,N_4043);
and U8913 (N_8913,N_840,N_1529);
or U8914 (N_8914,N_3519,N_915);
or U8915 (N_8915,N_2648,N_1146);
nor U8916 (N_8916,N_4611,N_1609);
nor U8917 (N_8917,N_3615,N_4305);
or U8918 (N_8918,N_2129,N_2765);
and U8919 (N_8919,N_736,N_3407);
nor U8920 (N_8920,N_572,N_2253);
or U8921 (N_8921,N_2894,N_1139);
nand U8922 (N_8922,N_3793,N_26);
or U8923 (N_8923,N_912,N_1487);
or U8924 (N_8924,N_3884,N_3474);
or U8925 (N_8925,N_4297,N_3802);
xor U8926 (N_8926,N_257,N_1065);
nor U8927 (N_8927,N_1810,N_2098);
nand U8928 (N_8928,N_740,N_217);
nand U8929 (N_8929,N_3496,N_1897);
and U8930 (N_8930,N_4479,N_10);
nor U8931 (N_8931,N_3633,N_3026);
or U8932 (N_8932,N_1834,N_1950);
nand U8933 (N_8933,N_3684,N_1745);
and U8934 (N_8934,N_3904,N_567);
nand U8935 (N_8935,N_223,N_1738);
nor U8936 (N_8936,N_4029,N_2189);
or U8937 (N_8937,N_4783,N_933);
nor U8938 (N_8938,N_1499,N_4020);
nor U8939 (N_8939,N_3931,N_2182);
nor U8940 (N_8940,N_3581,N_4971);
nor U8941 (N_8941,N_3421,N_677);
or U8942 (N_8942,N_1200,N_2673);
or U8943 (N_8943,N_4022,N_807);
nor U8944 (N_8944,N_1233,N_798);
nor U8945 (N_8945,N_1686,N_2359);
nand U8946 (N_8946,N_4941,N_794);
xnor U8947 (N_8947,N_2956,N_4485);
and U8948 (N_8948,N_4296,N_4871);
and U8949 (N_8949,N_678,N_4001);
nor U8950 (N_8950,N_2667,N_227);
and U8951 (N_8951,N_180,N_3095);
nor U8952 (N_8952,N_995,N_4930);
nor U8953 (N_8953,N_1546,N_3651);
and U8954 (N_8954,N_3848,N_1729);
and U8955 (N_8955,N_4170,N_2412);
nor U8956 (N_8956,N_1130,N_3523);
nand U8957 (N_8957,N_4104,N_2874);
and U8958 (N_8958,N_4142,N_2924);
nor U8959 (N_8959,N_4255,N_2400);
nor U8960 (N_8960,N_3140,N_71);
nand U8961 (N_8961,N_2042,N_2980);
nor U8962 (N_8962,N_2951,N_4732);
and U8963 (N_8963,N_4497,N_1944);
nor U8964 (N_8964,N_4507,N_2814);
or U8965 (N_8965,N_1215,N_3508);
and U8966 (N_8966,N_2430,N_3516);
or U8967 (N_8967,N_4733,N_4504);
or U8968 (N_8968,N_1552,N_3033);
and U8969 (N_8969,N_1953,N_3498);
nand U8970 (N_8970,N_3313,N_1796);
nand U8971 (N_8971,N_1917,N_3605);
nor U8972 (N_8972,N_3262,N_2858);
or U8973 (N_8973,N_296,N_1627);
or U8974 (N_8974,N_127,N_3592);
nor U8975 (N_8975,N_1901,N_1437);
and U8976 (N_8976,N_71,N_3815);
and U8977 (N_8977,N_2767,N_2714);
or U8978 (N_8978,N_2449,N_4039);
and U8979 (N_8979,N_3036,N_2269);
or U8980 (N_8980,N_1149,N_293);
nand U8981 (N_8981,N_53,N_845);
nor U8982 (N_8982,N_4513,N_4990);
or U8983 (N_8983,N_2578,N_2450);
or U8984 (N_8984,N_2853,N_3481);
or U8985 (N_8985,N_2514,N_525);
or U8986 (N_8986,N_1313,N_1011);
and U8987 (N_8987,N_2271,N_996);
nor U8988 (N_8988,N_3425,N_4528);
nand U8989 (N_8989,N_2924,N_480);
nand U8990 (N_8990,N_1224,N_2282);
nand U8991 (N_8991,N_3167,N_2501);
nand U8992 (N_8992,N_216,N_3591);
nor U8993 (N_8993,N_2504,N_2323);
xnor U8994 (N_8994,N_2391,N_4176);
or U8995 (N_8995,N_4272,N_2415);
nor U8996 (N_8996,N_403,N_3455);
or U8997 (N_8997,N_1727,N_2472);
and U8998 (N_8998,N_2457,N_3226);
and U8999 (N_8999,N_4504,N_288);
and U9000 (N_9000,N_2683,N_3013);
and U9001 (N_9001,N_2518,N_2725);
and U9002 (N_9002,N_69,N_2063);
and U9003 (N_9003,N_142,N_4390);
and U9004 (N_9004,N_370,N_3441);
or U9005 (N_9005,N_2710,N_3425);
nand U9006 (N_9006,N_4434,N_1023);
or U9007 (N_9007,N_1314,N_3400);
and U9008 (N_9008,N_3695,N_4388);
and U9009 (N_9009,N_3407,N_1650);
nand U9010 (N_9010,N_3500,N_4016);
nand U9011 (N_9011,N_2673,N_4048);
nand U9012 (N_9012,N_810,N_3);
nor U9013 (N_9013,N_1808,N_3476);
nor U9014 (N_9014,N_4988,N_2470);
or U9015 (N_9015,N_1288,N_4796);
nand U9016 (N_9016,N_2168,N_406);
and U9017 (N_9017,N_4452,N_3393);
and U9018 (N_9018,N_2822,N_2843);
or U9019 (N_9019,N_389,N_1664);
and U9020 (N_9020,N_228,N_3826);
nand U9021 (N_9021,N_978,N_4890);
nand U9022 (N_9022,N_3060,N_4756);
or U9023 (N_9023,N_3542,N_1665);
nor U9024 (N_9024,N_3519,N_506);
and U9025 (N_9025,N_229,N_4168);
or U9026 (N_9026,N_1490,N_3240);
nand U9027 (N_9027,N_310,N_1274);
nand U9028 (N_9028,N_3216,N_2465);
nor U9029 (N_9029,N_4777,N_2591);
nand U9030 (N_9030,N_1903,N_4009);
and U9031 (N_9031,N_2995,N_4372);
and U9032 (N_9032,N_2418,N_1090);
nand U9033 (N_9033,N_2873,N_1852);
nor U9034 (N_9034,N_4248,N_4147);
nor U9035 (N_9035,N_3928,N_2776);
nand U9036 (N_9036,N_2937,N_2602);
nand U9037 (N_9037,N_3651,N_988);
or U9038 (N_9038,N_670,N_3291);
and U9039 (N_9039,N_4727,N_2230);
nor U9040 (N_9040,N_4437,N_17);
nand U9041 (N_9041,N_299,N_2491);
nor U9042 (N_9042,N_2974,N_186);
or U9043 (N_9043,N_1953,N_3497);
or U9044 (N_9044,N_1249,N_4022);
and U9045 (N_9045,N_1958,N_4562);
and U9046 (N_9046,N_3688,N_2876);
nor U9047 (N_9047,N_2976,N_2440);
nor U9048 (N_9048,N_1161,N_1757);
or U9049 (N_9049,N_1068,N_1938);
and U9050 (N_9050,N_131,N_3484);
nor U9051 (N_9051,N_1189,N_1278);
or U9052 (N_9052,N_3819,N_1803);
nand U9053 (N_9053,N_4008,N_791);
nor U9054 (N_9054,N_129,N_271);
nand U9055 (N_9055,N_1498,N_1274);
and U9056 (N_9056,N_4962,N_56);
nand U9057 (N_9057,N_4464,N_703);
and U9058 (N_9058,N_2950,N_3769);
nor U9059 (N_9059,N_1000,N_4801);
nand U9060 (N_9060,N_1556,N_2676);
nor U9061 (N_9061,N_328,N_2001);
nand U9062 (N_9062,N_3592,N_4368);
nor U9063 (N_9063,N_292,N_2371);
or U9064 (N_9064,N_3110,N_3506);
nand U9065 (N_9065,N_255,N_2395);
nor U9066 (N_9066,N_4592,N_3139);
nor U9067 (N_9067,N_2600,N_2984);
and U9068 (N_9068,N_4551,N_668);
nor U9069 (N_9069,N_3548,N_4740);
nand U9070 (N_9070,N_3471,N_3892);
and U9071 (N_9071,N_944,N_2037);
nand U9072 (N_9072,N_1199,N_745);
or U9073 (N_9073,N_4063,N_2446);
nand U9074 (N_9074,N_1026,N_262);
nor U9075 (N_9075,N_2117,N_527);
and U9076 (N_9076,N_555,N_3831);
and U9077 (N_9077,N_3281,N_1510);
nor U9078 (N_9078,N_342,N_381);
nor U9079 (N_9079,N_984,N_2809);
or U9080 (N_9080,N_649,N_189);
nor U9081 (N_9081,N_3534,N_4091);
nor U9082 (N_9082,N_3857,N_4899);
nor U9083 (N_9083,N_1825,N_3017);
nand U9084 (N_9084,N_3858,N_3291);
and U9085 (N_9085,N_355,N_4488);
nand U9086 (N_9086,N_3770,N_3841);
nand U9087 (N_9087,N_641,N_1739);
and U9088 (N_9088,N_139,N_2614);
nand U9089 (N_9089,N_3019,N_3479);
and U9090 (N_9090,N_1756,N_2392);
and U9091 (N_9091,N_4499,N_119);
nand U9092 (N_9092,N_4364,N_427);
or U9093 (N_9093,N_4397,N_1416);
nor U9094 (N_9094,N_1063,N_1345);
nor U9095 (N_9095,N_3909,N_371);
or U9096 (N_9096,N_3469,N_4967);
or U9097 (N_9097,N_3336,N_640);
nand U9098 (N_9098,N_2092,N_1458);
nand U9099 (N_9099,N_889,N_4449);
nor U9100 (N_9100,N_370,N_1897);
nand U9101 (N_9101,N_4949,N_3509);
or U9102 (N_9102,N_1260,N_1464);
and U9103 (N_9103,N_2061,N_484);
or U9104 (N_9104,N_585,N_1282);
or U9105 (N_9105,N_2061,N_2240);
or U9106 (N_9106,N_4969,N_2061);
nor U9107 (N_9107,N_3686,N_1336);
nand U9108 (N_9108,N_461,N_3810);
or U9109 (N_9109,N_4982,N_2621);
or U9110 (N_9110,N_3954,N_2752);
nand U9111 (N_9111,N_1276,N_2027);
or U9112 (N_9112,N_4429,N_3737);
or U9113 (N_9113,N_4254,N_2822);
or U9114 (N_9114,N_4405,N_4668);
or U9115 (N_9115,N_2787,N_4782);
nand U9116 (N_9116,N_531,N_2952);
or U9117 (N_9117,N_866,N_4064);
and U9118 (N_9118,N_3718,N_1846);
nor U9119 (N_9119,N_2714,N_3938);
and U9120 (N_9120,N_2907,N_2128);
nand U9121 (N_9121,N_110,N_2620);
nand U9122 (N_9122,N_103,N_599);
or U9123 (N_9123,N_3743,N_2536);
nand U9124 (N_9124,N_2467,N_4278);
nand U9125 (N_9125,N_4916,N_4175);
and U9126 (N_9126,N_4912,N_2681);
and U9127 (N_9127,N_4233,N_2793);
or U9128 (N_9128,N_1506,N_4726);
nand U9129 (N_9129,N_3472,N_1943);
nor U9130 (N_9130,N_4044,N_4594);
or U9131 (N_9131,N_1117,N_509);
nand U9132 (N_9132,N_2752,N_3207);
nor U9133 (N_9133,N_4611,N_3457);
or U9134 (N_9134,N_2773,N_2544);
or U9135 (N_9135,N_2113,N_4528);
nor U9136 (N_9136,N_4971,N_1634);
nand U9137 (N_9137,N_2359,N_1800);
nor U9138 (N_9138,N_2403,N_4629);
nor U9139 (N_9139,N_4005,N_4026);
or U9140 (N_9140,N_2731,N_3152);
nor U9141 (N_9141,N_2784,N_1908);
nand U9142 (N_9142,N_175,N_478);
nand U9143 (N_9143,N_2905,N_1543);
or U9144 (N_9144,N_4410,N_1426);
and U9145 (N_9145,N_2691,N_2333);
nor U9146 (N_9146,N_4424,N_1028);
nand U9147 (N_9147,N_1826,N_4261);
or U9148 (N_9148,N_3311,N_1271);
or U9149 (N_9149,N_4813,N_4679);
and U9150 (N_9150,N_2796,N_1098);
and U9151 (N_9151,N_355,N_3608);
and U9152 (N_9152,N_2223,N_1902);
nand U9153 (N_9153,N_1318,N_3916);
nand U9154 (N_9154,N_1199,N_4351);
nand U9155 (N_9155,N_70,N_195);
nor U9156 (N_9156,N_2366,N_1365);
or U9157 (N_9157,N_3320,N_2545);
nand U9158 (N_9158,N_2486,N_3418);
nor U9159 (N_9159,N_2378,N_4995);
and U9160 (N_9160,N_3748,N_1357);
or U9161 (N_9161,N_2468,N_3661);
nor U9162 (N_9162,N_1315,N_4151);
and U9163 (N_9163,N_3878,N_4363);
nor U9164 (N_9164,N_3451,N_1253);
xor U9165 (N_9165,N_4929,N_291);
nor U9166 (N_9166,N_679,N_4070);
nand U9167 (N_9167,N_4930,N_1919);
nor U9168 (N_9168,N_4808,N_1200);
nor U9169 (N_9169,N_4523,N_4719);
nor U9170 (N_9170,N_1111,N_4487);
nor U9171 (N_9171,N_1,N_445);
and U9172 (N_9172,N_3713,N_4404);
and U9173 (N_9173,N_3874,N_4657);
nand U9174 (N_9174,N_1264,N_2276);
nand U9175 (N_9175,N_2844,N_43);
and U9176 (N_9176,N_1728,N_813);
and U9177 (N_9177,N_1969,N_2618);
or U9178 (N_9178,N_2607,N_110);
nor U9179 (N_9179,N_1407,N_3728);
nor U9180 (N_9180,N_2712,N_1103);
and U9181 (N_9181,N_3739,N_1760);
and U9182 (N_9182,N_2213,N_4305);
or U9183 (N_9183,N_2937,N_509);
nand U9184 (N_9184,N_1225,N_2913);
or U9185 (N_9185,N_4926,N_3872);
or U9186 (N_9186,N_2315,N_1697);
nor U9187 (N_9187,N_3715,N_2923);
nand U9188 (N_9188,N_165,N_1676);
nor U9189 (N_9189,N_2819,N_1176);
or U9190 (N_9190,N_1930,N_2483);
and U9191 (N_9191,N_31,N_1144);
and U9192 (N_9192,N_3895,N_3296);
and U9193 (N_9193,N_4322,N_4354);
or U9194 (N_9194,N_4561,N_3846);
nand U9195 (N_9195,N_696,N_1159);
nor U9196 (N_9196,N_98,N_508);
nand U9197 (N_9197,N_1599,N_364);
and U9198 (N_9198,N_938,N_4762);
and U9199 (N_9199,N_3297,N_969);
nand U9200 (N_9200,N_2166,N_4503);
nor U9201 (N_9201,N_437,N_2238);
or U9202 (N_9202,N_2775,N_1685);
nor U9203 (N_9203,N_417,N_4435);
and U9204 (N_9204,N_1736,N_3680);
or U9205 (N_9205,N_3582,N_389);
nor U9206 (N_9206,N_4152,N_1613);
or U9207 (N_9207,N_3819,N_180);
nand U9208 (N_9208,N_3726,N_3482);
nor U9209 (N_9209,N_3980,N_4360);
or U9210 (N_9210,N_706,N_3402);
nand U9211 (N_9211,N_1390,N_392);
nor U9212 (N_9212,N_1495,N_2442);
and U9213 (N_9213,N_2670,N_1009);
nand U9214 (N_9214,N_4978,N_4312);
and U9215 (N_9215,N_134,N_2283);
and U9216 (N_9216,N_3872,N_1889);
and U9217 (N_9217,N_4575,N_196);
nor U9218 (N_9218,N_901,N_4230);
and U9219 (N_9219,N_1622,N_4981);
or U9220 (N_9220,N_2518,N_1011);
nand U9221 (N_9221,N_1139,N_1498);
or U9222 (N_9222,N_1914,N_3371);
and U9223 (N_9223,N_2001,N_2643);
nand U9224 (N_9224,N_666,N_3620);
nand U9225 (N_9225,N_2248,N_4807);
nand U9226 (N_9226,N_2386,N_4517);
or U9227 (N_9227,N_3024,N_4389);
or U9228 (N_9228,N_648,N_1821);
nand U9229 (N_9229,N_493,N_2931);
nor U9230 (N_9230,N_3549,N_2465);
nand U9231 (N_9231,N_1732,N_2506);
and U9232 (N_9232,N_3942,N_3027);
nand U9233 (N_9233,N_4975,N_4961);
or U9234 (N_9234,N_585,N_2843);
nand U9235 (N_9235,N_2590,N_259);
or U9236 (N_9236,N_358,N_2340);
nor U9237 (N_9237,N_627,N_1122);
and U9238 (N_9238,N_1951,N_2802);
nand U9239 (N_9239,N_859,N_4434);
or U9240 (N_9240,N_2030,N_1716);
or U9241 (N_9241,N_1885,N_4122);
nand U9242 (N_9242,N_390,N_2703);
and U9243 (N_9243,N_240,N_137);
or U9244 (N_9244,N_2322,N_4088);
nand U9245 (N_9245,N_2123,N_1409);
nor U9246 (N_9246,N_4609,N_4839);
nand U9247 (N_9247,N_2549,N_514);
nand U9248 (N_9248,N_4976,N_2013);
nor U9249 (N_9249,N_4533,N_2836);
nand U9250 (N_9250,N_4420,N_1480);
or U9251 (N_9251,N_2959,N_4369);
or U9252 (N_9252,N_580,N_1106);
nor U9253 (N_9253,N_3448,N_1598);
and U9254 (N_9254,N_4005,N_1117);
or U9255 (N_9255,N_2990,N_463);
nand U9256 (N_9256,N_4888,N_529);
nand U9257 (N_9257,N_3467,N_1788);
xnor U9258 (N_9258,N_3720,N_1042);
or U9259 (N_9259,N_498,N_4429);
or U9260 (N_9260,N_3357,N_3297);
or U9261 (N_9261,N_3360,N_3601);
nand U9262 (N_9262,N_3239,N_968);
nand U9263 (N_9263,N_2062,N_769);
nor U9264 (N_9264,N_394,N_2318);
nor U9265 (N_9265,N_584,N_2266);
and U9266 (N_9266,N_1035,N_1242);
nand U9267 (N_9267,N_3521,N_1495);
nand U9268 (N_9268,N_4054,N_3066);
or U9269 (N_9269,N_4634,N_4290);
nor U9270 (N_9270,N_693,N_3828);
nand U9271 (N_9271,N_3698,N_2611);
nand U9272 (N_9272,N_588,N_1697);
or U9273 (N_9273,N_3301,N_4282);
nand U9274 (N_9274,N_629,N_2197);
nor U9275 (N_9275,N_4280,N_4526);
nand U9276 (N_9276,N_4397,N_4005);
and U9277 (N_9277,N_107,N_1011);
and U9278 (N_9278,N_2039,N_1392);
nand U9279 (N_9279,N_2131,N_2787);
nand U9280 (N_9280,N_3890,N_1670);
and U9281 (N_9281,N_3338,N_2126);
or U9282 (N_9282,N_4202,N_2435);
or U9283 (N_9283,N_3698,N_199);
nand U9284 (N_9284,N_1510,N_735);
and U9285 (N_9285,N_679,N_1984);
nand U9286 (N_9286,N_3578,N_2329);
and U9287 (N_9287,N_1888,N_1564);
and U9288 (N_9288,N_497,N_4969);
nand U9289 (N_9289,N_948,N_1280);
and U9290 (N_9290,N_639,N_50);
nor U9291 (N_9291,N_421,N_2664);
nand U9292 (N_9292,N_2257,N_2067);
nor U9293 (N_9293,N_447,N_3385);
nor U9294 (N_9294,N_3310,N_1425);
and U9295 (N_9295,N_4681,N_3881);
and U9296 (N_9296,N_1795,N_966);
or U9297 (N_9297,N_950,N_3199);
nor U9298 (N_9298,N_4418,N_1778);
xnor U9299 (N_9299,N_613,N_3825);
nor U9300 (N_9300,N_2586,N_3220);
nand U9301 (N_9301,N_1652,N_1160);
and U9302 (N_9302,N_4752,N_1481);
and U9303 (N_9303,N_1090,N_1866);
nand U9304 (N_9304,N_953,N_980);
nand U9305 (N_9305,N_4125,N_2616);
nor U9306 (N_9306,N_2896,N_1452);
nand U9307 (N_9307,N_2080,N_728);
nor U9308 (N_9308,N_3015,N_2317);
nand U9309 (N_9309,N_1107,N_3069);
and U9310 (N_9310,N_2064,N_2185);
or U9311 (N_9311,N_1190,N_235);
or U9312 (N_9312,N_1088,N_1749);
nand U9313 (N_9313,N_312,N_621);
and U9314 (N_9314,N_4634,N_1618);
nand U9315 (N_9315,N_1122,N_2320);
nand U9316 (N_9316,N_3858,N_2720);
and U9317 (N_9317,N_580,N_1878);
nor U9318 (N_9318,N_1873,N_3073);
nand U9319 (N_9319,N_1556,N_3424);
and U9320 (N_9320,N_2539,N_1850);
and U9321 (N_9321,N_2452,N_2450);
or U9322 (N_9322,N_3220,N_202);
nor U9323 (N_9323,N_3187,N_1116);
nor U9324 (N_9324,N_2607,N_250);
nand U9325 (N_9325,N_2096,N_1068);
nor U9326 (N_9326,N_1890,N_3503);
nor U9327 (N_9327,N_3942,N_1037);
or U9328 (N_9328,N_2016,N_4802);
or U9329 (N_9329,N_913,N_485);
and U9330 (N_9330,N_117,N_3384);
nand U9331 (N_9331,N_4286,N_3480);
and U9332 (N_9332,N_2278,N_2022);
nand U9333 (N_9333,N_29,N_4241);
nand U9334 (N_9334,N_689,N_2281);
nor U9335 (N_9335,N_1871,N_1435);
nand U9336 (N_9336,N_4290,N_3583);
nand U9337 (N_9337,N_2614,N_4822);
nor U9338 (N_9338,N_4619,N_2839);
nor U9339 (N_9339,N_1433,N_1808);
or U9340 (N_9340,N_2424,N_1504);
nand U9341 (N_9341,N_4026,N_3041);
nand U9342 (N_9342,N_3072,N_3611);
or U9343 (N_9343,N_69,N_387);
nor U9344 (N_9344,N_357,N_4419);
nand U9345 (N_9345,N_4697,N_1011);
or U9346 (N_9346,N_538,N_3196);
nor U9347 (N_9347,N_4689,N_3669);
or U9348 (N_9348,N_3905,N_1393);
nand U9349 (N_9349,N_3727,N_2559);
nor U9350 (N_9350,N_2603,N_1563);
nor U9351 (N_9351,N_695,N_4117);
and U9352 (N_9352,N_3702,N_4219);
nor U9353 (N_9353,N_184,N_4582);
and U9354 (N_9354,N_32,N_1007);
nor U9355 (N_9355,N_359,N_3041);
or U9356 (N_9356,N_2546,N_2103);
nand U9357 (N_9357,N_1615,N_1560);
nor U9358 (N_9358,N_2034,N_1864);
nor U9359 (N_9359,N_853,N_1981);
or U9360 (N_9360,N_541,N_1668);
xor U9361 (N_9361,N_903,N_3244);
nand U9362 (N_9362,N_4065,N_4889);
nand U9363 (N_9363,N_4132,N_4122);
nor U9364 (N_9364,N_1147,N_2959);
nor U9365 (N_9365,N_64,N_3172);
or U9366 (N_9366,N_1898,N_4729);
or U9367 (N_9367,N_4285,N_3640);
nand U9368 (N_9368,N_507,N_992);
nor U9369 (N_9369,N_4017,N_3436);
nand U9370 (N_9370,N_4717,N_74);
nor U9371 (N_9371,N_122,N_4399);
nand U9372 (N_9372,N_2768,N_3528);
nor U9373 (N_9373,N_2361,N_1702);
nor U9374 (N_9374,N_3234,N_2659);
and U9375 (N_9375,N_4443,N_648);
nand U9376 (N_9376,N_324,N_895);
nor U9377 (N_9377,N_316,N_3963);
nor U9378 (N_9378,N_472,N_4777);
and U9379 (N_9379,N_3134,N_2070);
nor U9380 (N_9380,N_4385,N_2961);
or U9381 (N_9381,N_1470,N_3220);
or U9382 (N_9382,N_4872,N_3124);
nand U9383 (N_9383,N_730,N_3718);
and U9384 (N_9384,N_3266,N_32);
nor U9385 (N_9385,N_191,N_1063);
or U9386 (N_9386,N_4320,N_245);
or U9387 (N_9387,N_860,N_2990);
or U9388 (N_9388,N_4901,N_3897);
and U9389 (N_9389,N_2944,N_2188);
and U9390 (N_9390,N_2419,N_1497);
or U9391 (N_9391,N_652,N_4305);
or U9392 (N_9392,N_2792,N_1334);
nand U9393 (N_9393,N_265,N_3147);
or U9394 (N_9394,N_239,N_3914);
nor U9395 (N_9395,N_78,N_695);
nand U9396 (N_9396,N_4007,N_3250);
nor U9397 (N_9397,N_1770,N_1241);
and U9398 (N_9398,N_1574,N_2885);
or U9399 (N_9399,N_3606,N_4133);
or U9400 (N_9400,N_1176,N_3782);
or U9401 (N_9401,N_2101,N_1767);
nand U9402 (N_9402,N_709,N_3196);
or U9403 (N_9403,N_2967,N_419);
nand U9404 (N_9404,N_3635,N_3537);
and U9405 (N_9405,N_2252,N_1551);
nor U9406 (N_9406,N_297,N_2551);
nand U9407 (N_9407,N_4380,N_2773);
and U9408 (N_9408,N_3243,N_4162);
nand U9409 (N_9409,N_2703,N_4145);
and U9410 (N_9410,N_4329,N_1686);
and U9411 (N_9411,N_4784,N_1393);
nor U9412 (N_9412,N_1672,N_3320);
and U9413 (N_9413,N_2576,N_3376);
nand U9414 (N_9414,N_3388,N_2603);
nand U9415 (N_9415,N_3221,N_2002);
or U9416 (N_9416,N_2474,N_2352);
nand U9417 (N_9417,N_4281,N_2865);
nand U9418 (N_9418,N_137,N_3781);
nand U9419 (N_9419,N_583,N_3175);
nor U9420 (N_9420,N_1869,N_3510);
nand U9421 (N_9421,N_456,N_1790);
or U9422 (N_9422,N_1183,N_1825);
and U9423 (N_9423,N_4310,N_451);
nor U9424 (N_9424,N_594,N_4286);
xor U9425 (N_9425,N_295,N_3501);
and U9426 (N_9426,N_3348,N_2050);
and U9427 (N_9427,N_4382,N_1681);
and U9428 (N_9428,N_3341,N_4106);
and U9429 (N_9429,N_3180,N_551);
xnor U9430 (N_9430,N_3967,N_3983);
or U9431 (N_9431,N_4538,N_169);
or U9432 (N_9432,N_3837,N_97);
nand U9433 (N_9433,N_4502,N_20);
or U9434 (N_9434,N_2578,N_3273);
or U9435 (N_9435,N_2802,N_1012);
nand U9436 (N_9436,N_2625,N_2142);
nor U9437 (N_9437,N_3731,N_1657);
and U9438 (N_9438,N_310,N_1878);
and U9439 (N_9439,N_3020,N_882);
and U9440 (N_9440,N_1230,N_2410);
xnor U9441 (N_9441,N_4738,N_3172);
nand U9442 (N_9442,N_4118,N_2353);
or U9443 (N_9443,N_2182,N_2769);
nand U9444 (N_9444,N_683,N_2358);
or U9445 (N_9445,N_3531,N_744);
nor U9446 (N_9446,N_3159,N_4419);
nor U9447 (N_9447,N_4100,N_1555);
nand U9448 (N_9448,N_3137,N_38);
or U9449 (N_9449,N_2216,N_624);
nor U9450 (N_9450,N_2998,N_1727);
and U9451 (N_9451,N_2637,N_448);
and U9452 (N_9452,N_1581,N_3970);
nand U9453 (N_9453,N_887,N_1330);
nand U9454 (N_9454,N_4910,N_2148);
and U9455 (N_9455,N_3951,N_3955);
or U9456 (N_9456,N_2885,N_2574);
nand U9457 (N_9457,N_1255,N_2826);
nor U9458 (N_9458,N_1145,N_1998);
nor U9459 (N_9459,N_551,N_1272);
nor U9460 (N_9460,N_1943,N_3904);
or U9461 (N_9461,N_2557,N_2976);
and U9462 (N_9462,N_4827,N_1532);
nand U9463 (N_9463,N_1695,N_300);
and U9464 (N_9464,N_2431,N_966);
nor U9465 (N_9465,N_2835,N_4863);
and U9466 (N_9466,N_1398,N_1851);
or U9467 (N_9467,N_798,N_4314);
or U9468 (N_9468,N_4151,N_404);
or U9469 (N_9469,N_2568,N_930);
nor U9470 (N_9470,N_379,N_650);
and U9471 (N_9471,N_3116,N_4763);
nand U9472 (N_9472,N_4954,N_4147);
or U9473 (N_9473,N_4064,N_1244);
or U9474 (N_9474,N_3544,N_3706);
or U9475 (N_9475,N_2723,N_2142);
nor U9476 (N_9476,N_1018,N_688);
nand U9477 (N_9477,N_3854,N_4301);
and U9478 (N_9478,N_4461,N_4254);
and U9479 (N_9479,N_4366,N_3525);
and U9480 (N_9480,N_3151,N_2877);
and U9481 (N_9481,N_3917,N_518);
and U9482 (N_9482,N_2726,N_4313);
and U9483 (N_9483,N_31,N_548);
nor U9484 (N_9484,N_4220,N_2713);
nor U9485 (N_9485,N_4767,N_3329);
nor U9486 (N_9486,N_2667,N_1107);
nor U9487 (N_9487,N_2054,N_391);
nand U9488 (N_9488,N_2655,N_4833);
or U9489 (N_9489,N_3485,N_1568);
and U9490 (N_9490,N_826,N_4419);
nand U9491 (N_9491,N_1303,N_3085);
nand U9492 (N_9492,N_2249,N_656);
nand U9493 (N_9493,N_4142,N_3296);
or U9494 (N_9494,N_4302,N_2116);
and U9495 (N_9495,N_4926,N_1726);
or U9496 (N_9496,N_444,N_2195);
nand U9497 (N_9497,N_3353,N_3136);
or U9498 (N_9498,N_2561,N_2275);
nor U9499 (N_9499,N_3501,N_1241);
nand U9500 (N_9500,N_1689,N_4967);
nand U9501 (N_9501,N_765,N_607);
or U9502 (N_9502,N_534,N_943);
and U9503 (N_9503,N_2446,N_3334);
and U9504 (N_9504,N_2370,N_2769);
nand U9505 (N_9505,N_3015,N_3921);
nand U9506 (N_9506,N_980,N_3028);
nor U9507 (N_9507,N_2666,N_3262);
nand U9508 (N_9508,N_3750,N_4987);
and U9509 (N_9509,N_2883,N_4947);
nor U9510 (N_9510,N_1064,N_617);
or U9511 (N_9511,N_3843,N_4268);
nor U9512 (N_9512,N_1168,N_1929);
nand U9513 (N_9513,N_3865,N_17);
nor U9514 (N_9514,N_1174,N_3819);
or U9515 (N_9515,N_4199,N_1849);
nor U9516 (N_9516,N_1199,N_3254);
nor U9517 (N_9517,N_4519,N_1536);
and U9518 (N_9518,N_4670,N_1024);
nor U9519 (N_9519,N_702,N_2162);
nand U9520 (N_9520,N_2726,N_4443);
nor U9521 (N_9521,N_642,N_2699);
or U9522 (N_9522,N_1974,N_3240);
nor U9523 (N_9523,N_3974,N_4127);
nor U9524 (N_9524,N_3688,N_4091);
nand U9525 (N_9525,N_4660,N_1156);
nand U9526 (N_9526,N_2723,N_3009);
nand U9527 (N_9527,N_3142,N_1636);
nand U9528 (N_9528,N_1613,N_3441);
and U9529 (N_9529,N_2090,N_4906);
and U9530 (N_9530,N_4614,N_3887);
nor U9531 (N_9531,N_4425,N_386);
nor U9532 (N_9532,N_3693,N_717);
nor U9533 (N_9533,N_1411,N_1991);
nor U9534 (N_9534,N_4964,N_2033);
nand U9535 (N_9535,N_2051,N_385);
and U9536 (N_9536,N_1838,N_484);
and U9537 (N_9537,N_1915,N_1282);
nand U9538 (N_9538,N_4176,N_4899);
nor U9539 (N_9539,N_1479,N_4034);
nand U9540 (N_9540,N_2776,N_1491);
or U9541 (N_9541,N_1898,N_2198);
or U9542 (N_9542,N_4426,N_1983);
and U9543 (N_9543,N_1362,N_2158);
and U9544 (N_9544,N_4800,N_3759);
nor U9545 (N_9545,N_4225,N_2426);
or U9546 (N_9546,N_110,N_2190);
nand U9547 (N_9547,N_1767,N_2993);
nor U9548 (N_9548,N_875,N_4125);
nand U9549 (N_9549,N_2843,N_3114);
or U9550 (N_9550,N_3442,N_3947);
or U9551 (N_9551,N_3746,N_4543);
or U9552 (N_9552,N_3661,N_3514);
nand U9553 (N_9553,N_3103,N_2206);
nor U9554 (N_9554,N_596,N_2889);
or U9555 (N_9555,N_4276,N_2572);
and U9556 (N_9556,N_810,N_4723);
nor U9557 (N_9557,N_2353,N_1542);
nand U9558 (N_9558,N_1159,N_4243);
nor U9559 (N_9559,N_2582,N_2071);
and U9560 (N_9560,N_4659,N_1087);
or U9561 (N_9561,N_236,N_3008);
nand U9562 (N_9562,N_1099,N_3080);
nor U9563 (N_9563,N_2724,N_203);
nor U9564 (N_9564,N_372,N_1346);
and U9565 (N_9565,N_703,N_1194);
nor U9566 (N_9566,N_2808,N_4896);
or U9567 (N_9567,N_1932,N_2681);
nand U9568 (N_9568,N_3874,N_4101);
nand U9569 (N_9569,N_3368,N_1875);
and U9570 (N_9570,N_1459,N_2802);
and U9571 (N_9571,N_2217,N_222);
and U9572 (N_9572,N_1918,N_3144);
xor U9573 (N_9573,N_3110,N_3450);
nor U9574 (N_9574,N_4458,N_1287);
or U9575 (N_9575,N_4091,N_2173);
nor U9576 (N_9576,N_1862,N_470);
nand U9577 (N_9577,N_3522,N_1609);
and U9578 (N_9578,N_4784,N_3652);
xnor U9579 (N_9579,N_1029,N_2714);
nor U9580 (N_9580,N_3832,N_3798);
or U9581 (N_9581,N_1868,N_1836);
nand U9582 (N_9582,N_956,N_2993);
and U9583 (N_9583,N_929,N_1970);
nor U9584 (N_9584,N_1663,N_3030);
nor U9585 (N_9585,N_1725,N_4216);
and U9586 (N_9586,N_2762,N_1714);
or U9587 (N_9587,N_1254,N_143);
and U9588 (N_9588,N_1862,N_2902);
and U9589 (N_9589,N_2089,N_4654);
nor U9590 (N_9590,N_1965,N_2539);
nor U9591 (N_9591,N_4603,N_1783);
nand U9592 (N_9592,N_2230,N_2176);
nand U9593 (N_9593,N_4632,N_2043);
nor U9594 (N_9594,N_4193,N_1117);
or U9595 (N_9595,N_1661,N_2765);
nor U9596 (N_9596,N_1425,N_2361);
and U9597 (N_9597,N_61,N_3058);
and U9598 (N_9598,N_1907,N_3143);
and U9599 (N_9599,N_2175,N_3096);
or U9600 (N_9600,N_4982,N_4198);
or U9601 (N_9601,N_4636,N_4803);
xor U9602 (N_9602,N_1638,N_4307);
or U9603 (N_9603,N_2660,N_1394);
nor U9604 (N_9604,N_2216,N_1452);
and U9605 (N_9605,N_1384,N_1370);
nor U9606 (N_9606,N_4807,N_3868);
nor U9607 (N_9607,N_1089,N_790);
nand U9608 (N_9608,N_612,N_1189);
or U9609 (N_9609,N_2486,N_3711);
xor U9610 (N_9610,N_4034,N_3700);
nor U9611 (N_9611,N_2469,N_794);
and U9612 (N_9612,N_4389,N_1324);
and U9613 (N_9613,N_1894,N_4724);
nand U9614 (N_9614,N_751,N_3452);
nor U9615 (N_9615,N_899,N_972);
and U9616 (N_9616,N_4877,N_4367);
and U9617 (N_9617,N_4240,N_1979);
nor U9618 (N_9618,N_2531,N_340);
or U9619 (N_9619,N_1892,N_1062);
or U9620 (N_9620,N_126,N_4635);
nor U9621 (N_9621,N_3534,N_4404);
nand U9622 (N_9622,N_3407,N_3427);
nor U9623 (N_9623,N_4562,N_2745);
and U9624 (N_9624,N_1684,N_3365);
and U9625 (N_9625,N_3481,N_2902);
and U9626 (N_9626,N_2136,N_858);
or U9627 (N_9627,N_4928,N_2051);
nor U9628 (N_9628,N_602,N_3598);
nor U9629 (N_9629,N_3999,N_2800);
xor U9630 (N_9630,N_3307,N_3714);
nand U9631 (N_9631,N_4506,N_630);
or U9632 (N_9632,N_4592,N_1714);
nor U9633 (N_9633,N_4128,N_2396);
nor U9634 (N_9634,N_858,N_2298);
xnor U9635 (N_9635,N_42,N_4290);
and U9636 (N_9636,N_2604,N_3448);
nand U9637 (N_9637,N_312,N_959);
nor U9638 (N_9638,N_858,N_3273);
nand U9639 (N_9639,N_3108,N_4520);
nand U9640 (N_9640,N_2047,N_836);
or U9641 (N_9641,N_3168,N_1869);
xor U9642 (N_9642,N_1596,N_277);
nor U9643 (N_9643,N_2247,N_3552);
and U9644 (N_9644,N_3027,N_4955);
and U9645 (N_9645,N_2756,N_685);
nor U9646 (N_9646,N_4826,N_1179);
nor U9647 (N_9647,N_83,N_2680);
nand U9648 (N_9648,N_747,N_3033);
or U9649 (N_9649,N_2805,N_3432);
and U9650 (N_9650,N_532,N_1623);
and U9651 (N_9651,N_3068,N_4628);
and U9652 (N_9652,N_398,N_4795);
nand U9653 (N_9653,N_3142,N_419);
and U9654 (N_9654,N_2218,N_3414);
nand U9655 (N_9655,N_4427,N_875);
and U9656 (N_9656,N_934,N_936);
nand U9657 (N_9657,N_1120,N_2640);
nor U9658 (N_9658,N_3171,N_4570);
or U9659 (N_9659,N_3012,N_1494);
nor U9660 (N_9660,N_1582,N_2452);
xnor U9661 (N_9661,N_2624,N_38);
and U9662 (N_9662,N_2023,N_3633);
nand U9663 (N_9663,N_4779,N_1095);
or U9664 (N_9664,N_1375,N_900);
or U9665 (N_9665,N_1753,N_1471);
or U9666 (N_9666,N_1896,N_2742);
nor U9667 (N_9667,N_1888,N_3430);
nand U9668 (N_9668,N_2812,N_4169);
or U9669 (N_9669,N_4215,N_1307);
nand U9670 (N_9670,N_1966,N_4805);
and U9671 (N_9671,N_1738,N_2591);
or U9672 (N_9672,N_2308,N_3911);
nor U9673 (N_9673,N_4249,N_1832);
or U9674 (N_9674,N_1506,N_4874);
nor U9675 (N_9675,N_498,N_4124);
and U9676 (N_9676,N_4098,N_1019);
nand U9677 (N_9677,N_991,N_4423);
and U9678 (N_9678,N_934,N_403);
or U9679 (N_9679,N_4375,N_1303);
nand U9680 (N_9680,N_927,N_4704);
nand U9681 (N_9681,N_4660,N_2122);
or U9682 (N_9682,N_473,N_3523);
nand U9683 (N_9683,N_4078,N_2983);
nor U9684 (N_9684,N_4822,N_1179);
nand U9685 (N_9685,N_1671,N_3445);
nor U9686 (N_9686,N_3929,N_1388);
or U9687 (N_9687,N_4814,N_1740);
and U9688 (N_9688,N_2956,N_4021);
and U9689 (N_9689,N_1867,N_3118);
nor U9690 (N_9690,N_1401,N_926);
nand U9691 (N_9691,N_4357,N_1717);
and U9692 (N_9692,N_2677,N_4082);
nor U9693 (N_9693,N_1873,N_3949);
and U9694 (N_9694,N_4925,N_1091);
and U9695 (N_9695,N_3383,N_3689);
nand U9696 (N_9696,N_3086,N_742);
nor U9697 (N_9697,N_3306,N_402);
nor U9698 (N_9698,N_1910,N_1330);
and U9699 (N_9699,N_4699,N_1865);
or U9700 (N_9700,N_3418,N_3051);
or U9701 (N_9701,N_2041,N_4922);
and U9702 (N_9702,N_3442,N_0);
or U9703 (N_9703,N_4746,N_1941);
or U9704 (N_9704,N_3433,N_3791);
nor U9705 (N_9705,N_1542,N_4039);
and U9706 (N_9706,N_3322,N_3568);
nand U9707 (N_9707,N_2787,N_213);
nand U9708 (N_9708,N_1462,N_2458);
nor U9709 (N_9709,N_580,N_4517);
or U9710 (N_9710,N_2483,N_1446);
nor U9711 (N_9711,N_989,N_1511);
or U9712 (N_9712,N_1910,N_3726);
and U9713 (N_9713,N_3380,N_674);
or U9714 (N_9714,N_1489,N_4002);
nor U9715 (N_9715,N_3575,N_2041);
and U9716 (N_9716,N_446,N_4212);
nand U9717 (N_9717,N_957,N_2980);
nor U9718 (N_9718,N_2473,N_133);
nand U9719 (N_9719,N_878,N_4966);
nand U9720 (N_9720,N_1264,N_1365);
nand U9721 (N_9721,N_4388,N_2671);
xor U9722 (N_9722,N_3207,N_576);
nand U9723 (N_9723,N_2541,N_825);
or U9724 (N_9724,N_2254,N_4144);
nor U9725 (N_9725,N_3824,N_2502);
or U9726 (N_9726,N_1725,N_285);
nor U9727 (N_9727,N_1406,N_2255);
or U9728 (N_9728,N_2230,N_1898);
nand U9729 (N_9729,N_692,N_489);
or U9730 (N_9730,N_756,N_4964);
nand U9731 (N_9731,N_2876,N_2396);
and U9732 (N_9732,N_1634,N_2356);
and U9733 (N_9733,N_3895,N_4935);
nor U9734 (N_9734,N_4669,N_431);
nor U9735 (N_9735,N_4101,N_1142);
and U9736 (N_9736,N_4461,N_4986);
nor U9737 (N_9737,N_2610,N_3954);
or U9738 (N_9738,N_2189,N_2445);
and U9739 (N_9739,N_2577,N_54);
nand U9740 (N_9740,N_4027,N_737);
or U9741 (N_9741,N_2023,N_2892);
or U9742 (N_9742,N_4500,N_3287);
and U9743 (N_9743,N_2292,N_2311);
and U9744 (N_9744,N_3205,N_3089);
nand U9745 (N_9745,N_3205,N_752);
nor U9746 (N_9746,N_4280,N_876);
nand U9747 (N_9747,N_2879,N_672);
or U9748 (N_9748,N_3368,N_1086);
and U9749 (N_9749,N_235,N_2139);
and U9750 (N_9750,N_1399,N_1486);
or U9751 (N_9751,N_1398,N_3526);
or U9752 (N_9752,N_2396,N_2080);
or U9753 (N_9753,N_1077,N_1461);
nor U9754 (N_9754,N_2650,N_3925);
nand U9755 (N_9755,N_2546,N_1676);
nor U9756 (N_9756,N_4043,N_4613);
nand U9757 (N_9757,N_2619,N_4639);
nand U9758 (N_9758,N_2527,N_1697);
or U9759 (N_9759,N_4215,N_2348);
and U9760 (N_9760,N_1468,N_3029);
nor U9761 (N_9761,N_4556,N_2042);
nor U9762 (N_9762,N_548,N_2995);
nor U9763 (N_9763,N_4857,N_2150);
or U9764 (N_9764,N_2772,N_537);
or U9765 (N_9765,N_4692,N_2322);
nand U9766 (N_9766,N_1232,N_2252);
or U9767 (N_9767,N_4699,N_2391);
nand U9768 (N_9768,N_1667,N_2730);
or U9769 (N_9769,N_4999,N_2802);
nor U9770 (N_9770,N_4899,N_2277);
nand U9771 (N_9771,N_693,N_4099);
nand U9772 (N_9772,N_1783,N_3120);
and U9773 (N_9773,N_2902,N_4765);
and U9774 (N_9774,N_2630,N_2248);
nand U9775 (N_9775,N_2588,N_3045);
and U9776 (N_9776,N_4385,N_4637);
and U9777 (N_9777,N_1938,N_146);
or U9778 (N_9778,N_2640,N_4452);
or U9779 (N_9779,N_907,N_2648);
and U9780 (N_9780,N_2517,N_2438);
nor U9781 (N_9781,N_3630,N_1200);
nor U9782 (N_9782,N_3462,N_4107);
nand U9783 (N_9783,N_2704,N_4841);
and U9784 (N_9784,N_279,N_329);
nand U9785 (N_9785,N_4234,N_3990);
nand U9786 (N_9786,N_1525,N_4496);
nor U9787 (N_9787,N_2260,N_2217);
nand U9788 (N_9788,N_2534,N_1714);
and U9789 (N_9789,N_3272,N_828);
nand U9790 (N_9790,N_4332,N_321);
nand U9791 (N_9791,N_3815,N_4752);
nor U9792 (N_9792,N_3203,N_2482);
nand U9793 (N_9793,N_579,N_1633);
or U9794 (N_9794,N_3331,N_3210);
nand U9795 (N_9795,N_1102,N_137);
and U9796 (N_9796,N_4854,N_3881);
nand U9797 (N_9797,N_3009,N_4072);
or U9798 (N_9798,N_1557,N_680);
and U9799 (N_9799,N_1278,N_254);
and U9800 (N_9800,N_4073,N_2869);
and U9801 (N_9801,N_2768,N_1162);
nor U9802 (N_9802,N_4817,N_4461);
or U9803 (N_9803,N_1598,N_1661);
nor U9804 (N_9804,N_3540,N_2617);
nor U9805 (N_9805,N_1689,N_1074);
and U9806 (N_9806,N_1456,N_3132);
or U9807 (N_9807,N_1149,N_1548);
or U9808 (N_9808,N_3839,N_859);
or U9809 (N_9809,N_2584,N_1071);
and U9810 (N_9810,N_4875,N_107);
or U9811 (N_9811,N_490,N_1336);
or U9812 (N_9812,N_4963,N_4495);
and U9813 (N_9813,N_1126,N_697);
nand U9814 (N_9814,N_4351,N_4049);
or U9815 (N_9815,N_3996,N_3870);
or U9816 (N_9816,N_3509,N_4529);
nor U9817 (N_9817,N_1241,N_1292);
nor U9818 (N_9818,N_1626,N_3767);
and U9819 (N_9819,N_4027,N_3855);
nor U9820 (N_9820,N_4522,N_1670);
nor U9821 (N_9821,N_415,N_2952);
and U9822 (N_9822,N_2695,N_3407);
and U9823 (N_9823,N_375,N_1906);
nand U9824 (N_9824,N_1063,N_3355);
nand U9825 (N_9825,N_3011,N_1107);
nor U9826 (N_9826,N_2063,N_4278);
nor U9827 (N_9827,N_3620,N_747);
nand U9828 (N_9828,N_3098,N_4531);
or U9829 (N_9829,N_882,N_876);
and U9830 (N_9830,N_2834,N_4498);
or U9831 (N_9831,N_4208,N_74);
or U9832 (N_9832,N_1209,N_3568);
and U9833 (N_9833,N_4550,N_4504);
or U9834 (N_9834,N_2359,N_722);
or U9835 (N_9835,N_1922,N_4814);
or U9836 (N_9836,N_1564,N_1797);
nor U9837 (N_9837,N_3059,N_2698);
or U9838 (N_9838,N_3217,N_1751);
and U9839 (N_9839,N_3271,N_3848);
or U9840 (N_9840,N_4168,N_3082);
nor U9841 (N_9841,N_1818,N_1251);
and U9842 (N_9842,N_3030,N_3322);
and U9843 (N_9843,N_4072,N_129);
nand U9844 (N_9844,N_212,N_2062);
nor U9845 (N_9845,N_2277,N_66);
nand U9846 (N_9846,N_1255,N_496);
nor U9847 (N_9847,N_2124,N_3581);
or U9848 (N_9848,N_3197,N_2187);
or U9849 (N_9849,N_3011,N_2446);
and U9850 (N_9850,N_2187,N_2362);
and U9851 (N_9851,N_1723,N_3256);
nand U9852 (N_9852,N_1789,N_1183);
nor U9853 (N_9853,N_923,N_1678);
nor U9854 (N_9854,N_2215,N_3914);
and U9855 (N_9855,N_2527,N_3998);
and U9856 (N_9856,N_3008,N_1633);
and U9857 (N_9857,N_245,N_2298);
nand U9858 (N_9858,N_317,N_3733);
or U9859 (N_9859,N_4335,N_932);
nand U9860 (N_9860,N_1963,N_4583);
or U9861 (N_9861,N_1268,N_166);
nor U9862 (N_9862,N_4239,N_2564);
or U9863 (N_9863,N_429,N_284);
nand U9864 (N_9864,N_2415,N_3311);
and U9865 (N_9865,N_3412,N_881);
and U9866 (N_9866,N_307,N_3880);
and U9867 (N_9867,N_370,N_3086);
and U9868 (N_9868,N_990,N_1212);
nor U9869 (N_9869,N_1213,N_2933);
nand U9870 (N_9870,N_4693,N_870);
nor U9871 (N_9871,N_2070,N_2053);
or U9872 (N_9872,N_2371,N_1298);
or U9873 (N_9873,N_2905,N_1259);
nor U9874 (N_9874,N_4732,N_3517);
xnor U9875 (N_9875,N_2494,N_2027);
nor U9876 (N_9876,N_4917,N_2841);
or U9877 (N_9877,N_1315,N_2924);
nand U9878 (N_9878,N_4411,N_2658);
and U9879 (N_9879,N_4977,N_1800);
nor U9880 (N_9880,N_4500,N_4185);
nand U9881 (N_9881,N_3579,N_2209);
nor U9882 (N_9882,N_3177,N_1899);
or U9883 (N_9883,N_2775,N_1463);
or U9884 (N_9884,N_2091,N_2565);
nand U9885 (N_9885,N_28,N_2457);
nand U9886 (N_9886,N_3481,N_2201);
nor U9887 (N_9887,N_3105,N_61);
nor U9888 (N_9888,N_575,N_876);
and U9889 (N_9889,N_1439,N_4345);
nor U9890 (N_9890,N_4341,N_4772);
nor U9891 (N_9891,N_3496,N_37);
or U9892 (N_9892,N_1878,N_624);
xnor U9893 (N_9893,N_4693,N_877);
or U9894 (N_9894,N_4296,N_2852);
nand U9895 (N_9895,N_417,N_573);
and U9896 (N_9896,N_3695,N_744);
nand U9897 (N_9897,N_1720,N_1243);
nand U9898 (N_9898,N_2286,N_2282);
or U9899 (N_9899,N_4168,N_2542);
nand U9900 (N_9900,N_4074,N_1386);
nor U9901 (N_9901,N_2105,N_1579);
and U9902 (N_9902,N_776,N_2215);
or U9903 (N_9903,N_53,N_4377);
nor U9904 (N_9904,N_4852,N_4388);
or U9905 (N_9905,N_3886,N_3804);
nand U9906 (N_9906,N_2493,N_2231);
nand U9907 (N_9907,N_2030,N_267);
or U9908 (N_9908,N_1823,N_3161);
nor U9909 (N_9909,N_3228,N_4818);
and U9910 (N_9910,N_4000,N_1588);
and U9911 (N_9911,N_338,N_4374);
or U9912 (N_9912,N_2693,N_4094);
and U9913 (N_9913,N_3376,N_1261);
or U9914 (N_9914,N_2201,N_4074);
nor U9915 (N_9915,N_4936,N_567);
or U9916 (N_9916,N_1050,N_4001);
nor U9917 (N_9917,N_3371,N_4555);
or U9918 (N_9918,N_1692,N_59);
or U9919 (N_9919,N_3233,N_1330);
nand U9920 (N_9920,N_3954,N_2338);
nand U9921 (N_9921,N_4230,N_489);
nor U9922 (N_9922,N_2010,N_130);
nor U9923 (N_9923,N_154,N_4453);
or U9924 (N_9924,N_406,N_2485);
nor U9925 (N_9925,N_1663,N_1020);
nand U9926 (N_9926,N_3893,N_4443);
or U9927 (N_9927,N_1941,N_4630);
and U9928 (N_9928,N_2224,N_1232);
and U9929 (N_9929,N_2112,N_3850);
nand U9930 (N_9930,N_177,N_3818);
nor U9931 (N_9931,N_4096,N_2637);
and U9932 (N_9932,N_4975,N_3458);
or U9933 (N_9933,N_705,N_4181);
nor U9934 (N_9934,N_3214,N_3372);
nor U9935 (N_9935,N_4930,N_186);
and U9936 (N_9936,N_1536,N_3342);
or U9937 (N_9937,N_3597,N_4801);
nand U9938 (N_9938,N_172,N_1636);
nor U9939 (N_9939,N_1184,N_2485);
and U9940 (N_9940,N_969,N_4404);
nor U9941 (N_9941,N_980,N_3634);
nor U9942 (N_9942,N_2817,N_666);
nor U9943 (N_9943,N_4570,N_3400);
nand U9944 (N_9944,N_921,N_2927);
and U9945 (N_9945,N_3092,N_2746);
nand U9946 (N_9946,N_464,N_1473);
nor U9947 (N_9947,N_1217,N_4066);
nand U9948 (N_9948,N_4234,N_1232);
or U9949 (N_9949,N_1306,N_4190);
and U9950 (N_9950,N_4916,N_818);
nand U9951 (N_9951,N_22,N_909);
or U9952 (N_9952,N_2994,N_3185);
nor U9953 (N_9953,N_2910,N_412);
or U9954 (N_9954,N_1365,N_184);
or U9955 (N_9955,N_1685,N_4416);
nor U9956 (N_9956,N_2203,N_4674);
nor U9957 (N_9957,N_3081,N_1674);
or U9958 (N_9958,N_4912,N_1782);
nand U9959 (N_9959,N_3068,N_2616);
nand U9960 (N_9960,N_2087,N_2230);
nor U9961 (N_9961,N_1429,N_2349);
and U9962 (N_9962,N_4812,N_8);
nand U9963 (N_9963,N_44,N_614);
or U9964 (N_9964,N_1295,N_3054);
and U9965 (N_9965,N_4858,N_4151);
or U9966 (N_9966,N_1248,N_3725);
or U9967 (N_9967,N_4176,N_3375);
and U9968 (N_9968,N_1338,N_4253);
nor U9969 (N_9969,N_771,N_1704);
nor U9970 (N_9970,N_4087,N_4663);
nand U9971 (N_9971,N_3548,N_2726);
or U9972 (N_9972,N_4725,N_3354);
and U9973 (N_9973,N_4495,N_2537);
nor U9974 (N_9974,N_3483,N_4255);
nor U9975 (N_9975,N_1360,N_2939);
nand U9976 (N_9976,N_4857,N_4667);
and U9977 (N_9977,N_4388,N_3413);
nand U9978 (N_9978,N_2201,N_3251);
nor U9979 (N_9979,N_4311,N_4723);
and U9980 (N_9980,N_4675,N_3237);
or U9981 (N_9981,N_1446,N_2219);
nor U9982 (N_9982,N_1482,N_4718);
or U9983 (N_9983,N_1744,N_3880);
xnor U9984 (N_9984,N_3362,N_542);
nor U9985 (N_9985,N_426,N_4905);
and U9986 (N_9986,N_2482,N_2644);
or U9987 (N_9987,N_3765,N_1407);
nand U9988 (N_9988,N_947,N_1441);
nor U9989 (N_9989,N_2833,N_3489);
and U9990 (N_9990,N_4971,N_3763);
or U9991 (N_9991,N_4502,N_193);
xor U9992 (N_9992,N_1592,N_906);
and U9993 (N_9993,N_2247,N_2885);
or U9994 (N_9994,N_2575,N_2040);
xnor U9995 (N_9995,N_3127,N_3162);
or U9996 (N_9996,N_1569,N_4442);
and U9997 (N_9997,N_3351,N_1240);
nor U9998 (N_9998,N_4619,N_1336);
nor U9999 (N_9999,N_1131,N_2991);
and U10000 (N_10000,N_9923,N_9494);
xor U10001 (N_10001,N_7235,N_8776);
nor U10002 (N_10002,N_8756,N_5833);
and U10003 (N_10003,N_8446,N_9193);
nor U10004 (N_10004,N_9035,N_9076);
and U10005 (N_10005,N_9134,N_6958);
or U10006 (N_10006,N_8634,N_5177);
nand U10007 (N_10007,N_6576,N_7975);
nand U10008 (N_10008,N_9855,N_6590);
xor U10009 (N_10009,N_7999,N_6179);
nand U10010 (N_10010,N_8622,N_7460);
nand U10011 (N_10011,N_5318,N_5386);
or U10012 (N_10012,N_8485,N_6905);
nand U10013 (N_10013,N_5630,N_8722);
nand U10014 (N_10014,N_5754,N_8917);
and U10015 (N_10015,N_9891,N_5108);
nor U10016 (N_10016,N_8124,N_8547);
nand U10017 (N_10017,N_9054,N_9295);
and U10018 (N_10018,N_8913,N_9612);
and U10019 (N_10019,N_5515,N_9146);
nor U10020 (N_10020,N_7545,N_6052);
nor U10021 (N_10021,N_9514,N_8886);
or U10022 (N_10022,N_5740,N_6318);
nand U10023 (N_10023,N_6066,N_7482);
nor U10024 (N_10024,N_5198,N_5942);
nor U10025 (N_10025,N_8516,N_7037);
or U10026 (N_10026,N_7862,N_7309);
or U10027 (N_10027,N_5076,N_9571);
nor U10028 (N_10028,N_8158,N_9633);
nor U10029 (N_10029,N_6860,N_6072);
nor U10030 (N_10030,N_9106,N_9277);
nor U10031 (N_10031,N_5300,N_5412);
or U10032 (N_10032,N_8080,N_8108);
nand U10033 (N_10033,N_6418,N_5557);
and U10034 (N_10034,N_6935,N_7569);
or U10035 (N_10035,N_9542,N_7288);
and U10036 (N_10036,N_8206,N_7636);
and U10037 (N_10037,N_7664,N_7003);
or U10038 (N_10038,N_6517,N_9750);
nor U10039 (N_10039,N_7702,N_7984);
and U10040 (N_10040,N_7479,N_6748);
or U10041 (N_10041,N_8298,N_7083);
or U10042 (N_10042,N_8311,N_8273);
nand U10043 (N_10043,N_5395,N_6080);
and U10044 (N_10044,N_6674,N_7819);
or U10045 (N_10045,N_6100,N_6839);
nor U10046 (N_10046,N_7938,N_7314);
or U10047 (N_10047,N_5968,N_9541);
or U10048 (N_10048,N_6106,N_8340);
nor U10049 (N_10049,N_9977,N_5438);
nor U10050 (N_10050,N_9397,N_5542);
nand U10051 (N_10051,N_8774,N_7867);
nor U10052 (N_10052,N_6127,N_6622);
or U10053 (N_10053,N_7173,N_5350);
nand U10054 (N_10054,N_7944,N_8971);
or U10055 (N_10055,N_7737,N_8543);
or U10056 (N_10056,N_7480,N_6594);
nand U10057 (N_10057,N_7035,N_7802);
nor U10058 (N_10058,N_8493,N_6280);
nor U10059 (N_10059,N_8805,N_8810);
and U10060 (N_10060,N_8209,N_9584);
and U10061 (N_10061,N_5577,N_7259);
nor U10062 (N_10062,N_7162,N_5582);
or U10063 (N_10063,N_7603,N_9298);
and U10064 (N_10064,N_8180,N_5232);
or U10065 (N_10065,N_8847,N_9203);
nor U10066 (N_10066,N_9044,N_9816);
nand U10067 (N_10067,N_8746,N_9671);
and U10068 (N_10068,N_8051,N_7074);
nor U10069 (N_10069,N_5421,N_6286);
nor U10070 (N_10070,N_5396,N_7231);
and U10071 (N_10071,N_9903,N_8266);
or U10072 (N_10072,N_8175,N_8222);
nand U10073 (N_10073,N_7658,N_8085);
and U10074 (N_10074,N_7902,N_5358);
nor U10075 (N_10075,N_9704,N_8713);
nand U10076 (N_10076,N_5408,N_6481);
and U10077 (N_10077,N_9254,N_8379);
and U10078 (N_10078,N_9045,N_8574);
nand U10079 (N_10079,N_7156,N_5510);
and U10080 (N_10080,N_5612,N_9937);
and U10081 (N_10081,N_5948,N_7567);
nand U10082 (N_10082,N_5399,N_9930);
nor U10083 (N_10083,N_6420,N_7222);
nor U10084 (N_10084,N_8058,N_6146);
and U10085 (N_10085,N_8252,N_9257);
nand U10086 (N_10086,N_8658,N_9466);
nor U10087 (N_10087,N_8787,N_9646);
and U10088 (N_10088,N_6483,N_6200);
nand U10089 (N_10089,N_7853,N_5082);
xnor U10090 (N_10090,N_6413,N_8223);
nor U10091 (N_10091,N_5261,N_9491);
or U10092 (N_10092,N_5727,N_5956);
or U10093 (N_10093,N_5661,N_7697);
nand U10094 (N_10094,N_8940,N_9345);
nand U10095 (N_10095,N_5138,N_5877);
and U10096 (N_10096,N_6714,N_5698);
nor U10097 (N_10097,N_6643,N_6512);
or U10098 (N_10098,N_7986,N_8237);
nand U10099 (N_10099,N_8136,N_8808);
or U10100 (N_10100,N_9877,N_5394);
and U10101 (N_10101,N_5625,N_9673);
nand U10102 (N_10102,N_7331,N_9757);
and U10103 (N_10103,N_8681,N_9288);
or U10104 (N_10104,N_6181,N_9115);
nor U10105 (N_10105,N_7315,N_6513);
and U10106 (N_10106,N_5519,N_9033);
nor U10107 (N_10107,N_7191,N_9668);
and U10108 (N_10108,N_7143,N_7170);
nand U10109 (N_10109,N_7544,N_8921);
xnor U10110 (N_10110,N_6299,N_8545);
or U10111 (N_10111,N_8985,N_9702);
nand U10112 (N_10112,N_6957,N_7209);
nor U10113 (N_10113,N_6550,N_9524);
or U10114 (N_10114,N_5590,N_7561);
or U10115 (N_10115,N_9791,N_6793);
nand U10116 (N_10116,N_5616,N_6601);
and U10117 (N_10117,N_5157,N_7915);
or U10118 (N_10118,N_5458,N_8075);
xor U10119 (N_10119,N_9404,N_8164);
or U10120 (N_10120,N_9970,N_9438);
or U10121 (N_10121,N_9934,N_6419);
and U10122 (N_10122,N_8523,N_7145);
nand U10123 (N_10123,N_7564,N_7889);
nor U10124 (N_10124,N_5331,N_5656);
nor U10125 (N_10125,N_9927,N_6995);
nand U10126 (N_10126,N_8304,N_5613);
nor U10127 (N_10127,N_8229,N_6068);
or U10128 (N_10128,N_6692,N_6983);
or U10129 (N_10129,N_8844,N_7007);
and U10130 (N_10130,N_7735,N_7001);
nand U10131 (N_10131,N_8149,N_5959);
nand U10132 (N_10132,N_5141,N_6619);
or U10133 (N_10133,N_7733,N_6926);
or U10134 (N_10134,N_5233,N_9174);
xor U10135 (N_10135,N_8081,N_8306);
nand U10136 (N_10136,N_8624,N_8026);
and U10137 (N_10137,N_7097,N_5192);
nand U10138 (N_10138,N_5549,N_6242);
and U10139 (N_10139,N_7112,N_8123);
nand U10140 (N_10140,N_9963,N_7842);
nand U10141 (N_10141,N_6224,N_9627);
nand U10142 (N_10142,N_5869,N_5212);
nor U10143 (N_10143,N_9716,N_6219);
and U10144 (N_10144,N_9332,N_6487);
and U10145 (N_10145,N_8356,N_8877);
nand U10146 (N_10146,N_8505,N_5724);
or U10147 (N_10147,N_5855,N_7640);
nand U10148 (N_10148,N_6821,N_6085);
and U10149 (N_10149,N_7776,N_6159);
and U10150 (N_10150,N_7106,N_8278);
or U10151 (N_10151,N_5801,N_9748);
nand U10152 (N_10152,N_5791,N_6193);
nand U10153 (N_10153,N_6621,N_8344);
nor U10154 (N_10154,N_7738,N_7005);
nor U10155 (N_10155,N_6618,N_7048);
nor U10156 (N_10156,N_8183,N_6469);
nand U10157 (N_10157,N_8529,N_5814);
nand U10158 (N_10158,N_9302,N_8062);
nand U10159 (N_10159,N_5788,N_6685);
nand U10160 (N_10160,N_5923,N_7255);
and U10161 (N_10161,N_5606,N_8064);
and U10162 (N_10162,N_6940,N_7413);
and U10163 (N_10163,N_9499,N_6694);
nor U10164 (N_10164,N_7916,N_7855);
nor U10165 (N_10165,N_7403,N_5132);
nand U10166 (N_10166,N_5250,N_9645);
nand U10167 (N_10167,N_8996,N_8795);
and U10168 (N_10168,N_7124,N_9608);
or U10169 (N_10169,N_8739,N_7472);
and U10170 (N_10170,N_6073,N_7087);
nand U10171 (N_10171,N_7948,N_5351);
and U10172 (N_10172,N_9261,N_8839);
nor U10173 (N_10173,N_7877,N_5707);
nor U10174 (N_10174,N_6447,N_9710);
nor U10175 (N_10175,N_8841,N_6352);
nand U10176 (N_10176,N_9082,N_6817);
nand U10177 (N_10177,N_7570,N_8439);
or U10178 (N_10178,N_7505,N_6400);
nor U10179 (N_10179,N_8637,N_6741);
or U10180 (N_10180,N_7650,N_7192);
or U10181 (N_10181,N_8046,N_8797);
and U10182 (N_10182,N_6520,N_8038);
and U10183 (N_10183,N_8927,N_7411);
or U10184 (N_10184,N_7681,N_7562);
nand U10185 (N_10185,N_9619,N_9249);
nor U10186 (N_10186,N_8732,N_8151);
and U10187 (N_10187,N_6051,N_5890);
or U10188 (N_10188,N_5185,N_9041);
or U10189 (N_10189,N_9961,N_6906);
nand U10190 (N_10190,N_6638,N_7942);
and U10191 (N_10191,N_8358,N_9665);
and U10192 (N_10192,N_5713,N_8381);
or U10193 (N_10193,N_8185,N_7150);
nor U10194 (N_10194,N_7523,N_9316);
nor U10195 (N_10195,N_9911,N_6644);
nand U10196 (N_10196,N_6546,N_9049);
nand U10197 (N_10197,N_6007,N_7987);
and U10198 (N_10198,N_6291,N_6366);
or U10199 (N_10199,N_5634,N_9053);
and U10200 (N_10200,N_5560,N_7361);
nand U10201 (N_10201,N_5011,N_7746);
nand U10202 (N_10202,N_8753,N_8845);
or U10203 (N_10203,N_9897,N_7438);
and U10204 (N_10204,N_6067,N_6683);
or U10205 (N_10205,N_6728,N_7201);
nor U10206 (N_10206,N_7581,N_9511);
nand U10207 (N_10207,N_8626,N_8250);
nand U10208 (N_10208,N_9264,N_6696);
nor U10209 (N_10209,N_7149,N_7435);
or U10210 (N_10210,N_7560,N_5312);
nor U10211 (N_10211,N_6202,N_5187);
and U10212 (N_10212,N_7270,N_8320);
and U10213 (N_10213,N_6723,N_6320);
and U10214 (N_10214,N_8672,N_7256);
nand U10215 (N_10215,N_6473,N_6165);
nor U10216 (N_10216,N_6725,N_7522);
nor U10217 (N_10217,N_6573,N_7787);
or U10218 (N_10218,N_9490,N_8950);
nor U10219 (N_10219,N_6604,N_8727);
or U10220 (N_10220,N_9197,N_6515);
nand U10221 (N_10221,N_7366,N_7506);
and U10222 (N_10222,N_5035,N_9539);
nor U10223 (N_10223,N_6902,N_9628);
and U10224 (N_10224,N_9084,N_7196);
or U10225 (N_10225,N_9370,N_9160);
nand U10226 (N_10226,N_6650,N_7417);
and U10227 (N_10227,N_9538,N_8550);
or U10228 (N_10228,N_9536,N_9521);
nand U10229 (N_10229,N_8508,N_8212);
or U10230 (N_10230,N_8494,N_6697);
nand U10231 (N_10231,N_6084,N_9582);
nor U10232 (N_10232,N_8625,N_7386);
or U10233 (N_10233,N_9417,N_5057);
nand U10234 (N_10234,N_8090,N_6936);
or U10235 (N_10235,N_6844,N_9530);
nand U10236 (N_10236,N_8554,N_8862);
nor U10237 (N_10237,N_5061,N_8415);
nor U10238 (N_10238,N_5089,N_6474);
nand U10239 (N_10239,N_5165,N_8919);
nor U10240 (N_10240,N_7293,N_6059);
or U10241 (N_10241,N_8734,N_6975);
nand U10242 (N_10242,N_5517,N_9075);
or U10243 (N_10243,N_9950,N_8486);
nand U10244 (N_10244,N_7897,N_9094);
nor U10245 (N_10245,N_9532,N_5059);
nand U10246 (N_10246,N_5533,N_6246);
nand U10247 (N_10247,N_8730,N_6880);
and U10248 (N_10248,N_5790,N_6614);
or U10249 (N_10249,N_7054,N_8643);
nor U10250 (N_10250,N_6810,N_7212);
and U10251 (N_10251,N_7613,N_8002);
nand U10252 (N_10252,N_5360,N_8050);
nand U10253 (N_10253,N_6626,N_6430);
and U10254 (N_10254,N_7113,N_5337);
or U10255 (N_10255,N_7009,N_7794);
nand U10256 (N_10256,N_5739,N_9730);
or U10257 (N_10257,N_9371,N_9064);
and U10258 (N_10258,N_5882,N_7120);
or U10259 (N_10259,N_7701,N_7558);
nand U10260 (N_10260,N_8611,N_6260);
nand U10261 (N_10261,N_9284,N_9439);
or U10262 (N_10262,N_8608,N_8113);
and U10263 (N_10263,N_7084,N_7808);
and U10264 (N_10264,N_8382,N_9005);
nor U10265 (N_10265,N_5040,N_6651);
nand U10266 (N_10266,N_5868,N_6130);
or U10267 (N_10267,N_9293,N_5984);
and U10268 (N_10268,N_7696,N_7800);
nand U10269 (N_10269,N_7548,N_7719);
nor U10270 (N_10270,N_7950,N_8308);
nor U10271 (N_10271,N_5960,N_9794);
nand U10272 (N_10272,N_9269,N_6225);
nor U10273 (N_10273,N_5704,N_6412);
nor U10274 (N_10274,N_7806,N_8587);
nor U10275 (N_10275,N_7684,N_5503);
nor U10276 (N_10276,N_8213,N_7549);
nand U10277 (N_10277,N_6682,N_9548);
nor U10278 (N_10278,N_6433,N_5988);
or U10279 (N_10279,N_7940,N_6319);
nand U10280 (N_10280,N_5274,N_8986);
and U10281 (N_10281,N_5531,N_7273);
or U10282 (N_10282,N_8639,N_8366);
nor U10283 (N_10283,N_9935,N_5334);
nor U10284 (N_10284,N_7898,N_6999);
or U10285 (N_10285,N_9596,N_8191);
nor U10286 (N_10286,N_7881,N_5512);
or U10287 (N_10287,N_8775,N_6139);
nand U10288 (N_10288,N_8453,N_8657);
nand U10289 (N_10289,N_5328,N_7875);
nand U10290 (N_10290,N_5211,N_6768);
and U10291 (N_10291,N_8910,N_8897);
nor U10292 (N_10292,N_8821,N_8436);
and U10293 (N_10293,N_7577,N_5899);
and U10294 (N_10294,N_6230,N_9344);
or U10295 (N_10295,N_8980,N_9839);
nor U10296 (N_10296,N_5993,N_6443);
and U10297 (N_10297,N_6209,N_5400);
nor U10298 (N_10298,N_5505,N_6307);
or U10299 (N_10299,N_8895,N_6060);
nand U10300 (N_10300,N_7789,N_8208);
nor U10301 (N_10301,N_5292,N_9881);
or U10302 (N_10302,N_5675,N_8771);
or U10303 (N_10303,N_6415,N_9159);
and U10304 (N_10304,N_5842,N_9800);
nor U10305 (N_10305,N_7531,N_5467);
nand U10306 (N_10306,N_6216,N_8408);
nand U10307 (N_10307,N_7409,N_9485);
nor U10308 (N_10308,N_5017,N_8735);
nand U10309 (N_10309,N_7611,N_6727);
or U10310 (N_10310,N_5348,N_8331);
nor U10311 (N_10311,N_9544,N_9003);
nor U10312 (N_10312,N_6029,N_5856);
or U10313 (N_10313,N_8025,N_8563);
nor U10314 (N_10314,N_5474,N_9402);
and U10315 (N_10315,N_9823,N_5402);
nor U10316 (N_10316,N_9523,N_7739);
nor U10317 (N_10317,N_8434,N_6018);
nor U10318 (N_10318,N_9932,N_8872);
and U10319 (N_10319,N_7704,N_7785);
nand U10320 (N_10320,N_6608,N_8219);
and U10321 (N_10321,N_9270,N_5784);
nor U10322 (N_10322,N_5246,N_9330);
or U10323 (N_10323,N_6251,N_8948);
and U10324 (N_10324,N_5841,N_9820);
and U10325 (N_10325,N_5139,N_9365);
and U10326 (N_10326,N_8642,N_5056);
or U10327 (N_10327,N_6630,N_6093);
nand U10328 (N_10328,N_9440,N_6972);
nand U10329 (N_10329,N_9243,N_7248);
nand U10330 (N_10330,N_8215,N_9576);
or U10331 (N_10331,N_9941,N_7547);
and U10332 (N_10332,N_6323,N_6409);
and U10333 (N_10333,N_5589,N_5593);
nor U10334 (N_10334,N_7706,N_8021);
nor U10335 (N_10335,N_7781,N_6993);
nor U10336 (N_10336,N_6452,N_5084);
nor U10337 (N_10337,N_5673,N_9692);
nand U10338 (N_10338,N_5973,N_7540);
or U10339 (N_10339,N_9395,N_6462);
nand U10340 (N_10340,N_6663,N_9423);
or U10341 (N_10341,N_5172,N_8930);
or U10342 (N_10342,N_6110,N_7878);
and U10343 (N_10343,N_7262,N_7014);
or U10344 (N_10344,N_7765,N_7555);
and U10345 (N_10345,N_9662,N_5946);
nand U10346 (N_10346,N_8375,N_8603);
and U10347 (N_10347,N_6348,N_7216);
and U10348 (N_10348,N_7410,N_5663);
and U10349 (N_10349,N_6990,N_9593);
or U10350 (N_10350,N_5794,N_7043);
nor U10351 (N_10351,N_9981,N_7982);
nor U10352 (N_10352,N_6818,N_5189);
nand U10353 (N_10353,N_5155,N_6949);
and U10354 (N_10354,N_8460,N_5540);
nor U10355 (N_10355,N_6729,N_7864);
nand U10356 (N_10356,N_7217,N_6317);
nor U10357 (N_10357,N_6392,N_9387);
and U10358 (N_10358,N_5140,N_8506);
nand U10359 (N_10359,N_5924,N_9091);
or U10360 (N_10360,N_7047,N_7179);
nand U10361 (N_10361,N_7020,N_5701);
nand U10362 (N_10362,N_5094,N_9926);
nand U10363 (N_10363,N_5870,N_7408);
and U10364 (N_10364,N_5283,N_6680);
or U10365 (N_10365,N_8429,N_6647);
nor U10366 (N_10366,N_8748,N_6706);
nand U10367 (N_10367,N_5525,N_9217);
nor U10368 (N_10368,N_9508,N_9207);
nand U10369 (N_10369,N_5369,N_7233);
nor U10370 (N_10370,N_7187,N_8777);
nand U10371 (N_10371,N_9079,N_8678);
nand U10372 (N_10372,N_7851,N_5119);
and U10373 (N_10373,N_6541,N_5532);
nand U10374 (N_10374,N_6509,N_9376);
nand U10375 (N_10375,N_9756,N_9696);
or U10376 (N_10376,N_7670,N_9434);
and U10377 (N_10377,N_6340,N_5846);
and U10378 (N_10378,N_9443,N_8095);
nor U10379 (N_10379,N_7443,N_7724);
and U10380 (N_10380,N_7762,N_9598);
xnor U10381 (N_10381,N_6411,N_9418);
and U10382 (N_10382,N_9265,N_9537);
or U10383 (N_10383,N_7763,N_8096);
nand U10384 (N_10384,N_7773,N_7535);
nand U10385 (N_10385,N_9066,N_7065);
and U10386 (N_10386,N_6569,N_7379);
nor U10387 (N_10387,N_6107,N_9113);
and U10388 (N_10388,N_9385,N_5278);
or U10389 (N_10389,N_6221,N_7079);
nand U10390 (N_10390,N_8758,N_5898);
nor U10391 (N_10391,N_6916,N_6386);
nor U10392 (N_10392,N_9830,N_8918);
nor U10393 (N_10393,N_9367,N_9414);
nor U10394 (N_10394,N_7356,N_6354);
nor U10395 (N_10395,N_6721,N_9343);
or U10396 (N_10396,N_8196,N_5535);
nand U10397 (N_10397,N_5863,N_5690);
nor U10398 (N_10398,N_8673,N_9703);
or U10399 (N_10399,N_8894,N_9336);
or U10400 (N_10400,N_9516,N_9080);
nor U10401 (N_10401,N_7101,N_6794);
nand U10402 (N_10402,N_9708,N_8182);
nor U10403 (N_10403,N_9606,N_9683);
nand U10404 (N_10404,N_7610,N_7537);
or U10405 (N_10405,N_6804,N_8314);
nand U10406 (N_10406,N_5390,N_7638);
nand U10407 (N_10407,N_5181,N_7213);
and U10408 (N_10408,N_8056,N_8251);
nor U10409 (N_10409,N_5928,N_5494);
nor U10410 (N_10410,N_6171,N_5915);
and U10411 (N_10411,N_6823,N_8765);
nand U10412 (N_10412,N_8707,N_5149);
nand U10413 (N_10413,N_5125,N_8107);
nor U10414 (N_10414,N_5464,N_9303);
or U10415 (N_10415,N_7521,N_5257);
nand U10416 (N_10416,N_6873,N_7936);
or U10417 (N_10417,N_6557,N_6013);
and U10418 (N_10418,N_8231,N_5776);
nor U10419 (N_10419,N_8034,N_8285);
nor U10420 (N_10420,N_9314,N_9520);
nand U10421 (N_10421,N_7458,N_6244);
and U10422 (N_10422,N_5805,N_5415);
and U10423 (N_10423,N_7520,N_8109);
or U10424 (N_10424,N_5156,N_5581);
nor U10425 (N_10425,N_8702,N_6910);
nand U10426 (N_10426,N_6668,N_5897);
nand U10427 (N_10427,N_9359,N_5619);
nor U10428 (N_10428,N_8833,N_9181);
or U10429 (N_10429,N_6887,N_9862);
nor U10430 (N_10430,N_5476,N_5439);
or U10431 (N_10431,N_5290,N_9420);
and U10432 (N_10432,N_6351,N_8135);
and U10433 (N_10433,N_9019,N_5072);
and U10434 (N_10434,N_5977,N_7990);
nor U10435 (N_10435,N_5470,N_6489);
nand U10436 (N_10436,N_6846,N_6233);
or U10437 (N_10437,N_7755,N_7727);
nand U10438 (N_10438,N_8651,N_7375);
and U10439 (N_10439,N_7418,N_6207);
nand U10440 (N_10440,N_5629,N_9459);
nand U10441 (N_10441,N_5038,N_7809);
nor U10442 (N_10442,N_6813,N_5340);
or U10443 (N_10443,N_6893,N_5669);
nand U10444 (N_10444,N_9728,N_5566);
nand U10445 (N_10445,N_5252,N_7596);
and U10446 (N_10446,N_7780,N_7903);
nand U10447 (N_10447,N_5325,N_7637);
or U10448 (N_10448,N_5098,N_7011);
nor U10449 (N_10449,N_7130,N_6820);
or U10450 (N_10450,N_5559,N_8165);
nand U10451 (N_10451,N_5910,N_6010);
and U10452 (N_10452,N_5743,N_5873);
or U10453 (N_10453,N_9654,N_8991);
xor U10454 (N_10454,N_6395,N_6878);
xor U10455 (N_10455,N_8271,N_8843);
nor U10456 (N_10456,N_8849,N_9108);
and U10457 (N_10457,N_9992,N_9380);
or U10458 (N_10458,N_6459,N_6273);
and U10459 (N_10459,N_8300,N_5883);
nor U10460 (N_10460,N_8110,N_7714);
nand U10461 (N_10461,N_7393,N_6020);
nor U10462 (N_10462,N_7451,N_5168);
nor U10463 (N_10463,N_8332,N_9004);
nand U10464 (N_10464,N_6756,N_7110);
or U10465 (N_10465,N_7931,N_7578);
nand U10466 (N_10466,N_7516,N_9859);
and U10467 (N_10467,N_5806,N_7811);
and U10468 (N_10468,N_9462,N_5384);
nand U10469 (N_10469,N_8201,N_8924);
nor U10470 (N_10470,N_7376,N_7499);
xor U10471 (N_10471,N_5808,N_7153);
and U10472 (N_10472,N_8683,N_8518);
nor U10473 (N_10473,N_6114,N_9153);
and U10474 (N_10474,N_9695,N_9630);
nand U10475 (N_10475,N_6258,N_7164);
or U10476 (N_10476,N_8176,N_9947);
nor U10477 (N_10477,N_6210,N_9954);
nand U10478 (N_10478,N_9586,N_7978);
nor U10479 (N_10479,N_7236,N_8526);
nor U10480 (N_10480,N_8613,N_6710);
nand U10481 (N_10481,N_5311,N_8449);
nor U10482 (N_10482,N_8261,N_5664);
and U10483 (N_10483,N_5809,N_5551);
nor U10484 (N_10484,N_8537,N_5618);
nor U10485 (N_10485,N_7707,N_5498);
nand U10486 (N_10486,N_7527,N_8536);
nand U10487 (N_10487,N_6488,N_9413);
or U10488 (N_10488,N_6777,N_7383);
nor U10489 (N_10489,N_6406,N_5881);
nor U10490 (N_10490,N_9095,N_5699);
nand U10491 (N_10491,N_5120,N_8593);
or U10492 (N_10492,N_7943,N_7350);
nor U10493 (N_10493,N_7258,N_8166);
or U10494 (N_10494,N_8424,N_8586);
or U10495 (N_10495,N_9856,N_9894);
or U10496 (N_10496,N_9635,N_6426);
nand U10497 (N_10497,N_8906,N_6002);
nand U10498 (N_10498,N_8852,N_6095);
and U10499 (N_10499,N_9872,N_8994);
or U10500 (N_10500,N_6915,N_8478);
nand U10501 (N_10501,N_5005,N_8083);
nand U10502 (N_10502,N_7859,N_7140);
nor U10503 (N_10503,N_6428,N_5989);
and U10504 (N_10504,N_6482,N_8579);
or U10505 (N_10505,N_6437,N_6397);
nor U10506 (N_10506,N_8091,N_9611);
nor U10507 (N_10507,N_9427,N_9237);
nand U10508 (N_10508,N_9623,N_9141);
or U10509 (N_10509,N_8708,N_9317);
and U10510 (N_10510,N_9943,N_9018);
nand U10511 (N_10511,N_6190,N_8482);
nor U10512 (N_10512,N_7817,N_7988);
xor U10513 (N_10513,N_5456,N_8115);
nand U10514 (N_10514,N_5570,N_9451);
and U10515 (N_10515,N_5832,N_9906);
xnor U10516 (N_10516,N_5703,N_7952);
and U10517 (N_10517,N_6627,N_9682);
or U10518 (N_10518,N_8635,N_8670);
and U10519 (N_10519,N_6889,N_9472);
and U10520 (N_10520,N_9476,N_6329);
and U10521 (N_10521,N_9813,N_9198);
or U10522 (N_10522,N_7364,N_6276);
and U10523 (N_10523,N_5054,N_8671);
nand U10524 (N_10524,N_9346,N_7325);
nor U10525 (N_10525,N_9808,N_6241);
nor U10526 (N_10526,N_5448,N_8343);
nand U10527 (N_10527,N_9067,N_8920);
nand U10528 (N_10528,N_7805,N_9874);
and U10529 (N_10529,N_6065,N_7454);
nand U10530 (N_10530,N_8294,N_5151);
and U10531 (N_10531,N_6253,N_5296);
or U10532 (N_10532,N_5117,N_9915);
nand U10533 (N_10533,N_5326,N_8905);
and U10534 (N_10534,N_7654,N_5939);
and U10535 (N_10535,N_7094,N_8772);
and U10536 (N_10536,N_7512,N_7951);
and U10537 (N_10537,N_5289,N_6301);
nand U10538 (N_10538,N_6290,N_9090);
nor U10539 (N_10539,N_7373,N_7059);
or U10540 (N_10540,N_7252,N_8339);
and U10541 (N_10541,N_5501,N_6503);
nand U10542 (N_10542,N_8692,N_5916);
or U10543 (N_10543,N_5904,N_9761);
and U10544 (N_10544,N_6929,N_8577);
nand U10545 (N_10545,N_5095,N_5452);
and U10546 (N_10546,N_7147,N_9484);
nor U10547 (N_10547,N_8901,N_6096);
nor U10548 (N_10548,N_9917,N_9362);
nor U10549 (N_10549,N_6575,N_5262);
nor U10550 (N_10550,N_7088,N_7363);
nor U10551 (N_10551,N_8401,N_8409);
or U10552 (N_10552,N_5478,N_9194);
nand U10553 (N_10553,N_6042,N_9426);
and U10554 (N_10554,N_7599,N_9123);
nand U10555 (N_10555,N_6152,N_6533);
and U10556 (N_10556,N_6671,N_8481);
or U10557 (N_10557,N_5689,N_8428);
and U10558 (N_10558,N_7374,N_7671);
and U10559 (N_10559,N_9470,N_6522);
or U10560 (N_10560,N_8057,N_9858);
and U10561 (N_10561,N_7462,N_6799);
and U10562 (N_10562,N_6504,N_8316);
and U10563 (N_10563,N_9251,N_5398);
nand U10564 (N_10564,N_5614,N_8441);
or U10565 (N_10565,N_5096,N_8630);
or U10566 (N_10566,N_9342,N_8641);
nor U10567 (N_10567,N_7461,N_5774);
or U10568 (N_10568,N_7426,N_9910);
nor U10569 (N_10569,N_9121,N_8893);
and U10570 (N_10570,N_6876,N_8814);
nand U10571 (N_10571,N_5720,N_7144);
nor U10572 (N_10572,N_7207,N_8187);
nand U10573 (N_10573,N_8818,N_5875);
nor U10574 (N_10574,N_5203,N_5305);
nand U10575 (N_10575,N_9191,N_6427);
nor U10576 (N_10576,N_8342,N_7899);
nor U10577 (N_10577,N_5541,N_8380);
nor U10578 (N_10578,N_8615,N_8988);
nor U10579 (N_10579,N_9510,N_8174);
and U10580 (N_10580,N_8662,N_7378);
nor U10581 (N_10581,N_9711,N_5162);
nor U10582 (N_10582,N_5787,N_7556);
and U10583 (N_10583,N_7703,N_7830);
nor U10584 (N_10584,N_9964,N_8891);
or U10585 (N_10585,N_5935,N_7991);
nand U10586 (N_10586,N_7989,N_8378);
and U10587 (N_10587,N_5217,N_6776);
nand U10588 (N_10588,N_8568,N_5816);
or U10589 (N_10589,N_5216,N_9789);
nand U10590 (N_10590,N_5712,N_6123);
nor U10591 (N_10591,N_6491,N_9805);
nor U10592 (N_10592,N_5838,N_9037);
nand U10593 (N_10593,N_9211,N_9384);
nor U10594 (N_10594,N_8071,N_5433);
nor U10595 (N_10595,N_9238,N_5555);
nand U10596 (N_10596,N_5886,N_5355);
nor U10597 (N_10597,N_8301,N_5810);
and U10598 (N_10598,N_6024,N_9364);
nor U10599 (N_10599,N_9998,N_6864);
xor U10600 (N_10600,N_6841,N_6800);
and U10601 (N_10601,N_8817,N_7471);
xor U10602 (N_10602,N_7463,N_7188);
xor U10603 (N_10603,N_7085,N_8602);
nand U10604 (N_10604,N_6559,N_8747);
nand U10605 (N_10605,N_5765,N_8770);
nand U10606 (N_10606,N_9827,N_9133);
nor U10607 (N_10607,N_7056,N_8721);
or U10608 (N_10608,N_6494,N_5769);
nand U10609 (N_10609,N_5976,N_6480);
and U10610 (N_10610,N_7313,N_7849);
nor U10611 (N_10611,N_8011,N_5163);
nor U10612 (N_10612,N_5909,N_6151);
and U10613 (N_10613,N_5428,N_5969);
or U10614 (N_10614,N_8575,N_9222);
nand U10615 (N_10615,N_8793,N_9129);
and U10616 (N_10616,N_6510,N_8495);
or U10617 (N_10617,N_5323,N_8357);
nand U10618 (N_10618,N_6595,N_9172);
nor U10619 (N_10619,N_6635,N_8426);
and U10620 (N_10620,N_9152,N_9622);
nor U10621 (N_10621,N_9252,N_6587);
and U10622 (N_10622,N_5996,N_9899);
or U10623 (N_10623,N_6035,N_6370);
or U10624 (N_10624,N_9241,N_8766);
nor U10625 (N_10625,N_6250,N_9766);
nor U10626 (N_10626,N_8835,N_7491);
nand U10627 (N_10627,N_6008,N_8445);
nand U10628 (N_10628,N_7370,N_6167);
and U10629 (N_10629,N_8937,N_9636);
or U10630 (N_10630,N_8100,N_7204);
and U10631 (N_10631,N_5580,N_9112);
and U10632 (N_10632,N_8389,N_9187);
nor U10633 (N_10633,N_5012,N_5357);
nand U10634 (N_10634,N_9672,N_6750);
nand U10635 (N_10635,N_6271,N_6620);
or U10636 (N_10636,N_7291,N_8978);
or U10637 (N_10637,N_5224,N_8618);
nor U10638 (N_10638,N_8871,N_9286);
or U10639 (N_10639,N_5564,N_5708);
and U10640 (N_10640,N_5496,N_6888);
or U10641 (N_10641,N_5425,N_6477);
or U10642 (N_10642,N_5714,N_5640);
or U10643 (N_10643,N_6537,N_6153);
nor U10644 (N_10644,N_9052,N_7563);
nand U10645 (N_10645,N_7066,N_9901);
or U10646 (N_10646,N_5941,N_6911);
nand U10647 (N_10647,N_8292,N_6819);
and U10648 (N_10648,N_7717,N_8022);
nor U10649 (N_10649,N_7937,N_9560);
nor U10650 (N_10650,N_8472,N_5142);
or U10651 (N_10651,N_9880,N_9256);
or U10652 (N_10652,N_7301,N_9898);
and U10653 (N_10653,N_8558,N_6956);
nor U10654 (N_10654,N_6709,N_9594);
nand U10655 (N_10655,N_6111,N_5925);
and U10656 (N_10656,N_6341,N_8858);
nor U10657 (N_10657,N_8598,N_9546);
and U10658 (N_10658,N_9833,N_6726);
and U10659 (N_10659,N_6965,N_9400);
nand U10660 (N_10660,N_7911,N_8355);
or U10661 (N_10661,N_9762,N_8228);
nand U10662 (N_10662,N_7169,N_6616);
nand U10663 (N_10663,N_8682,N_5330);
or U10664 (N_10664,N_5087,N_9613);
and U10665 (N_10665,N_9506,N_9739);
nor U10666 (N_10666,N_7385,N_9587);
or U10667 (N_10667,N_7260,N_9535);
and U10668 (N_10668,N_7496,N_7642);
nand U10669 (N_10669,N_7312,N_7396);
and U10670 (N_10670,N_8923,N_7025);
and U10671 (N_10671,N_7300,N_5136);
and U10672 (N_10672,N_8277,N_9392);
nor U10673 (N_10673,N_5196,N_7655);
nor U10674 (N_10674,N_5235,N_8812);
or U10675 (N_10675,N_7530,N_9111);
nor U10676 (N_10676,N_6865,N_9040);
nand U10677 (N_10677,N_9460,N_9481);
or U10678 (N_10678,N_9273,N_7021);
nand U10679 (N_10679,N_5892,N_5597);
nor U10680 (N_10680,N_9834,N_7041);
nand U10681 (N_10681,N_7039,N_5050);
nor U10682 (N_10682,N_6105,N_9562);
and U10683 (N_10683,N_7352,N_8719);
nand U10684 (N_10684,N_7711,N_6529);
or U10685 (N_10685,N_5818,N_9580);
or U10686 (N_10686,N_6897,N_5450);
or U10687 (N_10687,N_8741,N_5756);
or U10688 (N_10688,N_5554,N_7298);
nor U10689 (N_10689,N_7134,N_5081);
nand U10690 (N_10690,N_7353,N_6252);
nand U10691 (N_10691,N_8003,N_8195);
nand U10692 (N_10692,N_9088,N_9700);
and U10693 (N_10693,N_9745,N_7804);
nor U10694 (N_10694,N_6201,N_7218);
nand U10695 (N_10695,N_9431,N_5100);
or U10696 (N_10696,N_6539,N_5049);
nor U10697 (N_10697,N_7509,N_9185);
and U10698 (N_10698,N_6334,N_9908);
nand U10699 (N_10699,N_7810,N_5671);
nor U10700 (N_10700,N_9647,N_9436);
or U10701 (N_10701,N_8496,N_6641);
nor U10702 (N_10702,N_5729,N_9245);
nor U10703 (N_10703,N_9691,N_6538);
xor U10704 (N_10704,N_5778,N_8525);
and U10705 (N_10705,N_6755,N_5459);
and U10706 (N_10706,N_6545,N_5972);
nor U10707 (N_10707,N_8763,N_5302);
and U10708 (N_10708,N_7713,N_5697);
and U10709 (N_10709,N_5397,N_7928);
and U10710 (N_10710,N_7813,N_8589);
nand U10711 (N_10711,N_5295,N_7181);
or U10712 (N_10712,N_5840,N_6194);
nand U10713 (N_10713,N_5105,N_7401);
nand U10714 (N_10714,N_5380,N_5702);
nand U10715 (N_10715,N_9182,N_6454);
and U10716 (N_10716,N_7333,N_9381);
nor U10717 (N_10717,N_7442,N_7686);
nand U10718 (N_10718,N_8863,N_7276);
and U10719 (N_10719,N_9006,N_7573);
nor U10720 (N_10720,N_8726,N_8942);
and U10721 (N_10721,N_9792,N_5986);
and U10722 (N_10722,N_9713,N_8049);
or U10723 (N_10723,N_5123,N_7691);
and U10724 (N_10724,N_6868,N_7620);
and U10725 (N_10725,N_7661,N_6581);
and U10726 (N_10726,N_5711,N_5905);
nor U10727 (N_10727,N_7500,N_8995);
nor U10728 (N_10728,N_6277,N_9024);
or U10729 (N_10729,N_5491,N_7985);
or U10730 (N_10730,N_9030,N_8138);
nor U10731 (N_10731,N_6746,N_8870);
or U10732 (N_10732,N_6112,N_9824);
or U10733 (N_10733,N_6184,N_6585);
and U10734 (N_10734,N_6087,N_9565);
nand U10735 (N_10735,N_9637,N_5468);
nand U10736 (N_10736,N_6180,N_5407);
nor U10737 (N_10737,N_7533,N_9883);
or U10738 (N_10738,N_6056,N_6379);
nor U10739 (N_10739,N_8504,N_5159);
and U10740 (N_10740,N_7160,N_7771);
and U10741 (N_10741,N_7138,N_5241);
nor U10742 (N_10742,N_9738,N_7306);
or U10743 (N_10743,N_5521,N_6816);
or U10744 (N_10744,N_5116,N_9916);
or U10745 (N_10745,N_8235,N_8789);
nand U10746 (N_10746,N_9811,N_8477);
nor U10747 (N_10747,N_8674,N_5143);
and U10748 (N_10748,N_8580,N_9271);
and U10749 (N_10749,N_5426,N_8404);
and U10750 (N_10750,N_5277,N_7422);
nor U10751 (N_10751,N_5324,N_7337);
and U10752 (N_10752,N_8666,N_8904);
or U10753 (N_10753,N_9577,N_6044);
nand U10754 (N_10754,N_8302,N_8599);
nor U10755 (N_10755,N_8029,N_5586);
nor U10756 (N_10756,N_8470,N_9085);
and U10757 (N_10757,N_5365,N_5565);
nor U10758 (N_10758,N_5522,N_8153);
or U10759 (N_10759,N_9784,N_8520);
or U10760 (N_10760,N_5387,N_6667);
nand U10761 (N_10761,N_7096,N_8498);
or U10762 (N_10762,N_7816,N_7269);
or U10763 (N_10763,N_5624,N_7692);
and U10764 (N_10764,N_8647,N_8655);
nor U10765 (N_10765,N_6649,N_7914);
and U10766 (N_10766,N_7183,N_7660);
nor U10767 (N_10767,N_7447,N_9802);
nand U10768 (N_10768,N_9373,N_9719);
nand U10769 (N_10769,N_7559,N_7504);
nor U10770 (N_10770,N_5601,N_6182);
or U10771 (N_10771,N_9806,N_6971);
and U10772 (N_10772,N_5029,N_8245);
nor U10773 (N_10773,N_7172,N_9027);
and U10774 (N_10774,N_9324,N_7240);
nand U10775 (N_10775,N_8510,N_9688);
and U10776 (N_10776,N_5075,N_8112);
and U10777 (N_10777,N_7121,N_7604);
nor U10778 (N_10778,N_8488,N_6363);
nor U10779 (N_10779,N_7423,N_9588);
nor U10780 (N_10780,N_6178,N_8287);
or U10781 (N_10781,N_6467,N_8898);
or U10782 (N_10782,N_8804,N_8933);
and U10783 (N_10783,N_8167,N_5173);
or U10784 (N_10784,N_9764,N_8855);
or U10785 (N_10785,N_7525,N_8570);
nand U10786 (N_10786,N_9643,N_7060);
nor U10787 (N_10787,N_9837,N_5020);
or U10788 (N_10788,N_9305,N_7111);
nand U10789 (N_10789,N_7225,N_8976);
nor U10790 (N_10790,N_5569,N_5353);
nor U10791 (N_10791,N_7861,N_6872);
nor U10792 (N_10792,N_5599,N_9493);
or U10793 (N_10793,N_7489,N_8473);
nor U10794 (N_10794,N_6083,N_7964);
or U10795 (N_10795,N_6145,N_6941);
nand U10796 (N_10796,N_6312,N_7334);
xor U10797 (N_10797,N_6851,N_7641);
and U10798 (N_10798,N_9667,N_9478);
nor U10799 (N_10799,N_7814,N_8307);
nand U10800 (N_10800,N_9326,N_5546);
nand U10801 (N_10801,N_7687,N_7646);
nor U10802 (N_10802,N_5286,N_6362);
nand U10803 (N_10803,N_6061,N_8715);
and U10804 (N_10804,N_5513,N_8761);
and U10805 (N_10805,N_5636,N_6955);
nand U10806 (N_10806,N_5273,N_5696);
or U10807 (N_10807,N_5214,N_6837);
nor U10808 (N_10808,N_9658,N_8257);
and U10809 (N_10809,N_5025,N_7245);
or U10810 (N_10810,N_5733,N_5763);
nand U10811 (N_10811,N_7807,N_5186);
nand U10812 (N_10812,N_7507,N_5970);
or U10813 (N_10813,N_9602,N_6045);
and U10814 (N_10814,N_6571,N_7912);
nor U10815 (N_10815,N_5596,N_5160);
or U10816 (N_10816,N_7167,N_9008);
and U10817 (N_10817,N_5280,N_7710);
or U10818 (N_10818,N_9363,N_9852);
nand U10819 (N_10819,N_7767,N_7343);
nor U10820 (N_10820,N_5998,N_6040);
nor U10821 (N_10821,N_8116,N_7792);
or U10822 (N_10822,N_6939,N_6380);
or U10823 (N_10823,N_7529,N_7466);
xor U10824 (N_10824,N_6414,N_9483);
or U10825 (N_10825,N_6154,N_9215);
nor U10826 (N_10826,N_6828,N_6490);
nand U10827 (N_10827,N_5556,N_5639);
nor U10828 (N_10828,N_5230,N_8604);
nor U10829 (N_10829,N_6215,N_7682);
or U10830 (N_10830,N_7685,N_9664);
nor U10831 (N_10831,N_9442,N_6733);
and U10832 (N_10832,N_7329,N_8295);
nor U10833 (N_10833,N_6325,N_6542);
xor U10834 (N_10834,N_5850,N_8450);
nor U10835 (N_10835,N_6774,N_5553);
and U10836 (N_10836,N_7788,N_5480);
or U10837 (N_10837,N_9341,N_9338);
nor U10838 (N_10838,N_7223,N_7972);
or U10839 (N_10839,N_6531,N_9656);
and U10840 (N_10840,N_8929,N_7033);
nand U10841 (N_10841,N_7431,N_7148);
nand U10842 (N_10842,N_7514,N_9177);
and U10843 (N_10843,N_6032,N_5822);
nor U10844 (N_10844,N_8319,N_9617);
and U10845 (N_10845,N_8422,N_7070);
nand U10846 (N_10846,N_8646,N_6740);
and U10847 (N_10847,N_5176,N_9154);
and U10848 (N_10848,N_7107,N_5294);
or U10849 (N_10849,N_6997,N_5845);
nand U10850 (N_10850,N_7061,N_9465);
nand U10851 (N_10851,N_8769,N_7541);
or U10852 (N_10852,N_8609,N_8539);
and U10853 (N_10853,N_7042,N_7672);
and U10854 (N_10854,N_5288,N_9253);
or U10855 (N_10855,N_5796,N_5041);
or U10856 (N_10856,N_6764,N_5411);
and U10857 (N_10857,N_5179,N_8867);
and U10858 (N_10858,N_6701,N_8132);
or U10859 (N_10859,N_6724,N_5991);
and U10860 (N_10860,N_5502,N_9777);
or U10861 (N_10861,N_9218,N_7405);
or U10862 (N_10862,N_5583,N_6012);
nor U10863 (N_10863,N_7184,N_7016);
xor U10864 (N_10864,N_5950,N_5034);
nor U10865 (N_10865,N_5306,N_5341);
and U10866 (N_10866,N_7566,N_5455);
nor U10867 (N_10867,N_7663,N_8665);
and U10868 (N_10868,N_7015,N_8802);
nor U10869 (N_10869,N_6925,N_7860);
nand U10870 (N_10870,N_8427,N_5088);
and U10871 (N_10871,N_9969,N_8289);
nor U10872 (N_10872,N_7917,N_7801);
nor U10873 (N_10873,N_9534,N_9543);
nor U10874 (N_10874,N_9743,N_9157);
nand U10875 (N_10875,N_8086,N_8189);
nand U10876 (N_10876,N_6500,N_9996);
and U10877 (N_10877,N_8997,N_6185);
or U10878 (N_10878,N_7073,N_6247);
and U10879 (N_10879,N_9931,N_8616);
and U10880 (N_10880,N_6206,N_6381);
nand U10881 (N_10881,N_5975,N_7310);
and U10882 (N_10882,N_7090,N_5249);
nand U10883 (N_10883,N_6992,N_7920);
and U10884 (N_10884,N_9403,N_7645);
and U10885 (N_10885,N_6333,N_5537);
or U10886 (N_10886,N_8455,N_8564);
nand U10887 (N_10887,N_5723,N_8027);
nand U10888 (N_10888,N_8888,N_5807);
nand U10889 (N_10889,N_6234,N_6498);
nor U10890 (N_10890,N_9214,N_5401);
nand U10891 (N_10891,N_9686,N_5874);
xnor U10892 (N_10892,N_7494,N_9479);
or U10893 (N_10893,N_8521,N_7032);
nor U10894 (N_10894,N_8267,N_6014);
nor U10895 (N_10895,N_7302,N_9829);
and U10896 (N_10896,N_7297,N_9940);
or U10897 (N_10897,N_8963,N_5872);
nor U10898 (N_10898,N_5943,N_8490);
or U10899 (N_10899,N_9117,N_8966);
or U10900 (N_10900,N_9583,N_7764);
nor U10901 (N_10901,N_9818,N_6753);
and U10902 (N_10902,N_6578,N_6640);
and U10903 (N_10903,N_8561,N_5558);
nand U10904 (N_10904,N_6231,N_7414);
or U10905 (N_10905,N_5338,N_5248);
nand U10906 (N_10906,N_5304,N_5834);
nor U10907 (N_10907,N_5709,N_7323);
nand U10908 (N_10908,N_5770,N_7568);
and U10909 (N_10909,N_8806,N_5062);
or U10910 (N_10910,N_8199,N_7576);
nor U10911 (N_10911,N_5710,N_8784);
nor U10912 (N_10912,N_5259,N_8573);
or U10913 (N_10913,N_5240,N_9731);
and U10914 (N_10914,N_9232,N_9225);
nand U10915 (N_10915,N_6690,N_6326);
and U10916 (N_10916,N_8418,N_5687);
and U10917 (N_10917,N_6584,N_5490);
nand U10918 (N_10918,N_6497,N_5715);
or U10919 (N_10919,N_8479,N_7526);
nand U10920 (N_10920,N_9169,N_8535);
or U10921 (N_10921,N_8644,N_7475);
or U10922 (N_10922,N_7441,N_9896);
nand U10923 (N_10923,N_8111,N_6164);
nand U10924 (N_10924,N_8262,N_8465);
nor U10925 (N_10925,N_6786,N_9863);
nand U10926 (N_10926,N_5037,N_9983);
nand U10927 (N_10927,N_6293,N_6403);
and U10928 (N_10928,N_6212,N_7863);
nor U10929 (N_10929,N_6855,N_8048);
and U10930 (N_10930,N_7215,N_5004);
nand U10931 (N_10931,N_6946,N_6170);
and U10932 (N_10932,N_7468,N_5067);
and U10933 (N_10933,N_5462,N_8040);
or U10934 (N_10934,N_9575,N_7866);
and U10935 (N_10935,N_7769,N_5717);
and U10936 (N_10936,N_9718,N_6305);
and U10937 (N_10937,N_7824,N_9055);
nand U10938 (N_10938,N_9393,N_6795);
nor U10939 (N_10939,N_6797,N_5668);
or U10940 (N_10940,N_5051,N_9659);
nand U10941 (N_10941,N_8031,N_9437);
nand U10942 (N_10942,N_9482,N_6023);
and U10943 (N_10943,N_7137,N_6009);
or U10944 (N_10944,N_8423,N_6505);
nand U10945 (N_10945,N_5244,N_8259);
nor U10946 (N_10946,N_6806,N_5819);
nand U10947 (N_10947,N_8204,N_7818);
or U10948 (N_10948,N_6658,N_6176);
nand U10949 (N_10949,N_9137,N_9333);
nor U10950 (N_10950,N_6356,N_7029);
and U10951 (N_10951,N_9101,N_5388);
or U10952 (N_10952,N_7709,N_5219);
nand U10953 (N_10953,N_7367,N_8416);
or U10954 (N_10954,N_5995,N_7913);
nand U10955 (N_10955,N_7839,N_6217);
nor U10956 (N_10956,N_9036,N_6248);
nor U10957 (N_10957,N_7071,N_8881);
or U10958 (N_10958,N_8992,N_8947);
or U10959 (N_10959,N_7062,N_6552);
or U10960 (N_10960,N_6205,N_9771);
or U10961 (N_10961,N_8363,N_6775);
and U10962 (N_10962,N_5644,N_7141);
nor U10963 (N_10963,N_6432,N_8704);
nor U10964 (N_10964,N_6673,N_6960);
and U10965 (N_10965,N_5799,N_8128);
nor U10966 (N_10966,N_7159,N_9853);
and U10967 (N_10967,N_5753,N_5180);
and U10968 (N_10968,N_7498,N_5048);
nand U10969 (N_10969,N_9828,N_9760);
nor U10970 (N_10970,N_6648,N_6142);
or U10971 (N_10971,N_8288,N_5003);
nor U10972 (N_10972,N_9875,N_9058);
and U10973 (N_10973,N_9212,N_9201);
or U10974 (N_10974,N_6016,N_8661);
and U10975 (N_10975,N_8464,N_9751);
or U10976 (N_10976,N_8955,N_6809);
and U10977 (N_10977,N_9405,N_6458);
and U10978 (N_10978,N_7519,N_7619);
or U10979 (N_10979,N_7883,N_6937);
or U10980 (N_10980,N_5371,N_6254);
nor U10981 (N_10981,N_9838,N_6313);
or U10982 (N_10982,N_7688,N_8480);
nand U10983 (N_10983,N_8467,N_7621);
and U10984 (N_10984,N_6460,N_8152);
and U10985 (N_10985,N_6556,N_9292);
or U10986 (N_10986,N_6470,N_5803);
nor U10987 (N_10987,N_9569,N_5681);
or U10988 (N_10988,N_6530,N_6544);
or U10989 (N_10989,N_5405,N_8668);
nand U10990 (N_10990,N_7341,N_5958);
and U10991 (N_10991,N_6423,N_9631);
nor U10992 (N_10992,N_6589,N_6101);
nand U10993 (N_10993,N_8399,N_8544);
or U10994 (N_10994,N_5880,N_8501);
or U10995 (N_10995,N_9072,N_9723);
and U10996 (N_10996,N_8885,N_8016);
and U10997 (N_10997,N_5033,N_7019);
nor U10998 (N_10998,N_5130,N_6814);
nor U10999 (N_10999,N_6144,N_6404);
or U11000 (N_11000,N_8232,N_7299);
nand U11001 (N_11001,N_6967,N_6987);
nand U11002 (N_11002,N_6607,N_6834);
and U11003 (N_11003,N_6731,N_8813);
and U11004 (N_11004,N_9379,N_8338);
and U11005 (N_11005,N_9463,N_8612);
or U11006 (N_11006,N_9919,N_5101);
nor U11007 (N_11007,N_8264,N_7268);
nor U11008 (N_11008,N_8752,N_8840);
and U11009 (N_11009,N_5114,N_9002);
nand U11010 (N_11010,N_7552,N_6850);
nor U11011 (N_11011,N_7616,N_6006);
and U11012 (N_11012,N_8979,N_6173);
nand U11013 (N_11013,N_5069,N_5889);
and U11014 (N_11014,N_7133,N_7254);
nand U11015 (N_11015,N_7617,N_7338);
nor U11016 (N_11016,N_9502,N_5144);
or U11017 (N_11017,N_5750,N_8054);
or U11018 (N_11018,N_6953,N_8414);
and U11019 (N_11019,N_8519,N_5103);
or U11020 (N_11020,N_7241,N_6986);
nor U11021 (N_11021,N_9509,N_6543);
and U11022 (N_11022,N_8968,N_6036);
or U11023 (N_11023,N_5013,N_9933);
or U11024 (N_11024,N_5609,N_6295);
nand U11025 (N_11025,N_9790,N_9164);
nor U11026 (N_11026,N_7630,N_6448);
or U11027 (N_11027,N_6579,N_7354);
and U11028 (N_11028,N_8458,N_8860);
and U11029 (N_11029,N_9390,N_7407);
or U11030 (N_11030,N_6331,N_5682);
or U11031 (N_11031,N_7892,N_5666);
nand U11032 (N_11032,N_8440,N_9322);
or U11033 (N_11033,N_9353,N_8336);
or U11034 (N_11034,N_9461,N_7456);
or U11035 (N_11035,N_8951,N_8638);
or U11036 (N_11036,N_7190,N_6677);
and U11037 (N_11037,N_8044,N_9325);
nand U11038 (N_11038,N_9455,N_8636);
nor U11039 (N_11039,N_8181,N_8367);
and U11040 (N_11040,N_8911,N_9287);
nand U11041 (N_11041,N_9976,N_5738);
nand U11042 (N_11042,N_6166,N_9107);
nand U11043 (N_11043,N_8347,N_5285);
nor U11044 (N_11044,N_7469,N_5786);
and U11045 (N_11045,N_7828,N_9720);
nor U11046 (N_11046,N_8744,N_5479);
nor U11047 (N_11047,N_5449,N_5830);
nor U11048 (N_11048,N_8354,N_6296);
nand U11049 (N_11049,N_7797,N_5745);
or U11050 (N_11050,N_5766,N_5097);
nand U11051 (N_11051,N_8082,N_7834);
nor U11052 (N_11052,N_5732,N_5779);
nand U11053 (N_11053,N_7885,N_6199);
nand U11054 (N_11054,N_5914,N_6842);
xor U11055 (N_11055,N_5487,N_9677);
or U11056 (N_11056,N_6711,N_8648);
nand U11057 (N_11057,N_6950,N_9732);
nor U11058 (N_11058,N_8263,N_7970);
and U11059 (N_11059,N_9590,N_9999);
and U11060 (N_11060,N_7871,N_9301);
nand U11061 (N_11061,N_7266,N_8142);
nand U11062 (N_11062,N_8313,N_9737);
and U11063 (N_11063,N_6996,N_7588);
or U11064 (N_11064,N_8555,N_5633);
nand U11065 (N_11065,N_8178,N_9009);
and U11066 (N_11066,N_5073,N_8412);
and U11067 (N_11067,N_7927,N_7840);
or U11068 (N_11068,N_8827,N_5432);
and U11069 (N_11069,N_6698,N_6718);
nand U11070 (N_11070,N_5206,N_7659);
nor U11071 (N_11071,N_5955,N_6033);
nor U11072 (N_11072,N_5451,N_7332);
nand U11073 (N_11073,N_6963,N_5167);
nand U11074 (N_11074,N_8605,N_6297);
nor U11075 (N_11075,N_8764,N_6952);
nand U11076 (N_11076,N_8869,N_8977);
nand U11077 (N_11077,N_7715,N_8729);
or U11078 (N_11078,N_7959,N_6526);
nand U11079 (N_11079,N_6330,N_6133);
and U11080 (N_11080,N_9350,N_9229);
and U11081 (N_11081,N_8974,N_5587);
nor U11082 (N_11082,N_6597,N_8497);
or U11083 (N_11083,N_9616,N_6289);
or U11084 (N_11084,N_5982,N_5392);
and U11085 (N_11085,N_8689,N_9724);
or U11086 (N_11086,N_7053,N_7832);
and U11087 (N_11087,N_5523,N_7966);
nor U11088 (N_11088,N_9871,N_5764);
nand U11089 (N_11089,N_7751,N_7893);
or U11090 (N_11090,N_8394,N_9446);
and U11091 (N_11091,N_5674,N_6285);
and U11092 (N_11092,N_8359,N_9339);
nor U11093 (N_11093,N_6464,N_5315);
nand U11094 (N_11094,N_9528,N_5637);
nand U11095 (N_11095,N_7846,N_9895);
nand U11096 (N_11096,N_7285,N_9938);
or U11097 (N_11097,N_9801,N_6003);
nor U11098 (N_11098,N_5383,N_9032);
or U11099 (N_11099,N_5045,N_6877);
nor U11100 (N_11100,N_7459,N_6198);
nor U11101 (N_11101,N_6004,N_9953);
nand U11102 (N_11102,N_6693,N_8850);
nor U11103 (N_11103,N_9522,N_8017);
nand U11104 (N_11104,N_6303,N_5308);
nand U11105 (N_11105,N_6847,N_6349);
or U11106 (N_11106,N_7812,N_8964);
or U11107 (N_11107,N_9955,N_6966);
nand U11108 (N_11108,N_7993,N_8330);
nor U11109 (N_11109,N_6624,N_8310);
or U11110 (N_11110,N_9653,N_9966);
and U11111 (N_11111,N_7958,N_8785);
nand U11112 (N_11112,N_8385,N_8868);
and U11113 (N_11113,N_7072,N_5813);
nor U11114 (N_11114,N_8015,N_5831);
nand U11115 (N_11115,N_9624,N_6760);
nand U11116 (N_11116,N_8788,N_8392);
or U11117 (N_11117,N_6866,N_5298);
nor U11118 (N_11118,N_6315,N_7271);
nand U11119 (N_11119,N_6646,N_6962);
nand U11120 (N_11120,N_9957,N_7077);
and U11121 (N_11121,N_6121,N_9722);
nand U11122 (N_11122,N_8581,N_7953);
nor U11123 (N_11123,N_5070,N_6665);
nor U11124 (N_11124,N_7592,N_6565);
nor U11125 (N_11125,N_7208,N_8507);
or U11126 (N_11126,N_8061,N_9394);
nand U11127 (N_11127,N_7058,N_6075);
and U11128 (N_11128,N_5594,N_8596);
and U11129 (N_11129,N_9864,N_8258);
and U11130 (N_11130,N_6449,N_8837);
xnor U11131 (N_11131,N_9701,N_9914);
or U11132 (N_11132,N_9726,N_6377);
nor U11133 (N_11133,N_7036,N_7565);
or U11134 (N_11134,N_5752,N_9774);
nor U11135 (N_11135,N_6985,N_7869);
and U11136 (N_11136,N_9334,N_9697);
nor U11137 (N_11137,N_9092,N_5952);
nor U11138 (N_11138,N_9487,N_6735);
nand U11139 (N_11139,N_5166,N_8786);
nor U11140 (N_11140,N_9236,N_8282);
and U11141 (N_11141,N_6269,N_7852);
and U11142 (N_11142,N_7239,N_8349);
nand U11143 (N_11143,N_9625,N_9050);
nand U11144 (N_11144,N_6717,N_8621);
or U11145 (N_11145,N_7318,N_6302);
nand U11146 (N_11146,N_5603,N_5797);
or U11147 (N_11147,N_5234,N_5620);
or U11148 (N_11148,N_9266,N_8072);
and U11149 (N_11149,N_5659,N_6540);
nor U11150 (N_11150,N_9213,N_6979);
and U11151 (N_11151,N_5860,N_8965);
nand U11152 (N_11152,N_6183,N_8967);
nand U11153 (N_11153,N_5231,N_5228);
or U11154 (N_11154,N_5936,N_7608);
and U11155 (N_11155,N_7146,N_6832);
nor U11156 (N_11156,N_7126,N_5536);
or U11157 (N_11157,N_5333,N_8463);
nand U11158 (N_11158,N_7104,N_6506);
nand U11159 (N_11159,N_5858,N_8148);
nand U11160 (N_11160,N_9161,N_6431);
nor U11161 (N_11161,N_6298,N_9907);
nor U11162 (N_11162,N_7955,N_9268);
nor U11163 (N_11163,N_5043,N_5303);
or U11164 (N_11164,N_6948,N_6854);
nand U11165 (N_11165,N_6082,N_9531);
or U11166 (N_11166,N_8820,N_7976);
nor U11167 (N_11167,N_5651,N_8177);
and U11168 (N_11168,N_8782,N_9226);
xor U11169 (N_11169,N_6603,N_8122);
nor U11170 (N_11170,N_5251,N_7622);
nor U11171 (N_11171,N_8532,N_8312);
nand U11172 (N_11172,N_5475,N_5339);
nand U11173 (N_11173,N_8631,N_6399);
nor U11174 (N_11174,N_9729,N_5635);
or U11175 (N_11175,N_5178,N_7380);
and U11176 (N_11176,N_7752,N_9500);
and U11177 (N_11177,N_9978,N_6989);
and U11178 (N_11178,N_8101,N_8864);
or U11179 (N_11179,N_6339,N_6328);
nand U11180 (N_11180,N_5255,N_9515);
or U11181 (N_11181,N_7585,N_5992);
and U11182 (N_11182,N_5653,N_7394);
nor U11183 (N_11183,N_9096,N_8139);
nor U11184 (N_11184,N_9779,N_8990);
nand U11185 (N_11185,N_8104,N_8010);
or U11186 (N_11186,N_7495,N_5483);
or U11187 (N_11187,N_6120,N_7843);
nor U11188 (N_11188,N_8369,N_9803);
and U11189 (N_11189,N_5684,N_8315);
nor U11190 (N_11190,N_9661,N_8691);
and U11191 (N_11191,N_5660,N_7712);
and U11192 (N_11192,N_5828,N_8296);
and U11193 (N_11193,N_6451,N_9202);
or U11194 (N_11194,N_8945,N_9308);
and U11195 (N_11195,N_7197,N_9401);
nand U11196 (N_11196,N_6197,N_9860);
or U11197 (N_11197,N_5245,N_8710);
nand U11198 (N_11198,N_9031,N_8407);
or U11199 (N_11199,N_7052,N_6628);
nor U11200 (N_11200,N_5321,N_8368);
nand U11201 (N_11201,N_5042,N_9347);
nor U11202 (N_11202,N_5484,N_6263);
nand U11203 (N_11203,N_8815,N_5239);
nor U11204 (N_11204,N_9567,N_5751);
nor U11205 (N_11205,N_6562,N_5563);
and U11206 (N_11206,N_7669,N_7593);
and U11207 (N_11207,N_6852,N_6108);
and U11208 (N_11208,N_9651,N_7006);
nand U11209 (N_11209,N_9210,N_9679);
nor U11210 (N_11210,N_5893,N_5194);
and U11211 (N_11211,N_8623,N_8703);
and U11212 (N_11212,N_5945,N_5847);
and U11213 (N_11213,N_7135,N_8376);
nand U11214 (N_11214,N_6308,N_7647);
and U11215 (N_11215,N_9289,N_5127);
and U11216 (N_11216,N_9512,N_6904);
or U11217 (N_11217,N_9985,N_9707);
or U11218 (N_11218,N_6732,N_7369);
nand U11219 (N_11219,N_6090,N_8693);
nor U11220 (N_11220,N_6332,N_9550);
and U11221 (N_11221,N_9660,N_9960);
and U11222 (N_11222,N_8799,N_5256);
or U11223 (N_11223,N_9131,N_8249);
nand U11224 (N_11224,N_8926,N_7010);
or U11225 (N_11225,N_6446,N_5592);
or U11226 (N_11226,N_9698,N_9351);
and U11227 (N_11227,N_5667,N_8317);
or U11228 (N_11228,N_9984,N_6822);
nor U11229 (N_11229,N_8254,N_9070);
nand U11230 (N_11230,N_6688,N_9398);
nand U11231 (N_11231,N_6656,N_8226);
and U11232 (N_11232,N_6678,N_8514);
nor U11233 (N_11233,N_5862,N_9621);
or U11234 (N_11234,N_5431,N_5678);
and U11235 (N_11235,N_5099,N_8973);
or U11236 (N_11236,N_6240,N_8192);
nor U11237 (N_11237,N_5430,N_7510);
nor U11238 (N_11238,N_8972,N_8120);
or U11239 (N_11239,N_9282,N_6261);
xor U11240 (N_11240,N_9735,N_8400);
nor U11241 (N_11241,N_5627,N_9162);
or U11242 (N_11242,N_7177,N_9183);
nor U11243 (N_11243,N_7068,N_7997);
nand U11244 (N_11244,N_7742,N_9549);
nand U11245 (N_11245,N_6679,N_7923);
nand U11246 (N_11246,N_9233,N_8781);
nand U11247 (N_11247,N_5226,N_6278);
nor U11248 (N_11248,N_8438,N_8890);
or U11249 (N_11249,N_9821,N_8633);
nor U11250 (N_11250,N_9391,N_9819);
or U11251 (N_11251,N_8084,N_9997);
xnor U11252 (N_11252,N_8395,N_8341);
or U11253 (N_11253,N_7890,N_9093);
nand U11254 (N_11254,N_5281,N_6612);
or U11255 (N_11255,N_5588,N_9150);
nand U11256 (N_11256,N_9629,N_9850);
nor U11257 (N_11257,N_9545,N_9518);
and U11258 (N_11258,N_7844,N_9166);
nor U11259 (N_11259,N_9951,N_5418);
nor U11260 (N_11260,N_5762,N_9415);
and U11261 (N_11261,N_5865,N_6922);
nand U11262 (N_11262,N_7481,N_6662);
or U11263 (N_11263,N_6162,N_9320);
and U11264 (N_11264,N_6064,N_6281);
or U11265 (N_11265,N_6754,N_6335);
nor U11266 (N_11266,N_9601,N_5672);
and U11267 (N_11267,N_6577,N_8912);
nand U11268 (N_11268,N_5036,N_8738);
nand U11269 (N_11269,N_9069,N_8907);
nand U11270 (N_11270,N_7995,N_8328);
and U11271 (N_11271,N_9492,N_5372);
or U11272 (N_11272,N_7234,N_5481);
nor U11273 (N_11273,N_9815,N_7109);
nand U11274 (N_11274,N_5820,N_5363);
nand U11275 (N_11275,N_6687,N_6238);
nor U11276 (N_11276,N_6959,N_7579);
nor U11277 (N_11277,N_8687,N_5896);
or U11278 (N_11278,N_9020,N_5742);
and U11279 (N_11279,N_8896,N_8607);
and U11280 (N_11280,N_8653,N_6582);
nand U11281 (N_11281,N_7265,N_7511);
nand U11282 (N_11282,N_7732,N_8946);
and U11283 (N_11283,N_7591,N_7249);
nor U11284 (N_11284,N_5864,N_6306);
or U11285 (N_11285,N_7793,N_5578);
nor U11286 (N_11286,N_5906,N_7790);
nand U11287 (N_11287,N_5662,N_6444);
nor U11288 (N_11288,N_7674,N_7440);
nor U11289 (N_11289,N_5052,N_5477);
or U11290 (N_11290,N_6028,N_8822);
nand U11291 (N_11291,N_8419,N_9189);
nand U11292 (N_11292,N_7497,N_6829);
or U11293 (N_11293,N_7689,N_8773);
or U11294 (N_11294,N_7322,N_5679);
nand U11295 (N_11295,N_5547,N_9657);
nor U11296 (N_11296,N_6593,N_9776);
or U11297 (N_11297,N_7030,N_8242);
or U11298 (N_11298,N_5963,N_7433);
nor U11299 (N_11299,N_6907,N_8383);
nand U11300 (N_11300,N_7368,N_7633);
or U11301 (N_11301,N_8716,N_5344);
or U11302 (N_11302,N_8700,N_6267);
and U11303 (N_11303,N_8155,N_8437);
and U11304 (N_11304,N_8179,N_7662);
or U11305 (N_11305,N_5113,N_7895);
nor U11306 (N_11306,N_6081,N_8922);
nand U11307 (N_11307,N_6079,N_8350);
nor U11308 (N_11308,N_7831,N_9958);
nand U11309 (N_11309,N_9578,N_8754);
nor U11310 (N_11310,N_5210,N_6324);
nand U11311 (N_11311,N_9842,N_6213);
and U11312 (N_11312,N_5393,N_5965);
and U11313 (N_11313,N_9591,N_5891);
nor U11314 (N_11314,N_5471,N_5953);
and U11315 (N_11315,N_9204,N_5913);
or U11316 (N_11316,N_6981,N_8361);
nor U11317 (N_11317,N_6988,N_5243);
and U11318 (N_11318,N_8411,N_5327);
nor U11319 (N_11319,N_8873,N_9221);
nor U11320 (N_11320,N_6017,N_9179);
or U11321 (N_11321,N_8958,N_6243);
nor U11322 (N_11322,N_7355,N_9165);
or U11323 (N_11323,N_5530,N_7371);
or U11324 (N_11324,N_5917,N_6623);
nor U11325 (N_11325,N_5685,N_7754);
nor U11326 (N_11326,N_6288,N_5023);
nor U11327 (N_11327,N_6891,N_6343);
and U11328 (N_11328,N_8403,N_5562);
nand U11329 (N_11329,N_7835,N_7821);
nand U11330 (N_11330,N_6137,N_9632);
nand U11331 (N_11331,N_8829,N_5366);
nand U11332 (N_11332,N_8009,N_9884);
nor U11333 (N_11333,N_5795,N_6778);
or U11334 (N_11334,N_8337,N_7078);
nand U11335 (N_11335,N_7114,N_9307);
or U11336 (N_11336,N_5920,N_5486);
nand U11337 (N_11337,N_6041,N_8474);
nor U11338 (N_11338,N_6885,N_9377);
nor U11339 (N_11339,N_6886,N_5518);
nand U11340 (N_11340,N_5782,N_7093);
nor U11341 (N_11341,N_9135,N_6549);
and U11342 (N_11342,N_6767,N_9797);
and U11343 (N_11343,N_5495,N_7027);
nor U11344 (N_11344,N_5544,N_8193);
nor U11345 (N_11345,N_8290,N_6781);
nand U11346 (N_11346,N_6203,N_6632);
or U11347 (N_11347,N_9464,N_5437);
xnor U11348 (N_11348,N_7151,N_6091);
or U11349 (N_11349,N_5316,N_9016);
nand U11350 (N_11350,N_7328,N_7274);
and U11351 (N_11351,N_9893,N_8001);
nand U11352 (N_11352,N_7008,N_9558);
nand U11353 (N_11353,N_9062,N_8811);
nand U11354 (N_11354,N_8706,N_9556);
and U11355 (N_11355,N_8103,N_9557);
or U11356 (N_11356,N_6705,N_9195);
nor U11357 (N_11357,N_9952,N_6553);
or U11358 (N_11358,N_6149,N_6570);
nand U11359 (N_11359,N_9469,N_5721);
and U11360 (N_11360,N_6918,N_8690);
nor U11361 (N_11361,N_7609,N_6099);
nand U11362 (N_11362,N_9787,N_5317);
nor U11363 (N_11363,N_8220,N_7795);
nor U11364 (N_11364,N_8468,N_9231);
nand U11365 (N_11365,N_7117,N_7919);
and U11366 (N_11366,N_5444,N_5610);
nor U11367 (N_11367,N_9846,N_5416);
nand U11368 (N_11368,N_9290,N_5493);
and U11369 (N_11369,N_5741,N_6761);
and U11370 (N_11370,N_6011,N_9147);
or U11371 (N_11371,N_8717,N_7784);
or U11372 (N_11372,N_9474,N_5735);
nor U11373 (N_11373,N_6976,N_8335);
nor U11374 (N_11374,N_7947,N_9902);
and U11375 (N_11375,N_5007,N_5343);
nor U11376 (N_11376,N_9990,N_8800);
nor U11377 (N_11377,N_9428,N_8941);
or U11378 (N_11378,N_9973,N_6991);
or U11379 (N_11379,N_7799,N_8154);
or U11380 (N_11380,N_5926,N_7247);
or U11381 (N_11381,N_8859,N_9982);
and U11382 (N_11382,N_9319,N_6602);
nor U11383 (N_11383,N_6063,N_6994);
nand U11384 (N_11384,N_6408,N_5223);
and U11385 (N_11385,N_7116,N_6713);
or U11386 (N_11386,N_7246,N_5039);
nand U11387 (N_11387,N_6903,N_8397);
nand U11388 (N_11388,N_6441,N_6336);
or U11389 (N_11389,N_8141,N_7251);
nand U11390 (N_11390,N_5878,N_7163);
or U11391 (N_11391,N_6977,N_8551);
or U11392 (N_11392,N_6218,N_7152);
or U11393 (N_11393,N_6034,N_7199);
and U11394 (N_11394,N_5171,N_9847);
or U11395 (N_11395,N_6580,N_7758);
nor U11396 (N_11396,N_7057,N_8562);
nor U11397 (N_11397,N_8854,N_6613);
nor U11398 (N_11398,N_7210,N_8303);
and U11399 (N_11399,N_5670,N_9620);
nand U11400 (N_11400,N_6259,N_7740);
nor U11401 (N_11401,N_6934,N_6389);
or U11402 (N_11402,N_6782,N_7583);
or U11403 (N_11403,N_6391,N_7272);
nor U11404 (N_11404,N_9056,N_8534);
nand U11405 (N_11405,N_6070,N_9597);
or U11406 (N_11406,N_5417,N_7822);
and U11407 (N_11407,N_8956,N_6848);
and U11408 (N_11408,N_7736,N_6187);
nor U11409 (N_11409,N_8012,N_6747);
or U11410 (N_11410,N_6659,N_8565);
or U11411 (N_11411,N_6870,N_6062);
nor U11412 (N_11412,N_7095,N_7307);
or U11413 (N_11413,N_8186,N_9017);
nand U11414 (N_11414,N_6143,N_8572);
xor U11415 (N_11415,N_8546,N_9836);
and U11416 (N_11416,N_9059,N_5027);
and U11417 (N_11417,N_8724,N_7484);
nor U11418 (N_11418,N_7022,N_9354);
or U11419 (N_11419,N_9890,N_5199);
and U11420 (N_11420,N_6405,N_9458);
or U11421 (N_11421,N_9848,N_6375);
or U11422 (N_11422,N_5175,N_6558);
or U11423 (N_11423,N_8884,N_7894);
xnor U11424 (N_11424,N_6094,N_8346);
nand U11425 (N_11425,N_5031,N_6122);
nand U11426 (N_11426,N_7614,N_9844);
nor U11427 (N_11427,N_9349,N_9775);
nand U11428 (N_11428,N_5600,N_7518);
nand U11429 (N_11429,N_9471,N_6634);
or U11430 (N_11430,N_7320,N_9705);
nor U11431 (N_11431,N_6523,N_7398);
or U11432 (N_11432,N_8515,N_5543);
and U11433 (N_11433,N_6360,N_7503);
or U11434 (N_11434,N_7069,N_7777);
and U11435 (N_11435,N_8255,N_6076);
and U11436 (N_11436,N_7050,N_7345);
nor U11437 (N_11437,N_7168,N_9767);
nand U11438 (N_11438,N_7076,N_7775);
nor U11439 (N_11439,N_5561,N_6527);
or U11440 (N_11440,N_7994,N_5150);
and U11441 (N_11441,N_8807,N_6282);
nor U11442 (N_11442,N_5504,N_7305);
or U11443 (N_11443,N_5550,N_6751);
nand U11444 (N_11444,N_7729,N_5200);
nor U11445 (N_11445,N_7884,N_9073);
nand U11446 (N_11446,N_8790,N_7465);
nand U11447 (N_11447,N_9235,N_5006);
or U11448 (N_11448,N_5485,N_8063);
nand U11449 (N_11449,N_8949,N_9909);
or U11450 (N_11450,N_5903,N_6689);
xor U11451 (N_11451,N_6398,N_9145);
nand U11452 (N_11452,N_6126,N_7587);
nor U11453 (N_11453,N_5378,N_9143);
nor U11454 (N_11454,N_7961,N_8826);
xnor U11455 (N_11455,N_5301,N_6371);
nor U11456 (N_11456,N_7295,N_9527);
or U11457 (N_11457,N_5677,N_8531);
nand U11458 (N_11458,N_9709,N_6914);
nand U11459 (N_11459,N_5767,N_8329);
or U11460 (N_11460,N_7296,N_8327);
or U11461 (N_11461,N_7774,N_5445);
nand U11462 (N_11462,N_7845,N_9294);
and U11463 (N_11463,N_8270,N_6508);
nor U11464 (N_11464,N_8640,N_5737);
nand U11465 (N_11465,N_7198,N_6445);
nand U11466 (N_11466,N_8234,N_9968);
or U11467 (N_11467,N_5135,N_9281);
nor U11468 (N_11468,N_6765,N_6245);
and U11469 (N_11469,N_6811,N_5115);
nor U11470 (N_11470,N_8838,N_8221);
or U11471 (N_11471,N_8373,N_9886);
or U11472 (N_11472,N_7227,N_5146);
and U11473 (N_11473,N_9260,N_7253);
and U11474 (N_11474,N_9585,N_7557);
or U11475 (N_11475,N_7193,N_7779);
nor U11476 (N_11476,N_7316,N_9573);
nand U11477 (N_11477,N_5201,N_5680);
nand U11478 (N_11478,N_9878,N_9138);
nand U11479 (N_11479,N_9634,N_5573);
and U11480 (N_11480,N_9717,N_6563);
and U11481 (N_11481,N_8632,N_7648);
and U11482 (N_11482,N_5749,N_5413);
nor U11483 (N_11483,N_8969,N_6054);
or U11484 (N_11484,N_6393,N_8846);
and U11485 (N_11485,N_6894,N_8487);
and U11486 (N_11486,N_5665,N_5472);
and U11487 (N_11487,N_5242,N_6232);
and U11488 (N_11488,N_5346,N_7695);
or U11489 (N_11489,N_5264,N_8372);
or U11490 (N_11490,N_7750,N_7317);
nand U11491 (N_11491,N_6047,N_9046);
or U11492 (N_11492,N_8466,N_7154);
and U11493 (N_11493,N_5423,N_6350);
nand U11494 (N_11494,N_7283,N_8000);
nand U11495 (N_11495,N_5646,N_6759);
nor U11496 (N_11496,N_7597,N_7055);
nor U11497 (N_11497,N_9690,N_7716);
or U11498 (N_11498,N_6554,N_8511);
nand U11499 (N_11499,N_9885,N_5871);
and U11500 (N_11500,N_8305,N_8939);
and U11501 (N_11501,N_8583,N_7649);
nand U11502 (N_11502,N_6186,N_7232);
nor U11503 (N_11503,N_5859,N_9870);
or U11504 (N_11504,N_6015,N_5182);
nand U11505 (N_11505,N_5726,N_8324);
and U11506 (N_11506,N_5907,N_6773);
nor U11507 (N_11507,N_8205,N_7171);
or U11508 (N_11508,N_8433,N_7629);
nor U11509 (N_11509,N_5815,N_8649);
or U11510 (N_11510,N_8699,N_7136);
nand U11511 (N_11511,N_5538,N_7524);
or U11512 (N_11512,N_8077,N_9454);
xnor U11513 (N_11513,N_5747,N_7929);
nor U11514 (N_11514,N_6172,N_6532);
and U11515 (N_11515,N_8039,N_6763);
or U11516 (N_11516,N_6001,N_8492);
nand U11517 (N_11517,N_8851,N_9714);
and U11518 (N_11518,N_8866,N_7424);
or U11519 (N_11519,N_9807,N_8126);
and U11520 (N_11520,N_8425,N_6421);
nand U11521 (N_11521,N_6913,N_6394);
nand U11522 (N_11522,N_9409,N_7292);
nor U11523 (N_11523,N_8982,N_6268);
nand U11524 (N_11524,N_5436,N_8362);
nor U11525 (N_11525,N_8954,N_9854);
or U11526 (N_11526,N_6274,N_8459);
nor U11527 (N_11527,N_9553,N_6196);
nand U11528 (N_11528,N_6808,N_6770);
and U11529 (N_11529,N_6027,N_8902);
nand U11530 (N_11530,N_8041,N_9925);
and U11531 (N_11531,N_8512,N_8020);
and U11532 (N_11532,N_9563,N_8272);
or U11533 (N_11533,N_7321,N_7237);
or U11534 (N_11534,N_7905,N_9366);
or U11535 (N_11535,N_8092,N_7705);
nor U11536 (N_11536,N_8281,N_8117);
or U11537 (N_11537,N_8036,N_5827);
or U11538 (N_11538,N_5837,N_6796);
nand U11539 (N_11539,N_5347,N_6485);
nand U11540 (N_11540,N_6863,N_7517);
nor U11541 (N_11541,N_9944,N_6116);
nor U11542 (N_11542,N_6192,N_8694);
and U11543 (N_11543,N_5342,N_6125);
or U11544 (N_11544,N_9796,N_6373);
and U11545 (N_11545,N_5319,N_8291);
nand U11546 (N_11546,N_6875,N_9116);
and U11547 (N_11547,N_5356,N_9770);
and U11548 (N_11548,N_5849,N_9889);
nor U11549 (N_11549,N_5193,N_6425);
and U11550 (N_11550,N_9136,N_7979);
nor U11551 (N_11551,N_7091,N_6385);
or U11552 (N_11552,N_8778,N_9425);
and U11553 (N_11553,N_8931,N_9329);
and U11554 (N_11554,N_7783,N_8233);
nor U11555 (N_11555,N_6815,N_6049);
or U11556 (N_11556,N_9274,N_8169);
or U11557 (N_11557,N_6270,N_5572);
or U11558 (N_11558,N_8214,N_8779);
or U11559 (N_11559,N_8614,N_5954);
nor U11560 (N_11560,N_5204,N_5482);
nor U11561 (N_11561,N_8190,N_8420);
nand U11562 (N_11562,N_8731,N_5912);
and U11563 (N_11563,N_8203,N_9105);
nor U11564 (N_11564,N_8161,N_6316);
and U11565 (N_11565,N_9000,N_6739);
nor U11566 (N_11566,N_6455,N_5929);
and U11567 (N_11567,N_6970,N_8348);
nor U11568 (N_11568,N_5987,N_9196);
and U11569 (N_11569,N_9680,N_7720);
nor U11570 (N_11570,N_5800,N_8742);
or U11571 (N_11571,N_7602,N_7220);
nor U11572 (N_11572,N_9077,N_7430);
nand U11573 (N_11573,N_5761,N_5345);
nor U11574 (N_11574,N_9453,N_8456);
and U11575 (N_11575,N_8909,N_8390);
and U11576 (N_11576,N_5352,N_8047);
nand U11577 (N_11577,N_7628,N_6636);
nand U11578 (N_11578,N_5879,N_6978);
and U11579 (N_11579,N_9452,N_6801);
nor U11580 (N_11580,N_7759,N_7833);
and U11581 (N_11581,N_9263,N_9209);
nor U11582 (N_11582,N_6664,N_9975);
nand U11583 (N_11583,N_9276,N_8500);
and U11584 (N_11584,N_5579,N_6292);
nor U11585 (N_11585,N_9758,N_6896);
xor U11586 (N_11586,N_5469,N_5823);
or U11587 (N_11587,N_5944,N_5576);
and U11588 (N_11588,N_7428,N_9638);
and U11589 (N_11589,N_7063,N_8045);
or U11590 (N_11590,N_6493,N_7886);
or U11591 (N_11591,N_6309,N_6572);
or U11592 (N_11592,N_6364,N_6927);
nand U11593 (N_11593,N_5376,N_5911);
or U11594 (N_11594,N_5804,N_6272);
nand U11595 (N_11595,N_8168,N_7311);
and U11596 (N_11596,N_7365,N_8627);
or U11597 (N_11597,N_7123,N_9989);
xnor U11598 (N_11598,N_8617,N_9321);
nand U11599 (N_11599,N_6310,N_8830);
or U11600 (N_11600,N_6429,N_5091);
and U11601 (N_11601,N_5575,N_8645);
nand U11602 (N_11602,N_9765,N_5990);
and U11603 (N_11603,N_7980,N_5961);
and U11604 (N_11604,N_8140,N_8087);
and U11605 (N_11605,N_7412,N_5137);
and U11606 (N_11606,N_7024,N_7046);
nand U11607 (N_11607,N_6502,N_8834);
or U11608 (N_11608,N_7551,N_5602);
or U11609 (N_11609,N_6439,N_9987);
or U11610 (N_11610,N_9047,N_8679);
nand U11611 (N_11611,N_8792,N_6521);
or U11612 (N_11612,N_9015,N_9669);
and U11613 (N_11613,N_9312,N_5777);
or U11614 (N_11614,N_5197,N_7967);
nand U11615 (N_11615,N_9920,N_6525);
nand U11616 (N_11616,N_9922,N_5032);
nand U11617 (N_11617,N_6134,N_9693);
and U11618 (N_11618,N_9814,N_5461);
nor U11619 (N_11619,N_7387,N_5046);
and U11620 (N_11620,N_5454,N_9412);
nand U11621 (N_11621,N_5465,N_8751);
or U11622 (N_11622,N_5686,N_9867);
and U11623 (N_11623,N_5758,N_8351);
nand U11624 (N_11624,N_7229,N_7444);
or U11625 (N_11625,N_7949,N_7324);
nor U11626 (N_11626,N_8762,N_7099);
and U11627 (N_11627,N_8476,N_7452);
nand U11628 (N_11628,N_7018,N_5768);
and U11629 (N_11629,N_5457,N_5118);
or U11630 (N_11630,N_6157,N_8889);
or U11631 (N_11631,N_8216,N_8019);
or U11632 (N_11632,N_6478,N_6704);
and U11633 (N_11633,N_9173,N_6177);
and U11634 (N_11634,N_5134,N_5354);
or U11635 (N_11635,N_9945,N_8198);
and U11636 (N_11636,N_6229,N_5188);
nand U11637 (N_11637,N_5382,N_7189);
nand U11638 (N_11638,N_6920,N_6516);
nor U11639 (N_11639,N_5642,N_9285);
nand U11640 (N_11640,N_7768,N_8384);
and U11641 (N_11641,N_7708,N_5314);
nand U11642 (N_11642,N_5731,N_8957);
and U11643 (N_11643,N_9449,N_6660);
and U11644 (N_11644,N_9410,N_8714);
and U11645 (N_11645,N_9640,N_7741);
and U11646 (N_11646,N_5507,N_7049);
nand U11647 (N_11647,N_9267,N_6980);
nand U11648 (N_11648,N_9205,N_9368);
nor U11649 (N_11649,N_9759,N_8323);
nand U11650 (N_11650,N_8932,N_9533);
nor U11651 (N_11651,N_9175,N_7470);
or U11652 (N_11652,N_8318,N_7238);
and U11653 (N_11653,N_8610,N_8874);
and U11654 (N_11654,N_6387,N_7221);
nor U11655 (N_11655,N_6653,N_5373);
and U11656 (N_11656,N_7429,N_6798);
and U11657 (N_11657,N_9310,N_9965);
nor U11658 (N_11658,N_8386,N_9011);
nor U11659 (N_11659,N_7485,N_6484);
nor U11660 (N_11660,N_8013,N_8680);
and U11661 (N_11661,N_6135,N_6486);
nand U11662 (N_11662,N_5370,N_7700);
nand U11663 (N_11663,N_5509,N_6858);
nand U11664 (N_11664,N_9639,N_5781);
nor U11665 (N_11665,N_7837,N_5271);
or U11666 (N_11666,N_7930,N_5725);
nand U11667 (N_11667,N_9559,N_8998);
and U11668 (N_11668,N_8398,N_8865);
and U11669 (N_11669,N_6743,N_5994);
nand U11670 (N_11670,N_9156,N_8274);
and U11671 (N_11671,N_9025,N_8299);
nor U11672 (N_11672,N_7900,N_7693);
nor U11673 (N_11673,N_8280,N_9752);
nor U11674 (N_11674,N_5112,N_6861);
nor U11675 (N_11675,N_7957,N_8798);
and U11676 (N_11676,N_9513,N_6766);
and U11677 (N_11677,N_6881,N_5658);
or U11678 (N_11678,N_9674,N_5152);
or U11679 (N_11679,N_5435,N_9278);
nor U11680 (N_11680,N_9561,N_8989);
nor U11681 (N_11681,N_6730,N_7421);
nand U11682 (N_11682,N_8669,N_5002);
or U11683 (N_11683,N_7904,N_9074);
and U11684 (N_11684,N_8502,N_7051);
or U11685 (N_11685,N_6156,N_8194);
and U11686 (N_11686,N_9021,N_7081);
nand U11687 (N_11687,N_8157,N_9429);
nor U11688 (N_11688,N_7639,N_6402);
nand U11689 (N_11689,N_8936,N_6853);
nor U11690 (N_11690,N_5299,N_9786);
nand U11691 (N_11691,N_9876,N_5158);
or U11692 (N_11692,N_5826,N_9995);
or U11693 (N_11693,N_5545,N_8585);
and U11694 (N_11694,N_9299,N_5066);
and U11695 (N_11695,N_5867,N_9604);
or U11696 (N_11696,N_8908,N_8125);
nor U11697 (N_11697,N_7176,N_6422);
and U11698 (N_11698,N_8548,N_7284);
xnor U11699 (N_11699,N_9348,N_5529);
nand U11700 (N_11700,N_6942,N_5169);
nand U11701 (N_11701,N_6359,N_7214);
xnor U11702 (N_11702,N_8569,N_7600);
nand U11703 (N_11703,N_8240,N_9868);
and U11704 (N_11704,N_5121,N_6255);
nand U11705 (N_11705,N_6118,N_7478);
or U11706 (N_11706,N_9733,N_5221);
nand U11707 (N_11707,N_9110,N_6898);
or U11708 (N_11708,N_5126,N_5083);
nand U11709 (N_11709,N_9065,N_5692);
nand U11710 (N_11710,N_7910,N_7131);
and U11711 (N_11711,N_9122,N_7195);
nand U11712 (N_11712,N_7344,N_7673);
nor U11713 (N_11713,N_5938,N_9352);
or U11714 (N_11714,N_9741,N_5410);
and U11715 (N_11715,N_8697,N_6974);
nand U11716 (N_11716,N_5783,N_8993);
nand U11717 (N_11717,N_8007,N_8006);
or U11718 (N_11718,N_9297,N_8953);
nand U11719 (N_11719,N_7203,N_5074);
nor U11720 (N_11720,N_6703,N_9180);
or U11721 (N_11721,N_6722,N_7108);
or U11722 (N_11722,N_9061,N_6283);
and U11723 (N_11723,N_6655,N_9103);
xor U11724 (N_11724,N_5693,N_7166);
and U11725 (N_11725,N_9773,N_8444);
or U11726 (N_11726,N_6588,N_7102);
or U11727 (N_11727,N_5861,N_5133);
or U11728 (N_11728,N_5215,N_5272);
and U11729 (N_11729,N_9419,N_6642);
nand U11730 (N_11730,N_7921,N_8442);
nand U11731 (N_11731,N_7282,N_5329);
nor U11732 (N_11732,N_8239,N_5263);
nor U11733 (N_11733,N_9102,N_9184);
and U11734 (N_11734,N_9967,N_9013);
or U11735 (N_11735,N_5008,N_9851);
nor U11736 (N_11736,N_8952,N_9551);
nand U11737 (N_11737,N_5628,N_9832);
or U11738 (N_11738,N_6424,N_8286);
and U11739 (N_11739,N_9456,N_6189);
nor U11740 (N_11740,N_9230,N_8431);
nor U11741 (N_11741,N_6652,N_7275);
nand U11742 (N_11742,N_9335,N_6555);
nor U11743 (N_11743,N_9038,N_7397);
nand U11744 (N_11744,N_9715,N_8709);
and U11745 (N_11745,N_7850,N_6998);
nand U11746 (N_11746,N_7983,N_6938);
nor U11747 (N_11747,N_8405,N_9568);
nor U11748 (N_11748,N_6097,N_8098);
or U11749 (N_11749,N_9060,N_7657);
and U11750 (N_11750,N_8899,N_7635);
nor U11751 (N_11751,N_7289,N_7726);
nor U11752 (N_11752,N_6103,N_8066);
and U11753 (N_11753,N_6435,N_7362);
nand U11754 (N_11754,N_8760,N_5009);
nor U11755 (N_11755,N_6921,N_5368);
or U11756 (N_11756,N_8628,N_5443);
and U11757 (N_11757,N_8217,N_8230);
or U11758 (N_11758,N_9605,N_5000);
nor U11759 (N_11759,N_9519,N_6830);
or U11760 (N_11760,N_6737,N_8325);
xnor U11761 (N_11761,N_9140,N_5825);
nor U11762 (N_11762,N_5153,N_7105);
nand U11763 (N_11763,N_9125,N_5265);
nand U11764 (N_11764,N_7178,N_7743);
nand U11765 (N_11765,N_7157,N_8452);
nand U11766 (N_11766,N_5798,N_7194);
nand U11767 (N_11767,N_9959,N_6417);
and U11768 (N_11768,N_5110,N_6117);
and U11769 (N_11769,N_5124,N_8127);
nand U11770 (N_11770,N_5104,N_9763);
or U11771 (N_11771,N_8297,N_7668);
and U11772 (N_11772,N_9603,N_5894);
and U11773 (N_11773,N_5145,N_5902);
and U11774 (N_11774,N_8659,N_8723);
and U11775 (N_11775,N_9104,N_6327);
or U11776 (N_11776,N_7437,N_9128);
nor U11777 (N_11777,N_9939,N_8406);
and U11778 (N_11778,N_7508,N_5706);
nand U11779 (N_11779,N_7926,N_7643);
and U11780 (N_11780,N_9337,N_7870);
or U11781 (N_11781,N_9555,N_5885);
nand U11782 (N_11782,N_7128,N_9227);
nand U11783 (N_11783,N_8619,N_9259);
nor U11784 (N_11784,N_9655,N_8200);
and U11785 (N_11785,N_5683,N_7542);
and U11786 (N_11786,N_7267,N_6695);
and U11787 (N_11787,N_9843,N_6836);
and U11788 (N_11788,N_9188,N_8685);
nand U11789 (N_11789,N_7086,N_6785);
nor U11790 (N_11790,N_7934,N_6944);
or U11791 (N_11791,N_8227,N_6372);
or U11792 (N_11792,N_8857,N_5539);
and U11793 (N_11793,N_7115,N_6388);
nor U11794 (N_11794,N_7492,N_9809);
or U11795 (N_11795,N_5297,N_9595);
nand U11796 (N_11796,N_9517,N_9411);
and U11797 (N_11797,N_7575,N_7971);
nand U11798 (N_11798,N_7683,N_8584);
nor U11799 (N_11799,N_8944,N_5930);
nor U11800 (N_11800,N_7434,N_9744);
or U11801 (N_11801,N_6534,N_9433);
nor U11802 (N_11802,N_6744,N_8396);
and U11803 (N_11803,N_5429,N_5218);
and U11804 (N_11804,N_9007,N_9247);
nand U11805 (N_11805,N_8491,N_6547);
or U11806 (N_11806,N_7595,N_8560);
nand U11807 (N_11807,N_8078,N_6909);
and U11808 (N_11808,N_8068,N_5291);
and U11809 (N_11809,N_7449,N_9641);
or U11810 (N_11810,N_6838,N_9480);
nor U11811 (N_11811,N_6294,N_7922);
nor U11812 (N_11812,N_9042,N_7281);
nor U11813 (N_11813,N_7224,N_7625);
or U11814 (N_11814,N_8247,N_9607);
and U11815 (N_11815,N_9501,N_8284);
or U11816 (N_11816,N_6719,N_7908);
or U11817 (N_11817,N_8374,N_9496);
or U11818 (N_11818,N_7230,N_7453);
and U11819 (N_11819,N_9936,N_6712);
or U11820 (N_11820,N_8070,N_8093);
and U11821 (N_11821,N_7348,N_9126);
or U11822 (N_11822,N_5748,N_7627);
and U11823 (N_11823,N_8542,N_5237);
nor U11824 (N_11824,N_5236,N_5279);
nor U11825 (N_11825,N_9445,N_5700);
nor U11826 (N_11826,N_9754,N_8517);
and U11827 (N_11827,N_8848,N_8597);
and U11828 (N_11828,N_9826,N_5090);
and U11829 (N_11829,N_5058,N_8121);
nor U11830 (N_11830,N_5129,N_6102);
nand U11831 (N_11831,N_7909,N_5010);
nand U11832 (N_11832,N_7219,N_6338);
or U11833 (N_11833,N_5688,N_7666);
nor U11834 (N_11834,N_7034,N_7294);
nor U11835 (N_11835,N_9048,N_6772);
nor U11836 (N_11836,N_5848,N_6501);
nand U11837 (N_11837,N_5001,N_6676);
nor U11838 (N_11838,N_9681,N_9149);
or U11839 (N_11839,N_5313,N_6048);
xnor U11840 (N_11840,N_8005,N_7803);
and U11841 (N_11841,N_8321,N_5367);
nor U11842 (N_11842,N_9793,N_6030);
nand U11843 (N_11843,N_8767,N_9552);
nor U11844 (N_11844,N_7728,N_9132);
xnor U11845 (N_11845,N_5760,N_6353);
or U11846 (N_11846,N_7487,N_7829);
and U11847 (N_11847,N_8819,N_7381);
and U11848 (N_11848,N_5789,N_8471);
nor U11849 (N_11849,N_6337,N_6275);
and U11850 (N_11850,N_5643,N_6453);
nand U11851 (N_11851,N_7677,N_8733);
nand U11852 (N_11852,N_8074,N_6598);
and U11853 (N_11853,N_9171,N_9051);
nand U11854 (N_11854,N_7678,N_8391);
or U11855 (N_11855,N_7605,N_6908);
and U11856 (N_11856,N_9216,N_7601);
nor U11857 (N_11857,N_6053,N_6438);
nand U11858 (N_11858,N_8457,N_8283);
nor U11859 (N_11859,N_5792,N_9441);
nor U11860 (N_11860,N_6639,N_5026);
and U11861 (N_11861,N_7448,N_5500);
nor U11862 (N_11862,N_6615,N_6257);
and U11863 (N_11863,N_8588,N_7550);
and U11864 (N_11864,N_6346,N_9574);
xnor U11865 (N_11865,N_8594,N_7040);
xor U11866 (N_11866,N_6499,N_7303);
and U11867 (N_11867,N_6859,N_7319);
and U11868 (N_11868,N_7002,N_9663);
or U11869 (N_11869,N_5440,N_9224);
nand U11870 (N_11870,N_9949,N_6609);
xor U11871 (N_11871,N_5270,N_9652);
and U11872 (N_11872,N_6771,N_7206);
nor U11873 (N_11873,N_8879,N_9119);
nor U11874 (N_11874,N_6672,N_8959);
nor U11875 (N_11875,N_9845,N_8803);
or U11876 (N_11876,N_8144,N_6857);
or U11877 (N_11877,N_8530,N_8079);
xor U11878 (N_11878,N_6803,N_5999);
and U11879 (N_11879,N_7200,N_8364);
nand U11880 (N_11880,N_5385,N_5148);
nor U11881 (N_11881,N_5028,N_6390);
or U11882 (N_11882,N_8836,N_6311);
or U11883 (N_11883,N_6109,N_6314);
and U11884 (N_11884,N_6124,N_9355);
nor U11885 (N_11885,N_7612,N_6223);
or U11886 (N_11886,N_6961,N_6188);
nor U11887 (N_11887,N_9234,N_6104);
nand U11888 (N_11888,N_8032,N_5238);
and U11889 (N_11889,N_7747,N_7242);
nor U11890 (N_11890,N_6943,N_8377);
nand U11891 (N_11891,N_5746,N_8008);
nor U11892 (N_11892,N_5434,N_7634);
nor U11893 (N_11893,N_8701,N_7358);
and U11894 (N_11894,N_8557,N_7901);
nor U11895 (N_11895,N_7766,N_8134);
or U11896 (N_11896,N_5183,N_5364);
or U11897 (N_11897,N_5622,N_6882);
or U11898 (N_11898,N_9448,N_8556);
nor U11899 (N_11899,N_7782,N_7388);
nor U11900 (N_11900,N_9694,N_8004);
or U11901 (N_11901,N_8660,N_9430);
or U11902 (N_11902,N_5381,N_8503);
nor U11903 (N_11903,N_6237,N_6611);
or U11904 (N_11904,N_8780,N_6684);
nor U11905 (N_11905,N_8060,N_6802);
nand U11906 (N_11906,N_7770,N_6752);
nand U11907 (N_11907,N_9579,N_5514);
nand U11908 (N_11908,N_6088,N_9648);
or U11909 (N_11909,N_5647,N_6174);
and U11910 (N_11910,N_8549,N_7346);
nor U11911 (N_11911,N_5854,N_5887);
or U11912 (N_11912,N_8981,N_9913);
or U11913 (N_11913,N_9279,N_6899);
nand U11914 (N_11914,N_5391,N_6951);
nand U11915 (N_11915,N_5654,N_5018);
or U11916 (N_11916,N_9882,N_7888);
nor U11917 (N_11917,N_8172,N_5422);
nand U11918 (N_11918,N_7327,N_7590);
nand U11919 (N_11919,N_6236,N_7969);
nor U11920 (N_11920,N_8018,N_6069);
nand U11921 (N_11921,N_5079,N_9028);
and U11922 (N_11922,N_5649,N_7623);
nor U11923 (N_11923,N_7119,N_8975);
nor U11924 (N_11924,N_8842,N_8276);
nand U11925 (N_11925,N_5895,N_6840);
or U11926 (N_11926,N_9477,N_8828);
nor U11927 (N_11927,N_7731,N_5567);
or U11928 (N_11928,N_5528,N_6691);
nor U11929 (N_11929,N_8809,N_6456);
nor U11930 (N_11930,N_8173,N_6287);
or U11931 (N_11931,N_8900,N_7730);
or U11932 (N_11932,N_6917,N_6591);
nand U11933 (N_11933,N_8861,N_9250);
nor U11934 (N_11934,N_8590,N_5205);
or U11935 (N_11935,N_5111,N_6792);
nor U11936 (N_11936,N_9014,N_5811);
nor U11937 (N_11937,N_7607,N_6637);
and U11938 (N_11938,N_7935,N_6912);
or U11939 (N_11939,N_9473,N_6416);
nand U11940 (N_11940,N_5730,N_8711);
nand U11941 (N_11941,N_9921,N_6150);
and U11942 (N_11942,N_5574,N_7718);
or U11943 (N_11943,N_8053,N_6657);
nand U11944 (N_11944,N_9861,N_6700);
nor U11945 (N_11945,N_8043,N_9300);
nand U11946 (N_11946,N_9725,N_8755);
nor U11947 (N_11947,N_5086,N_5106);
nand U11948 (N_11948,N_9592,N_6833);
nor U11949 (N_11949,N_5406,N_7342);
nand U11950 (N_11950,N_9416,N_5548);
or U11951 (N_11951,N_7129,N_7574);
nor U11952 (N_11952,N_8728,N_7723);
and U11953 (N_11953,N_6825,N_5361);
nand U11954 (N_11954,N_8824,N_7082);
or U11955 (N_11955,N_9804,N_9327);
and U11956 (N_11956,N_9783,N_5853);
and U11957 (N_11957,N_5309,N_9980);
and U11958 (N_11958,N_6031,N_5947);
or U11959 (N_11959,N_7882,N_5269);
nor U11960 (N_11960,N_9386,N_9120);
nor U11961 (N_11961,N_7584,N_6140);
or U11962 (N_11962,N_8559,N_7304);
nor U11963 (N_11963,N_6050,N_9331);
and U11964 (N_11964,N_8129,N_6856);
and U11965 (N_11965,N_9948,N_5208);
or U11966 (N_11966,N_9781,N_9034);
and U11967 (N_11967,N_6617,N_8887);
and U11968 (N_11968,N_9670,N_9296);
nand U11969 (N_11969,N_5335,N_7017);
or U11970 (N_11970,N_5202,N_7626);
nor U11971 (N_11971,N_5077,N_9742);
or U11972 (N_11972,N_7653,N_8528);
nor U11973 (N_11973,N_8882,N_6610);
nand U11974 (N_11974,N_9525,N_7515);
or U11975 (N_11975,N_6119,N_8875);
nand U11976 (N_11976,N_6536,N_8483);
and U11977 (N_11977,N_8055,N_6901);
or U11978 (N_11978,N_7100,N_8293);
and U11979 (N_11979,N_8791,N_6879);
nor U11980 (N_11980,N_9857,N_6769);
nor U11981 (N_11981,N_9869,N_7028);
and U11982 (N_11982,N_6586,N_9206);
nand U11983 (N_11983,N_9753,N_6973);
nand U11984 (N_11984,N_9148,N_9498);
and U11985 (N_11985,N_7528,N_8984);
or U11986 (N_11986,N_6867,N_9817);
nor U11987 (N_11987,N_9768,N_9200);
nor U11988 (N_11988,N_6147,N_8745);
or U11989 (N_11989,N_5526,N_7656);
and U11990 (N_11990,N_5122,N_7907);
nor U11991 (N_11991,N_6169,N_7359);
or U11992 (N_11992,N_5966,N_9100);
nor U11993 (N_11993,N_6384,N_8073);
and U11994 (N_11994,N_6376,N_7896);
nand U11995 (N_11995,N_9650,N_9727);
or U11996 (N_11996,N_6262,N_6736);
or U11997 (N_11997,N_8876,N_8052);
and U11998 (N_11998,N_8759,N_9087);
nor U11999 (N_11999,N_7933,N_8606);
and U12000 (N_12000,N_5427,N_7906);
nor U12001 (N_12001,N_5918,N_8935);
nand U12002 (N_12002,N_7165,N_5060);
nand U12003 (N_12003,N_8207,N_6566);
or U12004 (N_12004,N_5824,N_9369);
or U12005 (N_12005,N_8353,N_7856);
nand U12006 (N_12006,N_7012,N_8225);
nor U12007 (N_12007,N_9127,N_9099);
and U12008 (N_12008,N_9083,N_7939);
or U12009 (N_12009,N_6479,N_8592);
or U12010 (N_12010,N_9291,N_9382);
nor U12011 (N_12011,N_7536,N_7571);
nor U12012 (N_12012,N_7389,N_7815);
nor U12013 (N_12013,N_9721,N_7432);
nor U12014 (N_12014,N_9244,N_5802);
or U12015 (N_12015,N_7631,N_5015);
nor U12016 (N_12016,N_5362,N_7080);
nor U12017 (N_12017,N_9676,N_5310);
and U12018 (N_12018,N_5460,N_7698);
nor U12019 (N_12019,N_9986,N_6524);
nor U12020 (N_12020,N_7925,N_6071);
nor U12021 (N_12021,N_7382,N_7290);
or U12022 (N_12022,N_6890,N_9699);
nor U12023 (N_12023,N_9010,N_8246);
or U12024 (N_12024,N_7330,N_7416);
and U12025 (N_12025,N_6560,N_7868);
nor U12026 (N_12026,N_7139,N_5293);
nand U12027 (N_12027,N_9356,N_5184);
nand U12028 (N_12028,N_6374,N_8684);
and U12029 (N_12029,N_8903,N_6805);
or U12030 (N_12030,N_5734,N_5927);
and U12031 (N_12031,N_7960,N_6790);
and U12032 (N_12032,N_9799,N_8541);
nand U12033 (N_12033,N_9489,N_7761);
nor U12034 (N_12034,N_8014,N_9086);
nand U12035 (N_12035,N_6115,N_7826);
nand U12036 (N_12036,N_7594,N_6666);
or U12037 (N_12037,N_7615,N_5974);
or U12038 (N_12038,N_7420,N_9503);
or U12039 (N_12039,N_6835,N_7390);
or U12040 (N_12040,N_6862,N_6789);
and U12041 (N_12041,N_8211,N_7415);
and U12042 (N_12042,N_8099,N_5591);
or U12043 (N_12043,N_7404,N_8094);
or U12044 (N_12044,N_7858,N_6158);
or U12045 (N_12045,N_5759,N_7439);
or U12046 (N_12046,N_7924,N_6396);
nand U12047 (N_12047,N_9572,N_5268);
nor U12048 (N_12048,N_5866,N_7865);
nand U12049 (N_12049,N_6599,N_7467);
or U12050 (N_12050,N_9280,N_6321);
and U12051 (N_12051,N_5908,N_6670);
and U12052 (N_12052,N_9825,N_5359);
nand U12053 (N_12053,N_6807,N_5835);
and U12054 (N_12054,N_5414,N_8540);
or U12055 (N_12055,N_7778,N_5014);
and U12056 (N_12056,N_8970,N_6128);
nand U12057 (N_12057,N_6239,N_7490);
nor U12058 (N_12058,N_6869,N_7243);
and U12059 (N_12059,N_7580,N_7501);
nor U12060 (N_12060,N_9746,N_5595);
nor U12061 (N_12061,N_6235,N_7339);
or U12062 (N_12062,N_6928,N_9849);
or U12063 (N_12063,N_6791,N_9904);
and U12064 (N_12064,N_8241,N_9309);
nor U12065 (N_12065,N_7918,N_6982);
and U12066 (N_12066,N_7175,N_6211);
or U12067 (N_12067,N_9078,N_5102);
nor U12068 (N_12068,N_8102,N_6592);
nand U12069 (N_12069,N_7257,N_7757);
nand U12070 (N_12070,N_5534,N_8664);
or U12071 (N_12071,N_6226,N_9554);
nand U12072 (N_12072,N_6923,N_9228);
and U12073 (N_12073,N_9081,N_5980);
nor U12074 (N_12074,N_8042,N_7823);
nand U12075 (N_12075,N_6365,N_5489);
nor U12076 (N_12076,N_7455,N_8718);
nor U12077 (N_12077,N_7286,N_5473);
nor U12078 (N_12078,N_5648,N_8238);
nand U12079 (N_12079,N_5951,N_7749);
or U12080 (N_12080,N_6933,N_7264);
nand U12081 (N_12081,N_5655,N_9991);
and U12082 (N_12082,N_7261,N_7873);
xor U12083 (N_12083,N_6633,N_8162);
and U12084 (N_12084,N_5584,N_7067);
and U12085 (N_12085,N_6092,N_6625);
or U12086 (N_12086,N_5967,N_6900);
nor U12087 (N_12087,N_7486,N_7690);
or U12088 (N_12088,N_9097,N_5332);
nand U12089 (N_12089,N_7064,N_5068);
nor U12090 (N_12090,N_8737,N_6000);
and U12091 (N_12091,N_9190,N_5213);
nand U12092 (N_12092,N_7745,N_8106);
and U12093 (N_12093,N_6884,N_7392);
or U12094 (N_12094,N_5552,N_8600);
nor U12095 (N_12095,N_6382,N_7891);
or U12096 (N_12096,N_9258,N_9246);
nor U12097 (N_12097,N_9547,N_5772);
or U12098 (N_12098,N_6279,N_7031);
and U12099 (N_12099,N_7606,N_5080);
and U12100 (N_12100,N_5030,N_7360);
and U12101 (N_12101,N_7744,N_5085);
or U12102 (N_12102,N_6758,N_8768);
or U12103 (N_12103,N_7384,N_7553);
and U12104 (N_12104,N_6883,N_9361);
nor U12105 (N_12105,N_5078,N_8489);
or U12106 (N_12106,N_8210,N_9614);
nand U12107 (N_12107,N_8816,N_9043);
or U12108 (N_12108,N_6564,N_5071);
or U12109 (N_12109,N_9315,N_6131);
or U12110 (N_12110,N_7721,N_8571);
and U12111 (N_12111,N_9026,N_9785);
and U12112 (N_12112,N_8448,N_8962);
nor U12113 (N_12113,N_6874,N_7211);
nor U12114 (N_12114,N_5047,N_7202);
nand U12115 (N_12115,N_6300,N_6026);
nor U12116 (N_12116,N_9071,N_6827);
and U12117 (N_12117,N_5626,N_8736);
and U12118 (N_12118,N_6675,N_9467);
nand U12119 (N_12119,N_5641,N_7848);
and U12120 (N_12120,N_7089,N_7277);
nor U12121 (N_12121,N_5981,N_5919);
nor U12122 (N_12122,N_5209,N_6368);
nor U12123 (N_12123,N_8794,N_9118);
and U12124 (N_12124,N_8878,N_8150);
nand U12125 (N_12125,N_8801,N_9993);
nand U12126 (N_12126,N_6968,N_7618);
or U12127 (N_12127,N_6699,N_9311);
nor U12128 (N_12128,N_9124,N_9313);
nor U12129 (N_12129,N_8582,N_8916);
or U12130 (N_12130,N_5147,N_5611);
nand U12131 (N_12131,N_9199,N_5598);
or U12132 (N_12132,N_7250,N_5092);
nand U12133 (N_12133,N_7748,N_6304);
and U12134 (N_12134,N_6845,N_7963);
or U12135 (N_12135,N_5389,N_9098);
nor U12136 (N_12136,N_5374,N_9865);
and U12137 (N_12137,N_8269,N_8443);
or U12138 (N_12138,N_7945,N_7174);
nand U12139 (N_12139,N_7098,N_5053);
nand U12140 (N_12140,N_8371,N_8105);
nand U12141 (N_12141,N_7180,N_8334);
xor U12142 (N_12142,N_5821,N_8509);
nor U12143 (N_12143,N_6043,N_9675);
nor U12144 (N_12144,N_5520,N_5225);
nand U12145 (N_12145,N_6496,N_8160);
and U12146 (N_12146,N_9974,N_7694);
nand U12147 (N_12147,N_7946,N_6155);
and U12148 (N_12148,N_9900,N_8620);
and U12149 (N_12149,N_5884,N_8522);
or U12150 (N_12150,N_7186,N_9734);
nand U12151 (N_12151,N_8676,N_5419);
nand U12152 (N_12152,N_5719,N_7675);
nand U12153 (N_12153,N_9001,N_7632);
or U12154 (N_12154,N_7425,N_7493);
nand U12155 (N_12155,N_9178,N_6984);
nor U12156 (N_12156,N_8712,N_8527);
nand U12157 (N_12157,N_7791,N_9421);
nand U12158 (N_12158,N_6410,N_7474);
nor U12159 (N_12159,N_9450,N_6932);
or U12160 (N_12160,N_6022,N_9130);
or U12161 (N_12161,N_7158,N_9151);
nor U12162 (N_12162,N_5254,N_5403);
and U12163 (N_12163,N_9589,N_6227);
nand U12164 (N_12164,N_8279,N_8663);
nand U12165 (N_12165,N_9971,N_6518);
nand U12166 (N_12166,N_7546,N_9109);
nand U12167 (N_12167,N_7857,N_7880);
nor U12168 (N_12168,N_5524,N_8601);
xnor U12169 (N_12169,N_6113,N_6138);
nor U12170 (N_12170,N_5409,N_8796);
nand U12171 (N_12171,N_5844,N_8076);
nor U12172 (N_12172,N_5128,N_6849);
nand U12173 (N_12173,N_5463,N_9615);
and U12174 (N_12174,N_7372,N_5190);
and U12175 (N_12175,N_7457,N_7589);
and U12176 (N_12176,N_9495,N_7879);
and U12177 (N_12177,N_7534,N_7513);
or U12178 (N_12178,N_5638,N_6463);
and U12179 (N_12179,N_6831,N_9163);
and U12180 (N_12180,N_5492,N_5284);
or U12181 (N_12181,N_7075,N_8243);
or U12182 (N_12182,N_5978,N_8462);
and U12183 (N_12183,N_7725,N_8832);
and U12184 (N_12184,N_8133,N_7598);
or U12185 (N_12185,N_9873,N_9566);
and U12186 (N_12186,N_5267,N_7847);
nor U12187 (N_12187,N_9022,N_9685);
and U12188 (N_12188,N_8097,N_8260);
nor U12189 (N_12189,N_5424,N_8675);
nand U12190 (N_12190,N_7399,N_5499);
and U12191 (N_12191,N_6222,N_7502);
nor U12192 (N_12192,N_5220,N_8591);
nor U12193 (N_12193,N_9504,N_6021);
and U12194 (N_12194,N_5605,N_6843);
nor U12195 (N_12195,N_8677,N_5705);
or U12196 (N_12196,N_9168,N_7992);
nor U12197 (N_12197,N_8750,N_6495);
or U12198 (N_12198,N_8333,N_9684);
nor U12199 (N_12199,N_8360,N_7825);
nand U12200 (N_12200,N_7667,N_6779);
and U12201 (N_12201,N_9089,N_8248);
or U12202 (N_12202,N_8365,N_5691);
or U12203 (N_12203,N_5191,N_7004);
xnor U12204 (N_12204,N_6055,N_9068);
or U12205 (N_12205,N_9570,N_5985);
nor U12206 (N_12206,N_9139,N_8188);
nor U12207 (N_12207,N_5957,N_6214);
and U12208 (N_12208,N_8553,N_9972);
nand U12209 (N_12209,N_9378,N_6078);
or U12210 (N_12210,N_6089,N_8629);
nor U12211 (N_12211,N_8943,N_6600);
nor U12212 (N_12212,N_9822,N_7554);
or U12213 (N_12213,N_9644,N_7436);
nand U12214 (N_12214,N_5453,N_6383);
or U12215 (N_12215,N_7820,N_9272);
and U12216 (N_12216,N_7427,N_9144);
and U12217 (N_12217,N_7278,N_8914);
nor U12218 (N_12218,N_5744,N_6284);
nand U12219 (N_12219,N_6465,N_5441);
nor U12220 (N_12220,N_5773,N_9323);
or U12221 (N_12221,N_6436,N_6969);
and U12222 (N_12222,N_8705,N_9782);
and U12223 (N_12223,N_5645,N_5227);
nor U12224 (N_12224,N_8244,N_7941);
nand U12225 (N_12225,N_9788,N_7340);
or U12226 (N_12226,N_8720,N_8370);
nor U12227 (N_12227,N_5379,N_8961);
nor U12228 (N_12228,N_5921,N_8067);
or U12229 (N_12229,N_8275,N_6708);
nand U12230 (N_12230,N_8118,N_7786);
nor U12231 (N_12231,N_9618,N_8119);
and U12232 (N_12232,N_6551,N_5931);
and U12233 (N_12233,N_9994,N_6361);
nor U12234 (N_12234,N_5608,N_8880);
nor U12235 (N_12235,N_8088,N_5222);
nor U12236 (N_12236,N_6954,N_6629);
and U12237 (N_12237,N_7038,N_8023);
nand U12238 (N_12238,N_9457,N_7680);
nand U12239 (N_12239,N_7977,N_9167);
nor U12240 (N_12240,N_5170,N_7013);
nor U12241 (N_12241,N_7956,N_6716);
nand U12242 (N_12242,N_8499,N_7699);
nor U12243 (N_12243,N_8960,N_9186);
or U12244 (N_12244,N_5044,N_8037);
or U12245 (N_12245,N_8853,N_7127);
and U12246 (N_12246,N_9468,N_5937);
and U12247 (N_12247,N_9918,N_6148);
nand U12248 (N_12248,N_6357,N_6720);
nand U12249 (N_12249,N_7676,N_6514);
nor U12250 (N_12250,N_5934,N_7651);
nor U12251 (N_12251,N_8928,N_6605);
nand U12252 (N_12252,N_9928,N_9942);
nand U12253 (N_12253,N_5375,N_9678);
nand U12254 (N_12254,N_9929,N_9155);
and U12255 (N_12255,N_6788,N_5857);
nor U12256 (N_12256,N_7722,N_5979);
and U12257 (N_12257,N_8454,N_9170);
and U12258 (N_12258,N_7473,N_8578);
nand U12259 (N_12259,N_6964,N_5718);
and U12260 (N_12260,N_6407,N_7122);
and U12261 (N_12261,N_5447,N_9262);
nand U12262 (N_12262,N_8576,N_8432);
or U12263 (N_12263,N_8402,N_5055);
nand U12264 (N_12264,N_5527,N_7932);
nor U12265 (N_12265,N_9242,N_6945);
nor U12266 (N_12266,N_6195,N_8934);
and U12267 (N_12267,N_6345,N_9712);
or U12268 (N_12268,N_8410,N_7263);
and U12269 (N_12269,N_8387,N_8059);
or U12270 (N_12270,N_9223,N_6098);
nand U12271 (N_12271,N_6568,N_8146);
and U12272 (N_12272,N_5516,N_6046);
and U12273 (N_12273,N_8256,N_6369);
or U12274 (N_12274,N_8566,N_8740);
or U12275 (N_12275,N_6702,N_7827);
nor U12276 (N_12276,N_9192,N_5093);
nand U12277 (N_12277,N_6077,N_7974);
and U12278 (N_12278,N_6228,N_8326);
and U12279 (N_12279,N_6440,N_7734);
and U12280 (N_12280,N_7395,N_7280);
and U12281 (N_12281,N_6037,N_8696);
nand U12282 (N_12282,N_9208,N_5404);
nor U12283 (N_12283,N_9841,N_9526);
nand U12284 (N_12284,N_8925,N_7326);
or U12285 (N_12285,N_9029,N_6567);
nor U12286 (N_12286,N_9497,N_8421);
nor U12287 (N_12287,N_7155,N_6787);
and U12288 (N_12288,N_7488,N_9304);
nor U12289 (N_12289,N_8667,N_9780);
and U12290 (N_12290,N_5420,N_8322);
nand U12291 (N_12291,N_7092,N_5063);
nor U12292 (N_12292,N_7351,N_8552);
or U12293 (N_12293,N_6507,N_7665);
or U12294 (N_12294,N_5940,N_5466);
nand U12295 (N_12295,N_5446,N_6892);
and U12296 (N_12296,N_9835,N_9063);
and U12297 (N_12297,N_5604,N_8131);
and U12298 (N_12298,N_5780,N_5632);
nand U12299 (N_12299,N_7045,N_7308);
nor U12300 (N_12300,N_8224,N_8130);
or U12301 (N_12301,N_6476,N_6924);
or U12302 (N_12302,N_5282,N_6519);
nor U12303 (N_12303,N_8749,N_7483);
or U12304 (N_12304,N_9422,N_7652);
or U12305 (N_12305,N_7103,N_6631);
nand U12306 (N_12306,N_8595,N_7132);
nand U12307 (N_12307,N_9374,N_9772);
nor U12308 (N_12308,N_9372,N_6358);
or U12309 (N_12309,N_9406,N_5971);
and U12310 (N_12310,N_7973,N_9012);
or U12311 (N_12311,N_9540,N_6707);
and U12312 (N_12312,N_8156,N_8309);
or U12313 (N_12313,N_5933,N_6322);
nor U12314 (N_12314,N_5755,N_5107);
nand U12315 (N_12315,N_5207,N_5024);
nand U12316 (N_12316,N_6266,N_9306);
and U12317 (N_12317,N_7679,N_6548);
or U12318 (N_12318,N_8461,N_6132);
or U12319 (N_12319,N_9505,N_9879);
nor U12320 (N_12320,N_9383,N_6204);
and U12321 (N_12321,N_9057,N_8184);
and U12322 (N_12322,N_8987,N_9220);
and U12323 (N_12323,N_6762,N_9486);
nand U12324 (N_12324,N_6669,N_6745);
or U12325 (N_12325,N_8698,N_5307);
nand U12326 (N_12326,N_7854,N_6715);
nor U12327 (N_12327,N_8114,N_6824);
or U12328 (N_12328,N_5260,N_8447);
or U12329 (N_12329,N_9435,N_6738);
nor U12330 (N_12330,N_9114,N_8069);
nand U12331 (N_12331,N_6661,N_5736);
nor U12332 (N_12332,N_5829,N_5852);
and U12333 (N_12333,N_7287,N_8475);
or U12334 (N_12334,N_5349,N_6757);
nor U12335 (N_12335,N_6947,N_5817);
and U12336 (N_12336,N_9581,N_5229);
nand U12337 (N_12337,N_8089,N_5266);
nand U12338 (N_12338,N_9023,N_5571);
and U12339 (N_12339,N_5623,N_7624);
xnor U12340 (N_12340,N_8524,N_8033);
or U12341 (N_12341,N_5621,N_8533);
or U12342 (N_12342,N_8352,N_7377);
nand U12343 (N_12343,N_7357,N_9649);
nor U12344 (N_12344,N_9142,N_6074);
or U12345 (N_12345,N_9599,N_9283);
nor U12346 (N_12346,N_5757,N_6025);
nand U12347 (N_12347,N_9778,N_7572);
and U12348 (N_12348,N_9962,N_5964);
nand U12349 (N_12349,N_9507,N_5650);
or U12350 (N_12350,N_7226,N_9740);
nor U12351 (N_12351,N_8999,N_9275);
nor U12352 (N_12352,N_7998,N_9039);
and U12353 (N_12353,N_5164,N_7279);
nor U12354 (N_12354,N_5607,N_8892);
nor U12355 (N_12355,N_6208,N_7532);
nand U12356 (N_12356,N_6367,N_8513);
nor U12357 (N_12357,N_6686,N_5109);
nand U12358 (N_12358,N_9239,N_8236);
nand U12359 (N_12359,N_9357,N_8218);
nand U12360 (N_12360,N_9988,N_5065);
nor U12361 (N_12361,N_5922,N_5676);
nand U12362 (N_12362,N_6784,N_6528);
nand U12363 (N_12363,N_7872,N_9769);
nand U12364 (N_12364,N_8484,N_9946);
nor U12365 (N_12365,N_6136,N_6265);
nand U12366 (N_12366,N_5722,N_6220);
nor U12367 (N_12367,N_7798,N_9798);
or U12368 (N_12368,N_5275,N_7981);
and U12369 (N_12369,N_5962,N_7539);
nor U12370 (N_12370,N_6161,N_8656);
nor U12371 (N_12371,N_7349,N_6347);
or U12372 (N_12372,N_9736,N_6871);
nor U12373 (N_12373,N_7968,N_6574);
or U12374 (N_12374,N_6931,N_8163);
nor U12375 (N_12375,N_7450,N_5497);
nor U12376 (N_12376,N_5019,N_7841);
and U12377 (N_12377,N_5657,N_6466);
nor U12378 (N_12378,N_5851,N_8197);
or U12379 (N_12379,N_5320,N_9887);
nor U12380 (N_12380,N_7476,N_7838);
nor U12381 (N_12381,N_9407,N_5983);
or U12382 (N_12382,N_5695,N_7962);
or U12383 (N_12383,N_8137,N_6191);
xnor U12384 (N_12384,N_9666,N_6826);
and U12385 (N_12385,N_5488,N_6344);
or U12386 (N_12386,N_9924,N_8417);
nor U12387 (N_12387,N_6783,N_5836);
nor U12388 (N_12388,N_7876,N_8856);
and U12389 (N_12389,N_7244,N_7586);
nor U12390 (N_12390,N_7026,N_6511);
nor U12391 (N_12391,N_6895,N_8145);
or U12392 (N_12392,N_9488,N_6019);
or U12393 (N_12393,N_6468,N_9389);
and U12394 (N_12394,N_5617,N_7446);
or U12395 (N_12395,N_5585,N_9626);
nand U12396 (N_12396,N_7000,N_7996);
and U12397 (N_12397,N_7477,N_5615);
or U12398 (N_12398,N_7205,N_7796);
nor U12399 (N_12399,N_7182,N_5901);
or U12400 (N_12400,N_7347,N_9642);
or U12401 (N_12401,N_8567,N_8430);
nor U12402 (N_12402,N_8268,N_6475);
or U12403 (N_12403,N_8652,N_6256);
or U12404 (N_12404,N_5876,N_8686);
and U12405 (N_12405,N_5021,N_9689);
and U12406 (N_12406,N_7406,N_5775);
and U12407 (N_12407,N_9358,N_9219);
nand U12408 (N_12408,N_7023,N_7445);
xor U12409 (N_12409,N_9956,N_9747);
nand U12410 (N_12410,N_5276,N_9444);
nor U12411 (N_12411,N_9388,N_5322);
nand U12412 (N_12412,N_8725,N_5997);
nor U12413 (N_12413,N_8345,N_8688);
nor U12414 (N_12414,N_8435,N_8143);
nand U12415 (N_12415,N_5716,N_5949);
nand U12416 (N_12416,N_7335,N_5652);
nand U12417 (N_12417,N_7400,N_9912);
nor U12418 (N_12418,N_5888,N_9432);
and U12419 (N_12419,N_5511,N_6461);
nand U12420 (N_12420,N_7836,N_8024);
nor U12421 (N_12421,N_5247,N_7125);
nor U12422 (N_12422,N_7402,N_8171);
or U12423 (N_12423,N_9687,N_5506);
and U12424 (N_12424,N_8028,N_6038);
nand U12425 (N_12425,N_7772,N_9564);
or U12426 (N_12426,N_7118,N_9248);
nor U12427 (N_12427,N_5195,N_8695);
nand U12428 (N_12428,N_9360,N_9831);
nand U12429 (N_12429,N_9866,N_5812);
nand U12430 (N_12430,N_5022,N_6129);
and U12431 (N_12431,N_6492,N_7044);
nor U12432 (N_12432,N_7887,N_6742);
and U12433 (N_12433,N_9396,N_7391);
or U12434 (N_12434,N_8831,N_6401);
or U12435 (N_12435,N_5287,N_8253);
nor U12436 (N_12436,N_9424,N_5785);
or U12437 (N_12437,N_5253,N_6342);
or U12438 (N_12438,N_5377,N_6450);
or U12439 (N_12439,N_8915,N_6058);
nor U12440 (N_12440,N_9749,N_7419);
nand U12441 (N_12441,N_5839,N_6168);
nor U12442 (N_12442,N_8469,N_7753);
xor U12443 (N_12443,N_8823,N_9176);
and U12444 (N_12444,N_6378,N_9810);
nand U12445 (N_12445,N_8170,N_7336);
and U12446 (N_12446,N_6264,N_5131);
nand U12447 (N_12447,N_7954,N_6442);
or U12448 (N_12448,N_5016,N_8388);
nor U12449 (N_12449,N_5932,N_9240);
and U12450 (N_12450,N_8983,N_9158);
and U12451 (N_12451,N_6681,N_6596);
or U12452 (N_12452,N_6249,N_6005);
or U12453 (N_12453,N_9255,N_5631);
nand U12454 (N_12454,N_7543,N_5161);
nand U12455 (N_12455,N_8035,N_7185);
and U12456 (N_12456,N_9795,N_8757);
or U12457 (N_12457,N_6086,N_6457);
nand U12458 (N_12458,N_6606,N_6163);
and U12459 (N_12459,N_6645,N_5064);
nand U12460 (N_12460,N_5508,N_9888);
and U12461 (N_12461,N_6141,N_9609);
nor U12462 (N_12462,N_8650,N_8825);
nand U12463 (N_12463,N_7582,N_7464);
nor U12464 (N_12464,N_8159,N_7161);
and U12465 (N_12465,N_8065,N_8743);
nand U12466 (N_12466,N_8030,N_5336);
nand U12467 (N_12467,N_8413,N_6175);
nor U12468 (N_12468,N_5442,N_5793);
and U12469 (N_12469,N_6812,N_5771);
nor U12470 (N_12470,N_7874,N_8883);
nand U12471 (N_12471,N_5694,N_5258);
nand U12472 (N_12472,N_7644,N_9475);
or U12473 (N_12473,N_9408,N_5843);
and U12474 (N_12474,N_9328,N_6471);
nand U12475 (N_12475,N_7142,N_7760);
nor U12476 (N_12476,N_6039,N_9399);
and U12477 (N_12477,N_8202,N_5728);
nor U12478 (N_12478,N_5154,N_9706);
nand U12479 (N_12479,N_6654,N_9600);
nand U12480 (N_12480,N_7538,N_7228);
or U12481 (N_12481,N_9905,N_9529);
nor U12482 (N_12482,N_6734,N_8451);
nand U12483 (N_12483,N_6930,N_9812);
or U12484 (N_12484,N_6472,N_6535);
and U12485 (N_12485,N_8147,N_6561);
or U12486 (N_12486,N_8265,N_6057);
and U12487 (N_12487,N_9318,N_9610);
nand U12488 (N_12488,N_8783,N_9892);
and U12489 (N_12489,N_9340,N_7965);
and U12490 (N_12490,N_8938,N_8538);
or U12491 (N_12491,N_5900,N_6160);
nor U12492 (N_12492,N_9375,N_9840);
nand U12493 (N_12493,N_6919,N_9447);
and U12494 (N_12494,N_5568,N_9755);
nand U12495 (N_12495,N_8393,N_6434);
or U12496 (N_12496,N_7756,N_6583);
nand U12497 (N_12497,N_6749,N_8654);
nand U12498 (N_12498,N_5174,N_6355);
nor U12499 (N_12499,N_6780,N_9979);
nand U12500 (N_12500,N_7642,N_6525);
or U12501 (N_12501,N_6503,N_6254);
and U12502 (N_12502,N_6313,N_8135);
nand U12503 (N_12503,N_8368,N_7566);
nand U12504 (N_12504,N_9103,N_7736);
nand U12505 (N_12505,N_8958,N_6826);
nand U12506 (N_12506,N_9330,N_9760);
or U12507 (N_12507,N_9776,N_7846);
nand U12508 (N_12508,N_9231,N_5236);
nor U12509 (N_12509,N_6828,N_5030);
nor U12510 (N_12510,N_6927,N_8212);
nand U12511 (N_12511,N_5661,N_9235);
nand U12512 (N_12512,N_6008,N_8919);
nand U12513 (N_12513,N_6646,N_6447);
or U12514 (N_12514,N_7998,N_9265);
or U12515 (N_12515,N_8799,N_5482);
nor U12516 (N_12516,N_9734,N_5029);
or U12517 (N_12517,N_8204,N_6691);
nand U12518 (N_12518,N_6459,N_5961);
or U12519 (N_12519,N_8049,N_8079);
or U12520 (N_12520,N_7362,N_7704);
or U12521 (N_12521,N_7517,N_5297);
nand U12522 (N_12522,N_9781,N_9778);
or U12523 (N_12523,N_5160,N_6356);
nor U12524 (N_12524,N_9398,N_5760);
nor U12525 (N_12525,N_8726,N_8547);
nor U12526 (N_12526,N_8824,N_9233);
nand U12527 (N_12527,N_5101,N_8543);
nor U12528 (N_12528,N_7278,N_5245);
nand U12529 (N_12529,N_8618,N_6727);
nor U12530 (N_12530,N_6364,N_9072);
nand U12531 (N_12531,N_7441,N_9697);
or U12532 (N_12532,N_6808,N_7321);
and U12533 (N_12533,N_7960,N_8592);
nor U12534 (N_12534,N_9200,N_7984);
nor U12535 (N_12535,N_8511,N_9270);
and U12536 (N_12536,N_5407,N_7998);
and U12537 (N_12537,N_5635,N_9876);
nor U12538 (N_12538,N_7494,N_7817);
and U12539 (N_12539,N_8703,N_5600);
nor U12540 (N_12540,N_6694,N_9304);
nand U12541 (N_12541,N_5414,N_7355);
nand U12542 (N_12542,N_8912,N_8039);
and U12543 (N_12543,N_7805,N_7521);
and U12544 (N_12544,N_9039,N_6551);
nand U12545 (N_12545,N_7093,N_6994);
nor U12546 (N_12546,N_9172,N_9238);
or U12547 (N_12547,N_6373,N_7497);
nor U12548 (N_12548,N_7896,N_8007);
nand U12549 (N_12549,N_7059,N_6514);
nand U12550 (N_12550,N_6587,N_9677);
nor U12551 (N_12551,N_5649,N_5059);
or U12552 (N_12552,N_9480,N_6389);
nor U12553 (N_12553,N_5326,N_9096);
or U12554 (N_12554,N_5759,N_9820);
nand U12555 (N_12555,N_7507,N_5133);
and U12556 (N_12556,N_5829,N_5850);
and U12557 (N_12557,N_8432,N_5798);
nand U12558 (N_12558,N_6803,N_8912);
nand U12559 (N_12559,N_5520,N_6589);
or U12560 (N_12560,N_5542,N_7152);
and U12561 (N_12561,N_5049,N_7774);
nor U12562 (N_12562,N_7977,N_9908);
nor U12563 (N_12563,N_9556,N_6219);
xnor U12564 (N_12564,N_9017,N_5131);
xnor U12565 (N_12565,N_5458,N_8770);
or U12566 (N_12566,N_9439,N_7968);
nand U12567 (N_12567,N_7463,N_8744);
nand U12568 (N_12568,N_7860,N_5757);
nor U12569 (N_12569,N_7335,N_6171);
nor U12570 (N_12570,N_9481,N_5844);
nand U12571 (N_12571,N_5817,N_8408);
nand U12572 (N_12572,N_7956,N_5277);
xnor U12573 (N_12573,N_8870,N_9425);
or U12574 (N_12574,N_9234,N_9747);
or U12575 (N_12575,N_8896,N_8534);
nand U12576 (N_12576,N_9666,N_7358);
or U12577 (N_12577,N_9126,N_7962);
and U12578 (N_12578,N_7865,N_9834);
and U12579 (N_12579,N_6455,N_9347);
and U12580 (N_12580,N_9330,N_5001);
and U12581 (N_12581,N_9168,N_8174);
and U12582 (N_12582,N_5222,N_9408);
or U12583 (N_12583,N_6556,N_9206);
nor U12584 (N_12584,N_5608,N_7440);
nand U12585 (N_12585,N_6477,N_6778);
nand U12586 (N_12586,N_9479,N_8060);
and U12587 (N_12587,N_9454,N_7422);
or U12588 (N_12588,N_7736,N_7255);
nand U12589 (N_12589,N_6717,N_5809);
and U12590 (N_12590,N_6682,N_6971);
and U12591 (N_12591,N_9797,N_7275);
and U12592 (N_12592,N_5888,N_6093);
nor U12593 (N_12593,N_6439,N_9494);
and U12594 (N_12594,N_6064,N_7934);
nand U12595 (N_12595,N_6575,N_8763);
or U12596 (N_12596,N_6157,N_8848);
xnor U12597 (N_12597,N_8532,N_5098);
and U12598 (N_12598,N_9237,N_9544);
and U12599 (N_12599,N_7582,N_7369);
nor U12600 (N_12600,N_7896,N_7488);
nor U12601 (N_12601,N_6052,N_8049);
or U12602 (N_12602,N_8064,N_8715);
or U12603 (N_12603,N_6660,N_7218);
nor U12604 (N_12604,N_6942,N_9001);
nor U12605 (N_12605,N_7900,N_7011);
nor U12606 (N_12606,N_7341,N_7030);
or U12607 (N_12607,N_7086,N_8379);
nor U12608 (N_12608,N_9923,N_9902);
nand U12609 (N_12609,N_6733,N_8644);
or U12610 (N_12610,N_5377,N_6544);
nand U12611 (N_12611,N_5633,N_9894);
nand U12612 (N_12612,N_7585,N_5403);
nand U12613 (N_12613,N_8335,N_7687);
nor U12614 (N_12614,N_9095,N_5000);
or U12615 (N_12615,N_8168,N_8912);
nor U12616 (N_12616,N_6931,N_6011);
or U12617 (N_12617,N_7650,N_8778);
nand U12618 (N_12618,N_8551,N_6556);
nand U12619 (N_12619,N_9133,N_7034);
nor U12620 (N_12620,N_9541,N_9398);
nor U12621 (N_12621,N_5192,N_6426);
or U12622 (N_12622,N_5162,N_7252);
and U12623 (N_12623,N_7500,N_7050);
nand U12624 (N_12624,N_9182,N_9559);
and U12625 (N_12625,N_6532,N_6702);
or U12626 (N_12626,N_5961,N_9002);
and U12627 (N_12627,N_6031,N_8581);
and U12628 (N_12628,N_9691,N_6395);
nand U12629 (N_12629,N_5866,N_9372);
and U12630 (N_12630,N_9698,N_8416);
and U12631 (N_12631,N_5871,N_5349);
nor U12632 (N_12632,N_5613,N_5626);
and U12633 (N_12633,N_6108,N_8390);
nand U12634 (N_12634,N_5471,N_6863);
and U12635 (N_12635,N_6810,N_8178);
or U12636 (N_12636,N_9860,N_5249);
xor U12637 (N_12637,N_6041,N_5915);
or U12638 (N_12638,N_8714,N_8937);
nand U12639 (N_12639,N_6949,N_8972);
and U12640 (N_12640,N_8857,N_8947);
nor U12641 (N_12641,N_7477,N_5691);
or U12642 (N_12642,N_8741,N_8357);
and U12643 (N_12643,N_8903,N_8818);
xor U12644 (N_12644,N_7023,N_9450);
or U12645 (N_12645,N_9857,N_5674);
or U12646 (N_12646,N_5856,N_5267);
nor U12647 (N_12647,N_9588,N_6507);
nand U12648 (N_12648,N_5138,N_7888);
and U12649 (N_12649,N_5740,N_5181);
or U12650 (N_12650,N_9841,N_8321);
or U12651 (N_12651,N_6035,N_7190);
nor U12652 (N_12652,N_9444,N_6494);
or U12653 (N_12653,N_9771,N_6350);
and U12654 (N_12654,N_9460,N_5606);
nor U12655 (N_12655,N_5815,N_7485);
nand U12656 (N_12656,N_9170,N_7749);
or U12657 (N_12657,N_7550,N_8401);
nor U12658 (N_12658,N_5553,N_6310);
or U12659 (N_12659,N_8332,N_5611);
or U12660 (N_12660,N_7765,N_6933);
nand U12661 (N_12661,N_9912,N_8746);
nor U12662 (N_12662,N_6383,N_6431);
or U12663 (N_12663,N_8083,N_6166);
and U12664 (N_12664,N_6518,N_6698);
nand U12665 (N_12665,N_9983,N_7904);
or U12666 (N_12666,N_6224,N_6701);
or U12667 (N_12667,N_6639,N_8957);
and U12668 (N_12668,N_9064,N_5842);
or U12669 (N_12669,N_5486,N_5072);
or U12670 (N_12670,N_7599,N_9772);
and U12671 (N_12671,N_8445,N_8595);
nand U12672 (N_12672,N_5901,N_8143);
nor U12673 (N_12673,N_8405,N_9776);
nand U12674 (N_12674,N_7925,N_6116);
and U12675 (N_12675,N_5357,N_9202);
and U12676 (N_12676,N_5012,N_6572);
nand U12677 (N_12677,N_6288,N_9943);
nand U12678 (N_12678,N_6731,N_6553);
xnor U12679 (N_12679,N_9965,N_7163);
and U12680 (N_12680,N_9816,N_8925);
nor U12681 (N_12681,N_5743,N_5547);
nand U12682 (N_12682,N_5679,N_5225);
nand U12683 (N_12683,N_9149,N_6939);
nand U12684 (N_12684,N_5323,N_8768);
nand U12685 (N_12685,N_8468,N_7920);
nand U12686 (N_12686,N_6506,N_5126);
nor U12687 (N_12687,N_9152,N_8467);
nor U12688 (N_12688,N_6938,N_6275);
or U12689 (N_12689,N_8218,N_8648);
or U12690 (N_12690,N_5270,N_9093);
nand U12691 (N_12691,N_7792,N_5291);
and U12692 (N_12692,N_9943,N_8081);
nand U12693 (N_12693,N_6338,N_5676);
nor U12694 (N_12694,N_9631,N_9821);
and U12695 (N_12695,N_8603,N_6468);
and U12696 (N_12696,N_8349,N_5692);
nor U12697 (N_12697,N_7149,N_8510);
or U12698 (N_12698,N_7635,N_6507);
and U12699 (N_12699,N_6611,N_6504);
or U12700 (N_12700,N_5007,N_7617);
and U12701 (N_12701,N_8129,N_7704);
or U12702 (N_12702,N_6981,N_5965);
nor U12703 (N_12703,N_5532,N_6157);
nand U12704 (N_12704,N_5788,N_9780);
nand U12705 (N_12705,N_9304,N_6411);
nor U12706 (N_12706,N_6536,N_7670);
or U12707 (N_12707,N_5007,N_6014);
and U12708 (N_12708,N_5247,N_5178);
nand U12709 (N_12709,N_6726,N_8139);
and U12710 (N_12710,N_6924,N_6767);
nor U12711 (N_12711,N_5397,N_8221);
nand U12712 (N_12712,N_5474,N_6812);
or U12713 (N_12713,N_7318,N_9160);
and U12714 (N_12714,N_6891,N_6628);
nand U12715 (N_12715,N_7784,N_6766);
nor U12716 (N_12716,N_6335,N_7047);
or U12717 (N_12717,N_9118,N_8322);
nand U12718 (N_12718,N_9350,N_9424);
nand U12719 (N_12719,N_5208,N_9595);
or U12720 (N_12720,N_6631,N_7195);
nand U12721 (N_12721,N_9005,N_7192);
or U12722 (N_12722,N_9529,N_8624);
and U12723 (N_12723,N_7061,N_6869);
and U12724 (N_12724,N_9096,N_5622);
or U12725 (N_12725,N_8414,N_5075);
nand U12726 (N_12726,N_8948,N_7645);
or U12727 (N_12727,N_7445,N_6073);
and U12728 (N_12728,N_7884,N_5586);
or U12729 (N_12729,N_7922,N_5639);
nand U12730 (N_12730,N_5543,N_6128);
nor U12731 (N_12731,N_5847,N_9962);
nor U12732 (N_12732,N_7540,N_9513);
nor U12733 (N_12733,N_6454,N_9913);
and U12734 (N_12734,N_9336,N_6984);
and U12735 (N_12735,N_6358,N_6892);
or U12736 (N_12736,N_7314,N_6339);
or U12737 (N_12737,N_8241,N_8326);
and U12738 (N_12738,N_8093,N_7785);
nor U12739 (N_12739,N_8746,N_7418);
nand U12740 (N_12740,N_7575,N_8672);
nand U12741 (N_12741,N_9349,N_9736);
nand U12742 (N_12742,N_5069,N_7972);
nor U12743 (N_12743,N_9641,N_8983);
nand U12744 (N_12744,N_5376,N_5607);
or U12745 (N_12745,N_8594,N_7782);
and U12746 (N_12746,N_9564,N_7740);
and U12747 (N_12747,N_5307,N_5513);
and U12748 (N_12748,N_8214,N_6347);
xnor U12749 (N_12749,N_9610,N_9842);
nand U12750 (N_12750,N_5183,N_5075);
and U12751 (N_12751,N_7405,N_9283);
nand U12752 (N_12752,N_6823,N_6034);
or U12753 (N_12753,N_5742,N_8502);
or U12754 (N_12754,N_7391,N_5511);
nand U12755 (N_12755,N_7655,N_6024);
nand U12756 (N_12756,N_6241,N_6028);
nand U12757 (N_12757,N_7473,N_7654);
xnor U12758 (N_12758,N_9650,N_6176);
or U12759 (N_12759,N_6225,N_7487);
or U12760 (N_12760,N_7219,N_9891);
nand U12761 (N_12761,N_8405,N_6562);
nand U12762 (N_12762,N_8991,N_5718);
nor U12763 (N_12763,N_5281,N_6671);
or U12764 (N_12764,N_9331,N_8280);
or U12765 (N_12765,N_8830,N_9310);
nand U12766 (N_12766,N_5000,N_5616);
and U12767 (N_12767,N_9163,N_6485);
or U12768 (N_12768,N_7871,N_9657);
nor U12769 (N_12769,N_6669,N_8466);
and U12770 (N_12770,N_6310,N_5568);
nor U12771 (N_12771,N_9290,N_7104);
and U12772 (N_12772,N_5586,N_8526);
or U12773 (N_12773,N_9118,N_5385);
or U12774 (N_12774,N_5870,N_8439);
or U12775 (N_12775,N_9493,N_7244);
nand U12776 (N_12776,N_6147,N_6835);
or U12777 (N_12777,N_7266,N_9335);
nand U12778 (N_12778,N_8634,N_6477);
and U12779 (N_12779,N_9634,N_9288);
and U12780 (N_12780,N_8321,N_6510);
and U12781 (N_12781,N_5525,N_9432);
nor U12782 (N_12782,N_8393,N_7474);
nor U12783 (N_12783,N_6674,N_5455);
or U12784 (N_12784,N_6304,N_9313);
or U12785 (N_12785,N_5034,N_8276);
and U12786 (N_12786,N_9976,N_7950);
nand U12787 (N_12787,N_5330,N_8031);
or U12788 (N_12788,N_9818,N_7411);
and U12789 (N_12789,N_7912,N_8217);
nor U12790 (N_12790,N_7786,N_6189);
nor U12791 (N_12791,N_8441,N_7706);
nor U12792 (N_12792,N_9515,N_5102);
nor U12793 (N_12793,N_6510,N_8930);
and U12794 (N_12794,N_8807,N_9641);
or U12795 (N_12795,N_7690,N_8843);
nand U12796 (N_12796,N_5110,N_7795);
or U12797 (N_12797,N_9315,N_8948);
nor U12798 (N_12798,N_7043,N_6200);
nand U12799 (N_12799,N_6957,N_7945);
and U12800 (N_12800,N_7916,N_8375);
or U12801 (N_12801,N_6791,N_7955);
nand U12802 (N_12802,N_6830,N_5818);
nor U12803 (N_12803,N_7968,N_6571);
nor U12804 (N_12804,N_9696,N_5645);
nand U12805 (N_12805,N_7505,N_6639);
and U12806 (N_12806,N_9432,N_8099);
and U12807 (N_12807,N_9880,N_6390);
or U12808 (N_12808,N_6697,N_8428);
and U12809 (N_12809,N_7867,N_5730);
nand U12810 (N_12810,N_5205,N_5543);
or U12811 (N_12811,N_6482,N_9227);
nor U12812 (N_12812,N_7164,N_7824);
or U12813 (N_12813,N_5768,N_5107);
nor U12814 (N_12814,N_6986,N_9679);
nor U12815 (N_12815,N_5311,N_9965);
or U12816 (N_12816,N_6408,N_8622);
and U12817 (N_12817,N_6347,N_5083);
nor U12818 (N_12818,N_9451,N_6839);
nand U12819 (N_12819,N_5593,N_7989);
nand U12820 (N_12820,N_8220,N_9640);
nand U12821 (N_12821,N_6888,N_9701);
and U12822 (N_12822,N_8366,N_5312);
nand U12823 (N_12823,N_8648,N_8798);
nand U12824 (N_12824,N_7607,N_5193);
nand U12825 (N_12825,N_7832,N_7830);
nor U12826 (N_12826,N_6621,N_6518);
and U12827 (N_12827,N_6464,N_7554);
nor U12828 (N_12828,N_7535,N_8359);
or U12829 (N_12829,N_5912,N_6431);
nor U12830 (N_12830,N_5109,N_5173);
and U12831 (N_12831,N_7347,N_9189);
or U12832 (N_12832,N_5250,N_6084);
or U12833 (N_12833,N_9629,N_5109);
nand U12834 (N_12834,N_6061,N_7015);
nor U12835 (N_12835,N_9210,N_8357);
and U12836 (N_12836,N_9308,N_6885);
or U12837 (N_12837,N_6051,N_9757);
and U12838 (N_12838,N_6994,N_8870);
or U12839 (N_12839,N_7155,N_5684);
or U12840 (N_12840,N_6303,N_8560);
nor U12841 (N_12841,N_9186,N_5253);
nor U12842 (N_12842,N_5093,N_6950);
nand U12843 (N_12843,N_5317,N_9416);
nor U12844 (N_12844,N_8324,N_8323);
nor U12845 (N_12845,N_5429,N_5144);
and U12846 (N_12846,N_5491,N_5302);
or U12847 (N_12847,N_9547,N_6121);
or U12848 (N_12848,N_5705,N_5925);
and U12849 (N_12849,N_9290,N_6318);
or U12850 (N_12850,N_7562,N_7748);
and U12851 (N_12851,N_7251,N_9021);
and U12852 (N_12852,N_9649,N_9985);
nor U12853 (N_12853,N_5468,N_6927);
and U12854 (N_12854,N_5156,N_7848);
nand U12855 (N_12855,N_9309,N_5182);
nand U12856 (N_12856,N_8444,N_5716);
and U12857 (N_12857,N_8269,N_6939);
nor U12858 (N_12858,N_6466,N_5741);
or U12859 (N_12859,N_8868,N_7086);
and U12860 (N_12860,N_8085,N_7290);
and U12861 (N_12861,N_9550,N_6097);
and U12862 (N_12862,N_5709,N_5661);
nor U12863 (N_12863,N_7996,N_5475);
nand U12864 (N_12864,N_7946,N_6293);
nor U12865 (N_12865,N_9108,N_9293);
or U12866 (N_12866,N_9373,N_8027);
nand U12867 (N_12867,N_8542,N_6250);
or U12868 (N_12868,N_5052,N_7118);
nand U12869 (N_12869,N_5345,N_7987);
or U12870 (N_12870,N_8329,N_6247);
and U12871 (N_12871,N_9059,N_8106);
or U12872 (N_12872,N_8754,N_8182);
nand U12873 (N_12873,N_5525,N_5300);
nor U12874 (N_12874,N_5755,N_6647);
nor U12875 (N_12875,N_6400,N_6232);
nand U12876 (N_12876,N_5258,N_7788);
or U12877 (N_12877,N_8657,N_9493);
nor U12878 (N_12878,N_8413,N_8285);
nor U12879 (N_12879,N_6537,N_7535);
nor U12880 (N_12880,N_7726,N_5077);
nor U12881 (N_12881,N_9695,N_8105);
xor U12882 (N_12882,N_9698,N_5208);
and U12883 (N_12883,N_9651,N_7572);
nor U12884 (N_12884,N_7111,N_5483);
nand U12885 (N_12885,N_9665,N_7208);
nand U12886 (N_12886,N_8539,N_8786);
or U12887 (N_12887,N_7837,N_5521);
and U12888 (N_12888,N_5573,N_9944);
nand U12889 (N_12889,N_5720,N_7414);
nand U12890 (N_12890,N_5310,N_9183);
or U12891 (N_12891,N_8009,N_8597);
nor U12892 (N_12892,N_5741,N_7894);
and U12893 (N_12893,N_9976,N_9211);
and U12894 (N_12894,N_7326,N_8748);
nor U12895 (N_12895,N_7555,N_6692);
nand U12896 (N_12896,N_6116,N_6750);
and U12897 (N_12897,N_9732,N_5933);
and U12898 (N_12898,N_6390,N_5806);
nor U12899 (N_12899,N_5652,N_7398);
nand U12900 (N_12900,N_7637,N_6449);
and U12901 (N_12901,N_8352,N_8278);
nor U12902 (N_12902,N_5086,N_8179);
nor U12903 (N_12903,N_6812,N_5588);
nor U12904 (N_12904,N_8722,N_5438);
nand U12905 (N_12905,N_7530,N_9601);
nand U12906 (N_12906,N_8928,N_7667);
nor U12907 (N_12907,N_6381,N_5400);
nand U12908 (N_12908,N_5402,N_7236);
or U12909 (N_12909,N_5030,N_8942);
nand U12910 (N_12910,N_5739,N_5285);
nand U12911 (N_12911,N_9396,N_6979);
nor U12912 (N_12912,N_9870,N_5548);
nor U12913 (N_12913,N_5796,N_7118);
and U12914 (N_12914,N_9011,N_8092);
nor U12915 (N_12915,N_6142,N_6610);
nand U12916 (N_12916,N_8309,N_6063);
nand U12917 (N_12917,N_9027,N_6643);
and U12918 (N_12918,N_5518,N_9823);
and U12919 (N_12919,N_5061,N_5107);
nand U12920 (N_12920,N_9360,N_7490);
nand U12921 (N_12921,N_5230,N_8841);
nor U12922 (N_12922,N_6435,N_8745);
and U12923 (N_12923,N_8573,N_7199);
and U12924 (N_12924,N_7164,N_5630);
or U12925 (N_12925,N_7160,N_9508);
nor U12926 (N_12926,N_8598,N_5013);
nor U12927 (N_12927,N_9943,N_5902);
and U12928 (N_12928,N_6939,N_7711);
and U12929 (N_12929,N_5310,N_7965);
nor U12930 (N_12930,N_7096,N_9152);
nor U12931 (N_12931,N_7323,N_7142);
xnor U12932 (N_12932,N_7481,N_5131);
nor U12933 (N_12933,N_5866,N_9734);
and U12934 (N_12934,N_8120,N_5687);
nand U12935 (N_12935,N_7901,N_6090);
nor U12936 (N_12936,N_7385,N_7092);
and U12937 (N_12937,N_8338,N_6893);
and U12938 (N_12938,N_8433,N_9186);
nand U12939 (N_12939,N_9734,N_8103);
nand U12940 (N_12940,N_7958,N_8409);
and U12941 (N_12941,N_6771,N_9704);
or U12942 (N_12942,N_6544,N_9719);
or U12943 (N_12943,N_7503,N_8064);
and U12944 (N_12944,N_7391,N_8216);
and U12945 (N_12945,N_8473,N_8600);
or U12946 (N_12946,N_6931,N_7093);
nor U12947 (N_12947,N_5792,N_9244);
nand U12948 (N_12948,N_6474,N_7293);
and U12949 (N_12949,N_7799,N_6962);
nand U12950 (N_12950,N_8412,N_9730);
or U12951 (N_12951,N_7727,N_8548);
and U12952 (N_12952,N_7883,N_6002);
or U12953 (N_12953,N_7158,N_9705);
xor U12954 (N_12954,N_5815,N_8885);
and U12955 (N_12955,N_5538,N_8486);
and U12956 (N_12956,N_8413,N_7719);
or U12957 (N_12957,N_9602,N_6831);
nand U12958 (N_12958,N_6766,N_7263);
and U12959 (N_12959,N_7667,N_8692);
nor U12960 (N_12960,N_6513,N_8987);
nand U12961 (N_12961,N_5927,N_7135);
nor U12962 (N_12962,N_5071,N_8988);
or U12963 (N_12963,N_6170,N_7949);
or U12964 (N_12964,N_5704,N_6342);
nor U12965 (N_12965,N_6640,N_9372);
nor U12966 (N_12966,N_5262,N_5967);
and U12967 (N_12967,N_6684,N_8476);
or U12968 (N_12968,N_8638,N_6082);
and U12969 (N_12969,N_6088,N_9434);
and U12970 (N_12970,N_6108,N_8207);
or U12971 (N_12971,N_5509,N_6185);
or U12972 (N_12972,N_6530,N_9571);
nand U12973 (N_12973,N_6108,N_5425);
nor U12974 (N_12974,N_9453,N_7395);
and U12975 (N_12975,N_8380,N_7415);
and U12976 (N_12976,N_9960,N_7905);
or U12977 (N_12977,N_6298,N_7675);
nor U12978 (N_12978,N_6932,N_6275);
nand U12979 (N_12979,N_5038,N_9016);
or U12980 (N_12980,N_8037,N_5793);
or U12981 (N_12981,N_7835,N_8924);
nor U12982 (N_12982,N_7292,N_9552);
or U12983 (N_12983,N_9954,N_6663);
or U12984 (N_12984,N_5194,N_5324);
or U12985 (N_12985,N_6679,N_6111);
nand U12986 (N_12986,N_8331,N_9208);
nor U12987 (N_12987,N_7640,N_6880);
nor U12988 (N_12988,N_5183,N_9368);
nor U12989 (N_12989,N_5542,N_5014);
nor U12990 (N_12990,N_8743,N_6316);
nand U12991 (N_12991,N_8945,N_8597);
nor U12992 (N_12992,N_8887,N_9322);
nand U12993 (N_12993,N_9325,N_5995);
and U12994 (N_12994,N_5978,N_6855);
nand U12995 (N_12995,N_5069,N_6187);
nand U12996 (N_12996,N_6931,N_8785);
nor U12997 (N_12997,N_9568,N_9464);
or U12998 (N_12998,N_5270,N_9567);
or U12999 (N_12999,N_9012,N_9667);
nor U13000 (N_13000,N_9858,N_7122);
and U13001 (N_13001,N_9775,N_9580);
nand U13002 (N_13002,N_6128,N_8029);
nand U13003 (N_13003,N_6318,N_7654);
nor U13004 (N_13004,N_8649,N_5118);
nand U13005 (N_13005,N_8251,N_9841);
or U13006 (N_13006,N_5877,N_7055);
and U13007 (N_13007,N_5625,N_9630);
or U13008 (N_13008,N_6746,N_9075);
nand U13009 (N_13009,N_9830,N_5283);
nand U13010 (N_13010,N_5490,N_7051);
nand U13011 (N_13011,N_8873,N_9674);
nor U13012 (N_13012,N_9403,N_9580);
nor U13013 (N_13013,N_8217,N_7181);
nand U13014 (N_13014,N_5726,N_7434);
nor U13015 (N_13015,N_8053,N_9094);
nand U13016 (N_13016,N_5503,N_8347);
nand U13017 (N_13017,N_5628,N_5802);
or U13018 (N_13018,N_6000,N_7757);
nand U13019 (N_13019,N_7178,N_9902);
or U13020 (N_13020,N_6968,N_8648);
and U13021 (N_13021,N_5698,N_8026);
or U13022 (N_13022,N_6447,N_5442);
or U13023 (N_13023,N_9477,N_9082);
nor U13024 (N_13024,N_6147,N_8155);
nand U13025 (N_13025,N_6416,N_6169);
nor U13026 (N_13026,N_7566,N_9573);
or U13027 (N_13027,N_7479,N_5951);
or U13028 (N_13028,N_9873,N_6360);
or U13029 (N_13029,N_6716,N_7826);
and U13030 (N_13030,N_5425,N_8213);
nand U13031 (N_13031,N_6339,N_6148);
nand U13032 (N_13032,N_6345,N_9971);
and U13033 (N_13033,N_6608,N_8087);
and U13034 (N_13034,N_5260,N_6566);
or U13035 (N_13035,N_6587,N_8323);
and U13036 (N_13036,N_8110,N_8309);
nand U13037 (N_13037,N_7383,N_6131);
or U13038 (N_13038,N_8859,N_5411);
or U13039 (N_13039,N_7610,N_8938);
nor U13040 (N_13040,N_5229,N_7782);
nor U13041 (N_13041,N_6551,N_8226);
and U13042 (N_13042,N_8000,N_5568);
nor U13043 (N_13043,N_8809,N_5811);
and U13044 (N_13044,N_9316,N_5224);
and U13045 (N_13045,N_7494,N_8403);
and U13046 (N_13046,N_7559,N_8327);
or U13047 (N_13047,N_6259,N_7472);
and U13048 (N_13048,N_9440,N_7851);
or U13049 (N_13049,N_7393,N_7159);
nand U13050 (N_13050,N_7877,N_7314);
nand U13051 (N_13051,N_6640,N_9629);
and U13052 (N_13052,N_8228,N_9898);
and U13053 (N_13053,N_9345,N_9080);
nor U13054 (N_13054,N_8071,N_8471);
nand U13055 (N_13055,N_5395,N_6400);
nor U13056 (N_13056,N_6481,N_8166);
and U13057 (N_13057,N_9420,N_6130);
nand U13058 (N_13058,N_5290,N_7973);
and U13059 (N_13059,N_9884,N_6567);
nor U13060 (N_13060,N_8861,N_8623);
nor U13061 (N_13061,N_5953,N_7792);
nor U13062 (N_13062,N_8319,N_8546);
or U13063 (N_13063,N_7602,N_8484);
nor U13064 (N_13064,N_6863,N_5103);
or U13065 (N_13065,N_5556,N_7347);
or U13066 (N_13066,N_5579,N_7858);
and U13067 (N_13067,N_6686,N_8344);
nor U13068 (N_13068,N_7094,N_6273);
and U13069 (N_13069,N_8225,N_8880);
or U13070 (N_13070,N_9897,N_8890);
nor U13071 (N_13071,N_6530,N_9596);
nor U13072 (N_13072,N_6238,N_6713);
nor U13073 (N_13073,N_9516,N_6713);
nor U13074 (N_13074,N_5328,N_5316);
or U13075 (N_13075,N_8486,N_7115);
or U13076 (N_13076,N_9363,N_7652);
and U13077 (N_13077,N_9846,N_6650);
nand U13078 (N_13078,N_5660,N_9410);
and U13079 (N_13079,N_9383,N_6389);
nand U13080 (N_13080,N_9265,N_6564);
or U13081 (N_13081,N_7515,N_5468);
nand U13082 (N_13082,N_8528,N_6340);
or U13083 (N_13083,N_9481,N_8013);
and U13084 (N_13084,N_9092,N_8129);
nor U13085 (N_13085,N_5399,N_6360);
nor U13086 (N_13086,N_8029,N_6462);
xnor U13087 (N_13087,N_6724,N_8197);
and U13088 (N_13088,N_5317,N_6490);
and U13089 (N_13089,N_6132,N_6312);
or U13090 (N_13090,N_9997,N_7476);
nor U13091 (N_13091,N_8766,N_9854);
or U13092 (N_13092,N_8714,N_5050);
and U13093 (N_13093,N_8801,N_9655);
nand U13094 (N_13094,N_8711,N_7430);
or U13095 (N_13095,N_6752,N_9851);
and U13096 (N_13096,N_6338,N_9506);
nand U13097 (N_13097,N_7307,N_6865);
nor U13098 (N_13098,N_6727,N_6870);
and U13099 (N_13099,N_8840,N_9299);
and U13100 (N_13100,N_5537,N_6233);
or U13101 (N_13101,N_9170,N_6658);
or U13102 (N_13102,N_8855,N_9653);
or U13103 (N_13103,N_8412,N_8568);
and U13104 (N_13104,N_7586,N_6434);
nand U13105 (N_13105,N_7043,N_8973);
nand U13106 (N_13106,N_5128,N_5503);
and U13107 (N_13107,N_9352,N_6356);
or U13108 (N_13108,N_7737,N_9939);
nand U13109 (N_13109,N_6661,N_8032);
nand U13110 (N_13110,N_7786,N_8346);
nand U13111 (N_13111,N_5412,N_6304);
nor U13112 (N_13112,N_7494,N_5712);
and U13113 (N_13113,N_8420,N_6662);
nor U13114 (N_13114,N_8970,N_9756);
and U13115 (N_13115,N_9309,N_9093);
nor U13116 (N_13116,N_8823,N_6162);
nand U13117 (N_13117,N_8363,N_5151);
and U13118 (N_13118,N_8602,N_6009);
or U13119 (N_13119,N_7111,N_5027);
or U13120 (N_13120,N_7369,N_7473);
nand U13121 (N_13121,N_6430,N_5626);
nor U13122 (N_13122,N_7511,N_6064);
nor U13123 (N_13123,N_7341,N_6914);
or U13124 (N_13124,N_6459,N_7632);
or U13125 (N_13125,N_5475,N_6041);
and U13126 (N_13126,N_8156,N_9498);
nand U13127 (N_13127,N_5004,N_6871);
and U13128 (N_13128,N_5475,N_5287);
nand U13129 (N_13129,N_9602,N_9512);
and U13130 (N_13130,N_9063,N_9776);
nand U13131 (N_13131,N_8935,N_9660);
and U13132 (N_13132,N_8218,N_5963);
nand U13133 (N_13133,N_9350,N_5035);
nand U13134 (N_13134,N_5332,N_7795);
nand U13135 (N_13135,N_9222,N_8534);
nand U13136 (N_13136,N_9884,N_6632);
and U13137 (N_13137,N_5061,N_5855);
or U13138 (N_13138,N_5272,N_9695);
nand U13139 (N_13139,N_8843,N_9642);
and U13140 (N_13140,N_7543,N_7796);
nand U13141 (N_13141,N_9261,N_9285);
and U13142 (N_13142,N_8761,N_6338);
and U13143 (N_13143,N_5181,N_7884);
nor U13144 (N_13144,N_7080,N_7329);
nand U13145 (N_13145,N_7782,N_6368);
nor U13146 (N_13146,N_6088,N_9994);
or U13147 (N_13147,N_7074,N_7358);
and U13148 (N_13148,N_5507,N_7733);
nand U13149 (N_13149,N_8685,N_8402);
or U13150 (N_13150,N_6702,N_9785);
nor U13151 (N_13151,N_7840,N_6788);
nor U13152 (N_13152,N_9453,N_7067);
and U13153 (N_13153,N_9958,N_8625);
nor U13154 (N_13154,N_6382,N_9222);
nand U13155 (N_13155,N_6860,N_9557);
and U13156 (N_13156,N_8753,N_8171);
and U13157 (N_13157,N_8948,N_9720);
nand U13158 (N_13158,N_9540,N_6649);
or U13159 (N_13159,N_5199,N_7819);
nand U13160 (N_13160,N_7170,N_9886);
nand U13161 (N_13161,N_7264,N_8005);
or U13162 (N_13162,N_9885,N_7551);
nand U13163 (N_13163,N_7392,N_5418);
or U13164 (N_13164,N_6510,N_6144);
or U13165 (N_13165,N_7423,N_7147);
or U13166 (N_13166,N_9984,N_5243);
and U13167 (N_13167,N_6975,N_6341);
xor U13168 (N_13168,N_6647,N_6964);
nand U13169 (N_13169,N_8421,N_9750);
and U13170 (N_13170,N_7357,N_5752);
and U13171 (N_13171,N_8230,N_9947);
or U13172 (N_13172,N_9692,N_6200);
or U13173 (N_13173,N_5213,N_9200);
and U13174 (N_13174,N_5619,N_7379);
nand U13175 (N_13175,N_6300,N_9523);
and U13176 (N_13176,N_7448,N_9226);
nor U13177 (N_13177,N_7905,N_8955);
xnor U13178 (N_13178,N_7607,N_7550);
and U13179 (N_13179,N_8975,N_6395);
nor U13180 (N_13180,N_6912,N_5469);
and U13181 (N_13181,N_5910,N_6345);
nand U13182 (N_13182,N_5362,N_7724);
nor U13183 (N_13183,N_8679,N_8026);
nor U13184 (N_13184,N_9914,N_7743);
or U13185 (N_13185,N_8202,N_6827);
or U13186 (N_13186,N_8595,N_9877);
nor U13187 (N_13187,N_9840,N_9915);
and U13188 (N_13188,N_5365,N_5955);
nor U13189 (N_13189,N_8759,N_5809);
nand U13190 (N_13190,N_5888,N_9365);
nand U13191 (N_13191,N_9769,N_9212);
or U13192 (N_13192,N_6587,N_7891);
or U13193 (N_13193,N_8575,N_9656);
and U13194 (N_13194,N_7131,N_9031);
and U13195 (N_13195,N_9476,N_8749);
and U13196 (N_13196,N_5758,N_5407);
nand U13197 (N_13197,N_9374,N_6321);
and U13198 (N_13198,N_9140,N_7803);
nor U13199 (N_13199,N_8977,N_6257);
nor U13200 (N_13200,N_8019,N_7643);
nor U13201 (N_13201,N_8316,N_6192);
nand U13202 (N_13202,N_9006,N_9127);
and U13203 (N_13203,N_9277,N_6802);
or U13204 (N_13204,N_9727,N_6915);
and U13205 (N_13205,N_8071,N_9205);
nand U13206 (N_13206,N_5754,N_6991);
nor U13207 (N_13207,N_8978,N_9328);
or U13208 (N_13208,N_8124,N_9962);
and U13209 (N_13209,N_9311,N_7476);
nor U13210 (N_13210,N_9800,N_9632);
nor U13211 (N_13211,N_7419,N_7672);
and U13212 (N_13212,N_8563,N_5772);
nand U13213 (N_13213,N_7454,N_5023);
nor U13214 (N_13214,N_9430,N_6569);
nand U13215 (N_13215,N_6156,N_8327);
and U13216 (N_13216,N_5845,N_5420);
nand U13217 (N_13217,N_8587,N_5800);
and U13218 (N_13218,N_9846,N_5342);
nand U13219 (N_13219,N_5852,N_7995);
nand U13220 (N_13220,N_8922,N_8291);
nand U13221 (N_13221,N_7104,N_7172);
or U13222 (N_13222,N_7959,N_9633);
or U13223 (N_13223,N_8692,N_9997);
or U13224 (N_13224,N_7986,N_5622);
nand U13225 (N_13225,N_9702,N_8156);
and U13226 (N_13226,N_9686,N_6152);
and U13227 (N_13227,N_7244,N_6414);
xor U13228 (N_13228,N_9964,N_6012);
nor U13229 (N_13229,N_6284,N_5146);
nor U13230 (N_13230,N_7829,N_7387);
or U13231 (N_13231,N_7186,N_8668);
and U13232 (N_13232,N_5908,N_6058);
and U13233 (N_13233,N_9147,N_8874);
or U13234 (N_13234,N_6906,N_6615);
or U13235 (N_13235,N_9987,N_9632);
nand U13236 (N_13236,N_6296,N_8973);
or U13237 (N_13237,N_5083,N_5033);
nand U13238 (N_13238,N_6376,N_6807);
or U13239 (N_13239,N_7735,N_5492);
nor U13240 (N_13240,N_5658,N_8005);
and U13241 (N_13241,N_5959,N_7018);
and U13242 (N_13242,N_8258,N_8506);
nand U13243 (N_13243,N_7534,N_5139);
nor U13244 (N_13244,N_9420,N_8027);
nand U13245 (N_13245,N_6622,N_9562);
and U13246 (N_13246,N_5991,N_7898);
and U13247 (N_13247,N_8341,N_9969);
or U13248 (N_13248,N_5731,N_9784);
nand U13249 (N_13249,N_7822,N_8052);
xor U13250 (N_13250,N_7975,N_9242);
and U13251 (N_13251,N_6972,N_9533);
nand U13252 (N_13252,N_7562,N_9862);
nor U13253 (N_13253,N_8920,N_9915);
and U13254 (N_13254,N_6278,N_7056);
nand U13255 (N_13255,N_6687,N_6451);
or U13256 (N_13256,N_8386,N_9138);
nand U13257 (N_13257,N_9188,N_8368);
and U13258 (N_13258,N_7414,N_8274);
nor U13259 (N_13259,N_7241,N_5207);
and U13260 (N_13260,N_8120,N_6629);
nor U13261 (N_13261,N_5430,N_6285);
or U13262 (N_13262,N_7617,N_8509);
nand U13263 (N_13263,N_6768,N_7096);
and U13264 (N_13264,N_8985,N_9140);
or U13265 (N_13265,N_9426,N_8362);
and U13266 (N_13266,N_7865,N_7293);
and U13267 (N_13267,N_6184,N_6753);
or U13268 (N_13268,N_6990,N_7432);
nand U13269 (N_13269,N_9835,N_7864);
and U13270 (N_13270,N_5970,N_6075);
nand U13271 (N_13271,N_5458,N_5728);
or U13272 (N_13272,N_8014,N_5447);
and U13273 (N_13273,N_9909,N_9403);
and U13274 (N_13274,N_5188,N_5049);
and U13275 (N_13275,N_8885,N_7134);
and U13276 (N_13276,N_9790,N_9806);
nand U13277 (N_13277,N_9732,N_7920);
or U13278 (N_13278,N_6778,N_9499);
nand U13279 (N_13279,N_8970,N_6688);
or U13280 (N_13280,N_6106,N_8527);
nor U13281 (N_13281,N_5538,N_7038);
and U13282 (N_13282,N_5819,N_5857);
or U13283 (N_13283,N_6217,N_7321);
nor U13284 (N_13284,N_9810,N_8415);
nand U13285 (N_13285,N_9480,N_9937);
and U13286 (N_13286,N_5293,N_7041);
and U13287 (N_13287,N_8781,N_7195);
or U13288 (N_13288,N_8312,N_9940);
and U13289 (N_13289,N_9176,N_5585);
nand U13290 (N_13290,N_6539,N_5067);
nor U13291 (N_13291,N_8824,N_5590);
nor U13292 (N_13292,N_6826,N_5658);
nor U13293 (N_13293,N_8908,N_6036);
nor U13294 (N_13294,N_6421,N_8416);
or U13295 (N_13295,N_7742,N_5962);
nand U13296 (N_13296,N_9975,N_9756);
and U13297 (N_13297,N_7975,N_5659);
nor U13298 (N_13298,N_7225,N_6378);
nor U13299 (N_13299,N_8062,N_7123);
and U13300 (N_13300,N_6399,N_6728);
xnor U13301 (N_13301,N_9883,N_5190);
nand U13302 (N_13302,N_6666,N_5870);
or U13303 (N_13303,N_9243,N_5934);
nand U13304 (N_13304,N_7733,N_5046);
and U13305 (N_13305,N_7505,N_5149);
and U13306 (N_13306,N_6974,N_9984);
nand U13307 (N_13307,N_7501,N_8305);
or U13308 (N_13308,N_9528,N_7178);
nor U13309 (N_13309,N_6967,N_7664);
or U13310 (N_13310,N_7076,N_8443);
nand U13311 (N_13311,N_8118,N_6041);
nor U13312 (N_13312,N_5367,N_7303);
nor U13313 (N_13313,N_8125,N_5897);
nand U13314 (N_13314,N_5808,N_8137);
or U13315 (N_13315,N_8323,N_5058);
nor U13316 (N_13316,N_5883,N_5226);
nor U13317 (N_13317,N_8700,N_9859);
or U13318 (N_13318,N_5884,N_6033);
or U13319 (N_13319,N_6506,N_9467);
nand U13320 (N_13320,N_9668,N_6080);
nor U13321 (N_13321,N_7225,N_7852);
nand U13322 (N_13322,N_6334,N_6369);
nor U13323 (N_13323,N_5051,N_6431);
nor U13324 (N_13324,N_9459,N_7849);
and U13325 (N_13325,N_9058,N_7421);
nand U13326 (N_13326,N_5815,N_7536);
nor U13327 (N_13327,N_6384,N_8275);
nand U13328 (N_13328,N_5914,N_9407);
nand U13329 (N_13329,N_6823,N_7450);
nor U13330 (N_13330,N_7945,N_6299);
and U13331 (N_13331,N_9726,N_5627);
and U13332 (N_13332,N_5625,N_5328);
nor U13333 (N_13333,N_8599,N_7099);
nor U13334 (N_13334,N_8047,N_6411);
nand U13335 (N_13335,N_9750,N_8489);
or U13336 (N_13336,N_9826,N_6864);
nor U13337 (N_13337,N_5564,N_6805);
or U13338 (N_13338,N_9712,N_5029);
nand U13339 (N_13339,N_7175,N_9229);
nand U13340 (N_13340,N_6347,N_8267);
or U13341 (N_13341,N_8006,N_6227);
nand U13342 (N_13342,N_7118,N_7910);
or U13343 (N_13343,N_9636,N_5687);
nand U13344 (N_13344,N_8612,N_9360);
nand U13345 (N_13345,N_6697,N_7167);
or U13346 (N_13346,N_9821,N_5331);
or U13347 (N_13347,N_7158,N_7532);
or U13348 (N_13348,N_6629,N_7348);
nand U13349 (N_13349,N_5149,N_9980);
or U13350 (N_13350,N_6193,N_8935);
or U13351 (N_13351,N_9819,N_6928);
and U13352 (N_13352,N_8945,N_8154);
and U13353 (N_13353,N_9220,N_9963);
nor U13354 (N_13354,N_7794,N_7719);
nor U13355 (N_13355,N_6512,N_6151);
nor U13356 (N_13356,N_9890,N_8186);
nand U13357 (N_13357,N_6154,N_7001);
and U13358 (N_13358,N_9526,N_7307);
and U13359 (N_13359,N_7251,N_7356);
or U13360 (N_13360,N_5506,N_5422);
and U13361 (N_13361,N_5434,N_7678);
nand U13362 (N_13362,N_5940,N_8574);
nor U13363 (N_13363,N_7271,N_8620);
nor U13364 (N_13364,N_9919,N_7429);
nor U13365 (N_13365,N_7661,N_7204);
or U13366 (N_13366,N_5241,N_9397);
or U13367 (N_13367,N_7386,N_7477);
nor U13368 (N_13368,N_8198,N_6227);
xor U13369 (N_13369,N_5344,N_5880);
and U13370 (N_13370,N_7109,N_7257);
nor U13371 (N_13371,N_5239,N_7556);
nor U13372 (N_13372,N_8734,N_9162);
nand U13373 (N_13373,N_5584,N_5104);
and U13374 (N_13374,N_6899,N_8647);
or U13375 (N_13375,N_5723,N_5842);
and U13376 (N_13376,N_5064,N_9666);
or U13377 (N_13377,N_5025,N_9460);
nand U13378 (N_13378,N_6017,N_7296);
and U13379 (N_13379,N_8182,N_5487);
or U13380 (N_13380,N_8110,N_9785);
or U13381 (N_13381,N_5191,N_9402);
or U13382 (N_13382,N_9679,N_5975);
nor U13383 (N_13383,N_7680,N_8334);
nor U13384 (N_13384,N_7674,N_5529);
or U13385 (N_13385,N_6792,N_9450);
nand U13386 (N_13386,N_5283,N_8667);
nand U13387 (N_13387,N_7098,N_5329);
and U13388 (N_13388,N_9807,N_6448);
nor U13389 (N_13389,N_9933,N_9811);
or U13390 (N_13390,N_9323,N_8742);
nor U13391 (N_13391,N_6826,N_8885);
nor U13392 (N_13392,N_8256,N_5319);
xor U13393 (N_13393,N_9744,N_5966);
or U13394 (N_13394,N_5350,N_8905);
and U13395 (N_13395,N_7477,N_5257);
and U13396 (N_13396,N_8695,N_9157);
nand U13397 (N_13397,N_6374,N_7494);
and U13398 (N_13398,N_8178,N_6385);
or U13399 (N_13399,N_9688,N_5085);
nor U13400 (N_13400,N_6199,N_8198);
or U13401 (N_13401,N_8004,N_8554);
nand U13402 (N_13402,N_9138,N_9525);
nand U13403 (N_13403,N_6686,N_9947);
or U13404 (N_13404,N_8191,N_7674);
and U13405 (N_13405,N_8654,N_7508);
nor U13406 (N_13406,N_5573,N_7518);
or U13407 (N_13407,N_9067,N_8510);
nor U13408 (N_13408,N_6851,N_7889);
nand U13409 (N_13409,N_9041,N_9645);
or U13410 (N_13410,N_8892,N_6215);
nand U13411 (N_13411,N_5666,N_7349);
nor U13412 (N_13412,N_7336,N_8621);
nor U13413 (N_13413,N_8417,N_9192);
nand U13414 (N_13414,N_8982,N_9650);
nand U13415 (N_13415,N_6082,N_7933);
nor U13416 (N_13416,N_8632,N_9739);
or U13417 (N_13417,N_7484,N_8351);
or U13418 (N_13418,N_8189,N_8117);
nor U13419 (N_13419,N_5423,N_9858);
nor U13420 (N_13420,N_8066,N_7877);
nand U13421 (N_13421,N_9150,N_7152);
nor U13422 (N_13422,N_9216,N_8792);
or U13423 (N_13423,N_8792,N_5293);
nand U13424 (N_13424,N_5929,N_9342);
nand U13425 (N_13425,N_6084,N_5302);
nand U13426 (N_13426,N_5663,N_7939);
nand U13427 (N_13427,N_6520,N_9297);
or U13428 (N_13428,N_6093,N_5533);
and U13429 (N_13429,N_5567,N_8151);
nand U13430 (N_13430,N_7590,N_6884);
nand U13431 (N_13431,N_7390,N_9422);
nand U13432 (N_13432,N_9919,N_7737);
or U13433 (N_13433,N_9799,N_9142);
nand U13434 (N_13434,N_8077,N_8480);
nor U13435 (N_13435,N_7133,N_9089);
nor U13436 (N_13436,N_7552,N_6597);
or U13437 (N_13437,N_7662,N_8713);
nand U13438 (N_13438,N_9516,N_9567);
and U13439 (N_13439,N_7930,N_9373);
nor U13440 (N_13440,N_8698,N_5865);
and U13441 (N_13441,N_6202,N_6587);
nor U13442 (N_13442,N_8339,N_7836);
nand U13443 (N_13443,N_8551,N_8550);
nor U13444 (N_13444,N_6005,N_6211);
nand U13445 (N_13445,N_6030,N_6432);
and U13446 (N_13446,N_9246,N_5965);
nand U13447 (N_13447,N_6165,N_5132);
or U13448 (N_13448,N_9040,N_8890);
nand U13449 (N_13449,N_7585,N_8187);
nor U13450 (N_13450,N_9066,N_6955);
or U13451 (N_13451,N_6304,N_9814);
nor U13452 (N_13452,N_6152,N_9685);
and U13453 (N_13453,N_6414,N_6826);
or U13454 (N_13454,N_5248,N_7954);
nand U13455 (N_13455,N_9444,N_9149);
or U13456 (N_13456,N_9558,N_8490);
or U13457 (N_13457,N_5644,N_5453);
nand U13458 (N_13458,N_5447,N_8107);
nor U13459 (N_13459,N_8296,N_9843);
or U13460 (N_13460,N_5729,N_7384);
nand U13461 (N_13461,N_7866,N_8607);
nand U13462 (N_13462,N_7196,N_7670);
or U13463 (N_13463,N_7922,N_8330);
nor U13464 (N_13464,N_5142,N_7310);
and U13465 (N_13465,N_7091,N_5477);
and U13466 (N_13466,N_9806,N_8683);
and U13467 (N_13467,N_9387,N_5081);
nor U13468 (N_13468,N_8323,N_5466);
nor U13469 (N_13469,N_9621,N_8363);
and U13470 (N_13470,N_9211,N_8395);
nand U13471 (N_13471,N_6177,N_8602);
nor U13472 (N_13472,N_8276,N_5542);
and U13473 (N_13473,N_7173,N_9618);
or U13474 (N_13474,N_8442,N_9644);
nand U13475 (N_13475,N_9510,N_5464);
nand U13476 (N_13476,N_8303,N_8982);
or U13477 (N_13477,N_9733,N_8013);
nor U13478 (N_13478,N_6045,N_6587);
nor U13479 (N_13479,N_5623,N_6080);
or U13480 (N_13480,N_9452,N_9647);
or U13481 (N_13481,N_7538,N_9069);
nor U13482 (N_13482,N_7180,N_5427);
nor U13483 (N_13483,N_8210,N_7021);
nor U13484 (N_13484,N_8527,N_7230);
nand U13485 (N_13485,N_9212,N_9640);
and U13486 (N_13486,N_8836,N_9458);
and U13487 (N_13487,N_9867,N_9280);
or U13488 (N_13488,N_8722,N_9675);
nand U13489 (N_13489,N_6615,N_7373);
or U13490 (N_13490,N_6718,N_8359);
or U13491 (N_13491,N_7926,N_5206);
nand U13492 (N_13492,N_7508,N_8877);
nor U13493 (N_13493,N_9686,N_5667);
nor U13494 (N_13494,N_8979,N_5522);
and U13495 (N_13495,N_5002,N_7560);
nor U13496 (N_13496,N_9662,N_5544);
or U13497 (N_13497,N_7271,N_8757);
nand U13498 (N_13498,N_5725,N_6946);
nor U13499 (N_13499,N_6662,N_8394);
nand U13500 (N_13500,N_5696,N_9423);
nor U13501 (N_13501,N_7003,N_6046);
or U13502 (N_13502,N_6678,N_8972);
or U13503 (N_13503,N_5472,N_6019);
or U13504 (N_13504,N_7226,N_6576);
and U13505 (N_13505,N_8260,N_6447);
and U13506 (N_13506,N_9143,N_5421);
nand U13507 (N_13507,N_5166,N_8533);
or U13508 (N_13508,N_6090,N_7115);
nor U13509 (N_13509,N_7210,N_9576);
and U13510 (N_13510,N_8959,N_9093);
and U13511 (N_13511,N_7290,N_5547);
or U13512 (N_13512,N_6815,N_6753);
or U13513 (N_13513,N_6655,N_8178);
nor U13514 (N_13514,N_6663,N_8940);
and U13515 (N_13515,N_7139,N_6027);
nor U13516 (N_13516,N_7401,N_6443);
nor U13517 (N_13517,N_9906,N_9590);
nand U13518 (N_13518,N_7434,N_6720);
and U13519 (N_13519,N_8983,N_6171);
nor U13520 (N_13520,N_7442,N_7116);
nand U13521 (N_13521,N_7549,N_6100);
nand U13522 (N_13522,N_5231,N_6977);
or U13523 (N_13523,N_8415,N_8037);
or U13524 (N_13524,N_8408,N_7843);
nand U13525 (N_13525,N_6208,N_7525);
and U13526 (N_13526,N_8635,N_6558);
nor U13527 (N_13527,N_9958,N_6191);
and U13528 (N_13528,N_9357,N_9080);
nor U13529 (N_13529,N_7719,N_6361);
and U13530 (N_13530,N_5952,N_8115);
nand U13531 (N_13531,N_9473,N_9283);
or U13532 (N_13532,N_6228,N_7905);
nor U13533 (N_13533,N_7758,N_8366);
and U13534 (N_13534,N_6114,N_6533);
nor U13535 (N_13535,N_9808,N_8925);
or U13536 (N_13536,N_8007,N_5842);
nor U13537 (N_13537,N_5693,N_5695);
and U13538 (N_13538,N_5218,N_5469);
and U13539 (N_13539,N_5578,N_8656);
nand U13540 (N_13540,N_9604,N_5553);
nand U13541 (N_13541,N_6414,N_7643);
xor U13542 (N_13542,N_7534,N_7808);
nor U13543 (N_13543,N_6501,N_5301);
nor U13544 (N_13544,N_6854,N_8674);
nor U13545 (N_13545,N_6417,N_9131);
or U13546 (N_13546,N_9888,N_9890);
nand U13547 (N_13547,N_6192,N_9212);
nor U13548 (N_13548,N_5505,N_9127);
nand U13549 (N_13549,N_5589,N_9191);
and U13550 (N_13550,N_6976,N_8983);
or U13551 (N_13551,N_6357,N_8908);
or U13552 (N_13552,N_6595,N_7706);
nand U13553 (N_13553,N_9560,N_8041);
nand U13554 (N_13554,N_8847,N_8112);
nand U13555 (N_13555,N_6260,N_9937);
nand U13556 (N_13556,N_5335,N_8303);
nor U13557 (N_13557,N_7698,N_9793);
and U13558 (N_13558,N_6736,N_6427);
or U13559 (N_13559,N_7602,N_5555);
or U13560 (N_13560,N_6328,N_6726);
or U13561 (N_13561,N_9885,N_7659);
nor U13562 (N_13562,N_8741,N_9074);
and U13563 (N_13563,N_9756,N_9243);
nor U13564 (N_13564,N_5996,N_5722);
nor U13565 (N_13565,N_9292,N_8657);
nor U13566 (N_13566,N_6503,N_6647);
and U13567 (N_13567,N_6814,N_9011);
nor U13568 (N_13568,N_9693,N_6252);
or U13569 (N_13569,N_9254,N_7443);
nand U13570 (N_13570,N_7433,N_6471);
nor U13571 (N_13571,N_8100,N_7992);
nor U13572 (N_13572,N_8525,N_8271);
and U13573 (N_13573,N_5908,N_5077);
nor U13574 (N_13574,N_5748,N_6778);
and U13575 (N_13575,N_9041,N_6159);
nor U13576 (N_13576,N_6109,N_7862);
and U13577 (N_13577,N_6752,N_6155);
nand U13578 (N_13578,N_7585,N_6177);
and U13579 (N_13579,N_7825,N_5042);
nor U13580 (N_13580,N_9863,N_7027);
and U13581 (N_13581,N_5165,N_7517);
nor U13582 (N_13582,N_5984,N_5009);
and U13583 (N_13583,N_8900,N_5568);
nor U13584 (N_13584,N_5505,N_9822);
nand U13585 (N_13585,N_5222,N_7216);
and U13586 (N_13586,N_5082,N_6601);
nor U13587 (N_13587,N_8190,N_8790);
or U13588 (N_13588,N_5251,N_8988);
xor U13589 (N_13589,N_9327,N_9937);
nand U13590 (N_13590,N_5160,N_8199);
and U13591 (N_13591,N_9251,N_5888);
and U13592 (N_13592,N_9843,N_7236);
or U13593 (N_13593,N_5545,N_7500);
or U13594 (N_13594,N_5002,N_9271);
or U13595 (N_13595,N_6675,N_6968);
nor U13596 (N_13596,N_7743,N_6532);
or U13597 (N_13597,N_9192,N_8632);
nand U13598 (N_13598,N_7278,N_9295);
nor U13599 (N_13599,N_5133,N_8920);
nor U13600 (N_13600,N_9593,N_6222);
nor U13601 (N_13601,N_9248,N_5616);
and U13602 (N_13602,N_5660,N_7395);
and U13603 (N_13603,N_6218,N_5035);
nor U13604 (N_13604,N_6908,N_8982);
or U13605 (N_13605,N_9775,N_7749);
or U13606 (N_13606,N_6145,N_9819);
nand U13607 (N_13607,N_7697,N_7623);
and U13608 (N_13608,N_7723,N_9322);
nand U13609 (N_13609,N_9374,N_5386);
and U13610 (N_13610,N_8308,N_7042);
nor U13611 (N_13611,N_5801,N_7869);
nand U13612 (N_13612,N_5625,N_6560);
nand U13613 (N_13613,N_7611,N_9955);
and U13614 (N_13614,N_8828,N_8306);
or U13615 (N_13615,N_6389,N_8560);
or U13616 (N_13616,N_7722,N_8386);
nand U13617 (N_13617,N_6870,N_7585);
and U13618 (N_13618,N_5492,N_8001);
nand U13619 (N_13619,N_7693,N_7248);
nand U13620 (N_13620,N_9305,N_5056);
nand U13621 (N_13621,N_9217,N_8757);
nand U13622 (N_13622,N_6599,N_9135);
and U13623 (N_13623,N_8447,N_9552);
nand U13624 (N_13624,N_9085,N_9453);
nand U13625 (N_13625,N_9559,N_6718);
and U13626 (N_13626,N_6938,N_6927);
nand U13627 (N_13627,N_7484,N_6628);
nand U13628 (N_13628,N_8806,N_7104);
nor U13629 (N_13629,N_7206,N_6441);
nand U13630 (N_13630,N_9422,N_7207);
and U13631 (N_13631,N_5314,N_5144);
and U13632 (N_13632,N_6344,N_9333);
and U13633 (N_13633,N_8152,N_5615);
and U13634 (N_13634,N_8465,N_6916);
or U13635 (N_13635,N_6877,N_9988);
and U13636 (N_13636,N_9868,N_8421);
and U13637 (N_13637,N_5100,N_8751);
and U13638 (N_13638,N_7710,N_9145);
nor U13639 (N_13639,N_9794,N_8856);
and U13640 (N_13640,N_9454,N_9055);
or U13641 (N_13641,N_7233,N_6685);
and U13642 (N_13642,N_8771,N_9420);
and U13643 (N_13643,N_5504,N_7742);
nor U13644 (N_13644,N_8580,N_8393);
and U13645 (N_13645,N_7906,N_8532);
xor U13646 (N_13646,N_7706,N_5571);
nor U13647 (N_13647,N_5238,N_9333);
or U13648 (N_13648,N_8052,N_9954);
nor U13649 (N_13649,N_9556,N_6077);
or U13650 (N_13650,N_5507,N_6241);
nor U13651 (N_13651,N_8531,N_8886);
and U13652 (N_13652,N_5860,N_9669);
nand U13653 (N_13653,N_5111,N_8719);
or U13654 (N_13654,N_6838,N_7529);
nand U13655 (N_13655,N_9067,N_8257);
nor U13656 (N_13656,N_9053,N_8310);
nor U13657 (N_13657,N_5390,N_8316);
or U13658 (N_13658,N_5148,N_7065);
and U13659 (N_13659,N_8293,N_6177);
or U13660 (N_13660,N_6655,N_9443);
nor U13661 (N_13661,N_6695,N_5235);
or U13662 (N_13662,N_5603,N_6621);
nand U13663 (N_13663,N_5369,N_5671);
and U13664 (N_13664,N_7679,N_9893);
and U13665 (N_13665,N_7142,N_6300);
or U13666 (N_13666,N_5559,N_6191);
or U13667 (N_13667,N_5169,N_6085);
or U13668 (N_13668,N_9982,N_6031);
and U13669 (N_13669,N_7190,N_8222);
nand U13670 (N_13670,N_9654,N_8400);
or U13671 (N_13671,N_9893,N_7211);
nand U13672 (N_13672,N_6396,N_6644);
nand U13673 (N_13673,N_9250,N_9689);
or U13674 (N_13674,N_6142,N_7201);
nand U13675 (N_13675,N_8380,N_7974);
nor U13676 (N_13676,N_9362,N_7074);
nand U13677 (N_13677,N_7622,N_8671);
and U13678 (N_13678,N_6348,N_9376);
nor U13679 (N_13679,N_6878,N_8672);
and U13680 (N_13680,N_8346,N_8406);
and U13681 (N_13681,N_6380,N_6482);
nand U13682 (N_13682,N_9348,N_9296);
nor U13683 (N_13683,N_7797,N_8558);
nor U13684 (N_13684,N_5130,N_9014);
nand U13685 (N_13685,N_7711,N_9601);
and U13686 (N_13686,N_7624,N_8717);
or U13687 (N_13687,N_6430,N_8764);
or U13688 (N_13688,N_7237,N_7260);
nor U13689 (N_13689,N_8004,N_8787);
nor U13690 (N_13690,N_6226,N_8763);
and U13691 (N_13691,N_6278,N_5626);
and U13692 (N_13692,N_8274,N_7591);
nor U13693 (N_13693,N_5893,N_5945);
and U13694 (N_13694,N_7520,N_6759);
nor U13695 (N_13695,N_5276,N_6203);
or U13696 (N_13696,N_5450,N_6696);
and U13697 (N_13697,N_7691,N_9315);
or U13698 (N_13698,N_7071,N_9818);
or U13699 (N_13699,N_5988,N_8927);
and U13700 (N_13700,N_6970,N_5839);
or U13701 (N_13701,N_6754,N_9259);
nor U13702 (N_13702,N_8586,N_7060);
nor U13703 (N_13703,N_8891,N_8126);
and U13704 (N_13704,N_8212,N_9478);
nor U13705 (N_13705,N_8586,N_5281);
and U13706 (N_13706,N_9343,N_5662);
nand U13707 (N_13707,N_9356,N_7988);
nand U13708 (N_13708,N_8135,N_5287);
and U13709 (N_13709,N_7951,N_8696);
and U13710 (N_13710,N_7817,N_9151);
and U13711 (N_13711,N_5742,N_6254);
nor U13712 (N_13712,N_5552,N_6632);
nor U13713 (N_13713,N_5851,N_5874);
nand U13714 (N_13714,N_5255,N_8485);
or U13715 (N_13715,N_5589,N_8148);
nor U13716 (N_13716,N_6012,N_7598);
and U13717 (N_13717,N_5976,N_7491);
and U13718 (N_13718,N_8423,N_7262);
or U13719 (N_13719,N_8787,N_6876);
nand U13720 (N_13720,N_5454,N_8522);
and U13721 (N_13721,N_5585,N_6996);
nand U13722 (N_13722,N_9696,N_9869);
nand U13723 (N_13723,N_7094,N_8124);
and U13724 (N_13724,N_6398,N_6818);
or U13725 (N_13725,N_5464,N_5948);
nor U13726 (N_13726,N_7854,N_9143);
nand U13727 (N_13727,N_6950,N_6070);
and U13728 (N_13728,N_5256,N_5716);
and U13729 (N_13729,N_7106,N_9760);
and U13730 (N_13730,N_9634,N_9653);
and U13731 (N_13731,N_7017,N_5424);
or U13732 (N_13732,N_9334,N_9900);
or U13733 (N_13733,N_7954,N_6878);
nor U13734 (N_13734,N_8786,N_7171);
and U13735 (N_13735,N_9817,N_8426);
xnor U13736 (N_13736,N_8574,N_8095);
nor U13737 (N_13737,N_8290,N_9108);
or U13738 (N_13738,N_8542,N_5849);
and U13739 (N_13739,N_9292,N_8588);
and U13740 (N_13740,N_5943,N_5171);
nand U13741 (N_13741,N_8272,N_6306);
or U13742 (N_13742,N_9710,N_9264);
nand U13743 (N_13743,N_6286,N_5518);
nand U13744 (N_13744,N_7111,N_6942);
nor U13745 (N_13745,N_7911,N_5075);
or U13746 (N_13746,N_9263,N_5070);
and U13747 (N_13747,N_9125,N_5814);
or U13748 (N_13748,N_8936,N_8809);
and U13749 (N_13749,N_5076,N_9943);
and U13750 (N_13750,N_5444,N_6577);
and U13751 (N_13751,N_8513,N_5575);
nand U13752 (N_13752,N_9162,N_6960);
or U13753 (N_13753,N_8956,N_7705);
or U13754 (N_13754,N_8507,N_8794);
nor U13755 (N_13755,N_6061,N_9916);
or U13756 (N_13756,N_9800,N_5439);
or U13757 (N_13757,N_6745,N_9742);
nor U13758 (N_13758,N_8465,N_5890);
nand U13759 (N_13759,N_9011,N_5063);
and U13760 (N_13760,N_8798,N_7809);
nand U13761 (N_13761,N_5839,N_7255);
nor U13762 (N_13762,N_5902,N_5039);
and U13763 (N_13763,N_5143,N_8941);
or U13764 (N_13764,N_7937,N_8556);
nand U13765 (N_13765,N_5620,N_9817);
or U13766 (N_13766,N_7052,N_9423);
nand U13767 (N_13767,N_6658,N_5104);
or U13768 (N_13768,N_5400,N_7400);
and U13769 (N_13769,N_7120,N_8035);
or U13770 (N_13770,N_9210,N_7874);
or U13771 (N_13771,N_8894,N_5742);
or U13772 (N_13772,N_6720,N_5432);
or U13773 (N_13773,N_5674,N_7594);
nand U13774 (N_13774,N_7822,N_8757);
nor U13775 (N_13775,N_8320,N_8588);
and U13776 (N_13776,N_8653,N_7984);
and U13777 (N_13777,N_9131,N_7855);
nor U13778 (N_13778,N_9082,N_7462);
nand U13779 (N_13779,N_7165,N_9174);
nand U13780 (N_13780,N_8560,N_8462);
nand U13781 (N_13781,N_8562,N_7258);
nand U13782 (N_13782,N_8624,N_7359);
and U13783 (N_13783,N_9240,N_7659);
nor U13784 (N_13784,N_7997,N_9741);
or U13785 (N_13785,N_5265,N_9219);
nor U13786 (N_13786,N_5877,N_7506);
nor U13787 (N_13787,N_5031,N_6080);
or U13788 (N_13788,N_5488,N_6530);
and U13789 (N_13789,N_8388,N_9846);
and U13790 (N_13790,N_6919,N_6307);
or U13791 (N_13791,N_7439,N_7242);
and U13792 (N_13792,N_9297,N_7642);
and U13793 (N_13793,N_5894,N_5594);
or U13794 (N_13794,N_5886,N_5616);
and U13795 (N_13795,N_8949,N_7779);
nor U13796 (N_13796,N_8435,N_9332);
and U13797 (N_13797,N_8688,N_6776);
nor U13798 (N_13798,N_6805,N_9873);
nor U13799 (N_13799,N_8140,N_9499);
and U13800 (N_13800,N_9819,N_6985);
nor U13801 (N_13801,N_7365,N_5415);
nand U13802 (N_13802,N_6161,N_7612);
nand U13803 (N_13803,N_5168,N_5750);
or U13804 (N_13804,N_5331,N_7327);
nand U13805 (N_13805,N_7823,N_7069);
or U13806 (N_13806,N_9589,N_5610);
nor U13807 (N_13807,N_6067,N_7446);
and U13808 (N_13808,N_8053,N_8944);
or U13809 (N_13809,N_5740,N_7514);
and U13810 (N_13810,N_6490,N_8044);
nand U13811 (N_13811,N_9430,N_9206);
and U13812 (N_13812,N_8326,N_8546);
or U13813 (N_13813,N_5009,N_9270);
and U13814 (N_13814,N_6728,N_7164);
and U13815 (N_13815,N_7946,N_9583);
or U13816 (N_13816,N_5897,N_6420);
nand U13817 (N_13817,N_6984,N_8470);
or U13818 (N_13818,N_7585,N_5723);
and U13819 (N_13819,N_5660,N_9672);
nor U13820 (N_13820,N_7254,N_9528);
and U13821 (N_13821,N_6156,N_8872);
nor U13822 (N_13822,N_5615,N_6981);
or U13823 (N_13823,N_7068,N_9480);
nand U13824 (N_13824,N_7534,N_5590);
nand U13825 (N_13825,N_5063,N_5500);
or U13826 (N_13826,N_8367,N_9368);
or U13827 (N_13827,N_8114,N_5251);
nand U13828 (N_13828,N_6094,N_6862);
or U13829 (N_13829,N_7419,N_5338);
nand U13830 (N_13830,N_6656,N_5665);
nand U13831 (N_13831,N_5970,N_8952);
nand U13832 (N_13832,N_9514,N_7750);
nor U13833 (N_13833,N_8317,N_6363);
nor U13834 (N_13834,N_6514,N_5362);
or U13835 (N_13835,N_5911,N_7855);
or U13836 (N_13836,N_6691,N_7151);
nor U13837 (N_13837,N_8737,N_8024);
or U13838 (N_13838,N_7352,N_5983);
nor U13839 (N_13839,N_5787,N_6159);
nor U13840 (N_13840,N_9010,N_5925);
or U13841 (N_13841,N_5705,N_6482);
nor U13842 (N_13842,N_7725,N_9568);
nand U13843 (N_13843,N_6796,N_7386);
or U13844 (N_13844,N_8485,N_5714);
or U13845 (N_13845,N_5193,N_6395);
nor U13846 (N_13846,N_8052,N_8199);
nand U13847 (N_13847,N_8004,N_8988);
nor U13848 (N_13848,N_8050,N_6496);
or U13849 (N_13849,N_7456,N_5570);
nand U13850 (N_13850,N_6559,N_8947);
nor U13851 (N_13851,N_7809,N_5185);
or U13852 (N_13852,N_9286,N_9851);
nor U13853 (N_13853,N_6612,N_8096);
or U13854 (N_13854,N_9058,N_6776);
nand U13855 (N_13855,N_8434,N_5887);
nor U13856 (N_13856,N_6085,N_7188);
nor U13857 (N_13857,N_8192,N_5634);
and U13858 (N_13858,N_7047,N_9666);
and U13859 (N_13859,N_6131,N_6569);
and U13860 (N_13860,N_9011,N_5130);
or U13861 (N_13861,N_7157,N_5104);
nor U13862 (N_13862,N_7728,N_9347);
nand U13863 (N_13863,N_8000,N_8759);
nor U13864 (N_13864,N_5824,N_5274);
nor U13865 (N_13865,N_5952,N_9364);
or U13866 (N_13866,N_7056,N_9623);
or U13867 (N_13867,N_9970,N_6295);
xnor U13868 (N_13868,N_7083,N_6972);
or U13869 (N_13869,N_6754,N_9409);
xor U13870 (N_13870,N_9796,N_7795);
or U13871 (N_13871,N_8466,N_5662);
nand U13872 (N_13872,N_7242,N_5257);
nand U13873 (N_13873,N_5353,N_6297);
nor U13874 (N_13874,N_9402,N_9683);
nor U13875 (N_13875,N_8009,N_9831);
or U13876 (N_13876,N_7640,N_5126);
and U13877 (N_13877,N_5091,N_6254);
and U13878 (N_13878,N_6927,N_9918);
and U13879 (N_13879,N_6596,N_8871);
nand U13880 (N_13880,N_6180,N_7147);
nor U13881 (N_13881,N_5377,N_7369);
or U13882 (N_13882,N_5031,N_6878);
and U13883 (N_13883,N_6981,N_9843);
or U13884 (N_13884,N_6974,N_5850);
nor U13885 (N_13885,N_5727,N_7197);
or U13886 (N_13886,N_5952,N_7060);
and U13887 (N_13887,N_9797,N_6992);
nor U13888 (N_13888,N_8290,N_6297);
nor U13889 (N_13889,N_9613,N_7244);
or U13890 (N_13890,N_9495,N_5231);
or U13891 (N_13891,N_5364,N_9250);
nor U13892 (N_13892,N_8439,N_8494);
nor U13893 (N_13893,N_9812,N_9276);
nand U13894 (N_13894,N_6999,N_8779);
or U13895 (N_13895,N_5196,N_5423);
or U13896 (N_13896,N_6709,N_9683);
and U13897 (N_13897,N_8377,N_7757);
or U13898 (N_13898,N_7649,N_7713);
or U13899 (N_13899,N_9597,N_8330);
nor U13900 (N_13900,N_9073,N_7370);
and U13901 (N_13901,N_5283,N_9161);
nand U13902 (N_13902,N_9039,N_6214);
nand U13903 (N_13903,N_8078,N_9858);
or U13904 (N_13904,N_6865,N_5317);
nand U13905 (N_13905,N_6986,N_5174);
nor U13906 (N_13906,N_9240,N_9851);
nand U13907 (N_13907,N_8744,N_5804);
or U13908 (N_13908,N_6681,N_5490);
nand U13909 (N_13909,N_6729,N_9827);
nor U13910 (N_13910,N_6392,N_9345);
nor U13911 (N_13911,N_6661,N_7284);
and U13912 (N_13912,N_8375,N_5972);
or U13913 (N_13913,N_5636,N_6973);
nand U13914 (N_13914,N_7769,N_7452);
or U13915 (N_13915,N_9625,N_6620);
nor U13916 (N_13916,N_5177,N_7615);
nand U13917 (N_13917,N_8892,N_9610);
or U13918 (N_13918,N_5431,N_7050);
or U13919 (N_13919,N_6941,N_5809);
nand U13920 (N_13920,N_8478,N_6575);
nor U13921 (N_13921,N_6032,N_9167);
nor U13922 (N_13922,N_7114,N_9331);
and U13923 (N_13923,N_6113,N_8957);
nand U13924 (N_13924,N_7196,N_9622);
nand U13925 (N_13925,N_7356,N_9287);
and U13926 (N_13926,N_6898,N_9258);
and U13927 (N_13927,N_8567,N_5080);
nor U13928 (N_13928,N_7078,N_6792);
or U13929 (N_13929,N_9387,N_5457);
nor U13930 (N_13930,N_7207,N_6167);
and U13931 (N_13931,N_6997,N_6744);
nor U13932 (N_13932,N_7295,N_8376);
and U13933 (N_13933,N_5100,N_5380);
and U13934 (N_13934,N_5955,N_7476);
nand U13935 (N_13935,N_6361,N_6700);
nand U13936 (N_13936,N_6507,N_5379);
nor U13937 (N_13937,N_6810,N_9565);
and U13938 (N_13938,N_6401,N_9566);
nand U13939 (N_13939,N_9725,N_6017);
nand U13940 (N_13940,N_5733,N_5780);
and U13941 (N_13941,N_6301,N_7035);
nand U13942 (N_13942,N_5394,N_9669);
nor U13943 (N_13943,N_6825,N_7704);
nand U13944 (N_13944,N_5210,N_7768);
nor U13945 (N_13945,N_6917,N_8621);
and U13946 (N_13946,N_5537,N_9961);
or U13947 (N_13947,N_6140,N_9093);
and U13948 (N_13948,N_5187,N_7706);
nand U13949 (N_13949,N_5159,N_8425);
or U13950 (N_13950,N_5751,N_9111);
nand U13951 (N_13951,N_9344,N_7089);
and U13952 (N_13952,N_9503,N_9522);
nor U13953 (N_13953,N_8242,N_6634);
and U13954 (N_13954,N_9307,N_8350);
and U13955 (N_13955,N_5486,N_9374);
nor U13956 (N_13956,N_5263,N_5562);
and U13957 (N_13957,N_8851,N_7209);
nand U13958 (N_13958,N_7687,N_8983);
or U13959 (N_13959,N_8808,N_7473);
nor U13960 (N_13960,N_6125,N_5555);
and U13961 (N_13961,N_6945,N_8146);
and U13962 (N_13962,N_8582,N_9540);
nor U13963 (N_13963,N_5779,N_6531);
or U13964 (N_13964,N_7134,N_7187);
nand U13965 (N_13965,N_6312,N_8009);
and U13966 (N_13966,N_6809,N_7754);
nor U13967 (N_13967,N_7988,N_9413);
nand U13968 (N_13968,N_8625,N_5558);
nand U13969 (N_13969,N_8060,N_9157);
xor U13970 (N_13970,N_7299,N_8941);
nand U13971 (N_13971,N_5568,N_5407);
and U13972 (N_13972,N_5986,N_6266);
nor U13973 (N_13973,N_8963,N_9750);
nand U13974 (N_13974,N_5830,N_5071);
nor U13975 (N_13975,N_5619,N_5342);
nor U13976 (N_13976,N_5237,N_5676);
nand U13977 (N_13977,N_9026,N_8848);
or U13978 (N_13978,N_6777,N_8346);
and U13979 (N_13979,N_7803,N_9744);
nor U13980 (N_13980,N_5942,N_6788);
nor U13981 (N_13981,N_8307,N_5893);
and U13982 (N_13982,N_9138,N_9539);
and U13983 (N_13983,N_5663,N_6024);
or U13984 (N_13984,N_6056,N_5113);
and U13985 (N_13985,N_8738,N_9498);
nor U13986 (N_13986,N_7867,N_9232);
nor U13987 (N_13987,N_9657,N_5325);
or U13988 (N_13988,N_9092,N_7044);
and U13989 (N_13989,N_8587,N_9181);
or U13990 (N_13990,N_9349,N_5748);
nand U13991 (N_13991,N_9971,N_7499);
xnor U13992 (N_13992,N_6265,N_8467);
or U13993 (N_13993,N_5390,N_5617);
nand U13994 (N_13994,N_8652,N_5952);
nand U13995 (N_13995,N_9765,N_7008);
nor U13996 (N_13996,N_5170,N_5742);
nand U13997 (N_13997,N_7542,N_9801);
or U13998 (N_13998,N_6057,N_5344);
nor U13999 (N_13999,N_8642,N_5943);
nor U14000 (N_14000,N_7914,N_7040);
nor U14001 (N_14001,N_5887,N_9228);
nor U14002 (N_14002,N_7634,N_5977);
or U14003 (N_14003,N_6820,N_7996);
nand U14004 (N_14004,N_7249,N_6884);
and U14005 (N_14005,N_6970,N_7557);
nand U14006 (N_14006,N_5108,N_5935);
nor U14007 (N_14007,N_7284,N_7610);
and U14008 (N_14008,N_8744,N_5135);
nor U14009 (N_14009,N_7350,N_6671);
or U14010 (N_14010,N_9903,N_8106);
or U14011 (N_14011,N_8270,N_8696);
nand U14012 (N_14012,N_7066,N_7318);
nand U14013 (N_14013,N_5622,N_8639);
or U14014 (N_14014,N_9366,N_7753);
and U14015 (N_14015,N_6945,N_7838);
nor U14016 (N_14016,N_6264,N_6392);
or U14017 (N_14017,N_7235,N_5300);
nand U14018 (N_14018,N_7182,N_8640);
nor U14019 (N_14019,N_5540,N_5766);
and U14020 (N_14020,N_6821,N_5674);
nor U14021 (N_14021,N_8592,N_7594);
and U14022 (N_14022,N_5362,N_7758);
nand U14023 (N_14023,N_9596,N_6501);
nor U14024 (N_14024,N_6833,N_6152);
and U14025 (N_14025,N_8852,N_9463);
nand U14026 (N_14026,N_9694,N_5650);
nand U14027 (N_14027,N_6124,N_8883);
and U14028 (N_14028,N_6061,N_7602);
and U14029 (N_14029,N_7207,N_8655);
and U14030 (N_14030,N_8293,N_8433);
or U14031 (N_14031,N_7164,N_7046);
nand U14032 (N_14032,N_5767,N_7007);
nor U14033 (N_14033,N_6644,N_7639);
nor U14034 (N_14034,N_6177,N_8627);
xor U14035 (N_14035,N_7016,N_9882);
or U14036 (N_14036,N_6152,N_6835);
and U14037 (N_14037,N_8543,N_5921);
nand U14038 (N_14038,N_8370,N_5649);
or U14039 (N_14039,N_5198,N_5606);
nand U14040 (N_14040,N_7545,N_6974);
nor U14041 (N_14041,N_6659,N_6834);
or U14042 (N_14042,N_9492,N_5367);
nor U14043 (N_14043,N_9445,N_7651);
or U14044 (N_14044,N_8307,N_5373);
nor U14045 (N_14045,N_7795,N_8563);
nor U14046 (N_14046,N_7557,N_5899);
nand U14047 (N_14047,N_9837,N_6088);
nand U14048 (N_14048,N_5167,N_7190);
nand U14049 (N_14049,N_7630,N_7918);
nor U14050 (N_14050,N_8015,N_8452);
nor U14051 (N_14051,N_6130,N_7072);
and U14052 (N_14052,N_6755,N_8012);
or U14053 (N_14053,N_6407,N_7572);
and U14054 (N_14054,N_9317,N_6321);
nor U14055 (N_14055,N_7817,N_8688);
nor U14056 (N_14056,N_7120,N_6568);
nand U14057 (N_14057,N_9957,N_8416);
nand U14058 (N_14058,N_6204,N_7723);
nand U14059 (N_14059,N_5228,N_8456);
or U14060 (N_14060,N_9346,N_8362);
nor U14061 (N_14061,N_6185,N_6325);
nand U14062 (N_14062,N_9525,N_5968);
nand U14063 (N_14063,N_5085,N_9908);
and U14064 (N_14064,N_7987,N_5595);
nor U14065 (N_14065,N_6010,N_7684);
nand U14066 (N_14066,N_8663,N_5750);
or U14067 (N_14067,N_5656,N_7558);
and U14068 (N_14068,N_6254,N_6586);
nor U14069 (N_14069,N_9816,N_5389);
nor U14070 (N_14070,N_9301,N_9450);
and U14071 (N_14071,N_5080,N_9453);
nand U14072 (N_14072,N_9944,N_5119);
or U14073 (N_14073,N_7530,N_8800);
or U14074 (N_14074,N_9115,N_5997);
or U14075 (N_14075,N_5120,N_8009);
or U14076 (N_14076,N_9236,N_8725);
or U14077 (N_14077,N_6628,N_7029);
and U14078 (N_14078,N_8131,N_7591);
nand U14079 (N_14079,N_9485,N_9398);
or U14080 (N_14080,N_8922,N_5810);
nor U14081 (N_14081,N_9919,N_6753);
nor U14082 (N_14082,N_7925,N_9940);
nand U14083 (N_14083,N_5189,N_6516);
xor U14084 (N_14084,N_6299,N_6991);
nor U14085 (N_14085,N_9059,N_7170);
and U14086 (N_14086,N_7390,N_9762);
and U14087 (N_14087,N_9383,N_9599);
or U14088 (N_14088,N_8339,N_5597);
nand U14089 (N_14089,N_6906,N_9231);
nor U14090 (N_14090,N_8403,N_8681);
nor U14091 (N_14091,N_6973,N_6341);
nand U14092 (N_14092,N_7038,N_8250);
or U14093 (N_14093,N_6756,N_6677);
or U14094 (N_14094,N_8385,N_7116);
or U14095 (N_14095,N_6728,N_5639);
nor U14096 (N_14096,N_5057,N_7574);
or U14097 (N_14097,N_6615,N_5349);
or U14098 (N_14098,N_7098,N_8158);
nor U14099 (N_14099,N_9817,N_7901);
and U14100 (N_14100,N_7911,N_8830);
nor U14101 (N_14101,N_5018,N_6826);
and U14102 (N_14102,N_9198,N_6063);
and U14103 (N_14103,N_5706,N_7867);
nand U14104 (N_14104,N_6688,N_6628);
and U14105 (N_14105,N_7955,N_8091);
and U14106 (N_14106,N_8596,N_7694);
or U14107 (N_14107,N_9390,N_8849);
or U14108 (N_14108,N_8225,N_8678);
and U14109 (N_14109,N_6824,N_8293);
nand U14110 (N_14110,N_7377,N_8190);
and U14111 (N_14111,N_5752,N_9689);
or U14112 (N_14112,N_8662,N_5550);
or U14113 (N_14113,N_7306,N_7767);
nand U14114 (N_14114,N_6152,N_7907);
nand U14115 (N_14115,N_9938,N_6720);
or U14116 (N_14116,N_8343,N_9020);
and U14117 (N_14117,N_9618,N_8381);
nand U14118 (N_14118,N_9491,N_9553);
nor U14119 (N_14119,N_9599,N_8616);
or U14120 (N_14120,N_8361,N_9770);
or U14121 (N_14121,N_5459,N_6412);
and U14122 (N_14122,N_6185,N_6949);
nor U14123 (N_14123,N_6021,N_5262);
or U14124 (N_14124,N_6990,N_6507);
and U14125 (N_14125,N_8139,N_7984);
nand U14126 (N_14126,N_9422,N_6117);
and U14127 (N_14127,N_6658,N_8155);
or U14128 (N_14128,N_5160,N_8583);
and U14129 (N_14129,N_7667,N_7948);
nand U14130 (N_14130,N_9971,N_9514);
and U14131 (N_14131,N_5488,N_5773);
or U14132 (N_14132,N_5505,N_7546);
and U14133 (N_14133,N_8903,N_7793);
nand U14134 (N_14134,N_8677,N_7265);
and U14135 (N_14135,N_9091,N_6444);
nand U14136 (N_14136,N_8017,N_8786);
or U14137 (N_14137,N_5390,N_8873);
or U14138 (N_14138,N_7643,N_5509);
nand U14139 (N_14139,N_5754,N_9874);
and U14140 (N_14140,N_8232,N_7753);
and U14141 (N_14141,N_8087,N_7412);
nand U14142 (N_14142,N_9092,N_5389);
or U14143 (N_14143,N_5719,N_9899);
nand U14144 (N_14144,N_8594,N_7182);
or U14145 (N_14145,N_7304,N_5660);
nand U14146 (N_14146,N_7406,N_7197);
nand U14147 (N_14147,N_9003,N_7106);
nand U14148 (N_14148,N_7829,N_7030);
nor U14149 (N_14149,N_7425,N_9991);
or U14150 (N_14150,N_5414,N_9115);
and U14151 (N_14151,N_8757,N_8921);
or U14152 (N_14152,N_8839,N_6484);
or U14153 (N_14153,N_9226,N_7000);
nand U14154 (N_14154,N_9323,N_5344);
or U14155 (N_14155,N_9420,N_7708);
nor U14156 (N_14156,N_6611,N_9484);
or U14157 (N_14157,N_5686,N_8267);
and U14158 (N_14158,N_7257,N_7584);
nand U14159 (N_14159,N_7987,N_9590);
or U14160 (N_14160,N_5308,N_8837);
and U14161 (N_14161,N_8772,N_8756);
xnor U14162 (N_14162,N_6673,N_5647);
nand U14163 (N_14163,N_6534,N_8314);
and U14164 (N_14164,N_6123,N_9178);
or U14165 (N_14165,N_7637,N_6133);
or U14166 (N_14166,N_5311,N_8516);
and U14167 (N_14167,N_8847,N_6156);
nor U14168 (N_14168,N_7325,N_7490);
or U14169 (N_14169,N_8192,N_5890);
nand U14170 (N_14170,N_7151,N_8598);
or U14171 (N_14171,N_6438,N_5053);
nand U14172 (N_14172,N_5776,N_8930);
nor U14173 (N_14173,N_9752,N_5407);
nand U14174 (N_14174,N_6758,N_6321);
nand U14175 (N_14175,N_8767,N_8109);
or U14176 (N_14176,N_9273,N_6484);
nand U14177 (N_14177,N_9481,N_6669);
or U14178 (N_14178,N_7473,N_7133);
nand U14179 (N_14179,N_5102,N_5953);
and U14180 (N_14180,N_5769,N_5136);
and U14181 (N_14181,N_8884,N_8574);
nor U14182 (N_14182,N_5361,N_5945);
or U14183 (N_14183,N_7258,N_8634);
or U14184 (N_14184,N_5542,N_8352);
or U14185 (N_14185,N_9485,N_5625);
and U14186 (N_14186,N_9086,N_7525);
and U14187 (N_14187,N_6110,N_8761);
nand U14188 (N_14188,N_7909,N_7934);
nand U14189 (N_14189,N_9645,N_6316);
or U14190 (N_14190,N_9988,N_6977);
and U14191 (N_14191,N_5624,N_5039);
and U14192 (N_14192,N_6353,N_5103);
nand U14193 (N_14193,N_5936,N_8215);
or U14194 (N_14194,N_6163,N_9687);
or U14195 (N_14195,N_5914,N_9708);
and U14196 (N_14196,N_7039,N_6214);
nor U14197 (N_14197,N_7043,N_8632);
nor U14198 (N_14198,N_9245,N_7277);
and U14199 (N_14199,N_7308,N_5533);
nand U14200 (N_14200,N_5712,N_6521);
or U14201 (N_14201,N_7708,N_5823);
and U14202 (N_14202,N_5352,N_8879);
or U14203 (N_14203,N_8953,N_7405);
nor U14204 (N_14204,N_8522,N_8851);
or U14205 (N_14205,N_9098,N_7042);
and U14206 (N_14206,N_8896,N_5707);
nor U14207 (N_14207,N_7700,N_9763);
nand U14208 (N_14208,N_9961,N_8931);
nand U14209 (N_14209,N_5587,N_7215);
nand U14210 (N_14210,N_7274,N_8186);
nor U14211 (N_14211,N_7960,N_6327);
and U14212 (N_14212,N_6759,N_7785);
nand U14213 (N_14213,N_5963,N_8705);
or U14214 (N_14214,N_8602,N_5925);
or U14215 (N_14215,N_8535,N_8328);
and U14216 (N_14216,N_9440,N_7301);
nor U14217 (N_14217,N_5351,N_7501);
nor U14218 (N_14218,N_9185,N_6853);
nand U14219 (N_14219,N_7391,N_7665);
nand U14220 (N_14220,N_5707,N_9432);
and U14221 (N_14221,N_6246,N_9441);
and U14222 (N_14222,N_9557,N_6748);
and U14223 (N_14223,N_8670,N_8463);
and U14224 (N_14224,N_9876,N_7648);
nand U14225 (N_14225,N_7215,N_9435);
nor U14226 (N_14226,N_9465,N_5313);
or U14227 (N_14227,N_7226,N_6458);
nor U14228 (N_14228,N_8131,N_8195);
and U14229 (N_14229,N_7519,N_8413);
nand U14230 (N_14230,N_8824,N_9135);
or U14231 (N_14231,N_8211,N_9850);
or U14232 (N_14232,N_7402,N_5365);
and U14233 (N_14233,N_5019,N_5791);
and U14234 (N_14234,N_7320,N_6448);
or U14235 (N_14235,N_7421,N_8458);
or U14236 (N_14236,N_5067,N_6230);
nand U14237 (N_14237,N_7797,N_7432);
and U14238 (N_14238,N_9906,N_7571);
and U14239 (N_14239,N_6983,N_6935);
and U14240 (N_14240,N_6733,N_6924);
nor U14241 (N_14241,N_8451,N_8768);
nor U14242 (N_14242,N_8739,N_6865);
or U14243 (N_14243,N_9818,N_6244);
nor U14244 (N_14244,N_5876,N_5134);
or U14245 (N_14245,N_8660,N_6211);
nand U14246 (N_14246,N_5486,N_6613);
nand U14247 (N_14247,N_6758,N_6231);
nor U14248 (N_14248,N_6073,N_5851);
and U14249 (N_14249,N_8495,N_8940);
or U14250 (N_14250,N_6123,N_5213);
nor U14251 (N_14251,N_5330,N_8011);
nand U14252 (N_14252,N_5567,N_6395);
or U14253 (N_14253,N_9858,N_9848);
nand U14254 (N_14254,N_5936,N_9538);
nand U14255 (N_14255,N_5830,N_6893);
nor U14256 (N_14256,N_8030,N_8856);
or U14257 (N_14257,N_8465,N_7916);
nand U14258 (N_14258,N_9508,N_7704);
nor U14259 (N_14259,N_6341,N_6911);
nand U14260 (N_14260,N_9015,N_5639);
or U14261 (N_14261,N_5926,N_6244);
or U14262 (N_14262,N_9332,N_6942);
or U14263 (N_14263,N_5915,N_9383);
nor U14264 (N_14264,N_5776,N_5571);
nand U14265 (N_14265,N_9094,N_9386);
nand U14266 (N_14266,N_6325,N_9213);
or U14267 (N_14267,N_6279,N_7706);
or U14268 (N_14268,N_8105,N_5036);
nor U14269 (N_14269,N_9778,N_7251);
nand U14270 (N_14270,N_6665,N_6115);
or U14271 (N_14271,N_7754,N_9852);
and U14272 (N_14272,N_8725,N_8084);
nand U14273 (N_14273,N_9429,N_5182);
and U14274 (N_14274,N_5364,N_5663);
nand U14275 (N_14275,N_5644,N_9888);
nand U14276 (N_14276,N_7232,N_7736);
nand U14277 (N_14277,N_5670,N_9188);
nor U14278 (N_14278,N_5569,N_6607);
or U14279 (N_14279,N_5750,N_6364);
nand U14280 (N_14280,N_9047,N_9199);
or U14281 (N_14281,N_7622,N_5366);
nand U14282 (N_14282,N_7204,N_8930);
and U14283 (N_14283,N_6755,N_9524);
or U14284 (N_14284,N_8640,N_7090);
nor U14285 (N_14285,N_5672,N_9290);
nand U14286 (N_14286,N_8874,N_5828);
or U14287 (N_14287,N_7609,N_9081);
and U14288 (N_14288,N_9963,N_6142);
or U14289 (N_14289,N_9940,N_5321);
and U14290 (N_14290,N_9056,N_8709);
nand U14291 (N_14291,N_8419,N_7884);
or U14292 (N_14292,N_5220,N_6187);
nor U14293 (N_14293,N_7612,N_8808);
or U14294 (N_14294,N_6267,N_5330);
or U14295 (N_14295,N_9474,N_7352);
nor U14296 (N_14296,N_7165,N_9696);
and U14297 (N_14297,N_8423,N_8282);
or U14298 (N_14298,N_7146,N_8512);
xor U14299 (N_14299,N_7418,N_8118);
and U14300 (N_14300,N_8142,N_5919);
and U14301 (N_14301,N_9814,N_6012);
nand U14302 (N_14302,N_5568,N_9563);
nor U14303 (N_14303,N_7452,N_9680);
nor U14304 (N_14304,N_9384,N_6943);
or U14305 (N_14305,N_8444,N_9823);
nor U14306 (N_14306,N_6455,N_9714);
nand U14307 (N_14307,N_7242,N_9392);
or U14308 (N_14308,N_6162,N_8089);
and U14309 (N_14309,N_7907,N_6972);
nor U14310 (N_14310,N_6470,N_7924);
and U14311 (N_14311,N_9795,N_9804);
nor U14312 (N_14312,N_6742,N_9928);
or U14313 (N_14313,N_6011,N_7843);
and U14314 (N_14314,N_9820,N_5980);
and U14315 (N_14315,N_5358,N_8580);
and U14316 (N_14316,N_7984,N_9611);
and U14317 (N_14317,N_7111,N_9762);
xor U14318 (N_14318,N_9243,N_9758);
or U14319 (N_14319,N_5204,N_5634);
or U14320 (N_14320,N_9487,N_7446);
and U14321 (N_14321,N_8242,N_9012);
xor U14322 (N_14322,N_5589,N_6293);
nor U14323 (N_14323,N_6878,N_5991);
and U14324 (N_14324,N_7159,N_8559);
nand U14325 (N_14325,N_9686,N_9579);
or U14326 (N_14326,N_5682,N_6301);
and U14327 (N_14327,N_8720,N_5490);
nand U14328 (N_14328,N_9615,N_8669);
or U14329 (N_14329,N_6398,N_6537);
or U14330 (N_14330,N_8797,N_7785);
and U14331 (N_14331,N_7957,N_7051);
nor U14332 (N_14332,N_9266,N_7388);
nand U14333 (N_14333,N_9994,N_9166);
nor U14334 (N_14334,N_7282,N_5111);
nand U14335 (N_14335,N_7038,N_8753);
nand U14336 (N_14336,N_6191,N_8566);
nor U14337 (N_14337,N_7238,N_7688);
or U14338 (N_14338,N_6648,N_5901);
or U14339 (N_14339,N_8780,N_5561);
xor U14340 (N_14340,N_9402,N_5414);
nand U14341 (N_14341,N_5319,N_6577);
nand U14342 (N_14342,N_5983,N_7867);
nor U14343 (N_14343,N_7099,N_9061);
nor U14344 (N_14344,N_8314,N_6855);
and U14345 (N_14345,N_8342,N_9872);
nor U14346 (N_14346,N_7755,N_7005);
nand U14347 (N_14347,N_9775,N_6165);
and U14348 (N_14348,N_5661,N_9936);
nand U14349 (N_14349,N_6823,N_7361);
nand U14350 (N_14350,N_8498,N_5829);
or U14351 (N_14351,N_8089,N_9813);
and U14352 (N_14352,N_7934,N_7066);
or U14353 (N_14353,N_7560,N_6465);
or U14354 (N_14354,N_5049,N_6213);
nor U14355 (N_14355,N_9556,N_8944);
or U14356 (N_14356,N_5564,N_9262);
or U14357 (N_14357,N_8404,N_6303);
and U14358 (N_14358,N_5436,N_7709);
or U14359 (N_14359,N_6477,N_8353);
and U14360 (N_14360,N_6079,N_7681);
or U14361 (N_14361,N_7693,N_6032);
or U14362 (N_14362,N_6450,N_8698);
and U14363 (N_14363,N_6167,N_7584);
nor U14364 (N_14364,N_8846,N_9170);
or U14365 (N_14365,N_5689,N_7206);
nor U14366 (N_14366,N_8565,N_5562);
nor U14367 (N_14367,N_9197,N_7322);
and U14368 (N_14368,N_8530,N_8622);
nor U14369 (N_14369,N_7528,N_8279);
and U14370 (N_14370,N_9068,N_5727);
nor U14371 (N_14371,N_6409,N_5650);
or U14372 (N_14372,N_8350,N_8487);
nand U14373 (N_14373,N_5822,N_8315);
nand U14374 (N_14374,N_8539,N_9613);
and U14375 (N_14375,N_8192,N_6247);
and U14376 (N_14376,N_7668,N_9882);
nor U14377 (N_14377,N_9781,N_5102);
nand U14378 (N_14378,N_9054,N_5393);
or U14379 (N_14379,N_8394,N_7807);
and U14380 (N_14380,N_8189,N_8144);
or U14381 (N_14381,N_6246,N_5939);
nor U14382 (N_14382,N_9964,N_5553);
nor U14383 (N_14383,N_6223,N_9964);
nor U14384 (N_14384,N_7842,N_6143);
and U14385 (N_14385,N_5049,N_7166);
nor U14386 (N_14386,N_5623,N_7487);
nand U14387 (N_14387,N_8062,N_7576);
or U14388 (N_14388,N_9709,N_6870);
and U14389 (N_14389,N_5804,N_7379);
nor U14390 (N_14390,N_9257,N_6585);
or U14391 (N_14391,N_7123,N_9493);
nand U14392 (N_14392,N_6913,N_6258);
nand U14393 (N_14393,N_8081,N_5580);
or U14394 (N_14394,N_6962,N_9877);
or U14395 (N_14395,N_8629,N_8901);
or U14396 (N_14396,N_7769,N_6468);
nand U14397 (N_14397,N_8982,N_8169);
nor U14398 (N_14398,N_9832,N_5382);
and U14399 (N_14399,N_9414,N_8863);
and U14400 (N_14400,N_9758,N_9845);
nor U14401 (N_14401,N_7648,N_5391);
and U14402 (N_14402,N_8173,N_6512);
and U14403 (N_14403,N_8108,N_8619);
and U14404 (N_14404,N_6166,N_8149);
or U14405 (N_14405,N_7906,N_8517);
or U14406 (N_14406,N_6343,N_5541);
nand U14407 (N_14407,N_8783,N_5350);
and U14408 (N_14408,N_5563,N_6010);
or U14409 (N_14409,N_6709,N_9959);
nor U14410 (N_14410,N_5526,N_9867);
nor U14411 (N_14411,N_6447,N_5698);
nand U14412 (N_14412,N_5249,N_7841);
and U14413 (N_14413,N_7225,N_6987);
nor U14414 (N_14414,N_8395,N_8186);
and U14415 (N_14415,N_6865,N_5686);
nand U14416 (N_14416,N_5906,N_7758);
or U14417 (N_14417,N_7141,N_5559);
nor U14418 (N_14418,N_9567,N_6245);
nand U14419 (N_14419,N_7768,N_8770);
nor U14420 (N_14420,N_6854,N_9636);
and U14421 (N_14421,N_7240,N_6427);
nand U14422 (N_14422,N_6860,N_9652);
and U14423 (N_14423,N_5726,N_7497);
or U14424 (N_14424,N_6485,N_6135);
nor U14425 (N_14425,N_5982,N_9582);
or U14426 (N_14426,N_9744,N_5050);
nand U14427 (N_14427,N_8168,N_8323);
nand U14428 (N_14428,N_6949,N_9334);
or U14429 (N_14429,N_8172,N_5224);
nor U14430 (N_14430,N_7707,N_5234);
or U14431 (N_14431,N_6336,N_6276);
or U14432 (N_14432,N_8413,N_6815);
nand U14433 (N_14433,N_9743,N_5999);
or U14434 (N_14434,N_9008,N_5152);
and U14435 (N_14435,N_8154,N_8786);
and U14436 (N_14436,N_8241,N_5512);
nor U14437 (N_14437,N_6086,N_8353);
nor U14438 (N_14438,N_9938,N_9148);
or U14439 (N_14439,N_5930,N_5943);
nand U14440 (N_14440,N_9975,N_7566);
and U14441 (N_14441,N_9552,N_7310);
nor U14442 (N_14442,N_5772,N_9536);
nand U14443 (N_14443,N_7364,N_7869);
or U14444 (N_14444,N_7578,N_7592);
nand U14445 (N_14445,N_9785,N_7574);
nand U14446 (N_14446,N_6464,N_8147);
nand U14447 (N_14447,N_7277,N_9747);
and U14448 (N_14448,N_5653,N_9082);
and U14449 (N_14449,N_5871,N_9242);
nor U14450 (N_14450,N_9469,N_8901);
nor U14451 (N_14451,N_6220,N_7739);
nand U14452 (N_14452,N_6111,N_7178);
nand U14453 (N_14453,N_9132,N_5433);
nor U14454 (N_14454,N_7607,N_7204);
or U14455 (N_14455,N_9806,N_8896);
nor U14456 (N_14456,N_9912,N_7475);
nor U14457 (N_14457,N_5355,N_8873);
and U14458 (N_14458,N_8561,N_7837);
or U14459 (N_14459,N_6073,N_9667);
or U14460 (N_14460,N_7159,N_7368);
nor U14461 (N_14461,N_7839,N_7112);
or U14462 (N_14462,N_8345,N_8420);
or U14463 (N_14463,N_6822,N_8849);
nand U14464 (N_14464,N_9404,N_8697);
and U14465 (N_14465,N_9203,N_6619);
and U14466 (N_14466,N_9366,N_7760);
nand U14467 (N_14467,N_6085,N_9151);
and U14468 (N_14468,N_6751,N_6333);
nand U14469 (N_14469,N_6077,N_7672);
or U14470 (N_14470,N_9471,N_6332);
nand U14471 (N_14471,N_9925,N_6376);
nand U14472 (N_14472,N_9674,N_5023);
nand U14473 (N_14473,N_8352,N_8700);
and U14474 (N_14474,N_9519,N_9946);
and U14475 (N_14475,N_5064,N_6599);
and U14476 (N_14476,N_9170,N_8820);
or U14477 (N_14477,N_6769,N_5549);
and U14478 (N_14478,N_9040,N_8663);
or U14479 (N_14479,N_8247,N_9858);
or U14480 (N_14480,N_6404,N_5173);
and U14481 (N_14481,N_8948,N_5539);
and U14482 (N_14482,N_9233,N_5089);
or U14483 (N_14483,N_7583,N_9519);
and U14484 (N_14484,N_5694,N_7858);
nor U14485 (N_14485,N_6844,N_5596);
or U14486 (N_14486,N_8678,N_9751);
nand U14487 (N_14487,N_7102,N_8214);
xor U14488 (N_14488,N_8162,N_5005);
and U14489 (N_14489,N_7177,N_8420);
nor U14490 (N_14490,N_9556,N_6717);
nor U14491 (N_14491,N_6065,N_9188);
nor U14492 (N_14492,N_9637,N_6492);
and U14493 (N_14493,N_5061,N_7641);
and U14494 (N_14494,N_5024,N_6090);
nand U14495 (N_14495,N_7067,N_7525);
nor U14496 (N_14496,N_5905,N_8009);
nand U14497 (N_14497,N_7467,N_9584);
or U14498 (N_14498,N_5511,N_5649);
and U14499 (N_14499,N_9634,N_9002);
and U14500 (N_14500,N_6645,N_8244);
and U14501 (N_14501,N_8184,N_8464);
nor U14502 (N_14502,N_6937,N_9911);
nor U14503 (N_14503,N_9158,N_8717);
nor U14504 (N_14504,N_7278,N_6109);
nand U14505 (N_14505,N_9660,N_8399);
or U14506 (N_14506,N_9301,N_8609);
and U14507 (N_14507,N_7015,N_5573);
nor U14508 (N_14508,N_7468,N_6545);
nand U14509 (N_14509,N_5312,N_5049);
or U14510 (N_14510,N_8694,N_9572);
or U14511 (N_14511,N_9906,N_9758);
nand U14512 (N_14512,N_7144,N_9620);
nor U14513 (N_14513,N_7299,N_7180);
nand U14514 (N_14514,N_8066,N_9878);
nor U14515 (N_14515,N_8421,N_9594);
nor U14516 (N_14516,N_5356,N_9270);
nor U14517 (N_14517,N_5481,N_5505);
nor U14518 (N_14518,N_8163,N_8806);
and U14519 (N_14519,N_8729,N_9745);
and U14520 (N_14520,N_6951,N_9600);
nor U14521 (N_14521,N_7659,N_9849);
or U14522 (N_14522,N_6619,N_7891);
nand U14523 (N_14523,N_7685,N_8205);
nand U14524 (N_14524,N_5814,N_9581);
and U14525 (N_14525,N_9246,N_7823);
nand U14526 (N_14526,N_7846,N_9729);
and U14527 (N_14527,N_8447,N_7875);
or U14528 (N_14528,N_8207,N_7349);
nand U14529 (N_14529,N_9286,N_6927);
and U14530 (N_14530,N_6682,N_5185);
nor U14531 (N_14531,N_6839,N_9826);
and U14532 (N_14532,N_8029,N_9254);
nor U14533 (N_14533,N_6010,N_8871);
or U14534 (N_14534,N_8057,N_9471);
and U14535 (N_14535,N_7906,N_7105);
nor U14536 (N_14536,N_8837,N_8176);
nor U14537 (N_14537,N_6574,N_6818);
or U14538 (N_14538,N_5658,N_6494);
nand U14539 (N_14539,N_9231,N_9272);
and U14540 (N_14540,N_6742,N_7338);
nor U14541 (N_14541,N_9790,N_5745);
nor U14542 (N_14542,N_9068,N_6620);
and U14543 (N_14543,N_5576,N_9807);
nor U14544 (N_14544,N_9313,N_9567);
nand U14545 (N_14545,N_6747,N_9012);
and U14546 (N_14546,N_7956,N_7997);
or U14547 (N_14547,N_9442,N_8057);
and U14548 (N_14548,N_9941,N_5406);
nor U14549 (N_14549,N_6462,N_7967);
nor U14550 (N_14550,N_8498,N_9825);
nand U14551 (N_14551,N_6317,N_6495);
nor U14552 (N_14552,N_5542,N_6594);
nor U14553 (N_14553,N_6188,N_9870);
and U14554 (N_14554,N_7038,N_6886);
or U14555 (N_14555,N_7794,N_9966);
nor U14556 (N_14556,N_9986,N_5770);
and U14557 (N_14557,N_6618,N_9916);
nand U14558 (N_14558,N_7404,N_7215);
nand U14559 (N_14559,N_8288,N_9784);
and U14560 (N_14560,N_8064,N_7860);
or U14561 (N_14561,N_7758,N_5361);
nand U14562 (N_14562,N_6508,N_6754);
nand U14563 (N_14563,N_7394,N_6656);
nor U14564 (N_14564,N_6804,N_8559);
or U14565 (N_14565,N_5930,N_9017);
nand U14566 (N_14566,N_8639,N_8243);
nor U14567 (N_14567,N_8190,N_6713);
nor U14568 (N_14568,N_7928,N_6953);
nor U14569 (N_14569,N_5384,N_8547);
and U14570 (N_14570,N_9484,N_7956);
or U14571 (N_14571,N_9841,N_9346);
or U14572 (N_14572,N_5993,N_8744);
or U14573 (N_14573,N_6096,N_7164);
nor U14574 (N_14574,N_6446,N_8423);
nor U14575 (N_14575,N_8443,N_7452);
nor U14576 (N_14576,N_7254,N_9151);
and U14577 (N_14577,N_7964,N_6380);
or U14578 (N_14578,N_6120,N_7531);
or U14579 (N_14579,N_8459,N_9928);
and U14580 (N_14580,N_9586,N_6241);
and U14581 (N_14581,N_5949,N_9043);
nand U14582 (N_14582,N_8168,N_5384);
nand U14583 (N_14583,N_6496,N_9943);
and U14584 (N_14584,N_9120,N_8914);
and U14585 (N_14585,N_8973,N_5251);
and U14586 (N_14586,N_6955,N_6539);
or U14587 (N_14587,N_8146,N_5896);
nand U14588 (N_14588,N_6467,N_7354);
and U14589 (N_14589,N_7832,N_9107);
nor U14590 (N_14590,N_7569,N_7909);
nor U14591 (N_14591,N_7076,N_5946);
and U14592 (N_14592,N_8205,N_6666);
and U14593 (N_14593,N_8497,N_8435);
and U14594 (N_14594,N_5594,N_6371);
and U14595 (N_14595,N_8173,N_5177);
and U14596 (N_14596,N_7701,N_8599);
nor U14597 (N_14597,N_6000,N_5218);
nor U14598 (N_14598,N_6018,N_8616);
and U14599 (N_14599,N_5525,N_7574);
or U14600 (N_14600,N_9551,N_5949);
nor U14601 (N_14601,N_9727,N_5554);
nor U14602 (N_14602,N_5375,N_6332);
nor U14603 (N_14603,N_5165,N_5530);
and U14604 (N_14604,N_5498,N_5315);
nor U14605 (N_14605,N_5992,N_6392);
and U14606 (N_14606,N_9421,N_7795);
and U14607 (N_14607,N_9327,N_6303);
nand U14608 (N_14608,N_7920,N_7099);
xnor U14609 (N_14609,N_5004,N_6048);
and U14610 (N_14610,N_9939,N_7183);
nand U14611 (N_14611,N_9565,N_6854);
or U14612 (N_14612,N_7545,N_5194);
nor U14613 (N_14613,N_8953,N_9390);
or U14614 (N_14614,N_7118,N_6838);
and U14615 (N_14615,N_7646,N_8593);
and U14616 (N_14616,N_6426,N_7518);
or U14617 (N_14617,N_5143,N_5494);
nand U14618 (N_14618,N_8243,N_6724);
nor U14619 (N_14619,N_6986,N_8817);
nor U14620 (N_14620,N_6427,N_5763);
nor U14621 (N_14621,N_9691,N_5324);
nand U14622 (N_14622,N_8626,N_7909);
and U14623 (N_14623,N_8991,N_8873);
or U14624 (N_14624,N_5918,N_9203);
nor U14625 (N_14625,N_8541,N_8040);
or U14626 (N_14626,N_8296,N_7418);
nand U14627 (N_14627,N_6766,N_7652);
xnor U14628 (N_14628,N_9207,N_7597);
and U14629 (N_14629,N_7149,N_6628);
or U14630 (N_14630,N_6067,N_6290);
nor U14631 (N_14631,N_6026,N_7962);
or U14632 (N_14632,N_8835,N_9149);
nand U14633 (N_14633,N_6152,N_7310);
nand U14634 (N_14634,N_5409,N_8974);
and U14635 (N_14635,N_7307,N_7754);
nor U14636 (N_14636,N_8580,N_6867);
nor U14637 (N_14637,N_8597,N_7323);
nor U14638 (N_14638,N_9756,N_5687);
or U14639 (N_14639,N_7563,N_5533);
nand U14640 (N_14640,N_6276,N_5590);
and U14641 (N_14641,N_7657,N_9561);
nand U14642 (N_14642,N_8785,N_7607);
nand U14643 (N_14643,N_5870,N_7974);
nor U14644 (N_14644,N_7488,N_5500);
nand U14645 (N_14645,N_7387,N_5629);
and U14646 (N_14646,N_9371,N_8976);
and U14647 (N_14647,N_8306,N_6523);
nor U14648 (N_14648,N_8178,N_6151);
nor U14649 (N_14649,N_8348,N_5323);
nor U14650 (N_14650,N_7991,N_8281);
and U14651 (N_14651,N_8828,N_9929);
or U14652 (N_14652,N_8376,N_5269);
and U14653 (N_14653,N_5508,N_7851);
nand U14654 (N_14654,N_8926,N_9406);
and U14655 (N_14655,N_5065,N_8982);
and U14656 (N_14656,N_9830,N_8053);
and U14657 (N_14657,N_5738,N_8497);
nand U14658 (N_14658,N_6497,N_7107);
nand U14659 (N_14659,N_6506,N_8435);
nor U14660 (N_14660,N_6087,N_6538);
nand U14661 (N_14661,N_6638,N_5825);
or U14662 (N_14662,N_7798,N_6402);
nor U14663 (N_14663,N_8602,N_9854);
nor U14664 (N_14664,N_7443,N_7742);
xor U14665 (N_14665,N_9207,N_7558);
or U14666 (N_14666,N_8716,N_7824);
nand U14667 (N_14667,N_6835,N_6125);
and U14668 (N_14668,N_7351,N_7702);
and U14669 (N_14669,N_7296,N_9859);
nand U14670 (N_14670,N_5627,N_8197);
or U14671 (N_14671,N_5874,N_5988);
or U14672 (N_14672,N_6899,N_9478);
and U14673 (N_14673,N_8918,N_7209);
and U14674 (N_14674,N_5903,N_5048);
nand U14675 (N_14675,N_8417,N_7157);
or U14676 (N_14676,N_5003,N_9488);
and U14677 (N_14677,N_7045,N_7372);
and U14678 (N_14678,N_8716,N_7901);
nor U14679 (N_14679,N_6495,N_8672);
and U14680 (N_14680,N_9944,N_8244);
nor U14681 (N_14681,N_6469,N_5880);
or U14682 (N_14682,N_7538,N_6119);
and U14683 (N_14683,N_9910,N_6263);
nand U14684 (N_14684,N_6052,N_8847);
nand U14685 (N_14685,N_9417,N_8358);
nor U14686 (N_14686,N_6911,N_8734);
nand U14687 (N_14687,N_8826,N_7631);
or U14688 (N_14688,N_5553,N_8447);
nand U14689 (N_14689,N_6553,N_8812);
nor U14690 (N_14690,N_5552,N_9231);
or U14691 (N_14691,N_8063,N_6574);
and U14692 (N_14692,N_7610,N_9175);
or U14693 (N_14693,N_8456,N_5477);
nand U14694 (N_14694,N_8072,N_9874);
or U14695 (N_14695,N_6232,N_9813);
nand U14696 (N_14696,N_9484,N_5406);
nand U14697 (N_14697,N_5443,N_9968);
and U14698 (N_14698,N_9145,N_6827);
nor U14699 (N_14699,N_8171,N_6687);
nor U14700 (N_14700,N_6269,N_8454);
nor U14701 (N_14701,N_5105,N_6723);
and U14702 (N_14702,N_6330,N_8537);
nor U14703 (N_14703,N_6983,N_6195);
xnor U14704 (N_14704,N_7828,N_9196);
nor U14705 (N_14705,N_7528,N_9781);
nand U14706 (N_14706,N_6349,N_9468);
and U14707 (N_14707,N_7759,N_7034);
nor U14708 (N_14708,N_9226,N_7840);
and U14709 (N_14709,N_9363,N_8599);
or U14710 (N_14710,N_9377,N_7217);
and U14711 (N_14711,N_8077,N_9924);
nand U14712 (N_14712,N_7327,N_8328);
nor U14713 (N_14713,N_9653,N_8736);
nand U14714 (N_14714,N_5674,N_7661);
or U14715 (N_14715,N_6154,N_5312);
or U14716 (N_14716,N_8447,N_7087);
nor U14717 (N_14717,N_9638,N_6976);
xor U14718 (N_14718,N_5005,N_8101);
nor U14719 (N_14719,N_7541,N_6674);
or U14720 (N_14720,N_5888,N_7578);
nand U14721 (N_14721,N_6264,N_8312);
or U14722 (N_14722,N_8715,N_8721);
nand U14723 (N_14723,N_7653,N_6126);
or U14724 (N_14724,N_5380,N_8972);
and U14725 (N_14725,N_5631,N_9709);
and U14726 (N_14726,N_8490,N_7425);
nor U14727 (N_14727,N_5148,N_5997);
and U14728 (N_14728,N_7696,N_5559);
or U14729 (N_14729,N_6206,N_7675);
nor U14730 (N_14730,N_9451,N_8103);
and U14731 (N_14731,N_5647,N_6250);
and U14732 (N_14732,N_8053,N_8019);
nand U14733 (N_14733,N_8992,N_7978);
nand U14734 (N_14734,N_9303,N_5754);
and U14735 (N_14735,N_7847,N_6140);
and U14736 (N_14736,N_6102,N_5643);
nand U14737 (N_14737,N_7835,N_6176);
nand U14738 (N_14738,N_6785,N_5974);
nor U14739 (N_14739,N_6254,N_6808);
and U14740 (N_14740,N_8798,N_9434);
and U14741 (N_14741,N_6683,N_9533);
nor U14742 (N_14742,N_6295,N_6396);
nor U14743 (N_14743,N_7463,N_5372);
or U14744 (N_14744,N_5346,N_8397);
and U14745 (N_14745,N_8306,N_5721);
nor U14746 (N_14746,N_9186,N_6805);
or U14747 (N_14747,N_6767,N_9938);
nor U14748 (N_14748,N_8486,N_6085);
nand U14749 (N_14749,N_8440,N_7590);
and U14750 (N_14750,N_6338,N_9724);
nand U14751 (N_14751,N_7278,N_8399);
nand U14752 (N_14752,N_8736,N_9615);
nor U14753 (N_14753,N_7284,N_7568);
nor U14754 (N_14754,N_8217,N_6067);
or U14755 (N_14755,N_9142,N_5982);
nand U14756 (N_14756,N_8964,N_6363);
and U14757 (N_14757,N_9100,N_8546);
nand U14758 (N_14758,N_9037,N_8821);
nor U14759 (N_14759,N_8581,N_7740);
nand U14760 (N_14760,N_5105,N_8096);
and U14761 (N_14761,N_8486,N_7374);
nand U14762 (N_14762,N_5061,N_7210);
nor U14763 (N_14763,N_8430,N_8376);
nor U14764 (N_14764,N_6569,N_9217);
nand U14765 (N_14765,N_8238,N_9910);
nor U14766 (N_14766,N_5098,N_9859);
nand U14767 (N_14767,N_5573,N_8482);
and U14768 (N_14768,N_9945,N_8842);
or U14769 (N_14769,N_7341,N_6304);
nor U14770 (N_14770,N_7731,N_7104);
nor U14771 (N_14771,N_7582,N_9459);
or U14772 (N_14772,N_5856,N_7791);
xnor U14773 (N_14773,N_9101,N_6275);
or U14774 (N_14774,N_5449,N_8280);
or U14775 (N_14775,N_8294,N_8784);
or U14776 (N_14776,N_9090,N_6058);
nand U14777 (N_14777,N_7018,N_9785);
nor U14778 (N_14778,N_6395,N_8779);
nand U14779 (N_14779,N_6300,N_8524);
or U14780 (N_14780,N_7434,N_8776);
and U14781 (N_14781,N_6289,N_6929);
nand U14782 (N_14782,N_8570,N_5561);
nor U14783 (N_14783,N_7701,N_8251);
nor U14784 (N_14784,N_7264,N_8971);
nand U14785 (N_14785,N_7295,N_9237);
nor U14786 (N_14786,N_7309,N_5119);
nand U14787 (N_14787,N_6123,N_8243);
nor U14788 (N_14788,N_8736,N_9724);
nor U14789 (N_14789,N_8417,N_8252);
and U14790 (N_14790,N_9737,N_7936);
and U14791 (N_14791,N_5861,N_7628);
and U14792 (N_14792,N_5015,N_6218);
or U14793 (N_14793,N_8886,N_8892);
and U14794 (N_14794,N_6925,N_7593);
and U14795 (N_14795,N_8832,N_7654);
nand U14796 (N_14796,N_5078,N_9970);
nand U14797 (N_14797,N_6265,N_8086);
or U14798 (N_14798,N_9180,N_7008);
nand U14799 (N_14799,N_7768,N_7622);
nor U14800 (N_14800,N_7874,N_9890);
or U14801 (N_14801,N_7791,N_9846);
and U14802 (N_14802,N_9408,N_5186);
or U14803 (N_14803,N_5686,N_6734);
nor U14804 (N_14804,N_8834,N_7605);
and U14805 (N_14805,N_7042,N_7300);
nand U14806 (N_14806,N_5055,N_5856);
or U14807 (N_14807,N_7493,N_6037);
nor U14808 (N_14808,N_7898,N_9016);
or U14809 (N_14809,N_7062,N_8648);
and U14810 (N_14810,N_8400,N_8772);
nor U14811 (N_14811,N_5436,N_5115);
and U14812 (N_14812,N_9235,N_9909);
or U14813 (N_14813,N_5608,N_7744);
nand U14814 (N_14814,N_8143,N_7167);
nand U14815 (N_14815,N_7029,N_5578);
or U14816 (N_14816,N_8797,N_8991);
and U14817 (N_14817,N_7560,N_8566);
nand U14818 (N_14818,N_7087,N_6286);
nand U14819 (N_14819,N_8051,N_7492);
nand U14820 (N_14820,N_9974,N_6981);
or U14821 (N_14821,N_7308,N_9340);
nand U14822 (N_14822,N_8441,N_6461);
nor U14823 (N_14823,N_5204,N_5139);
nor U14824 (N_14824,N_5709,N_7529);
and U14825 (N_14825,N_7884,N_5960);
and U14826 (N_14826,N_5854,N_9931);
nor U14827 (N_14827,N_6817,N_9377);
or U14828 (N_14828,N_8551,N_9769);
and U14829 (N_14829,N_8442,N_5949);
nor U14830 (N_14830,N_9552,N_8371);
or U14831 (N_14831,N_5226,N_8594);
and U14832 (N_14832,N_9121,N_8540);
nor U14833 (N_14833,N_9812,N_8724);
nand U14834 (N_14834,N_9264,N_8657);
and U14835 (N_14835,N_6566,N_7328);
or U14836 (N_14836,N_7684,N_5978);
nor U14837 (N_14837,N_7756,N_9536);
nor U14838 (N_14838,N_6246,N_9959);
or U14839 (N_14839,N_6881,N_5323);
or U14840 (N_14840,N_5925,N_7468);
and U14841 (N_14841,N_7772,N_6126);
and U14842 (N_14842,N_7124,N_5259);
and U14843 (N_14843,N_6861,N_9095);
and U14844 (N_14844,N_7352,N_8891);
nor U14845 (N_14845,N_7724,N_6452);
nor U14846 (N_14846,N_6904,N_5283);
nand U14847 (N_14847,N_6765,N_5824);
and U14848 (N_14848,N_8886,N_6537);
nor U14849 (N_14849,N_5542,N_6811);
nand U14850 (N_14850,N_6171,N_9628);
nand U14851 (N_14851,N_7753,N_6512);
and U14852 (N_14852,N_6624,N_6077);
nor U14853 (N_14853,N_7638,N_6403);
or U14854 (N_14854,N_8258,N_8550);
nand U14855 (N_14855,N_9921,N_9665);
or U14856 (N_14856,N_8505,N_5321);
nand U14857 (N_14857,N_5623,N_5920);
nand U14858 (N_14858,N_6350,N_5737);
or U14859 (N_14859,N_8326,N_6905);
nor U14860 (N_14860,N_9311,N_8671);
nor U14861 (N_14861,N_9815,N_8556);
nand U14862 (N_14862,N_7867,N_7719);
or U14863 (N_14863,N_7828,N_8602);
or U14864 (N_14864,N_9778,N_6868);
nor U14865 (N_14865,N_9488,N_5361);
nor U14866 (N_14866,N_7079,N_7742);
or U14867 (N_14867,N_9255,N_5129);
nand U14868 (N_14868,N_6540,N_8461);
or U14869 (N_14869,N_6272,N_6116);
xor U14870 (N_14870,N_5369,N_5926);
and U14871 (N_14871,N_8828,N_5914);
or U14872 (N_14872,N_8075,N_7841);
nor U14873 (N_14873,N_9789,N_5457);
nor U14874 (N_14874,N_6399,N_5923);
and U14875 (N_14875,N_9756,N_8075);
and U14876 (N_14876,N_8836,N_8317);
nand U14877 (N_14877,N_7515,N_5600);
or U14878 (N_14878,N_7836,N_5164);
or U14879 (N_14879,N_5393,N_5420);
nor U14880 (N_14880,N_8112,N_9236);
nand U14881 (N_14881,N_7053,N_8320);
nor U14882 (N_14882,N_8129,N_8051);
nor U14883 (N_14883,N_6163,N_8980);
nand U14884 (N_14884,N_8465,N_7817);
nor U14885 (N_14885,N_5982,N_9909);
and U14886 (N_14886,N_5088,N_6988);
nor U14887 (N_14887,N_9048,N_7417);
and U14888 (N_14888,N_5700,N_9313);
nand U14889 (N_14889,N_7822,N_6668);
and U14890 (N_14890,N_9231,N_8984);
xnor U14891 (N_14891,N_8714,N_5172);
and U14892 (N_14892,N_6980,N_8114);
and U14893 (N_14893,N_9317,N_8370);
and U14894 (N_14894,N_7323,N_6429);
or U14895 (N_14895,N_5803,N_5689);
nor U14896 (N_14896,N_9516,N_5780);
nand U14897 (N_14897,N_8020,N_6171);
nand U14898 (N_14898,N_7869,N_8604);
xnor U14899 (N_14899,N_8207,N_8399);
or U14900 (N_14900,N_5549,N_9816);
nand U14901 (N_14901,N_6381,N_7328);
nand U14902 (N_14902,N_8860,N_6923);
or U14903 (N_14903,N_9169,N_8132);
nand U14904 (N_14904,N_9927,N_8604);
and U14905 (N_14905,N_7590,N_5098);
and U14906 (N_14906,N_7058,N_5521);
nor U14907 (N_14907,N_6048,N_7313);
and U14908 (N_14908,N_8788,N_5061);
nor U14909 (N_14909,N_5367,N_6248);
and U14910 (N_14910,N_7632,N_5683);
nand U14911 (N_14911,N_5675,N_6356);
nand U14912 (N_14912,N_9987,N_9862);
nand U14913 (N_14913,N_7193,N_9827);
and U14914 (N_14914,N_7993,N_5613);
and U14915 (N_14915,N_7887,N_9644);
and U14916 (N_14916,N_5908,N_8609);
xor U14917 (N_14917,N_5487,N_5696);
and U14918 (N_14918,N_8767,N_5865);
and U14919 (N_14919,N_9335,N_5867);
nand U14920 (N_14920,N_5256,N_6465);
nor U14921 (N_14921,N_6742,N_6475);
nand U14922 (N_14922,N_7300,N_8989);
or U14923 (N_14923,N_9799,N_8404);
nor U14924 (N_14924,N_7232,N_7193);
or U14925 (N_14925,N_8328,N_9268);
or U14926 (N_14926,N_6145,N_5741);
nand U14927 (N_14927,N_7872,N_9169);
nor U14928 (N_14928,N_5676,N_8128);
nor U14929 (N_14929,N_9234,N_5185);
or U14930 (N_14930,N_6122,N_8271);
nor U14931 (N_14931,N_6083,N_9809);
and U14932 (N_14932,N_8323,N_5924);
and U14933 (N_14933,N_9502,N_5561);
and U14934 (N_14934,N_6475,N_8532);
nand U14935 (N_14935,N_6895,N_7930);
and U14936 (N_14936,N_7790,N_6044);
and U14937 (N_14937,N_5934,N_9946);
and U14938 (N_14938,N_8929,N_7585);
nor U14939 (N_14939,N_7738,N_5993);
or U14940 (N_14940,N_5617,N_9662);
nand U14941 (N_14941,N_9829,N_7266);
or U14942 (N_14942,N_6722,N_9885);
and U14943 (N_14943,N_8205,N_6601);
or U14944 (N_14944,N_5421,N_6784);
and U14945 (N_14945,N_7002,N_6990);
or U14946 (N_14946,N_7794,N_6612);
or U14947 (N_14947,N_8961,N_6620);
and U14948 (N_14948,N_8732,N_6053);
or U14949 (N_14949,N_8981,N_6184);
nand U14950 (N_14950,N_7104,N_6068);
or U14951 (N_14951,N_7586,N_6655);
or U14952 (N_14952,N_9853,N_8903);
or U14953 (N_14953,N_6632,N_9260);
and U14954 (N_14954,N_8148,N_5869);
or U14955 (N_14955,N_6380,N_5287);
nor U14956 (N_14956,N_5784,N_9712);
nand U14957 (N_14957,N_9329,N_5262);
nor U14958 (N_14958,N_7656,N_8837);
nor U14959 (N_14959,N_6289,N_8097);
nor U14960 (N_14960,N_5243,N_9455);
and U14961 (N_14961,N_6788,N_6983);
nor U14962 (N_14962,N_9805,N_6027);
nand U14963 (N_14963,N_8070,N_5738);
nand U14964 (N_14964,N_6427,N_6971);
and U14965 (N_14965,N_6505,N_9084);
nand U14966 (N_14966,N_6082,N_8564);
nor U14967 (N_14967,N_5753,N_8927);
nor U14968 (N_14968,N_9213,N_8415);
or U14969 (N_14969,N_5450,N_9519);
and U14970 (N_14970,N_8727,N_8182);
nor U14971 (N_14971,N_6697,N_5468);
nor U14972 (N_14972,N_5027,N_8608);
or U14973 (N_14973,N_6756,N_6122);
and U14974 (N_14974,N_7721,N_7999);
and U14975 (N_14975,N_9687,N_9973);
or U14976 (N_14976,N_8329,N_9347);
nand U14977 (N_14977,N_9354,N_6074);
nand U14978 (N_14978,N_9193,N_5938);
nand U14979 (N_14979,N_9871,N_7904);
and U14980 (N_14980,N_5281,N_9599);
nand U14981 (N_14981,N_8714,N_9382);
nand U14982 (N_14982,N_6890,N_6111);
and U14983 (N_14983,N_6834,N_7747);
nand U14984 (N_14984,N_5365,N_8039);
or U14985 (N_14985,N_7434,N_7402);
and U14986 (N_14986,N_5825,N_8856);
nor U14987 (N_14987,N_7778,N_9138);
or U14988 (N_14988,N_9375,N_9711);
or U14989 (N_14989,N_9368,N_8402);
and U14990 (N_14990,N_8385,N_7734);
or U14991 (N_14991,N_8195,N_7142);
nor U14992 (N_14992,N_6435,N_5409);
nor U14993 (N_14993,N_5329,N_5791);
and U14994 (N_14994,N_9136,N_7036);
nor U14995 (N_14995,N_6903,N_5461);
or U14996 (N_14996,N_7045,N_6634);
xor U14997 (N_14997,N_6141,N_8750);
nand U14998 (N_14998,N_7819,N_7150);
or U14999 (N_14999,N_5578,N_9791);
nand UO_0 (O_0,N_14621,N_10063);
nor UO_1 (O_1,N_11751,N_13041);
and UO_2 (O_2,N_14449,N_12657);
or UO_3 (O_3,N_11067,N_14413);
and UO_4 (O_4,N_14527,N_10509);
nand UO_5 (O_5,N_12180,N_14182);
and UO_6 (O_6,N_14942,N_11155);
or UO_7 (O_7,N_11034,N_14478);
nand UO_8 (O_8,N_11695,N_10416);
nor UO_9 (O_9,N_10668,N_12623);
and UO_10 (O_10,N_11427,N_13474);
and UO_11 (O_11,N_14195,N_12149);
nand UO_12 (O_12,N_14596,N_13832);
and UO_13 (O_13,N_13482,N_10938);
or UO_14 (O_14,N_11259,N_14678);
xor UO_15 (O_15,N_13451,N_11534);
and UO_16 (O_16,N_13711,N_11422);
or UO_17 (O_17,N_13740,N_11026);
and UO_18 (O_18,N_11805,N_11320);
or UO_19 (O_19,N_14444,N_12058);
and UO_20 (O_20,N_12888,N_14907);
nand UO_21 (O_21,N_13085,N_11540);
nand UO_22 (O_22,N_10201,N_12636);
nor UO_23 (O_23,N_10500,N_11296);
nor UO_24 (O_24,N_12785,N_13863);
and UO_25 (O_25,N_13860,N_11410);
or UO_26 (O_26,N_14177,N_14381);
or UO_27 (O_27,N_13647,N_11232);
nor UO_28 (O_28,N_12231,N_12729);
or UO_29 (O_29,N_14622,N_13859);
and UO_30 (O_30,N_13987,N_13389);
nand UO_31 (O_31,N_10343,N_11527);
nand UO_32 (O_32,N_13761,N_10324);
nor UO_33 (O_33,N_10433,N_10771);
nand UO_34 (O_34,N_12800,N_14467);
nand UO_35 (O_35,N_11045,N_11866);
nor UO_36 (O_36,N_14610,N_10196);
or UO_37 (O_37,N_13927,N_11475);
and UO_38 (O_38,N_12304,N_12196);
xor UO_39 (O_39,N_11097,N_11716);
and UO_40 (O_40,N_14530,N_10559);
nand UO_41 (O_41,N_14924,N_12339);
and UO_42 (O_42,N_10532,N_13469);
nand UO_43 (O_43,N_13931,N_10318);
nor UO_44 (O_44,N_12583,N_13967);
nand UO_45 (O_45,N_12336,N_14531);
nand UO_46 (O_46,N_11501,N_14109);
and UO_47 (O_47,N_11450,N_13108);
or UO_48 (O_48,N_14783,N_14434);
or UO_49 (O_49,N_10138,N_14296);
nand UO_50 (O_50,N_10161,N_11869);
xor UO_51 (O_51,N_10592,N_13536);
and UO_52 (O_52,N_13962,N_14380);
nand UO_53 (O_53,N_14710,N_11612);
or UO_54 (O_54,N_13112,N_12014);
nor UO_55 (O_55,N_12588,N_11190);
nand UO_56 (O_56,N_13964,N_12876);
or UO_57 (O_57,N_12215,N_11928);
or UO_58 (O_58,N_14994,N_14266);
or UO_59 (O_59,N_11400,N_12438);
and UO_60 (O_60,N_10855,N_10317);
nor UO_61 (O_61,N_11056,N_13159);
or UO_62 (O_62,N_10437,N_11680);
nand UO_63 (O_63,N_13485,N_11003);
and UO_64 (O_64,N_14702,N_11878);
and UO_65 (O_65,N_10417,N_10849);
nand UO_66 (O_66,N_11614,N_14362);
or UO_67 (O_67,N_14323,N_13192);
or UO_68 (O_68,N_12227,N_12786);
and UO_69 (O_69,N_14164,N_11474);
or UO_70 (O_70,N_10399,N_12598);
nor UO_71 (O_71,N_14893,N_13988);
and UO_72 (O_72,N_11014,N_13201);
and UO_73 (O_73,N_11967,N_10402);
nand UO_74 (O_74,N_14800,N_12504);
nand UO_75 (O_75,N_13925,N_12272);
nor UO_76 (O_76,N_13605,N_11033);
and UO_77 (O_77,N_14423,N_10734);
and UO_78 (O_78,N_14570,N_12854);
and UO_79 (O_79,N_12021,N_11754);
and UO_80 (O_80,N_11094,N_12124);
and UO_81 (O_81,N_10803,N_14421);
or UO_82 (O_82,N_11797,N_11982);
xor UO_83 (O_83,N_12698,N_13214);
and UO_84 (O_84,N_13680,N_10154);
and UO_85 (O_85,N_13454,N_14768);
nand UO_86 (O_86,N_13720,N_12942);
or UO_87 (O_87,N_10413,N_10242);
or UO_88 (O_88,N_13488,N_10095);
or UO_89 (O_89,N_14680,N_13417);
and UO_90 (O_90,N_12517,N_12479);
and UO_91 (O_91,N_12714,N_14754);
nand UO_92 (O_92,N_10332,N_14488);
or UO_93 (O_93,N_14244,N_14432);
or UO_94 (O_94,N_10877,N_10105);
or UO_95 (O_95,N_12743,N_12594);
nand UO_96 (O_96,N_14493,N_10140);
nand UO_97 (O_97,N_10330,N_12547);
and UO_98 (O_98,N_11550,N_10932);
or UO_99 (O_99,N_12857,N_10542);
and UO_100 (O_100,N_13833,N_12917);
nand UO_101 (O_101,N_11576,N_14455);
nand UO_102 (O_102,N_13718,N_11502);
nor UO_103 (O_103,N_13447,N_10456);
nor UO_104 (O_104,N_13480,N_11404);
nor UO_105 (O_105,N_12461,N_10582);
nand UO_106 (O_106,N_14275,N_11807);
or UO_107 (O_107,N_10223,N_12884);
nor UO_108 (O_108,N_10577,N_10455);
nor UO_109 (O_109,N_10011,N_10584);
nand UO_110 (O_110,N_13500,N_12817);
and UO_111 (O_111,N_14854,N_13935);
xor UO_112 (O_112,N_13478,N_13137);
nand UO_113 (O_113,N_14750,N_10609);
nand UO_114 (O_114,N_11770,N_14874);
or UO_115 (O_115,N_11916,N_11592);
nor UO_116 (O_116,N_11909,N_12205);
nand UO_117 (O_117,N_10810,N_11420);
and UO_118 (O_118,N_14262,N_11511);
nor UO_119 (O_119,N_10867,N_11029);
and UO_120 (O_120,N_14869,N_11949);
nor UO_121 (O_121,N_13800,N_14221);
or UO_122 (O_122,N_12390,N_12125);
nand UO_123 (O_123,N_13932,N_12839);
nor UO_124 (O_124,N_12522,N_14475);
nor UO_125 (O_125,N_12428,N_11104);
nor UO_126 (O_126,N_12984,N_10664);
and UO_127 (O_127,N_13381,N_12142);
or UO_128 (O_128,N_10558,N_10380);
and UO_129 (O_129,N_11268,N_14339);
or UO_130 (O_130,N_14709,N_10238);
and UO_131 (O_131,N_11374,N_13830);
nor UO_132 (O_132,N_13788,N_11719);
and UO_133 (O_133,N_12943,N_14405);
nor UO_134 (O_134,N_11039,N_12110);
nand UO_135 (O_135,N_10436,N_12643);
and UO_136 (O_136,N_11713,N_13261);
nand UO_137 (O_137,N_14976,N_13604);
nor UO_138 (O_138,N_12858,N_14480);
or UO_139 (O_139,N_10106,N_12118);
and UO_140 (O_140,N_11922,N_10439);
or UO_141 (O_141,N_13246,N_10370);
and UO_142 (O_142,N_14400,N_10697);
nand UO_143 (O_143,N_11962,N_14500);
nand UO_144 (O_144,N_14201,N_14495);
and UO_145 (O_145,N_11961,N_14818);
nor UO_146 (O_146,N_12503,N_14028);
or UO_147 (O_147,N_10367,N_14473);
nor UO_148 (O_148,N_12027,N_14871);
nor UO_149 (O_149,N_14850,N_13467);
nor UO_150 (O_150,N_12426,N_10146);
and UO_151 (O_151,N_14767,N_13837);
or UO_152 (O_152,N_11447,N_14592);
or UO_153 (O_153,N_14061,N_11757);
or UO_154 (O_154,N_14199,N_13651);
or UO_155 (O_155,N_11759,N_13323);
or UO_156 (O_156,N_13687,N_13899);
nand UO_157 (O_157,N_13065,N_13911);
or UO_158 (O_158,N_10199,N_14411);
or UO_159 (O_159,N_14327,N_10818);
nand UO_160 (O_160,N_13476,N_14008);
or UO_161 (O_161,N_10192,N_12606);
and UO_162 (O_162,N_12085,N_11388);
nand UO_163 (O_163,N_14471,N_13385);
nor UO_164 (O_164,N_12105,N_11654);
and UO_165 (O_165,N_13477,N_13360);
and UO_166 (O_166,N_14312,N_11459);
nand UO_167 (O_167,N_10198,N_14903);
and UO_168 (O_168,N_11358,N_12431);
or UO_169 (O_169,N_13363,N_14052);
nand UO_170 (O_170,N_14066,N_12945);
and UO_171 (O_171,N_11547,N_14016);
or UO_172 (O_172,N_10236,N_10164);
nand UO_173 (O_173,N_13742,N_12930);
xnor UO_174 (O_174,N_11860,N_13048);
or UO_175 (O_175,N_11673,N_12368);
nand UO_176 (O_176,N_11817,N_10895);
nand UO_177 (O_177,N_12006,N_13691);
and UO_178 (O_178,N_10638,N_13587);
and UO_179 (O_179,N_10406,N_12948);
or UO_180 (O_180,N_11477,N_13876);
or UO_181 (O_181,N_14307,N_12007);
nor UO_182 (O_182,N_12892,N_13044);
nand UO_183 (O_183,N_12312,N_11121);
and UO_184 (O_184,N_12031,N_12561);
nand UO_185 (O_185,N_10117,N_14820);
nor UO_186 (O_186,N_10982,N_11216);
nor UO_187 (O_187,N_13103,N_12832);
and UO_188 (O_188,N_12315,N_11563);
or UO_189 (O_189,N_11266,N_13064);
nor UO_190 (O_190,N_12274,N_14890);
or UO_191 (O_191,N_14420,N_10615);
nor UO_192 (O_192,N_14576,N_14574);
nand UO_193 (O_193,N_10457,N_12516);
and UO_194 (O_194,N_10791,N_14360);
nand UO_195 (O_195,N_11015,N_10873);
and UO_196 (O_196,N_10156,N_13423);
or UO_197 (O_197,N_10919,N_12655);
and UO_198 (O_198,N_10915,N_13151);
or UO_199 (O_199,N_13255,N_12760);
nand UO_200 (O_200,N_13063,N_14039);
nand UO_201 (O_201,N_12557,N_10033);
nor UO_202 (O_202,N_13353,N_14704);
nand UO_203 (O_203,N_12033,N_12870);
nand UO_204 (O_204,N_12960,N_13050);
nor UO_205 (O_205,N_11519,N_11762);
and UO_206 (O_206,N_12060,N_11679);
nor UO_207 (O_207,N_10487,N_13525);
or UO_208 (O_208,N_12335,N_13529);
nand UO_209 (O_209,N_12696,N_10352);
or UO_210 (O_210,N_14886,N_12863);
or UO_211 (O_211,N_10431,N_12615);
nor UO_212 (O_212,N_11398,N_12267);
or UO_213 (O_213,N_13682,N_11628);
nand UO_214 (O_214,N_12477,N_10913);
and UO_215 (O_215,N_13708,N_11060);
or UO_216 (O_216,N_13554,N_13387);
or UO_217 (O_217,N_13713,N_12508);
nor UO_218 (O_218,N_11930,N_14218);
nor UO_219 (O_219,N_14660,N_14494);
or UO_220 (O_220,N_11304,N_11743);
nand UO_221 (O_221,N_10353,N_14552);
nor UO_222 (O_222,N_12741,N_13562);
or UO_223 (O_223,N_12932,N_10188);
and UO_224 (O_224,N_11513,N_10741);
and UO_225 (O_225,N_14819,N_12806);
nand UO_226 (O_226,N_12061,N_10221);
or UO_227 (O_227,N_10498,N_12975);
or UO_228 (O_228,N_12486,N_13015);
and UO_229 (O_229,N_13564,N_11171);
nor UO_230 (O_230,N_10490,N_12373);
and UO_231 (O_231,N_10764,N_13514);
and UO_232 (O_232,N_13093,N_11802);
or UO_233 (O_233,N_11629,N_12911);
and UO_234 (O_234,N_10709,N_12704);
nand UO_235 (O_235,N_11537,N_11745);
nor UO_236 (O_236,N_10514,N_11917);
nand UO_237 (O_237,N_14388,N_13494);
nand UO_238 (O_238,N_12777,N_10049);
and UO_239 (O_239,N_10361,N_12514);
and UO_240 (O_240,N_10286,N_11299);
nand UO_241 (O_241,N_13940,N_10789);
and UO_242 (O_242,N_13726,N_14748);
or UO_243 (O_243,N_12718,N_13664);
and UO_244 (O_244,N_13432,N_12025);
or UO_245 (O_245,N_12902,N_10871);
nor UO_246 (O_246,N_12661,N_12918);
nor UO_247 (O_247,N_10633,N_13779);
or UO_248 (O_248,N_10842,N_12332);
nand UO_249 (O_249,N_12228,N_12880);
nor UO_250 (O_250,N_10645,N_11234);
nor UO_251 (O_251,N_12976,N_14200);
nand UO_252 (O_252,N_10249,N_13592);
and UO_253 (O_253,N_10969,N_11764);
xor UO_254 (O_254,N_13487,N_14983);
nor UO_255 (O_255,N_14127,N_13908);
and UO_256 (O_256,N_11282,N_11413);
or UO_257 (O_257,N_14281,N_14946);
or UO_258 (O_258,N_13884,N_13977);
or UO_259 (O_259,N_12120,N_14264);
nand UO_260 (O_260,N_13570,N_14456);
nand UO_261 (O_261,N_11533,N_14761);
nor UO_262 (O_262,N_11934,N_10174);
nand UO_263 (O_263,N_10703,N_10419);
nor UO_264 (O_264,N_12881,N_10129);
nor UO_265 (O_265,N_12997,N_11984);
nor UO_266 (O_266,N_11077,N_13663);
and UO_267 (O_267,N_13346,N_10048);
or UO_268 (O_268,N_14283,N_12451);
nor UO_269 (O_269,N_14346,N_14721);
nor UO_270 (O_270,N_10470,N_10491);
nor UO_271 (O_271,N_11657,N_14825);
or UO_272 (O_272,N_11063,N_11437);
or UO_273 (O_273,N_13505,N_12130);
nor UO_274 (O_274,N_11880,N_12411);
nand UO_275 (O_275,N_14701,N_10018);
nor UO_276 (O_276,N_12866,N_10257);
and UO_277 (O_277,N_14569,N_12250);
nand UO_278 (O_278,N_11389,N_11898);
and UO_279 (O_279,N_10694,N_14450);
nand UO_280 (O_280,N_11042,N_14625);
nand UO_281 (O_281,N_13721,N_13149);
or UO_282 (O_282,N_13997,N_12402);
or UO_283 (O_283,N_12834,N_14258);
nor UO_284 (O_284,N_13163,N_11196);
xor UO_285 (O_285,N_14846,N_13565);
and UO_286 (O_286,N_11524,N_10131);
nor UO_287 (O_287,N_10134,N_10122);
nor UO_288 (O_288,N_10551,N_11622);
nor UO_289 (O_289,N_14588,N_13823);
and UO_290 (O_290,N_12784,N_12952);
or UO_291 (O_291,N_11470,N_10692);
and UO_292 (O_292,N_12466,N_14502);
nor UO_293 (O_293,N_11061,N_10831);
or UO_294 (O_294,N_13208,N_14382);
nor UO_295 (O_295,N_10721,N_10879);
and UO_296 (O_296,N_13948,N_13867);
and UO_297 (O_297,N_12494,N_14171);
nor UO_298 (O_298,N_11717,N_14344);
nand UO_299 (O_299,N_14259,N_13216);
nand UO_300 (O_300,N_11431,N_11311);
nand UO_301 (O_301,N_10561,N_13731);
nor UO_302 (O_302,N_12422,N_13256);
and UO_303 (O_303,N_13182,N_12822);
nor UO_304 (O_304,N_14377,N_10837);
nand UO_305 (O_305,N_10477,N_10102);
and UO_306 (O_306,N_10099,N_12664);
or UO_307 (O_307,N_14082,N_11073);
nand UO_308 (O_308,N_13463,N_12263);
nor UO_309 (O_309,N_12172,N_14898);
nor UO_310 (O_310,N_12998,N_13507);
nand UO_311 (O_311,N_13073,N_11955);
nor UO_312 (O_312,N_12389,N_14566);
nor UO_313 (O_313,N_13922,N_14212);
or UO_314 (O_314,N_10412,N_12986);
or UO_315 (O_315,N_12302,N_14410);
and UO_316 (O_316,N_13298,N_13052);
nor UO_317 (O_317,N_12654,N_10881);
nand UO_318 (O_318,N_13645,N_14011);
nand UO_319 (O_319,N_14628,N_12558);
or UO_320 (O_320,N_10450,N_14796);
and UO_321 (O_321,N_12885,N_12971);
or UO_322 (O_322,N_14022,N_14554);
nor UO_323 (O_323,N_13366,N_11394);
or UO_324 (O_324,N_11292,N_12738);
and UO_325 (O_325,N_13576,N_13597);
and UO_326 (O_326,N_13882,N_12889);
nor UO_327 (O_327,N_11911,N_14017);
or UO_328 (O_328,N_11889,N_11062);
nor UO_329 (O_329,N_13760,N_13743);
nand UO_330 (O_330,N_10679,N_14241);
nor UO_331 (O_331,N_14149,N_13627);
and UO_332 (O_332,N_12452,N_13710);
nand UO_333 (O_333,N_10543,N_14828);
xor UO_334 (O_334,N_12780,N_14406);
and UO_335 (O_335,N_10846,N_13247);
or UO_336 (O_336,N_11151,N_10724);
nand UO_337 (O_337,N_14665,N_12487);
nand UO_338 (O_338,N_12417,N_11446);
nand UO_339 (O_339,N_11854,N_14533);
nor UO_340 (O_340,N_14140,N_12645);
or UO_341 (O_341,N_12382,N_12859);
or UO_342 (O_342,N_12089,N_14373);
or UO_343 (O_343,N_11146,N_12955);
and UO_344 (O_344,N_11112,N_11371);
and UO_345 (O_345,N_10340,N_14209);
or UO_346 (O_346,N_12099,N_12166);
nand UO_347 (O_347,N_12893,N_12963);
and UO_348 (O_348,N_11862,N_10628);
nand UO_349 (O_349,N_10512,N_14743);
or UO_350 (O_350,N_14785,N_11637);
nand UO_351 (O_351,N_10172,N_12811);
and UO_352 (O_352,N_10363,N_14633);
and UO_353 (O_353,N_13993,N_13074);
and UO_354 (O_354,N_11627,N_10998);
nor UO_355 (O_355,N_12506,N_11338);
and UO_356 (O_356,N_12418,N_10847);
and UO_357 (O_357,N_12107,N_13276);
and UO_358 (O_358,N_11438,N_12183);
or UO_359 (O_359,N_14490,N_10601);
nand UO_360 (O_360,N_11321,N_10935);
or UO_361 (O_361,N_11465,N_10097);
or UO_362 (O_362,N_13378,N_11835);
and UO_363 (O_363,N_12281,N_10123);
or UO_364 (O_364,N_14401,N_14294);
nor UO_365 (O_365,N_10306,N_14289);
nand UO_366 (O_366,N_12471,N_12515);
nand UO_367 (O_367,N_11009,N_13571);
and UO_368 (O_368,N_10596,N_10273);
or UO_369 (O_369,N_11460,N_10497);
nand UO_370 (O_370,N_11824,N_13880);
nand UO_371 (O_371,N_10891,N_11523);
and UO_372 (O_372,N_13668,N_11783);
or UO_373 (O_373,N_14615,N_13465);
nand UO_374 (O_374,N_13459,N_12243);
and UO_375 (O_375,N_10655,N_13162);
nor UO_376 (O_376,N_14692,N_11123);
nand UO_377 (O_377,N_12603,N_14799);
nor UO_378 (O_378,N_11670,N_11913);
or UO_379 (O_379,N_12816,N_14431);
or UO_380 (O_380,N_13755,N_14412);
and UO_381 (O_381,N_11180,N_11906);
nand UO_382 (O_382,N_12407,N_11541);
nor UO_383 (O_383,N_12016,N_11254);
nand UO_384 (O_384,N_10053,N_14358);
nor UO_385 (O_385,N_12549,N_11444);
or UO_386 (O_386,N_12102,N_13235);
nor UO_387 (O_387,N_11994,N_14836);
and UO_388 (O_388,N_12725,N_14097);
or UO_389 (O_389,N_14371,N_11908);
nand UO_390 (O_390,N_14085,N_14013);
nand UO_391 (O_391,N_12961,N_13952);
nor UO_392 (O_392,N_13382,N_12282);
nand UO_393 (O_393,N_14445,N_10686);
nor UO_394 (O_394,N_12841,N_10147);
nand UO_395 (O_395,N_11324,N_10203);
or UO_396 (O_396,N_11392,N_12609);
and UO_397 (O_397,N_11047,N_14073);
and UO_398 (O_398,N_12585,N_12057);
and UO_399 (O_399,N_11215,N_11309);
and UO_400 (O_400,N_11750,N_10357);
and UO_401 (O_401,N_10008,N_12254);
nand UO_402 (O_402,N_10379,N_13681);
nand UO_403 (O_403,N_11035,N_12193);
or UO_404 (O_404,N_13157,N_12724);
or UO_405 (O_405,N_13446,N_13013);
or UO_406 (O_406,N_12469,N_13342);
nand UO_407 (O_407,N_14069,N_14600);
nor UO_408 (O_408,N_13563,N_12179);
or UO_409 (O_409,N_11018,N_11200);
or UO_410 (O_410,N_10677,N_12734);
nor UO_411 (O_411,N_10209,N_14526);
or UO_412 (O_412,N_13766,N_11618);
nor UO_413 (O_413,N_14481,N_13544);
or UO_414 (O_414,N_14324,N_10162);
nor UO_415 (O_415,N_13858,N_11594);
nand UO_416 (O_416,N_14667,N_11493);
and UO_417 (O_417,N_11977,N_10564);
nor UO_418 (O_418,N_13213,N_11865);
nor UO_419 (O_419,N_12823,N_10687);
nor UO_420 (O_420,N_14263,N_12496);
or UO_421 (O_421,N_11555,N_10917);
and UO_422 (O_422,N_12393,N_13448);
or UO_423 (O_423,N_13702,N_12462);
nand UO_424 (O_424,N_11409,N_12872);
nor UO_425 (O_425,N_10319,N_13040);
and UO_426 (O_426,N_13338,N_12765);
or UO_427 (O_427,N_10591,N_14370);
and UO_428 (O_428,N_14080,N_14782);
or UO_429 (O_429,N_12013,N_10443);
nand UO_430 (O_430,N_13704,N_12219);
nand UO_431 (O_431,N_14973,N_11838);
and UO_432 (O_432,N_12776,N_13316);
nand UO_433 (O_433,N_11344,N_14943);
and UO_434 (O_434,N_10816,N_10783);
nand UO_435 (O_435,N_12737,N_11126);
and UO_436 (O_436,N_14595,N_13331);
and UO_437 (O_437,N_11515,N_10549);
nand UO_438 (O_438,N_10795,N_14860);
nand UO_439 (O_439,N_11333,N_11132);
or UO_440 (O_440,N_12275,N_13491);
nor UO_441 (O_441,N_12305,N_10535);
nand UO_442 (O_442,N_10280,N_11451);
nor UO_443 (O_443,N_12989,N_10976);
or UO_444 (O_444,N_10075,N_13251);
and UO_445 (O_445,N_11167,N_14673);
and UO_446 (O_446,N_12008,N_12604);
nor UO_447 (O_447,N_14389,N_13580);
nor UO_448 (O_448,N_13079,N_13603);
nand UO_449 (O_449,N_10312,N_11342);
nand UO_450 (O_450,N_13436,N_13111);
or UO_451 (O_451,N_12860,N_14181);
or UO_452 (O_452,N_10220,N_14912);
and UO_453 (O_453,N_11191,N_14997);
nand UO_454 (O_454,N_12886,N_10260);
and UO_455 (O_455,N_10817,N_12868);
and UO_456 (O_456,N_11635,N_14580);
nand UO_457 (O_457,N_13841,N_13513);
and UO_458 (O_458,N_13080,N_13613);
or UO_459 (O_459,N_10304,N_14563);
nand UO_460 (O_460,N_13104,N_10571);
nand UO_461 (O_461,N_12326,N_11965);
nand UO_462 (O_462,N_11490,N_13509);
nand UO_463 (O_463,N_11620,N_13812);
nand UO_464 (O_464,N_12084,N_13107);
nand UO_465 (O_465,N_12185,N_13795);
nor UO_466 (O_466,N_11483,N_11904);
and UO_467 (O_467,N_11815,N_11871);
nand UO_468 (O_468,N_14713,N_13835);
nand UO_469 (O_469,N_11467,N_13657);
and UO_470 (O_470,N_13379,N_13177);
or UO_471 (O_471,N_11731,N_10387);
or UO_472 (O_472,N_12261,N_10135);
nand UO_473 (O_473,N_12656,N_10294);
nor UO_474 (O_474,N_13471,N_10113);
or UO_475 (O_475,N_12420,N_10518);
nand UO_476 (O_476,N_12882,N_10865);
nor UO_477 (O_477,N_13976,N_14184);
nor UO_478 (O_478,N_10481,N_13171);
and UO_479 (O_479,N_12491,N_14577);
and UO_480 (O_480,N_11359,N_11631);
nand UO_481 (O_481,N_13411,N_12280);
nor UO_482 (O_482,N_13686,N_10956);
or UO_483 (O_483,N_11578,N_11090);
nor UO_484 (O_484,N_12298,N_12248);
nand UO_485 (O_485,N_11454,N_10723);
or UO_486 (O_486,N_12233,N_14775);
nand UO_487 (O_487,N_10282,N_10300);
nand UO_488 (O_488,N_10921,N_10510);
and UO_489 (O_489,N_12632,N_10887);
and UO_490 (O_490,N_11755,N_11863);
nand UO_491 (O_491,N_11825,N_11380);
or UO_492 (O_492,N_14965,N_12330);
nor UO_493 (O_493,N_12595,N_14112);
nor UO_494 (O_494,N_10963,N_11782);
or UO_495 (O_495,N_12157,N_14207);
nand UO_496 (O_496,N_12802,N_10365);
nand UO_497 (O_497,N_13336,N_13971);
nand UO_498 (O_498,N_13715,N_12761);
and UO_499 (O_499,N_10043,N_13153);
and UO_500 (O_500,N_11587,N_10926);
and UO_501 (O_501,N_14277,N_10767);
nand UO_502 (O_502,N_10944,N_14483);
nor UO_503 (O_503,N_12246,N_12216);
nand UO_504 (O_504,N_10689,N_12094);
and UO_505 (O_505,N_14341,N_11125);
or UO_506 (O_506,N_11726,N_12098);
nor UO_507 (O_507,N_13909,N_10176);
and UO_508 (O_508,N_14252,N_13945);
nand UO_509 (O_509,N_13101,N_10109);
and UO_510 (O_510,N_11597,N_14310);
nor UO_511 (O_511,N_11789,N_12059);
nand UO_512 (O_512,N_13874,N_10572);
or UO_513 (O_513,N_12512,N_10792);
nand UO_514 (O_514,N_13689,N_12377);
or UO_515 (O_515,N_11894,N_12276);
nand UO_516 (O_516,N_11998,N_11030);
and UO_517 (O_517,N_11096,N_10583);
nor UO_518 (O_518,N_11675,N_14586);
and UO_519 (O_519,N_10373,N_11987);
or UO_520 (O_520,N_14248,N_13281);
and UO_521 (O_521,N_11315,N_11066);
nand UO_522 (O_522,N_14253,N_11682);
nor UO_523 (O_523,N_11507,N_12095);
nor UO_524 (O_524,N_11310,N_11369);
nand UO_525 (O_525,N_12790,N_12821);
nor UO_526 (O_526,N_12751,N_11544);
or UO_527 (O_527,N_13160,N_13005);
nand UO_528 (O_528,N_14485,N_11117);
or UO_529 (O_529,N_14808,N_12828);
nor UO_530 (O_530,N_11022,N_10732);
and UO_531 (O_531,N_11518,N_12711);
or UO_532 (O_532,N_11781,N_13764);
or UO_533 (O_533,N_13706,N_11621);
xnor UO_534 (O_534,N_12397,N_10082);
nor UO_535 (O_535,N_14198,N_10955);
and UO_536 (O_536,N_14498,N_12383);
or UO_537 (O_537,N_12812,N_14009);
or UO_538 (O_538,N_12175,N_11793);
nand UO_539 (O_539,N_11417,N_11231);
nand UO_540 (O_540,N_10016,N_10426);
and UO_541 (O_541,N_13732,N_10553);
nand UO_542 (O_542,N_12253,N_10711);
nand UO_543 (O_543,N_11122,N_11411);
or UO_544 (O_544,N_13754,N_10036);
nand UO_545 (O_545,N_11630,N_12223);
or UO_546 (O_546,N_13409,N_12245);
nand UO_547 (O_547,N_10626,N_13662);
or UO_548 (O_548,N_14050,N_13453);
nor UO_549 (O_549,N_10844,N_10284);
or UO_550 (O_550,N_12987,N_10139);
nor UO_551 (O_551,N_14730,N_13280);
and UO_552 (O_552,N_11463,N_12768);
nor UO_553 (O_553,N_13730,N_14786);
nand UO_554 (O_554,N_13059,N_13337);
or UO_555 (O_555,N_14823,N_12526);
nor UO_556 (O_556,N_11382,N_10012);
nor UO_557 (O_557,N_14096,N_14553);
or UO_558 (O_558,N_12981,N_11536);
nand UO_559 (O_559,N_12174,N_10093);
or UO_560 (O_560,N_11345,N_11971);
nand UO_561 (O_561,N_10067,N_10947);
or UO_562 (O_562,N_14234,N_13039);
xnor UO_563 (O_563,N_10667,N_12173);
nor UO_564 (O_564,N_14409,N_13941);
or UO_565 (O_565,N_11432,N_14882);
nor UO_566 (O_566,N_11508,N_10605);
nor UO_567 (O_567,N_13905,N_12907);
and UO_568 (O_568,N_14115,N_13386);
nor UO_569 (O_569,N_10620,N_14845);
and UO_570 (O_570,N_14396,N_14763);
and UO_571 (O_571,N_11288,N_12053);
and UO_572 (O_572,N_14316,N_14732);
and UO_573 (O_573,N_12542,N_12257);
and UO_574 (O_574,N_13838,N_13271);
nand UO_575 (O_575,N_14661,N_14581);
nand UO_576 (O_576,N_14546,N_12347);
and UO_577 (O_577,N_14931,N_13545);
nor UO_578 (O_578,N_11884,N_14697);
and UO_579 (O_579,N_10997,N_12427);
nand UO_580 (O_580,N_14392,N_10781);
or UO_581 (O_581,N_11152,N_12460);
or UO_582 (O_582,N_13868,N_11546);
nand UO_583 (O_583,N_11829,N_12565);
nand UO_584 (O_584,N_14309,N_13913);
nand UO_585 (O_585,N_10945,N_12064);
nor UO_586 (O_586,N_14242,N_14105);
nor UO_587 (O_587,N_13560,N_13590);
and UO_588 (O_588,N_11937,N_13985);
and UO_589 (O_589,N_10625,N_14865);
and UO_590 (O_590,N_14876,N_14851);
and UO_591 (O_591,N_10952,N_10882);
nand UO_592 (O_592,N_14414,N_13426);
and UO_593 (O_593,N_14638,N_10194);
or UO_594 (O_594,N_13367,N_10204);
and UO_595 (O_595,N_11895,N_11876);
and UO_596 (O_596,N_13690,N_10602);
nand UO_597 (O_597,N_13365,N_14522);
nand UO_598 (O_598,N_14535,N_10641);
nand UO_599 (O_599,N_13460,N_12959);
or UO_600 (O_600,N_14376,N_10854);
nor UO_601 (O_601,N_11888,N_14217);
nor UO_602 (O_602,N_11300,N_14384);
or UO_603 (O_603,N_10793,N_11363);
nand UO_604 (O_604,N_12663,N_10555);
or UO_605 (O_605,N_10757,N_14988);
and UO_606 (O_606,N_12307,N_10788);
nor UO_607 (O_607,N_14774,N_14330);
or UO_608 (O_608,N_11833,N_14908);
and UO_609 (O_609,N_10020,N_12212);
and UO_610 (O_610,N_10118,N_12674);
nor UO_611 (O_611,N_13575,N_10640);
nor UO_612 (O_612,N_14157,N_10039);
and UO_613 (O_613,N_11848,N_12082);
and UO_614 (O_614,N_14107,N_10950);
and UO_615 (O_615,N_14053,N_14427);
and UO_616 (O_616,N_10924,N_12345);
and UO_617 (O_617,N_13124,N_10445);
and UO_618 (O_618,N_13953,N_14086);
nand UO_619 (O_619,N_10814,N_11974);
or UO_620 (O_620,N_10245,N_13831);
or UO_621 (O_621,N_14760,N_11262);
nor UO_622 (O_622,N_10144,N_13032);
and UO_623 (O_623,N_14276,N_14245);
and UO_624 (O_624,N_11600,N_12198);
and UO_625 (O_625,N_12559,N_11059);
nand UO_626 (O_626,N_14295,N_11852);
nor UO_627 (O_627,N_12629,N_11615);
or UO_628 (O_628,N_13011,N_12747);
or UO_629 (O_629,N_14594,N_12079);
nand UO_630 (O_630,N_10254,N_12296);
and UO_631 (O_631,N_10405,N_13930);
or UO_632 (O_632,N_14632,N_13914);
and UO_633 (O_633,N_14547,N_10088);
or UO_634 (O_634,N_14194,N_11832);
or UO_635 (O_635,N_14403,N_14254);
nand UO_636 (O_636,N_12056,N_13511);
or UO_637 (O_637,N_10393,N_11267);
or UO_638 (O_638,N_12092,N_12803);
nor UO_639 (O_639,N_10305,N_14320);
or UO_640 (O_640,N_10647,N_13031);
nand UO_641 (O_641,N_14805,N_12808);
nor UO_642 (O_642,N_11853,N_11859);
or UO_643 (O_643,N_10568,N_13441);
xnor UO_644 (O_644,N_10089,N_10971);
and UO_645 (O_645,N_12300,N_13288);
or UO_646 (O_646,N_12111,N_10101);
nand UO_647 (O_647,N_13669,N_13550);
nand UO_648 (O_648,N_12938,N_11864);
nor UO_649 (O_649,N_10408,N_12301);
or UO_650 (O_650,N_14881,N_10446);
or UO_651 (O_651,N_10737,N_12659);
and UO_652 (O_652,N_11734,N_11071);
or UO_653 (O_653,N_13632,N_12232);
nand UO_654 (O_654,N_10167,N_12820);
or UO_655 (O_655,N_14790,N_11901);
nand UO_656 (O_656,N_10580,N_11946);
nor UO_657 (O_657,N_11074,N_10107);
nand UO_658 (O_658,N_13412,N_13685);
nand UO_659 (O_659,N_10907,N_11771);
and UO_660 (O_660,N_11964,N_11372);
and UO_661 (O_661,N_13789,N_10511);
and UO_662 (O_662,N_10676,N_12241);
and UO_663 (O_663,N_12269,N_10086);
nor UO_664 (O_664,N_11704,N_13675);
or UO_665 (O_665,N_12386,N_13626);
nor UO_666 (O_666,N_14271,N_11529);
nor UO_667 (O_667,N_10349,N_14875);
nor UO_668 (O_668,N_14832,N_12753);
nor UO_669 (O_669,N_11186,N_11367);
or UO_670 (O_670,N_14542,N_12314);
nor UO_671 (O_671,N_13806,N_11585);
or UO_672 (O_672,N_13763,N_11678);
nor UO_673 (O_673,N_10484,N_12708);
nand UO_674 (O_674,N_12456,N_13649);
or UO_675 (O_675,N_11811,N_14512);
nand UO_676 (O_676,N_12523,N_13056);
and UO_677 (O_677,N_10964,N_10494);
and UO_678 (O_678,N_11676,N_12745);
nand UO_679 (O_679,N_11773,N_13141);
nand UO_680 (O_680,N_13705,N_11116);
or UO_681 (O_681,N_11305,N_10184);
and UO_682 (O_682,N_10875,N_11706);
nor UO_683 (O_683,N_10243,N_13236);
or UO_684 (O_684,N_14335,N_12927);
nand UO_685 (O_685,N_10988,N_13181);
nand UO_686 (O_686,N_12464,N_13456);
nand UO_687 (O_687,N_13699,N_12824);
or UO_688 (O_688,N_13569,N_13630);
or UO_689 (O_689,N_12238,N_14781);
and UO_690 (O_690,N_10461,N_13756);
or UO_691 (O_691,N_14005,N_14826);
nand UO_692 (O_692,N_11176,N_14123);
and UO_693 (O_693,N_11336,N_12631);
nor UO_694 (O_694,N_13197,N_12641);
nand UO_695 (O_695,N_11253,N_13933);
xnor UO_696 (O_696,N_10136,N_13733);
and UO_697 (O_697,N_12896,N_10278);
and UO_698 (O_698,N_11735,N_12810);
or UO_699 (O_699,N_14185,N_10465);
nor UO_700 (O_700,N_14506,N_13295);
nand UO_701 (O_701,N_10453,N_14286);
and UO_702 (O_702,N_12625,N_12691);
and UO_703 (O_703,N_14919,N_13173);
nand UO_704 (O_704,N_14930,N_11051);
and UO_705 (O_705,N_10733,N_12484);
nor UO_706 (O_706,N_12537,N_10768);
nand UO_707 (O_707,N_14803,N_14191);
or UO_708 (O_708,N_13998,N_14447);
nand UO_709 (O_709,N_12865,N_12414);
nor UO_710 (O_710,N_11181,N_14399);
or UO_711 (O_711,N_12543,N_11590);
or UO_712 (O_712,N_12207,N_10930);
nor UO_713 (O_713,N_12985,N_11918);
or UO_714 (O_714,N_11158,N_13944);
and UO_715 (O_715,N_13826,N_14345);
nand UO_716 (O_716,N_14419,N_14688);
nand UO_717 (O_717,N_14913,N_10472);
nor UO_718 (O_718,N_12221,N_10290);
nand UO_719 (O_719,N_12485,N_12012);
and UO_720 (O_720,N_12836,N_14379);
nor UO_721 (O_721,N_12972,N_13573);
or UO_722 (O_722,N_11792,N_11416);
and UO_723 (O_723,N_12308,N_11166);
and UO_724 (O_724,N_10648,N_10622);
and UO_725 (O_725,N_14597,N_10941);
nor UO_726 (O_726,N_10064,N_13618);
and UO_727 (O_727,N_14036,N_13134);
or UO_728 (O_728,N_12791,N_13257);
or UO_729 (O_729,N_14971,N_11821);
or UO_730 (O_730,N_11258,N_14952);
and UO_731 (O_731,N_14664,N_13566);
nor UO_732 (O_732,N_12727,N_11108);
nor UO_733 (O_733,N_13915,N_13608);
nand UO_734 (O_734,N_13629,N_13254);
nor UO_735 (O_735,N_10336,N_10180);
or UO_736 (O_736,N_10342,N_10862);
nor UO_737 (O_737,N_10307,N_10507);
nand UO_738 (O_738,N_12855,N_13844);
nand UO_739 (O_739,N_13440,N_14470);
or UO_740 (O_740,N_10504,N_14278);
or UO_741 (O_741,N_14429,N_11696);
or UO_742 (O_742,N_11439,N_12122);
and UO_743 (O_743,N_11655,N_12967);
and UO_744 (O_744,N_11102,N_12717);
or UO_745 (O_745,N_10372,N_13292);
and UO_746 (O_746,N_12775,N_12341);
and UO_747 (O_747,N_10874,N_14029);
or UO_748 (O_748,N_11354,N_12353);
and UO_749 (O_749,N_13883,N_10375);
nand UO_750 (O_750,N_12845,N_12399);
and UO_751 (O_751,N_10121,N_13464);
nand UO_752 (O_752,N_14837,N_13278);
nand UO_753 (O_753,N_13522,N_12169);
or UO_754 (O_754,N_12853,N_14020);
nand UO_755 (O_755,N_11319,N_14404);
nand UO_756 (O_756,N_14203,N_12070);
nor UO_757 (O_757,N_12217,N_10228);
nand UO_758 (O_758,N_12381,N_12334);
nand UO_759 (O_759,N_11775,N_13109);
or UO_760 (O_760,N_14962,N_14368);
or UO_761 (O_761,N_11851,N_14319);
or UO_762 (O_762,N_14655,N_14000);
and UO_763 (O_763,N_11275,N_14703);
nand UO_764 (O_764,N_13739,N_13495);
nand UO_765 (O_765,N_10821,N_11020);
or UO_766 (O_766,N_13445,N_10909);
nor UO_767 (O_767,N_11397,N_11421);
nand UO_768 (O_768,N_14896,N_12093);
or UO_769 (O_769,N_12699,N_12188);
nor UO_770 (O_770,N_12778,N_10607);
nand UO_771 (O_771,N_11129,N_12167);
or UO_772 (O_772,N_12141,N_10575);
and UO_773 (O_773,N_10524,N_13327);
and UO_774 (O_774,N_11224,N_13016);
or UO_775 (O_775,N_12758,N_10922);
nor UO_776 (O_776,N_10321,N_10427);
nor UO_777 (O_777,N_12081,N_10414);
nand UO_778 (O_778,N_11244,N_10742);
nand UO_779 (O_779,N_12042,N_13792);
nor UO_780 (O_780,N_13875,N_10975);
nand UO_781 (O_781,N_12020,N_12627);
and UO_782 (O_782,N_12589,N_14398);
nand UO_783 (O_783,N_13008,N_13753);
nand UO_784 (O_784,N_13805,N_11093);
nand UO_785 (O_785,N_13989,N_10295);
nor UO_786 (O_786,N_11660,N_10566);
and UO_787 (O_787,N_14090,N_14056);
nor UO_788 (O_788,N_12290,N_13019);
nand UO_789 (O_789,N_11149,N_13273);
or UO_790 (O_790,N_14274,N_10508);
and UO_791 (O_791,N_11885,N_11070);
nand UO_792 (O_792,N_10636,N_11243);
and UO_793 (O_793,N_12797,N_14857);
nand UO_794 (O_794,N_10884,N_12436);
nor UO_795 (O_795,N_10074,N_12668);
and UO_796 (O_796,N_12848,N_12483);
and UO_797 (O_797,N_10702,N_11187);
or UO_798 (O_798,N_10388,N_12694);
or UO_799 (O_799,N_13775,N_12447);
and UO_800 (O_800,N_13264,N_14887);
or UO_801 (O_801,N_13279,N_12687);
nand UO_802 (O_802,N_13879,N_13200);
or UO_803 (O_803,N_14418,N_10348);
nand UO_804 (O_804,N_10534,N_12346);
nor UO_805 (O_805,N_12990,N_12165);
nand UO_806 (O_806,N_14113,N_11378);
and UO_807 (O_807,N_11883,N_13489);
or UO_808 (O_808,N_13362,N_14922);
nand UO_809 (O_809,N_14350,N_12676);
or UO_810 (O_810,N_13588,N_11956);
or UO_811 (O_811,N_12613,N_10247);
or UO_812 (O_812,N_10251,N_12320);
nand UO_813 (O_813,N_13828,N_11820);
nand UO_814 (O_814,N_14102,N_10462);
nand UO_815 (O_815,N_13259,N_14288);
nor UO_816 (O_816,N_13421,N_10360);
or UO_817 (O_817,N_12475,N_14590);
and UO_818 (O_818,N_12533,N_10684);
nand UO_819 (O_819,N_10428,N_14163);
or UO_820 (O_820,N_13694,N_14416);
nand UO_821 (O_821,N_10186,N_12922);
nor UO_822 (O_822,N_12450,N_14734);
nor UO_823 (O_823,N_14187,N_10669);
and UO_824 (O_824,N_11506,N_10157);
or UO_825 (O_825,N_14202,N_11040);
nor UO_826 (O_826,N_11023,N_13226);
and UO_827 (O_827,N_14567,N_14121);
nor UO_828 (O_828,N_11645,N_12408);
or UO_829 (O_829,N_14100,N_12540);
and UO_830 (O_830,N_14618,N_12109);
nand UO_831 (O_831,N_13658,N_14934);
nor UO_832 (O_832,N_10731,N_13122);
and UO_833 (O_833,N_14044,N_11535);
nand UO_834 (O_834,N_10656,N_14176);
or UO_835 (O_835,N_11156,N_11160);
nor UO_836 (O_836,N_12003,N_12560);
and UO_837 (O_837,N_14969,N_12647);
nor UO_838 (O_838,N_13116,N_11443);
and UO_839 (O_839,N_13719,N_10371);
and UO_840 (O_840,N_12392,N_10246);
nor UO_841 (O_841,N_14463,N_13548);
and UO_842 (O_842,N_11351,N_12618);
or UO_843 (O_843,N_13816,N_13615);
nor UO_844 (O_844,N_14422,N_10652);
and UO_845 (O_845,N_13321,N_14441);
nand UO_846 (O_846,N_12178,N_13593);
and UO_847 (O_847,N_13431,N_14822);
nand UO_848 (O_848,N_11698,N_14981);
and UO_849 (O_849,N_12391,N_13286);
and UO_850 (O_850,N_10070,N_10786);
nor UO_851 (O_851,N_12028,N_13781);
nand UO_852 (O_852,N_10713,N_11613);
nor UO_853 (O_853,N_14479,N_11945);
nor UO_854 (O_854,N_14466,N_11099);
nand UO_855 (O_855,N_14970,N_14866);
nor UO_856 (O_856,N_14830,N_12037);
nor UO_857 (O_857,N_13473,N_10191);
nor UO_858 (O_858,N_14848,N_10780);
and UO_859 (O_859,N_10646,N_10747);
nand UO_860 (O_860,N_14126,N_11842);
and UO_861 (O_861,N_13496,N_11512);
nand UO_862 (O_862,N_11114,N_12200);
nor UO_863 (O_863,N_10755,N_12349);
nand UO_864 (O_864,N_14605,N_14476);
nand UO_865 (O_865,N_10738,N_13811);
and UO_866 (O_866,N_13245,N_14669);
and UO_867 (O_867,N_11900,N_13150);
or UO_868 (O_868,N_14706,N_10859);
or UO_869 (O_869,N_14996,N_13845);
nand UO_870 (O_870,N_10991,N_14679);
or UO_871 (O_871,N_12591,N_14809);
and UO_872 (O_872,N_14749,N_13023);
nand UO_873 (O_873,N_11286,N_13285);
nor UO_874 (O_874,N_12370,N_14745);
or UO_875 (O_875,N_11449,N_13077);
nor UO_876 (O_876,N_13889,N_10597);
nand UO_877 (O_877,N_10076,N_13364);
nand UO_878 (O_878,N_10447,N_12069);
nand UO_879 (O_879,N_13991,N_14145);
nand UO_880 (O_880,N_13503,N_11008);
or UO_881 (O_881,N_13345,N_14031);
nand UO_882 (O_882,N_12009,N_10314);
and UO_883 (O_883,N_14708,N_12369);
and UO_884 (O_884,N_12256,N_12240);
nand UO_885 (O_885,N_10858,N_13022);
nand UO_886 (O_886,N_14003,N_14173);
and UO_887 (O_887,N_11335,N_12168);
nor UO_888 (O_888,N_10739,N_14351);
and UO_889 (O_889,N_10383,N_10612);
nand UO_890 (O_890,N_11225,N_13589);
and UO_891 (O_891,N_10823,N_10271);
nor UO_892 (O_892,N_12356,N_12572);
and UO_893 (O_893,N_12505,N_12544);
or UO_894 (O_894,N_14391,N_10420);
or UO_895 (O_895,N_11105,N_12497);
or UO_896 (O_896,N_10025,N_10451);
nor UO_897 (O_897,N_10301,N_11572);
nand UO_898 (O_898,N_12049,N_13371);
nor UO_899 (O_899,N_11796,N_12814);
nand UO_900 (O_900,N_11276,N_11957);
nor UO_901 (O_901,N_14239,N_11738);
and UO_902 (O_902,N_11038,N_14839);
and UO_903 (O_903,N_10554,N_14804);
nand UO_904 (O_904,N_11150,N_13036);
and UO_905 (O_905,N_10397,N_11415);
or UO_906 (O_906,N_14844,N_11203);
and UO_907 (O_907,N_11779,N_12562);
or UO_908 (O_908,N_13921,N_14304);
or UO_909 (O_909,N_10992,N_12830);
and UO_910 (O_910,N_11999,N_11691);
nand UO_911 (O_911,N_12712,N_11287);
and UO_912 (O_912,N_13067,N_14523);
or UO_913 (O_913,N_11744,N_11100);
and UO_914 (O_914,N_14647,N_12550);
and UO_915 (O_915,N_13524,N_13862);
and UO_916 (O_916,N_13186,N_10760);
and UO_917 (O_917,N_12265,N_12612);
and UO_918 (O_918,N_11837,N_11261);
or UO_919 (O_919,N_13060,N_12423);
nand UO_920 (O_920,N_10513,N_11752);
nand UO_921 (O_921,N_10981,N_11646);
nor UO_922 (O_922,N_10632,N_13510);
nand UO_923 (O_923,N_12726,N_14682);
xnor UO_924 (O_924,N_14439,N_12781);
nand UO_925 (O_925,N_10272,N_11666);
or UO_926 (O_926,N_13302,N_14047);
or UO_927 (O_927,N_13119,N_11935);
nor UO_928 (O_928,N_14402,N_12313);
and UO_929 (O_929,N_11365,N_11222);
and UO_930 (O_930,N_14657,N_12137);
nor UO_931 (O_931,N_11983,N_10374);
nor UO_932 (O_932,N_13033,N_14675);
nor UO_933 (O_933,N_13395,N_10505);
or UO_934 (O_934,N_14920,N_12213);
nand UO_935 (O_935,N_11356,N_13678);
and UO_936 (O_936,N_12103,N_11144);
nor UO_937 (O_937,N_10866,N_12262);
or UO_938 (O_938,N_12914,N_14075);
or UO_939 (O_939,N_11131,N_14153);
nor UO_940 (O_940,N_10448,N_12129);
nor UO_941 (O_941,N_13856,N_11858);
or UO_942 (O_942,N_13258,N_12363);
nand UO_943 (O_943,N_12038,N_12638);
nor UO_944 (O_944,N_12974,N_10335);
nor UO_945 (O_945,N_14656,N_14899);
nand UO_946 (O_946,N_13918,N_14759);
or UO_947 (O_947,N_14991,N_13054);
and UO_948 (O_948,N_12570,N_13852);
or UO_949 (O_949,N_14771,N_12988);
nand UO_950 (O_950,N_12709,N_13152);
and UO_951 (O_951,N_11462,N_11668);
nor UO_952 (O_952,N_11103,N_10464);
nor UO_953 (O_953,N_10007,N_13824);
and UO_954 (O_954,N_14645,N_10722);
and UO_955 (O_955,N_11887,N_11043);
and UO_956 (O_956,N_10119,N_10163);
nor UO_957 (O_957,N_11237,N_10369);
or UO_958 (O_958,N_11740,N_10649);
nand UO_959 (O_959,N_12877,N_12088);
and UO_960 (O_960,N_11936,N_13986);
nor UO_961 (O_961,N_12671,N_10631);
and UO_962 (O_962,N_13846,N_10310);
and UO_963 (O_963,N_14624,N_10046);
nand UO_964 (O_964,N_14895,N_12576);
nor UO_965 (O_965,N_14630,N_11142);
or UO_966 (O_966,N_10068,N_14635);
and UO_967 (O_967,N_11663,N_13340);
and UO_968 (O_968,N_13322,N_14611);
nor UO_969 (O_969,N_11348,N_10889);
nand UO_970 (O_970,N_11772,N_10654);
or UO_971 (O_971,N_11791,N_14070);
and UO_972 (O_972,N_11905,N_13897);
nor UO_973 (O_973,N_13420,N_13350);
and UO_974 (O_974,N_13239,N_12343);
or UO_975 (O_975,N_10225,N_13318);
and UO_976 (O_976,N_11632,N_10219);
nand UO_977 (O_977,N_11733,N_11826);
or UO_978 (O_978,N_14634,N_10666);
nand UO_979 (O_979,N_12513,N_14674);
and UO_980 (O_980,N_14446,N_11478);
and UO_981 (O_981,N_12571,N_10143);
and UO_982 (O_982,N_14921,N_13368);
nand UO_983 (O_983,N_11701,N_11845);
and UO_984 (O_984,N_14613,N_11521);
nor UO_985 (O_985,N_13574,N_11279);
and UO_986 (O_986,N_12639,N_12443);
or UO_987 (O_987,N_10993,N_10750);
and UO_988 (O_988,N_11530,N_11135);
nor UO_989 (O_989,N_13966,N_14462);
xnor UO_990 (O_990,N_12563,N_14491);
and UO_991 (O_991,N_12968,N_11714);
nand UO_992 (O_992,N_11297,N_13549);
nor UO_993 (O_993,N_10062,N_12910);
and UO_994 (O_994,N_14568,N_12651);
or UO_995 (O_995,N_13652,N_14180);
nor UO_996 (O_996,N_12043,N_11727);
nor UO_997 (O_997,N_11407,N_13521);
and UO_998 (O_998,N_13504,N_10619);
nor UO_999 (O_999,N_10562,N_10525);
nor UO_1000 (O_1000,N_10717,N_12701);
or UO_1001 (O_1001,N_12002,N_13193);
or UO_1002 (O_1002,N_11314,N_12316);
and UO_1003 (O_1003,N_14603,N_13762);
nand UO_1004 (O_1004,N_11992,N_10486);
nand UO_1005 (O_1005,N_11128,N_11002);
nand UO_1006 (O_1006,N_13045,N_13771);
nand UO_1007 (O_1007,N_10806,N_14363);
and UO_1008 (O_1008,N_10942,N_12851);
nand UO_1009 (O_1009,N_10090,N_11313);
or UO_1010 (O_1010,N_12579,N_10804);
or UO_1011 (O_1011,N_10683,N_10759);
and UO_1012 (O_1012,N_13616,N_14489);
and UO_1013 (O_1013,N_11159,N_12833);
nor UO_1014 (O_1014,N_14321,N_12351);
and UO_1015 (O_1015,N_14914,N_11430);
or UO_1016 (O_1016,N_14838,N_12991);
or UO_1017 (O_1017,N_10411,N_12191);
or UO_1018 (O_1018,N_11808,N_11814);
nor UO_1019 (O_1019,N_13132,N_11509);
and UO_1020 (O_1020,N_14131,N_14452);
nor UO_1021 (O_1021,N_12658,N_12278);
or UO_1022 (O_1022,N_11370,N_12683);
or UO_1023 (O_1023,N_12412,N_12628);
nor UO_1024 (O_1024,N_14948,N_10538);
and UO_1025 (O_1025,N_14918,N_12176);
and UO_1026 (O_1026,N_10966,N_14861);
or UO_1027 (O_1027,N_14142,N_13335);
nand UO_1028 (O_1028,N_10496,N_10878);
nor UO_1029 (O_1029,N_14408,N_10418);
and UO_1030 (O_1030,N_14021,N_14561);
nand UO_1031 (O_1031,N_14723,N_11756);
nor UO_1032 (O_1032,N_10480,N_10252);
nand UO_1033 (O_1033,N_11019,N_14672);
or UO_1034 (O_1034,N_14074,N_11328);
or UO_1035 (O_1035,N_13746,N_13185);
and UO_1036 (O_1036,N_10281,N_10813);
nand UO_1037 (O_1037,N_13787,N_14385);
or UO_1038 (O_1038,N_13120,N_14905);
nand UO_1039 (O_1039,N_10841,N_14987);
and UO_1040 (O_1040,N_12119,N_13878);
and UO_1041 (O_1041,N_14356,N_11143);
nor UO_1042 (O_1042,N_13218,N_10227);
nand UO_1043 (O_1043,N_12468,N_14357);
xnor UO_1044 (O_1044,N_11823,N_11395);
or UO_1045 (O_1045,N_14507,N_13798);
nor UO_1046 (O_1046,N_14720,N_11985);
nand UO_1047 (O_1047,N_10213,N_10933);
nand UO_1048 (O_1048,N_11643,N_11036);
and UO_1049 (O_1049,N_14197,N_12361);
nor UO_1050 (O_1050,N_11564,N_11500);
nand UO_1051 (O_1051,N_11959,N_14654);
and UO_1052 (O_1052,N_13375,N_11174);
or UO_1053 (O_1053,N_14451,N_12921);
and UO_1054 (O_1054,N_13404,N_12255);
nor UO_1055 (O_1055,N_14811,N_12568);
and UO_1056 (O_1056,N_11303,N_14870);
nor UO_1057 (O_1057,N_10864,N_14953);
or UO_1058 (O_1058,N_11777,N_10995);
nand UO_1059 (O_1059,N_14813,N_14864);
or UO_1060 (O_1060,N_14663,N_14440);
nand UO_1061 (O_1061,N_11649,N_11154);
or UO_1062 (O_1062,N_11239,N_11334);
and UO_1063 (O_1063,N_10539,N_11147);
or UO_1064 (O_1064,N_11877,N_13803);
nand UO_1065 (O_1065,N_10704,N_10230);
and UO_1066 (O_1066,N_14099,N_11768);
and UO_1067 (O_1067,N_14428,N_14609);
and UO_1068 (O_1068,N_11923,N_14034);
nand UO_1069 (O_1069,N_11075,N_12873);
or UO_1070 (O_1070,N_11798,N_10799);
nand UO_1071 (O_1071,N_14753,N_12380);
nand UO_1072 (O_1072,N_13354,N_14303);
xnor UO_1073 (O_1073,N_10103,N_13659);
and UO_1074 (O_1074,N_10610,N_11291);
nor UO_1075 (O_1075,N_10744,N_14814);
and UO_1076 (O_1076,N_12083,N_12626);
or UO_1077 (O_1077,N_14947,N_14023);
nor UO_1078 (O_1078,N_10211,N_14019);
or UO_1079 (O_1079,N_13427,N_12144);
nor UO_1080 (O_1080,N_14904,N_10503);
nand UO_1081 (O_1081,N_11861,N_14602);
nand UO_1082 (O_1082,N_10288,N_14130);
or UO_1083 (O_1083,N_11403,N_13165);
nand UO_1084 (O_1084,N_13154,N_10769);
or UO_1085 (O_1085,N_10044,N_13808);
or UO_1086 (O_1086,N_14599,N_11769);
nor UO_1087 (O_1087,N_14048,N_10132);
or UO_1088 (O_1088,N_12548,N_12966);
and UO_1089 (O_1089,N_12949,N_11347);
nor UO_1090 (O_1090,N_13466,N_13490);
nor UO_1091 (O_1091,N_10745,N_14517);
and UO_1092 (O_1092,N_14833,N_12546);
nor UO_1093 (O_1093,N_14161,N_12323);
and UO_1094 (O_1094,N_12681,N_12620);
nor UO_1095 (O_1095,N_12716,N_14550);
or UO_1096 (O_1096,N_11611,N_10673);
nand UO_1097 (O_1097,N_11197,N_10479);
xor UO_1098 (O_1098,N_12601,N_10544);
nand UO_1099 (O_1099,N_12982,N_11434);
or UO_1100 (O_1100,N_12317,N_11041);
and UO_1101 (O_1101,N_14700,N_14224);
nand UO_1102 (O_1102,N_13888,N_10912);
or UO_1103 (O_1103,N_12446,N_10634);
nand UO_1104 (O_1104,N_10699,N_10754);
nor UO_1105 (O_1105,N_12536,N_11525);
and UO_1106 (O_1106,N_13822,N_13533);
or UO_1107 (O_1107,N_11625,N_12970);
and UO_1108 (O_1108,N_14146,N_12964);
and UO_1109 (O_1109,N_13907,N_12667);
or UO_1110 (O_1110,N_14033,N_13847);
nand UO_1111 (O_1111,N_12161,N_10547);
or UO_1112 (O_1112,N_11050,N_14190);
or UO_1113 (O_1113,N_12145,N_13105);
nand UO_1114 (O_1114,N_11428,N_13737);
and UO_1115 (O_1115,N_10351,N_13268);
nor UO_1116 (O_1116,N_14686,N_11703);
nand UO_1117 (O_1117,N_14394,N_13047);
or UO_1118 (O_1118,N_11387,N_13738);
nor UO_1119 (O_1119,N_14251,N_12891);
nand UO_1120 (O_1120,N_12879,N_10526);
and UO_1121 (O_1121,N_10401,N_12457);
or UO_1122 (O_1122,N_11273,N_13747);
nand UO_1123 (O_1123,N_13861,N_12689);
or UO_1124 (O_1124,N_14247,N_11510);
and UO_1125 (O_1125,N_12396,N_11711);
and UO_1126 (O_1126,N_14035,N_14642);
nor UO_1127 (O_1127,N_13091,N_14778);
nand UO_1128 (O_1128,N_11376,N_11795);
or UO_1129 (O_1129,N_12406,N_14272);
nor UO_1130 (O_1130,N_11165,N_14095);
and UO_1131 (O_1131,N_14280,N_13179);
nor UO_1132 (O_1132,N_13347,N_12433);
or UO_1133 (O_1133,N_12480,N_14961);
or UO_1134 (O_1134,N_12920,N_12495);
nor UO_1135 (O_1135,N_11264,N_12733);
and UO_1136 (O_1136,N_10459,N_14231);
nor UO_1137 (O_1137,N_14765,N_13783);
nand UO_1138 (O_1138,N_11001,N_10277);
or UO_1139 (O_1139,N_10111,N_13376);
and UO_1140 (O_1140,N_11179,N_14015);
nor UO_1141 (O_1141,N_12713,N_13146);
nand UO_1142 (O_1142,N_13439,N_12831);
or UO_1143 (O_1143,N_13636,N_13919);
or UO_1144 (O_1144,N_13405,N_11442);
and UO_1145 (O_1145,N_12686,N_11175);
nor UO_1146 (O_1146,N_13187,N_13640);
and UO_1147 (O_1147,N_12962,N_13126);
or UO_1148 (O_1148,N_10905,N_13903);
nand UO_1149 (O_1149,N_13419,N_12826);
and UO_1150 (O_1150,N_14659,N_12430);
or UO_1151 (O_1151,N_14925,N_13572);
and UO_1152 (O_1152,N_13729,N_10822);
and UO_1153 (O_1153,N_11920,N_13871);
xnor UO_1154 (O_1154,N_12472,N_10034);
or UO_1155 (O_1155,N_11423,N_13483);
nand UO_1156 (O_1156,N_13425,N_13559);
nor UO_1157 (O_1157,N_13942,N_14582);
or UO_1158 (O_1158,N_13557,N_11910);
nor UO_1159 (O_1159,N_11661,N_12688);
and UO_1160 (O_1160,N_14313,N_12004);
or UO_1161 (O_1161,N_10234,N_12782);
or UO_1162 (O_1162,N_14054,N_14484);
or UO_1163 (O_1163,N_14539,N_10208);
nand UO_1164 (O_1164,N_14780,N_12587);
or UO_1165 (O_1165,N_12371,N_11375);
and UO_1166 (O_1166,N_10948,N_12292);
nor UO_1167 (O_1167,N_13188,N_14359);
nand UO_1168 (O_1168,N_10545,N_13130);
or UO_1169 (O_1169,N_11058,N_14696);
and UO_1170 (O_1170,N_11979,N_13144);
nand UO_1171 (O_1171,N_13314,N_14442);
nor UO_1172 (O_1172,N_10579,N_10784);
nor UO_1173 (O_1173,N_10567,N_14972);
nor UO_1174 (O_1174,N_10327,N_11966);
or UO_1175 (O_1175,N_13770,N_12752);
nand UO_1176 (O_1176,N_10714,N_10515);
nor UO_1177 (O_1177,N_12026,N_14584);
or UO_1178 (O_1178,N_13975,N_13499);
nor UO_1179 (O_1179,N_10590,N_12425);
nand UO_1180 (O_1180,N_12856,N_10087);
and UO_1181 (O_1181,N_11241,N_12735);
nand UO_1182 (O_1182,N_10094,N_11183);
nor UO_1183 (O_1183,N_14482,N_10302);
nand UO_1184 (O_1184,N_11065,N_14862);
and UO_1185 (O_1185,N_13424,N_11331);
nor UO_1186 (O_1186,N_14237,N_14226);
or UO_1187 (O_1187,N_11294,N_14843);
or UO_1188 (O_1188,N_13620,N_11584);
nor UO_1189 (O_1189,N_12101,N_12903);
nand UO_1190 (O_1190,N_14165,N_12375);
nor UO_1191 (O_1191,N_13076,N_10128);
nor UO_1192 (O_1192,N_11571,N_10552);
and UO_1193 (O_1193,N_12771,N_11715);
nor UO_1194 (O_1194,N_11697,N_11556);
nor UO_1195 (O_1195,N_13534,N_10743);
nand UO_1196 (O_1196,N_13191,N_13553);
and UO_1197 (O_1197,N_10506,N_14508);
nand UO_1198 (O_1198,N_13328,N_11306);
nor UO_1199 (O_1199,N_12600,N_10285);
and UO_1200 (O_1200,N_11185,N_13745);
or UO_1201 (O_1201,N_10444,N_14397);
and UO_1202 (O_1202,N_12331,N_12220);
or UO_1203 (O_1203,N_10557,N_11339);
nor UO_1204 (O_1204,N_14644,N_13996);
nand UO_1205 (O_1205,N_13004,N_14916);
nand UO_1206 (O_1206,N_11776,N_13894);
or UO_1207 (O_1207,N_13638,N_13249);
nand UO_1208 (O_1208,N_10537,N_10391);
nor UO_1209 (O_1209,N_10796,N_10060);
nand UO_1210 (O_1210,N_10698,N_10421);
nor UO_1211 (O_1211,N_10037,N_11327);
nor UO_1212 (O_1212,N_11440,N_11976);
and UO_1213 (O_1213,N_13584,N_12979);
nand UO_1214 (O_1214,N_13438,N_10356);
or UO_1215 (O_1215,N_11127,N_11709);
or UO_1216 (O_1216,N_14636,N_11607);
nor UO_1217 (O_1217,N_11867,N_10377);
and UO_1218 (O_1218,N_10398,N_12388);
or UO_1219 (O_1219,N_14847,N_14134);
nand UO_1220 (O_1220,N_12635,N_11212);
and UO_1221 (O_1221,N_13000,N_14728);
or UO_1222 (O_1222,N_14727,N_14878);
and UO_1223 (O_1223,N_10259,N_13660);
nor UO_1224 (O_1224,N_10925,N_12121);
nand UO_1225 (O_1225,N_11349,N_14329);
nand UO_1226 (O_1226,N_14741,N_14718);
or UO_1227 (O_1227,N_13317,N_14712);
and UO_1228 (O_1228,N_11566,N_10303);
nor UO_1229 (O_1229,N_10961,N_14980);
nor UO_1230 (O_1230,N_13917,N_10530);
and UO_1231 (O_1231,N_10263,N_10084);
and UO_1232 (O_1232,N_11565,N_14269);
nor UO_1233 (O_1233,N_11652,N_12076);
nand UO_1234 (O_1234,N_12730,N_11931);
nor UO_1235 (O_1235,N_12901,N_10587);
nand UO_1236 (O_1236,N_12235,N_14300);
nand UO_1237 (O_1237,N_10805,N_14111);
nand UO_1238 (O_1238,N_10127,N_14355);
nor UO_1239 (O_1239,N_10495,N_12352);
nand UO_1240 (O_1240,N_10345,N_14042);
nand UO_1241 (O_1241,N_13289,N_14940);
or UO_1242 (O_1242,N_14742,N_13757);
nor UO_1243 (O_1243,N_11110,N_10385);
nand UO_1244 (O_1244,N_13890,N_11765);
nand UO_1245 (O_1245,N_12285,N_13958);
or UO_1246 (O_1246,N_12905,N_14670);
nand UO_1247 (O_1247,N_12387,N_11708);
nor UO_1248 (O_1248,N_11010,N_13943);
nand UO_1249 (O_1249,N_14435,N_10868);
and UO_1250 (O_1250,N_14469,N_11658);
nand UO_1251 (O_1251,N_14888,N_11366);
nand UO_1252 (O_1252,N_10815,N_13100);
or UO_1253 (O_1253,N_10283,N_14162);
or UO_1254 (O_1254,N_10790,N_10297);
nand UO_1255 (O_1255,N_10836,N_14332);
or UO_1256 (O_1256,N_11406,N_10151);
and UO_1257 (O_1257,N_11881,N_12018);
and UO_1258 (O_1258,N_11803,N_10027);
nor UO_1259 (O_1259,N_13772,N_12710);
nand UO_1260 (O_1260,N_14430,N_10869);
xnor UO_1261 (O_1261,N_10644,N_10962);
nand UO_1262 (O_1262,N_12288,N_14699);
or UO_1263 (O_1263,N_10173,N_10079);
or UO_1264 (O_1264,N_14027,N_13969);
nor UO_1265 (O_1265,N_14564,N_10965);
and UO_1266 (O_1266,N_11169,N_11656);
nand UO_1267 (O_1267,N_10328,N_13954);
and UO_1268 (O_1268,N_13069,N_10071);
and UO_1269 (O_1269,N_11933,N_14935);
nand UO_1270 (O_1270,N_13750,N_10706);
nand UO_1271 (O_1271,N_12206,N_14910);
and UO_1272 (O_1272,N_14206,N_10115);
or UO_1273 (O_1273,N_13444,N_14318);
nand UO_1274 (O_1274,N_13692,N_10206);
or UO_1275 (O_1275,N_14687,N_12624);
nand UO_1276 (O_1276,N_10040,N_14284);
and UO_1277 (O_1277,N_13671,N_11856);
nand UO_1278 (O_1278,N_12134,N_13380);
and UO_1279 (O_1279,N_14606,N_10827);
and UO_1280 (O_1280,N_11623,N_12759);
nand UO_1281 (O_1281,N_11596,N_10331);
and UO_1282 (O_1282,N_11551,N_13057);
nor UO_1283 (O_1283,N_11256,N_13399);
or UO_1284 (O_1284,N_14957,N_11879);
nand UO_1285 (O_1285,N_14333,N_10031);
xor UO_1286 (O_1286,N_10523,N_10005);
nand UO_1287 (O_1287,N_10137,N_10600);
nand UO_1288 (O_1288,N_13999,N_11408);
and UO_1289 (O_1289,N_14079,N_12861);
or UO_1290 (O_1290,N_14110,N_13628);
or UO_1291 (O_1291,N_14238,N_11830);
nand UO_1292 (O_1292,N_12139,N_11849);
and UO_1293 (O_1293,N_14477,N_11098);
nand UO_1294 (O_1294,N_13683,N_11581);
nor UO_1295 (O_1295,N_10972,N_12695);
and UO_1296 (O_1296,N_13284,N_13458);
and UO_1297 (O_1297,N_12519,N_13818);
and UO_1298 (O_1298,N_11816,N_13241);
and UO_1299 (O_1299,N_13416,N_12010);
xnor UO_1300 (O_1300,N_13895,N_11240);
nor UO_1301 (O_1301,N_11317,N_12535);
or UO_1302 (O_1302,N_14071,N_14978);
or UO_1303 (O_1303,N_11651,N_12000);
and UO_1304 (O_1304,N_10586,N_13530);
or UO_1305 (O_1305,N_10073,N_14758);
nor UO_1306 (O_1306,N_10395,N_14496);
nor UO_1307 (O_1307,N_12394,N_11497);
and UO_1308 (O_1308,N_14210,N_10700);
nor UO_1309 (O_1309,N_12524,N_12091);
or UO_1310 (O_1310,N_10996,N_13709);
nor UO_1311 (O_1311,N_12441,N_11195);
nor UO_1312 (O_1312,N_11377,N_12531);
or UO_1313 (O_1313,N_11280,N_13881);
nand UO_1314 (O_1314,N_10430,N_10072);
and UO_1315 (O_1315,N_14092,N_13639);
and UO_1316 (O_1316,N_12465,N_12919);
and UO_1317 (O_1317,N_11886,N_13204);
nand UO_1318 (O_1318,N_11120,N_12819);
nand UO_1319 (O_1319,N_14268,N_12622);
nand UO_1320 (O_1320,N_11942,N_14492);
and UO_1321 (O_1321,N_13407,N_14094);
nand UO_1322 (O_1322,N_13972,N_13595);
xnor UO_1323 (O_1323,N_14872,N_11271);
or UO_1324 (O_1324,N_14829,N_10359);
nor UO_1325 (O_1325,N_11385,N_13297);
and UO_1326 (O_1326,N_11872,N_13117);
and UO_1327 (O_1327,N_11504,N_11659);
and UO_1328 (O_1328,N_13646,N_14315);
and UO_1329 (O_1329,N_13714,N_12135);
nand UO_1330 (O_1330,N_14938,N_12459);
nor UO_1331 (O_1331,N_12432,N_12054);
or UO_1332 (O_1332,N_14714,N_12424);
xor UO_1333 (O_1333,N_12398,N_13384);
or UO_1334 (O_1334,N_14155,N_11890);
nand UO_1335 (O_1335,N_11284,N_14014);
nor UO_1336 (O_1336,N_10914,N_10627);
or UO_1337 (O_1337,N_14125,N_13751);
nor UO_1338 (O_1338,N_11617,N_13030);
or UO_1339 (O_1339,N_10190,N_12087);
and UO_1340 (O_1340,N_11648,N_14894);
nor UO_1341 (O_1341,N_13391,N_12805);
and UO_1342 (O_1342,N_11312,N_10727);
nor UO_1343 (O_1343,N_14937,N_11800);
nor UO_1344 (O_1344,N_14168,N_13135);
and UO_1345 (O_1345,N_13648,N_10197);
or UO_1346 (O_1346,N_13774,N_13558);
or UO_1347 (O_1347,N_12453,N_10378);
nor UO_1348 (O_1348,N_11368,N_13979);
and UO_1349 (O_1349,N_10155,N_11766);
nand UO_1350 (O_1350,N_14298,N_11381);
and UO_1351 (O_1351,N_14228,N_10876);
nor UO_1352 (O_1352,N_12171,N_10522);
or UO_1353 (O_1353,N_11178,N_13523);
and UO_1354 (O_1354,N_11013,N_11788);
nand UO_1355 (O_1355,N_10292,N_12342);
and UO_1356 (O_1356,N_11583,N_10269);
or UO_1357 (O_1357,N_11870,N_12528);
and UO_1358 (O_1358,N_11499,N_10594);
nand UO_1359 (O_1359,N_10797,N_10287);
nor UO_1360 (O_1360,N_11316,N_12994);
nor UO_1361 (O_1361,N_10801,N_10017);
or UO_1362 (O_1362,N_10368,N_12593);
and UO_1363 (O_1363,N_13736,N_12983);
and UO_1364 (O_1364,N_13515,N_10045);
nor UO_1365 (O_1365,N_13538,N_10390);
nand UO_1366 (O_1366,N_11694,N_10298);
nand UO_1367 (O_1367,N_13672,N_12525);
nand UO_1368 (O_1368,N_10315,N_10181);
nand UO_1369 (O_1369,N_14949,N_12827);
and UO_1370 (O_1370,N_10756,N_14215);
or UO_1371 (O_1371,N_11926,N_14689);
nand UO_1372 (O_1372,N_12160,N_11599);
or UO_1373 (O_1373,N_11285,N_12788);
and UO_1374 (O_1374,N_11289,N_13403);
nor UO_1375 (O_1375,N_14002,N_13602);
nand UO_1376 (O_1376,N_12566,N_14059);
and UO_1377 (O_1377,N_14108,N_11722);
nand UO_1378 (O_1378,N_14695,N_14222);
or UO_1379 (O_1379,N_13155,N_10309);
nor UO_1380 (O_1380,N_12329,N_12077);
nand UO_1381 (O_1381,N_13158,N_13778);
nor UO_1382 (O_1382,N_11025,N_11847);
or UO_1383 (O_1383,N_12744,N_12706);
nor UO_1384 (O_1384,N_11665,N_10216);
nand UO_1385 (O_1385,N_13330,N_13125);
or UO_1386 (O_1386,N_11068,N_13827);
or UO_1387 (O_1387,N_13674,N_11575);
nor UO_1388 (O_1388,N_13901,N_10604);
nand UO_1389 (O_1389,N_10765,N_10499);
nor UO_1390 (O_1390,N_10166,N_13099);
nor UO_1391 (O_1391,N_10104,N_12474);
nand UO_1392 (O_1392,N_11549,N_12419);
nand UO_1393 (O_1393,N_10150,N_13369);
nor UO_1394 (O_1394,N_10014,N_13728);
nand UO_1395 (O_1395,N_10334,N_10435);
and UO_1396 (O_1396,N_10880,N_12355);
and UO_1397 (O_1397,N_14927,N_14292);
and UO_1398 (O_1398,N_12825,N_12792);
or UO_1399 (O_1399,N_12030,N_12883);
or UO_1400 (O_1400,N_12529,N_14867);
xnor UO_1401 (O_1401,N_13293,N_13633);
nor UO_1402 (O_1402,N_13075,N_13864);
or UO_1403 (O_1403,N_14417,N_11414);
or UO_1404 (O_1404,N_12041,N_14729);
or UO_1405 (O_1405,N_13518,N_10276);
or UO_1406 (O_1406,N_13068,N_14025);
nand UO_1407 (O_1407,N_11220,N_14255);
nand UO_1408 (O_1408,N_11488,N_11806);
and UO_1409 (O_1409,N_12787,N_12939);
and UO_1410 (O_1410,N_13227,N_10158);
nand UO_1411 (O_1411,N_11995,N_13252);
and UO_1412 (O_1412,N_13070,N_13343);
nand UO_1413 (O_1413,N_10028,N_10231);
and UO_1414 (O_1414,N_14311,N_13947);
nand UO_1415 (O_1415,N_14486,N_10096);
or UO_1416 (O_1416,N_13707,N_10171);
nor UO_1417 (O_1417,N_11461,N_13568);
and UO_1418 (O_1418,N_13963,N_14196);
and UO_1419 (O_1419,N_10886,N_11855);
and UO_1420 (O_1420,N_11874,N_13857);
nor UO_1421 (O_1421,N_12071,N_14717);
and UO_1422 (O_1422,N_13612,N_10585);
nor UO_1423 (O_1423,N_14573,N_11188);
or UO_1424 (O_1424,N_10404,N_11148);
or UO_1425 (O_1425,N_12607,N_12039);
or UO_1426 (O_1426,N_11642,N_12748);
nand UO_1427 (O_1427,N_10896,N_12502);
and UO_1428 (O_1428,N_14990,N_13842);
and UO_1429 (O_1429,N_12908,N_12953);
or UO_1430 (O_1430,N_13949,N_13637);
nand UO_1431 (O_1431,N_12348,N_10691);
nor UO_1432 (O_1432,N_13303,N_11520);
or UO_1433 (O_1433,N_10758,N_12367);
nand UO_1434 (O_1434,N_11466,N_10556);
nand UO_1435 (O_1435,N_11479,N_14909);
or UO_1436 (O_1436,N_13129,N_11078);
and UO_1437 (O_1437,N_14010,N_10261);
and UO_1438 (O_1438,N_13248,N_13853);
nor UO_1439 (O_1439,N_10193,N_14361);
and UO_1440 (O_1440,N_14571,N_12319);
and UO_1441 (O_1441,N_13872,N_14966);
and UO_1442 (O_1442,N_11472,N_12322);
and UO_1443 (O_1443,N_11586,N_10681);
nand UO_1444 (O_1444,N_14607,N_12211);
nand UO_1445 (O_1445,N_13351,N_11211);
and UO_1446 (O_1446,N_13413,N_14213);
and UO_1447 (O_1447,N_14179,N_13081);
nand UO_1448 (O_1448,N_10953,N_13090);
nand UO_1449 (O_1449,N_12078,N_14156);
nand UO_1450 (O_1450,N_11846,N_12429);
and UO_1451 (O_1451,N_11579,N_11265);
or UO_1452 (O_1452,N_13609,N_12992);
and UO_1453 (O_1453,N_13136,N_14088);
and UO_1454 (O_1454,N_14144,N_11737);
and UO_1455 (O_1455,N_14366,N_11136);
nand UO_1456 (O_1456,N_11963,N_10520);
nor UO_1457 (O_1457,N_13012,N_10029);
nand UO_1458 (O_1458,N_11080,N_12950);
nor UO_1459 (O_1459,N_12732,N_13266);
or UO_1460 (O_1460,N_11476,N_14835);
and UO_1461 (O_1461,N_13873,N_13097);
nor UO_1462 (O_1462,N_12444,N_11489);
and UO_1463 (O_1463,N_11758,N_11707);
nand UO_1464 (O_1464,N_11950,N_10474);
nor UO_1465 (O_1465,N_10069,N_12956);
and UO_1466 (O_1466,N_13184,N_10574);
and UO_1467 (O_1467,N_13665,N_10748);
and UO_1468 (O_1468,N_11402,N_13939);
or UO_1469 (O_1469,N_10661,N_11640);
nor UO_1470 (O_1470,N_14738,N_11924);
nor UO_1471 (O_1471,N_10384,N_14652);
or UO_1472 (O_1472,N_13601,N_11570);
and UO_1473 (O_1473,N_11140,N_13886);
and UO_1474 (O_1474,N_10392,N_12596);
nor UO_1475 (O_1475,N_12762,N_10794);
nand UO_1476 (O_1476,N_11246,N_12194);
and UO_1477 (O_1477,N_14807,N_14058);
nand UO_1478 (O_1478,N_12234,N_10092);
nand UO_1479 (O_1479,N_12770,N_11786);
nand UO_1480 (O_1480,N_11868,N_13232);
or UO_1481 (O_1481,N_13349,N_10010);
nand UO_1482 (O_1482,N_11353,N_13243);
or UO_1483 (O_1483,N_10316,N_14849);
or UO_1484 (O_1484,N_10078,N_14087);
nor UO_1485 (O_1485,N_12156,N_10949);
and UO_1486 (O_1486,N_14138,N_10364);
or UO_1487 (O_1487,N_14167,N_10322);
nand UO_1488 (O_1488,N_13517,N_14504);
nor UO_1489 (O_1489,N_14776,N_13725);
nand UO_1490 (O_1490,N_14293,N_11940);
nor UO_1491 (O_1491,N_12029,N_14369);
and UO_1492 (O_1492,N_12500,N_11087);
nor UO_1493 (O_1493,N_12138,N_10977);
nand UO_1494 (O_1494,N_12034,N_13229);
nor UO_1495 (O_1495,N_12842,N_13929);
nor UO_1496 (O_1496,N_10032,N_13430);
nor UO_1497 (O_1497,N_10165,N_11528);
and UO_1498 (O_1498,N_12592,N_10659);
nand UO_1499 (O_1499,N_13497,N_11302);
or UO_1500 (O_1500,N_12126,N_13098);
and UO_1501 (O_1501,N_13083,N_14106);
nor UO_1502 (O_1502,N_12153,N_13531);
and UO_1503 (O_1503,N_13392,N_10458);
nand UO_1504 (O_1504,N_11343,N_11687);
nand UO_1505 (O_1505,N_13673,N_14148);
nor UO_1506 (O_1506,N_14525,N_10980);
nor UO_1507 (O_1507,N_10149,N_11981);
and UO_1508 (O_1508,N_12435,N_13142);
or UO_1509 (O_1509,N_13282,N_10715);
nor UO_1510 (O_1510,N_12630,N_11494);
or UO_1511 (O_1511,N_11559,N_10482);
and UO_1512 (O_1512,N_14348,N_13294);
and UO_1513 (O_1513,N_12019,N_13512);
or UO_1514 (O_1514,N_13147,N_12294);
nand UO_1515 (O_1515,N_11496,N_11069);
nor UO_1516 (O_1516,N_12679,N_14879);
nor UO_1517 (O_1517,N_13965,N_12520);
and UO_1518 (O_1518,N_11052,N_11552);
nor UO_1519 (O_1519,N_10425,N_13210);
and UO_1520 (O_1520,N_10023,N_13506);
nor UO_1521 (O_1521,N_11545,N_13552);
or UO_1522 (O_1522,N_11574,N_12362);
or UO_1523 (O_1523,N_11053,N_12291);
nand UO_1524 (O_1524,N_10237,N_13748);
nor UO_1525 (O_1525,N_13053,N_14065);
nand UO_1526 (O_1526,N_14999,N_13357);
and UO_1527 (O_1527,N_11184,N_11048);
and UO_1528 (O_1528,N_13203,N_14789);
and UO_1529 (O_1529,N_10178,N_11341);
or UO_1530 (O_1530,N_10215,N_10798);
and UO_1531 (O_1531,N_10904,N_13734);
nand UO_1532 (O_1532,N_11193,N_13263);
or UO_1533 (O_1533,N_10787,N_11486);
or UO_1534 (O_1534,N_14891,N_14998);
or UO_1535 (O_1535,N_13433,N_11812);
and UO_1536 (O_1536,N_11223,N_13359);
and UO_1537 (O_1537,N_13170,N_12977);
nand UO_1538 (O_1538,N_13131,N_12794);
or UO_1539 (O_1539,N_13199,N_14038);
or UO_1540 (O_1540,N_11991,N_11145);
and UO_1541 (O_1541,N_12555,N_13981);
or UO_1542 (O_1542,N_10749,N_12074);
or UO_1543 (O_1543,N_14619,N_13920);
nand UO_1544 (O_1544,N_11226,N_13174);
and UO_1545 (O_1545,N_10885,N_11558);
or UO_1546 (O_1546,N_11610,N_14383);
nand UO_1547 (O_1547,N_11857,N_10042);
nor UO_1548 (O_1548,N_11141,N_14956);
nand UO_1549 (O_1549,N_10989,N_10624);
or UO_1550 (O_1550,N_11608,N_11705);
or UO_1551 (O_1551,N_10978,N_14989);
nand UO_1552 (O_1552,N_12923,N_11763);
nor UO_1553 (O_1553,N_14443,N_12251);
or UO_1554 (O_1554,N_13807,N_10460);
or UO_1555 (O_1555,N_11790,N_12186);
and UO_1556 (O_1556,N_11373,N_14260);
and UO_1557 (O_1557,N_11531,N_10250);
or UO_1558 (O_1558,N_10983,N_12270);
and UO_1559 (O_1559,N_11318,N_14551);
and UO_1560 (O_1560,N_14617,N_14448);
or UO_1561 (O_1561,N_10133,N_11208);
nor UO_1562 (O_1562,N_10642,N_10984);
or UO_1563 (O_1563,N_12539,N_10710);
or UO_1564 (O_1564,N_12835,N_12066);
or UO_1565 (O_1565,N_13270,N_14072);
and UO_1566 (O_1566,N_14084,N_13820);
nand UO_1567 (O_1567,N_13310,N_13887);
and UO_1568 (O_1568,N_14766,N_13021);
nand UO_1569 (O_1569,N_13885,N_13902);
or UO_1570 (O_1570,N_14902,N_13304);
and UO_1571 (O_1571,N_13250,N_10051);
and UO_1572 (O_1572,N_13434,N_10888);
xor UO_1573 (O_1573,N_13078,N_10434);
nand UO_1574 (O_1574,N_14812,N_11589);
nand UO_1575 (O_1575,N_14698,N_11669);
and UO_1576 (O_1576,N_13697,N_12749);
nor UO_1577 (O_1577,N_11538,N_14270);
nand UO_1578 (O_1578,N_11323,N_11173);
and UO_1579 (O_1579,N_10593,N_11194);
nor UO_1580 (O_1580,N_10588,N_14534);
nor UO_1581 (O_1581,N_10746,N_12476);
nor UO_1582 (O_1582,N_10047,N_14892);
nand UO_1583 (O_1583,N_10705,N_14683);
and UO_1584 (O_1584,N_13614,N_13148);
and UO_1585 (O_1585,N_14076,N_11753);
nand UO_1586 (O_1586,N_11213,N_13468);
nor UO_1587 (O_1587,N_14306,N_14387);
or UO_1588 (O_1588,N_14118,N_13300);
nand UO_1589 (O_1589,N_10808,N_12225);
nand UO_1590 (O_1590,N_10066,N_14616);
nor UO_1591 (O_1591,N_14433,N_10970);
nand UO_1592 (O_1592,N_11182,N_11996);
and UO_1593 (O_1593,N_10833,N_14233);
nor UO_1594 (O_1594,N_10205,N_10690);
nor UO_1595 (O_1595,N_11526,N_14043);
or UO_1596 (O_1596,N_14175,N_13906);
nand UO_1597 (O_1597,N_11329,N_10852);
and UO_1598 (O_1598,N_13062,N_13212);
or UO_1599 (O_1599,N_14511,N_12481);
and UO_1600 (O_1600,N_10344,N_13127);
nand UO_1601 (O_1601,N_12203,N_12545);
and UO_1602 (O_1602,N_12541,N_14499);
nor UO_1603 (O_1603,N_10536,N_12065);
and UO_1604 (O_1604,N_14257,N_12114);
nand UO_1605 (O_1605,N_11384,N_14193);
or UO_1606 (O_1606,N_10779,N_10311);
nor UO_1607 (O_1607,N_10726,N_12707);
or UO_1608 (O_1608,N_12106,N_10541);
or UO_1609 (O_1609,N_11699,N_14917);
nor UO_1610 (O_1610,N_13156,N_14540);
and UO_1611 (O_1611,N_12490,N_14317);
or UO_1612 (O_1612,N_10608,N_14842);
or UO_1613 (O_1613,N_12644,N_11907);
and UO_1614 (O_1614,N_10394,N_12454);
nor UO_1615 (O_1615,N_12366,N_12660);
nor UO_1616 (O_1616,N_13355,N_13973);
nor UO_1617 (O_1617,N_14225,N_10527);
nor UO_1618 (O_1618,N_12439,N_13356);
nor UO_1619 (O_1619,N_12214,N_13084);
nand UO_1620 (O_1620,N_12047,N_13829);
or UO_1621 (O_1621,N_14192,N_14250);
nor UO_1622 (O_1622,N_14364,N_13666);
nand UO_1623 (O_1623,N_13813,N_11624);
nand UO_1624 (O_1624,N_13532,N_10735);
nand UO_1625 (O_1625,N_14791,N_13009);
and UO_1626 (O_1626,N_13287,N_10603);
or UO_1627 (O_1627,N_14468,N_12310);
or UO_1628 (O_1628,N_11688,N_10521);
nand UO_1629 (O_1629,N_13851,N_12779);
nor UO_1630 (O_1630,N_14119,N_10616);
nand UO_1631 (O_1631,N_11542,N_14137);
or UO_1632 (O_1632,N_13418,N_13006);
nand UO_1633 (O_1633,N_13115,N_12552);
nand UO_1634 (O_1634,N_13164,N_12333);
or UO_1635 (O_1635,N_13133,N_14183);
or UO_1636 (O_1636,N_10674,N_14343);
nand UO_1637 (O_1637,N_11278,N_13290);
and UO_1638 (O_1638,N_11810,N_11850);
and UO_1639 (O_1639,N_11573,N_12132);
nand UO_1640 (O_1640,N_10112,N_14815);
nor UO_1641 (O_1641,N_12133,N_11557);
nand UO_1642 (O_1642,N_13002,N_14651);
or UO_1643 (O_1643,N_10785,N_11198);
nor UO_1644 (O_1644,N_12796,N_11157);
nand UO_1645 (O_1645,N_13299,N_10531);
and UO_1646 (O_1646,N_13020,N_14273);
nand UO_1647 (O_1647,N_13370,N_11748);
or UO_1648 (O_1648,N_12492,N_14548);
or UO_1649 (O_1649,N_14959,N_11247);
or UO_1650 (O_1650,N_13622,N_13027);
nor UO_1651 (O_1651,N_10241,N_10685);
or UO_1652 (O_1652,N_11162,N_11739);
and UO_1653 (O_1653,N_13676,N_10233);
nor UO_1654 (O_1654,N_10145,N_14885);
nor UO_1655 (O_1655,N_13189,N_12470);
nand UO_1656 (O_1656,N_14378,N_10894);
and UO_1657 (O_1657,N_13198,N_11892);
and UO_1658 (O_1658,N_11780,N_13429);
or UO_1659 (O_1659,N_11801,N_14950);
and UO_1660 (O_1660,N_14232,N_13670);
and UO_1661 (O_1661,N_14936,N_12669);
and UO_1662 (O_1662,N_13175,N_14159);
nor UO_1663 (O_1663,N_14984,N_10617);
nor UO_1664 (O_1664,N_14578,N_11749);
nand UO_1665 (O_1665,N_11774,N_11448);
nor UO_1666 (O_1666,N_10485,N_10264);
nand UO_1667 (O_1667,N_12344,N_11948);
and UO_1668 (O_1668,N_14236,N_10918);
nor UO_1669 (O_1669,N_13551,N_14974);
or UO_1670 (O_1670,N_11107,N_13308);
nand UO_1671 (O_1671,N_12947,N_14915);
nor UO_1672 (O_1672,N_14060,N_11638);
or UO_1673 (O_1673,N_13910,N_12358);
or UO_1674 (O_1674,N_10124,N_12236);
nor UO_1675 (O_1675,N_10488,N_11233);
or UO_1676 (O_1676,N_13642,N_13980);
and UO_1677 (O_1677,N_13797,N_11970);
and UO_1678 (O_1678,N_13819,N_10835);
nand UO_1679 (O_1679,N_10772,N_14291);
or UO_1680 (O_1680,N_12783,N_10346);
nand UO_1681 (O_1681,N_14979,N_14639);
nand UO_1682 (O_1682,N_12666,N_12197);
and UO_1683 (O_1683,N_11516,N_10929);
and UO_1684 (O_1684,N_13228,N_14243);
nor UO_1685 (O_1685,N_14587,N_12840);
or UO_1686 (O_1686,N_12756,N_11839);
nand UO_1687 (O_1687,N_12619,N_10381);
and UO_1688 (O_1688,N_13698,N_14063);
nand UO_1689 (O_1689,N_10142,N_10452);
or UO_1690 (O_1690,N_11134,N_12755);
and UO_1691 (O_1691,N_12403,N_10670);
or UO_1692 (O_1692,N_11006,N_11498);
and UO_1693 (O_1693,N_10003,N_14543);
nor UO_1694 (O_1694,N_14436,N_11251);
nand UO_1695 (O_1695,N_11054,N_12266);
or UO_1696 (O_1696,N_11988,N_11747);
and UO_1697 (O_1697,N_14690,N_12774);
and UO_1698 (O_1698,N_12616,N_10291);
nor UO_1699 (O_1699,N_12289,N_11567);
or UO_1700 (O_1700,N_12416,N_12757);
nand UO_1701 (O_1701,N_13843,N_14120);
or UO_1702 (O_1702,N_10908,N_11016);
nor UO_1703 (O_1703,N_10362,N_12852);
and UO_1704 (O_1704,N_10934,N_13968);
or UO_1705 (O_1705,N_10901,N_10224);
nor UO_1706 (O_1706,N_12050,N_10761);
or UO_1707 (O_1707,N_12415,N_12055);
and UO_1708 (O_1708,N_12442,N_12324);
or UO_1709 (O_1709,N_11210,N_12032);
nor UO_1710 (O_1710,N_12799,N_12913);
or UO_1711 (O_1711,N_10126,N_12062);
and UO_1712 (O_1712,N_11954,N_11064);
or UO_1713 (O_1713,N_12510,N_10440);
nand UO_1714 (O_1714,N_12239,N_10678);
or UO_1715 (O_1715,N_10897,N_12209);
xor UO_1716 (O_1716,N_12569,N_13950);
nand UO_1717 (O_1717,N_10471,N_10442);
and UO_1718 (O_1718,N_12746,N_10838);
and UO_1719 (O_1719,N_12201,N_12736);
nor UO_1720 (O_1720,N_10483,N_11257);
nor UO_1721 (O_1721,N_10774,N_12247);
and UO_1722 (O_1722,N_11609,N_11172);
nand UO_1723 (O_1723,N_12022,N_10212);
nor UO_1724 (O_1724,N_10595,N_11124);
or UO_1725 (O_1725,N_12151,N_10812);
nor UO_1726 (O_1726,N_10333,N_13325);
and UO_1727 (O_1727,N_13567,N_14827);
nand UO_1728 (O_1728,N_11383,N_10540);
nor UO_1729 (O_1729,N_11350,N_13408);
or UO_1730 (O_1730,N_11199,N_10546);
nor UO_1731 (O_1731,N_10424,N_11227);
or UO_1732 (O_1732,N_13926,N_13654);
or UO_1733 (O_1733,N_13442,N_10091);
or UO_1734 (O_1734,N_11601,N_13625);
nand UO_1735 (O_1735,N_14707,N_12410);
or UO_1736 (O_1736,N_10098,N_10856);
and UO_1737 (O_1737,N_13617,N_13937);
or UO_1738 (O_1738,N_14178,N_14932);
nor UO_1739 (O_1739,N_12530,N_10693);
and UO_1740 (O_1740,N_11274,N_11281);
nor UO_1741 (O_1741,N_13007,N_14694);
nand UO_1742 (O_1742,N_10148,N_12847);
and UO_1743 (O_1743,N_14122,N_10850);
and UO_1744 (O_1744,N_13801,N_12048);
nand UO_1745 (O_1745,N_14007,N_12297);
xnor UO_1746 (O_1746,N_14559,N_13722);
nand UO_1747 (O_1747,N_12614,N_10175);
nor UO_1748 (O_1748,N_14081,N_13470);
nand UO_1749 (O_1749,N_14205,N_13825);
and UO_1750 (O_1750,N_11503,N_13703);
or UO_1751 (O_1751,N_11352,N_14204);
nor UO_1752 (O_1752,N_10766,N_13089);
nand UO_1753 (O_1753,N_14545,N_14579);
or UO_1754 (O_1754,N_14792,N_11990);
and UO_1755 (O_1755,N_14640,N_13624);
and UO_1756 (O_1756,N_12080,N_13688);
nor UO_1757 (O_1757,N_10820,N_12925);
nor UO_1758 (O_1758,N_11007,N_10467);
and UO_1759 (O_1759,N_11939,N_14933);
and UO_1760 (O_1760,N_12720,N_13390);
nand UO_1761 (O_1761,N_12999,N_11554);
nand UO_1762 (O_1762,N_11480,N_10860);
nor UO_1763 (O_1763,N_13026,N_11456);
or UO_1764 (O_1764,N_14681,N_10432);
nand UO_1765 (O_1765,N_11364,N_12813);
or UO_1766 (O_1766,N_13814,N_10339);
and UO_1767 (O_1767,N_10183,N_11604);
and UO_1768 (O_1768,N_12642,N_10323);
nand UO_1769 (O_1769,N_14457,N_10022);
nor UO_1770 (O_1770,N_12874,N_14046);
or UO_1771 (O_1771,N_14285,N_14653);
nand UO_1772 (O_1772,N_12597,N_13656);
nand UO_1773 (O_1773,N_14746,N_11978);
nand UO_1774 (O_1774,N_13312,N_12862);
and UO_1775 (O_1775,N_11418,N_10195);
nand UO_1776 (O_1776,N_14858,N_10903);
and UO_1777 (O_1777,N_10169,N_10959);
and UO_1778 (O_1778,N_11595,N_13984);
or UO_1779 (O_1779,N_10130,N_12599);
and UO_1780 (O_1780,N_14855,N_10832);
nand UO_1781 (O_1781,N_13414,N_13319);
nor UO_1782 (O_1782,N_13087,N_11106);
nor UO_1783 (O_1783,N_10890,N_14037);
or UO_1784 (O_1784,N_12900,N_13611);
nor UO_1785 (O_1785,N_14305,N_14801);
nand UO_1786 (O_1786,N_11553,N_13267);
or UO_1787 (O_1787,N_12401,N_11799);
or UO_1788 (O_1788,N_10701,N_13377);
or UO_1789 (O_1789,N_11944,N_12286);
nand UO_1790 (O_1790,N_12934,N_12350);
nand UO_1791 (O_1791,N_13028,N_11252);
nand UO_1792 (O_1792,N_12764,N_14012);
or UO_1793 (O_1793,N_13836,N_14133);
and UO_1794 (O_1794,N_11891,N_11634);
or UO_1795 (O_1795,N_10639,N_14968);
nand UO_1796 (O_1796,N_11089,N_12036);
nand UO_1797 (O_1797,N_12128,N_10187);
and UO_1798 (O_1798,N_12226,N_10080);
and UO_1799 (O_1799,N_11720,N_13619);
and UO_1800 (O_1800,N_12897,N_10239);
nand UO_1801 (O_1801,N_13786,N_11742);
or UO_1802 (O_1802,N_10729,N_14117);
and UO_1803 (O_1803,N_13581,N_13916);
and UO_1804 (O_1804,N_11283,N_13329);
nand UO_1805 (O_1805,N_13934,N_14518);
nor UO_1806 (O_1806,N_13145,N_14216);
nand UO_1807 (O_1807,N_14170,N_11836);
nand UO_1808 (O_1808,N_12675,N_14648);
nor UO_1809 (O_1809,N_13790,N_10960);
nand UO_1810 (O_1810,N_11667,N_11357);
or UO_1811 (O_1811,N_12152,N_11396);
and UO_1812 (O_1812,N_11693,N_11221);
and UO_1813 (O_1813,N_12621,N_10548);
nor UO_1814 (O_1814,N_10598,N_12944);
or UO_1815 (O_1815,N_10840,N_14299);
nor UO_1816 (O_1816,N_14897,N_11986);
nor UO_1817 (O_1817,N_12357,N_14868);
nor UO_1818 (O_1818,N_13653,N_14279);
or UO_1819 (O_1819,N_10185,N_14724);
nand UO_1820 (O_1820,N_10778,N_12649);
nor UO_1821 (O_1821,N_14834,N_12521);
nor UO_1822 (O_1822,N_14372,N_12328);
nand UO_1823 (O_1823,N_11337,N_12602);
nand UO_1824 (O_1824,N_13402,N_12958);
and UO_1825 (O_1825,N_13594,N_14958);
or UO_1826 (O_1826,N_11809,N_13269);
nor UO_1827 (O_1827,N_13994,N_10581);
or UO_1828 (O_1828,N_13406,N_14328);
or UO_1829 (O_1829,N_11647,N_11681);
nor UO_1830 (O_1830,N_11582,N_12409);
and UO_1831 (O_1831,N_14929,N_13502);
nand UO_1832 (O_1832,N_12584,N_14057);
nand UO_1833 (O_1833,N_12303,N_10338);
or UO_1834 (O_1834,N_11662,N_14824);
nor UO_1835 (O_1835,N_12150,N_13183);
or UO_1836 (O_1836,N_14166,N_12488);
nor UO_1837 (O_1837,N_14773,N_11340);
nand UO_1838 (O_1838,N_10614,N_14223);
and UO_1839 (O_1839,N_13802,N_11138);
nor UO_1840 (O_1840,N_12445,N_13462);
or UO_1841 (O_1841,N_13118,N_13951);
and UO_1842 (O_1842,N_14795,N_14208);
or UO_1843 (O_1843,N_12740,N_14026);
and UO_1844 (O_1844,N_10728,N_10222);
and UO_1845 (O_1845,N_14465,N_11914);
nand UO_1846 (O_1846,N_11548,N_10968);
and UO_1847 (O_1847,N_11072,N_11272);
nand UO_1848 (O_1848,N_13849,N_10217);
or UO_1849 (O_1849,N_11818,N_11037);
or UO_1850 (O_1850,N_13623,N_11028);
nor UO_1851 (O_1851,N_12273,N_13082);
and UO_1852 (O_1852,N_12731,N_12035);
and UO_1853 (O_1853,N_10325,N_10911);
and UO_1854 (O_1854,N_14684,N_12067);
nand UO_1855 (O_1855,N_11938,N_13810);
or UO_1856 (O_1856,N_11897,N_14128);
nand UO_1857 (O_1857,N_11137,N_10054);
or UO_1858 (O_1858,N_14719,N_12650);
or UO_1859 (O_1859,N_11433,N_10776);
nand UO_1860 (O_1860,N_10712,N_13238);
and UO_1861 (O_1861,N_14352,N_10410);
nor UO_1862 (O_1862,N_11391,N_11325);
and UO_1863 (O_1863,N_14532,N_13956);
and UO_1864 (O_1864,N_14614,N_11718);
and UO_1865 (O_1865,N_10753,N_14151);
and UO_1866 (O_1866,N_14629,N_13029);
nor UO_1867 (O_1867,N_14114,N_11202);
or UO_1868 (O_1868,N_11457,N_13928);
nand UO_1869 (O_1869,N_11577,N_12933);
and UO_1870 (O_1870,N_13123,N_12264);
and UO_1871 (O_1871,N_14516,N_11362);
and UO_1872 (O_1872,N_12113,N_10116);
nand UO_1873 (O_1873,N_14227,N_12155);
or UO_1874 (O_1874,N_10606,N_13461);
or UO_1875 (O_1875,N_14152,N_14322);
or UO_1876 (O_1876,N_12742,N_13110);
nand UO_1877 (O_1877,N_10341,N_13037);
and UO_1878 (O_1878,N_14365,N_11813);
nand UO_1879 (O_1879,N_12017,N_14737);
and UO_1880 (O_1880,N_12473,N_14685);
and UO_1881 (O_1881,N_12693,N_14521);
and UO_1882 (O_1882,N_14030,N_11674);
nand UO_1883 (O_1883,N_10226,N_14646);
and UO_1884 (O_1884,N_10920,N_11298);
and UO_1885 (O_1885,N_13220,N_12909);
and UO_1886 (O_1886,N_13961,N_13695);
and UO_1887 (O_1887,N_10152,N_12365);
nand UO_1888 (O_1888,N_14004,N_10182);
or UO_1889 (O_1889,N_11912,N_10389);
and UO_1890 (O_1890,N_11639,N_13190);
nand UO_1891 (O_1891,N_10936,N_12309);
nand UO_1892 (O_1892,N_11206,N_14711);
nor UO_1893 (O_1893,N_14816,N_12046);
and UO_1894 (O_1894,N_12844,N_13373);
and UO_1895 (O_1895,N_13765,N_14982);
and UO_1896 (O_1896,N_10857,N_11027);
nand UO_1897 (O_1897,N_14464,N_10258);
nand UO_1898 (O_1898,N_11686,N_14497);
nor UO_1899 (O_1899,N_10650,N_14214);
nand UO_1900 (O_1900,N_14337,N_13501);
nor UO_1901 (O_1901,N_10529,N_11361);
and UO_1902 (O_1902,N_13233,N_11204);
and UO_1903 (O_1903,N_11794,N_13821);
or UO_1904 (O_1904,N_10382,N_14572);
or UO_1905 (O_1905,N_14631,N_10730);
nand UO_1906 (O_1906,N_14798,N_13741);
nand UO_1907 (O_1907,N_10957,N_14461);
nor UO_1908 (O_1908,N_13896,N_13450);
or UO_1909 (O_1909,N_13428,N_10839);
and UO_1910 (O_1910,N_13540,N_11326);
or UO_1911 (O_1911,N_12143,N_12146);
nand UO_1912 (O_1912,N_13455,N_14301);
nor UO_1913 (O_1913,N_11588,N_10235);
or UO_1914 (O_1914,N_11249,N_13840);
nand UO_1915 (O_1915,N_14794,N_13457);
nor UO_1916 (O_1916,N_12177,N_11484);
nor UO_1917 (O_1917,N_13799,N_11641);
nor UO_1918 (O_1918,N_12673,N_12159);
nor UO_1919 (O_1919,N_11760,N_11230);
nand UO_1920 (O_1920,N_13231,N_13017);
and UO_1921 (O_1921,N_14764,N_14437);
and UO_1922 (O_1922,N_12360,N_13121);
nor UO_1923 (O_1923,N_14777,N_11569);
nand UO_1924 (O_1924,N_13415,N_11346);
or UO_1925 (O_1925,N_12617,N_14650);
nand UO_1926 (O_1926,N_14220,N_14116);
and UO_1927 (O_1927,N_11139,N_13661);
nand UO_1928 (O_1928,N_13024,N_11784);
and UO_1929 (O_1929,N_13767,N_12846);
and UO_1930 (O_1930,N_13644,N_13443);
and UO_1931 (O_1931,N_12359,N_14693);
nor UO_1932 (O_1932,N_11021,N_12680);
or UO_1933 (O_1933,N_12582,N_13809);
nor UO_1934 (O_1934,N_14537,N_11875);
nand UO_1935 (O_1935,N_11445,N_14438);
and UO_1936 (O_1936,N_14018,N_13621);
nor UO_1937 (O_1937,N_13001,N_14340);
nor UO_1938 (O_1938,N_14219,N_14752);
and UO_1939 (O_1939,N_11619,N_13936);
or UO_1940 (O_1940,N_10589,N_11636);
or UO_1941 (O_1941,N_10056,N_14536);
nor UO_1942 (O_1942,N_14725,N_13982);
nand UO_1943 (O_1943,N_10629,N_11633);
nor UO_1944 (O_1944,N_14460,N_10623);
nand UO_1945 (O_1945,N_10695,N_13839);
or UO_1946 (O_1946,N_13202,N_12928);
nor UO_1947 (O_1947,N_11044,N_14555);
nand UO_1948 (O_1948,N_13361,N_11005);
nor UO_1949 (O_1949,N_10279,N_12170);
nand UO_1950 (O_1950,N_11972,N_12804);
nor UO_1951 (O_1951,N_12553,N_12073);
and UO_1952 (O_1952,N_11086,N_10999);
and UO_1953 (O_1953,N_12926,N_10900);
and UO_1954 (O_1954,N_13527,N_12670);
and UO_1955 (O_1955,N_10248,N_11079);
and UO_1956 (O_1956,N_11017,N_10266);
or UO_1957 (O_1957,N_10635,N_11293);
or UO_1958 (O_1958,N_11412,N_14906);
nand UO_1959 (O_1959,N_13034,N_13475);
nand UO_1960 (O_1960,N_10516,N_14503);
and UO_1961 (O_1961,N_14472,N_14787);
and UO_1962 (O_1962,N_12878,N_13422);
nand UO_1963 (O_1963,N_10763,N_12564);
nand UO_1964 (O_1964,N_12140,N_12045);
or UO_1965 (O_1965,N_10015,N_12184);
or UO_1966 (O_1966,N_12325,N_10630);
or UO_1967 (O_1967,N_13955,N_10848);
and UO_1968 (O_1968,N_12773,N_11522);
or UO_1969 (O_1969,N_11263,N_11778);
and UO_1970 (O_1970,N_14873,N_12754);
nor UO_1971 (O_1971,N_13855,N_14926);
nand UO_1972 (O_1972,N_12405,N_12108);
nand UO_1973 (O_1973,N_10255,N_11736);
and UO_1974 (O_1974,N_13205,N_13555);
nand UO_1975 (O_1975,N_10475,N_13291);
and UO_1976 (O_1976,N_10100,N_12187);
nor UO_1977 (O_1977,N_13749,N_12912);
and UO_1978 (O_1978,N_13784,N_14041);
and UO_1979 (O_1979,N_12260,N_12940);
nor UO_1980 (O_1980,N_13785,N_13556);
and UO_1981 (O_1981,N_12097,N_14515);
or UO_1982 (O_1982,N_14375,N_14995);
nand UO_1983 (O_1983,N_12767,N_12973);
or UO_1984 (O_1984,N_13519,N_11119);
nor UO_1985 (O_1985,N_13042,N_12763);
or UO_1986 (O_1986,N_12702,N_11505);
or UO_1987 (O_1987,N_14802,N_10893);
or UO_1988 (O_1988,N_10329,N_10708);
and UO_1989 (O_1989,N_12195,N_14784);
or UO_1990 (O_1990,N_13272,N_11153);
and UO_1991 (O_1991,N_10489,N_12574);
and UO_1992 (O_1992,N_12063,N_10643);
or UO_1993 (O_1993,N_13061,N_10354);
nand UO_1994 (O_1994,N_11004,N_14637);
or UO_1995 (O_1995,N_11032,N_14104);
and UO_1996 (O_1996,N_13168,N_12665);
nor UO_1997 (O_1997,N_11710,N_12662);
and UO_1998 (O_1998,N_14261,N_14977);
and UO_1999 (O_1999,N_12954,N_13498);
endmodule