module basic_500_3000_500_60_levels_5xor_2(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
or U0 (N_0,In_430,In_122);
and U1 (N_1,In_135,In_455);
nand U2 (N_2,In_294,In_95);
nor U3 (N_3,In_8,In_87);
and U4 (N_4,In_249,In_285);
and U5 (N_5,In_219,In_327);
nor U6 (N_6,In_382,In_470);
xnor U7 (N_7,In_319,In_291);
nand U8 (N_8,In_460,In_148);
or U9 (N_9,In_245,In_224);
or U10 (N_10,In_447,In_258);
nor U11 (N_11,In_69,In_203);
nor U12 (N_12,In_488,In_215);
nand U13 (N_13,In_45,In_247);
or U14 (N_14,In_237,In_263);
or U15 (N_15,In_453,In_162);
nor U16 (N_16,In_474,In_50);
nand U17 (N_17,In_201,In_322);
or U18 (N_18,In_329,In_7);
nand U19 (N_19,In_265,In_317);
or U20 (N_20,In_53,In_281);
or U21 (N_21,In_138,In_226);
xor U22 (N_22,In_487,In_164);
or U23 (N_23,In_129,In_229);
nand U24 (N_24,In_288,In_289);
and U25 (N_25,In_283,In_255);
xnor U26 (N_26,In_494,In_275);
xor U27 (N_27,In_57,In_132);
nand U28 (N_28,In_19,In_480);
and U29 (N_29,In_457,In_368);
or U30 (N_30,In_101,In_114);
xnor U31 (N_31,In_104,In_91);
nor U32 (N_32,In_436,In_12);
nand U33 (N_33,In_34,In_15);
and U34 (N_34,In_166,In_261);
nor U35 (N_35,In_153,In_360);
nand U36 (N_36,In_223,In_313);
and U37 (N_37,In_102,In_9);
and U38 (N_38,In_0,In_358);
nand U39 (N_39,In_344,In_268);
nand U40 (N_40,In_168,In_343);
and U41 (N_41,In_5,In_364);
or U42 (N_42,In_48,In_361);
nor U43 (N_43,In_394,In_303);
and U44 (N_44,In_362,In_46);
and U45 (N_45,In_434,In_80);
and U46 (N_46,In_190,In_276);
and U47 (N_47,In_120,In_2);
or U48 (N_48,In_254,In_318);
and U49 (N_49,In_170,In_188);
nand U50 (N_50,N_7,In_330);
and U51 (N_51,In_356,N_33);
and U52 (N_52,In_11,In_85);
nor U53 (N_53,In_137,In_30);
nand U54 (N_54,In_279,In_159);
xnor U55 (N_55,In_408,In_181);
xnor U56 (N_56,In_131,In_495);
xor U57 (N_57,In_174,In_77);
and U58 (N_58,In_435,In_272);
nor U59 (N_59,In_139,In_476);
and U60 (N_60,In_336,In_88);
xor U61 (N_61,N_37,In_419);
xor U62 (N_62,In_482,In_340);
nand U63 (N_63,In_301,In_209);
nand U64 (N_64,In_412,In_115);
nor U65 (N_65,In_172,In_179);
or U66 (N_66,In_230,In_378);
nor U67 (N_67,In_388,In_269);
nor U68 (N_68,In_380,In_267);
nor U69 (N_69,In_489,In_176);
nand U70 (N_70,N_21,In_103);
nand U71 (N_71,In_257,In_297);
nor U72 (N_72,In_227,In_234);
nor U73 (N_73,In_220,In_189);
and U74 (N_74,In_441,N_6);
and U75 (N_75,In_497,N_22);
or U76 (N_76,N_32,In_149);
or U77 (N_77,In_280,In_42);
xnor U78 (N_78,In_61,In_338);
and U79 (N_79,In_262,In_473);
or U80 (N_80,In_182,In_105);
xnor U81 (N_81,N_48,In_490);
and U82 (N_82,N_20,In_199);
nor U83 (N_83,N_28,In_130);
and U84 (N_84,In_16,In_242);
or U85 (N_85,In_461,In_421);
nor U86 (N_86,In_18,In_373);
nand U87 (N_87,In_55,In_399);
or U88 (N_88,In_161,N_41);
and U89 (N_89,In_180,In_450);
nor U90 (N_90,In_354,In_266);
nor U91 (N_91,In_391,In_331);
and U92 (N_92,In_143,In_32);
xor U93 (N_93,In_481,In_54);
or U94 (N_94,In_411,In_33);
and U95 (N_95,In_312,In_405);
nor U96 (N_96,In_35,In_328);
nand U97 (N_97,In_410,In_194);
nand U98 (N_98,In_60,In_156);
nor U99 (N_99,In_370,In_438);
or U100 (N_100,In_376,In_251);
nor U101 (N_101,In_66,In_377);
xor U102 (N_102,In_81,In_459);
and U103 (N_103,In_348,In_345);
or U104 (N_104,In_27,N_40);
and U105 (N_105,In_456,In_25);
and U106 (N_106,In_432,N_2);
xor U107 (N_107,In_82,In_195);
and U108 (N_108,In_483,In_24);
or U109 (N_109,N_77,In_347);
nor U110 (N_110,In_468,In_386);
nor U111 (N_111,In_284,In_260);
nand U112 (N_112,In_454,In_420);
nand U113 (N_113,In_274,N_59);
xnor U114 (N_114,In_4,N_26);
nor U115 (N_115,In_379,In_165);
nor U116 (N_116,In_425,In_145);
nor U117 (N_117,In_383,N_71);
nor U118 (N_118,N_70,In_28);
nand U119 (N_119,N_90,In_31);
nor U120 (N_120,In_499,In_416);
nor U121 (N_121,In_37,In_236);
or U122 (N_122,In_295,N_9);
xnor U123 (N_123,In_466,In_211);
nor U124 (N_124,In_116,In_21);
or U125 (N_125,N_73,In_350);
or U126 (N_126,In_372,In_365);
xnor U127 (N_127,In_302,In_47);
and U128 (N_128,In_369,In_307);
or U129 (N_129,N_23,N_83);
nor U130 (N_130,In_415,In_93);
and U131 (N_131,In_171,In_73);
nand U132 (N_132,In_185,In_100);
nor U133 (N_133,In_467,N_66);
nor U134 (N_134,In_29,In_332);
nand U135 (N_135,In_306,N_13);
or U136 (N_136,N_18,In_452);
nor U137 (N_137,In_205,In_134);
and U138 (N_138,N_82,In_406);
and U139 (N_139,In_3,In_250);
and U140 (N_140,In_68,N_95);
and U141 (N_141,In_207,In_496);
nor U142 (N_142,In_469,In_397);
xnor U143 (N_143,In_197,In_385);
nor U144 (N_144,In_67,In_20);
and U145 (N_145,N_3,In_426);
and U146 (N_146,In_51,In_106);
nand U147 (N_147,In_125,N_47);
and U148 (N_148,In_191,In_244);
xnor U149 (N_149,In_259,In_335);
or U150 (N_150,N_148,N_129);
xor U151 (N_151,In_56,In_124);
or U152 (N_152,In_71,In_225);
and U153 (N_153,N_143,N_78);
nor U154 (N_154,In_392,N_87);
and U155 (N_155,In_63,In_186);
or U156 (N_156,In_217,In_300);
nand U157 (N_157,In_290,N_135);
and U158 (N_158,N_62,N_24);
or U159 (N_159,In_401,In_58);
nor U160 (N_160,N_116,In_393);
nand U161 (N_161,In_173,In_374);
nand U162 (N_162,In_359,N_46);
nand U163 (N_163,N_4,In_38);
nand U164 (N_164,N_85,In_310);
or U165 (N_165,N_76,In_167);
nand U166 (N_166,N_128,In_144);
nor U167 (N_167,N_106,In_158);
nor U168 (N_168,N_38,In_112);
nor U169 (N_169,In_70,In_273);
and U170 (N_170,N_112,In_41);
or U171 (N_171,In_418,In_314);
and U172 (N_172,N_127,In_342);
and U173 (N_173,In_427,N_88);
or U174 (N_174,In_346,In_187);
and U175 (N_175,N_75,In_395);
or U176 (N_176,In_6,N_145);
nor U177 (N_177,In_271,In_121);
nor U178 (N_178,N_35,In_155);
and U179 (N_179,In_320,In_212);
nor U180 (N_180,In_353,In_398);
nor U181 (N_181,In_216,N_60);
nor U182 (N_182,N_117,In_142);
xnor U183 (N_183,N_146,In_221);
xor U184 (N_184,In_52,In_118);
and U185 (N_185,N_57,N_121);
and U186 (N_186,In_484,In_133);
or U187 (N_187,In_475,In_107);
or U188 (N_188,N_93,In_315);
nor U189 (N_189,In_357,In_127);
nand U190 (N_190,N_119,In_471);
nor U191 (N_191,In_384,N_29);
nand U192 (N_192,In_444,In_65);
nor U193 (N_193,N_125,In_140);
nand U194 (N_194,In_177,In_407);
or U195 (N_195,N_36,In_367);
or U196 (N_196,In_10,In_49);
xnor U197 (N_197,In_94,In_443);
nor U198 (N_198,In_208,In_477);
and U199 (N_199,In_198,In_429);
or U200 (N_200,In_286,In_351);
nand U201 (N_201,In_13,N_14);
nand U202 (N_202,In_123,In_375);
or U203 (N_203,N_5,In_64);
or U204 (N_204,In_472,N_132);
and U205 (N_205,N_199,N_155);
nor U206 (N_206,In_409,In_14);
and U207 (N_207,N_110,In_293);
nand U208 (N_208,In_113,N_54);
xor U209 (N_209,N_149,In_163);
or U210 (N_210,N_154,N_140);
and U211 (N_211,In_193,N_190);
or U212 (N_212,In_431,In_72);
xor U213 (N_213,N_120,N_94);
and U214 (N_214,In_462,N_172);
xnor U215 (N_215,N_138,N_182);
nor U216 (N_216,In_491,In_59);
xnor U217 (N_217,In_43,In_445);
nor U218 (N_218,In_109,In_1);
or U219 (N_219,In_248,In_23);
xor U220 (N_220,In_108,N_107);
xor U221 (N_221,N_72,In_126);
xnor U222 (N_222,N_197,In_228);
and U223 (N_223,N_166,N_187);
xor U224 (N_224,N_109,N_27);
nand U225 (N_225,N_1,In_98);
nor U226 (N_226,In_119,In_324);
and U227 (N_227,In_465,In_381);
nor U228 (N_228,In_192,In_110);
nor U229 (N_229,N_8,N_180);
and U230 (N_230,In_175,In_389);
and U231 (N_231,In_252,N_139);
and U232 (N_232,In_264,In_287);
nand U233 (N_233,N_58,In_270);
nand U234 (N_234,In_240,In_246);
or U235 (N_235,N_165,N_185);
xor U236 (N_236,In_62,In_39);
or U237 (N_237,In_439,In_213);
xor U238 (N_238,In_233,In_363);
nand U239 (N_239,In_222,In_89);
and U240 (N_240,N_174,N_89);
nand U241 (N_241,N_34,N_43);
xor U242 (N_242,N_25,N_150);
nand U243 (N_243,In_117,In_84);
or U244 (N_244,In_352,In_17);
nor U245 (N_245,In_423,In_256);
xnor U246 (N_246,In_334,N_167);
and U247 (N_247,In_278,In_136);
xor U248 (N_248,In_243,In_316);
nor U249 (N_249,In_424,N_56);
nand U250 (N_250,In_387,In_323);
or U251 (N_251,In_241,In_413);
and U252 (N_252,In_337,N_30);
nor U253 (N_253,N_136,N_10);
and U254 (N_254,N_134,In_196);
and U255 (N_255,N_209,In_325);
nor U256 (N_256,N_68,N_195);
nand U257 (N_257,N_194,N_49);
and U258 (N_258,N_161,In_451);
or U259 (N_259,In_151,In_304);
and U260 (N_260,N_211,In_349);
and U261 (N_261,In_355,N_17);
and U262 (N_262,In_437,In_183);
nor U263 (N_263,N_188,In_404);
or U264 (N_264,In_321,N_213);
and U265 (N_265,N_240,In_305);
xor U266 (N_266,N_204,N_176);
or U267 (N_267,In_178,N_162);
or U268 (N_268,N_151,N_232);
and U269 (N_269,N_198,N_79);
or U270 (N_270,N_130,N_126);
or U271 (N_271,In_239,In_485);
xor U272 (N_272,In_83,N_243);
nor U273 (N_273,N_249,In_128);
nand U274 (N_274,In_97,N_235);
and U275 (N_275,N_241,In_44);
or U276 (N_276,In_154,N_152);
nand U277 (N_277,N_215,In_282);
or U278 (N_278,N_84,N_242);
or U279 (N_279,In_449,In_232);
or U280 (N_280,In_402,N_101);
and U281 (N_281,In_296,In_40);
nor U282 (N_282,N_31,N_246);
and U283 (N_283,N_202,In_210);
and U284 (N_284,In_341,N_158);
nor U285 (N_285,N_192,In_169);
and U286 (N_286,In_90,In_458);
nor U287 (N_287,N_98,In_339);
nand U288 (N_288,N_51,In_292);
or U289 (N_289,N_173,In_333);
and U290 (N_290,N_86,N_16);
xnor U291 (N_291,In_428,In_150);
nor U292 (N_292,N_178,N_102);
or U293 (N_293,In_74,N_227);
xnor U294 (N_294,In_371,N_184);
nor U295 (N_295,In_311,N_238);
nor U296 (N_296,N_233,N_168);
nor U297 (N_297,In_464,In_214);
nor U298 (N_298,In_204,N_175);
nor U299 (N_299,N_189,N_186);
and U300 (N_300,N_264,In_390);
or U301 (N_301,N_63,N_74);
nand U302 (N_302,N_44,N_277);
xnor U303 (N_303,N_269,N_45);
or U304 (N_304,N_208,N_123);
nor U305 (N_305,In_326,N_133);
nor U306 (N_306,In_78,N_299);
or U307 (N_307,N_212,N_257);
nor U308 (N_308,In_202,In_76);
nand U309 (N_309,N_11,N_19);
or U310 (N_310,N_141,N_97);
or U311 (N_311,In_446,N_214);
or U312 (N_312,N_224,N_295);
or U313 (N_313,In_238,N_171);
and U314 (N_314,N_105,In_253);
or U315 (N_315,N_293,In_235);
and U316 (N_316,N_292,N_92);
or U317 (N_317,N_262,N_266);
nor U318 (N_318,N_160,N_39);
or U319 (N_319,In_160,N_272);
and U320 (N_320,N_222,N_144);
nor U321 (N_321,N_260,N_291);
or U322 (N_322,N_279,N_285);
xor U323 (N_323,N_247,N_294);
nor U324 (N_324,In_92,N_50);
or U325 (N_325,N_163,N_297);
or U326 (N_326,N_137,In_417);
or U327 (N_327,N_256,N_142);
and U328 (N_328,N_157,In_200);
nand U329 (N_329,In_231,In_396);
or U330 (N_330,N_64,N_289);
or U331 (N_331,N_99,N_164);
and U332 (N_332,In_414,In_146);
or U333 (N_333,N_225,N_177);
nor U334 (N_334,N_252,N_221);
or U335 (N_335,N_263,In_96);
xor U336 (N_336,N_201,N_118);
or U337 (N_337,In_493,In_86);
or U338 (N_338,N_170,N_55);
and U339 (N_339,In_22,N_276);
nor U340 (N_340,N_298,In_218);
xor U341 (N_341,N_271,N_65);
nand U342 (N_342,N_255,N_216);
xnor U343 (N_343,N_124,N_275);
nand U344 (N_344,In_111,N_230);
and U345 (N_345,In_184,N_122);
nor U346 (N_346,N_245,N_218);
nand U347 (N_347,N_52,N_228);
or U348 (N_348,N_274,N_205);
or U349 (N_349,N_159,In_366);
or U350 (N_350,N_229,N_287);
and U351 (N_351,In_26,N_283);
nor U352 (N_352,N_223,N_231);
xor U353 (N_353,N_332,N_335);
nor U354 (N_354,N_301,N_67);
and U355 (N_355,In_298,N_111);
or U356 (N_356,N_191,N_270);
and U357 (N_357,N_267,In_463);
nor U358 (N_358,N_345,N_273);
nand U359 (N_359,N_203,N_282);
nand U360 (N_360,N_349,In_79);
or U361 (N_361,N_343,N_113);
and U362 (N_362,N_254,N_304);
nor U363 (N_363,N_303,N_324);
and U364 (N_364,N_325,N_114);
nand U365 (N_365,N_53,N_217);
nand U366 (N_366,N_69,In_277);
nand U367 (N_367,N_319,N_342);
nand U368 (N_368,N_336,N_210);
xor U369 (N_369,N_250,N_296);
and U370 (N_370,N_341,N_80);
or U371 (N_371,N_196,In_492);
or U372 (N_372,N_346,N_333);
nor U373 (N_373,N_0,In_152);
and U374 (N_374,N_331,N_348);
and U375 (N_375,N_15,In_433);
xor U376 (N_376,N_207,N_244);
nor U377 (N_377,In_157,In_478);
and U378 (N_378,N_339,N_305);
nor U379 (N_379,N_330,In_299);
or U380 (N_380,N_312,N_104);
nor U381 (N_381,N_81,N_147);
and U382 (N_382,N_236,N_259);
and U383 (N_383,In_206,N_309);
nand U384 (N_384,In_403,N_347);
nand U385 (N_385,N_239,N_334);
nand U386 (N_386,N_237,N_181);
or U387 (N_387,N_317,N_311);
nand U388 (N_388,N_308,N_313);
and U389 (N_389,N_226,N_220);
xnor U390 (N_390,N_310,N_280);
nor U391 (N_391,N_251,N_108);
nand U392 (N_392,In_309,In_440);
and U393 (N_393,N_265,N_321);
nor U394 (N_394,N_96,N_278);
nor U395 (N_395,N_314,N_131);
or U396 (N_396,N_326,In_479);
xnor U397 (N_397,N_284,N_300);
nand U398 (N_398,In_486,N_318);
and U399 (N_399,N_302,N_248);
or U400 (N_400,N_366,N_288);
nand U401 (N_401,N_367,N_383);
nand U402 (N_402,N_354,N_393);
nor U403 (N_403,N_386,N_365);
nor U404 (N_404,In_75,N_281);
nor U405 (N_405,N_327,N_61);
xnor U406 (N_406,N_307,N_315);
or U407 (N_407,N_379,N_350);
nand U408 (N_408,N_357,N_156);
nor U409 (N_409,N_322,N_375);
and U410 (N_410,N_395,N_286);
nor U411 (N_411,N_115,N_389);
or U412 (N_412,N_179,N_398);
nor U413 (N_413,N_153,N_234);
nand U414 (N_414,N_361,N_320);
and U415 (N_415,N_364,N_363);
nor U416 (N_416,N_382,N_370);
xor U417 (N_417,In_147,N_368);
nor U418 (N_418,N_394,In_442);
or U419 (N_419,N_200,N_392);
nor U420 (N_420,N_377,N_397);
and U421 (N_421,N_374,N_344);
and U422 (N_422,N_380,N_328);
nor U423 (N_423,N_329,N_359);
nor U424 (N_424,N_219,N_396);
nand U425 (N_425,N_362,N_206);
and U426 (N_426,N_388,N_384);
and U427 (N_427,N_316,N_340);
and U428 (N_428,N_369,N_100);
or U429 (N_429,N_372,N_358);
or U430 (N_430,N_261,N_42);
xnor U431 (N_431,In_400,N_373);
nand U432 (N_432,N_290,In_308);
or U433 (N_433,N_371,N_353);
or U434 (N_434,N_356,In_422);
nand U435 (N_435,N_306,N_381);
nand U436 (N_436,N_360,In_99);
nor U437 (N_437,N_391,In_448);
or U438 (N_438,N_169,N_390);
nand U439 (N_439,In_36,N_385);
nand U440 (N_440,In_141,N_12);
nand U441 (N_441,N_91,N_399);
or U442 (N_442,N_193,N_323);
and U443 (N_443,N_183,N_253);
nor U444 (N_444,N_338,In_498);
nand U445 (N_445,N_378,N_103);
or U446 (N_446,N_352,N_268);
nor U447 (N_447,N_351,N_376);
and U448 (N_448,N_355,N_337);
and U449 (N_449,N_387,N_258);
and U450 (N_450,N_441,N_418);
nand U451 (N_451,N_427,N_422);
and U452 (N_452,N_438,N_403);
and U453 (N_453,N_442,N_421);
and U454 (N_454,N_433,N_401);
xor U455 (N_455,N_449,N_426);
xnor U456 (N_456,N_439,N_434);
and U457 (N_457,N_443,N_416);
nor U458 (N_458,N_440,N_447);
nor U459 (N_459,N_400,N_425);
nand U460 (N_460,N_405,N_430);
xor U461 (N_461,N_431,N_412);
nand U462 (N_462,N_404,N_437);
nor U463 (N_463,N_406,N_429);
and U464 (N_464,N_435,N_402);
and U465 (N_465,N_446,N_423);
nand U466 (N_466,N_444,N_445);
and U467 (N_467,N_409,N_419);
xnor U468 (N_468,N_436,N_420);
or U469 (N_469,N_448,N_407);
nand U470 (N_470,N_413,N_417);
and U471 (N_471,N_410,N_411);
nor U472 (N_472,N_408,N_432);
nand U473 (N_473,N_414,N_415);
and U474 (N_474,N_424,N_428);
and U475 (N_475,N_409,N_420);
and U476 (N_476,N_433,N_436);
or U477 (N_477,N_420,N_418);
and U478 (N_478,N_408,N_418);
nand U479 (N_479,N_435,N_445);
xnor U480 (N_480,N_402,N_425);
xor U481 (N_481,N_404,N_442);
nor U482 (N_482,N_428,N_402);
nor U483 (N_483,N_423,N_436);
nand U484 (N_484,N_448,N_409);
or U485 (N_485,N_437,N_429);
nand U486 (N_486,N_443,N_412);
and U487 (N_487,N_444,N_431);
xor U488 (N_488,N_410,N_431);
and U489 (N_489,N_428,N_449);
or U490 (N_490,N_429,N_408);
xor U491 (N_491,N_449,N_421);
nor U492 (N_492,N_414,N_428);
nor U493 (N_493,N_413,N_433);
nor U494 (N_494,N_447,N_445);
nor U495 (N_495,N_431,N_448);
nor U496 (N_496,N_421,N_433);
nand U497 (N_497,N_447,N_414);
xnor U498 (N_498,N_439,N_420);
nand U499 (N_499,N_439,N_417);
nand U500 (N_500,N_483,N_465);
nand U501 (N_501,N_455,N_498);
or U502 (N_502,N_497,N_487);
and U503 (N_503,N_451,N_450);
nand U504 (N_504,N_493,N_469);
or U505 (N_505,N_452,N_476);
nand U506 (N_506,N_492,N_464);
or U507 (N_507,N_478,N_470);
or U508 (N_508,N_480,N_473);
or U509 (N_509,N_471,N_482);
nand U510 (N_510,N_467,N_490);
xor U511 (N_511,N_457,N_496);
nor U512 (N_512,N_499,N_484);
nand U513 (N_513,N_486,N_481);
nor U514 (N_514,N_485,N_459);
or U515 (N_515,N_454,N_453);
and U516 (N_516,N_489,N_461);
or U517 (N_517,N_456,N_495);
nor U518 (N_518,N_463,N_477);
nor U519 (N_519,N_460,N_466);
nand U520 (N_520,N_488,N_472);
nand U521 (N_521,N_475,N_479);
or U522 (N_522,N_474,N_494);
nand U523 (N_523,N_462,N_468);
nor U524 (N_524,N_491,N_458);
or U525 (N_525,N_471,N_486);
or U526 (N_526,N_480,N_460);
or U527 (N_527,N_451,N_478);
xor U528 (N_528,N_498,N_462);
or U529 (N_529,N_456,N_493);
and U530 (N_530,N_465,N_467);
and U531 (N_531,N_498,N_491);
or U532 (N_532,N_481,N_475);
and U533 (N_533,N_453,N_494);
nand U534 (N_534,N_493,N_460);
or U535 (N_535,N_468,N_459);
or U536 (N_536,N_484,N_450);
xnor U537 (N_537,N_491,N_474);
or U538 (N_538,N_461,N_471);
nor U539 (N_539,N_493,N_451);
or U540 (N_540,N_459,N_492);
nand U541 (N_541,N_499,N_494);
nand U542 (N_542,N_462,N_463);
xor U543 (N_543,N_471,N_490);
and U544 (N_544,N_473,N_459);
nor U545 (N_545,N_452,N_455);
xnor U546 (N_546,N_462,N_478);
xnor U547 (N_547,N_481,N_483);
or U548 (N_548,N_495,N_461);
xor U549 (N_549,N_451,N_476);
xor U550 (N_550,N_508,N_506);
or U551 (N_551,N_512,N_548);
nand U552 (N_552,N_526,N_531);
or U553 (N_553,N_510,N_537);
and U554 (N_554,N_545,N_502);
nand U555 (N_555,N_538,N_517);
nand U556 (N_556,N_500,N_521);
nor U557 (N_557,N_549,N_543);
or U558 (N_558,N_518,N_504);
nand U559 (N_559,N_507,N_528);
nor U560 (N_560,N_519,N_525);
and U561 (N_561,N_513,N_534);
nand U562 (N_562,N_501,N_532);
or U563 (N_563,N_515,N_544);
or U564 (N_564,N_514,N_527);
nor U565 (N_565,N_547,N_503);
xnor U566 (N_566,N_533,N_546);
nor U567 (N_567,N_530,N_516);
nor U568 (N_568,N_542,N_535);
or U569 (N_569,N_524,N_509);
and U570 (N_570,N_520,N_522);
and U571 (N_571,N_540,N_529);
nor U572 (N_572,N_505,N_539);
or U573 (N_573,N_523,N_536);
nor U574 (N_574,N_511,N_541);
nand U575 (N_575,N_527,N_542);
nor U576 (N_576,N_504,N_529);
nand U577 (N_577,N_549,N_534);
nand U578 (N_578,N_515,N_548);
nand U579 (N_579,N_517,N_541);
or U580 (N_580,N_518,N_522);
and U581 (N_581,N_500,N_509);
nand U582 (N_582,N_536,N_538);
nand U583 (N_583,N_522,N_549);
and U584 (N_584,N_537,N_506);
nor U585 (N_585,N_513,N_518);
nor U586 (N_586,N_543,N_501);
xnor U587 (N_587,N_529,N_535);
and U588 (N_588,N_518,N_536);
nor U589 (N_589,N_541,N_532);
nand U590 (N_590,N_500,N_536);
nand U591 (N_591,N_509,N_525);
nand U592 (N_592,N_528,N_543);
or U593 (N_593,N_538,N_523);
and U594 (N_594,N_517,N_526);
nand U595 (N_595,N_518,N_542);
and U596 (N_596,N_512,N_501);
and U597 (N_597,N_506,N_513);
and U598 (N_598,N_530,N_547);
nor U599 (N_599,N_548,N_501);
xor U600 (N_600,N_573,N_586);
and U601 (N_601,N_595,N_575);
and U602 (N_602,N_582,N_580);
or U603 (N_603,N_568,N_561);
or U604 (N_604,N_598,N_555);
or U605 (N_605,N_597,N_599);
xor U606 (N_606,N_590,N_557);
or U607 (N_607,N_566,N_594);
nor U608 (N_608,N_574,N_579);
xnor U609 (N_609,N_571,N_559);
nand U610 (N_610,N_591,N_572);
nand U611 (N_611,N_570,N_593);
nor U612 (N_612,N_558,N_576);
and U613 (N_613,N_584,N_553);
and U614 (N_614,N_592,N_551);
and U615 (N_615,N_583,N_564);
nor U616 (N_616,N_562,N_554);
or U617 (N_617,N_585,N_589);
xor U618 (N_618,N_588,N_569);
xnor U619 (N_619,N_567,N_556);
xnor U620 (N_620,N_587,N_563);
xnor U621 (N_621,N_596,N_560);
or U622 (N_622,N_565,N_552);
nor U623 (N_623,N_581,N_578);
or U624 (N_624,N_550,N_577);
nor U625 (N_625,N_556,N_584);
or U626 (N_626,N_581,N_565);
nand U627 (N_627,N_554,N_591);
xnor U628 (N_628,N_575,N_596);
nor U629 (N_629,N_566,N_565);
nor U630 (N_630,N_587,N_576);
nand U631 (N_631,N_568,N_555);
nor U632 (N_632,N_598,N_566);
nand U633 (N_633,N_592,N_574);
xor U634 (N_634,N_553,N_552);
or U635 (N_635,N_565,N_572);
or U636 (N_636,N_551,N_570);
and U637 (N_637,N_583,N_559);
or U638 (N_638,N_564,N_550);
nor U639 (N_639,N_595,N_588);
nor U640 (N_640,N_568,N_597);
and U641 (N_641,N_564,N_555);
xor U642 (N_642,N_559,N_564);
nand U643 (N_643,N_592,N_570);
nand U644 (N_644,N_586,N_553);
nand U645 (N_645,N_589,N_565);
nand U646 (N_646,N_591,N_567);
or U647 (N_647,N_554,N_571);
or U648 (N_648,N_550,N_581);
nor U649 (N_649,N_565,N_556);
and U650 (N_650,N_648,N_626);
nand U651 (N_651,N_623,N_621);
nand U652 (N_652,N_634,N_633);
xor U653 (N_653,N_610,N_612);
nand U654 (N_654,N_645,N_602);
or U655 (N_655,N_613,N_630);
nand U656 (N_656,N_609,N_608);
nor U657 (N_657,N_639,N_636);
or U658 (N_658,N_649,N_622);
or U659 (N_659,N_637,N_641);
nand U660 (N_660,N_625,N_604);
nor U661 (N_661,N_644,N_607);
nand U662 (N_662,N_638,N_640);
or U663 (N_663,N_642,N_616);
nor U664 (N_664,N_606,N_614);
or U665 (N_665,N_611,N_628);
xor U666 (N_666,N_615,N_635);
nor U667 (N_667,N_619,N_643);
nor U668 (N_668,N_600,N_603);
nand U669 (N_669,N_647,N_620);
or U670 (N_670,N_629,N_617);
and U671 (N_671,N_605,N_624);
nand U672 (N_672,N_627,N_618);
or U673 (N_673,N_601,N_631);
and U674 (N_674,N_632,N_646);
nor U675 (N_675,N_627,N_630);
nand U676 (N_676,N_615,N_612);
nor U677 (N_677,N_602,N_637);
nor U678 (N_678,N_628,N_624);
nand U679 (N_679,N_616,N_620);
and U680 (N_680,N_607,N_612);
or U681 (N_681,N_612,N_632);
or U682 (N_682,N_641,N_638);
nand U683 (N_683,N_612,N_634);
and U684 (N_684,N_611,N_642);
or U685 (N_685,N_631,N_642);
or U686 (N_686,N_623,N_640);
xor U687 (N_687,N_623,N_649);
nand U688 (N_688,N_619,N_623);
or U689 (N_689,N_611,N_624);
nor U690 (N_690,N_646,N_628);
and U691 (N_691,N_608,N_632);
xnor U692 (N_692,N_634,N_625);
and U693 (N_693,N_628,N_605);
xnor U694 (N_694,N_640,N_625);
nand U695 (N_695,N_634,N_604);
nand U696 (N_696,N_648,N_620);
and U697 (N_697,N_634,N_615);
nor U698 (N_698,N_606,N_601);
nor U699 (N_699,N_635,N_644);
or U700 (N_700,N_653,N_680);
nand U701 (N_701,N_692,N_675);
or U702 (N_702,N_693,N_697);
and U703 (N_703,N_658,N_696);
or U704 (N_704,N_672,N_682);
nor U705 (N_705,N_689,N_683);
and U706 (N_706,N_694,N_677);
and U707 (N_707,N_690,N_659);
and U708 (N_708,N_691,N_666);
nor U709 (N_709,N_685,N_674);
and U710 (N_710,N_655,N_676);
nor U711 (N_711,N_657,N_681);
nand U712 (N_712,N_687,N_652);
and U713 (N_713,N_662,N_684);
nor U714 (N_714,N_686,N_660);
nor U715 (N_715,N_695,N_656);
nand U716 (N_716,N_671,N_698);
or U717 (N_717,N_651,N_654);
nor U718 (N_718,N_679,N_667);
or U719 (N_719,N_673,N_664);
and U720 (N_720,N_665,N_661);
nor U721 (N_721,N_650,N_678);
or U722 (N_722,N_699,N_669);
nor U723 (N_723,N_668,N_670);
nand U724 (N_724,N_688,N_663);
xor U725 (N_725,N_656,N_670);
nand U726 (N_726,N_654,N_689);
xor U727 (N_727,N_664,N_683);
xnor U728 (N_728,N_694,N_680);
and U729 (N_729,N_650,N_686);
and U730 (N_730,N_685,N_652);
or U731 (N_731,N_654,N_678);
and U732 (N_732,N_694,N_670);
or U733 (N_733,N_655,N_695);
nor U734 (N_734,N_666,N_675);
nor U735 (N_735,N_661,N_670);
nor U736 (N_736,N_682,N_651);
or U737 (N_737,N_693,N_667);
xnor U738 (N_738,N_699,N_668);
nand U739 (N_739,N_674,N_683);
or U740 (N_740,N_677,N_688);
or U741 (N_741,N_656,N_685);
or U742 (N_742,N_650,N_690);
nor U743 (N_743,N_692,N_657);
and U744 (N_744,N_652,N_650);
nand U745 (N_745,N_666,N_683);
xnor U746 (N_746,N_669,N_664);
and U747 (N_747,N_677,N_685);
xnor U748 (N_748,N_676,N_692);
and U749 (N_749,N_654,N_673);
or U750 (N_750,N_716,N_711);
or U751 (N_751,N_728,N_722);
nand U752 (N_752,N_739,N_745);
nor U753 (N_753,N_726,N_707);
nand U754 (N_754,N_717,N_734);
nand U755 (N_755,N_708,N_703);
xor U756 (N_756,N_732,N_720);
nor U757 (N_757,N_741,N_747);
and U758 (N_758,N_710,N_737);
or U759 (N_759,N_719,N_733);
nand U760 (N_760,N_721,N_718);
or U761 (N_761,N_702,N_723);
nand U762 (N_762,N_700,N_749);
and U763 (N_763,N_738,N_748);
or U764 (N_764,N_731,N_742);
or U765 (N_765,N_715,N_725);
or U766 (N_766,N_713,N_709);
and U767 (N_767,N_735,N_743);
and U768 (N_768,N_746,N_724);
and U769 (N_769,N_712,N_706);
or U770 (N_770,N_729,N_744);
and U771 (N_771,N_704,N_705);
nor U772 (N_772,N_727,N_736);
or U773 (N_773,N_730,N_714);
nand U774 (N_774,N_740,N_701);
or U775 (N_775,N_742,N_734);
or U776 (N_776,N_749,N_739);
or U777 (N_777,N_746,N_743);
nor U778 (N_778,N_736,N_718);
nor U779 (N_779,N_707,N_747);
nand U780 (N_780,N_749,N_706);
nand U781 (N_781,N_736,N_700);
xor U782 (N_782,N_732,N_703);
xor U783 (N_783,N_701,N_707);
nand U784 (N_784,N_735,N_712);
or U785 (N_785,N_748,N_718);
and U786 (N_786,N_720,N_716);
and U787 (N_787,N_704,N_741);
nor U788 (N_788,N_728,N_704);
and U789 (N_789,N_709,N_701);
nand U790 (N_790,N_736,N_714);
nor U791 (N_791,N_731,N_716);
and U792 (N_792,N_733,N_716);
and U793 (N_793,N_731,N_748);
or U794 (N_794,N_728,N_725);
or U795 (N_795,N_742,N_706);
and U796 (N_796,N_739,N_715);
or U797 (N_797,N_725,N_703);
nor U798 (N_798,N_746,N_717);
and U799 (N_799,N_731,N_718);
nor U800 (N_800,N_755,N_769);
nor U801 (N_801,N_754,N_787);
nand U802 (N_802,N_773,N_760);
and U803 (N_803,N_782,N_774);
and U804 (N_804,N_776,N_753);
or U805 (N_805,N_770,N_777);
nor U806 (N_806,N_795,N_788);
xor U807 (N_807,N_772,N_771);
or U808 (N_808,N_768,N_765);
xor U809 (N_809,N_761,N_752);
and U810 (N_810,N_751,N_796);
and U811 (N_811,N_767,N_759);
or U812 (N_812,N_764,N_758);
and U813 (N_813,N_781,N_779);
nand U814 (N_814,N_798,N_757);
nand U815 (N_815,N_766,N_756);
nor U816 (N_816,N_763,N_784);
nor U817 (N_817,N_791,N_783);
xnor U818 (N_818,N_750,N_789);
nand U819 (N_819,N_775,N_797);
xor U820 (N_820,N_762,N_799);
nand U821 (N_821,N_785,N_793);
xor U822 (N_822,N_790,N_778);
and U823 (N_823,N_792,N_786);
nor U824 (N_824,N_794,N_780);
and U825 (N_825,N_754,N_777);
nor U826 (N_826,N_789,N_761);
and U827 (N_827,N_760,N_752);
nand U828 (N_828,N_773,N_761);
or U829 (N_829,N_755,N_780);
or U830 (N_830,N_778,N_799);
or U831 (N_831,N_774,N_780);
nand U832 (N_832,N_778,N_785);
nand U833 (N_833,N_790,N_751);
or U834 (N_834,N_778,N_767);
nand U835 (N_835,N_778,N_753);
nand U836 (N_836,N_771,N_766);
or U837 (N_837,N_785,N_762);
and U838 (N_838,N_762,N_763);
or U839 (N_839,N_771,N_788);
xor U840 (N_840,N_768,N_776);
and U841 (N_841,N_787,N_779);
xor U842 (N_842,N_752,N_774);
or U843 (N_843,N_779,N_796);
nor U844 (N_844,N_770,N_763);
nand U845 (N_845,N_772,N_769);
nand U846 (N_846,N_782,N_798);
nor U847 (N_847,N_761,N_775);
nor U848 (N_848,N_798,N_764);
and U849 (N_849,N_768,N_756);
nor U850 (N_850,N_838,N_814);
nor U851 (N_851,N_848,N_839);
and U852 (N_852,N_836,N_816);
nor U853 (N_853,N_807,N_826);
nor U854 (N_854,N_815,N_837);
and U855 (N_855,N_802,N_810);
nor U856 (N_856,N_833,N_813);
nand U857 (N_857,N_821,N_847);
and U858 (N_858,N_824,N_834);
nor U859 (N_859,N_846,N_849);
or U860 (N_860,N_844,N_841);
and U861 (N_861,N_830,N_800);
nand U862 (N_862,N_842,N_819);
nor U863 (N_863,N_809,N_806);
or U864 (N_864,N_805,N_840);
nand U865 (N_865,N_820,N_827);
and U866 (N_866,N_804,N_822);
nor U867 (N_867,N_825,N_801);
and U868 (N_868,N_808,N_817);
and U869 (N_869,N_835,N_831);
xnor U870 (N_870,N_845,N_832);
or U871 (N_871,N_803,N_823);
and U872 (N_872,N_828,N_829);
or U873 (N_873,N_843,N_812);
and U874 (N_874,N_811,N_818);
nand U875 (N_875,N_806,N_808);
nand U876 (N_876,N_832,N_808);
nand U877 (N_877,N_828,N_846);
or U878 (N_878,N_832,N_822);
xor U879 (N_879,N_847,N_846);
or U880 (N_880,N_827,N_816);
or U881 (N_881,N_828,N_820);
xnor U882 (N_882,N_818,N_829);
and U883 (N_883,N_823,N_843);
nor U884 (N_884,N_836,N_807);
nand U885 (N_885,N_838,N_800);
nand U886 (N_886,N_830,N_822);
or U887 (N_887,N_822,N_821);
or U888 (N_888,N_844,N_827);
or U889 (N_889,N_816,N_806);
or U890 (N_890,N_845,N_806);
nor U891 (N_891,N_821,N_836);
or U892 (N_892,N_835,N_830);
nand U893 (N_893,N_820,N_809);
or U894 (N_894,N_845,N_800);
nand U895 (N_895,N_841,N_805);
or U896 (N_896,N_817,N_846);
nand U897 (N_897,N_819,N_814);
nor U898 (N_898,N_802,N_814);
nand U899 (N_899,N_818,N_819);
xor U900 (N_900,N_853,N_878);
nand U901 (N_901,N_852,N_893);
and U902 (N_902,N_875,N_885);
xnor U903 (N_903,N_899,N_898);
nand U904 (N_904,N_865,N_870);
nor U905 (N_905,N_869,N_851);
and U906 (N_906,N_873,N_874);
or U907 (N_907,N_880,N_889);
and U908 (N_908,N_891,N_864);
and U909 (N_909,N_850,N_887);
nand U910 (N_910,N_882,N_890);
or U911 (N_911,N_867,N_895);
and U912 (N_912,N_866,N_860);
nand U913 (N_913,N_897,N_884);
nand U914 (N_914,N_868,N_859);
or U915 (N_915,N_888,N_857);
nand U916 (N_916,N_883,N_894);
nor U917 (N_917,N_879,N_892);
nand U918 (N_918,N_876,N_886);
nand U919 (N_919,N_896,N_871);
or U920 (N_920,N_877,N_863);
nand U921 (N_921,N_872,N_862);
and U922 (N_922,N_854,N_881);
nor U923 (N_923,N_855,N_861);
and U924 (N_924,N_858,N_856);
and U925 (N_925,N_894,N_855);
nor U926 (N_926,N_856,N_890);
or U927 (N_927,N_860,N_861);
and U928 (N_928,N_887,N_884);
and U929 (N_929,N_868,N_898);
nor U930 (N_930,N_871,N_876);
and U931 (N_931,N_850,N_851);
or U932 (N_932,N_899,N_858);
or U933 (N_933,N_882,N_891);
nand U934 (N_934,N_858,N_870);
nor U935 (N_935,N_863,N_876);
or U936 (N_936,N_862,N_882);
and U937 (N_937,N_870,N_880);
or U938 (N_938,N_876,N_864);
nor U939 (N_939,N_874,N_885);
and U940 (N_940,N_878,N_888);
nand U941 (N_941,N_875,N_883);
nor U942 (N_942,N_879,N_868);
xnor U943 (N_943,N_859,N_888);
nor U944 (N_944,N_882,N_868);
or U945 (N_945,N_883,N_878);
or U946 (N_946,N_868,N_892);
xor U947 (N_947,N_887,N_854);
or U948 (N_948,N_887,N_888);
and U949 (N_949,N_879,N_881);
and U950 (N_950,N_924,N_923);
and U951 (N_951,N_946,N_904);
and U952 (N_952,N_942,N_936);
nor U953 (N_953,N_913,N_908);
and U954 (N_954,N_945,N_939);
nand U955 (N_955,N_921,N_938);
and U956 (N_956,N_903,N_914);
nand U957 (N_957,N_920,N_933);
and U958 (N_958,N_944,N_912);
and U959 (N_959,N_948,N_909);
nand U960 (N_960,N_922,N_943);
nand U961 (N_961,N_925,N_931);
nor U962 (N_962,N_937,N_900);
xor U963 (N_963,N_947,N_917);
or U964 (N_964,N_934,N_902);
or U965 (N_965,N_919,N_907);
or U966 (N_966,N_901,N_910);
and U967 (N_967,N_935,N_928);
and U968 (N_968,N_915,N_932);
and U969 (N_969,N_906,N_930);
and U970 (N_970,N_929,N_949);
or U971 (N_971,N_940,N_918);
xnor U972 (N_972,N_905,N_941);
xor U973 (N_973,N_926,N_916);
or U974 (N_974,N_927,N_911);
xnor U975 (N_975,N_916,N_923);
nor U976 (N_976,N_929,N_937);
and U977 (N_977,N_909,N_908);
or U978 (N_978,N_947,N_944);
nor U979 (N_979,N_928,N_929);
and U980 (N_980,N_911,N_941);
and U981 (N_981,N_918,N_919);
nand U982 (N_982,N_933,N_926);
xnor U983 (N_983,N_922,N_910);
and U984 (N_984,N_933,N_927);
and U985 (N_985,N_930,N_948);
or U986 (N_986,N_904,N_909);
nand U987 (N_987,N_925,N_928);
or U988 (N_988,N_940,N_927);
nand U989 (N_989,N_942,N_934);
nor U990 (N_990,N_924,N_920);
or U991 (N_991,N_944,N_906);
nor U992 (N_992,N_911,N_916);
and U993 (N_993,N_911,N_914);
or U994 (N_994,N_928,N_937);
nor U995 (N_995,N_930,N_938);
nor U996 (N_996,N_902,N_927);
nand U997 (N_997,N_926,N_923);
nand U998 (N_998,N_908,N_901);
nor U999 (N_999,N_944,N_942);
nand U1000 (N_1000,N_962,N_988);
and U1001 (N_1001,N_956,N_989);
and U1002 (N_1002,N_986,N_992);
nand U1003 (N_1003,N_974,N_981);
nor U1004 (N_1004,N_983,N_982);
or U1005 (N_1005,N_995,N_967);
or U1006 (N_1006,N_964,N_961);
and U1007 (N_1007,N_978,N_994);
nand U1008 (N_1008,N_960,N_963);
nand U1009 (N_1009,N_951,N_998);
xor U1010 (N_1010,N_950,N_972);
and U1011 (N_1011,N_966,N_996);
xor U1012 (N_1012,N_990,N_984);
or U1013 (N_1013,N_952,N_977);
xor U1014 (N_1014,N_999,N_968);
nor U1015 (N_1015,N_959,N_975);
and U1016 (N_1016,N_973,N_991);
nor U1017 (N_1017,N_971,N_987);
nand U1018 (N_1018,N_953,N_969);
and U1019 (N_1019,N_957,N_979);
nor U1020 (N_1020,N_955,N_997);
or U1021 (N_1021,N_980,N_985);
nand U1022 (N_1022,N_970,N_965);
and U1023 (N_1023,N_958,N_993);
nor U1024 (N_1024,N_976,N_954);
xor U1025 (N_1025,N_952,N_989);
nand U1026 (N_1026,N_961,N_970);
nand U1027 (N_1027,N_974,N_970);
and U1028 (N_1028,N_968,N_967);
nand U1029 (N_1029,N_984,N_969);
and U1030 (N_1030,N_964,N_960);
nand U1031 (N_1031,N_969,N_970);
nor U1032 (N_1032,N_963,N_969);
nand U1033 (N_1033,N_964,N_969);
and U1034 (N_1034,N_982,N_956);
or U1035 (N_1035,N_992,N_975);
nor U1036 (N_1036,N_964,N_975);
and U1037 (N_1037,N_975,N_970);
and U1038 (N_1038,N_974,N_991);
nand U1039 (N_1039,N_997,N_999);
nor U1040 (N_1040,N_983,N_955);
and U1041 (N_1041,N_966,N_981);
and U1042 (N_1042,N_987,N_955);
and U1043 (N_1043,N_963,N_973);
nor U1044 (N_1044,N_961,N_966);
nand U1045 (N_1045,N_962,N_972);
and U1046 (N_1046,N_986,N_975);
and U1047 (N_1047,N_964,N_991);
nor U1048 (N_1048,N_960,N_966);
nor U1049 (N_1049,N_953,N_950);
and U1050 (N_1050,N_1010,N_1002);
nor U1051 (N_1051,N_1024,N_1019);
nand U1052 (N_1052,N_1034,N_1039);
and U1053 (N_1053,N_1022,N_1036);
and U1054 (N_1054,N_1044,N_1016);
xnor U1055 (N_1055,N_1001,N_1009);
nor U1056 (N_1056,N_1037,N_1032);
nand U1057 (N_1057,N_1003,N_1033);
and U1058 (N_1058,N_1047,N_1004);
or U1059 (N_1059,N_1020,N_1000);
or U1060 (N_1060,N_1005,N_1029);
or U1061 (N_1061,N_1025,N_1030);
or U1062 (N_1062,N_1006,N_1015);
and U1063 (N_1063,N_1028,N_1017);
and U1064 (N_1064,N_1048,N_1035);
or U1065 (N_1065,N_1011,N_1040);
and U1066 (N_1066,N_1012,N_1046);
nor U1067 (N_1067,N_1031,N_1027);
or U1068 (N_1068,N_1049,N_1045);
or U1069 (N_1069,N_1023,N_1021);
nor U1070 (N_1070,N_1018,N_1043);
and U1071 (N_1071,N_1042,N_1007);
or U1072 (N_1072,N_1013,N_1008);
nor U1073 (N_1073,N_1014,N_1038);
nand U1074 (N_1074,N_1041,N_1026);
nand U1075 (N_1075,N_1026,N_1049);
and U1076 (N_1076,N_1036,N_1037);
and U1077 (N_1077,N_1015,N_1017);
or U1078 (N_1078,N_1010,N_1014);
nand U1079 (N_1079,N_1039,N_1041);
or U1080 (N_1080,N_1030,N_1001);
nor U1081 (N_1081,N_1011,N_1031);
nand U1082 (N_1082,N_1043,N_1014);
nor U1083 (N_1083,N_1042,N_1027);
and U1084 (N_1084,N_1028,N_1003);
nor U1085 (N_1085,N_1035,N_1032);
nor U1086 (N_1086,N_1004,N_1008);
xor U1087 (N_1087,N_1011,N_1018);
nand U1088 (N_1088,N_1029,N_1037);
nand U1089 (N_1089,N_1024,N_1048);
and U1090 (N_1090,N_1039,N_1016);
nand U1091 (N_1091,N_1010,N_1046);
and U1092 (N_1092,N_1026,N_1030);
and U1093 (N_1093,N_1038,N_1043);
nand U1094 (N_1094,N_1048,N_1047);
nand U1095 (N_1095,N_1045,N_1003);
xnor U1096 (N_1096,N_1038,N_1046);
nand U1097 (N_1097,N_1011,N_1020);
or U1098 (N_1098,N_1039,N_1019);
nor U1099 (N_1099,N_1039,N_1023);
xnor U1100 (N_1100,N_1073,N_1068);
or U1101 (N_1101,N_1072,N_1061);
nand U1102 (N_1102,N_1094,N_1079);
or U1103 (N_1103,N_1075,N_1097);
nor U1104 (N_1104,N_1083,N_1089);
nor U1105 (N_1105,N_1057,N_1064);
and U1106 (N_1106,N_1086,N_1081);
or U1107 (N_1107,N_1058,N_1095);
nand U1108 (N_1108,N_1090,N_1066);
nor U1109 (N_1109,N_1078,N_1091);
and U1110 (N_1110,N_1050,N_1055);
nand U1111 (N_1111,N_1065,N_1070);
nor U1112 (N_1112,N_1092,N_1099);
nor U1113 (N_1113,N_1098,N_1059);
or U1114 (N_1114,N_1051,N_1074);
or U1115 (N_1115,N_1084,N_1054);
or U1116 (N_1116,N_1080,N_1088);
and U1117 (N_1117,N_1071,N_1063);
nand U1118 (N_1118,N_1053,N_1093);
or U1119 (N_1119,N_1077,N_1069);
and U1120 (N_1120,N_1056,N_1087);
xnor U1121 (N_1121,N_1076,N_1085);
nor U1122 (N_1122,N_1082,N_1062);
nor U1123 (N_1123,N_1060,N_1052);
or U1124 (N_1124,N_1067,N_1096);
or U1125 (N_1125,N_1054,N_1069);
or U1126 (N_1126,N_1077,N_1066);
nand U1127 (N_1127,N_1096,N_1064);
nand U1128 (N_1128,N_1075,N_1073);
and U1129 (N_1129,N_1069,N_1073);
or U1130 (N_1130,N_1076,N_1082);
nor U1131 (N_1131,N_1069,N_1081);
nor U1132 (N_1132,N_1091,N_1071);
and U1133 (N_1133,N_1094,N_1082);
nor U1134 (N_1134,N_1094,N_1057);
nor U1135 (N_1135,N_1092,N_1074);
nand U1136 (N_1136,N_1053,N_1064);
or U1137 (N_1137,N_1099,N_1065);
nor U1138 (N_1138,N_1087,N_1069);
nand U1139 (N_1139,N_1090,N_1055);
nor U1140 (N_1140,N_1077,N_1085);
and U1141 (N_1141,N_1073,N_1057);
or U1142 (N_1142,N_1074,N_1065);
nand U1143 (N_1143,N_1075,N_1061);
xor U1144 (N_1144,N_1085,N_1092);
nand U1145 (N_1145,N_1057,N_1069);
xnor U1146 (N_1146,N_1099,N_1074);
nand U1147 (N_1147,N_1078,N_1053);
or U1148 (N_1148,N_1077,N_1059);
nor U1149 (N_1149,N_1072,N_1086);
nor U1150 (N_1150,N_1117,N_1149);
and U1151 (N_1151,N_1141,N_1128);
nor U1152 (N_1152,N_1106,N_1148);
or U1153 (N_1153,N_1146,N_1107);
nand U1154 (N_1154,N_1124,N_1113);
or U1155 (N_1155,N_1108,N_1136);
and U1156 (N_1156,N_1143,N_1104);
and U1157 (N_1157,N_1119,N_1138);
nor U1158 (N_1158,N_1121,N_1134);
nor U1159 (N_1159,N_1116,N_1140);
nor U1160 (N_1160,N_1127,N_1142);
or U1161 (N_1161,N_1137,N_1133);
or U1162 (N_1162,N_1132,N_1145);
and U1163 (N_1163,N_1129,N_1131);
and U1164 (N_1164,N_1118,N_1130);
xor U1165 (N_1165,N_1125,N_1144);
or U1166 (N_1166,N_1126,N_1102);
nand U1167 (N_1167,N_1115,N_1111);
or U1168 (N_1168,N_1101,N_1105);
and U1169 (N_1169,N_1110,N_1147);
nor U1170 (N_1170,N_1120,N_1114);
or U1171 (N_1171,N_1100,N_1139);
xnor U1172 (N_1172,N_1122,N_1109);
or U1173 (N_1173,N_1123,N_1135);
and U1174 (N_1174,N_1112,N_1103);
nand U1175 (N_1175,N_1111,N_1126);
nand U1176 (N_1176,N_1103,N_1145);
nand U1177 (N_1177,N_1123,N_1107);
nand U1178 (N_1178,N_1138,N_1112);
nand U1179 (N_1179,N_1129,N_1130);
or U1180 (N_1180,N_1134,N_1140);
or U1181 (N_1181,N_1138,N_1135);
xnor U1182 (N_1182,N_1128,N_1131);
or U1183 (N_1183,N_1127,N_1120);
nor U1184 (N_1184,N_1121,N_1127);
or U1185 (N_1185,N_1147,N_1114);
xnor U1186 (N_1186,N_1132,N_1120);
and U1187 (N_1187,N_1132,N_1100);
or U1188 (N_1188,N_1108,N_1130);
or U1189 (N_1189,N_1121,N_1116);
xor U1190 (N_1190,N_1101,N_1126);
and U1191 (N_1191,N_1128,N_1121);
and U1192 (N_1192,N_1147,N_1132);
nand U1193 (N_1193,N_1104,N_1130);
nor U1194 (N_1194,N_1107,N_1124);
and U1195 (N_1195,N_1126,N_1143);
and U1196 (N_1196,N_1138,N_1139);
and U1197 (N_1197,N_1144,N_1145);
nor U1198 (N_1198,N_1120,N_1128);
nor U1199 (N_1199,N_1119,N_1117);
xor U1200 (N_1200,N_1158,N_1194);
or U1201 (N_1201,N_1155,N_1186);
or U1202 (N_1202,N_1189,N_1183);
or U1203 (N_1203,N_1157,N_1177);
xor U1204 (N_1204,N_1171,N_1175);
xor U1205 (N_1205,N_1153,N_1193);
nand U1206 (N_1206,N_1167,N_1184);
or U1207 (N_1207,N_1181,N_1163);
or U1208 (N_1208,N_1170,N_1162);
nor U1209 (N_1209,N_1169,N_1195);
nor U1210 (N_1210,N_1160,N_1187);
nand U1211 (N_1211,N_1159,N_1173);
nand U1212 (N_1212,N_1168,N_1179);
and U1213 (N_1213,N_1188,N_1190);
or U1214 (N_1214,N_1174,N_1182);
nor U1215 (N_1215,N_1192,N_1152);
or U1216 (N_1216,N_1164,N_1151);
and U1217 (N_1217,N_1154,N_1161);
nand U1218 (N_1218,N_1172,N_1199);
nor U1219 (N_1219,N_1198,N_1156);
nand U1220 (N_1220,N_1165,N_1197);
or U1221 (N_1221,N_1191,N_1166);
and U1222 (N_1222,N_1196,N_1185);
nand U1223 (N_1223,N_1150,N_1176);
or U1224 (N_1224,N_1180,N_1178);
nor U1225 (N_1225,N_1183,N_1170);
nor U1226 (N_1226,N_1175,N_1156);
nand U1227 (N_1227,N_1163,N_1174);
and U1228 (N_1228,N_1190,N_1176);
nor U1229 (N_1229,N_1152,N_1160);
nor U1230 (N_1230,N_1188,N_1169);
nand U1231 (N_1231,N_1164,N_1152);
nand U1232 (N_1232,N_1153,N_1150);
or U1233 (N_1233,N_1192,N_1164);
xor U1234 (N_1234,N_1168,N_1178);
nor U1235 (N_1235,N_1178,N_1161);
nand U1236 (N_1236,N_1171,N_1176);
nand U1237 (N_1237,N_1150,N_1178);
nand U1238 (N_1238,N_1160,N_1185);
and U1239 (N_1239,N_1182,N_1168);
or U1240 (N_1240,N_1182,N_1155);
nor U1241 (N_1241,N_1198,N_1174);
or U1242 (N_1242,N_1172,N_1187);
or U1243 (N_1243,N_1180,N_1163);
nand U1244 (N_1244,N_1176,N_1156);
nand U1245 (N_1245,N_1168,N_1189);
nand U1246 (N_1246,N_1184,N_1152);
nor U1247 (N_1247,N_1181,N_1180);
xnor U1248 (N_1248,N_1189,N_1171);
nor U1249 (N_1249,N_1159,N_1178);
or U1250 (N_1250,N_1233,N_1230);
or U1251 (N_1251,N_1229,N_1223);
or U1252 (N_1252,N_1226,N_1225);
nand U1253 (N_1253,N_1232,N_1219);
and U1254 (N_1254,N_1244,N_1222);
xnor U1255 (N_1255,N_1203,N_1205);
nor U1256 (N_1256,N_1211,N_1204);
xor U1257 (N_1257,N_1220,N_1201);
or U1258 (N_1258,N_1240,N_1242);
or U1259 (N_1259,N_1208,N_1200);
nand U1260 (N_1260,N_1218,N_1227);
nand U1261 (N_1261,N_1209,N_1207);
and U1262 (N_1262,N_1239,N_1231);
or U1263 (N_1263,N_1234,N_1247);
or U1264 (N_1264,N_1206,N_1241);
nor U1265 (N_1265,N_1224,N_1210);
nor U1266 (N_1266,N_1215,N_1214);
and U1267 (N_1267,N_1216,N_1202);
and U1268 (N_1268,N_1245,N_1217);
nor U1269 (N_1269,N_1237,N_1238);
or U1270 (N_1270,N_1236,N_1212);
nand U1271 (N_1271,N_1243,N_1235);
or U1272 (N_1272,N_1248,N_1246);
nor U1273 (N_1273,N_1228,N_1213);
and U1274 (N_1274,N_1221,N_1249);
or U1275 (N_1275,N_1219,N_1235);
or U1276 (N_1276,N_1202,N_1208);
nand U1277 (N_1277,N_1221,N_1245);
and U1278 (N_1278,N_1216,N_1247);
or U1279 (N_1279,N_1208,N_1224);
xor U1280 (N_1280,N_1242,N_1229);
xor U1281 (N_1281,N_1204,N_1227);
or U1282 (N_1282,N_1230,N_1208);
and U1283 (N_1283,N_1214,N_1228);
nand U1284 (N_1284,N_1243,N_1248);
nand U1285 (N_1285,N_1239,N_1205);
nor U1286 (N_1286,N_1248,N_1201);
or U1287 (N_1287,N_1221,N_1224);
nor U1288 (N_1288,N_1206,N_1238);
or U1289 (N_1289,N_1202,N_1238);
xor U1290 (N_1290,N_1219,N_1213);
and U1291 (N_1291,N_1246,N_1217);
or U1292 (N_1292,N_1220,N_1231);
xor U1293 (N_1293,N_1223,N_1235);
nand U1294 (N_1294,N_1222,N_1243);
nor U1295 (N_1295,N_1231,N_1224);
nor U1296 (N_1296,N_1216,N_1219);
nand U1297 (N_1297,N_1226,N_1227);
or U1298 (N_1298,N_1228,N_1234);
and U1299 (N_1299,N_1218,N_1231);
nor U1300 (N_1300,N_1297,N_1270);
and U1301 (N_1301,N_1298,N_1258);
nand U1302 (N_1302,N_1289,N_1268);
or U1303 (N_1303,N_1257,N_1277);
nor U1304 (N_1304,N_1259,N_1255);
nand U1305 (N_1305,N_1263,N_1287);
or U1306 (N_1306,N_1296,N_1251);
nand U1307 (N_1307,N_1285,N_1292);
nor U1308 (N_1308,N_1269,N_1282);
nand U1309 (N_1309,N_1275,N_1256);
and U1310 (N_1310,N_1286,N_1266);
or U1311 (N_1311,N_1284,N_1279);
and U1312 (N_1312,N_1272,N_1254);
nand U1313 (N_1313,N_1264,N_1280);
or U1314 (N_1314,N_1288,N_1291);
and U1315 (N_1315,N_1262,N_1299);
or U1316 (N_1316,N_1252,N_1294);
nor U1317 (N_1317,N_1265,N_1267);
nor U1318 (N_1318,N_1273,N_1250);
or U1319 (N_1319,N_1281,N_1271);
or U1320 (N_1320,N_1290,N_1261);
and U1321 (N_1321,N_1276,N_1295);
xnor U1322 (N_1322,N_1274,N_1260);
or U1323 (N_1323,N_1253,N_1293);
or U1324 (N_1324,N_1283,N_1278);
nand U1325 (N_1325,N_1266,N_1263);
xor U1326 (N_1326,N_1279,N_1280);
or U1327 (N_1327,N_1278,N_1284);
nand U1328 (N_1328,N_1292,N_1280);
and U1329 (N_1329,N_1298,N_1281);
and U1330 (N_1330,N_1296,N_1261);
xor U1331 (N_1331,N_1299,N_1261);
nor U1332 (N_1332,N_1273,N_1277);
xnor U1333 (N_1333,N_1281,N_1282);
nand U1334 (N_1334,N_1288,N_1261);
and U1335 (N_1335,N_1294,N_1267);
and U1336 (N_1336,N_1253,N_1276);
nand U1337 (N_1337,N_1290,N_1295);
nor U1338 (N_1338,N_1261,N_1284);
or U1339 (N_1339,N_1299,N_1256);
or U1340 (N_1340,N_1269,N_1250);
nand U1341 (N_1341,N_1285,N_1288);
or U1342 (N_1342,N_1257,N_1258);
or U1343 (N_1343,N_1269,N_1252);
nand U1344 (N_1344,N_1276,N_1262);
or U1345 (N_1345,N_1257,N_1295);
nand U1346 (N_1346,N_1266,N_1265);
nor U1347 (N_1347,N_1279,N_1285);
xnor U1348 (N_1348,N_1277,N_1266);
and U1349 (N_1349,N_1287,N_1284);
nand U1350 (N_1350,N_1347,N_1309);
nand U1351 (N_1351,N_1312,N_1343);
or U1352 (N_1352,N_1306,N_1331);
and U1353 (N_1353,N_1327,N_1319);
or U1354 (N_1354,N_1346,N_1333);
or U1355 (N_1355,N_1308,N_1305);
nor U1356 (N_1356,N_1338,N_1314);
nand U1357 (N_1357,N_1302,N_1301);
xor U1358 (N_1358,N_1320,N_1317);
or U1359 (N_1359,N_1307,N_1315);
or U1360 (N_1360,N_1325,N_1300);
nor U1361 (N_1361,N_1336,N_1334);
or U1362 (N_1362,N_1310,N_1329);
nor U1363 (N_1363,N_1326,N_1313);
or U1364 (N_1364,N_1349,N_1328);
nand U1365 (N_1365,N_1332,N_1324);
or U1366 (N_1366,N_1345,N_1344);
and U1367 (N_1367,N_1330,N_1318);
or U1368 (N_1368,N_1311,N_1341);
or U1369 (N_1369,N_1337,N_1303);
and U1370 (N_1370,N_1335,N_1342);
xor U1371 (N_1371,N_1323,N_1316);
nand U1372 (N_1372,N_1321,N_1304);
nand U1373 (N_1373,N_1322,N_1340);
nor U1374 (N_1374,N_1339,N_1348);
or U1375 (N_1375,N_1328,N_1318);
or U1376 (N_1376,N_1345,N_1328);
nand U1377 (N_1377,N_1325,N_1349);
nand U1378 (N_1378,N_1326,N_1328);
nand U1379 (N_1379,N_1325,N_1319);
xnor U1380 (N_1380,N_1300,N_1344);
nand U1381 (N_1381,N_1348,N_1330);
or U1382 (N_1382,N_1349,N_1336);
nand U1383 (N_1383,N_1341,N_1301);
and U1384 (N_1384,N_1320,N_1331);
nor U1385 (N_1385,N_1335,N_1319);
or U1386 (N_1386,N_1320,N_1323);
and U1387 (N_1387,N_1314,N_1329);
and U1388 (N_1388,N_1346,N_1342);
and U1389 (N_1389,N_1319,N_1331);
and U1390 (N_1390,N_1342,N_1331);
xnor U1391 (N_1391,N_1348,N_1304);
or U1392 (N_1392,N_1301,N_1326);
and U1393 (N_1393,N_1326,N_1322);
and U1394 (N_1394,N_1340,N_1323);
nor U1395 (N_1395,N_1307,N_1310);
xor U1396 (N_1396,N_1332,N_1319);
and U1397 (N_1397,N_1322,N_1315);
or U1398 (N_1398,N_1311,N_1302);
xor U1399 (N_1399,N_1322,N_1329);
nand U1400 (N_1400,N_1377,N_1354);
nand U1401 (N_1401,N_1365,N_1355);
or U1402 (N_1402,N_1375,N_1399);
or U1403 (N_1403,N_1385,N_1396);
xnor U1404 (N_1404,N_1384,N_1394);
nand U1405 (N_1405,N_1352,N_1368);
nand U1406 (N_1406,N_1380,N_1391);
nor U1407 (N_1407,N_1363,N_1398);
nand U1408 (N_1408,N_1361,N_1366);
or U1409 (N_1409,N_1357,N_1389);
nor U1410 (N_1410,N_1351,N_1392);
nor U1411 (N_1411,N_1358,N_1359);
xor U1412 (N_1412,N_1353,N_1371);
and U1413 (N_1413,N_1376,N_1390);
and U1414 (N_1414,N_1393,N_1397);
nor U1415 (N_1415,N_1370,N_1356);
and U1416 (N_1416,N_1387,N_1381);
nor U1417 (N_1417,N_1378,N_1364);
nand U1418 (N_1418,N_1388,N_1360);
nor U1419 (N_1419,N_1350,N_1395);
and U1420 (N_1420,N_1374,N_1369);
or U1421 (N_1421,N_1362,N_1379);
nand U1422 (N_1422,N_1373,N_1383);
or U1423 (N_1423,N_1386,N_1372);
nand U1424 (N_1424,N_1382,N_1367);
and U1425 (N_1425,N_1395,N_1370);
and U1426 (N_1426,N_1379,N_1355);
xnor U1427 (N_1427,N_1368,N_1353);
nor U1428 (N_1428,N_1395,N_1375);
or U1429 (N_1429,N_1356,N_1371);
and U1430 (N_1430,N_1385,N_1376);
nor U1431 (N_1431,N_1397,N_1399);
xnor U1432 (N_1432,N_1392,N_1379);
or U1433 (N_1433,N_1352,N_1372);
or U1434 (N_1434,N_1350,N_1352);
nand U1435 (N_1435,N_1399,N_1398);
nor U1436 (N_1436,N_1387,N_1357);
or U1437 (N_1437,N_1372,N_1380);
and U1438 (N_1438,N_1359,N_1382);
and U1439 (N_1439,N_1353,N_1351);
or U1440 (N_1440,N_1374,N_1356);
nand U1441 (N_1441,N_1398,N_1354);
nor U1442 (N_1442,N_1372,N_1371);
nor U1443 (N_1443,N_1399,N_1354);
nor U1444 (N_1444,N_1381,N_1378);
nor U1445 (N_1445,N_1372,N_1382);
nor U1446 (N_1446,N_1365,N_1387);
nor U1447 (N_1447,N_1354,N_1375);
and U1448 (N_1448,N_1352,N_1392);
and U1449 (N_1449,N_1391,N_1394);
or U1450 (N_1450,N_1440,N_1426);
or U1451 (N_1451,N_1415,N_1448);
nand U1452 (N_1452,N_1449,N_1401);
nand U1453 (N_1453,N_1400,N_1443);
or U1454 (N_1454,N_1421,N_1420);
nor U1455 (N_1455,N_1422,N_1434);
and U1456 (N_1456,N_1429,N_1445);
xnor U1457 (N_1457,N_1404,N_1431);
nor U1458 (N_1458,N_1444,N_1413);
nand U1459 (N_1459,N_1414,N_1433);
and U1460 (N_1460,N_1417,N_1405);
nand U1461 (N_1461,N_1439,N_1423);
and U1462 (N_1462,N_1424,N_1410);
nor U1463 (N_1463,N_1425,N_1416);
nor U1464 (N_1464,N_1402,N_1438);
and U1465 (N_1465,N_1427,N_1411);
and U1466 (N_1466,N_1428,N_1447);
nand U1467 (N_1467,N_1441,N_1435);
or U1468 (N_1468,N_1446,N_1408);
and U1469 (N_1469,N_1403,N_1419);
nand U1470 (N_1470,N_1436,N_1437);
or U1471 (N_1471,N_1406,N_1412);
xnor U1472 (N_1472,N_1418,N_1409);
xor U1473 (N_1473,N_1430,N_1442);
nor U1474 (N_1474,N_1407,N_1432);
or U1475 (N_1475,N_1411,N_1407);
and U1476 (N_1476,N_1428,N_1411);
nor U1477 (N_1477,N_1433,N_1423);
or U1478 (N_1478,N_1441,N_1407);
nor U1479 (N_1479,N_1428,N_1432);
nand U1480 (N_1480,N_1433,N_1417);
or U1481 (N_1481,N_1423,N_1401);
xor U1482 (N_1482,N_1425,N_1418);
nor U1483 (N_1483,N_1416,N_1431);
xnor U1484 (N_1484,N_1448,N_1438);
nand U1485 (N_1485,N_1447,N_1430);
nand U1486 (N_1486,N_1437,N_1441);
nor U1487 (N_1487,N_1434,N_1449);
nor U1488 (N_1488,N_1404,N_1408);
nor U1489 (N_1489,N_1435,N_1431);
or U1490 (N_1490,N_1422,N_1420);
and U1491 (N_1491,N_1404,N_1406);
nand U1492 (N_1492,N_1433,N_1427);
xor U1493 (N_1493,N_1404,N_1419);
nor U1494 (N_1494,N_1426,N_1438);
nand U1495 (N_1495,N_1421,N_1433);
and U1496 (N_1496,N_1416,N_1403);
nor U1497 (N_1497,N_1446,N_1417);
xor U1498 (N_1498,N_1437,N_1420);
xnor U1499 (N_1499,N_1414,N_1429);
and U1500 (N_1500,N_1489,N_1493);
and U1501 (N_1501,N_1498,N_1499);
or U1502 (N_1502,N_1484,N_1474);
or U1503 (N_1503,N_1466,N_1453);
nor U1504 (N_1504,N_1462,N_1496);
nand U1505 (N_1505,N_1480,N_1457);
nor U1506 (N_1506,N_1476,N_1471);
or U1507 (N_1507,N_1454,N_1488);
or U1508 (N_1508,N_1468,N_1495);
nor U1509 (N_1509,N_1491,N_1452);
or U1510 (N_1510,N_1473,N_1475);
or U1511 (N_1511,N_1450,N_1463);
and U1512 (N_1512,N_1479,N_1464);
nand U1513 (N_1513,N_1478,N_1460);
nor U1514 (N_1514,N_1459,N_1458);
nor U1515 (N_1515,N_1477,N_1451);
nand U1516 (N_1516,N_1481,N_1470);
nor U1517 (N_1517,N_1467,N_1465);
or U1518 (N_1518,N_1497,N_1494);
nor U1519 (N_1519,N_1482,N_1486);
or U1520 (N_1520,N_1461,N_1455);
or U1521 (N_1521,N_1469,N_1485);
nor U1522 (N_1522,N_1492,N_1472);
nand U1523 (N_1523,N_1456,N_1483);
nand U1524 (N_1524,N_1490,N_1487);
and U1525 (N_1525,N_1455,N_1495);
or U1526 (N_1526,N_1497,N_1487);
or U1527 (N_1527,N_1451,N_1463);
nor U1528 (N_1528,N_1464,N_1459);
nand U1529 (N_1529,N_1493,N_1458);
or U1530 (N_1530,N_1460,N_1472);
xor U1531 (N_1531,N_1451,N_1462);
or U1532 (N_1532,N_1459,N_1493);
or U1533 (N_1533,N_1462,N_1463);
nor U1534 (N_1534,N_1490,N_1474);
and U1535 (N_1535,N_1468,N_1496);
xnor U1536 (N_1536,N_1463,N_1490);
and U1537 (N_1537,N_1499,N_1460);
and U1538 (N_1538,N_1451,N_1494);
and U1539 (N_1539,N_1464,N_1460);
nor U1540 (N_1540,N_1495,N_1465);
or U1541 (N_1541,N_1475,N_1491);
xnor U1542 (N_1542,N_1494,N_1465);
nor U1543 (N_1543,N_1486,N_1496);
nor U1544 (N_1544,N_1491,N_1472);
nor U1545 (N_1545,N_1461,N_1479);
or U1546 (N_1546,N_1483,N_1454);
and U1547 (N_1547,N_1451,N_1496);
xnor U1548 (N_1548,N_1475,N_1453);
or U1549 (N_1549,N_1458,N_1457);
and U1550 (N_1550,N_1502,N_1542);
nand U1551 (N_1551,N_1538,N_1507);
nor U1552 (N_1552,N_1522,N_1535);
nor U1553 (N_1553,N_1521,N_1524);
and U1554 (N_1554,N_1548,N_1503);
and U1555 (N_1555,N_1516,N_1529);
nand U1556 (N_1556,N_1540,N_1518);
and U1557 (N_1557,N_1517,N_1539);
and U1558 (N_1558,N_1505,N_1547);
and U1559 (N_1559,N_1501,N_1541);
nand U1560 (N_1560,N_1536,N_1512);
nand U1561 (N_1561,N_1549,N_1526);
nor U1562 (N_1562,N_1515,N_1506);
nand U1563 (N_1563,N_1523,N_1509);
xnor U1564 (N_1564,N_1533,N_1510);
or U1565 (N_1565,N_1520,N_1528);
xor U1566 (N_1566,N_1500,N_1525);
nand U1567 (N_1567,N_1532,N_1545);
or U1568 (N_1568,N_1527,N_1537);
nor U1569 (N_1569,N_1530,N_1543);
nor U1570 (N_1570,N_1546,N_1519);
or U1571 (N_1571,N_1544,N_1514);
xor U1572 (N_1572,N_1508,N_1513);
xnor U1573 (N_1573,N_1531,N_1534);
and U1574 (N_1574,N_1511,N_1504);
and U1575 (N_1575,N_1522,N_1546);
nand U1576 (N_1576,N_1500,N_1519);
nand U1577 (N_1577,N_1508,N_1545);
nand U1578 (N_1578,N_1546,N_1529);
nand U1579 (N_1579,N_1530,N_1537);
or U1580 (N_1580,N_1531,N_1547);
nor U1581 (N_1581,N_1543,N_1503);
or U1582 (N_1582,N_1523,N_1537);
nand U1583 (N_1583,N_1544,N_1545);
and U1584 (N_1584,N_1531,N_1502);
xnor U1585 (N_1585,N_1510,N_1530);
or U1586 (N_1586,N_1515,N_1537);
nand U1587 (N_1587,N_1516,N_1524);
xnor U1588 (N_1588,N_1526,N_1516);
and U1589 (N_1589,N_1545,N_1513);
or U1590 (N_1590,N_1517,N_1536);
nand U1591 (N_1591,N_1538,N_1519);
or U1592 (N_1592,N_1549,N_1519);
and U1593 (N_1593,N_1514,N_1519);
nand U1594 (N_1594,N_1547,N_1546);
nor U1595 (N_1595,N_1539,N_1512);
and U1596 (N_1596,N_1547,N_1537);
nand U1597 (N_1597,N_1520,N_1508);
or U1598 (N_1598,N_1517,N_1541);
and U1599 (N_1599,N_1517,N_1531);
or U1600 (N_1600,N_1560,N_1586);
or U1601 (N_1601,N_1552,N_1550);
nor U1602 (N_1602,N_1562,N_1554);
and U1603 (N_1603,N_1565,N_1585);
nand U1604 (N_1604,N_1580,N_1551);
or U1605 (N_1605,N_1587,N_1564);
or U1606 (N_1606,N_1574,N_1573);
xor U1607 (N_1607,N_1572,N_1569);
nor U1608 (N_1608,N_1584,N_1567);
or U1609 (N_1609,N_1591,N_1563);
and U1610 (N_1610,N_1557,N_1579);
or U1611 (N_1611,N_1553,N_1568);
nand U1612 (N_1612,N_1556,N_1596);
and U1613 (N_1613,N_1576,N_1582);
and U1614 (N_1614,N_1597,N_1555);
nand U1615 (N_1615,N_1598,N_1592);
and U1616 (N_1616,N_1590,N_1571);
and U1617 (N_1617,N_1588,N_1583);
nand U1618 (N_1618,N_1593,N_1575);
or U1619 (N_1619,N_1581,N_1559);
and U1620 (N_1620,N_1561,N_1578);
and U1621 (N_1621,N_1595,N_1570);
nand U1622 (N_1622,N_1558,N_1589);
or U1623 (N_1623,N_1594,N_1599);
nand U1624 (N_1624,N_1566,N_1577);
nor U1625 (N_1625,N_1558,N_1591);
nor U1626 (N_1626,N_1592,N_1594);
nand U1627 (N_1627,N_1572,N_1562);
and U1628 (N_1628,N_1555,N_1598);
nor U1629 (N_1629,N_1551,N_1577);
nand U1630 (N_1630,N_1578,N_1583);
nand U1631 (N_1631,N_1598,N_1574);
or U1632 (N_1632,N_1582,N_1573);
nand U1633 (N_1633,N_1583,N_1577);
and U1634 (N_1634,N_1562,N_1590);
or U1635 (N_1635,N_1588,N_1567);
nor U1636 (N_1636,N_1598,N_1587);
xnor U1637 (N_1637,N_1557,N_1574);
and U1638 (N_1638,N_1593,N_1562);
and U1639 (N_1639,N_1585,N_1588);
nand U1640 (N_1640,N_1588,N_1566);
nor U1641 (N_1641,N_1575,N_1597);
and U1642 (N_1642,N_1597,N_1589);
or U1643 (N_1643,N_1584,N_1591);
xor U1644 (N_1644,N_1599,N_1597);
and U1645 (N_1645,N_1595,N_1577);
or U1646 (N_1646,N_1568,N_1585);
and U1647 (N_1647,N_1565,N_1556);
and U1648 (N_1648,N_1599,N_1566);
nand U1649 (N_1649,N_1586,N_1598);
and U1650 (N_1650,N_1611,N_1620);
nand U1651 (N_1651,N_1631,N_1619);
or U1652 (N_1652,N_1630,N_1616);
xnor U1653 (N_1653,N_1608,N_1639);
or U1654 (N_1654,N_1626,N_1621);
nor U1655 (N_1655,N_1636,N_1622);
or U1656 (N_1656,N_1640,N_1642);
nand U1657 (N_1657,N_1644,N_1646);
and U1658 (N_1658,N_1605,N_1629);
nor U1659 (N_1659,N_1632,N_1618);
and U1660 (N_1660,N_1614,N_1623);
and U1661 (N_1661,N_1613,N_1635);
nor U1662 (N_1662,N_1638,N_1625);
and U1663 (N_1663,N_1606,N_1602);
nand U1664 (N_1664,N_1643,N_1607);
nor U1665 (N_1665,N_1624,N_1634);
nor U1666 (N_1666,N_1601,N_1641);
nand U1667 (N_1667,N_1648,N_1609);
or U1668 (N_1668,N_1633,N_1612);
xor U1669 (N_1669,N_1627,N_1628);
and U1670 (N_1670,N_1604,N_1647);
nand U1671 (N_1671,N_1645,N_1617);
nand U1672 (N_1672,N_1600,N_1603);
nand U1673 (N_1673,N_1615,N_1637);
nor U1674 (N_1674,N_1649,N_1610);
nor U1675 (N_1675,N_1641,N_1614);
or U1676 (N_1676,N_1631,N_1641);
and U1677 (N_1677,N_1643,N_1602);
and U1678 (N_1678,N_1604,N_1623);
xor U1679 (N_1679,N_1614,N_1615);
nand U1680 (N_1680,N_1614,N_1620);
or U1681 (N_1681,N_1611,N_1623);
xnor U1682 (N_1682,N_1621,N_1642);
xnor U1683 (N_1683,N_1603,N_1619);
or U1684 (N_1684,N_1630,N_1610);
nor U1685 (N_1685,N_1601,N_1600);
xnor U1686 (N_1686,N_1621,N_1624);
xnor U1687 (N_1687,N_1611,N_1628);
xnor U1688 (N_1688,N_1612,N_1604);
nor U1689 (N_1689,N_1626,N_1623);
or U1690 (N_1690,N_1612,N_1603);
nor U1691 (N_1691,N_1637,N_1626);
nand U1692 (N_1692,N_1636,N_1629);
or U1693 (N_1693,N_1641,N_1638);
or U1694 (N_1694,N_1618,N_1645);
or U1695 (N_1695,N_1638,N_1616);
nor U1696 (N_1696,N_1609,N_1608);
or U1697 (N_1697,N_1600,N_1640);
or U1698 (N_1698,N_1643,N_1629);
and U1699 (N_1699,N_1643,N_1646);
nand U1700 (N_1700,N_1660,N_1696);
or U1701 (N_1701,N_1659,N_1693);
nand U1702 (N_1702,N_1682,N_1699);
nor U1703 (N_1703,N_1684,N_1652);
nor U1704 (N_1704,N_1677,N_1692);
and U1705 (N_1705,N_1686,N_1663);
and U1706 (N_1706,N_1683,N_1678);
nand U1707 (N_1707,N_1689,N_1695);
or U1708 (N_1708,N_1657,N_1674);
nor U1709 (N_1709,N_1673,N_1688);
nand U1710 (N_1710,N_1681,N_1654);
and U1711 (N_1711,N_1680,N_1666);
nand U1712 (N_1712,N_1658,N_1690);
nor U1713 (N_1713,N_1656,N_1668);
or U1714 (N_1714,N_1665,N_1698);
and U1715 (N_1715,N_1653,N_1671);
nor U1716 (N_1716,N_1669,N_1697);
xor U1717 (N_1717,N_1672,N_1662);
and U1718 (N_1718,N_1676,N_1667);
or U1719 (N_1719,N_1664,N_1675);
or U1720 (N_1720,N_1685,N_1655);
and U1721 (N_1721,N_1691,N_1650);
and U1722 (N_1722,N_1687,N_1694);
nand U1723 (N_1723,N_1661,N_1670);
and U1724 (N_1724,N_1679,N_1651);
nand U1725 (N_1725,N_1693,N_1669);
or U1726 (N_1726,N_1660,N_1654);
and U1727 (N_1727,N_1655,N_1679);
xnor U1728 (N_1728,N_1683,N_1691);
nor U1729 (N_1729,N_1663,N_1674);
nor U1730 (N_1730,N_1671,N_1650);
or U1731 (N_1731,N_1659,N_1668);
nand U1732 (N_1732,N_1678,N_1694);
or U1733 (N_1733,N_1667,N_1690);
nand U1734 (N_1734,N_1697,N_1680);
xor U1735 (N_1735,N_1695,N_1687);
nand U1736 (N_1736,N_1679,N_1665);
and U1737 (N_1737,N_1677,N_1679);
or U1738 (N_1738,N_1670,N_1689);
and U1739 (N_1739,N_1682,N_1692);
or U1740 (N_1740,N_1671,N_1660);
or U1741 (N_1741,N_1664,N_1696);
and U1742 (N_1742,N_1652,N_1682);
and U1743 (N_1743,N_1657,N_1698);
nor U1744 (N_1744,N_1688,N_1690);
or U1745 (N_1745,N_1661,N_1654);
or U1746 (N_1746,N_1681,N_1659);
nand U1747 (N_1747,N_1662,N_1654);
or U1748 (N_1748,N_1683,N_1693);
nand U1749 (N_1749,N_1681,N_1651);
nor U1750 (N_1750,N_1724,N_1722);
nor U1751 (N_1751,N_1738,N_1720);
or U1752 (N_1752,N_1742,N_1711);
nand U1753 (N_1753,N_1740,N_1739);
nor U1754 (N_1754,N_1716,N_1730);
and U1755 (N_1755,N_1732,N_1706);
nor U1756 (N_1756,N_1744,N_1712);
nand U1757 (N_1757,N_1714,N_1709);
or U1758 (N_1758,N_1704,N_1705);
nand U1759 (N_1759,N_1715,N_1719);
nand U1760 (N_1760,N_1701,N_1726);
nand U1761 (N_1761,N_1735,N_1746);
nor U1762 (N_1762,N_1736,N_1728);
nand U1763 (N_1763,N_1710,N_1708);
nand U1764 (N_1764,N_1723,N_1745);
or U1765 (N_1765,N_1734,N_1748);
nor U1766 (N_1766,N_1703,N_1737);
nand U1767 (N_1767,N_1733,N_1727);
or U1768 (N_1768,N_1749,N_1743);
nor U1769 (N_1769,N_1700,N_1717);
nor U1770 (N_1770,N_1725,N_1718);
nand U1771 (N_1771,N_1741,N_1731);
nor U1772 (N_1772,N_1702,N_1707);
or U1773 (N_1773,N_1713,N_1729);
nand U1774 (N_1774,N_1721,N_1747);
nor U1775 (N_1775,N_1734,N_1718);
nand U1776 (N_1776,N_1744,N_1717);
nor U1777 (N_1777,N_1704,N_1739);
nor U1778 (N_1778,N_1741,N_1712);
or U1779 (N_1779,N_1748,N_1732);
and U1780 (N_1780,N_1702,N_1741);
or U1781 (N_1781,N_1743,N_1720);
xor U1782 (N_1782,N_1719,N_1730);
nor U1783 (N_1783,N_1735,N_1704);
nor U1784 (N_1784,N_1722,N_1705);
nor U1785 (N_1785,N_1708,N_1721);
or U1786 (N_1786,N_1728,N_1742);
nor U1787 (N_1787,N_1725,N_1742);
nand U1788 (N_1788,N_1717,N_1738);
and U1789 (N_1789,N_1748,N_1704);
nand U1790 (N_1790,N_1727,N_1705);
and U1791 (N_1791,N_1746,N_1744);
nor U1792 (N_1792,N_1739,N_1713);
nand U1793 (N_1793,N_1745,N_1707);
and U1794 (N_1794,N_1709,N_1740);
nand U1795 (N_1795,N_1706,N_1748);
or U1796 (N_1796,N_1733,N_1740);
nor U1797 (N_1797,N_1710,N_1718);
or U1798 (N_1798,N_1709,N_1719);
xnor U1799 (N_1799,N_1702,N_1745);
nor U1800 (N_1800,N_1788,N_1750);
xnor U1801 (N_1801,N_1789,N_1774);
nor U1802 (N_1802,N_1777,N_1759);
or U1803 (N_1803,N_1781,N_1798);
or U1804 (N_1804,N_1796,N_1764);
nand U1805 (N_1805,N_1770,N_1756);
nor U1806 (N_1806,N_1799,N_1773);
and U1807 (N_1807,N_1758,N_1790);
and U1808 (N_1808,N_1780,N_1787);
nor U1809 (N_1809,N_1775,N_1782);
or U1810 (N_1810,N_1754,N_1783);
and U1811 (N_1811,N_1761,N_1795);
and U1812 (N_1812,N_1769,N_1786);
nor U1813 (N_1813,N_1765,N_1793);
nor U1814 (N_1814,N_1763,N_1766);
nor U1815 (N_1815,N_1755,N_1753);
or U1816 (N_1816,N_1767,N_1760);
nand U1817 (N_1817,N_1772,N_1776);
nor U1818 (N_1818,N_1779,N_1792);
nor U1819 (N_1819,N_1784,N_1751);
or U1820 (N_1820,N_1791,N_1771);
nand U1821 (N_1821,N_1778,N_1797);
or U1822 (N_1822,N_1768,N_1794);
nor U1823 (N_1823,N_1757,N_1752);
and U1824 (N_1824,N_1785,N_1762);
nand U1825 (N_1825,N_1781,N_1791);
and U1826 (N_1826,N_1794,N_1760);
and U1827 (N_1827,N_1794,N_1767);
xor U1828 (N_1828,N_1753,N_1765);
and U1829 (N_1829,N_1766,N_1783);
and U1830 (N_1830,N_1795,N_1794);
nand U1831 (N_1831,N_1776,N_1754);
or U1832 (N_1832,N_1750,N_1755);
nor U1833 (N_1833,N_1755,N_1777);
or U1834 (N_1834,N_1750,N_1762);
nand U1835 (N_1835,N_1781,N_1751);
and U1836 (N_1836,N_1779,N_1761);
and U1837 (N_1837,N_1779,N_1754);
nand U1838 (N_1838,N_1766,N_1768);
nand U1839 (N_1839,N_1778,N_1789);
or U1840 (N_1840,N_1799,N_1790);
xor U1841 (N_1841,N_1787,N_1770);
or U1842 (N_1842,N_1799,N_1780);
and U1843 (N_1843,N_1754,N_1784);
or U1844 (N_1844,N_1790,N_1798);
xnor U1845 (N_1845,N_1787,N_1756);
and U1846 (N_1846,N_1783,N_1781);
nor U1847 (N_1847,N_1756,N_1774);
xnor U1848 (N_1848,N_1780,N_1763);
and U1849 (N_1849,N_1791,N_1766);
or U1850 (N_1850,N_1817,N_1818);
nand U1851 (N_1851,N_1833,N_1809);
nand U1852 (N_1852,N_1839,N_1838);
and U1853 (N_1853,N_1831,N_1848);
nand U1854 (N_1854,N_1843,N_1846);
nor U1855 (N_1855,N_1805,N_1812);
nor U1856 (N_1856,N_1822,N_1814);
nand U1857 (N_1857,N_1824,N_1813);
and U1858 (N_1858,N_1832,N_1802);
and U1859 (N_1859,N_1845,N_1835);
xnor U1860 (N_1860,N_1841,N_1801);
nor U1861 (N_1861,N_1811,N_1826);
and U1862 (N_1862,N_1800,N_1815);
nand U1863 (N_1863,N_1840,N_1834);
nor U1864 (N_1864,N_1844,N_1808);
or U1865 (N_1865,N_1806,N_1829);
nand U1866 (N_1866,N_1820,N_1836);
and U1867 (N_1867,N_1842,N_1803);
nand U1868 (N_1868,N_1849,N_1804);
nand U1869 (N_1869,N_1847,N_1825);
nand U1870 (N_1870,N_1823,N_1821);
or U1871 (N_1871,N_1830,N_1828);
and U1872 (N_1872,N_1807,N_1819);
xor U1873 (N_1873,N_1816,N_1827);
and U1874 (N_1874,N_1837,N_1810);
xnor U1875 (N_1875,N_1818,N_1826);
or U1876 (N_1876,N_1828,N_1823);
or U1877 (N_1877,N_1835,N_1836);
or U1878 (N_1878,N_1803,N_1846);
or U1879 (N_1879,N_1838,N_1844);
nor U1880 (N_1880,N_1801,N_1802);
and U1881 (N_1881,N_1810,N_1836);
nor U1882 (N_1882,N_1849,N_1818);
and U1883 (N_1883,N_1848,N_1830);
and U1884 (N_1884,N_1810,N_1815);
xnor U1885 (N_1885,N_1829,N_1812);
xor U1886 (N_1886,N_1814,N_1838);
xor U1887 (N_1887,N_1849,N_1845);
and U1888 (N_1888,N_1843,N_1832);
xnor U1889 (N_1889,N_1809,N_1820);
nand U1890 (N_1890,N_1843,N_1809);
nor U1891 (N_1891,N_1812,N_1823);
or U1892 (N_1892,N_1825,N_1808);
and U1893 (N_1893,N_1840,N_1825);
and U1894 (N_1894,N_1800,N_1834);
and U1895 (N_1895,N_1803,N_1811);
and U1896 (N_1896,N_1826,N_1802);
or U1897 (N_1897,N_1843,N_1812);
and U1898 (N_1898,N_1823,N_1826);
and U1899 (N_1899,N_1814,N_1834);
nand U1900 (N_1900,N_1883,N_1861);
nor U1901 (N_1901,N_1889,N_1891);
and U1902 (N_1902,N_1873,N_1871);
nor U1903 (N_1903,N_1879,N_1864);
nand U1904 (N_1904,N_1850,N_1869);
nand U1905 (N_1905,N_1888,N_1868);
nor U1906 (N_1906,N_1886,N_1867);
and U1907 (N_1907,N_1874,N_1866);
nand U1908 (N_1908,N_1855,N_1892);
nand U1909 (N_1909,N_1897,N_1858);
nand U1910 (N_1910,N_1881,N_1857);
xor U1911 (N_1911,N_1893,N_1876);
and U1912 (N_1912,N_1862,N_1865);
or U1913 (N_1913,N_1887,N_1894);
or U1914 (N_1914,N_1884,N_1896);
nand U1915 (N_1915,N_1860,N_1875);
nor U1916 (N_1916,N_1853,N_1880);
or U1917 (N_1917,N_1870,N_1872);
or U1918 (N_1918,N_1890,N_1852);
and U1919 (N_1919,N_1898,N_1878);
or U1920 (N_1920,N_1863,N_1854);
or U1921 (N_1921,N_1877,N_1851);
nand U1922 (N_1922,N_1885,N_1882);
or U1923 (N_1923,N_1895,N_1899);
and U1924 (N_1924,N_1856,N_1859);
nor U1925 (N_1925,N_1884,N_1870);
nor U1926 (N_1926,N_1862,N_1875);
and U1927 (N_1927,N_1895,N_1853);
nand U1928 (N_1928,N_1865,N_1851);
nor U1929 (N_1929,N_1888,N_1877);
or U1930 (N_1930,N_1884,N_1895);
nor U1931 (N_1931,N_1851,N_1898);
and U1932 (N_1932,N_1855,N_1877);
nand U1933 (N_1933,N_1883,N_1866);
nor U1934 (N_1934,N_1865,N_1894);
and U1935 (N_1935,N_1880,N_1870);
xor U1936 (N_1936,N_1851,N_1882);
or U1937 (N_1937,N_1880,N_1896);
nand U1938 (N_1938,N_1899,N_1869);
or U1939 (N_1939,N_1854,N_1857);
and U1940 (N_1940,N_1891,N_1865);
and U1941 (N_1941,N_1885,N_1891);
or U1942 (N_1942,N_1877,N_1854);
nand U1943 (N_1943,N_1881,N_1877);
and U1944 (N_1944,N_1862,N_1867);
nor U1945 (N_1945,N_1859,N_1891);
xor U1946 (N_1946,N_1868,N_1853);
nand U1947 (N_1947,N_1874,N_1870);
nand U1948 (N_1948,N_1857,N_1855);
nor U1949 (N_1949,N_1898,N_1853);
or U1950 (N_1950,N_1922,N_1939);
nor U1951 (N_1951,N_1933,N_1943);
xnor U1952 (N_1952,N_1940,N_1936);
and U1953 (N_1953,N_1900,N_1944);
or U1954 (N_1954,N_1920,N_1945);
nor U1955 (N_1955,N_1923,N_1915);
and U1956 (N_1956,N_1902,N_1901);
and U1957 (N_1957,N_1937,N_1914);
nor U1958 (N_1958,N_1931,N_1906);
or U1959 (N_1959,N_1910,N_1916);
nand U1960 (N_1960,N_1941,N_1924);
nor U1961 (N_1961,N_1930,N_1904);
and U1962 (N_1962,N_1911,N_1919);
nor U1963 (N_1963,N_1947,N_1918);
nor U1964 (N_1964,N_1913,N_1927);
xor U1965 (N_1965,N_1948,N_1942);
and U1966 (N_1966,N_1912,N_1932);
and U1967 (N_1967,N_1935,N_1909);
nand U1968 (N_1968,N_1905,N_1949);
nor U1969 (N_1969,N_1925,N_1938);
nand U1970 (N_1970,N_1907,N_1917);
and U1971 (N_1971,N_1926,N_1934);
and U1972 (N_1972,N_1929,N_1946);
nand U1973 (N_1973,N_1908,N_1928);
xnor U1974 (N_1974,N_1903,N_1921);
xnor U1975 (N_1975,N_1912,N_1902);
nor U1976 (N_1976,N_1949,N_1930);
nor U1977 (N_1977,N_1927,N_1914);
and U1978 (N_1978,N_1911,N_1943);
and U1979 (N_1979,N_1943,N_1922);
or U1980 (N_1980,N_1939,N_1903);
and U1981 (N_1981,N_1949,N_1908);
or U1982 (N_1982,N_1942,N_1909);
xor U1983 (N_1983,N_1927,N_1900);
nor U1984 (N_1984,N_1922,N_1904);
and U1985 (N_1985,N_1941,N_1948);
nor U1986 (N_1986,N_1908,N_1906);
xnor U1987 (N_1987,N_1901,N_1918);
and U1988 (N_1988,N_1929,N_1949);
or U1989 (N_1989,N_1906,N_1947);
nor U1990 (N_1990,N_1910,N_1948);
xor U1991 (N_1991,N_1908,N_1901);
nor U1992 (N_1992,N_1935,N_1932);
nand U1993 (N_1993,N_1920,N_1903);
or U1994 (N_1994,N_1921,N_1927);
nor U1995 (N_1995,N_1900,N_1911);
or U1996 (N_1996,N_1932,N_1929);
nor U1997 (N_1997,N_1934,N_1947);
nor U1998 (N_1998,N_1915,N_1905);
nand U1999 (N_1999,N_1908,N_1947);
xor U2000 (N_2000,N_1993,N_1953);
and U2001 (N_2001,N_1983,N_1977);
and U2002 (N_2002,N_1986,N_1963);
nand U2003 (N_2003,N_1984,N_1992);
or U2004 (N_2004,N_1995,N_1965);
nand U2005 (N_2005,N_1985,N_1970);
or U2006 (N_2006,N_1969,N_1966);
xor U2007 (N_2007,N_1959,N_1968);
nor U2008 (N_2008,N_1955,N_1978);
nor U2009 (N_2009,N_1981,N_1975);
nand U2010 (N_2010,N_1964,N_1961);
nand U2011 (N_2011,N_1994,N_1971);
nand U2012 (N_2012,N_1950,N_1954);
and U2013 (N_2013,N_1958,N_1987);
or U2014 (N_2014,N_1956,N_1957);
nor U2015 (N_2015,N_1972,N_1973);
nor U2016 (N_2016,N_1952,N_1999);
and U2017 (N_2017,N_1967,N_1979);
nor U2018 (N_2018,N_1951,N_1991);
nand U2019 (N_2019,N_1997,N_1990);
or U2020 (N_2020,N_1960,N_1980);
nand U2021 (N_2021,N_1982,N_1996);
nand U2022 (N_2022,N_1989,N_1998);
nand U2023 (N_2023,N_1962,N_1974);
nor U2024 (N_2024,N_1976,N_1988);
and U2025 (N_2025,N_1999,N_1992);
or U2026 (N_2026,N_1960,N_1971);
nand U2027 (N_2027,N_1983,N_1989);
and U2028 (N_2028,N_1986,N_1997);
nand U2029 (N_2029,N_1962,N_1999);
and U2030 (N_2030,N_1978,N_1984);
nand U2031 (N_2031,N_1981,N_1989);
nor U2032 (N_2032,N_1988,N_1951);
or U2033 (N_2033,N_1961,N_1966);
nand U2034 (N_2034,N_1976,N_1961);
nand U2035 (N_2035,N_1980,N_1953);
nand U2036 (N_2036,N_1957,N_1967);
or U2037 (N_2037,N_1987,N_1972);
nand U2038 (N_2038,N_1973,N_1952);
nand U2039 (N_2039,N_1996,N_1952);
or U2040 (N_2040,N_1960,N_1954);
and U2041 (N_2041,N_1952,N_1953);
or U2042 (N_2042,N_1961,N_1977);
xnor U2043 (N_2043,N_1952,N_1983);
nor U2044 (N_2044,N_1964,N_1959);
and U2045 (N_2045,N_1966,N_1958);
and U2046 (N_2046,N_1983,N_1963);
nor U2047 (N_2047,N_1969,N_1987);
nor U2048 (N_2048,N_1999,N_1954);
and U2049 (N_2049,N_1979,N_1954);
nor U2050 (N_2050,N_2001,N_2017);
nand U2051 (N_2051,N_2036,N_2028);
or U2052 (N_2052,N_2010,N_2015);
and U2053 (N_2053,N_2027,N_2006);
or U2054 (N_2054,N_2023,N_2049);
xnor U2055 (N_2055,N_2022,N_2030);
nand U2056 (N_2056,N_2013,N_2011);
xnor U2057 (N_2057,N_2031,N_2008);
nor U2058 (N_2058,N_2002,N_2009);
nor U2059 (N_2059,N_2020,N_2007);
or U2060 (N_2060,N_2037,N_2043);
and U2061 (N_2061,N_2025,N_2040);
nor U2062 (N_2062,N_2038,N_2019);
xnor U2063 (N_2063,N_2046,N_2029);
and U2064 (N_2064,N_2004,N_2039);
or U2065 (N_2065,N_2034,N_2035);
nor U2066 (N_2066,N_2044,N_2033);
xor U2067 (N_2067,N_2021,N_2041);
and U2068 (N_2068,N_2018,N_2012);
and U2069 (N_2069,N_2000,N_2014);
nand U2070 (N_2070,N_2045,N_2024);
nor U2071 (N_2071,N_2042,N_2016);
nor U2072 (N_2072,N_2003,N_2026);
and U2073 (N_2073,N_2048,N_2005);
nand U2074 (N_2074,N_2032,N_2047);
xor U2075 (N_2075,N_2015,N_2039);
nor U2076 (N_2076,N_2021,N_2005);
and U2077 (N_2077,N_2049,N_2015);
nand U2078 (N_2078,N_2000,N_2041);
nor U2079 (N_2079,N_2044,N_2007);
nor U2080 (N_2080,N_2001,N_2034);
xor U2081 (N_2081,N_2049,N_2000);
nand U2082 (N_2082,N_2041,N_2004);
nor U2083 (N_2083,N_2041,N_2043);
nor U2084 (N_2084,N_2039,N_2040);
nand U2085 (N_2085,N_2049,N_2014);
or U2086 (N_2086,N_2001,N_2015);
nand U2087 (N_2087,N_2006,N_2042);
xnor U2088 (N_2088,N_2046,N_2009);
nor U2089 (N_2089,N_2018,N_2045);
nor U2090 (N_2090,N_2043,N_2004);
nand U2091 (N_2091,N_2002,N_2000);
and U2092 (N_2092,N_2045,N_2025);
or U2093 (N_2093,N_2033,N_2012);
xor U2094 (N_2094,N_2029,N_2010);
nor U2095 (N_2095,N_2000,N_2033);
nand U2096 (N_2096,N_2035,N_2019);
or U2097 (N_2097,N_2046,N_2026);
nand U2098 (N_2098,N_2047,N_2048);
nand U2099 (N_2099,N_2006,N_2020);
and U2100 (N_2100,N_2072,N_2091);
or U2101 (N_2101,N_2057,N_2052);
or U2102 (N_2102,N_2094,N_2063);
or U2103 (N_2103,N_2070,N_2065);
or U2104 (N_2104,N_2078,N_2069);
nor U2105 (N_2105,N_2058,N_2080);
and U2106 (N_2106,N_2050,N_2095);
xor U2107 (N_2107,N_2060,N_2062);
or U2108 (N_2108,N_2081,N_2073);
and U2109 (N_2109,N_2067,N_2076);
nor U2110 (N_2110,N_2097,N_2059);
and U2111 (N_2111,N_2083,N_2061);
or U2112 (N_2112,N_2088,N_2053);
nor U2113 (N_2113,N_2092,N_2084);
nand U2114 (N_2114,N_2066,N_2074);
nand U2115 (N_2115,N_2071,N_2090);
or U2116 (N_2116,N_2089,N_2096);
or U2117 (N_2117,N_2075,N_2098);
or U2118 (N_2118,N_2082,N_2054);
xnor U2119 (N_2119,N_2077,N_2064);
nand U2120 (N_2120,N_2099,N_2056);
nor U2121 (N_2121,N_2068,N_2079);
nor U2122 (N_2122,N_2085,N_2051);
nand U2123 (N_2123,N_2055,N_2086);
nand U2124 (N_2124,N_2093,N_2087);
nand U2125 (N_2125,N_2088,N_2055);
xnor U2126 (N_2126,N_2080,N_2075);
and U2127 (N_2127,N_2069,N_2077);
or U2128 (N_2128,N_2094,N_2080);
nor U2129 (N_2129,N_2058,N_2085);
xor U2130 (N_2130,N_2072,N_2078);
or U2131 (N_2131,N_2082,N_2080);
nand U2132 (N_2132,N_2086,N_2073);
and U2133 (N_2133,N_2093,N_2064);
nand U2134 (N_2134,N_2059,N_2096);
or U2135 (N_2135,N_2061,N_2098);
and U2136 (N_2136,N_2090,N_2098);
xor U2137 (N_2137,N_2073,N_2067);
nor U2138 (N_2138,N_2073,N_2091);
and U2139 (N_2139,N_2076,N_2088);
and U2140 (N_2140,N_2059,N_2083);
nor U2141 (N_2141,N_2082,N_2084);
nor U2142 (N_2142,N_2090,N_2096);
nor U2143 (N_2143,N_2067,N_2053);
nor U2144 (N_2144,N_2050,N_2091);
nor U2145 (N_2145,N_2080,N_2052);
nor U2146 (N_2146,N_2074,N_2085);
and U2147 (N_2147,N_2065,N_2056);
or U2148 (N_2148,N_2078,N_2093);
and U2149 (N_2149,N_2076,N_2064);
or U2150 (N_2150,N_2124,N_2125);
and U2151 (N_2151,N_2145,N_2119);
nor U2152 (N_2152,N_2123,N_2131);
nor U2153 (N_2153,N_2129,N_2105);
nor U2154 (N_2154,N_2141,N_2132);
nand U2155 (N_2155,N_2111,N_2133);
or U2156 (N_2156,N_2147,N_2121);
and U2157 (N_2157,N_2107,N_2112);
and U2158 (N_2158,N_2118,N_2114);
nor U2159 (N_2159,N_2122,N_2146);
and U2160 (N_2160,N_2137,N_2148);
nand U2161 (N_2161,N_2115,N_2143);
or U2162 (N_2162,N_2110,N_2106);
nor U2163 (N_2163,N_2100,N_2130);
and U2164 (N_2164,N_2103,N_2117);
nor U2165 (N_2165,N_2116,N_2108);
and U2166 (N_2166,N_2134,N_2135);
or U2167 (N_2167,N_2138,N_2127);
nand U2168 (N_2168,N_2102,N_2142);
nand U2169 (N_2169,N_2104,N_2144);
nand U2170 (N_2170,N_2140,N_2101);
and U2171 (N_2171,N_2120,N_2149);
nand U2172 (N_2172,N_2113,N_2126);
nor U2173 (N_2173,N_2109,N_2136);
or U2174 (N_2174,N_2128,N_2139);
nor U2175 (N_2175,N_2110,N_2112);
or U2176 (N_2176,N_2125,N_2115);
nor U2177 (N_2177,N_2148,N_2145);
nor U2178 (N_2178,N_2136,N_2130);
xor U2179 (N_2179,N_2108,N_2130);
nor U2180 (N_2180,N_2123,N_2133);
and U2181 (N_2181,N_2140,N_2106);
and U2182 (N_2182,N_2120,N_2128);
or U2183 (N_2183,N_2148,N_2113);
nand U2184 (N_2184,N_2128,N_2142);
or U2185 (N_2185,N_2138,N_2140);
xor U2186 (N_2186,N_2136,N_2106);
and U2187 (N_2187,N_2149,N_2147);
and U2188 (N_2188,N_2141,N_2115);
nor U2189 (N_2189,N_2109,N_2130);
nor U2190 (N_2190,N_2140,N_2105);
nand U2191 (N_2191,N_2115,N_2129);
nor U2192 (N_2192,N_2134,N_2108);
nor U2193 (N_2193,N_2105,N_2117);
nand U2194 (N_2194,N_2126,N_2125);
or U2195 (N_2195,N_2117,N_2137);
xor U2196 (N_2196,N_2108,N_2112);
nor U2197 (N_2197,N_2115,N_2106);
nand U2198 (N_2198,N_2112,N_2138);
xnor U2199 (N_2199,N_2104,N_2128);
and U2200 (N_2200,N_2167,N_2163);
xor U2201 (N_2201,N_2159,N_2157);
nor U2202 (N_2202,N_2194,N_2160);
or U2203 (N_2203,N_2177,N_2193);
nor U2204 (N_2204,N_2153,N_2184);
nand U2205 (N_2205,N_2189,N_2161);
nor U2206 (N_2206,N_2171,N_2178);
xor U2207 (N_2207,N_2185,N_2176);
or U2208 (N_2208,N_2162,N_2172);
and U2209 (N_2209,N_2175,N_2197);
or U2210 (N_2210,N_2179,N_2181);
and U2211 (N_2211,N_2199,N_2165);
xnor U2212 (N_2212,N_2166,N_2150);
and U2213 (N_2213,N_2188,N_2196);
nor U2214 (N_2214,N_2174,N_2187);
nand U2215 (N_2215,N_2152,N_2154);
nor U2216 (N_2216,N_2195,N_2151);
nand U2217 (N_2217,N_2183,N_2164);
and U2218 (N_2218,N_2169,N_2170);
and U2219 (N_2219,N_2198,N_2182);
and U2220 (N_2220,N_2190,N_2156);
or U2221 (N_2221,N_2168,N_2155);
nand U2222 (N_2222,N_2191,N_2192);
and U2223 (N_2223,N_2158,N_2186);
and U2224 (N_2224,N_2173,N_2180);
and U2225 (N_2225,N_2170,N_2198);
nand U2226 (N_2226,N_2186,N_2155);
and U2227 (N_2227,N_2188,N_2160);
xor U2228 (N_2228,N_2191,N_2176);
or U2229 (N_2229,N_2150,N_2174);
xor U2230 (N_2230,N_2175,N_2177);
xor U2231 (N_2231,N_2151,N_2193);
nand U2232 (N_2232,N_2169,N_2154);
xnor U2233 (N_2233,N_2185,N_2192);
nor U2234 (N_2234,N_2198,N_2195);
nand U2235 (N_2235,N_2166,N_2187);
nor U2236 (N_2236,N_2157,N_2173);
or U2237 (N_2237,N_2152,N_2185);
and U2238 (N_2238,N_2183,N_2151);
nand U2239 (N_2239,N_2184,N_2179);
or U2240 (N_2240,N_2198,N_2151);
xor U2241 (N_2241,N_2186,N_2181);
nand U2242 (N_2242,N_2155,N_2194);
nand U2243 (N_2243,N_2178,N_2189);
or U2244 (N_2244,N_2152,N_2163);
nor U2245 (N_2245,N_2165,N_2168);
or U2246 (N_2246,N_2183,N_2181);
nor U2247 (N_2247,N_2173,N_2198);
nor U2248 (N_2248,N_2184,N_2190);
nand U2249 (N_2249,N_2181,N_2163);
and U2250 (N_2250,N_2243,N_2233);
nor U2251 (N_2251,N_2220,N_2227);
and U2252 (N_2252,N_2204,N_2209);
and U2253 (N_2253,N_2230,N_2235);
nor U2254 (N_2254,N_2248,N_2213);
nand U2255 (N_2255,N_2226,N_2228);
nand U2256 (N_2256,N_2216,N_2242);
xor U2257 (N_2257,N_2203,N_2232);
or U2258 (N_2258,N_2231,N_2218);
or U2259 (N_2259,N_2229,N_2249);
or U2260 (N_2260,N_2222,N_2237);
nand U2261 (N_2261,N_2240,N_2206);
nand U2262 (N_2262,N_2239,N_2221);
nor U2263 (N_2263,N_2205,N_2201);
nor U2264 (N_2264,N_2241,N_2236);
nor U2265 (N_2265,N_2219,N_2207);
and U2266 (N_2266,N_2224,N_2215);
nor U2267 (N_2267,N_2225,N_2214);
or U2268 (N_2268,N_2211,N_2238);
nor U2269 (N_2269,N_2244,N_2247);
nor U2270 (N_2270,N_2223,N_2208);
and U2271 (N_2271,N_2217,N_2200);
nand U2272 (N_2272,N_2210,N_2202);
or U2273 (N_2273,N_2246,N_2212);
nor U2274 (N_2274,N_2245,N_2234);
and U2275 (N_2275,N_2245,N_2241);
or U2276 (N_2276,N_2211,N_2248);
nand U2277 (N_2277,N_2213,N_2206);
nand U2278 (N_2278,N_2213,N_2211);
nand U2279 (N_2279,N_2249,N_2237);
xor U2280 (N_2280,N_2212,N_2237);
and U2281 (N_2281,N_2232,N_2238);
and U2282 (N_2282,N_2237,N_2233);
or U2283 (N_2283,N_2240,N_2205);
nand U2284 (N_2284,N_2242,N_2240);
nand U2285 (N_2285,N_2221,N_2242);
or U2286 (N_2286,N_2227,N_2245);
nor U2287 (N_2287,N_2230,N_2220);
xnor U2288 (N_2288,N_2216,N_2221);
nor U2289 (N_2289,N_2219,N_2243);
or U2290 (N_2290,N_2206,N_2237);
or U2291 (N_2291,N_2246,N_2205);
or U2292 (N_2292,N_2224,N_2210);
and U2293 (N_2293,N_2230,N_2216);
nor U2294 (N_2294,N_2222,N_2225);
xnor U2295 (N_2295,N_2245,N_2204);
nor U2296 (N_2296,N_2216,N_2210);
and U2297 (N_2297,N_2238,N_2245);
and U2298 (N_2298,N_2246,N_2235);
nor U2299 (N_2299,N_2200,N_2212);
nand U2300 (N_2300,N_2269,N_2266);
xor U2301 (N_2301,N_2274,N_2294);
and U2302 (N_2302,N_2261,N_2251);
or U2303 (N_2303,N_2283,N_2270);
and U2304 (N_2304,N_2268,N_2272);
nor U2305 (N_2305,N_2260,N_2299);
and U2306 (N_2306,N_2263,N_2291);
and U2307 (N_2307,N_2276,N_2284);
or U2308 (N_2308,N_2255,N_2277);
nor U2309 (N_2309,N_2292,N_2256);
and U2310 (N_2310,N_2287,N_2282);
nor U2311 (N_2311,N_2295,N_2265);
nor U2312 (N_2312,N_2257,N_2288);
or U2313 (N_2313,N_2275,N_2289);
nand U2314 (N_2314,N_2267,N_2296);
nand U2315 (N_2315,N_2290,N_2252);
nor U2316 (N_2316,N_2278,N_2298);
or U2317 (N_2317,N_2253,N_2271);
xnor U2318 (N_2318,N_2285,N_2293);
nor U2319 (N_2319,N_2264,N_2259);
nor U2320 (N_2320,N_2297,N_2254);
nor U2321 (N_2321,N_2286,N_2262);
or U2322 (N_2322,N_2281,N_2250);
xor U2323 (N_2323,N_2279,N_2273);
nor U2324 (N_2324,N_2258,N_2280);
and U2325 (N_2325,N_2296,N_2299);
or U2326 (N_2326,N_2299,N_2263);
nor U2327 (N_2327,N_2297,N_2287);
nand U2328 (N_2328,N_2279,N_2251);
nor U2329 (N_2329,N_2255,N_2269);
and U2330 (N_2330,N_2273,N_2263);
nor U2331 (N_2331,N_2262,N_2275);
xnor U2332 (N_2332,N_2274,N_2293);
nor U2333 (N_2333,N_2271,N_2287);
or U2334 (N_2334,N_2287,N_2286);
xor U2335 (N_2335,N_2299,N_2271);
and U2336 (N_2336,N_2294,N_2279);
or U2337 (N_2337,N_2254,N_2279);
and U2338 (N_2338,N_2277,N_2275);
or U2339 (N_2339,N_2294,N_2281);
or U2340 (N_2340,N_2255,N_2257);
nor U2341 (N_2341,N_2277,N_2283);
nand U2342 (N_2342,N_2262,N_2267);
or U2343 (N_2343,N_2289,N_2287);
or U2344 (N_2344,N_2286,N_2260);
nor U2345 (N_2345,N_2277,N_2290);
nor U2346 (N_2346,N_2261,N_2286);
nand U2347 (N_2347,N_2250,N_2267);
or U2348 (N_2348,N_2256,N_2250);
nand U2349 (N_2349,N_2280,N_2270);
xnor U2350 (N_2350,N_2325,N_2343);
nor U2351 (N_2351,N_2332,N_2314);
nor U2352 (N_2352,N_2311,N_2331);
xnor U2353 (N_2353,N_2321,N_2315);
and U2354 (N_2354,N_2320,N_2341);
nand U2355 (N_2355,N_2328,N_2330);
xor U2356 (N_2356,N_2313,N_2333);
and U2357 (N_2357,N_2317,N_2309);
and U2358 (N_2358,N_2308,N_2340);
nand U2359 (N_2359,N_2324,N_2334);
nand U2360 (N_2360,N_2329,N_2339);
nor U2361 (N_2361,N_2319,N_2344);
nand U2362 (N_2362,N_2303,N_2304);
or U2363 (N_2363,N_2302,N_2306);
or U2364 (N_2364,N_2316,N_2347);
nand U2365 (N_2365,N_2318,N_2322);
and U2366 (N_2366,N_2346,N_2305);
nor U2367 (N_2367,N_2338,N_2300);
xor U2368 (N_2368,N_2349,N_2342);
or U2369 (N_2369,N_2345,N_2337);
or U2370 (N_2370,N_2336,N_2310);
and U2371 (N_2371,N_2348,N_2335);
nand U2372 (N_2372,N_2307,N_2312);
or U2373 (N_2373,N_2301,N_2327);
or U2374 (N_2374,N_2326,N_2323);
and U2375 (N_2375,N_2306,N_2327);
nor U2376 (N_2376,N_2305,N_2306);
nor U2377 (N_2377,N_2304,N_2344);
or U2378 (N_2378,N_2322,N_2320);
nand U2379 (N_2379,N_2337,N_2332);
or U2380 (N_2380,N_2348,N_2310);
nand U2381 (N_2381,N_2323,N_2336);
xnor U2382 (N_2382,N_2349,N_2317);
nand U2383 (N_2383,N_2334,N_2319);
xnor U2384 (N_2384,N_2302,N_2347);
or U2385 (N_2385,N_2342,N_2309);
and U2386 (N_2386,N_2343,N_2318);
nor U2387 (N_2387,N_2304,N_2333);
or U2388 (N_2388,N_2304,N_2332);
and U2389 (N_2389,N_2301,N_2343);
nand U2390 (N_2390,N_2349,N_2340);
nor U2391 (N_2391,N_2311,N_2338);
nand U2392 (N_2392,N_2312,N_2333);
nand U2393 (N_2393,N_2311,N_2337);
or U2394 (N_2394,N_2344,N_2335);
or U2395 (N_2395,N_2318,N_2301);
nand U2396 (N_2396,N_2331,N_2334);
nor U2397 (N_2397,N_2323,N_2348);
xnor U2398 (N_2398,N_2316,N_2335);
or U2399 (N_2399,N_2314,N_2301);
or U2400 (N_2400,N_2356,N_2392);
nand U2401 (N_2401,N_2393,N_2362);
nand U2402 (N_2402,N_2387,N_2355);
or U2403 (N_2403,N_2351,N_2354);
and U2404 (N_2404,N_2363,N_2373);
nor U2405 (N_2405,N_2369,N_2388);
and U2406 (N_2406,N_2391,N_2397);
and U2407 (N_2407,N_2377,N_2361);
or U2408 (N_2408,N_2395,N_2360);
nor U2409 (N_2409,N_2379,N_2353);
nand U2410 (N_2410,N_2357,N_2350);
and U2411 (N_2411,N_2365,N_2383);
and U2412 (N_2412,N_2396,N_2384);
and U2413 (N_2413,N_2385,N_2380);
nor U2414 (N_2414,N_2371,N_2368);
nand U2415 (N_2415,N_2389,N_2386);
or U2416 (N_2416,N_2375,N_2390);
nand U2417 (N_2417,N_2398,N_2378);
or U2418 (N_2418,N_2376,N_2381);
and U2419 (N_2419,N_2399,N_2382);
and U2420 (N_2420,N_2359,N_2358);
and U2421 (N_2421,N_2366,N_2364);
xor U2422 (N_2422,N_2352,N_2370);
xnor U2423 (N_2423,N_2372,N_2394);
and U2424 (N_2424,N_2374,N_2367);
nand U2425 (N_2425,N_2366,N_2356);
nor U2426 (N_2426,N_2386,N_2376);
or U2427 (N_2427,N_2358,N_2374);
nand U2428 (N_2428,N_2373,N_2396);
nor U2429 (N_2429,N_2376,N_2385);
nor U2430 (N_2430,N_2360,N_2355);
and U2431 (N_2431,N_2374,N_2351);
and U2432 (N_2432,N_2390,N_2353);
and U2433 (N_2433,N_2381,N_2355);
and U2434 (N_2434,N_2383,N_2387);
nand U2435 (N_2435,N_2358,N_2352);
nand U2436 (N_2436,N_2381,N_2378);
or U2437 (N_2437,N_2390,N_2393);
or U2438 (N_2438,N_2386,N_2360);
xnor U2439 (N_2439,N_2352,N_2356);
nor U2440 (N_2440,N_2355,N_2383);
and U2441 (N_2441,N_2399,N_2396);
or U2442 (N_2442,N_2365,N_2398);
nor U2443 (N_2443,N_2379,N_2371);
nor U2444 (N_2444,N_2397,N_2350);
nand U2445 (N_2445,N_2375,N_2389);
nand U2446 (N_2446,N_2386,N_2385);
and U2447 (N_2447,N_2380,N_2378);
or U2448 (N_2448,N_2375,N_2395);
or U2449 (N_2449,N_2379,N_2365);
and U2450 (N_2450,N_2421,N_2426);
nor U2451 (N_2451,N_2431,N_2406);
or U2452 (N_2452,N_2403,N_2402);
nand U2453 (N_2453,N_2415,N_2427);
and U2454 (N_2454,N_2408,N_2407);
nand U2455 (N_2455,N_2449,N_2423);
nor U2456 (N_2456,N_2438,N_2443);
nor U2457 (N_2457,N_2412,N_2400);
nand U2458 (N_2458,N_2404,N_2417);
nand U2459 (N_2459,N_2432,N_2428);
and U2460 (N_2460,N_2410,N_2413);
nand U2461 (N_2461,N_2422,N_2434);
nor U2462 (N_2462,N_2424,N_2436);
nand U2463 (N_2463,N_2429,N_2430);
or U2464 (N_2464,N_2419,N_2405);
nand U2465 (N_2465,N_2416,N_2409);
and U2466 (N_2466,N_2420,N_2418);
and U2467 (N_2467,N_2414,N_2440);
and U2468 (N_2468,N_2425,N_2448);
and U2469 (N_2469,N_2445,N_2444);
and U2470 (N_2470,N_2433,N_2447);
nand U2471 (N_2471,N_2437,N_2441);
nand U2472 (N_2472,N_2401,N_2411);
nand U2473 (N_2473,N_2446,N_2439);
or U2474 (N_2474,N_2435,N_2442);
nand U2475 (N_2475,N_2423,N_2435);
or U2476 (N_2476,N_2438,N_2441);
and U2477 (N_2477,N_2433,N_2430);
and U2478 (N_2478,N_2438,N_2406);
xnor U2479 (N_2479,N_2422,N_2407);
nor U2480 (N_2480,N_2436,N_2402);
nor U2481 (N_2481,N_2416,N_2412);
and U2482 (N_2482,N_2436,N_2429);
and U2483 (N_2483,N_2438,N_2442);
and U2484 (N_2484,N_2445,N_2439);
nor U2485 (N_2485,N_2446,N_2406);
or U2486 (N_2486,N_2443,N_2433);
xor U2487 (N_2487,N_2403,N_2431);
or U2488 (N_2488,N_2435,N_2429);
nor U2489 (N_2489,N_2416,N_2418);
and U2490 (N_2490,N_2415,N_2428);
nor U2491 (N_2491,N_2442,N_2418);
and U2492 (N_2492,N_2420,N_2438);
nand U2493 (N_2493,N_2405,N_2430);
and U2494 (N_2494,N_2400,N_2411);
or U2495 (N_2495,N_2448,N_2428);
nor U2496 (N_2496,N_2407,N_2405);
nor U2497 (N_2497,N_2409,N_2425);
nand U2498 (N_2498,N_2448,N_2435);
nand U2499 (N_2499,N_2434,N_2426);
or U2500 (N_2500,N_2459,N_2454);
and U2501 (N_2501,N_2499,N_2465);
nor U2502 (N_2502,N_2480,N_2489);
nand U2503 (N_2503,N_2486,N_2485);
nand U2504 (N_2504,N_2456,N_2479);
nand U2505 (N_2505,N_2455,N_2464);
or U2506 (N_2506,N_2470,N_2460);
nor U2507 (N_2507,N_2496,N_2493);
nand U2508 (N_2508,N_2488,N_2450);
and U2509 (N_2509,N_2487,N_2477);
and U2510 (N_2510,N_2492,N_2457);
nor U2511 (N_2511,N_2466,N_2476);
or U2512 (N_2512,N_2472,N_2494);
nand U2513 (N_2513,N_2481,N_2451);
nand U2514 (N_2514,N_2490,N_2483);
nor U2515 (N_2515,N_2461,N_2453);
or U2516 (N_2516,N_2484,N_2463);
or U2517 (N_2517,N_2468,N_2478);
xnor U2518 (N_2518,N_2462,N_2474);
or U2519 (N_2519,N_2471,N_2491);
or U2520 (N_2520,N_2475,N_2497);
or U2521 (N_2521,N_2482,N_2467);
or U2522 (N_2522,N_2458,N_2469);
nand U2523 (N_2523,N_2452,N_2473);
and U2524 (N_2524,N_2495,N_2498);
and U2525 (N_2525,N_2491,N_2494);
and U2526 (N_2526,N_2455,N_2493);
nor U2527 (N_2527,N_2469,N_2450);
nand U2528 (N_2528,N_2466,N_2467);
nor U2529 (N_2529,N_2477,N_2455);
or U2530 (N_2530,N_2486,N_2487);
or U2531 (N_2531,N_2494,N_2486);
and U2532 (N_2532,N_2459,N_2494);
nand U2533 (N_2533,N_2492,N_2453);
or U2534 (N_2534,N_2452,N_2482);
or U2535 (N_2535,N_2476,N_2486);
xnor U2536 (N_2536,N_2493,N_2483);
and U2537 (N_2537,N_2457,N_2476);
or U2538 (N_2538,N_2451,N_2493);
or U2539 (N_2539,N_2475,N_2450);
nand U2540 (N_2540,N_2455,N_2463);
or U2541 (N_2541,N_2495,N_2482);
or U2542 (N_2542,N_2482,N_2471);
or U2543 (N_2543,N_2494,N_2460);
and U2544 (N_2544,N_2486,N_2462);
and U2545 (N_2545,N_2478,N_2490);
nand U2546 (N_2546,N_2494,N_2475);
nand U2547 (N_2547,N_2497,N_2483);
nand U2548 (N_2548,N_2475,N_2461);
and U2549 (N_2549,N_2492,N_2496);
and U2550 (N_2550,N_2544,N_2541);
nand U2551 (N_2551,N_2548,N_2505);
nand U2552 (N_2552,N_2539,N_2515);
and U2553 (N_2553,N_2522,N_2516);
and U2554 (N_2554,N_2526,N_2514);
and U2555 (N_2555,N_2540,N_2537);
nor U2556 (N_2556,N_2525,N_2546);
nand U2557 (N_2557,N_2535,N_2545);
xnor U2558 (N_2558,N_2506,N_2512);
or U2559 (N_2559,N_2501,N_2538);
nor U2560 (N_2560,N_2542,N_2533);
and U2561 (N_2561,N_2502,N_2517);
nand U2562 (N_2562,N_2510,N_2529);
and U2563 (N_2563,N_2534,N_2531);
nand U2564 (N_2564,N_2523,N_2527);
and U2565 (N_2565,N_2524,N_2513);
nand U2566 (N_2566,N_2549,N_2521);
nor U2567 (N_2567,N_2518,N_2504);
nor U2568 (N_2568,N_2511,N_2503);
and U2569 (N_2569,N_2508,N_2520);
nand U2570 (N_2570,N_2543,N_2536);
and U2571 (N_2571,N_2530,N_2532);
or U2572 (N_2572,N_2519,N_2507);
nand U2573 (N_2573,N_2509,N_2500);
and U2574 (N_2574,N_2528,N_2547);
xor U2575 (N_2575,N_2506,N_2534);
or U2576 (N_2576,N_2523,N_2536);
or U2577 (N_2577,N_2528,N_2515);
nand U2578 (N_2578,N_2517,N_2504);
xnor U2579 (N_2579,N_2540,N_2525);
or U2580 (N_2580,N_2530,N_2528);
or U2581 (N_2581,N_2542,N_2524);
nand U2582 (N_2582,N_2530,N_2521);
nor U2583 (N_2583,N_2527,N_2531);
and U2584 (N_2584,N_2534,N_2501);
and U2585 (N_2585,N_2540,N_2506);
xor U2586 (N_2586,N_2535,N_2501);
and U2587 (N_2587,N_2521,N_2525);
or U2588 (N_2588,N_2511,N_2520);
xnor U2589 (N_2589,N_2510,N_2516);
nor U2590 (N_2590,N_2509,N_2522);
nand U2591 (N_2591,N_2537,N_2539);
nor U2592 (N_2592,N_2514,N_2506);
nand U2593 (N_2593,N_2528,N_2526);
nand U2594 (N_2594,N_2533,N_2501);
nor U2595 (N_2595,N_2505,N_2515);
nand U2596 (N_2596,N_2543,N_2523);
or U2597 (N_2597,N_2526,N_2527);
xnor U2598 (N_2598,N_2524,N_2536);
nand U2599 (N_2599,N_2549,N_2502);
or U2600 (N_2600,N_2555,N_2596);
or U2601 (N_2601,N_2560,N_2598);
nand U2602 (N_2602,N_2550,N_2585);
or U2603 (N_2603,N_2576,N_2586);
or U2604 (N_2604,N_2574,N_2591);
nor U2605 (N_2605,N_2557,N_2595);
nor U2606 (N_2606,N_2593,N_2592);
nand U2607 (N_2607,N_2567,N_2583);
nand U2608 (N_2608,N_2566,N_2572);
nor U2609 (N_2609,N_2589,N_2556);
and U2610 (N_2610,N_2579,N_2554);
nand U2611 (N_2611,N_2564,N_2573);
nand U2612 (N_2612,N_2581,N_2565);
or U2613 (N_2613,N_2561,N_2551);
and U2614 (N_2614,N_2590,N_2559);
nand U2615 (N_2615,N_2552,N_2575);
nor U2616 (N_2616,N_2578,N_2584);
nand U2617 (N_2617,N_2562,N_2568);
and U2618 (N_2618,N_2571,N_2580);
and U2619 (N_2619,N_2553,N_2594);
nor U2620 (N_2620,N_2558,N_2577);
and U2621 (N_2621,N_2588,N_2563);
nand U2622 (N_2622,N_2569,N_2582);
nor U2623 (N_2623,N_2570,N_2597);
and U2624 (N_2624,N_2599,N_2587);
xnor U2625 (N_2625,N_2554,N_2551);
or U2626 (N_2626,N_2572,N_2579);
nand U2627 (N_2627,N_2590,N_2573);
or U2628 (N_2628,N_2560,N_2592);
nor U2629 (N_2629,N_2553,N_2597);
xor U2630 (N_2630,N_2582,N_2564);
nand U2631 (N_2631,N_2594,N_2596);
nand U2632 (N_2632,N_2590,N_2564);
and U2633 (N_2633,N_2575,N_2558);
nand U2634 (N_2634,N_2562,N_2579);
or U2635 (N_2635,N_2569,N_2593);
or U2636 (N_2636,N_2585,N_2570);
or U2637 (N_2637,N_2558,N_2568);
nor U2638 (N_2638,N_2567,N_2597);
nor U2639 (N_2639,N_2570,N_2586);
nor U2640 (N_2640,N_2591,N_2558);
or U2641 (N_2641,N_2599,N_2584);
nor U2642 (N_2642,N_2578,N_2589);
and U2643 (N_2643,N_2588,N_2570);
nand U2644 (N_2644,N_2550,N_2588);
xnor U2645 (N_2645,N_2555,N_2575);
nand U2646 (N_2646,N_2557,N_2585);
or U2647 (N_2647,N_2576,N_2582);
or U2648 (N_2648,N_2550,N_2587);
nor U2649 (N_2649,N_2584,N_2568);
nor U2650 (N_2650,N_2612,N_2604);
xor U2651 (N_2651,N_2623,N_2639);
nor U2652 (N_2652,N_2627,N_2608);
and U2653 (N_2653,N_2637,N_2640);
nor U2654 (N_2654,N_2633,N_2602);
and U2655 (N_2655,N_2624,N_2648);
or U2656 (N_2656,N_2638,N_2646);
xor U2657 (N_2657,N_2603,N_2605);
nand U2658 (N_2658,N_2635,N_2642);
or U2659 (N_2659,N_2647,N_2601);
nor U2660 (N_2660,N_2618,N_2621);
and U2661 (N_2661,N_2606,N_2610);
and U2662 (N_2662,N_2600,N_2630);
nor U2663 (N_2663,N_2649,N_2634);
and U2664 (N_2664,N_2644,N_2613);
or U2665 (N_2665,N_2615,N_2619);
nand U2666 (N_2666,N_2631,N_2643);
and U2667 (N_2667,N_2645,N_2611);
nand U2668 (N_2668,N_2626,N_2614);
nor U2669 (N_2669,N_2628,N_2625);
or U2670 (N_2670,N_2620,N_2622);
nand U2671 (N_2671,N_2641,N_2632);
xnor U2672 (N_2672,N_2609,N_2607);
nand U2673 (N_2673,N_2636,N_2616);
nand U2674 (N_2674,N_2617,N_2629);
nor U2675 (N_2675,N_2648,N_2606);
nand U2676 (N_2676,N_2641,N_2622);
nor U2677 (N_2677,N_2608,N_2617);
xor U2678 (N_2678,N_2623,N_2633);
nand U2679 (N_2679,N_2617,N_2645);
nor U2680 (N_2680,N_2601,N_2611);
and U2681 (N_2681,N_2631,N_2645);
or U2682 (N_2682,N_2626,N_2627);
xor U2683 (N_2683,N_2637,N_2622);
xor U2684 (N_2684,N_2647,N_2606);
xor U2685 (N_2685,N_2628,N_2632);
nor U2686 (N_2686,N_2623,N_2646);
nand U2687 (N_2687,N_2628,N_2630);
or U2688 (N_2688,N_2608,N_2609);
and U2689 (N_2689,N_2616,N_2602);
nor U2690 (N_2690,N_2649,N_2617);
and U2691 (N_2691,N_2632,N_2606);
and U2692 (N_2692,N_2635,N_2634);
and U2693 (N_2693,N_2634,N_2643);
nand U2694 (N_2694,N_2640,N_2626);
nand U2695 (N_2695,N_2618,N_2630);
and U2696 (N_2696,N_2617,N_2604);
nor U2697 (N_2697,N_2609,N_2604);
or U2698 (N_2698,N_2645,N_2649);
nor U2699 (N_2699,N_2645,N_2607);
nor U2700 (N_2700,N_2678,N_2683);
nand U2701 (N_2701,N_2688,N_2689);
and U2702 (N_2702,N_2679,N_2667);
xnor U2703 (N_2703,N_2677,N_2697);
nand U2704 (N_2704,N_2674,N_2693);
and U2705 (N_2705,N_2650,N_2666);
and U2706 (N_2706,N_2669,N_2661);
or U2707 (N_2707,N_2668,N_2696);
and U2708 (N_2708,N_2673,N_2699);
xor U2709 (N_2709,N_2692,N_2663);
xor U2710 (N_2710,N_2690,N_2682);
xnor U2711 (N_2711,N_2654,N_2657);
nand U2712 (N_2712,N_2694,N_2671);
and U2713 (N_2713,N_2662,N_2675);
nand U2714 (N_2714,N_2676,N_2686);
nand U2715 (N_2715,N_2698,N_2653);
and U2716 (N_2716,N_2658,N_2685);
and U2717 (N_2717,N_2659,N_2687);
nand U2718 (N_2718,N_2651,N_2656);
nand U2719 (N_2719,N_2680,N_2655);
or U2720 (N_2720,N_2664,N_2670);
xor U2721 (N_2721,N_2691,N_2660);
nand U2722 (N_2722,N_2665,N_2695);
xnor U2723 (N_2723,N_2681,N_2672);
and U2724 (N_2724,N_2652,N_2684);
nor U2725 (N_2725,N_2651,N_2660);
nand U2726 (N_2726,N_2653,N_2699);
and U2727 (N_2727,N_2690,N_2694);
or U2728 (N_2728,N_2654,N_2666);
or U2729 (N_2729,N_2656,N_2677);
nor U2730 (N_2730,N_2688,N_2661);
nor U2731 (N_2731,N_2680,N_2679);
nor U2732 (N_2732,N_2695,N_2653);
and U2733 (N_2733,N_2651,N_2671);
nor U2734 (N_2734,N_2679,N_2670);
nand U2735 (N_2735,N_2652,N_2678);
xnor U2736 (N_2736,N_2655,N_2682);
and U2737 (N_2737,N_2661,N_2651);
or U2738 (N_2738,N_2678,N_2696);
nor U2739 (N_2739,N_2696,N_2673);
nand U2740 (N_2740,N_2661,N_2674);
and U2741 (N_2741,N_2663,N_2653);
or U2742 (N_2742,N_2661,N_2695);
xor U2743 (N_2743,N_2685,N_2677);
and U2744 (N_2744,N_2668,N_2699);
nor U2745 (N_2745,N_2668,N_2652);
and U2746 (N_2746,N_2698,N_2663);
or U2747 (N_2747,N_2682,N_2683);
nor U2748 (N_2748,N_2655,N_2663);
and U2749 (N_2749,N_2695,N_2694);
and U2750 (N_2750,N_2749,N_2704);
xor U2751 (N_2751,N_2706,N_2746);
and U2752 (N_2752,N_2702,N_2747);
nand U2753 (N_2753,N_2726,N_2740);
or U2754 (N_2754,N_2703,N_2730);
xnor U2755 (N_2755,N_2722,N_2738);
and U2756 (N_2756,N_2719,N_2723);
nand U2757 (N_2757,N_2737,N_2733);
nor U2758 (N_2758,N_2743,N_2729);
or U2759 (N_2759,N_2715,N_2731);
or U2760 (N_2760,N_2744,N_2700);
or U2761 (N_2761,N_2712,N_2701);
or U2762 (N_2762,N_2709,N_2708);
and U2763 (N_2763,N_2720,N_2728);
or U2764 (N_2764,N_2741,N_2705);
and U2765 (N_2765,N_2724,N_2736);
or U2766 (N_2766,N_2710,N_2739);
and U2767 (N_2767,N_2727,N_2718);
nand U2768 (N_2768,N_2734,N_2745);
and U2769 (N_2769,N_2714,N_2735);
nor U2770 (N_2770,N_2717,N_2748);
xnor U2771 (N_2771,N_2732,N_2716);
nand U2772 (N_2772,N_2742,N_2713);
or U2773 (N_2773,N_2725,N_2721);
nand U2774 (N_2774,N_2711,N_2707);
nand U2775 (N_2775,N_2747,N_2739);
xor U2776 (N_2776,N_2712,N_2705);
and U2777 (N_2777,N_2736,N_2719);
nand U2778 (N_2778,N_2706,N_2703);
nand U2779 (N_2779,N_2721,N_2712);
nor U2780 (N_2780,N_2734,N_2703);
xnor U2781 (N_2781,N_2716,N_2726);
and U2782 (N_2782,N_2733,N_2735);
or U2783 (N_2783,N_2741,N_2715);
nand U2784 (N_2784,N_2732,N_2729);
or U2785 (N_2785,N_2745,N_2700);
and U2786 (N_2786,N_2702,N_2703);
and U2787 (N_2787,N_2720,N_2733);
nor U2788 (N_2788,N_2739,N_2709);
or U2789 (N_2789,N_2723,N_2711);
or U2790 (N_2790,N_2701,N_2744);
nor U2791 (N_2791,N_2722,N_2743);
nor U2792 (N_2792,N_2717,N_2732);
nor U2793 (N_2793,N_2732,N_2708);
nand U2794 (N_2794,N_2736,N_2703);
nor U2795 (N_2795,N_2748,N_2736);
or U2796 (N_2796,N_2741,N_2701);
nor U2797 (N_2797,N_2724,N_2721);
or U2798 (N_2798,N_2728,N_2749);
or U2799 (N_2799,N_2747,N_2700);
nand U2800 (N_2800,N_2787,N_2768);
nor U2801 (N_2801,N_2774,N_2756);
xnor U2802 (N_2802,N_2795,N_2757);
nand U2803 (N_2803,N_2789,N_2773);
xor U2804 (N_2804,N_2752,N_2797);
nand U2805 (N_2805,N_2750,N_2780);
nor U2806 (N_2806,N_2767,N_2771);
nor U2807 (N_2807,N_2755,N_2786);
nand U2808 (N_2808,N_2776,N_2791);
nand U2809 (N_2809,N_2763,N_2758);
xnor U2810 (N_2810,N_2777,N_2759);
and U2811 (N_2811,N_2762,N_2785);
nor U2812 (N_2812,N_2790,N_2760);
xor U2813 (N_2813,N_2753,N_2772);
xnor U2814 (N_2814,N_2796,N_2799);
and U2815 (N_2815,N_2782,N_2793);
and U2816 (N_2816,N_2751,N_2761);
nand U2817 (N_2817,N_2783,N_2794);
and U2818 (N_2818,N_2779,N_2764);
and U2819 (N_2819,N_2788,N_2792);
or U2820 (N_2820,N_2754,N_2766);
or U2821 (N_2821,N_2775,N_2784);
nand U2822 (N_2822,N_2765,N_2778);
nand U2823 (N_2823,N_2770,N_2798);
nor U2824 (N_2824,N_2769,N_2781);
xor U2825 (N_2825,N_2796,N_2779);
and U2826 (N_2826,N_2795,N_2799);
or U2827 (N_2827,N_2764,N_2795);
nand U2828 (N_2828,N_2760,N_2767);
and U2829 (N_2829,N_2789,N_2762);
and U2830 (N_2830,N_2754,N_2753);
nand U2831 (N_2831,N_2764,N_2771);
nand U2832 (N_2832,N_2776,N_2783);
nand U2833 (N_2833,N_2763,N_2767);
or U2834 (N_2834,N_2767,N_2780);
nor U2835 (N_2835,N_2757,N_2771);
and U2836 (N_2836,N_2769,N_2795);
or U2837 (N_2837,N_2771,N_2750);
nor U2838 (N_2838,N_2770,N_2751);
and U2839 (N_2839,N_2781,N_2758);
and U2840 (N_2840,N_2793,N_2756);
nand U2841 (N_2841,N_2763,N_2785);
or U2842 (N_2842,N_2756,N_2795);
nand U2843 (N_2843,N_2771,N_2762);
or U2844 (N_2844,N_2773,N_2768);
nor U2845 (N_2845,N_2779,N_2785);
and U2846 (N_2846,N_2760,N_2787);
or U2847 (N_2847,N_2761,N_2750);
nand U2848 (N_2848,N_2788,N_2759);
and U2849 (N_2849,N_2773,N_2770);
nor U2850 (N_2850,N_2839,N_2836);
and U2851 (N_2851,N_2816,N_2806);
and U2852 (N_2852,N_2849,N_2846);
nand U2853 (N_2853,N_2848,N_2812);
or U2854 (N_2854,N_2817,N_2834);
nor U2855 (N_2855,N_2804,N_2831);
and U2856 (N_2856,N_2819,N_2838);
nor U2857 (N_2857,N_2818,N_2820);
and U2858 (N_2858,N_2815,N_2833);
and U2859 (N_2859,N_2829,N_2801);
or U2860 (N_2860,N_2845,N_2809);
and U2861 (N_2861,N_2830,N_2840);
and U2862 (N_2862,N_2813,N_2814);
or U2863 (N_2863,N_2837,N_2823);
and U2864 (N_2864,N_2825,N_2808);
and U2865 (N_2865,N_2844,N_2832);
nand U2866 (N_2866,N_2810,N_2847);
or U2867 (N_2867,N_2842,N_2802);
nor U2868 (N_2868,N_2843,N_2800);
or U2869 (N_2869,N_2824,N_2821);
nor U2870 (N_2870,N_2822,N_2835);
and U2871 (N_2871,N_2841,N_2811);
or U2872 (N_2872,N_2807,N_2827);
nand U2873 (N_2873,N_2826,N_2805);
and U2874 (N_2874,N_2828,N_2803);
and U2875 (N_2875,N_2807,N_2841);
or U2876 (N_2876,N_2845,N_2847);
nor U2877 (N_2877,N_2825,N_2843);
xor U2878 (N_2878,N_2839,N_2823);
xnor U2879 (N_2879,N_2804,N_2832);
nor U2880 (N_2880,N_2816,N_2845);
nor U2881 (N_2881,N_2804,N_2843);
xor U2882 (N_2882,N_2819,N_2802);
and U2883 (N_2883,N_2842,N_2834);
nand U2884 (N_2884,N_2808,N_2842);
xnor U2885 (N_2885,N_2812,N_2849);
nor U2886 (N_2886,N_2818,N_2841);
nor U2887 (N_2887,N_2832,N_2811);
nand U2888 (N_2888,N_2834,N_2818);
nand U2889 (N_2889,N_2829,N_2812);
nand U2890 (N_2890,N_2818,N_2833);
and U2891 (N_2891,N_2817,N_2807);
nand U2892 (N_2892,N_2836,N_2846);
nor U2893 (N_2893,N_2820,N_2805);
nor U2894 (N_2894,N_2846,N_2847);
or U2895 (N_2895,N_2800,N_2841);
nand U2896 (N_2896,N_2825,N_2834);
or U2897 (N_2897,N_2836,N_2834);
nand U2898 (N_2898,N_2806,N_2807);
xnor U2899 (N_2899,N_2824,N_2813);
nand U2900 (N_2900,N_2858,N_2875);
nor U2901 (N_2901,N_2855,N_2851);
nand U2902 (N_2902,N_2864,N_2870);
or U2903 (N_2903,N_2868,N_2854);
nand U2904 (N_2904,N_2883,N_2880);
or U2905 (N_2905,N_2890,N_2886);
nand U2906 (N_2906,N_2862,N_2884);
xor U2907 (N_2907,N_2893,N_2882);
xor U2908 (N_2908,N_2850,N_2881);
xnor U2909 (N_2909,N_2898,N_2876);
and U2910 (N_2910,N_2856,N_2866);
nand U2911 (N_2911,N_2891,N_2853);
and U2912 (N_2912,N_2896,N_2895);
nor U2913 (N_2913,N_2888,N_2877);
or U2914 (N_2914,N_2873,N_2859);
or U2915 (N_2915,N_2871,N_2889);
and U2916 (N_2916,N_2867,N_2860);
and U2917 (N_2917,N_2879,N_2857);
and U2918 (N_2918,N_2892,N_2865);
or U2919 (N_2919,N_2894,N_2863);
nand U2920 (N_2920,N_2897,N_2885);
nand U2921 (N_2921,N_2861,N_2852);
nor U2922 (N_2922,N_2874,N_2887);
and U2923 (N_2923,N_2899,N_2869);
or U2924 (N_2924,N_2878,N_2872);
nand U2925 (N_2925,N_2898,N_2890);
xnor U2926 (N_2926,N_2898,N_2874);
or U2927 (N_2927,N_2887,N_2851);
and U2928 (N_2928,N_2850,N_2867);
and U2929 (N_2929,N_2867,N_2884);
nor U2930 (N_2930,N_2857,N_2889);
nand U2931 (N_2931,N_2863,N_2850);
and U2932 (N_2932,N_2879,N_2893);
or U2933 (N_2933,N_2888,N_2887);
and U2934 (N_2934,N_2891,N_2877);
or U2935 (N_2935,N_2850,N_2869);
and U2936 (N_2936,N_2872,N_2899);
xor U2937 (N_2937,N_2885,N_2891);
and U2938 (N_2938,N_2862,N_2892);
or U2939 (N_2939,N_2864,N_2894);
and U2940 (N_2940,N_2882,N_2861);
and U2941 (N_2941,N_2862,N_2895);
and U2942 (N_2942,N_2857,N_2867);
and U2943 (N_2943,N_2873,N_2890);
and U2944 (N_2944,N_2861,N_2862);
nor U2945 (N_2945,N_2880,N_2866);
nor U2946 (N_2946,N_2881,N_2862);
or U2947 (N_2947,N_2874,N_2854);
nor U2948 (N_2948,N_2853,N_2856);
or U2949 (N_2949,N_2877,N_2861);
xor U2950 (N_2950,N_2916,N_2915);
nand U2951 (N_2951,N_2925,N_2923);
xor U2952 (N_2952,N_2910,N_2909);
nor U2953 (N_2953,N_2921,N_2933);
nand U2954 (N_2954,N_2901,N_2913);
nor U2955 (N_2955,N_2907,N_2906);
nand U2956 (N_2956,N_2926,N_2940);
and U2957 (N_2957,N_2914,N_2918);
and U2958 (N_2958,N_2908,N_2927);
nor U2959 (N_2959,N_2945,N_2922);
or U2960 (N_2960,N_2929,N_2930);
or U2961 (N_2961,N_2946,N_2920);
nand U2962 (N_2962,N_2941,N_2900);
nand U2963 (N_2963,N_2902,N_2931);
nand U2964 (N_2964,N_2934,N_2917);
nor U2965 (N_2965,N_2932,N_2911);
nor U2966 (N_2966,N_2936,N_2935);
nand U2967 (N_2967,N_2943,N_2939);
and U2968 (N_2968,N_2903,N_2924);
nor U2969 (N_2969,N_2904,N_2948);
nand U2970 (N_2970,N_2937,N_2919);
nor U2971 (N_2971,N_2947,N_2912);
or U2972 (N_2972,N_2928,N_2905);
nand U2973 (N_2973,N_2938,N_2949);
nand U2974 (N_2974,N_2942,N_2944);
or U2975 (N_2975,N_2931,N_2932);
and U2976 (N_2976,N_2946,N_2917);
or U2977 (N_2977,N_2947,N_2932);
and U2978 (N_2978,N_2946,N_2936);
nand U2979 (N_2979,N_2920,N_2909);
nand U2980 (N_2980,N_2909,N_2933);
xor U2981 (N_2981,N_2929,N_2910);
and U2982 (N_2982,N_2930,N_2947);
and U2983 (N_2983,N_2909,N_2926);
nor U2984 (N_2984,N_2945,N_2929);
xnor U2985 (N_2985,N_2925,N_2921);
and U2986 (N_2986,N_2906,N_2924);
and U2987 (N_2987,N_2907,N_2905);
xor U2988 (N_2988,N_2923,N_2920);
or U2989 (N_2989,N_2933,N_2944);
xnor U2990 (N_2990,N_2935,N_2944);
and U2991 (N_2991,N_2924,N_2914);
or U2992 (N_2992,N_2925,N_2915);
nand U2993 (N_2993,N_2900,N_2923);
and U2994 (N_2994,N_2916,N_2926);
nor U2995 (N_2995,N_2945,N_2947);
xor U2996 (N_2996,N_2917,N_2913);
and U2997 (N_2997,N_2935,N_2904);
and U2998 (N_2998,N_2911,N_2941);
xor U2999 (N_2999,N_2932,N_2940);
and UO_0 (O_0,N_2974,N_2994);
nor UO_1 (O_1,N_2992,N_2977);
nand UO_2 (O_2,N_2951,N_2962);
or UO_3 (O_3,N_2995,N_2993);
and UO_4 (O_4,N_2964,N_2961);
or UO_5 (O_5,N_2980,N_2952);
nand UO_6 (O_6,N_2967,N_2996);
or UO_7 (O_7,N_2986,N_2987);
or UO_8 (O_8,N_2968,N_2997);
nor UO_9 (O_9,N_2959,N_2960);
nand UO_10 (O_10,N_2976,N_2985);
nor UO_11 (O_11,N_2956,N_2950);
nor UO_12 (O_12,N_2990,N_2989);
or UO_13 (O_13,N_2955,N_2999);
or UO_14 (O_14,N_2983,N_2971);
xnor UO_15 (O_15,N_2969,N_2963);
nand UO_16 (O_16,N_2979,N_2957);
or UO_17 (O_17,N_2981,N_2988);
nand UO_18 (O_18,N_2954,N_2978);
nor UO_19 (O_19,N_2973,N_2965);
xor UO_20 (O_20,N_2953,N_2958);
or UO_21 (O_21,N_2998,N_2966);
and UO_22 (O_22,N_2984,N_2970);
or UO_23 (O_23,N_2991,N_2982);
nand UO_24 (O_24,N_2972,N_2975);
or UO_25 (O_25,N_2964,N_2987);
nor UO_26 (O_26,N_2998,N_2977);
nor UO_27 (O_27,N_2978,N_2950);
nand UO_28 (O_28,N_2989,N_2993);
nand UO_29 (O_29,N_2990,N_2966);
and UO_30 (O_30,N_2966,N_2981);
nor UO_31 (O_31,N_2970,N_2953);
or UO_32 (O_32,N_2996,N_2986);
nand UO_33 (O_33,N_2999,N_2978);
xor UO_34 (O_34,N_2957,N_2990);
nor UO_35 (O_35,N_2981,N_2968);
and UO_36 (O_36,N_2997,N_2989);
and UO_37 (O_37,N_2957,N_2996);
and UO_38 (O_38,N_2957,N_2987);
or UO_39 (O_39,N_2970,N_2963);
and UO_40 (O_40,N_2994,N_2988);
nand UO_41 (O_41,N_2973,N_2980);
or UO_42 (O_42,N_2972,N_2954);
or UO_43 (O_43,N_2995,N_2985);
nor UO_44 (O_44,N_2970,N_2996);
nand UO_45 (O_45,N_2955,N_2979);
and UO_46 (O_46,N_2989,N_2977);
and UO_47 (O_47,N_2962,N_2985);
nor UO_48 (O_48,N_2997,N_2990);
nor UO_49 (O_49,N_2972,N_2957);
and UO_50 (O_50,N_2976,N_2982);
nor UO_51 (O_51,N_2989,N_2953);
or UO_52 (O_52,N_2982,N_2966);
and UO_53 (O_53,N_2978,N_2976);
or UO_54 (O_54,N_2968,N_2965);
xnor UO_55 (O_55,N_2960,N_2999);
or UO_56 (O_56,N_2983,N_2990);
nand UO_57 (O_57,N_2953,N_2990);
and UO_58 (O_58,N_2988,N_2983);
nand UO_59 (O_59,N_2964,N_2967);
xor UO_60 (O_60,N_2972,N_2965);
nor UO_61 (O_61,N_2967,N_2973);
nand UO_62 (O_62,N_2953,N_2954);
and UO_63 (O_63,N_2978,N_2968);
xnor UO_64 (O_64,N_2973,N_2985);
and UO_65 (O_65,N_2953,N_2976);
nor UO_66 (O_66,N_2989,N_2964);
nor UO_67 (O_67,N_2995,N_2953);
and UO_68 (O_68,N_2996,N_2995);
and UO_69 (O_69,N_2999,N_2980);
nand UO_70 (O_70,N_2995,N_2963);
nor UO_71 (O_71,N_2992,N_2950);
or UO_72 (O_72,N_2990,N_2975);
nor UO_73 (O_73,N_2976,N_2967);
xnor UO_74 (O_74,N_2950,N_2963);
nand UO_75 (O_75,N_2997,N_2956);
or UO_76 (O_76,N_2982,N_2964);
and UO_77 (O_77,N_2969,N_2984);
nor UO_78 (O_78,N_2983,N_2996);
xor UO_79 (O_79,N_2970,N_2967);
and UO_80 (O_80,N_2953,N_2956);
xor UO_81 (O_81,N_2979,N_2960);
nor UO_82 (O_82,N_2967,N_2951);
nor UO_83 (O_83,N_2990,N_2950);
and UO_84 (O_84,N_2961,N_2975);
xor UO_85 (O_85,N_2991,N_2983);
nor UO_86 (O_86,N_2964,N_2992);
or UO_87 (O_87,N_2951,N_2985);
nor UO_88 (O_88,N_2984,N_2960);
or UO_89 (O_89,N_2973,N_2952);
xnor UO_90 (O_90,N_2954,N_2960);
xnor UO_91 (O_91,N_2999,N_2952);
and UO_92 (O_92,N_2982,N_2995);
nor UO_93 (O_93,N_2994,N_2976);
nor UO_94 (O_94,N_2969,N_2958);
nor UO_95 (O_95,N_2964,N_2981);
nor UO_96 (O_96,N_2952,N_2953);
or UO_97 (O_97,N_2975,N_2956);
xor UO_98 (O_98,N_2981,N_2955);
or UO_99 (O_99,N_2984,N_2977);
nand UO_100 (O_100,N_2974,N_2979);
nand UO_101 (O_101,N_2978,N_2956);
or UO_102 (O_102,N_2981,N_2965);
or UO_103 (O_103,N_2959,N_2975);
or UO_104 (O_104,N_2950,N_2988);
and UO_105 (O_105,N_2976,N_2983);
or UO_106 (O_106,N_2979,N_2967);
and UO_107 (O_107,N_2983,N_2980);
and UO_108 (O_108,N_2967,N_2995);
and UO_109 (O_109,N_2956,N_2973);
nand UO_110 (O_110,N_2981,N_2979);
and UO_111 (O_111,N_2969,N_2972);
nand UO_112 (O_112,N_2959,N_2963);
and UO_113 (O_113,N_2982,N_2983);
nand UO_114 (O_114,N_2959,N_2954);
nand UO_115 (O_115,N_2951,N_2996);
nor UO_116 (O_116,N_2967,N_2982);
nor UO_117 (O_117,N_2958,N_2950);
and UO_118 (O_118,N_2965,N_2971);
xnor UO_119 (O_119,N_2958,N_2985);
and UO_120 (O_120,N_2962,N_2979);
or UO_121 (O_121,N_2983,N_2987);
or UO_122 (O_122,N_2991,N_2968);
nor UO_123 (O_123,N_2952,N_2975);
and UO_124 (O_124,N_2995,N_2987);
nand UO_125 (O_125,N_2996,N_2984);
nand UO_126 (O_126,N_2996,N_2958);
nand UO_127 (O_127,N_2992,N_2985);
nand UO_128 (O_128,N_2963,N_2977);
nor UO_129 (O_129,N_2960,N_2997);
nor UO_130 (O_130,N_2990,N_2993);
nor UO_131 (O_131,N_2998,N_2984);
nor UO_132 (O_132,N_2976,N_2958);
xor UO_133 (O_133,N_2979,N_2958);
nor UO_134 (O_134,N_2952,N_2955);
and UO_135 (O_135,N_2969,N_2978);
or UO_136 (O_136,N_2969,N_2983);
nor UO_137 (O_137,N_2984,N_2975);
nand UO_138 (O_138,N_2998,N_2993);
or UO_139 (O_139,N_2958,N_2999);
and UO_140 (O_140,N_2991,N_2967);
xor UO_141 (O_141,N_2996,N_2998);
or UO_142 (O_142,N_2967,N_2955);
and UO_143 (O_143,N_2990,N_2959);
and UO_144 (O_144,N_2961,N_2965);
and UO_145 (O_145,N_2958,N_2954);
and UO_146 (O_146,N_2965,N_2976);
xnor UO_147 (O_147,N_2994,N_2996);
or UO_148 (O_148,N_2994,N_2979);
or UO_149 (O_149,N_2988,N_2970);
nor UO_150 (O_150,N_2971,N_2993);
or UO_151 (O_151,N_2953,N_2950);
or UO_152 (O_152,N_2957,N_2998);
or UO_153 (O_153,N_2960,N_2963);
or UO_154 (O_154,N_2985,N_2952);
and UO_155 (O_155,N_2987,N_2990);
or UO_156 (O_156,N_2998,N_2968);
or UO_157 (O_157,N_2987,N_2950);
nand UO_158 (O_158,N_2958,N_2984);
or UO_159 (O_159,N_2981,N_2982);
nor UO_160 (O_160,N_2999,N_2959);
or UO_161 (O_161,N_2966,N_2967);
xnor UO_162 (O_162,N_2958,N_2980);
nand UO_163 (O_163,N_2992,N_2954);
or UO_164 (O_164,N_2996,N_2963);
and UO_165 (O_165,N_2959,N_2987);
nand UO_166 (O_166,N_2961,N_2953);
or UO_167 (O_167,N_2985,N_2984);
nand UO_168 (O_168,N_2985,N_2969);
nor UO_169 (O_169,N_2996,N_2993);
nand UO_170 (O_170,N_2953,N_2998);
nand UO_171 (O_171,N_2993,N_2953);
and UO_172 (O_172,N_2982,N_2980);
and UO_173 (O_173,N_2965,N_2977);
nand UO_174 (O_174,N_2973,N_2996);
and UO_175 (O_175,N_2951,N_2952);
or UO_176 (O_176,N_2998,N_2987);
nand UO_177 (O_177,N_2979,N_2976);
and UO_178 (O_178,N_2990,N_2985);
and UO_179 (O_179,N_2978,N_2960);
and UO_180 (O_180,N_2982,N_2986);
or UO_181 (O_181,N_2965,N_2985);
nor UO_182 (O_182,N_2959,N_2957);
and UO_183 (O_183,N_2950,N_2957);
or UO_184 (O_184,N_2989,N_2999);
and UO_185 (O_185,N_2974,N_2952);
nor UO_186 (O_186,N_2950,N_2986);
and UO_187 (O_187,N_2994,N_2992);
nor UO_188 (O_188,N_2999,N_2997);
and UO_189 (O_189,N_2977,N_2961);
and UO_190 (O_190,N_2958,N_2987);
nor UO_191 (O_191,N_2986,N_2978);
or UO_192 (O_192,N_2980,N_2998);
nand UO_193 (O_193,N_2978,N_2966);
nor UO_194 (O_194,N_2992,N_2972);
or UO_195 (O_195,N_2983,N_2994);
or UO_196 (O_196,N_2966,N_2976);
or UO_197 (O_197,N_2974,N_2978);
nand UO_198 (O_198,N_2969,N_2977);
or UO_199 (O_199,N_2986,N_2994);
xor UO_200 (O_200,N_2968,N_2993);
nor UO_201 (O_201,N_2999,N_2969);
nor UO_202 (O_202,N_2977,N_2975);
or UO_203 (O_203,N_2979,N_2951);
nand UO_204 (O_204,N_2954,N_2988);
nor UO_205 (O_205,N_2966,N_2965);
or UO_206 (O_206,N_2958,N_2952);
nand UO_207 (O_207,N_2974,N_2987);
and UO_208 (O_208,N_2992,N_2999);
nor UO_209 (O_209,N_2999,N_2982);
nand UO_210 (O_210,N_2970,N_2960);
or UO_211 (O_211,N_2985,N_2959);
nor UO_212 (O_212,N_2956,N_2958);
or UO_213 (O_213,N_2985,N_2967);
nor UO_214 (O_214,N_2970,N_2954);
and UO_215 (O_215,N_2968,N_2985);
or UO_216 (O_216,N_2974,N_2998);
or UO_217 (O_217,N_2970,N_2993);
or UO_218 (O_218,N_2971,N_2973);
nor UO_219 (O_219,N_2972,N_2996);
nand UO_220 (O_220,N_2987,N_2956);
nand UO_221 (O_221,N_2966,N_2950);
nand UO_222 (O_222,N_2984,N_2989);
xor UO_223 (O_223,N_2958,N_2957);
nand UO_224 (O_224,N_2963,N_2984);
nor UO_225 (O_225,N_2997,N_2971);
or UO_226 (O_226,N_2961,N_2954);
nor UO_227 (O_227,N_2974,N_2959);
nand UO_228 (O_228,N_2990,N_2999);
or UO_229 (O_229,N_2968,N_2954);
or UO_230 (O_230,N_2957,N_2974);
nand UO_231 (O_231,N_2968,N_2976);
and UO_232 (O_232,N_2990,N_2956);
nor UO_233 (O_233,N_2973,N_2950);
nand UO_234 (O_234,N_2980,N_2989);
and UO_235 (O_235,N_2977,N_2997);
or UO_236 (O_236,N_2973,N_2997);
or UO_237 (O_237,N_2973,N_2955);
and UO_238 (O_238,N_2994,N_2978);
and UO_239 (O_239,N_2984,N_2951);
nor UO_240 (O_240,N_2988,N_2989);
nand UO_241 (O_241,N_2999,N_2962);
nand UO_242 (O_242,N_2961,N_2997);
and UO_243 (O_243,N_2983,N_2973);
and UO_244 (O_244,N_2984,N_2950);
nor UO_245 (O_245,N_2993,N_2987);
nand UO_246 (O_246,N_2951,N_2992);
xor UO_247 (O_247,N_2962,N_2995);
xor UO_248 (O_248,N_2999,N_2957);
nand UO_249 (O_249,N_2964,N_2968);
nor UO_250 (O_250,N_2952,N_2978);
nand UO_251 (O_251,N_2999,N_2951);
and UO_252 (O_252,N_2969,N_2965);
and UO_253 (O_253,N_2960,N_2971);
nor UO_254 (O_254,N_2964,N_2965);
nand UO_255 (O_255,N_2969,N_2951);
nand UO_256 (O_256,N_2959,N_2982);
nand UO_257 (O_257,N_2969,N_2986);
nor UO_258 (O_258,N_2968,N_2988);
or UO_259 (O_259,N_2965,N_2994);
and UO_260 (O_260,N_2988,N_2998);
nor UO_261 (O_261,N_2962,N_2980);
nand UO_262 (O_262,N_2970,N_2969);
xnor UO_263 (O_263,N_2972,N_2956);
nor UO_264 (O_264,N_2994,N_2969);
nor UO_265 (O_265,N_2956,N_2999);
or UO_266 (O_266,N_2956,N_2982);
and UO_267 (O_267,N_2965,N_2997);
nand UO_268 (O_268,N_2968,N_2982);
nand UO_269 (O_269,N_2990,N_2962);
xnor UO_270 (O_270,N_2957,N_2986);
and UO_271 (O_271,N_2973,N_2981);
or UO_272 (O_272,N_2979,N_2959);
or UO_273 (O_273,N_2969,N_2967);
or UO_274 (O_274,N_2999,N_2994);
nor UO_275 (O_275,N_2991,N_2979);
xnor UO_276 (O_276,N_2992,N_2971);
nand UO_277 (O_277,N_2985,N_2966);
and UO_278 (O_278,N_2955,N_2954);
and UO_279 (O_279,N_2954,N_2951);
and UO_280 (O_280,N_2961,N_2999);
and UO_281 (O_281,N_2984,N_2999);
nor UO_282 (O_282,N_2973,N_2987);
xor UO_283 (O_283,N_2988,N_2962);
xnor UO_284 (O_284,N_2950,N_2955);
xor UO_285 (O_285,N_2962,N_2970);
nor UO_286 (O_286,N_2962,N_2961);
nor UO_287 (O_287,N_2982,N_2957);
nand UO_288 (O_288,N_2983,N_2997);
nor UO_289 (O_289,N_2955,N_2959);
nand UO_290 (O_290,N_2969,N_2962);
or UO_291 (O_291,N_2995,N_2986);
nand UO_292 (O_292,N_2954,N_2977);
nor UO_293 (O_293,N_2987,N_2972);
and UO_294 (O_294,N_2978,N_2995);
nor UO_295 (O_295,N_2996,N_2965);
or UO_296 (O_296,N_2974,N_2976);
xnor UO_297 (O_297,N_2995,N_2988);
xnor UO_298 (O_298,N_2986,N_2984);
nor UO_299 (O_299,N_2980,N_2971);
or UO_300 (O_300,N_2952,N_2960);
nor UO_301 (O_301,N_2956,N_2954);
nand UO_302 (O_302,N_2953,N_2999);
or UO_303 (O_303,N_2951,N_2980);
nor UO_304 (O_304,N_2957,N_2984);
or UO_305 (O_305,N_2991,N_2964);
nand UO_306 (O_306,N_2975,N_2987);
and UO_307 (O_307,N_2974,N_2970);
nand UO_308 (O_308,N_2961,N_2994);
nand UO_309 (O_309,N_2991,N_2960);
nand UO_310 (O_310,N_2960,N_2988);
xnor UO_311 (O_311,N_2993,N_2961);
nor UO_312 (O_312,N_2972,N_2961);
nor UO_313 (O_313,N_2962,N_2992);
or UO_314 (O_314,N_2959,N_2951);
or UO_315 (O_315,N_2960,N_2982);
nor UO_316 (O_316,N_2957,N_2965);
nand UO_317 (O_317,N_2955,N_2960);
nand UO_318 (O_318,N_2951,N_2988);
nor UO_319 (O_319,N_2979,N_2966);
or UO_320 (O_320,N_2996,N_2968);
nor UO_321 (O_321,N_2980,N_2996);
and UO_322 (O_322,N_2966,N_2962);
nor UO_323 (O_323,N_2990,N_2991);
and UO_324 (O_324,N_2980,N_2956);
or UO_325 (O_325,N_2954,N_2974);
and UO_326 (O_326,N_2955,N_2982);
nand UO_327 (O_327,N_2979,N_2997);
or UO_328 (O_328,N_2984,N_2992);
and UO_329 (O_329,N_2999,N_2975);
nor UO_330 (O_330,N_2988,N_2976);
and UO_331 (O_331,N_2957,N_2985);
and UO_332 (O_332,N_2979,N_2998);
nor UO_333 (O_333,N_2976,N_2996);
nor UO_334 (O_334,N_2980,N_2957);
nor UO_335 (O_335,N_2967,N_2980);
or UO_336 (O_336,N_2978,N_2963);
nand UO_337 (O_337,N_2963,N_2998);
or UO_338 (O_338,N_2978,N_2982);
nor UO_339 (O_339,N_2975,N_2971);
xnor UO_340 (O_340,N_2964,N_2952);
nand UO_341 (O_341,N_2998,N_2961);
and UO_342 (O_342,N_2988,N_2979);
and UO_343 (O_343,N_2968,N_2975);
nor UO_344 (O_344,N_2980,N_2992);
or UO_345 (O_345,N_2988,N_2972);
and UO_346 (O_346,N_2974,N_2985);
and UO_347 (O_347,N_2986,N_2989);
or UO_348 (O_348,N_2993,N_2988);
nand UO_349 (O_349,N_2993,N_2957);
nand UO_350 (O_350,N_2991,N_2957);
nor UO_351 (O_351,N_2981,N_2990);
nor UO_352 (O_352,N_2983,N_2954);
nand UO_353 (O_353,N_2965,N_2988);
or UO_354 (O_354,N_2955,N_2953);
or UO_355 (O_355,N_2966,N_2960);
nor UO_356 (O_356,N_2973,N_2961);
nor UO_357 (O_357,N_2987,N_2982);
nand UO_358 (O_358,N_2956,N_2965);
and UO_359 (O_359,N_2970,N_2997);
or UO_360 (O_360,N_2962,N_2976);
nor UO_361 (O_361,N_2962,N_2952);
nor UO_362 (O_362,N_2950,N_2997);
and UO_363 (O_363,N_2997,N_2967);
or UO_364 (O_364,N_2965,N_2990);
or UO_365 (O_365,N_2990,N_2961);
and UO_366 (O_366,N_2950,N_2954);
and UO_367 (O_367,N_2963,N_2972);
nand UO_368 (O_368,N_2996,N_2966);
or UO_369 (O_369,N_2977,N_2987);
and UO_370 (O_370,N_2952,N_2997);
nor UO_371 (O_371,N_2978,N_2979);
or UO_372 (O_372,N_2958,N_2967);
nand UO_373 (O_373,N_2976,N_2995);
and UO_374 (O_374,N_2966,N_2991);
xor UO_375 (O_375,N_2974,N_2951);
nand UO_376 (O_376,N_2977,N_2990);
nor UO_377 (O_377,N_2962,N_2964);
xor UO_378 (O_378,N_2959,N_2972);
or UO_379 (O_379,N_2963,N_2992);
xnor UO_380 (O_380,N_2996,N_2960);
nand UO_381 (O_381,N_2960,N_2986);
nor UO_382 (O_382,N_2960,N_2977);
and UO_383 (O_383,N_2983,N_2977);
or UO_384 (O_384,N_2988,N_2952);
or UO_385 (O_385,N_2958,N_2974);
or UO_386 (O_386,N_2956,N_2957);
nand UO_387 (O_387,N_2986,N_2956);
nand UO_388 (O_388,N_2976,N_2971);
or UO_389 (O_389,N_2950,N_2981);
and UO_390 (O_390,N_2961,N_2981);
and UO_391 (O_391,N_2957,N_2975);
nand UO_392 (O_392,N_2974,N_2967);
and UO_393 (O_393,N_2960,N_2965);
nand UO_394 (O_394,N_2979,N_2970);
xor UO_395 (O_395,N_2968,N_2971);
nand UO_396 (O_396,N_2975,N_2950);
or UO_397 (O_397,N_2958,N_2990);
and UO_398 (O_398,N_2989,N_2954);
and UO_399 (O_399,N_2987,N_2999);
nand UO_400 (O_400,N_2995,N_2954);
and UO_401 (O_401,N_2953,N_2997);
nand UO_402 (O_402,N_2987,N_2962);
and UO_403 (O_403,N_2958,N_2977);
and UO_404 (O_404,N_2983,N_2960);
and UO_405 (O_405,N_2957,N_2952);
and UO_406 (O_406,N_2974,N_2988);
or UO_407 (O_407,N_2980,N_2986);
and UO_408 (O_408,N_2994,N_2962);
nor UO_409 (O_409,N_2987,N_2969);
nand UO_410 (O_410,N_2963,N_2966);
nor UO_411 (O_411,N_2978,N_2961);
or UO_412 (O_412,N_2973,N_2999);
or UO_413 (O_413,N_2974,N_2972);
or UO_414 (O_414,N_2951,N_2994);
nand UO_415 (O_415,N_2956,N_2993);
nor UO_416 (O_416,N_2980,N_2990);
or UO_417 (O_417,N_2988,N_2967);
or UO_418 (O_418,N_2966,N_2980);
nor UO_419 (O_419,N_2959,N_2973);
and UO_420 (O_420,N_2987,N_2971);
nand UO_421 (O_421,N_2998,N_2981);
nor UO_422 (O_422,N_2984,N_2980);
nand UO_423 (O_423,N_2975,N_2983);
nand UO_424 (O_424,N_2959,N_2992);
nand UO_425 (O_425,N_2965,N_2993);
nor UO_426 (O_426,N_2961,N_2988);
or UO_427 (O_427,N_2991,N_2993);
or UO_428 (O_428,N_2965,N_2991);
and UO_429 (O_429,N_2981,N_2971);
nor UO_430 (O_430,N_2985,N_2961);
nor UO_431 (O_431,N_2989,N_2972);
or UO_432 (O_432,N_2970,N_2999);
or UO_433 (O_433,N_2955,N_2996);
and UO_434 (O_434,N_2953,N_2980);
and UO_435 (O_435,N_2977,N_2976);
or UO_436 (O_436,N_2971,N_2994);
and UO_437 (O_437,N_2974,N_2991);
nor UO_438 (O_438,N_2963,N_2980);
xor UO_439 (O_439,N_2987,N_2988);
nand UO_440 (O_440,N_2989,N_2960);
and UO_441 (O_441,N_2989,N_2985);
xnor UO_442 (O_442,N_2997,N_2964);
and UO_443 (O_443,N_2972,N_2971);
nor UO_444 (O_444,N_2954,N_2999);
and UO_445 (O_445,N_2952,N_2959);
nand UO_446 (O_446,N_2969,N_2950);
nand UO_447 (O_447,N_2976,N_2991);
nand UO_448 (O_448,N_2978,N_2997);
nand UO_449 (O_449,N_2964,N_2972);
or UO_450 (O_450,N_2978,N_2989);
nor UO_451 (O_451,N_2971,N_2966);
or UO_452 (O_452,N_2969,N_2966);
and UO_453 (O_453,N_2977,N_2982);
or UO_454 (O_454,N_2977,N_2993);
or UO_455 (O_455,N_2986,N_2983);
nor UO_456 (O_456,N_2974,N_2975);
or UO_457 (O_457,N_2958,N_2995);
and UO_458 (O_458,N_2950,N_2976);
nand UO_459 (O_459,N_2963,N_2993);
nand UO_460 (O_460,N_2968,N_2999);
nor UO_461 (O_461,N_2957,N_2963);
and UO_462 (O_462,N_2952,N_2963);
nor UO_463 (O_463,N_2982,N_2952);
nor UO_464 (O_464,N_2953,N_2959);
and UO_465 (O_465,N_2986,N_2981);
or UO_466 (O_466,N_2976,N_2989);
nor UO_467 (O_467,N_2994,N_2966);
nor UO_468 (O_468,N_2960,N_2987);
and UO_469 (O_469,N_2991,N_2989);
and UO_470 (O_470,N_2957,N_2962);
xnor UO_471 (O_471,N_2951,N_2963);
or UO_472 (O_472,N_2962,N_2959);
nor UO_473 (O_473,N_2956,N_2983);
and UO_474 (O_474,N_2966,N_2959);
or UO_475 (O_475,N_2953,N_2985);
nand UO_476 (O_476,N_2970,N_2952);
and UO_477 (O_477,N_2956,N_2991);
nand UO_478 (O_478,N_2961,N_2960);
nor UO_479 (O_479,N_2995,N_2999);
nor UO_480 (O_480,N_2992,N_2970);
and UO_481 (O_481,N_2958,N_2965);
or UO_482 (O_482,N_2955,N_2984);
and UO_483 (O_483,N_2991,N_2970);
nand UO_484 (O_484,N_2972,N_2994);
nor UO_485 (O_485,N_2997,N_2980);
nor UO_486 (O_486,N_2989,N_2959);
or UO_487 (O_487,N_2957,N_2977);
and UO_488 (O_488,N_2996,N_2991);
and UO_489 (O_489,N_2989,N_2973);
or UO_490 (O_490,N_2990,N_2976);
nand UO_491 (O_491,N_2991,N_2959);
nor UO_492 (O_492,N_2972,N_2981);
and UO_493 (O_493,N_2967,N_2962);
or UO_494 (O_494,N_2978,N_2958);
nor UO_495 (O_495,N_2975,N_2963);
nor UO_496 (O_496,N_2960,N_2956);
nand UO_497 (O_497,N_2993,N_2974);
nor UO_498 (O_498,N_2979,N_2993);
xnor UO_499 (O_499,N_2963,N_2983);
endmodule