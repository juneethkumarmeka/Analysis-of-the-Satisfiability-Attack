module basic_500_3000_500_3_levels_5xor_8(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
xor U0 (N_0,In_322,In_80);
or U1 (N_1,In_319,In_251);
nor U2 (N_2,In_459,In_320);
or U3 (N_3,In_308,In_128);
nand U4 (N_4,In_480,In_197);
and U5 (N_5,In_187,In_254);
xnor U6 (N_6,In_160,In_272);
nand U7 (N_7,In_81,In_140);
nor U8 (N_8,In_49,In_38);
nor U9 (N_9,In_397,In_407);
nand U10 (N_10,In_321,In_178);
or U11 (N_11,In_203,In_284);
nand U12 (N_12,In_446,In_399);
and U13 (N_13,In_478,In_441);
and U14 (N_14,In_117,In_358);
nor U15 (N_15,In_253,In_483);
and U16 (N_16,In_70,In_157);
and U17 (N_17,In_278,In_408);
and U18 (N_18,In_40,In_427);
nand U19 (N_19,In_375,In_204);
nand U20 (N_20,In_115,In_12);
nand U21 (N_21,In_467,In_41);
and U22 (N_22,In_156,In_108);
nor U23 (N_23,In_418,In_307);
nand U24 (N_24,In_468,In_136);
nand U25 (N_25,In_63,In_111);
nand U26 (N_26,In_221,In_443);
nand U27 (N_27,In_166,In_464);
nor U28 (N_28,In_71,In_199);
or U29 (N_29,In_335,In_8);
nand U30 (N_30,In_231,In_410);
xnor U31 (N_31,In_9,In_318);
xnor U32 (N_32,In_305,In_444);
nor U33 (N_33,In_28,In_433);
xor U34 (N_34,In_473,In_466);
nor U35 (N_35,In_123,In_497);
xnor U36 (N_36,In_277,In_35);
nand U37 (N_37,In_104,In_499);
nand U38 (N_38,In_384,In_475);
and U39 (N_39,In_51,In_376);
nand U40 (N_40,In_202,In_491);
nand U41 (N_41,In_481,In_230);
xor U42 (N_42,In_207,In_2);
nand U43 (N_43,In_354,In_133);
nor U44 (N_44,In_243,In_169);
nor U45 (N_45,In_118,In_310);
xnor U46 (N_46,In_406,In_280);
or U47 (N_47,In_312,In_409);
and U48 (N_48,In_373,In_218);
and U49 (N_49,In_476,In_260);
nor U50 (N_50,In_292,In_14);
nor U51 (N_51,In_105,In_240);
nor U52 (N_52,In_442,In_485);
nand U53 (N_53,In_270,In_294);
xor U54 (N_54,In_90,In_282);
xnor U55 (N_55,In_364,In_402);
nand U56 (N_56,In_267,In_296);
and U57 (N_57,In_212,In_29);
or U58 (N_58,In_205,In_264);
nand U59 (N_59,In_227,In_55);
and U60 (N_60,In_224,In_208);
xnor U61 (N_61,In_153,In_439);
or U62 (N_62,In_216,In_431);
nand U63 (N_63,In_370,In_337);
and U64 (N_64,In_167,In_130);
or U65 (N_65,In_383,In_343);
and U66 (N_66,In_438,In_357);
nor U67 (N_67,In_366,In_299);
xnor U68 (N_68,In_365,In_0);
nor U69 (N_69,In_451,In_58);
or U70 (N_70,In_4,In_311);
nand U71 (N_71,In_33,In_26);
xor U72 (N_72,In_374,In_198);
and U73 (N_73,In_450,In_239);
or U74 (N_74,In_419,In_93);
and U75 (N_75,In_79,In_54);
nand U76 (N_76,In_263,In_132);
and U77 (N_77,In_392,In_189);
or U78 (N_78,In_182,In_168);
and U79 (N_79,In_349,In_31);
xnor U80 (N_80,In_414,In_64);
nand U81 (N_81,In_163,In_330);
or U82 (N_82,In_137,In_447);
nand U83 (N_83,In_423,In_211);
and U84 (N_84,In_200,In_440);
and U85 (N_85,In_285,In_269);
and U86 (N_86,In_43,In_185);
or U87 (N_87,In_302,In_390);
nand U88 (N_88,In_316,In_403);
xor U89 (N_89,In_232,In_395);
nand U90 (N_90,In_462,In_345);
nand U91 (N_91,In_146,In_323);
and U92 (N_92,In_449,In_333);
nand U93 (N_93,In_73,In_86);
or U94 (N_94,In_385,In_434);
xor U95 (N_95,In_255,In_44);
xnor U96 (N_96,In_192,In_77);
and U97 (N_97,In_448,In_340);
nand U98 (N_98,In_210,In_180);
nand U99 (N_99,In_122,In_252);
xnor U100 (N_100,In_469,In_68);
and U101 (N_101,In_482,In_454);
xor U102 (N_102,In_13,In_151);
nor U103 (N_103,In_334,In_114);
and U104 (N_104,In_6,In_173);
and U105 (N_105,In_209,In_194);
nor U106 (N_106,In_362,In_179);
nand U107 (N_107,In_184,In_257);
or U108 (N_108,In_386,In_304);
nand U109 (N_109,In_164,In_367);
nor U110 (N_110,In_155,In_486);
nor U111 (N_111,In_109,In_353);
xnor U112 (N_112,In_53,In_176);
or U113 (N_113,In_474,In_248);
or U114 (N_114,In_259,In_430);
or U115 (N_115,In_484,In_372);
nand U116 (N_116,In_127,In_15);
xor U117 (N_117,In_236,In_148);
or U118 (N_118,In_492,In_225);
nor U119 (N_119,In_351,In_181);
and U120 (N_120,In_88,In_387);
and U121 (N_121,In_400,In_341);
nand U122 (N_122,In_3,In_265);
or U123 (N_123,In_244,In_295);
or U124 (N_124,In_396,In_103);
nand U125 (N_125,In_107,In_241);
and U126 (N_126,In_139,In_289);
nor U127 (N_127,In_424,In_405);
and U128 (N_128,In_350,In_288);
nor U129 (N_129,In_287,In_315);
and U130 (N_130,In_411,In_471);
nand U131 (N_131,In_344,In_112);
or U132 (N_132,In_401,In_174);
nor U133 (N_133,In_61,In_177);
nand U134 (N_134,In_170,In_417);
nand U135 (N_135,In_477,In_391);
nand U136 (N_136,In_235,In_152);
and U137 (N_137,In_377,In_234);
nor U138 (N_138,In_47,In_124);
nand U139 (N_139,In_291,In_494);
or U140 (N_140,In_16,In_453);
and U141 (N_141,In_144,In_62);
nor U142 (N_142,In_110,In_456);
nor U143 (N_143,In_191,In_279);
xnor U144 (N_144,In_328,In_125);
and U145 (N_145,In_188,In_325);
and U146 (N_146,In_24,In_195);
and U147 (N_147,In_404,In_245);
or U148 (N_148,In_143,In_238);
nand U149 (N_149,In_247,In_416);
and U150 (N_150,In_332,In_298);
xnor U151 (N_151,In_271,In_363);
or U152 (N_152,In_92,In_313);
nand U153 (N_153,In_452,In_493);
nor U154 (N_154,In_134,In_129);
nor U155 (N_155,In_94,In_233);
nor U156 (N_156,In_57,In_22);
nand U157 (N_157,In_46,In_317);
or U158 (N_158,In_67,In_201);
or U159 (N_159,In_356,In_286);
or U160 (N_160,In_457,In_119);
nand U161 (N_161,In_488,In_72);
nand U162 (N_162,In_381,In_432);
xnor U163 (N_163,In_83,In_324);
and U164 (N_164,In_361,In_82);
nand U165 (N_165,In_135,In_470);
nor U166 (N_166,In_425,In_314);
nand U167 (N_167,In_283,In_226);
and U168 (N_168,In_274,In_113);
nor U169 (N_169,In_186,In_214);
or U170 (N_170,In_306,In_300);
nand U171 (N_171,In_25,In_266);
or U172 (N_172,In_309,In_102);
nand U173 (N_173,In_426,In_435);
nand U174 (N_174,In_37,In_489);
and U175 (N_175,In_19,In_23);
or U176 (N_176,In_355,In_27);
nand U177 (N_177,In_331,In_150);
nand U178 (N_178,In_219,In_99);
or U179 (N_179,In_162,In_45);
or U180 (N_180,In_342,In_360);
and U181 (N_181,In_420,In_159);
nor U182 (N_182,In_258,In_215);
nand U183 (N_183,In_217,In_290);
and U184 (N_184,In_172,In_413);
or U185 (N_185,In_141,In_213);
or U186 (N_186,In_422,In_154);
nand U187 (N_187,In_100,In_326);
nand U188 (N_188,In_175,In_59);
and U189 (N_189,In_429,In_242);
nand U190 (N_190,In_487,In_98);
nor U191 (N_191,In_145,In_281);
and U192 (N_192,In_412,In_495);
nor U193 (N_193,In_463,In_389);
and U194 (N_194,In_347,In_48);
or U195 (N_195,In_97,In_196);
nor U196 (N_196,In_398,In_50);
or U197 (N_197,In_415,In_7);
nand U198 (N_198,In_352,In_131);
nand U199 (N_199,In_479,In_262);
and U200 (N_200,In_327,In_348);
and U201 (N_201,In_297,In_78);
and U202 (N_202,In_303,In_490);
or U203 (N_203,In_445,In_149);
nand U204 (N_204,In_222,In_116);
or U205 (N_205,In_379,In_138);
and U206 (N_206,In_96,In_458);
nand U207 (N_207,In_436,In_5);
and U208 (N_208,In_74,In_18);
nand U209 (N_209,In_261,In_346);
nor U210 (N_210,In_34,In_101);
nand U211 (N_211,In_394,In_273);
and U212 (N_212,In_95,In_293);
and U213 (N_213,In_496,In_52);
nand U214 (N_214,In_21,In_11);
or U215 (N_215,In_223,In_369);
and U216 (N_216,In_87,In_190);
nand U217 (N_217,In_75,In_268);
or U218 (N_218,In_359,In_249);
nor U219 (N_219,In_371,In_161);
nor U220 (N_220,In_461,In_17);
or U221 (N_221,In_437,In_32);
xor U222 (N_222,In_142,In_421);
xnor U223 (N_223,In_76,In_1);
or U224 (N_224,In_339,In_158);
and U225 (N_225,In_256,In_193);
nor U226 (N_226,In_66,In_206);
nand U227 (N_227,In_380,In_65);
and U228 (N_228,In_10,In_120);
or U229 (N_229,In_147,In_84);
and U230 (N_230,In_121,In_36);
nand U231 (N_231,In_228,In_393);
xor U232 (N_232,In_378,In_338);
nand U233 (N_233,In_220,In_183);
nand U234 (N_234,In_165,In_498);
xor U235 (N_235,In_368,In_382);
xnor U236 (N_236,In_336,In_246);
nand U237 (N_237,In_237,In_42);
nor U238 (N_238,In_20,In_455);
or U239 (N_239,In_171,In_250);
nand U240 (N_240,In_301,In_465);
xnor U241 (N_241,In_60,In_460);
nand U242 (N_242,In_126,In_329);
nor U243 (N_243,In_85,In_275);
and U244 (N_244,In_276,In_428);
or U245 (N_245,In_229,In_91);
nor U246 (N_246,In_30,In_56);
or U247 (N_247,In_472,In_89);
nand U248 (N_248,In_69,In_388);
xor U249 (N_249,In_106,In_39);
or U250 (N_250,In_285,In_355);
nand U251 (N_251,In_52,In_224);
nor U252 (N_252,In_11,In_453);
nor U253 (N_253,In_373,In_383);
nor U254 (N_254,In_141,In_464);
xnor U255 (N_255,In_31,In_392);
or U256 (N_256,In_179,In_74);
or U257 (N_257,In_348,In_198);
nand U258 (N_258,In_55,In_122);
or U259 (N_259,In_480,In_343);
and U260 (N_260,In_451,In_394);
xnor U261 (N_261,In_2,In_74);
xor U262 (N_262,In_475,In_196);
nor U263 (N_263,In_62,In_235);
or U264 (N_264,In_155,In_139);
nand U265 (N_265,In_287,In_273);
nor U266 (N_266,In_32,In_373);
and U267 (N_267,In_294,In_157);
nor U268 (N_268,In_114,In_178);
nor U269 (N_269,In_494,In_142);
or U270 (N_270,In_134,In_82);
nor U271 (N_271,In_192,In_308);
xor U272 (N_272,In_97,In_285);
nand U273 (N_273,In_242,In_340);
or U274 (N_274,In_156,In_60);
nor U275 (N_275,In_283,In_196);
nand U276 (N_276,In_160,In_17);
or U277 (N_277,In_74,In_144);
or U278 (N_278,In_396,In_318);
nand U279 (N_279,In_294,In_258);
nor U280 (N_280,In_112,In_275);
xor U281 (N_281,In_462,In_156);
nand U282 (N_282,In_436,In_448);
nor U283 (N_283,In_379,In_260);
nand U284 (N_284,In_494,In_107);
or U285 (N_285,In_125,In_264);
xor U286 (N_286,In_126,In_283);
or U287 (N_287,In_51,In_46);
or U288 (N_288,In_392,In_302);
nand U289 (N_289,In_65,In_389);
or U290 (N_290,In_124,In_447);
nor U291 (N_291,In_185,In_322);
or U292 (N_292,In_179,In_434);
nor U293 (N_293,In_462,In_169);
nor U294 (N_294,In_335,In_250);
nor U295 (N_295,In_260,In_98);
nor U296 (N_296,In_215,In_424);
xor U297 (N_297,In_41,In_256);
nor U298 (N_298,In_428,In_400);
or U299 (N_299,In_45,In_383);
nand U300 (N_300,In_272,In_352);
or U301 (N_301,In_340,In_33);
xor U302 (N_302,In_191,In_185);
or U303 (N_303,In_332,In_376);
nand U304 (N_304,In_498,In_456);
and U305 (N_305,In_47,In_28);
and U306 (N_306,In_219,In_1);
xor U307 (N_307,In_20,In_192);
nor U308 (N_308,In_159,In_61);
and U309 (N_309,In_205,In_142);
nand U310 (N_310,In_13,In_339);
and U311 (N_311,In_287,In_382);
or U312 (N_312,In_214,In_314);
nand U313 (N_313,In_402,In_288);
xnor U314 (N_314,In_354,In_192);
and U315 (N_315,In_308,In_458);
xnor U316 (N_316,In_152,In_297);
and U317 (N_317,In_2,In_247);
or U318 (N_318,In_377,In_454);
nor U319 (N_319,In_492,In_29);
and U320 (N_320,In_327,In_42);
nand U321 (N_321,In_331,In_210);
and U322 (N_322,In_107,In_121);
or U323 (N_323,In_248,In_480);
nand U324 (N_324,In_422,In_200);
nor U325 (N_325,In_303,In_386);
nor U326 (N_326,In_1,In_488);
and U327 (N_327,In_472,In_65);
and U328 (N_328,In_414,In_405);
or U329 (N_329,In_73,In_117);
nor U330 (N_330,In_344,In_40);
nor U331 (N_331,In_307,In_217);
or U332 (N_332,In_343,In_42);
nor U333 (N_333,In_189,In_198);
or U334 (N_334,In_349,In_209);
nor U335 (N_335,In_365,In_2);
nand U336 (N_336,In_430,In_471);
or U337 (N_337,In_132,In_294);
and U338 (N_338,In_494,In_0);
and U339 (N_339,In_496,In_207);
and U340 (N_340,In_297,In_328);
nand U341 (N_341,In_340,In_430);
xor U342 (N_342,In_54,In_351);
and U343 (N_343,In_171,In_388);
nor U344 (N_344,In_2,In_246);
nand U345 (N_345,In_454,In_449);
nand U346 (N_346,In_6,In_299);
or U347 (N_347,In_63,In_349);
nor U348 (N_348,In_489,In_478);
nand U349 (N_349,In_320,In_238);
nor U350 (N_350,In_332,In_79);
or U351 (N_351,In_166,In_136);
or U352 (N_352,In_326,In_17);
nand U353 (N_353,In_423,In_310);
nor U354 (N_354,In_120,In_452);
nand U355 (N_355,In_268,In_197);
nor U356 (N_356,In_18,In_405);
nor U357 (N_357,In_24,In_138);
or U358 (N_358,In_5,In_234);
or U359 (N_359,In_488,In_185);
and U360 (N_360,In_376,In_342);
nor U361 (N_361,In_499,In_227);
xnor U362 (N_362,In_176,In_477);
and U363 (N_363,In_36,In_62);
nor U364 (N_364,In_328,In_251);
nand U365 (N_365,In_120,In_86);
and U366 (N_366,In_103,In_384);
xnor U367 (N_367,In_138,In_449);
nand U368 (N_368,In_212,In_23);
nor U369 (N_369,In_335,In_209);
or U370 (N_370,In_215,In_71);
nor U371 (N_371,In_185,In_360);
xnor U372 (N_372,In_346,In_52);
nor U373 (N_373,In_345,In_386);
nand U374 (N_374,In_321,In_487);
nand U375 (N_375,In_454,In_240);
nor U376 (N_376,In_351,In_466);
and U377 (N_377,In_94,In_85);
and U378 (N_378,In_316,In_89);
or U379 (N_379,In_482,In_165);
and U380 (N_380,In_326,In_210);
and U381 (N_381,In_331,In_322);
nor U382 (N_382,In_221,In_454);
nor U383 (N_383,In_486,In_183);
xnor U384 (N_384,In_168,In_67);
or U385 (N_385,In_291,In_269);
and U386 (N_386,In_399,In_331);
or U387 (N_387,In_159,In_126);
nand U388 (N_388,In_379,In_345);
nor U389 (N_389,In_481,In_152);
or U390 (N_390,In_301,In_398);
nand U391 (N_391,In_130,In_229);
nand U392 (N_392,In_69,In_14);
and U393 (N_393,In_231,In_258);
nor U394 (N_394,In_94,In_446);
nor U395 (N_395,In_194,In_21);
or U396 (N_396,In_398,In_35);
nand U397 (N_397,In_220,In_198);
or U398 (N_398,In_455,In_496);
nand U399 (N_399,In_16,In_254);
and U400 (N_400,In_254,In_326);
or U401 (N_401,In_310,In_384);
or U402 (N_402,In_482,In_43);
nand U403 (N_403,In_312,In_442);
or U404 (N_404,In_368,In_52);
and U405 (N_405,In_344,In_82);
or U406 (N_406,In_406,In_178);
and U407 (N_407,In_268,In_158);
nor U408 (N_408,In_428,In_3);
nor U409 (N_409,In_15,In_61);
nand U410 (N_410,In_103,In_177);
or U411 (N_411,In_472,In_334);
or U412 (N_412,In_38,In_295);
or U413 (N_413,In_431,In_150);
nand U414 (N_414,In_24,In_482);
xor U415 (N_415,In_288,In_343);
nor U416 (N_416,In_122,In_187);
or U417 (N_417,In_451,In_168);
nand U418 (N_418,In_437,In_158);
or U419 (N_419,In_129,In_410);
nor U420 (N_420,In_392,In_393);
and U421 (N_421,In_465,In_285);
nor U422 (N_422,In_113,In_360);
or U423 (N_423,In_325,In_261);
nand U424 (N_424,In_170,In_356);
nand U425 (N_425,In_298,In_351);
xnor U426 (N_426,In_284,In_80);
and U427 (N_427,In_202,In_88);
nand U428 (N_428,In_316,In_458);
nand U429 (N_429,In_249,In_167);
xnor U430 (N_430,In_141,In_126);
nand U431 (N_431,In_429,In_145);
and U432 (N_432,In_35,In_158);
nand U433 (N_433,In_28,In_56);
nor U434 (N_434,In_196,In_143);
nor U435 (N_435,In_241,In_487);
nor U436 (N_436,In_148,In_228);
and U437 (N_437,In_278,In_425);
xnor U438 (N_438,In_366,In_475);
nor U439 (N_439,In_334,In_162);
nand U440 (N_440,In_339,In_113);
or U441 (N_441,In_90,In_315);
nand U442 (N_442,In_397,In_457);
xnor U443 (N_443,In_76,In_6);
or U444 (N_444,In_407,In_376);
and U445 (N_445,In_231,In_455);
nor U446 (N_446,In_179,In_428);
or U447 (N_447,In_80,In_96);
nor U448 (N_448,In_449,In_298);
and U449 (N_449,In_239,In_276);
nor U450 (N_450,In_56,In_95);
nor U451 (N_451,In_131,In_65);
nor U452 (N_452,In_99,In_290);
and U453 (N_453,In_308,In_21);
or U454 (N_454,In_133,In_224);
and U455 (N_455,In_82,In_310);
or U456 (N_456,In_354,In_149);
nand U457 (N_457,In_449,In_306);
nand U458 (N_458,In_380,In_68);
or U459 (N_459,In_469,In_488);
nor U460 (N_460,In_196,In_485);
nor U461 (N_461,In_195,In_466);
nand U462 (N_462,In_72,In_218);
or U463 (N_463,In_266,In_381);
or U464 (N_464,In_351,In_468);
xnor U465 (N_465,In_310,In_140);
nor U466 (N_466,In_434,In_209);
nor U467 (N_467,In_112,In_176);
xnor U468 (N_468,In_360,In_274);
nor U469 (N_469,In_215,In_222);
nor U470 (N_470,In_476,In_413);
xor U471 (N_471,In_224,In_59);
nand U472 (N_472,In_137,In_201);
nand U473 (N_473,In_294,In_349);
xnor U474 (N_474,In_284,In_142);
and U475 (N_475,In_478,In_39);
or U476 (N_476,In_365,In_144);
nor U477 (N_477,In_290,In_11);
and U478 (N_478,In_30,In_80);
or U479 (N_479,In_266,In_101);
nor U480 (N_480,In_482,In_484);
or U481 (N_481,In_485,In_188);
nor U482 (N_482,In_390,In_19);
and U483 (N_483,In_472,In_132);
and U484 (N_484,In_116,In_136);
nor U485 (N_485,In_301,In_25);
nor U486 (N_486,In_402,In_422);
or U487 (N_487,In_263,In_177);
nand U488 (N_488,In_488,In_251);
nand U489 (N_489,In_494,In_394);
nor U490 (N_490,In_497,In_291);
xnor U491 (N_491,In_294,In_484);
and U492 (N_492,In_204,In_80);
nand U493 (N_493,In_35,In_206);
nor U494 (N_494,In_270,In_265);
xor U495 (N_495,In_25,In_42);
or U496 (N_496,In_391,In_378);
and U497 (N_497,In_371,In_257);
and U498 (N_498,In_209,In_228);
xnor U499 (N_499,In_404,In_63);
or U500 (N_500,In_396,In_120);
and U501 (N_501,In_370,In_183);
nor U502 (N_502,In_179,In_157);
and U503 (N_503,In_444,In_223);
or U504 (N_504,In_375,In_455);
xor U505 (N_505,In_132,In_89);
and U506 (N_506,In_257,In_297);
nand U507 (N_507,In_322,In_410);
nor U508 (N_508,In_277,In_107);
nor U509 (N_509,In_120,In_57);
nor U510 (N_510,In_120,In_198);
or U511 (N_511,In_77,In_22);
nand U512 (N_512,In_251,In_359);
xnor U513 (N_513,In_278,In_94);
or U514 (N_514,In_339,In_413);
and U515 (N_515,In_471,In_68);
or U516 (N_516,In_393,In_15);
nand U517 (N_517,In_213,In_340);
nand U518 (N_518,In_161,In_451);
nor U519 (N_519,In_87,In_204);
nor U520 (N_520,In_25,In_136);
and U521 (N_521,In_324,In_60);
or U522 (N_522,In_378,In_45);
and U523 (N_523,In_342,In_225);
or U524 (N_524,In_432,In_5);
nor U525 (N_525,In_483,In_192);
and U526 (N_526,In_450,In_336);
nand U527 (N_527,In_337,In_186);
xor U528 (N_528,In_230,In_459);
nor U529 (N_529,In_199,In_197);
nor U530 (N_530,In_475,In_402);
nand U531 (N_531,In_455,In_197);
nor U532 (N_532,In_357,In_467);
or U533 (N_533,In_291,In_157);
or U534 (N_534,In_87,In_150);
nand U535 (N_535,In_116,In_66);
xnor U536 (N_536,In_70,In_76);
or U537 (N_537,In_479,In_312);
nor U538 (N_538,In_305,In_121);
or U539 (N_539,In_24,In_336);
or U540 (N_540,In_106,In_121);
nand U541 (N_541,In_139,In_156);
or U542 (N_542,In_335,In_444);
nor U543 (N_543,In_82,In_473);
or U544 (N_544,In_327,In_401);
or U545 (N_545,In_381,In_51);
nor U546 (N_546,In_106,In_42);
xor U547 (N_547,In_484,In_492);
or U548 (N_548,In_425,In_20);
and U549 (N_549,In_65,In_2);
or U550 (N_550,In_425,In_198);
nor U551 (N_551,In_90,In_349);
or U552 (N_552,In_369,In_340);
nor U553 (N_553,In_279,In_299);
nand U554 (N_554,In_242,In_399);
or U555 (N_555,In_427,In_463);
and U556 (N_556,In_333,In_496);
nor U557 (N_557,In_104,In_114);
nor U558 (N_558,In_450,In_375);
or U559 (N_559,In_464,In_189);
nand U560 (N_560,In_175,In_185);
and U561 (N_561,In_360,In_33);
and U562 (N_562,In_457,In_427);
nand U563 (N_563,In_263,In_37);
nor U564 (N_564,In_4,In_140);
or U565 (N_565,In_466,In_34);
or U566 (N_566,In_407,In_201);
or U567 (N_567,In_295,In_313);
xnor U568 (N_568,In_43,In_237);
or U569 (N_569,In_58,In_487);
and U570 (N_570,In_219,In_303);
nor U571 (N_571,In_442,In_23);
nand U572 (N_572,In_173,In_165);
nor U573 (N_573,In_317,In_349);
nand U574 (N_574,In_492,In_72);
or U575 (N_575,In_266,In_45);
or U576 (N_576,In_360,In_111);
nand U577 (N_577,In_57,In_182);
nand U578 (N_578,In_405,In_199);
nor U579 (N_579,In_59,In_367);
and U580 (N_580,In_110,In_57);
and U581 (N_581,In_295,In_57);
nor U582 (N_582,In_189,In_142);
or U583 (N_583,In_487,In_82);
xnor U584 (N_584,In_194,In_349);
and U585 (N_585,In_464,In_136);
nor U586 (N_586,In_476,In_79);
nand U587 (N_587,In_203,In_186);
or U588 (N_588,In_438,In_137);
nand U589 (N_589,In_323,In_257);
nand U590 (N_590,In_189,In_37);
xor U591 (N_591,In_159,In_119);
nor U592 (N_592,In_75,In_32);
nor U593 (N_593,In_303,In_464);
nor U594 (N_594,In_165,In_373);
and U595 (N_595,In_275,In_374);
nor U596 (N_596,In_415,In_27);
or U597 (N_597,In_14,In_195);
and U598 (N_598,In_67,In_313);
nor U599 (N_599,In_281,In_102);
and U600 (N_600,In_340,In_142);
nand U601 (N_601,In_410,In_172);
and U602 (N_602,In_126,In_229);
or U603 (N_603,In_130,In_44);
nor U604 (N_604,In_483,In_190);
nor U605 (N_605,In_273,In_410);
nand U606 (N_606,In_204,In_21);
xor U607 (N_607,In_314,In_450);
nand U608 (N_608,In_27,In_65);
nor U609 (N_609,In_52,In_477);
xnor U610 (N_610,In_48,In_60);
or U611 (N_611,In_89,In_51);
and U612 (N_612,In_478,In_272);
nor U613 (N_613,In_436,In_413);
or U614 (N_614,In_273,In_438);
and U615 (N_615,In_27,In_345);
xor U616 (N_616,In_201,In_335);
or U617 (N_617,In_468,In_319);
nor U618 (N_618,In_339,In_119);
or U619 (N_619,In_299,In_4);
and U620 (N_620,In_174,In_128);
xor U621 (N_621,In_379,In_238);
nor U622 (N_622,In_443,In_72);
and U623 (N_623,In_22,In_13);
and U624 (N_624,In_221,In_164);
xnor U625 (N_625,In_110,In_297);
nor U626 (N_626,In_61,In_30);
and U627 (N_627,In_78,In_37);
nor U628 (N_628,In_422,In_403);
xnor U629 (N_629,In_74,In_260);
and U630 (N_630,In_423,In_55);
and U631 (N_631,In_299,In_26);
xor U632 (N_632,In_205,In_155);
nor U633 (N_633,In_57,In_215);
or U634 (N_634,In_200,In_56);
nand U635 (N_635,In_294,In_59);
nor U636 (N_636,In_483,In_74);
xnor U637 (N_637,In_145,In_407);
or U638 (N_638,In_259,In_138);
xnor U639 (N_639,In_365,In_318);
or U640 (N_640,In_94,In_181);
and U641 (N_641,In_42,In_206);
nand U642 (N_642,In_299,In_35);
nor U643 (N_643,In_139,In_462);
or U644 (N_644,In_379,In_241);
or U645 (N_645,In_451,In_45);
nor U646 (N_646,In_466,In_469);
xor U647 (N_647,In_22,In_336);
or U648 (N_648,In_430,In_135);
nand U649 (N_649,In_167,In_310);
or U650 (N_650,In_245,In_292);
nand U651 (N_651,In_444,In_330);
and U652 (N_652,In_469,In_498);
xnor U653 (N_653,In_134,In_108);
nor U654 (N_654,In_183,In_41);
or U655 (N_655,In_10,In_84);
nor U656 (N_656,In_455,In_441);
nand U657 (N_657,In_77,In_205);
nand U658 (N_658,In_370,In_342);
or U659 (N_659,In_161,In_458);
or U660 (N_660,In_250,In_170);
nand U661 (N_661,In_264,In_284);
xnor U662 (N_662,In_418,In_80);
or U663 (N_663,In_105,In_422);
and U664 (N_664,In_404,In_414);
or U665 (N_665,In_13,In_159);
nand U666 (N_666,In_355,In_167);
and U667 (N_667,In_383,In_410);
and U668 (N_668,In_103,In_397);
nor U669 (N_669,In_330,In_392);
and U670 (N_670,In_264,In_461);
nor U671 (N_671,In_443,In_194);
or U672 (N_672,In_424,In_286);
or U673 (N_673,In_157,In_419);
or U674 (N_674,In_370,In_485);
and U675 (N_675,In_168,In_178);
and U676 (N_676,In_218,In_417);
nand U677 (N_677,In_294,In_111);
nand U678 (N_678,In_222,In_173);
nor U679 (N_679,In_450,In_410);
and U680 (N_680,In_412,In_320);
nor U681 (N_681,In_398,In_207);
nand U682 (N_682,In_68,In_218);
nand U683 (N_683,In_280,In_129);
nand U684 (N_684,In_274,In_498);
nor U685 (N_685,In_266,In_94);
nor U686 (N_686,In_423,In_471);
nor U687 (N_687,In_428,In_5);
nor U688 (N_688,In_127,In_231);
nor U689 (N_689,In_423,In_54);
nand U690 (N_690,In_54,In_265);
nand U691 (N_691,In_282,In_273);
nand U692 (N_692,In_328,In_387);
nand U693 (N_693,In_158,In_252);
nand U694 (N_694,In_497,In_45);
nor U695 (N_695,In_255,In_4);
and U696 (N_696,In_368,In_196);
nor U697 (N_697,In_36,In_282);
or U698 (N_698,In_348,In_417);
or U699 (N_699,In_138,In_316);
and U700 (N_700,In_279,In_318);
and U701 (N_701,In_380,In_295);
nor U702 (N_702,In_417,In_443);
nand U703 (N_703,In_15,In_252);
or U704 (N_704,In_284,In_115);
nand U705 (N_705,In_46,In_493);
or U706 (N_706,In_486,In_467);
and U707 (N_707,In_378,In_191);
and U708 (N_708,In_268,In_238);
nand U709 (N_709,In_45,In_310);
and U710 (N_710,In_128,In_19);
nand U711 (N_711,In_425,In_326);
nor U712 (N_712,In_464,In_48);
and U713 (N_713,In_387,In_449);
and U714 (N_714,In_301,In_66);
nor U715 (N_715,In_10,In_317);
or U716 (N_716,In_265,In_167);
or U717 (N_717,In_143,In_477);
or U718 (N_718,In_485,In_191);
and U719 (N_719,In_90,In_305);
nand U720 (N_720,In_51,In_216);
or U721 (N_721,In_400,In_44);
or U722 (N_722,In_80,In_389);
and U723 (N_723,In_354,In_336);
nor U724 (N_724,In_412,In_286);
and U725 (N_725,In_410,In_266);
and U726 (N_726,In_445,In_208);
nand U727 (N_727,In_464,In_455);
and U728 (N_728,In_278,In_361);
nand U729 (N_729,In_27,In_184);
nand U730 (N_730,In_315,In_103);
nand U731 (N_731,In_493,In_485);
or U732 (N_732,In_267,In_158);
nor U733 (N_733,In_237,In_300);
nand U734 (N_734,In_235,In_105);
xor U735 (N_735,In_384,In_143);
xnor U736 (N_736,In_441,In_148);
nor U737 (N_737,In_320,In_170);
or U738 (N_738,In_444,In_70);
nor U739 (N_739,In_101,In_186);
or U740 (N_740,In_8,In_107);
nor U741 (N_741,In_352,In_290);
nor U742 (N_742,In_94,In_257);
and U743 (N_743,In_97,In_490);
and U744 (N_744,In_372,In_171);
nand U745 (N_745,In_419,In_159);
and U746 (N_746,In_318,In_31);
and U747 (N_747,In_313,In_432);
nand U748 (N_748,In_198,In_493);
nor U749 (N_749,In_54,In_137);
or U750 (N_750,In_388,In_15);
xor U751 (N_751,In_227,In_11);
nor U752 (N_752,In_164,In_440);
and U753 (N_753,In_92,In_36);
or U754 (N_754,In_47,In_110);
or U755 (N_755,In_41,In_234);
or U756 (N_756,In_238,In_171);
or U757 (N_757,In_116,In_64);
or U758 (N_758,In_168,In_317);
and U759 (N_759,In_343,In_214);
xnor U760 (N_760,In_361,In_83);
xor U761 (N_761,In_456,In_215);
nor U762 (N_762,In_198,In_209);
and U763 (N_763,In_406,In_155);
nand U764 (N_764,In_476,In_191);
nor U765 (N_765,In_29,In_419);
or U766 (N_766,In_365,In_253);
nor U767 (N_767,In_426,In_239);
nor U768 (N_768,In_16,In_108);
nand U769 (N_769,In_351,In_463);
nor U770 (N_770,In_17,In_488);
nor U771 (N_771,In_300,In_262);
nor U772 (N_772,In_196,In_460);
nand U773 (N_773,In_194,In_364);
and U774 (N_774,In_268,In_3);
nand U775 (N_775,In_216,In_263);
or U776 (N_776,In_285,In_150);
nor U777 (N_777,In_435,In_389);
or U778 (N_778,In_391,In_14);
or U779 (N_779,In_38,In_31);
xnor U780 (N_780,In_2,In_115);
and U781 (N_781,In_82,In_327);
nor U782 (N_782,In_158,In_33);
nand U783 (N_783,In_185,In_197);
nor U784 (N_784,In_446,In_69);
nor U785 (N_785,In_307,In_141);
or U786 (N_786,In_366,In_481);
and U787 (N_787,In_8,In_482);
nor U788 (N_788,In_96,In_210);
or U789 (N_789,In_183,In_12);
nand U790 (N_790,In_213,In_116);
and U791 (N_791,In_315,In_12);
xor U792 (N_792,In_325,In_165);
xnor U793 (N_793,In_28,In_305);
nor U794 (N_794,In_233,In_125);
and U795 (N_795,In_11,In_361);
and U796 (N_796,In_330,In_173);
nor U797 (N_797,In_246,In_350);
and U798 (N_798,In_254,In_41);
nor U799 (N_799,In_121,In_202);
nor U800 (N_800,In_345,In_434);
xor U801 (N_801,In_277,In_56);
nand U802 (N_802,In_472,In_307);
and U803 (N_803,In_169,In_111);
nor U804 (N_804,In_75,In_150);
or U805 (N_805,In_329,In_444);
nor U806 (N_806,In_422,In_77);
xnor U807 (N_807,In_427,In_291);
and U808 (N_808,In_22,In_145);
xor U809 (N_809,In_342,In_455);
nor U810 (N_810,In_300,In_271);
xor U811 (N_811,In_204,In_333);
and U812 (N_812,In_421,In_63);
nand U813 (N_813,In_252,In_434);
and U814 (N_814,In_355,In_441);
or U815 (N_815,In_55,In_497);
or U816 (N_816,In_2,In_88);
or U817 (N_817,In_287,In_421);
nor U818 (N_818,In_294,In_321);
or U819 (N_819,In_44,In_180);
nand U820 (N_820,In_31,In_49);
or U821 (N_821,In_488,In_485);
or U822 (N_822,In_181,In_168);
nand U823 (N_823,In_394,In_290);
and U824 (N_824,In_339,In_474);
nor U825 (N_825,In_437,In_216);
nor U826 (N_826,In_80,In_274);
nor U827 (N_827,In_81,In_166);
nand U828 (N_828,In_53,In_359);
nor U829 (N_829,In_122,In_291);
or U830 (N_830,In_342,In_89);
xnor U831 (N_831,In_31,In_198);
and U832 (N_832,In_88,In_173);
and U833 (N_833,In_451,In_68);
nand U834 (N_834,In_456,In_197);
and U835 (N_835,In_45,In_138);
nor U836 (N_836,In_393,In_287);
and U837 (N_837,In_325,In_209);
nand U838 (N_838,In_367,In_439);
nand U839 (N_839,In_2,In_471);
or U840 (N_840,In_316,In_320);
nand U841 (N_841,In_152,In_248);
nor U842 (N_842,In_477,In_227);
or U843 (N_843,In_398,In_477);
nor U844 (N_844,In_446,In_313);
nor U845 (N_845,In_73,In_15);
and U846 (N_846,In_396,In_434);
and U847 (N_847,In_178,In_20);
xor U848 (N_848,In_140,In_133);
nand U849 (N_849,In_97,In_241);
or U850 (N_850,In_123,In_179);
nand U851 (N_851,In_236,In_167);
and U852 (N_852,In_445,In_465);
nand U853 (N_853,In_420,In_381);
nor U854 (N_854,In_74,In_33);
nand U855 (N_855,In_401,In_143);
or U856 (N_856,In_436,In_454);
nor U857 (N_857,In_282,In_28);
or U858 (N_858,In_284,In_247);
and U859 (N_859,In_414,In_191);
and U860 (N_860,In_177,In_389);
or U861 (N_861,In_100,In_156);
or U862 (N_862,In_161,In_1);
and U863 (N_863,In_314,In_252);
or U864 (N_864,In_193,In_213);
nand U865 (N_865,In_10,In_186);
and U866 (N_866,In_398,In_376);
or U867 (N_867,In_348,In_122);
nand U868 (N_868,In_459,In_227);
nand U869 (N_869,In_432,In_286);
or U870 (N_870,In_69,In_332);
and U871 (N_871,In_428,In_333);
or U872 (N_872,In_434,In_494);
nor U873 (N_873,In_230,In_348);
and U874 (N_874,In_474,In_257);
or U875 (N_875,In_140,In_275);
nand U876 (N_876,In_243,In_284);
or U877 (N_877,In_80,In_482);
or U878 (N_878,In_382,In_358);
nor U879 (N_879,In_375,In_103);
or U880 (N_880,In_144,In_468);
nand U881 (N_881,In_241,In_495);
and U882 (N_882,In_122,In_104);
nor U883 (N_883,In_236,In_307);
nand U884 (N_884,In_269,In_304);
or U885 (N_885,In_90,In_17);
or U886 (N_886,In_222,In_317);
nor U887 (N_887,In_204,In_91);
or U888 (N_888,In_396,In_348);
or U889 (N_889,In_323,In_431);
nor U890 (N_890,In_490,In_92);
nor U891 (N_891,In_420,In_459);
xnor U892 (N_892,In_202,In_209);
or U893 (N_893,In_140,In_304);
nor U894 (N_894,In_419,In_258);
xnor U895 (N_895,In_33,In_346);
and U896 (N_896,In_167,In_469);
and U897 (N_897,In_313,In_183);
and U898 (N_898,In_322,In_128);
nor U899 (N_899,In_85,In_411);
or U900 (N_900,In_434,In_459);
nor U901 (N_901,In_431,In_303);
nor U902 (N_902,In_458,In_214);
xor U903 (N_903,In_114,In_256);
xor U904 (N_904,In_468,In_15);
xor U905 (N_905,In_434,In_399);
nand U906 (N_906,In_67,In_408);
and U907 (N_907,In_19,In_306);
and U908 (N_908,In_281,In_436);
nand U909 (N_909,In_293,In_118);
and U910 (N_910,In_193,In_353);
or U911 (N_911,In_49,In_280);
or U912 (N_912,In_483,In_399);
and U913 (N_913,In_254,In_376);
nand U914 (N_914,In_277,In_62);
nor U915 (N_915,In_8,In_201);
or U916 (N_916,In_265,In_451);
xor U917 (N_917,In_389,In_484);
or U918 (N_918,In_80,In_383);
nand U919 (N_919,In_457,In_262);
and U920 (N_920,In_346,In_0);
or U921 (N_921,In_340,In_444);
nor U922 (N_922,In_9,In_123);
or U923 (N_923,In_424,In_149);
or U924 (N_924,In_456,In_149);
nand U925 (N_925,In_196,In_49);
or U926 (N_926,In_8,In_499);
nor U927 (N_927,In_78,In_412);
and U928 (N_928,In_176,In_413);
or U929 (N_929,In_405,In_176);
nor U930 (N_930,In_208,In_298);
or U931 (N_931,In_71,In_20);
or U932 (N_932,In_309,In_483);
xnor U933 (N_933,In_357,In_124);
nand U934 (N_934,In_107,In_257);
or U935 (N_935,In_160,In_156);
xnor U936 (N_936,In_291,In_473);
and U937 (N_937,In_55,In_337);
or U938 (N_938,In_287,In_229);
nor U939 (N_939,In_157,In_45);
nor U940 (N_940,In_373,In_102);
nor U941 (N_941,In_291,In_387);
or U942 (N_942,In_279,In_314);
nor U943 (N_943,In_73,In_491);
nor U944 (N_944,In_164,In_498);
and U945 (N_945,In_216,In_131);
nor U946 (N_946,In_426,In_3);
and U947 (N_947,In_268,In_370);
or U948 (N_948,In_58,In_125);
and U949 (N_949,In_47,In_440);
or U950 (N_950,In_61,In_367);
nor U951 (N_951,In_343,In_193);
nor U952 (N_952,In_200,In_469);
or U953 (N_953,In_405,In_61);
nor U954 (N_954,In_237,In_219);
and U955 (N_955,In_45,In_87);
or U956 (N_956,In_272,In_156);
nand U957 (N_957,In_469,In_208);
and U958 (N_958,In_334,In_466);
and U959 (N_959,In_465,In_175);
nor U960 (N_960,In_487,In_290);
and U961 (N_961,In_383,In_200);
and U962 (N_962,In_233,In_389);
and U963 (N_963,In_151,In_117);
nand U964 (N_964,In_401,In_57);
and U965 (N_965,In_129,In_175);
and U966 (N_966,In_43,In_335);
nand U967 (N_967,In_332,In_102);
or U968 (N_968,In_208,In_423);
nand U969 (N_969,In_447,In_326);
nand U970 (N_970,In_82,In_434);
nand U971 (N_971,In_63,In_356);
or U972 (N_972,In_362,In_349);
nand U973 (N_973,In_334,In_141);
nor U974 (N_974,In_414,In_166);
and U975 (N_975,In_228,In_417);
or U976 (N_976,In_52,In_473);
nor U977 (N_977,In_64,In_452);
or U978 (N_978,In_323,In_205);
nor U979 (N_979,In_364,In_426);
nor U980 (N_980,In_314,In_477);
or U981 (N_981,In_91,In_451);
nor U982 (N_982,In_368,In_436);
nor U983 (N_983,In_163,In_315);
or U984 (N_984,In_224,In_142);
nand U985 (N_985,In_408,In_47);
nor U986 (N_986,In_401,In_29);
or U987 (N_987,In_348,In_183);
nor U988 (N_988,In_214,In_451);
nand U989 (N_989,In_326,In_352);
and U990 (N_990,In_92,In_334);
or U991 (N_991,In_407,In_452);
and U992 (N_992,In_202,In_487);
nor U993 (N_993,In_50,In_305);
xor U994 (N_994,In_346,In_355);
nand U995 (N_995,In_467,In_426);
nand U996 (N_996,In_254,In_344);
nand U997 (N_997,In_5,In_275);
or U998 (N_998,In_243,In_31);
nor U999 (N_999,In_241,In_142);
nand U1000 (N_1000,N_590,N_287);
or U1001 (N_1001,N_88,N_481);
xnor U1002 (N_1002,N_114,N_189);
nand U1003 (N_1003,N_636,N_520);
nand U1004 (N_1004,N_126,N_196);
nand U1005 (N_1005,N_978,N_664);
nor U1006 (N_1006,N_312,N_187);
and U1007 (N_1007,N_282,N_412);
nor U1008 (N_1008,N_25,N_902);
nor U1009 (N_1009,N_401,N_610);
or U1010 (N_1010,N_491,N_709);
or U1011 (N_1011,N_713,N_324);
or U1012 (N_1012,N_885,N_293);
or U1013 (N_1013,N_766,N_23);
or U1014 (N_1014,N_964,N_962);
or U1015 (N_1015,N_302,N_743);
nand U1016 (N_1016,N_638,N_209);
nor U1017 (N_1017,N_784,N_987);
and U1018 (N_1018,N_525,N_202);
nand U1019 (N_1019,N_516,N_977);
and U1020 (N_1020,N_304,N_912);
nor U1021 (N_1021,N_795,N_315);
nor U1022 (N_1022,N_266,N_283);
nand U1023 (N_1023,N_71,N_53);
nor U1024 (N_1024,N_985,N_618);
or U1025 (N_1025,N_915,N_949);
xor U1026 (N_1026,N_583,N_191);
nor U1027 (N_1027,N_635,N_518);
nor U1028 (N_1028,N_899,N_205);
nor U1029 (N_1029,N_248,N_591);
or U1030 (N_1030,N_323,N_46);
nor U1031 (N_1031,N_983,N_757);
nand U1032 (N_1032,N_980,N_846);
nor U1033 (N_1033,N_68,N_767);
nor U1034 (N_1034,N_479,N_810);
and U1035 (N_1035,N_670,N_627);
and U1036 (N_1036,N_808,N_519);
nand U1037 (N_1037,N_931,N_448);
nand U1038 (N_1038,N_669,N_44);
nor U1039 (N_1039,N_845,N_415);
xor U1040 (N_1040,N_442,N_177);
and U1041 (N_1041,N_373,N_891);
and U1042 (N_1042,N_629,N_914);
or U1043 (N_1043,N_489,N_511);
and U1044 (N_1044,N_19,N_622);
or U1045 (N_1045,N_289,N_830);
or U1046 (N_1046,N_486,N_544);
nand U1047 (N_1047,N_600,N_298);
nor U1048 (N_1048,N_819,N_596);
and U1049 (N_1049,N_361,N_309);
and U1050 (N_1050,N_346,N_395);
nor U1051 (N_1051,N_505,N_894);
or U1052 (N_1052,N_477,N_545);
nor U1053 (N_1053,N_413,N_913);
nor U1054 (N_1054,N_90,N_443);
nor U1055 (N_1055,N_50,N_769);
xnor U1056 (N_1056,N_929,N_497);
nand U1057 (N_1057,N_955,N_39);
nand U1058 (N_1058,N_563,N_349);
or U1059 (N_1059,N_762,N_946);
and U1060 (N_1060,N_262,N_49);
or U1061 (N_1061,N_982,N_848);
and U1062 (N_1062,N_554,N_786);
nand U1063 (N_1063,N_728,N_605);
and U1064 (N_1064,N_437,N_716);
or U1065 (N_1065,N_421,N_33);
xor U1066 (N_1066,N_774,N_83);
nand U1067 (N_1067,N_110,N_753);
nand U1068 (N_1068,N_847,N_75);
nor U1069 (N_1069,N_6,N_495);
nor U1070 (N_1070,N_671,N_738);
nand U1071 (N_1071,N_934,N_700);
xor U1072 (N_1072,N_678,N_322);
nor U1073 (N_1073,N_707,N_739);
or U1074 (N_1074,N_483,N_514);
and U1075 (N_1075,N_295,N_211);
nor U1076 (N_1076,N_195,N_103);
or U1077 (N_1077,N_122,N_811);
nand U1078 (N_1078,N_468,N_536);
nand U1079 (N_1079,N_956,N_156);
or U1080 (N_1080,N_697,N_508);
nand U1081 (N_1081,N_952,N_278);
nand U1082 (N_1082,N_95,N_470);
xnor U1083 (N_1083,N_105,N_822);
nand U1084 (N_1084,N_300,N_372);
nor U1085 (N_1085,N_921,N_216);
or U1086 (N_1086,N_995,N_67);
nor U1087 (N_1087,N_759,N_609);
and U1088 (N_1088,N_788,N_364);
or U1089 (N_1089,N_318,N_267);
nand U1090 (N_1090,N_127,N_906);
and U1091 (N_1091,N_20,N_532);
or U1092 (N_1092,N_128,N_258);
xor U1093 (N_1093,N_623,N_782);
nand U1094 (N_1094,N_389,N_192);
nor U1095 (N_1095,N_938,N_166);
and U1096 (N_1096,N_581,N_953);
xnor U1097 (N_1097,N_65,N_644);
nand U1098 (N_1098,N_310,N_319);
nand U1099 (N_1099,N_332,N_221);
or U1100 (N_1100,N_367,N_746);
nand U1101 (N_1101,N_555,N_909);
or U1102 (N_1102,N_675,N_719);
or U1103 (N_1103,N_425,N_167);
nand U1104 (N_1104,N_129,N_223);
and U1105 (N_1105,N_186,N_15);
nand U1106 (N_1106,N_578,N_735);
nand U1107 (N_1107,N_377,N_106);
nand U1108 (N_1108,N_341,N_198);
nor U1109 (N_1109,N_390,N_557);
nor U1110 (N_1110,N_246,N_732);
and U1111 (N_1111,N_397,N_427);
and U1112 (N_1112,N_131,N_445);
xnor U1113 (N_1113,N_659,N_577);
or U1114 (N_1114,N_244,N_641);
and U1115 (N_1115,N_856,N_776);
nor U1116 (N_1116,N_14,N_572);
or U1117 (N_1117,N_604,N_547);
and U1118 (N_1118,N_475,N_918);
or U1119 (N_1119,N_273,N_500);
and U1120 (N_1120,N_523,N_614);
xor U1121 (N_1121,N_376,N_344);
nand U1122 (N_1122,N_967,N_869);
or U1123 (N_1123,N_958,N_797);
nor U1124 (N_1124,N_923,N_417);
and U1125 (N_1125,N_109,N_630);
nand U1126 (N_1126,N_657,N_889);
nor U1127 (N_1127,N_580,N_676);
and U1128 (N_1128,N_893,N_998);
or U1129 (N_1129,N_5,N_655);
nor U1130 (N_1130,N_613,N_506);
nand U1131 (N_1131,N_271,N_907);
nand U1132 (N_1132,N_8,N_140);
nor U1133 (N_1133,N_194,N_729);
nor U1134 (N_1134,N_997,N_854);
nor U1135 (N_1135,N_178,N_540);
xnor U1136 (N_1136,N_690,N_803);
nand U1137 (N_1137,N_683,N_102);
nor U1138 (N_1138,N_615,N_538);
or U1139 (N_1139,N_818,N_74);
and U1140 (N_1140,N_203,N_992);
and U1141 (N_1141,N_450,N_237);
or U1142 (N_1142,N_134,N_524);
and U1143 (N_1143,N_159,N_825);
or U1144 (N_1144,N_687,N_496);
and U1145 (N_1145,N_616,N_763);
or U1146 (N_1146,N_552,N_502);
nand U1147 (N_1147,N_317,N_787);
and U1148 (N_1148,N_994,N_688);
nand U1149 (N_1149,N_841,N_488);
nor U1150 (N_1150,N_418,N_601);
and U1151 (N_1151,N_84,N_794);
or U1152 (N_1152,N_135,N_227);
xnor U1153 (N_1153,N_255,N_404);
nand U1154 (N_1154,N_462,N_781);
or U1155 (N_1155,N_214,N_241);
nor U1156 (N_1156,N_245,N_594);
and U1157 (N_1157,N_408,N_16);
and U1158 (N_1158,N_922,N_990);
nor U1159 (N_1159,N_272,N_467);
and U1160 (N_1160,N_370,N_855);
nor U1161 (N_1161,N_213,N_316);
nand U1162 (N_1162,N_951,N_175);
nand U1163 (N_1163,N_9,N_829);
or U1164 (N_1164,N_78,N_446);
and U1165 (N_1165,N_558,N_228);
xor U1166 (N_1166,N_111,N_896);
and U1167 (N_1167,N_264,N_858);
or U1168 (N_1168,N_619,N_490);
or U1169 (N_1169,N_568,N_865);
nor U1170 (N_1170,N_62,N_459);
and U1171 (N_1171,N_147,N_586);
nor U1172 (N_1172,N_606,N_0);
or U1173 (N_1173,N_1,N_742);
xor U1174 (N_1174,N_338,N_832);
nor U1175 (N_1175,N_268,N_851);
or U1176 (N_1176,N_56,N_363);
nand U1177 (N_1177,N_179,N_275);
nand U1178 (N_1178,N_441,N_579);
nor U1179 (N_1179,N_764,N_259);
or U1180 (N_1180,N_703,N_222);
and U1181 (N_1181,N_457,N_335);
xnor U1182 (N_1182,N_919,N_232);
or U1183 (N_1183,N_464,N_809);
nand U1184 (N_1184,N_996,N_679);
xor U1185 (N_1185,N_837,N_460);
or U1186 (N_1186,N_790,N_651);
nor U1187 (N_1187,N_770,N_513);
nand U1188 (N_1188,N_650,N_307);
and U1189 (N_1189,N_368,N_168);
or U1190 (N_1190,N_597,N_559);
and U1191 (N_1191,N_589,N_362);
or U1192 (N_1192,N_151,N_603);
and U1193 (N_1193,N_296,N_119);
and U1194 (N_1194,N_94,N_354);
nor U1195 (N_1195,N_290,N_720);
nor U1196 (N_1196,N_561,N_176);
nor U1197 (N_1197,N_291,N_173);
xnor U1198 (N_1198,N_117,N_836);
nand U1199 (N_1199,N_874,N_806);
or U1200 (N_1200,N_706,N_939);
xnor U1201 (N_1201,N_29,N_643);
and U1202 (N_1202,N_416,N_940);
nand U1203 (N_1203,N_576,N_55);
or U1204 (N_1204,N_252,N_394);
nor U1205 (N_1205,N_21,N_886);
or U1206 (N_1206,N_485,N_469);
nor U1207 (N_1207,N_433,N_101);
nor U1208 (N_1208,N_682,N_972);
xor U1209 (N_1209,N_286,N_263);
nor U1210 (N_1210,N_727,N_903);
nand U1211 (N_1211,N_123,N_36);
or U1212 (N_1212,N_748,N_3);
xor U1213 (N_1213,N_331,N_593);
and U1214 (N_1214,N_645,N_718);
or U1215 (N_1215,N_747,N_717);
and U1216 (N_1216,N_43,N_814);
or U1217 (N_1217,N_393,N_58);
xor U1218 (N_1218,N_897,N_342);
nor U1219 (N_1219,N_145,N_699);
and U1220 (N_1220,N_306,N_327);
nor U1221 (N_1221,N_183,N_498);
nand U1222 (N_1222,N_761,N_235);
nor U1223 (N_1223,N_208,N_440);
or U1224 (N_1224,N_883,N_715);
nand U1225 (N_1225,N_569,N_64);
nand U1226 (N_1226,N_878,N_862);
nor U1227 (N_1227,N_741,N_207);
or U1228 (N_1228,N_725,N_24);
or U1229 (N_1229,N_924,N_799);
nand U1230 (N_1230,N_269,N_69);
or U1231 (N_1231,N_824,N_672);
xor U1232 (N_1232,N_900,N_705);
nor U1233 (N_1233,N_857,N_981);
or U1234 (N_1234,N_936,N_750);
xnor U1235 (N_1235,N_432,N_60);
and U1236 (N_1236,N_154,N_438);
and U1237 (N_1237,N_484,N_882);
nand U1238 (N_1238,N_113,N_100);
and U1239 (N_1239,N_772,N_850);
or U1240 (N_1240,N_652,N_257);
or U1241 (N_1241,N_371,N_355);
nand U1242 (N_1242,N_261,N_815);
nand U1243 (N_1243,N_337,N_551);
nand U1244 (N_1244,N_311,N_11);
nor U1245 (N_1245,N_584,N_963);
nor U1246 (N_1246,N_108,N_30);
xnor U1247 (N_1247,N_308,N_968);
nor U1248 (N_1248,N_736,N_796);
nand U1249 (N_1249,N_357,N_334);
nor U1250 (N_1250,N_861,N_454);
and U1251 (N_1251,N_740,N_82);
nor U1252 (N_1252,N_144,N_439);
or U1253 (N_1253,N_132,N_904);
xor U1254 (N_1254,N_190,N_633);
or U1255 (N_1255,N_365,N_860);
xnor U1256 (N_1256,N_231,N_107);
nand U1257 (N_1257,N_637,N_406);
nor U1258 (N_1258,N_866,N_838);
nand U1259 (N_1259,N_428,N_158);
nor U1260 (N_1260,N_778,N_667);
or U1261 (N_1261,N_476,N_564);
nor U1262 (N_1262,N_98,N_607);
and U1263 (N_1263,N_386,N_353);
nor U1264 (N_1264,N_141,N_930);
and U1265 (N_1265,N_169,N_546);
xnor U1266 (N_1266,N_116,N_164);
or U1267 (N_1267,N_292,N_431);
nor U1268 (N_1268,N_347,N_971);
xor U1269 (N_1269,N_754,N_149);
and U1270 (N_1270,N_384,N_723);
nor U1271 (N_1271,N_876,N_321);
xnor U1272 (N_1272,N_798,N_553);
nand U1273 (N_1273,N_711,N_396);
nand U1274 (N_1274,N_943,N_684);
nand U1275 (N_1275,N_649,N_693);
or U1276 (N_1276,N_225,N_61);
nand U1277 (N_1277,N_961,N_674);
and U1278 (N_1278,N_574,N_239);
or U1279 (N_1279,N_453,N_420);
or U1280 (N_1280,N_828,N_632);
xnor U1281 (N_1281,N_256,N_812);
and U1282 (N_1282,N_330,N_369);
nor U1283 (N_1283,N_621,N_602);
and U1284 (N_1284,N_382,N_260);
or U1285 (N_1285,N_592,N_12);
or U1286 (N_1286,N_45,N_533);
nand U1287 (N_1287,N_28,N_405);
nand U1288 (N_1288,N_480,N_165);
or U1289 (N_1289,N_712,N_426);
or U1290 (N_1290,N_136,N_96);
xnor U1291 (N_1291,N_388,N_285);
nor U1292 (N_1292,N_531,N_66);
or U1293 (N_1293,N_451,N_539);
nand U1294 (N_1294,N_756,N_463);
nor U1295 (N_1295,N_240,N_352);
and U1296 (N_1296,N_104,N_343);
and U1297 (N_1297,N_152,N_724);
and U1298 (N_1298,N_146,N_137);
nor U1299 (N_1299,N_242,N_701);
nand U1300 (N_1300,N_698,N_400);
or U1301 (N_1301,N_387,N_410);
or U1302 (N_1302,N_466,N_336);
and U1303 (N_1303,N_562,N_91);
and U1304 (N_1304,N_625,N_379);
or U1305 (N_1305,N_478,N_646);
and U1306 (N_1306,N_22,N_853);
and U1307 (N_1307,N_901,N_399);
and U1308 (N_1308,N_38,N_932);
nand U1309 (N_1309,N_2,N_270);
and U1310 (N_1310,N_251,N_328);
or U1311 (N_1311,N_570,N_305);
or U1312 (N_1312,N_966,N_93);
nor U1313 (N_1313,N_503,N_473);
and U1314 (N_1314,N_366,N_668);
and U1315 (N_1315,N_945,N_429);
and U1316 (N_1316,N_247,N_92);
or U1317 (N_1317,N_7,N_608);
nor U1318 (N_1318,N_991,N_455);
nor U1319 (N_1319,N_849,N_771);
or U1320 (N_1320,N_360,N_765);
nand U1321 (N_1321,N_188,N_157);
nand U1322 (N_1322,N_805,N_686);
nand U1323 (N_1323,N_121,N_863);
nor U1324 (N_1324,N_494,N_634);
nand U1325 (N_1325,N_517,N_72);
nor U1326 (N_1326,N_734,N_654);
or U1327 (N_1327,N_656,N_695);
nor U1328 (N_1328,N_910,N_345);
nand U1329 (N_1329,N_976,N_852);
xor U1330 (N_1330,N_378,N_582);
nand U1331 (N_1331,N_447,N_556);
nor U1332 (N_1332,N_884,N_947);
nand U1333 (N_1333,N_138,N_325);
nand U1334 (N_1334,N_521,N_880);
and U1335 (N_1335,N_827,N_660);
or U1336 (N_1336,N_139,N_927);
or U1337 (N_1337,N_435,N_409);
or U1338 (N_1338,N_444,N_752);
nand U1339 (N_1339,N_391,N_665);
or U1340 (N_1340,N_612,N_969);
or U1341 (N_1341,N_744,N_957);
nand U1342 (N_1342,N_181,N_522);
nor U1343 (N_1343,N_833,N_230);
or U1344 (N_1344,N_161,N_908);
nand U1345 (N_1345,N_661,N_472);
and U1346 (N_1346,N_233,N_509);
or U1347 (N_1347,N_143,N_804);
or U1348 (N_1348,N_380,N_204);
nor U1349 (N_1349,N_218,N_737);
or U1350 (N_1350,N_507,N_595);
nor U1351 (N_1351,N_780,N_10);
xor U1352 (N_1352,N_130,N_471);
nor U1353 (N_1353,N_768,N_877);
xor U1354 (N_1354,N_351,N_155);
nor U1355 (N_1355,N_702,N_696);
and U1356 (N_1356,N_986,N_492);
xor U1357 (N_1357,N_197,N_97);
nor U1358 (N_1358,N_115,N_419);
and U1359 (N_1359,N_493,N_639);
or U1360 (N_1360,N_162,N_501);
nand U1361 (N_1361,N_430,N_959);
or U1362 (N_1362,N_449,N_714);
or U1363 (N_1363,N_541,N_274);
nand U1364 (N_1364,N_18,N_560);
nor U1365 (N_1365,N_76,N_864);
nand U1366 (N_1366,N_873,N_694);
or U1367 (N_1367,N_689,N_37);
and U1368 (N_1368,N_57,N_436);
or U1369 (N_1369,N_905,N_793);
nor U1370 (N_1370,N_785,N_41);
nand U1371 (N_1371,N_773,N_170);
or U1372 (N_1372,N_499,N_895);
and U1373 (N_1373,N_530,N_733);
nor U1374 (N_1374,N_571,N_374);
and U1375 (N_1375,N_730,N_817);
and U1376 (N_1376,N_465,N_692);
or U1377 (N_1377,N_642,N_26);
and U1378 (N_1378,N_284,N_585);
nand U1379 (N_1379,N_120,N_348);
and U1380 (N_1380,N_802,N_775);
xnor U1381 (N_1381,N_4,N_704);
nor U1382 (N_1382,N_407,N_281);
nor U1383 (N_1383,N_73,N_681);
or U1384 (N_1384,N_801,N_277);
or U1385 (N_1385,N_112,N_823);
nor U1386 (N_1386,N_171,N_926);
and U1387 (N_1387,N_356,N_456);
and U1388 (N_1388,N_79,N_973);
or U1389 (N_1389,N_474,N_31);
nand U1390 (N_1390,N_182,N_617);
nor U1391 (N_1391,N_792,N_17);
xor U1392 (N_1392,N_219,N_965);
and U1393 (N_1393,N_820,N_47);
or U1394 (N_1394,N_89,N_917);
and U1395 (N_1395,N_303,N_821);
and U1396 (N_1396,N_70,N_550);
nand U1397 (N_1397,N_662,N_77);
and U1398 (N_1398,N_350,N_320);
nand U1399 (N_1399,N_726,N_868);
nor U1400 (N_1400,N_800,N_527);
and U1401 (N_1401,N_482,N_434);
xnor U1402 (N_1402,N_708,N_193);
nand U1403 (N_1403,N_423,N_892);
and U1404 (N_1404,N_174,N_339);
and U1405 (N_1405,N_185,N_549);
and U1406 (N_1406,N_381,N_941);
or U1407 (N_1407,N_979,N_647);
and U1408 (N_1408,N_870,N_993);
or U1409 (N_1409,N_80,N_839);
nor U1410 (N_1410,N_526,N_620);
nand U1411 (N_1411,N_631,N_510);
and U1412 (N_1412,N_212,N_535);
nor U1413 (N_1413,N_265,N_294);
and U1414 (N_1414,N_691,N_515);
nor U1415 (N_1415,N_831,N_640);
nor U1416 (N_1416,N_911,N_916);
nor U1417 (N_1417,N_249,N_751);
nor U1418 (N_1418,N_34,N_124);
and U1419 (N_1419,N_999,N_512);
and U1420 (N_1420,N_937,N_314);
nor U1421 (N_1421,N_85,N_890);
and U1422 (N_1422,N_359,N_150);
xnor U1423 (N_1423,N_236,N_180);
xor U1424 (N_1424,N_789,N_898);
and U1425 (N_1425,N_35,N_835);
or U1426 (N_1426,N_411,N_42);
and U1427 (N_1427,N_458,N_59);
nor U1428 (N_1428,N_872,N_859);
nor U1429 (N_1429,N_238,N_279);
nand U1430 (N_1430,N_628,N_301);
or U1431 (N_1431,N_529,N_358);
nand U1432 (N_1432,N_745,N_875);
nand U1433 (N_1433,N_888,N_276);
and U1434 (N_1434,N_148,N_504);
nor U1435 (N_1435,N_133,N_567);
nand U1436 (N_1436,N_611,N_13);
nand U1437 (N_1437,N_220,N_950);
nor U1438 (N_1438,N_954,N_81);
and U1439 (N_1439,N_598,N_243);
nor U1440 (N_1440,N_253,N_226);
xnor U1441 (N_1441,N_297,N_206);
or U1442 (N_1442,N_313,N_653);
nand U1443 (N_1443,N_51,N_807);
nand U1444 (N_1444,N_210,N_199);
or U1445 (N_1445,N_624,N_542);
and U1446 (N_1446,N_673,N_537);
nand U1447 (N_1447,N_666,N_783);
and U1448 (N_1448,N_215,N_975);
nor U1449 (N_1449,N_721,N_777);
nor U1450 (N_1450,N_333,N_142);
and U1451 (N_1451,N_528,N_398);
nand U1452 (N_1452,N_160,N_534);
or U1453 (N_1453,N_988,N_543);
nand U1454 (N_1454,N_840,N_779);
or U1455 (N_1455,N_414,N_329);
xor U1456 (N_1456,N_989,N_710);
and U1457 (N_1457,N_834,N_224);
nor U1458 (N_1458,N_933,N_867);
nand U1459 (N_1459,N_566,N_153);
and U1460 (N_1460,N_27,N_487);
and U1461 (N_1461,N_63,N_280);
and U1462 (N_1462,N_588,N_250);
nor U1463 (N_1463,N_826,N_648);
or U1464 (N_1464,N_87,N_843);
or U1465 (N_1465,N_685,N_200);
nand U1466 (N_1466,N_383,N_86);
or U1467 (N_1467,N_599,N_40);
or U1468 (N_1468,N_879,N_422);
nand U1469 (N_1469,N_920,N_928);
or U1470 (N_1470,N_731,N_461);
and U1471 (N_1471,N_758,N_680);
nor U1472 (N_1472,N_626,N_54);
nor U1473 (N_1473,N_163,N_125);
or U1474 (N_1474,N_974,N_944);
xor U1475 (N_1475,N_658,N_184);
nor U1476 (N_1476,N_288,N_970);
nand U1477 (N_1477,N_844,N_925);
or U1478 (N_1478,N_229,N_587);
nand U1479 (N_1479,N_842,N_548);
or U1480 (N_1480,N_948,N_663);
nand U1481 (N_1481,N_403,N_881);
nor U1482 (N_1482,N_118,N_749);
and U1483 (N_1483,N_760,N_32);
nor U1484 (N_1484,N_791,N_887);
and U1485 (N_1485,N_52,N_402);
and U1486 (N_1486,N_813,N_234);
and U1487 (N_1487,N_392,N_201);
nor U1488 (N_1488,N_254,N_722);
and U1489 (N_1489,N_935,N_299);
and U1490 (N_1490,N_871,N_942);
or U1491 (N_1491,N_960,N_424);
and U1492 (N_1492,N_677,N_340);
and U1493 (N_1493,N_573,N_172);
nand U1494 (N_1494,N_816,N_217);
xor U1495 (N_1495,N_375,N_575);
nand U1496 (N_1496,N_99,N_452);
nand U1497 (N_1497,N_984,N_755);
nor U1498 (N_1498,N_565,N_48);
nor U1499 (N_1499,N_326,N_385);
or U1500 (N_1500,N_412,N_318);
or U1501 (N_1501,N_124,N_622);
nor U1502 (N_1502,N_610,N_228);
nor U1503 (N_1503,N_335,N_514);
and U1504 (N_1504,N_83,N_305);
xor U1505 (N_1505,N_276,N_194);
or U1506 (N_1506,N_954,N_241);
and U1507 (N_1507,N_24,N_325);
nor U1508 (N_1508,N_494,N_838);
nand U1509 (N_1509,N_286,N_284);
nand U1510 (N_1510,N_744,N_358);
or U1511 (N_1511,N_177,N_738);
nand U1512 (N_1512,N_794,N_780);
xnor U1513 (N_1513,N_277,N_142);
xor U1514 (N_1514,N_319,N_803);
and U1515 (N_1515,N_696,N_970);
and U1516 (N_1516,N_790,N_769);
or U1517 (N_1517,N_152,N_1);
or U1518 (N_1518,N_391,N_806);
or U1519 (N_1519,N_897,N_888);
nand U1520 (N_1520,N_353,N_476);
xnor U1521 (N_1521,N_438,N_526);
nand U1522 (N_1522,N_793,N_318);
and U1523 (N_1523,N_865,N_585);
nand U1524 (N_1524,N_994,N_484);
and U1525 (N_1525,N_353,N_129);
nand U1526 (N_1526,N_294,N_563);
nor U1527 (N_1527,N_866,N_28);
and U1528 (N_1528,N_149,N_132);
or U1529 (N_1529,N_675,N_285);
and U1530 (N_1530,N_198,N_606);
or U1531 (N_1531,N_805,N_598);
xnor U1532 (N_1532,N_810,N_940);
or U1533 (N_1533,N_29,N_733);
nor U1534 (N_1534,N_756,N_326);
nand U1535 (N_1535,N_300,N_506);
nor U1536 (N_1536,N_805,N_395);
and U1537 (N_1537,N_514,N_166);
and U1538 (N_1538,N_606,N_884);
and U1539 (N_1539,N_615,N_460);
or U1540 (N_1540,N_413,N_579);
and U1541 (N_1541,N_44,N_844);
xnor U1542 (N_1542,N_541,N_635);
or U1543 (N_1543,N_302,N_364);
and U1544 (N_1544,N_854,N_43);
or U1545 (N_1545,N_498,N_49);
and U1546 (N_1546,N_14,N_756);
or U1547 (N_1547,N_967,N_29);
or U1548 (N_1548,N_369,N_446);
nand U1549 (N_1549,N_280,N_724);
and U1550 (N_1550,N_337,N_930);
or U1551 (N_1551,N_936,N_542);
and U1552 (N_1552,N_100,N_660);
xor U1553 (N_1553,N_109,N_713);
or U1554 (N_1554,N_857,N_553);
nand U1555 (N_1555,N_1,N_63);
nor U1556 (N_1556,N_87,N_630);
or U1557 (N_1557,N_38,N_591);
or U1558 (N_1558,N_903,N_374);
nand U1559 (N_1559,N_375,N_251);
nor U1560 (N_1560,N_499,N_792);
and U1561 (N_1561,N_5,N_556);
nand U1562 (N_1562,N_749,N_706);
and U1563 (N_1563,N_858,N_343);
and U1564 (N_1564,N_609,N_846);
and U1565 (N_1565,N_734,N_139);
or U1566 (N_1566,N_124,N_612);
and U1567 (N_1567,N_193,N_587);
nand U1568 (N_1568,N_150,N_771);
or U1569 (N_1569,N_784,N_702);
nor U1570 (N_1570,N_661,N_538);
or U1571 (N_1571,N_164,N_341);
nor U1572 (N_1572,N_368,N_248);
or U1573 (N_1573,N_286,N_619);
or U1574 (N_1574,N_578,N_876);
nor U1575 (N_1575,N_693,N_947);
xnor U1576 (N_1576,N_529,N_194);
and U1577 (N_1577,N_816,N_505);
or U1578 (N_1578,N_675,N_303);
nor U1579 (N_1579,N_432,N_5);
nor U1580 (N_1580,N_765,N_441);
nand U1581 (N_1581,N_629,N_153);
and U1582 (N_1582,N_928,N_687);
nor U1583 (N_1583,N_186,N_932);
nand U1584 (N_1584,N_841,N_471);
and U1585 (N_1585,N_584,N_344);
nand U1586 (N_1586,N_819,N_423);
nand U1587 (N_1587,N_687,N_568);
or U1588 (N_1588,N_147,N_806);
xnor U1589 (N_1589,N_915,N_736);
and U1590 (N_1590,N_763,N_474);
and U1591 (N_1591,N_810,N_814);
nor U1592 (N_1592,N_621,N_859);
and U1593 (N_1593,N_648,N_39);
and U1594 (N_1594,N_453,N_3);
and U1595 (N_1595,N_811,N_906);
nand U1596 (N_1596,N_127,N_192);
nand U1597 (N_1597,N_947,N_725);
nor U1598 (N_1598,N_529,N_208);
or U1599 (N_1599,N_49,N_240);
and U1600 (N_1600,N_950,N_45);
nor U1601 (N_1601,N_424,N_932);
nand U1602 (N_1602,N_981,N_990);
nor U1603 (N_1603,N_207,N_627);
or U1604 (N_1604,N_52,N_193);
nor U1605 (N_1605,N_900,N_203);
or U1606 (N_1606,N_731,N_742);
and U1607 (N_1607,N_156,N_759);
and U1608 (N_1608,N_41,N_346);
or U1609 (N_1609,N_90,N_463);
or U1610 (N_1610,N_523,N_686);
xor U1611 (N_1611,N_608,N_409);
nor U1612 (N_1612,N_982,N_818);
and U1613 (N_1613,N_458,N_608);
or U1614 (N_1614,N_443,N_258);
nand U1615 (N_1615,N_991,N_952);
xnor U1616 (N_1616,N_852,N_524);
or U1617 (N_1617,N_723,N_126);
nor U1618 (N_1618,N_782,N_687);
nor U1619 (N_1619,N_360,N_211);
nand U1620 (N_1620,N_286,N_829);
nor U1621 (N_1621,N_318,N_419);
nand U1622 (N_1622,N_551,N_272);
or U1623 (N_1623,N_259,N_989);
xnor U1624 (N_1624,N_578,N_708);
nand U1625 (N_1625,N_30,N_143);
nor U1626 (N_1626,N_421,N_663);
and U1627 (N_1627,N_614,N_305);
nand U1628 (N_1628,N_819,N_882);
nor U1629 (N_1629,N_573,N_769);
and U1630 (N_1630,N_500,N_181);
and U1631 (N_1631,N_472,N_647);
nor U1632 (N_1632,N_298,N_916);
nor U1633 (N_1633,N_110,N_409);
or U1634 (N_1634,N_926,N_743);
or U1635 (N_1635,N_980,N_970);
xnor U1636 (N_1636,N_745,N_630);
xnor U1637 (N_1637,N_623,N_968);
nand U1638 (N_1638,N_502,N_643);
xor U1639 (N_1639,N_622,N_208);
or U1640 (N_1640,N_634,N_669);
or U1641 (N_1641,N_71,N_124);
nand U1642 (N_1642,N_745,N_163);
nor U1643 (N_1643,N_725,N_116);
nand U1644 (N_1644,N_500,N_12);
or U1645 (N_1645,N_619,N_599);
nand U1646 (N_1646,N_556,N_879);
nand U1647 (N_1647,N_298,N_100);
nand U1648 (N_1648,N_582,N_260);
or U1649 (N_1649,N_942,N_686);
xnor U1650 (N_1650,N_411,N_317);
and U1651 (N_1651,N_327,N_702);
or U1652 (N_1652,N_745,N_810);
xnor U1653 (N_1653,N_417,N_566);
nand U1654 (N_1654,N_343,N_602);
nand U1655 (N_1655,N_899,N_306);
xnor U1656 (N_1656,N_615,N_769);
or U1657 (N_1657,N_639,N_626);
xnor U1658 (N_1658,N_531,N_992);
nor U1659 (N_1659,N_882,N_195);
nand U1660 (N_1660,N_435,N_127);
or U1661 (N_1661,N_845,N_239);
nand U1662 (N_1662,N_306,N_552);
nand U1663 (N_1663,N_228,N_774);
xor U1664 (N_1664,N_910,N_475);
and U1665 (N_1665,N_741,N_516);
nor U1666 (N_1666,N_899,N_602);
nand U1667 (N_1667,N_588,N_213);
or U1668 (N_1668,N_437,N_339);
xnor U1669 (N_1669,N_676,N_66);
or U1670 (N_1670,N_265,N_54);
nand U1671 (N_1671,N_770,N_424);
or U1672 (N_1672,N_665,N_801);
or U1673 (N_1673,N_829,N_391);
or U1674 (N_1674,N_940,N_215);
nand U1675 (N_1675,N_126,N_165);
and U1676 (N_1676,N_62,N_572);
xor U1677 (N_1677,N_311,N_252);
nand U1678 (N_1678,N_120,N_652);
xnor U1679 (N_1679,N_223,N_673);
and U1680 (N_1680,N_776,N_965);
nor U1681 (N_1681,N_787,N_694);
and U1682 (N_1682,N_63,N_147);
and U1683 (N_1683,N_275,N_219);
and U1684 (N_1684,N_988,N_814);
and U1685 (N_1685,N_264,N_232);
nor U1686 (N_1686,N_833,N_941);
nand U1687 (N_1687,N_874,N_271);
nand U1688 (N_1688,N_39,N_629);
nor U1689 (N_1689,N_567,N_135);
nor U1690 (N_1690,N_825,N_170);
or U1691 (N_1691,N_730,N_407);
nand U1692 (N_1692,N_467,N_168);
and U1693 (N_1693,N_806,N_769);
nor U1694 (N_1694,N_509,N_442);
and U1695 (N_1695,N_198,N_16);
nand U1696 (N_1696,N_848,N_698);
or U1697 (N_1697,N_796,N_912);
or U1698 (N_1698,N_765,N_685);
nand U1699 (N_1699,N_719,N_295);
and U1700 (N_1700,N_459,N_719);
and U1701 (N_1701,N_438,N_187);
and U1702 (N_1702,N_859,N_191);
nand U1703 (N_1703,N_255,N_858);
or U1704 (N_1704,N_684,N_578);
nor U1705 (N_1705,N_136,N_772);
xnor U1706 (N_1706,N_161,N_654);
or U1707 (N_1707,N_160,N_34);
or U1708 (N_1708,N_321,N_130);
or U1709 (N_1709,N_950,N_962);
and U1710 (N_1710,N_572,N_413);
xor U1711 (N_1711,N_342,N_310);
or U1712 (N_1712,N_496,N_786);
nor U1713 (N_1713,N_42,N_918);
nand U1714 (N_1714,N_543,N_956);
or U1715 (N_1715,N_301,N_992);
nand U1716 (N_1716,N_109,N_617);
and U1717 (N_1717,N_112,N_248);
xor U1718 (N_1718,N_781,N_533);
and U1719 (N_1719,N_419,N_413);
and U1720 (N_1720,N_858,N_386);
or U1721 (N_1721,N_312,N_593);
nand U1722 (N_1722,N_97,N_284);
and U1723 (N_1723,N_539,N_105);
xor U1724 (N_1724,N_742,N_270);
or U1725 (N_1725,N_184,N_818);
and U1726 (N_1726,N_241,N_835);
and U1727 (N_1727,N_910,N_347);
and U1728 (N_1728,N_302,N_859);
and U1729 (N_1729,N_52,N_314);
nor U1730 (N_1730,N_287,N_144);
and U1731 (N_1731,N_402,N_939);
nand U1732 (N_1732,N_876,N_467);
or U1733 (N_1733,N_883,N_213);
nand U1734 (N_1734,N_176,N_486);
xor U1735 (N_1735,N_131,N_766);
nand U1736 (N_1736,N_961,N_492);
or U1737 (N_1737,N_676,N_853);
xnor U1738 (N_1738,N_890,N_926);
xnor U1739 (N_1739,N_774,N_962);
or U1740 (N_1740,N_345,N_736);
nor U1741 (N_1741,N_473,N_711);
nor U1742 (N_1742,N_505,N_893);
and U1743 (N_1743,N_555,N_185);
nand U1744 (N_1744,N_673,N_915);
or U1745 (N_1745,N_924,N_82);
and U1746 (N_1746,N_982,N_749);
nor U1747 (N_1747,N_28,N_228);
nand U1748 (N_1748,N_210,N_784);
xor U1749 (N_1749,N_66,N_980);
and U1750 (N_1750,N_390,N_454);
and U1751 (N_1751,N_453,N_38);
xnor U1752 (N_1752,N_416,N_916);
or U1753 (N_1753,N_301,N_897);
nor U1754 (N_1754,N_654,N_576);
nand U1755 (N_1755,N_789,N_833);
nor U1756 (N_1756,N_879,N_959);
nor U1757 (N_1757,N_265,N_272);
or U1758 (N_1758,N_84,N_542);
xnor U1759 (N_1759,N_230,N_246);
or U1760 (N_1760,N_984,N_534);
or U1761 (N_1761,N_734,N_946);
xnor U1762 (N_1762,N_71,N_252);
and U1763 (N_1763,N_685,N_117);
and U1764 (N_1764,N_962,N_500);
xnor U1765 (N_1765,N_697,N_404);
nand U1766 (N_1766,N_379,N_632);
or U1767 (N_1767,N_829,N_349);
and U1768 (N_1768,N_472,N_562);
or U1769 (N_1769,N_263,N_730);
nor U1770 (N_1770,N_846,N_855);
and U1771 (N_1771,N_696,N_321);
nor U1772 (N_1772,N_545,N_199);
xnor U1773 (N_1773,N_449,N_484);
nand U1774 (N_1774,N_338,N_358);
nand U1775 (N_1775,N_146,N_436);
or U1776 (N_1776,N_71,N_739);
xor U1777 (N_1777,N_384,N_323);
nor U1778 (N_1778,N_133,N_944);
xnor U1779 (N_1779,N_805,N_708);
nand U1780 (N_1780,N_206,N_87);
nand U1781 (N_1781,N_445,N_457);
or U1782 (N_1782,N_999,N_983);
and U1783 (N_1783,N_5,N_207);
nor U1784 (N_1784,N_426,N_265);
xnor U1785 (N_1785,N_135,N_210);
nor U1786 (N_1786,N_724,N_860);
and U1787 (N_1787,N_178,N_635);
or U1788 (N_1788,N_523,N_629);
nand U1789 (N_1789,N_521,N_267);
or U1790 (N_1790,N_201,N_330);
or U1791 (N_1791,N_71,N_581);
nor U1792 (N_1792,N_216,N_462);
nand U1793 (N_1793,N_424,N_912);
or U1794 (N_1794,N_486,N_672);
and U1795 (N_1795,N_407,N_536);
or U1796 (N_1796,N_223,N_860);
nand U1797 (N_1797,N_49,N_379);
and U1798 (N_1798,N_445,N_996);
nand U1799 (N_1799,N_825,N_867);
or U1800 (N_1800,N_288,N_195);
nand U1801 (N_1801,N_732,N_498);
or U1802 (N_1802,N_948,N_385);
nor U1803 (N_1803,N_367,N_705);
nand U1804 (N_1804,N_123,N_430);
or U1805 (N_1805,N_681,N_379);
or U1806 (N_1806,N_265,N_722);
xnor U1807 (N_1807,N_564,N_604);
nand U1808 (N_1808,N_79,N_98);
nand U1809 (N_1809,N_798,N_756);
nand U1810 (N_1810,N_473,N_914);
nand U1811 (N_1811,N_326,N_40);
and U1812 (N_1812,N_847,N_365);
nor U1813 (N_1813,N_334,N_214);
and U1814 (N_1814,N_426,N_791);
or U1815 (N_1815,N_337,N_437);
nand U1816 (N_1816,N_774,N_394);
nor U1817 (N_1817,N_565,N_765);
and U1818 (N_1818,N_271,N_326);
or U1819 (N_1819,N_287,N_40);
or U1820 (N_1820,N_925,N_40);
nand U1821 (N_1821,N_205,N_230);
nand U1822 (N_1822,N_801,N_966);
and U1823 (N_1823,N_131,N_449);
nand U1824 (N_1824,N_819,N_951);
or U1825 (N_1825,N_226,N_116);
or U1826 (N_1826,N_120,N_491);
or U1827 (N_1827,N_848,N_64);
or U1828 (N_1828,N_352,N_107);
and U1829 (N_1829,N_261,N_843);
nor U1830 (N_1830,N_578,N_799);
or U1831 (N_1831,N_167,N_265);
nand U1832 (N_1832,N_750,N_688);
nor U1833 (N_1833,N_815,N_211);
nor U1834 (N_1834,N_375,N_56);
nand U1835 (N_1835,N_589,N_825);
nor U1836 (N_1836,N_974,N_987);
or U1837 (N_1837,N_745,N_24);
or U1838 (N_1838,N_317,N_895);
and U1839 (N_1839,N_52,N_115);
and U1840 (N_1840,N_674,N_41);
nor U1841 (N_1841,N_770,N_402);
nor U1842 (N_1842,N_879,N_159);
nand U1843 (N_1843,N_414,N_217);
and U1844 (N_1844,N_112,N_703);
xor U1845 (N_1845,N_450,N_877);
or U1846 (N_1846,N_920,N_369);
nor U1847 (N_1847,N_959,N_461);
and U1848 (N_1848,N_94,N_540);
xor U1849 (N_1849,N_17,N_332);
nor U1850 (N_1850,N_802,N_623);
xor U1851 (N_1851,N_233,N_690);
and U1852 (N_1852,N_257,N_998);
nor U1853 (N_1853,N_672,N_348);
and U1854 (N_1854,N_491,N_745);
and U1855 (N_1855,N_466,N_263);
nor U1856 (N_1856,N_483,N_650);
nand U1857 (N_1857,N_809,N_871);
nand U1858 (N_1858,N_635,N_865);
nor U1859 (N_1859,N_287,N_428);
nand U1860 (N_1860,N_83,N_391);
nor U1861 (N_1861,N_663,N_968);
nand U1862 (N_1862,N_794,N_914);
and U1863 (N_1863,N_442,N_828);
nor U1864 (N_1864,N_246,N_612);
nand U1865 (N_1865,N_144,N_112);
nand U1866 (N_1866,N_266,N_675);
nor U1867 (N_1867,N_388,N_225);
nand U1868 (N_1868,N_462,N_42);
and U1869 (N_1869,N_176,N_180);
xnor U1870 (N_1870,N_432,N_636);
nor U1871 (N_1871,N_137,N_547);
or U1872 (N_1872,N_406,N_462);
nor U1873 (N_1873,N_123,N_10);
or U1874 (N_1874,N_763,N_532);
nand U1875 (N_1875,N_336,N_639);
nand U1876 (N_1876,N_701,N_315);
or U1877 (N_1877,N_895,N_362);
and U1878 (N_1878,N_665,N_664);
nor U1879 (N_1879,N_636,N_495);
nand U1880 (N_1880,N_379,N_982);
nor U1881 (N_1881,N_737,N_298);
nor U1882 (N_1882,N_696,N_522);
and U1883 (N_1883,N_701,N_153);
or U1884 (N_1884,N_100,N_199);
nor U1885 (N_1885,N_71,N_100);
nor U1886 (N_1886,N_278,N_381);
and U1887 (N_1887,N_417,N_950);
and U1888 (N_1888,N_527,N_39);
nor U1889 (N_1889,N_228,N_822);
or U1890 (N_1890,N_310,N_863);
nand U1891 (N_1891,N_236,N_32);
and U1892 (N_1892,N_125,N_824);
nor U1893 (N_1893,N_56,N_286);
nand U1894 (N_1894,N_167,N_229);
nand U1895 (N_1895,N_403,N_664);
or U1896 (N_1896,N_474,N_30);
nor U1897 (N_1897,N_679,N_700);
nor U1898 (N_1898,N_284,N_13);
or U1899 (N_1899,N_543,N_855);
or U1900 (N_1900,N_146,N_130);
nand U1901 (N_1901,N_549,N_99);
nor U1902 (N_1902,N_504,N_913);
nor U1903 (N_1903,N_7,N_853);
nand U1904 (N_1904,N_743,N_854);
nor U1905 (N_1905,N_570,N_862);
nand U1906 (N_1906,N_947,N_79);
or U1907 (N_1907,N_621,N_891);
nor U1908 (N_1908,N_27,N_472);
nor U1909 (N_1909,N_616,N_144);
or U1910 (N_1910,N_540,N_302);
and U1911 (N_1911,N_118,N_34);
nor U1912 (N_1912,N_970,N_899);
and U1913 (N_1913,N_341,N_26);
or U1914 (N_1914,N_909,N_31);
nor U1915 (N_1915,N_416,N_265);
and U1916 (N_1916,N_813,N_591);
nor U1917 (N_1917,N_406,N_435);
and U1918 (N_1918,N_568,N_90);
xnor U1919 (N_1919,N_476,N_500);
nand U1920 (N_1920,N_147,N_25);
xnor U1921 (N_1921,N_471,N_968);
and U1922 (N_1922,N_411,N_712);
nor U1923 (N_1923,N_901,N_867);
nor U1924 (N_1924,N_151,N_223);
nor U1925 (N_1925,N_171,N_612);
nand U1926 (N_1926,N_537,N_17);
nand U1927 (N_1927,N_130,N_117);
and U1928 (N_1928,N_695,N_891);
nand U1929 (N_1929,N_452,N_629);
nand U1930 (N_1930,N_54,N_215);
nor U1931 (N_1931,N_16,N_424);
nand U1932 (N_1932,N_276,N_474);
or U1933 (N_1933,N_984,N_966);
or U1934 (N_1934,N_493,N_970);
nor U1935 (N_1935,N_510,N_11);
nand U1936 (N_1936,N_376,N_540);
nor U1937 (N_1937,N_802,N_929);
nand U1938 (N_1938,N_294,N_806);
or U1939 (N_1939,N_490,N_391);
nor U1940 (N_1940,N_574,N_661);
xor U1941 (N_1941,N_71,N_341);
or U1942 (N_1942,N_775,N_936);
and U1943 (N_1943,N_351,N_204);
nand U1944 (N_1944,N_604,N_0);
or U1945 (N_1945,N_116,N_404);
xor U1946 (N_1946,N_967,N_879);
and U1947 (N_1947,N_937,N_716);
and U1948 (N_1948,N_110,N_825);
and U1949 (N_1949,N_788,N_70);
or U1950 (N_1950,N_583,N_145);
nor U1951 (N_1951,N_588,N_320);
or U1952 (N_1952,N_762,N_942);
nand U1953 (N_1953,N_363,N_634);
or U1954 (N_1954,N_298,N_946);
nor U1955 (N_1955,N_535,N_977);
and U1956 (N_1956,N_635,N_944);
nor U1957 (N_1957,N_11,N_701);
and U1958 (N_1958,N_805,N_10);
and U1959 (N_1959,N_48,N_905);
nand U1960 (N_1960,N_275,N_478);
nor U1961 (N_1961,N_214,N_862);
or U1962 (N_1962,N_77,N_718);
and U1963 (N_1963,N_338,N_306);
and U1964 (N_1964,N_437,N_371);
and U1965 (N_1965,N_838,N_19);
or U1966 (N_1966,N_344,N_781);
nand U1967 (N_1967,N_696,N_801);
nand U1968 (N_1968,N_113,N_43);
and U1969 (N_1969,N_731,N_956);
xnor U1970 (N_1970,N_945,N_362);
and U1971 (N_1971,N_74,N_352);
nand U1972 (N_1972,N_39,N_845);
xor U1973 (N_1973,N_825,N_81);
nand U1974 (N_1974,N_980,N_189);
or U1975 (N_1975,N_895,N_607);
nand U1976 (N_1976,N_681,N_61);
nor U1977 (N_1977,N_557,N_117);
and U1978 (N_1978,N_227,N_772);
or U1979 (N_1979,N_635,N_81);
nand U1980 (N_1980,N_407,N_859);
nand U1981 (N_1981,N_238,N_18);
or U1982 (N_1982,N_215,N_317);
nand U1983 (N_1983,N_86,N_321);
and U1984 (N_1984,N_615,N_86);
nor U1985 (N_1985,N_60,N_943);
nand U1986 (N_1986,N_563,N_913);
nor U1987 (N_1987,N_550,N_985);
and U1988 (N_1988,N_653,N_611);
nor U1989 (N_1989,N_249,N_113);
and U1990 (N_1990,N_957,N_175);
nor U1991 (N_1991,N_75,N_226);
nand U1992 (N_1992,N_356,N_887);
nor U1993 (N_1993,N_18,N_161);
nand U1994 (N_1994,N_858,N_253);
xor U1995 (N_1995,N_986,N_517);
nor U1996 (N_1996,N_307,N_937);
nor U1997 (N_1997,N_321,N_521);
nor U1998 (N_1998,N_189,N_962);
xor U1999 (N_1999,N_85,N_139);
xor U2000 (N_2000,N_1119,N_1170);
nand U2001 (N_2001,N_1889,N_1174);
or U2002 (N_2002,N_1704,N_1568);
and U2003 (N_2003,N_1812,N_1600);
or U2004 (N_2004,N_1724,N_1909);
nand U2005 (N_2005,N_1826,N_1437);
or U2006 (N_2006,N_1795,N_1647);
nand U2007 (N_2007,N_1792,N_1341);
nor U2008 (N_2008,N_1538,N_1066);
and U2009 (N_2009,N_1523,N_1630);
xor U2010 (N_2010,N_1971,N_1895);
and U2011 (N_2011,N_1569,N_1782);
nor U2012 (N_2012,N_1198,N_1722);
and U2013 (N_2013,N_1653,N_1186);
nand U2014 (N_2014,N_1698,N_1089);
nand U2015 (N_2015,N_1034,N_1990);
and U2016 (N_2016,N_1804,N_1528);
and U2017 (N_2017,N_1395,N_1199);
nor U2018 (N_2018,N_1354,N_1861);
nand U2019 (N_2019,N_1469,N_1539);
and U2020 (N_2020,N_1373,N_1043);
nand U2021 (N_2021,N_1381,N_1711);
or U2022 (N_2022,N_1945,N_1326);
nand U2023 (N_2023,N_1693,N_1480);
or U2024 (N_2024,N_1218,N_1321);
nor U2025 (N_2025,N_1825,N_1735);
nand U2026 (N_2026,N_1271,N_1232);
nand U2027 (N_2027,N_1108,N_1473);
or U2028 (N_2028,N_1947,N_1422);
nand U2029 (N_2029,N_1509,N_1963);
and U2030 (N_2030,N_1930,N_1579);
nand U2031 (N_2031,N_1876,N_1486);
nor U2032 (N_2032,N_1823,N_1520);
nor U2033 (N_2033,N_1334,N_1896);
nand U2034 (N_2034,N_1856,N_1346);
nand U2035 (N_2035,N_1261,N_1496);
nor U2036 (N_2036,N_1684,N_1942);
nand U2037 (N_2037,N_1970,N_1940);
nor U2038 (N_2038,N_1993,N_1254);
and U2039 (N_2039,N_1512,N_1585);
and U2040 (N_2040,N_1831,N_1086);
nand U2041 (N_2041,N_1873,N_1529);
or U2042 (N_2042,N_1537,N_1582);
nand U2043 (N_2043,N_1293,N_1927);
nor U2044 (N_2044,N_1713,N_1629);
nand U2045 (N_2045,N_1239,N_1706);
nand U2046 (N_2046,N_1998,N_1263);
nand U2047 (N_2047,N_1828,N_1885);
and U2048 (N_2048,N_1367,N_1617);
and U2049 (N_2049,N_1421,N_1734);
and U2050 (N_2050,N_1608,N_1903);
nand U2051 (N_2051,N_1181,N_1841);
or U2052 (N_2052,N_1316,N_1266);
nand U2053 (N_2053,N_1039,N_1370);
or U2054 (N_2054,N_1598,N_1914);
nor U2055 (N_2055,N_1465,N_1808);
nand U2056 (N_2056,N_1526,N_1589);
nand U2057 (N_2057,N_1456,N_1967);
or U2058 (N_2058,N_1965,N_1671);
xor U2059 (N_2059,N_1069,N_1228);
and U2060 (N_2060,N_1223,N_1285);
nand U2061 (N_2061,N_1615,N_1681);
and U2062 (N_2062,N_1661,N_1888);
or U2063 (N_2063,N_1461,N_1987);
or U2064 (N_2064,N_1624,N_1287);
nor U2065 (N_2065,N_1148,N_1769);
xnor U2066 (N_2066,N_1616,N_1028);
nand U2067 (N_2067,N_1201,N_1476);
and U2068 (N_2068,N_1121,N_1962);
nand U2069 (N_2069,N_1430,N_1580);
and U2070 (N_2070,N_1319,N_1205);
nor U2071 (N_2071,N_1351,N_1923);
and U2072 (N_2072,N_1144,N_1216);
nand U2073 (N_2073,N_1590,N_1871);
or U2074 (N_2074,N_1510,N_1785);
nand U2075 (N_2075,N_1749,N_1938);
and U2076 (N_2076,N_1961,N_1152);
and U2077 (N_2077,N_1125,N_1561);
and U2078 (N_2078,N_1442,N_1296);
or U2079 (N_2079,N_1423,N_1892);
nand U2080 (N_2080,N_1002,N_1359);
xor U2081 (N_2081,N_1564,N_1439);
and U2082 (N_2082,N_1837,N_1050);
nor U2083 (N_2083,N_1950,N_1699);
nand U2084 (N_2084,N_1434,N_1409);
nand U2085 (N_2085,N_1744,N_1061);
nand U2086 (N_2086,N_1406,N_1168);
or U2087 (N_2087,N_1774,N_1867);
nand U2088 (N_2088,N_1605,N_1779);
nand U2089 (N_2089,N_1384,N_1010);
nor U2090 (N_2090,N_1918,N_1401);
or U2091 (N_2091,N_1672,N_1543);
nor U2092 (N_2092,N_1103,N_1030);
nand U2093 (N_2093,N_1195,N_1435);
nor U2094 (N_2094,N_1275,N_1265);
nand U2095 (N_2095,N_1488,N_1768);
nand U2096 (N_2096,N_1448,N_1431);
or U2097 (N_2097,N_1462,N_1182);
or U2098 (N_2098,N_1820,N_1881);
nand U2099 (N_2099,N_1207,N_1491);
nor U2100 (N_2100,N_1008,N_1660);
and U2101 (N_2101,N_1169,N_1798);
xnor U2102 (N_2102,N_1709,N_1677);
or U2103 (N_2103,N_1802,N_1413);
and U2104 (N_2104,N_1594,N_1806);
nor U2105 (N_2105,N_1504,N_1872);
nand U2106 (N_2106,N_1011,N_1137);
nor U2107 (N_2107,N_1732,N_1308);
and U2108 (N_2108,N_1811,N_1708);
or U2109 (N_2109,N_1131,N_1953);
or U2110 (N_2110,N_1757,N_1386);
nor U2111 (N_2111,N_1356,N_1247);
nor U2112 (N_2112,N_1358,N_1130);
and U2113 (N_2113,N_1071,N_1333);
xnor U2114 (N_2114,N_1816,N_1101);
nor U2115 (N_2115,N_1482,N_1076);
and U2116 (N_2116,N_1584,N_1485);
xor U2117 (N_2117,N_1767,N_1555);
nand U2118 (N_2118,N_1911,N_1475);
xnor U2119 (N_2119,N_1338,N_1560);
nand U2120 (N_2120,N_1666,N_1443);
or U2121 (N_2121,N_1094,N_1638);
nor U2122 (N_2122,N_1748,N_1851);
nand U2123 (N_2123,N_1946,N_1105);
nand U2124 (N_2124,N_1695,N_1570);
nor U2125 (N_2125,N_1747,N_1236);
and U2126 (N_2126,N_1284,N_1890);
or U2127 (N_2127,N_1606,N_1801);
nand U2128 (N_2128,N_1141,N_1315);
or U2129 (N_2129,N_1793,N_1112);
or U2130 (N_2130,N_1226,N_1328);
and U2131 (N_2131,N_1139,N_1353);
xnor U2132 (N_2132,N_1268,N_1074);
or U2133 (N_2133,N_1032,N_1360);
and U2134 (N_2134,N_1493,N_1024);
nand U2135 (N_2135,N_1751,N_1175);
nand U2136 (N_2136,N_1759,N_1276);
nor U2137 (N_2137,N_1490,N_1879);
and U2138 (N_2138,N_1348,N_1920);
nor U2139 (N_2139,N_1634,N_1545);
and U2140 (N_2140,N_1730,N_1781);
and U2141 (N_2141,N_1057,N_1291);
nor U2142 (N_2142,N_1257,N_1116);
or U2143 (N_2143,N_1780,N_1639);
nor U2144 (N_2144,N_1642,N_1952);
nand U2145 (N_2145,N_1815,N_1127);
nor U2146 (N_2146,N_1149,N_1068);
xnor U2147 (N_2147,N_1988,N_1158);
nor U2148 (N_2148,N_1040,N_1824);
nor U2149 (N_2149,N_1622,N_1736);
or U2150 (N_2150,N_1863,N_1729);
or U2151 (N_2151,N_1391,N_1805);
and U2152 (N_2152,N_1613,N_1562);
and U2153 (N_2153,N_1797,N_1796);
nor U2154 (N_2154,N_1541,N_1789);
xor U2155 (N_2155,N_1368,N_1702);
or U2156 (N_2156,N_1436,N_1095);
nor U2157 (N_2157,N_1106,N_1450);
nand U2158 (N_2158,N_1227,N_1311);
and U2159 (N_2159,N_1627,N_1016);
or U2160 (N_2160,N_1870,N_1459);
nor U2161 (N_2161,N_1472,N_1836);
nand U2162 (N_2162,N_1534,N_1689);
or U2163 (N_2163,N_1314,N_1573);
nand U2164 (N_2164,N_1760,N_1013);
and U2165 (N_2165,N_1077,N_1173);
or U2166 (N_2166,N_1648,N_1344);
nand U2167 (N_2167,N_1256,N_1164);
nand U2168 (N_2168,N_1567,N_1775);
and U2169 (N_2169,N_1157,N_1756);
nor U2170 (N_2170,N_1309,N_1745);
and U2171 (N_2171,N_1269,N_1283);
nand U2172 (N_2172,N_1458,N_1065);
nand U2173 (N_2173,N_1934,N_1324);
and U2174 (N_2174,N_1166,N_1766);
nand U2175 (N_2175,N_1716,N_1571);
xnor U2176 (N_2176,N_1984,N_1156);
nor U2177 (N_2177,N_1038,N_1958);
nand U2178 (N_2178,N_1982,N_1093);
nand U2179 (N_2179,N_1104,N_1398);
nor U2180 (N_2180,N_1933,N_1669);
nand U2181 (N_2181,N_1471,N_1320);
nor U2182 (N_2182,N_1126,N_1411);
nand U2183 (N_2183,N_1073,N_1884);
xor U2184 (N_2184,N_1463,N_1814);
and U2185 (N_2185,N_1492,N_1047);
or U2186 (N_2186,N_1712,N_1803);
and U2187 (N_2187,N_1058,N_1162);
nor U2188 (N_2188,N_1402,N_1551);
or U2189 (N_2189,N_1649,N_1901);
or U2190 (N_2190,N_1455,N_1318);
and U2191 (N_2191,N_1847,N_1021);
xnor U2192 (N_2192,N_1978,N_1741);
nand U2193 (N_2193,N_1053,N_1260);
or U2194 (N_2194,N_1536,N_1300);
or U2195 (N_2195,N_1457,N_1165);
or U2196 (N_2196,N_1596,N_1403);
and U2197 (N_2197,N_1621,N_1111);
nor U2198 (N_2198,N_1989,N_1379);
and U2199 (N_2199,N_1549,N_1091);
or U2200 (N_2200,N_1396,N_1694);
and U2201 (N_2201,N_1894,N_1481);
nand U2202 (N_2202,N_1214,N_1146);
or U2203 (N_2203,N_1500,N_1022);
nand U2204 (N_2204,N_1676,N_1874);
and U2205 (N_2205,N_1683,N_1846);
or U2206 (N_2206,N_1385,N_1686);
or U2207 (N_2207,N_1117,N_1720);
and U2208 (N_2208,N_1150,N_1184);
nor U2209 (N_2209,N_1502,N_1827);
and U2210 (N_2210,N_1290,N_1371);
nand U2211 (N_2211,N_1453,N_1682);
nand U2212 (N_2212,N_1864,N_1794);
nand U2213 (N_2213,N_1147,N_1176);
nor U2214 (N_2214,N_1540,N_1429);
and U2215 (N_2215,N_1067,N_1675);
and U2216 (N_2216,N_1707,N_1160);
nand U2217 (N_2217,N_1244,N_1483);
and U2218 (N_2218,N_1817,N_1288);
nor U2219 (N_2219,N_1503,N_1614);
nor U2220 (N_2220,N_1020,N_1979);
and U2221 (N_2221,N_1737,N_1419);
nor U2222 (N_2222,N_1041,N_1096);
or U2223 (N_2223,N_1964,N_1136);
nor U2224 (N_2224,N_1188,N_1511);
nand U2225 (N_2225,N_1151,N_1045);
xnor U2226 (N_2226,N_1926,N_1948);
nand U2227 (N_2227,N_1187,N_1240);
nor U2228 (N_2228,N_1866,N_1656);
and U2229 (N_2229,N_1612,N_1939);
nand U2230 (N_2230,N_1644,N_1432);
nand U2231 (N_2231,N_1897,N_1611);
or U2232 (N_2232,N_1618,N_1468);
nand U2233 (N_2233,N_1765,N_1088);
nand U2234 (N_2234,N_1143,N_1394);
or U2235 (N_2235,N_1878,N_1597);
or U2236 (N_2236,N_1212,N_1025);
nor U2237 (N_2237,N_1393,N_1410);
nand U2238 (N_2238,N_1714,N_1109);
and U2239 (N_2239,N_1085,N_1548);
or U2240 (N_2240,N_1110,N_1916);
nor U2241 (N_2241,N_1754,N_1996);
nor U2242 (N_2242,N_1124,N_1771);
or U2243 (N_2243,N_1688,N_1154);
and U2244 (N_2244,N_1849,N_1908);
and U2245 (N_2245,N_1977,N_1850);
or U2246 (N_2246,N_1286,N_1222);
and U2247 (N_2247,N_1924,N_1762);
nand U2248 (N_2248,N_1397,N_1533);
nand U2249 (N_2249,N_1635,N_1886);
nand U2250 (N_2250,N_1913,N_1563);
nor U2251 (N_2251,N_1052,N_1327);
xnor U2252 (N_2252,N_1070,N_1578);
nor U2253 (N_2253,N_1378,N_1636);
or U2254 (N_2254,N_1830,N_1262);
or U2255 (N_2255,N_1023,N_1026);
or U2256 (N_2256,N_1784,N_1667);
nand U2257 (N_2257,N_1248,N_1113);
nand U2258 (N_2258,N_1005,N_1506);
nor U2259 (N_2259,N_1377,N_1976);
xnor U2260 (N_2260,N_1650,N_1389);
nand U2261 (N_2261,N_1731,N_1936);
nor U2262 (N_2262,N_1525,N_1799);
nand U2263 (N_2263,N_1625,N_1860);
or U2264 (N_2264,N_1554,N_1438);
nand U2265 (N_2265,N_1786,N_1044);
and U2266 (N_2266,N_1031,N_1210);
xnor U2267 (N_2267,N_1003,N_1331);
and U2268 (N_2268,N_1915,N_1547);
xnor U2269 (N_2269,N_1834,N_1738);
nor U2270 (N_2270,N_1508,N_1906);
or U2271 (N_2271,N_1992,N_1444);
nor U2272 (N_2272,N_1000,N_1209);
xor U2273 (N_2273,N_1420,N_1832);
nor U2274 (N_2274,N_1274,N_1535);
and U2275 (N_2275,N_1898,N_1242);
nand U2276 (N_2276,N_1279,N_1733);
or U2277 (N_2277,N_1033,N_1783);
or U2278 (N_2278,N_1362,N_1728);
or U2279 (N_2279,N_1544,N_1907);
xnor U2280 (N_2280,N_1084,N_1855);
or U2281 (N_2281,N_1788,N_1479);
and U2282 (N_2282,N_1342,N_1776);
and U2283 (N_2283,N_1626,N_1441);
or U2284 (N_2284,N_1721,N_1822);
nor U2285 (N_2285,N_1739,N_1138);
nand U2286 (N_2286,N_1224,N_1282);
or U2287 (N_2287,N_1376,N_1631);
nand U2288 (N_2288,N_1001,N_1668);
and U2289 (N_2289,N_1542,N_1763);
or U2290 (N_2290,N_1078,N_1514);
and U2291 (N_2291,N_1054,N_1657);
and U2292 (N_2292,N_1347,N_1951);
or U2293 (N_2293,N_1400,N_1446);
nand U2294 (N_2294,N_1957,N_1703);
and U2295 (N_2295,N_1552,N_1937);
or U2296 (N_2296,N_1383,N_1531);
nand U2297 (N_2297,N_1887,N_1451);
and U2298 (N_2298,N_1727,N_1405);
nand U2299 (N_2299,N_1659,N_1229);
or U2300 (N_2300,N_1035,N_1679);
nand U2301 (N_2301,N_1225,N_1064);
or U2302 (N_2302,N_1129,N_1691);
and U2303 (N_2303,N_1726,N_1601);
or U2304 (N_2304,N_1845,N_1407);
or U2305 (N_2305,N_1252,N_1417);
and U2306 (N_2306,N_1325,N_1098);
nor U2307 (N_2307,N_1857,N_1858);
or U2308 (N_2308,N_1470,N_1235);
or U2309 (N_2309,N_1883,N_1997);
nor U2310 (N_2310,N_1440,N_1029);
nor U2311 (N_2311,N_1390,N_1991);
nand U2312 (N_2312,N_1498,N_1464);
and U2313 (N_2313,N_1973,N_1840);
nand U2314 (N_2314,N_1452,N_1079);
and U2315 (N_2315,N_1340,N_1087);
or U2316 (N_2316,N_1234,N_1194);
or U2317 (N_2317,N_1289,N_1807);
or U2318 (N_2318,N_1004,N_1221);
or U2319 (N_2319,N_1418,N_1048);
or U2320 (N_2320,N_1416,N_1424);
nand U2321 (N_2321,N_1270,N_1576);
and U2322 (N_2322,N_1049,N_1685);
nand U2323 (N_2323,N_1852,N_1297);
nor U2324 (N_2324,N_1055,N_1322);
or U2325 (N_2325,N_1574,N_1355);
xor U2326 (N_2326,N_1009,N_1556);
or U2327 (N_2327,N_1056,N_1519);
nand U2328 (N_2328,N_1843,N_1761);
xnor U2329 (N_2329,N_1128,N_1272);
xor U2330 (N_2330,N_1838,N_1445);
and U2331 (N_2331,N_1875,N_1298);
nor U2332 (N_2332,N_1123,N_1818);
or U2333 (N_2333,N_1652,N_1306);
nor U2334 (N_2334,N_1932,N_1929);
nand U2335 (N_2335,N_1692,N_1809);
nand U2336 (N_2336,N_1524,N_1607);
nand U2337 (N_2337,N_1253,N_1246);
nor U2338 (N_2338,N_1980,N_1835);
nor U2339 (N_2339,N_1477,N_1259);
and U2340 (N_2340,N_1292,N_1277);
or U2341 (N_2341,N_1191,N_1099);
nand U2342 (N_2342,N_1425,N_1211);
or U2343 (N_2343,N_1036,N_1238);
xor U2344 (N_2344,N_1891,N_1610);
xnor U2345 (N_2345,N_1755,N_1854);
nand U2346 (N_2346,N_1842,N_1100);
or U2347 (N_2347,N_1335,N_1859);
nor U2348 (N_2348,N_1821,N_1140);
nor U2349 (N_2349,N_1294,N_1900);
nor U2350 (N_2350,N_1161,N_1975);
xor U2351 (N_2351,N_1499,N_1081);
xnor U2352 (N_2352,N_1696,N_1332);
nor U2353 (N_2353,N_1281,N_1723);
nand U2354 (N_2354,N_1591,N_1955);
nand U2355 (N_2355,N_1880,N_1893);
xor U2356 (N_2356,N_1905,N_1641);
xor U2357 (N_2357,N_1018,N_1633);
or U2358 (N_2358,N_1848,N_1717);
and U2359 (N_2359,N_1213,N_1267);
or U2360 (N_2360,N_1925,N_1742);
and U2361 (N_2361,N_1200,N_1778);
xnor U2362 (N_2362,N_1619,N_1178);
nor U2363 (N_2363,N_1142,N_1701);
or U2364 (N_2364,N_1329,N_1609);
and U2365 (N_2365,N_1972,N_1674);
nor U2366 (N_2366,N_1323,N_1575);
nand U2367 (N_2367,N_1273,N_1586);
or U2368 (N_2368,N_1364,N_1303);
nand U2369 (N_2369,N_1643,N_1250);
and U2370 (N_2370,N_1145,N_1999);
and U2371 (N_2371,N_1985,N_1190);
nand U2372 (N_2372,N_1375,N_1966);
and U2373 (N_2373,N_1447,N_1902);
and U2374 (N_2374,N_1899,N_1532);
or U2375 (N_2375,N_1467,N_1427);
and U2376 (N_2376,N_1877,N_1167);
and U2377 (N_2377,N_1336,N_1374);
nand U2378 (N_2378,N_1494,N_1245);
nor U2379 (N_2379,N_1299,N_1515);
xor U2380 (N_2380,N_1921,N_1193);
nand U2381 (N_2381,N_1460,N_1628);
and U2382 (N_2382,N_1388,N_1454);
xnor U2383 (N_2383,N_1361,N_1654);
or U2384 (N_2384,N_1904,N_1632);
and U2385 (N_2385,N_1772,N_1670);
nand U2386 (N_2386,N_1994,N_1132);
xnor U2387 (N_2387,N_1219,N_1865);
and U2388 (N_2388,N_1495,N_1505);
nor U2389 (N_2389,N_1697,N_1352);
nand U2390 (N_2390,N_1604,N_1264);
and U2391 (N_2391,N_1301,N_1719);
nand U2392 (N_2392,N_1662,N_1197);
nor U2393 (N_2393,N_1412,N_1295);
or U2394 (N_2394,N_1019,N_1387);
nor U2395 (N_2395,N_1546,N_1337);
and U2396 (N_2396,N_1983,N_1350);
and U2397 (N_2397,N_1092,N_1700);
nand U2398 (N_2398,N_1810,N_1839);
nor U2399 (N_2399,N_1083,N_1059);
and U2400 (N_2400,N_1037,N_1380);
or U2401 (N_2401,N_1192,N_1928);
nand U2402 (N_2402,N_1233,N_1912);
or U2403 (N_2403,N_1941,N_1725);
nor U2404 (N_2404,N_1082,N_1317);
nand U2405 (N_2405,N_1550,N_1183);
nor U2406 (N_2406,N_1172,N_1449);
nor U2407 (N_2407,N_1665,N_1415);
or U2408 (N_2408,N_1118,N_1790);
or U2409 (N_2409,N_1414,N_1466);
or U2410 (N_2410,N_1710,N_1527);
nand U2411 (N_2411,N_1366,N_1690);
nand U2412 (N_2412,N_1968,N_1120);
nor U2413 (N_2413,N_1557,N_1949);
xor U2414 (N_2414,N_1399,N_1497);
nand U2415 (N_2415,N_1758,N_1922);
nor U2416 (N_2416,N_1255,N_1583);
nand U2417 (N_2417,N_1006,N_1558);
nand U2418 (N_2418,N_1237,N_1062);
nand U2419 (N_2419,N_1718,N_1770);
and U2420 (N_2420,N_1599,N_1080);
nand U2421 (N_2421,N_1051,N_1773);
and U2422 (N_2422,N_1566,N_1122);
nand U2423 (N_2423,N_1487,N_1217);
nor U2424 (N_2424,N_1114,N_1640);
or U2425 (N_2425,N_1474,N_1365);
nand U2426 (N_2426,N_1844,N_1135);
and U2427 (N_2427,N_1102,N_1658);
and U2428 (N_2428,N_1369,N_1258);
or U2429 (N_2429,N_1577,N_1740);
nor U2430 (N_2430,N_1302,N_1813);
and U2431 (N_2431,N_1678,N_1313);
or U2432 (N_2432,N_1995,N_1981);
or U2433 (N_2433,N_1251,N_1959);
or U2434 (N_2434,N_1862,N_1345);
and U2435 (N_2435,N_1133,N_1944);
nor U2436 (N_2436,N_1097,N_1787);
or U2437 (N_2437,N_1581,N_1382);
nand U2438 (N_2438,N_1046,N_1042);
nand U2439 (N_2439,N_1651,N_1339);
nand U2440 (N_2440,N_1231,N_1163);
nand U2441 (N_2441,N_1956,N_1517);
nor U2442 (N_2442,N_1075,N_1588);
nor U2443 (N_2443,N_1203,N_1433);
or U2444 (N_2444,N_1960,N_1372);
nor U2445 (N_2445,N_1159,N_1954);
or U2446 (N_2446,N_1969,N_1655);
xor U2447 (N_2447,N_1516,N_1185);
nand U2448 (N_2448,N_1155,N_1645);
nand U2449 (N_2449,N_1180,N_1349);
nor U2450 (N_2450,N_1408,N_1743);
and U2451 (N_2451,N_1829,N_1646);
nand U2452 (N_2452,N_1060,N_1012);
and U2453 (N_2453,N_1663,N_1664);
xnor U2454 (N_2454,N_1521,N_1637);
nand U2455 (N_2455,N_1974,N_1017);
and U2456 (N_2456,N_1853,N_1986);
and U2457 (N_2457,N_1522,N_1014);
nand U2458 (N_2458,N_1910,N_1868);
and U2459 (N_2459,N_1015,N_1177);
xnor U2460 (N_2460,N_1620,N_1603);
and U2461 (N_2461,N_1764,N_1935);
and U2462 (N_2462,N_1530,N_1007);
nor U2463 (N_2463,N_1196,N_1595);
xnor U2464 (N_2464,N_1392,N_1241);
or U2465 (N_2465,N_1363,N_1134);
nand U2466 (N_2466,N_1882,N_1819);
nand U2467 (N_2467,N_1107,N_1592);
nand U2468 (N_2468,N_1063,N_1602);
or U2469 (N_2469,N_1484,N_1746);
and U2470 (N_2470,N_1189,N_1171);
nand U2471 (N_2471,N_1278,N_1204);
nand U2472 (N_2472,N_1518,N_1215);
and U2473 (N_2473,N_1673,N_1753);
or U2474 (N_2474,N_1305,N_1553);
and U2475 (N_2475,N_1249,N_1705);
or U2476 (N_2476,N_1404,N_1202);
xor U2477 (N_2477,N_1800,N_1752);
or U2478 (N_2478,N_1572,N_1513);
nor U2479 (N_2479,N_1357,N_1623);
and U2480 (N_2480,N_1791,N_1027);
nand U2481 (N_2481,N_1565,N_1777);
nand U2482 (N_2482,N_1179,N_1206);
nand U2483 (N_2483,N_1833,N_1478);
or U2484 (N_2484,N_1343,N_1559);
and U2485 (N_2485,N_1501,N_1307);
or U2486 (N_2486,N_1072,N_1428);
nor U2487 (N_2487,N_1115,N_1919);
nor U2488 (N_2488,N_1680,N_1304);
nand U2489 (N_2489,N_1687,N_1090);
and U2490 (N_2490,N_1243,N_1220);
nor U2491 (N_2491,N_1230,N_1869);
nor U2492 (N_2492,N_1931,N_1310);
or U2493 (N_2493,N_1330,N_1917);
nor U2494 (N_2494,N_1312,N_1489);
and U2495 (N_2495,N_1943,N_1153);
nand U2496 (N_2496,N_1715,N_1587);
nor U2497 (N_2497,N_1750,N_1208);
nor U2498 (N_2498,N_1507,N_1280);
and U2499 (N_2499,N_1426,N_1593);
and U2500 (N_2500,N_1909,N_1147);
or U2501 (N_2501,N_1902,N_1529);
and U2502 (N_2502,N_1310,N_1603);
xor U2503 (N_2503,N_1613,N_1614);
nor U2504 (N_2504,N_1507,N_1105);
nor U2505 (N_2505,N_1033,N_1671);
and U2506 (N_2506,N_1449,N_1662);
or U2507 (N_2507,N_1298,N_1192);
nand U2508 (N_2508,N_1170,N_1212);
and U2509 (N_2509,N_1655,N_1083);
nand U2510 (N_2510,N_1139,N_1573);
nand U2511 (N_2511,N_1765,N_1788);
or U2512 (N_2512,N_1849,N_1739);
nand U2513 (N_2513,N_1739,N_1870);
nor U2514 (N_2514,N_1143,N_1617);
nand U2515 (N_2515,N_1190,N_1706);
and U2516 (N_2516,N_1104,N_1463);
or U2517 (N_2517,N_1019,N_1361);
or U2518 (N_2518,N_1484,N_1698);
nor U2519 (N_2519,N_1332,N_1760);
xnor U2520 (N_2520,N_1705,N_1414);
nor U2521 (N_2521,N_1864,N_1077);
and U2522 (N_2522,N_1648,N_1567);
nor U2523 (N_2523,N_1980,N_1458);
nand U2524 (N_2524,N_1907,N_1397);
and U2525 (N_2525,N_1607,N_1579);
nand U2526 (N_2526,N_1250,N_1817);
nand U2527 (N_2527,N_1400,N_1545);
nand U2528 (N_2528,N_1930,N_1919);
and U2529 (N_2529,N_1133,N_1906);
nand U2530 (N_2530,N_1524,N_1799);
or U2531 (N_2531,N_1053,N_1786);
nor U2532 (N_2532,N_1545,N_1516);
or U2533 (N_2533,N_1356,N_1432);
xor U2534 (N_2534,N_1014,N_1434);
nand U2535 (N_2535,N_1740,N_1672);
xnor U2536 (N_2536,N_1624,N_1836);
nand U2537 (N_2537,N_1760,N_1060);
nor U2538 (N_2538,N_1957,N_1489);
xor U2539 (N_2539,N_1930,N_1897);
nor U2540 (N_2540,N_1136,N_1750);
nor U2541 (N_2541,N_1389,N_1515);
xor U2542 (N_2542,N_1396,N_1355);
or U2543 (N_2543,N_1122,N_1752);
or U2544 (N_2544,N_1167,N_1379);
or U2545 (N_2545,N_1209,N_1530);
or U2546 (N_2546,N_1580,N_1669);
and U2547 (N_2547,N_1116,N_1792);
or U2548 (N_2548,N_1167,N_1714);
nor U2549 (N_2549,N_1155,N_1353);
or U2550 (N_2550,N_1930,N_1052);
nor U2551 (N_2551,N_1994,N_1471);
xnor U2552 (N_2552,N_1039,N_1481);
nor U2553 (N_2553,N_1385,N_1355);
or U2554 (N_2554,N_1639,N_1862);
nand U2555 (N_2555,N_1879,N_1930);
xor U2556 (N_2556,N_1651,N_1461);
or U2557 (N_2557,N_1050,N_1063);
or U2558 (N_2558,N_1806,N_1778);
nand U2559 (N_2559,N_1002,N_1110);
nor U2560 (N_2560,N_1268,N_1967);
xnor U2561 (N_2561,N_1444,N_1420);
nor U2562 (N_2562,N_1538,N_1768);
xnor U2563 (N_2563,N_1470,N_1732);
nand U2564 (N_2564,N_1525,N_1277);
nand U2565 (N_2565,N_1718,N_1128);
nor U2566 (N_2566,N_1154,N_1752);
nor U2567 (N_2567,N_1446,N_1582);
or U2568 (N_2568,N_1327,N_1316);
xor U2569 (N_2569,N_1230,N_1127);
nor U2570 (N_2570,N_1222,N_1971);
or U2571 (N_2571,N_1123,N_1168);
nand U2572 (N_2572,N_1557,N_1090);
and U2573 (N_2573,N_1979,N_1298);
nor U2574 (N_2574,N_1645,N_1324);
or U2575 (N_2575,N_1683,N_1911);
nor U2576 (N_2576,N_1889,N_1150);
xnor U2577 (N_2577,N_1801,N_1939);
nor U2578 (N_2578,N_1400,N_1216);
or U2579 (N_2579,N_1877,N_1671);
xor U2580 (N_2580,N_1731,N_1853);
nand U2581 (N_2581,N_1286,N_1295);
nand U2582 (N_2582,N_1896,N_1236);
nand U2583 (N_2583,N_1237,N_1348);
xnor U2584 (N_2584,N_1800,N_1141);
and U2585 (N_2585,N_1744,N_1606);
and U2586 (N_2586,N_1574,N_1604);
nand U2587 (N_2587,N_1323,N_1794);
nand U2588 (N_2588,N_1890,N_1285);
and U2589 (N_2589,N_1067,N_1193);
and U2590 (N_2590,N_1676,N_1420);
nand U2591 (N_2591,N_1385,N_1899);
nor U2592 (N_2592,N_1047,N_1498);
and U2593 (N_2593,N_1181,N_1393);
xnor U2594 (N_2594,N_1703,N_1444);
and U2595 (N_2595,N_1894,N_1921);
nor U2596 (N_2596,N_1562,N_1851);
nand U2597 (N_2597,N_1819,N_1672);
nor U2598 (N_2598,N_1571,N_1590);
xor U2599 (N_2599,N_1721,N_1536);
and U2600 (N_2600,N_1185,N_1255);
nor U2601 (N_2601,N_1561,N_1042);
or U2602 (N_2602,N_1348,N_1981);
nor U2603 (N_2603,N_1455,N_1634);
and U2604 (N_2604,N_1865,N_1479);
xor U2605 (N_2605,N_1487,N_1277);
nor U2606 (N_2606,N_1908,N_1527);
nand U2607 (N_2607,N_1853,N_1328);
and U2608 (N_2608,N_1458,N_1236);
or U2609 (N_2609,N_1141,N_1136);
nor U2610 (N_2610,N_1979,N_1292);
nor U2611 (N_2611,N_1221,N_1096);
or U2612 (N_2612,N_1918,N_1520);
or U2613 (N_2613,N_1598,N_1962);
nor U2614 (N_2614,N_1254,N_1053);
nand U2615 (N_2615,N_1514,N_1470);
nor U2616 (N_2616,N_1636,N_1598);
nor U2617 (N_2617,N_1206,N_1718);
nand U2618 (N_2618,N_1881,N_1716);
nand U2619 (N_2619,N_1430,N_1243);
nor U2620 (N_2620,N_1500,N_1015);
nand U2621 (N_2621,N_1161,N_1438);
or U2622 (N_2622,N_1707,N_1672);
nor U2623 (N_2623,N_1949,N_1382);
and U2624 (N_2624,N_1295,N_1515);
and U2625 (N_2625,N_1052,N_1240);
nor U2626 (N_2626,N_1172,N_1657);
or U2627 (N_2627,N_1976,N_1063);
and U2628 (N_2628,N_1848,N_1873);
or U2629 (N_2629,N_1413,N_1031);
nor U2630 (N_2630,N_1750,N_1253);
or U2631 (N_2631,N_1456,N_1875);
nand U2632 (N_2632,N_1800,N_1847);
nand U2633 (N_2633,N_1126,N_1644);
nand U2634 (N_2634,N_1704,N_1786);
or U2635 (N_2635,N_1621,N_1990);
nor U2636 (N_2636,N_1861,N_1404);
and U2637 (N_2637,N_1561,N_1750);
or U2638 (N_2638,N_1093,N_1107);
or U2639 (N_2639,N_1732,N_1347);
nor U2640 (N_2640,N_1809,N_1059);
or U2641 (N_2641,N_1137,N_1270);
nor U2642 (N_2642,N_1383,N_1738);
nor U2643 (N_2643,N_1268,N_1408);
or U2644 (N_2644,N_1548,N_1090);
or U2645 (N_2645,N_1497,N_1776);
and U2646 (N_2646,N_1534,N_1199);
xor U2647 (N_2647,N_1975,N_1003);
and U2648 (N_2648,N_1408,N_1869);
xor U2649 (N_2649,N_1104,N_1790);
xnor U2650 (N_2650,N_1519,N_1851);
xor U2651 (N_2651,N_1790,N_1943);
and U2652 (N_2652,N_1285,N_1570);
xor U2653 (N_2653,N_1330,N_1391);
and U2654 (N_2654,N_1632,N_1129);
nand U2655 (N_2655,N_1637,N_1907);
nor U2656 (N_2656,N_1907,N_1842);
nor U2657 (N_2657,N_1185,N_1271);
xnor U2658 (N_2658,N_1870,N_1542);
nand U2659 (N_2659,N_1728,N_1716);
nand U2660 (N_2660,N_1021,N_1925);
or U2661 (N_2661,N_1385,N_1888);
or U2662 (N_2662,N_1804,N_1380);
xnor U2663 (N_2663,N_1003,N_1123);
or U2664 (N_2664,N_1360,N_1050);
and U2665 (N_2665,N_1890,N_1470);
nand U2666 (N_2666,N_1913,N_1343);
nand U2667 (N_2667,N_1746,N_1124);
and U2668 (N_2668,N_1227,N_1850);
or U2669 (N_2669,N_1376,N_1917);
or U2670 (N_2670,N_1596,N_1710);
and U2671 (N_2671,N_1837,N_1902);
or U2672 (N_2672,N_1084,N_1945);
nand U2673 (N_2673,N_1200,N_1788);
and U2674 (N_2674,N_1082,N_1961);
or U2675 (N_2675,N_1748,N_1929);
nand U2676 (N_2676,N_1953,N_1179);
nand U2677 (N_2677,N_1286,N_1072);
nand U2678 (N_2678,N_1199,N_1417);
nor U2679 (N_2679,N_1142,N_1984);
and U2680 (N_2680,N_1740,N_1616);
nand U2681 (N_2681,N_1456,N_1007);
nor U2682 (N_2682,N_1960,N_1539);
nand U2683 (N_2683,N_1890,N_1899);
nor U2684 (N_2684,N_1292,N_1073);
or U2685 (N_2685,N_1465,N_1951);
nor U2686 (N_2686,N_1264,N_1684);
nand U2687 (N_2687,N_1956,N_1054);
nor U2688 (N_2688,N_1239,N_1939);
or U2689 (N_2689,N_1400,N_1214);
xnor U2690 (N_2690,N_1878,N_1157);
nand U2691 (N_2691,N_1171,N_1771);
and U2692 (N_2692,N_1788,N_1227);
xor U2693 (N_2693,N_1662,N_1271);
and U2694 (N_2694,N_1185,N_1480);
nor U2695 (N_2695,N_1601,N_1446);
and U2696 (N_2696,N_1478,N_1904);
and U2697 (N_2697,N_1064,N_1830);
and U2698 (N_2698,N_1251,N_1080);
nand U2699 (N_2699,N_1910,N_1153);
or U2700 (N_2700,N_1924,N_1348);
nand U2701 (N_2701,N_1735,N_1506);
or U2702 (N_2702,N_1450,N_1677);
and U2703 (N_2703,N_1899,N_1572);
or U2704 (N_2704,N_1510,N_1731);
nor U2705 (N_2705,N_1199,N_1112);
and U2706 (N_2706,N_1626,N_1544);
and U2707 (N_2707,N_1171,N_1954);
nor U2708 (N_2708,N_1795,N_1438);
and U2709 (N_2709,N_1779,N_1019);
or U2710 (N_2710,N_1571,N_1350);
or U2711 (N_2711,N_1345,N_1610);
and U2712 (N_2712,N_1348,N_1107);
nor U2713 (N_2713,N_1769,N_1136);
xor U2714 (N_2714,N_1864,N_1369);
nor U2715 (N_2715,N_1391,N_1010);
and U2716 (N_2716,N_1872,N_1604);
nor U2717 (N_2717,N_1381,N_1694);
or U2718 (N_2718,N_1891,N_1248);
xnor U2719 (N_2719,N_1036,N_1550);
nand U2720 (N_2720,N_1730,N_1160);
xnor U2721 (N_2721,N_1554,N_1269);
and U2722 (N_2722,N_1755,N_1227);
nand U2723 (N_2723,N_1229,N_1958);
or U2724 (N_2724,N_1970,N_1774);
nor U2725 (N_2725,N_1396,N_1618);
nand U2726 (N_2726,N_1043,N_1092);
and U2727 (N_2727,N_1175,N_1695);
nor U2728 (N_2728,N_1402,N_1434);
and U2729 (N_2729,N_1263,N_1236);
or U2730 (N_2730,N_1818,N_1495);
nor U2731 (N_2731,N_1183,N_1826);
and U2732 (N_2732,N_1123,N_1161);
nor U2733 (N_2733,N_1785,N_1849);
nand U2734 (N_2734,N_1081,N_1546);
nor U2735 (N_2735,N_1846,N_1180);
nor U2736 (N_2736,N_1476,N_1309);
and U2737 (N_2737,N_1164,N_1980);
or U2738 (N_2738,N_1309,N_1805);
nand U2739 (N_2739,N_1249,N_1348);
or U2740 (N_2740,N_1873,N_1163);
nand U2741 (N_2741,N_1155,N_1795);
nand U2742 (N_2742,N_1285,N_1408);
and U2743 (N_2743,N_1138,N_1160);
or U2744 (N_2744,N_1809,N_1552);
nand U2745 (N_2745,N_1306,N_1600);
or U2746 (N_2746,N_1023,N_1544);
nor U2747 (N_2747,N_1030,N_1578);
or U2748 (N_2748,N_1875,N_1357);
or U2749 (N_2749,N_1639,N_1843);
and U2750 (N_2750,N_1043,N_1819);
or U2751 (N_2751,N_1641,N_1302);
nor U2752 (N_2752,N_1251,N_1297);
nand U2753 (N_2753,N_1205,N_1760);
nor U2754 (N_2754,N_1298,N_1218);
and U2755 (N_2755,N_1599,N_1668);
nand U2756 (N_2756,N_1531,N_1572);
and U2757 (N_2757,N_1225,N_1608);
or U2758 (N_2758,N_1822,N_1576);
nor U2759 (N_2759,N_1109,N_1498);
nand U2760 (N_2760,N_1479,N_1594);
nor U2761 (N_2761,N_1047,N_1327);
and U2762 (N_2762,N_1588,N_1460);
nor U2763 (N_2763,N_1714,N_1801);
or U2764 (N_2764,N_1922,N_1975);
nor U2765 (N_2765,N_1161,N_1108);
nand U2766 (N_2766,N_1652,N_1491);
or U2767 (N_2767,N_1227,N_1488);
or U2768 (N_2768,N_1429,N_1918);
or U2769 (N_2769,N_1467,N_1025);
xor U2770 (N_2770,N_1232,N_1673);
nor U2771 (N_2771,N_1450,N_1570);
nand U2772 (N_2772,N_1084,N_1190);
and U2773 (N_2773,N_1667,N_1546);
nor U2774 (N_2774,N_1837,N_1765);
or U2775 (N_2775,N_1853,N_1826);
and U2776 (N_2776,N_1377,N_1839);
or U2777 (N_2777,N_1495,N_1593);
nand U2778 (N_2778,N_1509,N_1999);
xor U2779 (N_2779,N_1416,N_1758);
or U2780 (N_2780,N_1182,N_1920);
nand U2781 (N_2781,N_1163,N_1147);
and U2782 (N_2782,N_1469,N_1821);
and U2783 (N_2783,N_1791,N_1599);
or U2784 (N_2784,N_1590,N_1695);
nand U2785 (N_2785,N_1547,N_1710);
or U2786 (N_2786,N_1734,N_1586);
nand U2787 (N_2787,N_1018,N_1034);
nand U2788 (N_2788,N_1777,N_1971);
or U2789 (N_2789,N_1695,N_1319);
nor U2790 (N_2790,N_1608,N_1138);
nand U2791 (N_2791,N_1180,N_1602);
or U2792 (N_2792,N_1494,N_1750);
and U2793 (N_2793,N_1897,N_1603);
and U2794 (N_2794,N_1627,N_1292);
nand U2795 (N_2795,N_1162,N_1663);
nor U2796 (N_2796,N_1541,N_1638);
nand U2797 (N_2797,N_1215,N_1178);
xnor U2798 (N_2798,N_1158,N_1397);
or U2799 (N_2799,N_1783,N_1814);
nand U2800 (N_2800,N_1222,N_1543);
or U2801 (N_2801,N_1556,N_1689);
nor U2802 (N_2802,N_1950,N_1583);
nand U2803 (N_2803,N_1544,N_1620);
nand U2804 (N_2804,N_1983,N_1451);
nor U2805 (N_2805,N_1080,N_1810);
and U2806 (N_2806,N_1048,N_1556);
xnor U2807 (N_2807,N_1369,N_1132);
and U2808 (N_2808,N_1174,N_1556);
nor U2809 (N_2809,N_1935,N_1803);
or U2810 (N_2810,N_1770,N_1246);
nand U2811 (N_2811,N_1520,N_1113);
and U2812 (N_2812,N_1894,N_1222);
xnor U2813 (N_2813,N_1761,N_1365);
or U2814 (N_2814,N_1441,N_1950);
or U2815 (N_2815,N_1209,N_1018);
xor U2816 (N_2816,N_1626,N_1546);
nor U2817 (N_2817,N_1331,N_1658);
and U2818 (N_2818,N_1506,N_1092);
nand U2819 (N_2819,N_1101,N_1690);
xnor U2820 (N_2820,N_1678,N_1696);
and U2821 (N_2821,N_1789,N_1280);
nor U2822 (N_2822,N_1918,N_1666);
and U2823 (N_2823,N_1154,N_1038);
xor U2824 (N_2824,N_1985,N_1948);
nand U2825 (N_2825,N_1168,N_1947);
or U2826 (N_2826,N_1770,N_1332);
nand U2827 (N_2827,N_1249,N_1273);
xnor U2828 (N_2828,N_1540,N_1059);
xnor U2829 (N_2829,N_1725,N_1243);
and U2830 (N_2830,N_1449,N_1896);
nand U2831 (N_2831,N_1040,N_1909);
nand U2832 (N_2832,N_1783,N_1081);
and U2833 (N_2833,N_1944,N_1912);
or U2834 (N_2834,N_1501,N_1706);
nand U2835 (N_2835,N_1185,N_1966);
nor U2836 (N_2836,N_1714,N_1214);
nor U2837 (N_2837,N_1714,N_1587);
nor U2838 (N_2838,N_1142,N_1004);
and U2839 (N_2839,N_1511,N_1437);
and U2840 (N_2840,N_1813,N_1022);
or U2841 (N_2841,N_1818,N_1757);
nand U2842 (N_2842,N_1223,N_1502);
and U2843 (N_2843,N_1206,N_1912);
nand U2844 (N_2844,N_1434,N_1520);
nor U2845 (N_2845,N_1624,N_1648);
nor U2846 (N_2846,N_1094,N_1977);
nor U2847 (N_2847,N_1031,N_1170);
and U2848 (N_2848,N_1271,N_1191);
and U2849 (N_2849,N_1810,N_1252);
or U2850 (N_2850,N_1481,N_1802);
nand U2851 (N_2851,N_1019,N_1773);
nand U2852 (N_2852,N_1256,N_1411);
xnor U2853 (N_2853,N_1717,N_1771);
and U2854 (N_2854,N_1813,N_1077);
nand U2855 (N_2855,N_1935,N_1870);
nor U2856 (N_2856,N_1715,N_1002);
and U2857 (N_2857,N_1595,N_1163);
or U2858 (N_2858,N_1604,N_1061);
nor U2859 (N_2859,N_1131,N_1783);
and U2860 (N_2860,N_1552,N_1917);
and U2861 (N_2861,N_1677,N_1345);
or U2862 (N_2862,N_1492,N_1324);
or U2863 (N_2863,N_1913,N_1648);
xor U2864 (N_2864,N_1060,N_1884);
nor U2865 (N_2865,N_1467,N_1676);
nand U2866 (N_2866,N_1659,N_1119);
nand U2867 (N_2867,N_1760,N_1807);
nand U2868 (N_2868,N_1146,N_1219);
nand U2869 (N_2869,N_1349,N_1586);
and U2870 (N_2870,N_1806,N_1901);
and U2871 (N_2871,N_1567,N_1322);
nand U2872 (N_2872,N_1394,N_1356);
xnor U2873 (N_2873,N_1656,N_1770);
or U2874 (N_2874,N_1385,N_1054);
nor U2875 (N_2875,N_1251,N_1456);
nor U2876 (N_2876,N_1960,N_1894);
nand U2877 (N_2877,N_1338,N_1841);
nand U2878 (N_2878,N_1890,N_1446);
nand U2879 (N_2879,N_1729,N_1681);
nor U2880 (N_2880,N_1066,N_1277);
or U2881 (N_2881,N_1165,N_1992);
nand U2882 (N_2882,N_1410,N_1439);
or U2883 (N_2883,N_1805,N_1408);
or U2884 (N_2884,N_1616,N_1794);
or U2885 (N_2885,N_1459,N_1771);
nand U2886 (N_2886,N_1899,N_1813);
nand U2887 (N_2887,N_1578,N_1327);
nand U2888 (N_2888,N_1321,N_1731);
nand U2889 (N_2889,N_1167,N_1285);
nor U2890 (N_2890,N_1816,N_1010);
and U2891 (N_2891,N_1284,N_1100);
and U2892 (N_2892,N_1067,N_1399);
nand U2893 (N_2893,N_1472,N_1522);
and U2894 (N_2894,N_1723,N_1043);
or U2895 (N_2895,N_1747,N_1084);
or U2896 (N_2896,N_1222,N_1795);
nand U2897 (N_2897,N_1856,N_1186);
or U2898 (N_2898,N_1499,N_1545);
or U2899 (N_2899,N_1018,N_1768);
nor U2900 (N_2900,N_1086,N_1398);
and U2901 (N_2901,N_1125,N_1172);
nor U2902 (N_2902,N_1738,N_1897);
or U2903 (N_2903,N_1756,N_1339);
xor U2904 (N_2904,N_1468,N_1164);
or U2905 (N_2905,N_1674,N_1714);
and U2906 (N_2906,N_1967,N_1309);
nor U2907 (N_2907,N_1828,N_1469);
or U2908 (N_2908,N_1893,N_1219);
and U2909 (N_2909,N_1048,N_1975);
or U2910 (N_2910,N_1604,N_1380);
nand U2911 (N_2911,N_1432,N_1871);
xor U2912 (N_2912,N_1321,N_1178);
nand U2913 (N_2913,N_1845,N_1796);
or U2914 (N_2914,N_1423,N_1911);
nand U2915 (N_2915,N_1209,N_1276);
nand U2916 (N_2916,N_1399,N_1767);
nand U2917 (N_2917,N_1428,N_1190);
and U2918 (N_2918,N_1381,N_1612);
and U2919 (N_2919,N_1155,N_1047);
or U2920 (N_2920,N_1878,N_1529);
nand U2921 (N_2921,N_1024,N_1505);
nor U2922 (N_2922,N_1071,N_1647);
and U2923 (N_2923,N_1057,N_1433);
xor U2924 (N_2924,N_1178,N_1591);
and U2925 (N_2925,N_1108,N_1470);
and U2926 (N_2926,N_1469,N_1749);
xor U2927 (N_2927,N_1235,N_1521);
and U2928 (N_2928,N_1416,N_1991);
or U2929 (N_2929,N_1221,N_1273);
or U2930 (N_2930,N_1194,N_1686);
and U2931 (N_2931,N_1230,N_1269);
nand U2932 (N_2932,N_1413,N_1039);
nand U2933 (N_2933,N_1333,N_1452);
and U2934 (N_2934,N_1017,N_1625);
nor U2935 (N_2935,N_1578,N_1658);
or U2936 (N_2936,N_1685,N_1080);
or U2937 (N_2937,N_1634,N_1907);
and U2938 (N_2938,N_1314,N_1614);
or U2939 (N_2939,N_1927,N_1610);
xor U2940 (N_2940,N_1162,N_1130);
and U2941 (N_2941,N_1382,N_1958);
nor U2942 (N_2942,N_1337,N_1267);
and U2943 (N_2943,N_1047,N_1001);
or U2944 (N_2944,N_1760,N_1781);
or U2945 (N_2945,N_1824,N_1408);
and U2946 (N_2946,N_1723,N_1393);
nor U2947 (N_2947,N_1164,N_1429);
nand U2948 (N_2948,N_1721,N_1167);
nand U2949 (N_2949,N_1272,N_1758);
and U2950 (N_2950,N_1614,N_1554);
and U2951 (N_2951,N_1177,N_1578);
or U2952 (N_2952,N_1426,N_1177);
nand U2953 (N_2953,N_1906,N_1450);
nor U2954 (N_2954,N_1575,N_1238);
or U2955 (N_2955,N_1021,N_1593);
xnor U2956 (N_2956,N_1783,N_1823);
and U2957 (N_2957,N_1937,N_1501);
xnor U2958 (N_2958,N_1159,N_1956);
or U2959 (N_2959,N_1082,N_1457);
and U2960 (N_2960,N_1116,N_1651);
and U2961 (N_2961,N_1237,N_1880);
or U2962 (N_2962,N_1287,N_1528);
or U2963 (N_2963,N_1562,N_1802);
and U2964 (N_2964,N_1354,N_1046);
nand U2965 (N_2965,N_1210,N_1545);
and U2966 (N_2966,N_1945,N_1859);
or U2967 (N_2967,N_1580,N_1897);
nand U2968 (N_2968,N_1605,N_1881);
or U2969 (N_2969,N_1725,N_1805);
or U2970 (N_2970,N_1392,N_1513);
nor U2971 (N_2971,N_1129,N_1438);
nor U2972 (N_2972,N_1995,N_1437);
xnor U2973 (N_2973,N_1158,N_1656);
nand U2974 (N_2974,N_1920,N_1030);
nor U2975 (N_2975,N_1155,N_1196);
nand U2976 (N_2976,N_1150,N_1993);
nor U2977 (N_2977,N_1193,N_1184);
or U2978 (N_2978,N_1174,N_1045);
nor U2979 (N_2979,N_1449,N_1063);
xor U2980 (N_2980,N_1422,N_1852);
nor U2981 (N_2981,N_1806,N_1796);
nand U2982 (N_2982,N_1094,N_1719);
nand U2983 (N_2983,N_1700,N_1326);
and U2984 (N_2984,N_1120,N_1195);
and U2985 (N_2985,N_1996,N_1584);
nand U2986 (N_2986,N_1282,N_1674);
or U2987 (N_2987,N_1541,N_1043);
xnor U2988 (N_2988,N_1841,N_1007);
nor U2989 (N_2989,N_1495,N_1848);
or U2990 (N_2990,N_1432,N_1887);
nand U2991 (N_2991,N_1211,N_1913);
nor U2992 (N_2992,N_1323,N_1233);
nand U2993 (N_2993,N_1335,N_1808);
or U2994 (N_2994,N_1045,N_1197);
nor U2995 (N_2995,N_1332,N_1172);
nor U2996 (N_2996,N_1785,N_1276);
nand U2997 (N_2997,N_1578,N_1541);
nand U2998 (N_2998,N_1961,N_1398);
or U2999 (N_2999,N_1209,N_1168);
xor UO_0 (O_0,N_2062,N_2567);
and UO_1 (O_1,N_2940,N_2626);
or UO_2 (O_2,N_2256,N_2067);
or UO_3 (O_3,N_2370,N_2772);
and UO_4 (O_4,N_2112,N_2205);
or UO_5 (O_5,N_2391,N_2155);
nor UO_6 (O_6,N_2100,N_2470);
or UO_7 (O_7,N_2573,N_2635);
nor UO_8 (O_8,N_2545,N_2597);
nand UO_9 (O_9,N_2342,N_2608);
or UO_10 (O_10,N_2394,N_2739);
nand UO_11 (O_11,N_2510,N_2787);
and UO_12 (O_12,N_2263,N_2761);
and UO_13 (O_13,N_2847,N_2704);
or UO_14 (O_14,N_2238,N_2583);
and UO_15 (O_15,N_2601,N_2233);
nand UO_16 (O_16,N_2445,N_2329);
nand UO_17 (O_17,N_2364,N_2544);
nand UO_18 (O_18,N_2165,N_2886);
nor UO_19 (O_19,N_2482,N_2507);
nor UO_20 (O_20,N_2616,N_2582);
and UO_21 (O_21,N_2865,N_2564);
nor UO_22 (O_22,N_2160,N_2110);
nor UO_23 (O_23,N_2088,N_2326);
nand UO_24 (O_24,N_2817,N_2453);
or UO_25 (O_25,N_2887,N_2462);
xor UO_26 (O_26,N_2141,N_2953);
xnor UO_27 (O_27,N_2825,N_2296);
and UO_28 (O_28,N_2841,N_2820);
and UO_29 (O_29,N_2192,N_2011);
or UO_30 (O_30,N_2099,N_2487);
nor UO_31 (O_31,N_2667,N_2810);
or UO_32 (O_32,N_2656,N_2882);
nor UO_33 (O_33,N_2707,N_2036);
or UO_34 (O_34,N_2410,N_2786);
and UO_35 (O_35,N_2148,N_2409);
or UO_36 (O_36,N_2388,N_2383);
nand UO_37 (O_37,N_2389,N_2004);
or UO_38 (O_38,N_2987,N_2982);
nand UO_39 (O_39,N_2999,N_2915);
and UO_40 (O_40,N_2513,N_2625);
nand UO_41 (O_41,N_2857,N_2368);
or UO_42 (O_42,N_2254,N_2925);
nand UO_43 (O_43,N_2087,N_2900);
or UO_44 (O_44,N_2349,N_2217);
xor UO_45 (O_45,N_2423,N_2691);
nor UO_46 (O_46,N_2203,N_2279);
or UO_47 (O_47,N_2491,N_2788);
nor UO_48 (O_48,N_2541,N_2064);
and UO_49 (O_49,N_2251,N_2655);
or UO_50 (O_50,N_2873,N_2901);
xor UO_51 (O_51,N_2271,N_2629);
and UO_52 (O_52,N_2664,N_2645);
xnor UO_53 (O_53,N_2435,N_2913);
nor UO_54 (O_54,N_2752,N_2669);
and UO_55 (O_55,N_2014,N_2909);
and UO_56 (O_56,N_2027,N_2756);
nand UO_57 (O_57,N_2800,N_2056);
nor UO_58 (O_58,N_2240,N_2869);
nor UO_59 (O_59,N_2313,N_2749);
xor UO_60 (O_60,N_2399,N_2611);
nand UO_61 (O_61,N_2016,N_2047);
or UO_62 (O_62,N_2782,N_2805);
nor UO_63 (O_63,N_2366,N_2017);
nand UO_64 (O_64,N_2277,N_2535);
nand UO_65 (O_65,N_2990,N_2652);
and UO_66 (O_66,N_2429,N_2317);
nand UO_67 (O_67,N_2996,N_2098);
nor UO_68 (O_68,N_2194,N_2933);
or UO_69 (O_69,N_2292,N_2357);
nor UO_70 (O_70,N_2499,N_2159);
nor UO_71 (O_71,N_2741,N_2730);
xor UO_72 (O_72,N_2815,N_2559);
nand UO_73 (O_73,N_2289,N_2031);
nor UO_74 (O_74,N_2469,N_2145);
nand UO_75 (O_75,N_2034,N_2899);
nand UO_76 (O_76,N_2187,N_2729);
and UO_77 (O_77,N_2848,N_2673);
nand UO_78 (O_78,N_2533,N_2236);
and UO_79 (O_79,N_2662,N_2688);
nand UO_80 (O_80,N_2035,N_2526);
or UO_81 (O_81,N_2924,N_2089);
nand UO_82 (O_82,N_2705,N_2387);
and UO_83 (O_83,N_2699,N_2127);
nand UO_84 (O_84,N_2576,N_2044);
nand UO_85 (O_85,N_2717,N_2854);
and UO_86 (O_86,N_2527,N_2822);
or UO_87 (O_87,N_2651,N_2604);
nand UO_88 (O_88,N_2703,N_2781);
or UO_89 (O_89,N_2091,N_2823);
or UO_90 (O_90,N_2128,N_2419);
nor UO_91 (O_91,N_2175,N_2740);
and UO_92 (O_92,N_2613,N_2144);
nand UO_93 (O_93,N_2392,N_2341);
and UO_94 (O_94,N_2606,N_2109);
nor UO_95 (O_95,N_2328,N_2577);
xor UO_96 (O_96,N_2977,N_2884);
nor UO_97 (O_97,N_2006,N_2138);
nor UO_98 (O_98,N_2026,N_2037);
nand UO_99 (O_99,N_2280,N_2104);
and UO_100 (O_100,N_2492,N_2167);
or UO_101 (O_101,N_2428,N_2307);
nor UO_102 (O_102,N_2022,N_2182);
or UO_103 (O_103,N_2695,N_2442);
and UO_104 (O_104,N_2605,N_2052);
or UO_105 (O_105,N_2747,N_2952);
and UO_106 (O_106,N_2369,N_2090);
or UO_107 (O_107,N_2759,N_2065);
xnor UO_108 (O_108,N_2665,N_2614);
or UO_109 (O_109,N_2060,N_2731);
and UO_110 (O_110,N_2550,N_2157);
and UO_111 (O_111,N_2654,N_2690);
nor UO_112 (O_112,N_2556,N_2287);
and UO_113 (O_113,N_2201,N_2745);
xor UO_114 (O_114,N_2166,N_2255);
nor UO_115 (O_115,N_2393,N_2769);
nand UO_116 (O_116,N_2072,N_2261);
nor UO_117 (O_117,N_2496,N_2177);
nor UO_118 (O_118,N_2042,N_2129);
and UO_119 (O_119,N_2984,N_2571);
or UO_120 (O_120,N_2385,N_2627);
and UO_121 (O_121,N_2743,N_2454);
and UO_122 (O_122,N_2966,N_2078);
or UO_123 (O_123,N_2168,N_2400);
and UO_124 (O_124,N_2404,N_2632);
and UO_125 (O_125,N_2637,N_2408);
nor UO_126 (O_126,N_2927,N_2377);
nor UO_127 (O_127,N_2944,N_2702);
nand UO_128 (O_128,N_2093,N_2914);
nand UO_129 (O_129,N_2521,N_2838);
xor UO_130 (O_130,N_2005,N_2790);
nand UO_131 (O_131,N_2003,N_2681);
nand UO_132 (O_132,N_2578,N_2241);
or UO_133 (O_133,N_2951,N_2242);
and UO_134 (O_134,N_2970,N_2853);
nand UO_135 (O_135,N_2860,N_2198);
nor UO_136 (O_136,N_2350,N_2497);
or UO_137 (O_137,N_2131,N_2053);
and UO_138 (O_138,N_2223,N_2552);
and UO_139 (O_139,N_2413,N_2542);
and UO_140 (O_140,N_2305,N_2284);
and UO_141 (O_141,N_2283,N_2232);
or UO_142 (O_142,N_2620,N_2967);
nand UO_143 (O_143,N_2602,N_2501);
or UO_144 (O_144,N_2579,N_2515);
nor UO_145 (O_145,N_2714,N_2495);
or UO_146 (O_146,N_2265,N_2021);
or UO_147 (O_147,N_2309,N_2178);
nand UO_148 (O_148,N_2939,N_2700);
nand UO_149 (O_149,N_2116,N_2184);
nor UO_150 (O_150,N_2123,N_2671);
and UO_151 (O_151,N_2845,N_2758);
nor UO_152 (O_152,N_2075,N_2268);
nand UO_153 (O_153,N_2360,N_2905);
nor UO_154 (O_154,N_2250,N_2523);
nor UO_155 (O_155,N_2776,N_2174);
and UO_156 (O_156,N_2694,N_2126);
nor UO_157 (O_157,N_2806,N_2051);
nand UO_158 (O_158,N_2992,N_2059);
and UO_159 (O_159,N_2932,N_2054);
nor UO_160 (O_160,N_2080,N_2386);
and UO_161 (O_161,N_2019,N_2903);
nand UO_162 (O_162,N_2281,N_2524);
nand UO_163 (O_163,N_2560,N_2146);
nand UO_164 (O_164,N_2612,N_2998);
or UO_165 (O_165,N_2343,N_2548);
nor UO_166 (O_166,N_2711,N_2956);
nor UO_167 (O_167,N_2594,N_2864);
xnor UO_168 (O_168,N_2319,N_2153);
and UO_169 (O_169,N_2898,N_2621);
nor UO_170 (O_170,N_2111,N_2101);
nor UO_171 (O_171,N_2529,N_2672);
nand UO_172 (O_172,N_2685,N_2460);
and UO_173 (O_173,N_2422,N_2249);
nor UO_174 (O_174,N_2757,N_2452);
nor UO_175 (O_175,N_2378,N_2512);
or UO_176 (O_176,N_2121,N_2530);
and UO_177 (O_177,N_2471,N_2943);
xnor UO_178 (O_178,N_2475,N_2798);
nand UO_179 (O_179,N_2143,N_2472);
and UO_180 (O_180,N_2151,N_2216);
nand UO_181 (O_181,N_2636,N_2096);
and UO_182 (O_182,N_2993,N_2013);
and UO_183 (O_183,N_2528,N_2816);
and UO_184 (O_184,N_2880,N_2398);
nor UO_185 (O_185,N_2630,N_2156);
and UO_186 (O_186,N_2963,N_2312);
and UO_187 (O_187,N_2457,N_2405);
or UO_188 (O_188,N_2338,N_2180);
nor UO_189 (O_189,N_2244,N_2683);
xnor UO_190 (O_190,N_2219,N_2796);
nor UO_191 (O_191,N_2354,N_2986);
nand UO_192 (O_192,N_2995,N_2546);
nor UO_193 (O_193,N_2768,N_2862);
and UO_194 (O_194,N_2079,N_2868);
xnor UO_195 (O_195,N_2975,N_2298);
or UO_196 (O_196,N_2193,N_2426);
or UO_197 (O_197,N_2981,N_2518);
nand UO_198 (O_198,N_2789,N_2103);
nand UO_199 (O_199,N_2808,N_2585);
xor UO_200 (O_200,N_2937,N_2173);
and UO_201 (O_201,N_2693,N_2359);
nor UO_202 (O_202,N_2425,N_2245);
xnor UO_203 (O_203,N_2661,N_2584);
and UO_204 (O_204,N_2874,N_2779);
nor UO_205 (O_205,N_2829,N_2553);
nor UO_206 (O_206,N_2588,N_2804);
or UO_207 (O_207,N_2765,N_2353);
nor UO_208 (O_208,N_2417,N_2696);
nand UO_209 (O_209,N_2437,N_2723);
or UO_210 (O_210,N_2911,N_2751);
nor UO_211 (O_211,N_2449,N_2498);
or UO_212 (O_212,N_2493,N_2722);
or UO_213 (O_213,N_2055,N_2340);
and UO_214 (O_214,N_2335,N_2839);
nor UO_215 (O_215,N_2861,N_2007);
nor UO_216 (O_216,N_2709,N_2331);
and UO_217 (O_217,N_2163,N_2412);
nor UO_218 (O_218,N_2916,N_2362);
or UO_219 (O_219,N_2118,N_2406);
xnor UO_220 (O_220,N_2397,N_2725);
or UO_221 (O_221,N_2721,N_2814);
or UO_222 (O_222,N_2226,N_2883);
xnor UO_223 (O_223,N_2907,N_2648);
xor UO_224 (O_224,N_2879,N_2274);
and UO_225 (O_225,N_2183,N_2234);
or UO_226 (O_226,N_2403,N_2070);
nand UO_227 (O_227,N_2023,N_2214);
xnor UO_228 (O_228,N_2971,N_2538);
nor UO_229 (O_229,N_2424,N_2554);
nor UO_230 (O_230,N_2311,N_2259);
or UO_231 (O_231,N_2285,N_2766);
nor UO_232 (O_232,N_2081,N_2069);
or UO_233 (O_233,N_2872,N_2902);
nor UO_234 (O_234,N_2888,N_2124);
nand UO_235 (O_235,N_2511,N_2107);
and UO_236 (O_236,N_2276,N_2117);
nand UO_237 (O_237,N_2633,N_2771);
or UO_238 (O_238,N_2959,N_2039);
and UO_239 (O_239,N_2945,N_2623);
nor UO_240 (O_240,N_2321,N_2459);
nor UO_241 (O_241,N_2742,N_2185);
nor UO_242 (O_242,N_2735,N_2622);
nor UO_243 (O_243,N_2097,N_2337);
nand UO_244 (O_244,N_2780,N_2955);
or UO_245 (O_245,N_2774,N_2293);
or UO_246 (O_246,N_2895,N_2172);
or UO_247 (O_247,N_2572,N_2674);
or UO_248 (O_248,N_2272,N_2028);
nand UO_249 (O_249,N_2962,N_2641);
xnor UO_250 (O_250,N_2969,N_2803);
nand UO_251 (O_251,N_2589,N_2720);
nor UO_252 (O_252,N_2684,N_2418);
or UO_253 (O_253,N_2303,N_2744);
xor UO_254 (O_254,N_2746,N_2231);
nor UO_255 (O_255,N_2777,N_2295);
nor UO_256 (O_256,N_2302,N_2191);
nand UO_257 (O_257,N_2373,N_2132);
nor UO_258 (O_258,N_2773,N_2033);
nand UO_259 (O_259,N_2867,N_2040);
or UO_260 (O_260,N_2140,N_2371);
and UO_261 (O_261,N_2767,N_2351);
nand UO_262 (O_262,N_2525,N_2610);
or UO_263 (O_263,N_2235,N_2195);
or UO_264 (O_264,N_2534,N_2164);
and UO_265 (O_265,N_2658,N_2018);
or UO_266 (O_266,N_2522,N_2257);
nor UO_267 (O_267,N_2586,N_2481);
and UO_268 (O_268,N_2108,N_2068);
or UO_269 (O_269,N_2802,N_2930);
or UO_270 (O_270,N_2569,N_2421);
and UO_271 (O_271,N_2954,N_2912);
and UO_272 (O_272,N_2269,N_2361);
nand UO_273 (O_273,N_2624,N_2563);
nor UO_274 (O_274,N_2300,N_2811);
nand UO_275 (O_275,N_2514,N_2414);
nor UO_276 (O_276,N_2503,N_2225);
nor UO_277 (O_277,N_2894,N_2716);
and UO_278 (O_278,N_2325,N_2537);
nand UO_279 (O_279,N_2327,N_2189);
nor UO_280 (O_280,N_2532,N_2119);
nor UO_281 (O_281,N_2352,N_2314);
nand UO_282 (O_282,N_2222,N_2439);
or UO_283 (O_283,N_2562,N_2575);
nand UO_284 (O_284,N_2607,N_2974);
xor UO_285 (O_285,N_2030,N_2032);
and UO_286 (O_286,N_2600,N_2543);
and UO_287 (O_287,N_2595,N_2547);
nand UO_288 (O_288,N_2920,N_2473);
nor UO_289 (O_289,N_2897,N_2540);
and UO_290 (O_290,N_2785,N_2456);
nand UO_291 (O_291,N_2332,N_2797);
nand UO_292 (O_292,N_2964,N_2836);
or UO_293 (O_293,N_2728,N_2947);
or UO_294 (O_294,N_2451,N_2137);
nand UO_295 (O_295,N_2881,N_2488);
xnor UO_296 (O_296,N_2994,N_2551);
or UO_297 (O_297,N_2666,N_2446);
and UO_298 (O_298,N_2390,N_2247);
nor UO_299 (O_299,N_2395,N_2372);
or UO_300 (O_300,N_2738,N_2643);
and UO_301 (O_301,N_2288,N_2381);
or UO_302 (O_302,N_2826,N_2972);
and UO_303 (O_303,N_2239,N_2008);
nor UO_304 (O_304,N_2015,N_2136);
or UO_305 (O_305,N_2082,N_2889);
nor UO_306 (O_306,N_2049,N_2443);
nand UO_307 (O_307,N_2447,N_2697);
nand UO_308 (O_308,N_2631,N_2983);
xor UO_309 (O_309,N_2850,N_2753);
or UO_310 (O_310,N_2333,N_2380);
nand UO_311 (O_311,N_2727,N_2149);
nor UO_312 (O_312,N_2948,N_2480);
or UO_313 (O_313,N_2230,N_2855);
nand UO_314 (O_314,N_2991,N_2025);
nand UO_315 (O_315,N_2593,N_2267);
nand UO_316 (O_316,N_2258,N_2336);
and UO_317 (O_317,N_2484,N_2890);
and UO_318 (O_318,N_2921,N_2659);
or UO_319 (O_319,N_2734,N_2286);
nor UO_320 (O_320,N_2415,N_2647);
nor UO_321 (O_321,N_2590,N_2821);
and UO_322 (O_322,N_2147,N_2807);
and UO_323 (O_323,N_2046,N_2210);
xnor UO_324 (O_324,N_2938,N_2570);
or UO_325 (O_325,N_2339,N_2878);
nand UO_326 (O_326,N_2464,N_2701);
or UO_327 (O_327,N_2928,N_2906);
xor UO_328 (O_328,N_2813,N_2162);
nand UO_329 (O_329,N_2215,N_2197);
and UO_330 (O_330,N_2468,N_2246);
and UO_331 (O_331,N_2270,N_2367);
and UO_332 (O_332,N_2133,N_2436);
nand UO_333 (O_333,N_2085,N_2638);
nand UO_334 (O_334,N_2919,N_2346);
and UO_335 (O_335,N_2334,N_2849);
or UO_336 (O_336,N_2396,N_2827);
xnor UO_337 (O_337,N_2615,N_2084);
nor UO_338 (O_338,N_2842,N_2646);
nand UO_339 (O_339,N_2871,N_2050);
nor UO_340 (O_340,N_2718,N_2726);
or UO_341 (O_341,N_2837,N_2732);
or UO_342 (O_342,N_2455,N_2427);
and UO_343 (O_343,N_2264,N_2950);
nand UO_344 (O_344,N_2748,N_2762);
nand UO_345 (O_345,N_2253,N_2844);
nor UO_346 (O_346,N_2278,N_2763);
or UO_347 (O_347,N_2207,N_2778);
nand UO_348 (O_348,N_2152,N_2891);
nand UO_349 (O_349,N_2965,N_2073);
nand UO_350 (O_350,N_2401,N_2158);
and UO_351 (O_351,N_2358,N_2074);
nor UO_352 (O_352,N_2833,N_2566);
or UO_353 (O_353,N_2934,N_2619);
nor UO_354 (O_354,N_2976,N_2171);
or UO_355 (O_355,N_2043,N_2676);
nor UO_356 (O_356,N_2262,N_2750);
and UO_357 (O_357,N_2299,N_2775);
or UO_358 (O_358,N_2824,N_2946);
or UO_359 (O_359,N_2663,N_2686);
nand UO_360 (O_360,N_2675,N_2509);
nor UO_361 (O_361,N_2910,N_2440);
or UO_362 (O_362,N_2851,N_2355);
xor UO_363 (O_363,N_2114,N_2519);
nor UO_364 (O_364,N_2106,N_2580);
or UO_365 (O_365,N_2852,N_2122);
nor UO_366 (O_366,N_2448,N_2791);
nor UO_367 (O_367,N_2649,N_2029);
or UO_368 (O_368,N_2083,N_2282);
nor UO_369 (O_369,N_2783,N_2557);
or UO_370 (O_370,N_2923,N_2561);
nand UO_371 (O_371,N_2348,N_2680);
and UO_372 (O_372,N_2458,N_2988);
or UO_373 (O_373,N_2628,N_2196);
nand UO_374 (O_374,N_2416,N_2057);
nor UO_375 (O_375,N_2120,N_2179);
or UO_376 (O_376,N_2504,N_2379);
nand UO_377 (O_377,N_2908,N_2708);
or UO_378 (O_378,N_2486,N_2224);
and UO_379 (O_379,N_2161,N_2715);
nand UO_380 (O_380,N_2870,N_2961);
and UO_381 (O_381,N_2323,N_2985);
nand UO_382 (O_382,N_2859,N_2476);
or UO_383 (O_383,N_2793,N_2592);
nand UO_384 (O_384,N_2220,N_2431);
or UO_385 (O_385,N_2181,N_2463);
or UO_386 (O_386,N_2294,N_2061);
nand UO_387 (O_387,N_2483,N_2689);
or UO_388 (O_388,N_2434,N_2794);
or UO_389 (O_389,N_2795,N_2831);
xnor UO_390 (O_390,N_2819,N_2713);
nor UO_391 (O_391,N_2830,N_2188);
nor UO_392 (O_392,N_2678,N_2558);
and UO_393 (O_393,N_2935,N_2002);
and UO_394 (O_394,N_2076,N_2958);
nor UO_395 (O_395,N_2045,N_2587);
xor UO_396 (O_396,N_2818,N_2402);
nor UO_397 (O_397,N_2375,N_2012);
or UO_398 (O_398,N_2324,N_2450);
and UO_399 (O_399,N_2211,N_2041);
or UO_400 (O_400,N_2634,N_2330);
and UO_401 (O_401,N_2308,N_2531);
nor UO_402 (O_402,N_2444,N_2549);
or UO_403 (O_403,N_2834,N_2318);
nor UO_404 (O_404,N_2420,N_2698);
or UO_405 (O_405,N_2202,N_2186);
nand UO_406 (O_406,N_2679,N_2135);
or UO_407 (O_407,N_2310,N_2828);
nor UO_408 (O_408,N_2154,N_2115);
or UO_409 (O_409,N_2520,N_2382);
xor UO_410 (O_410,N_2266,N_2596);
nor UO_411 (O_411,N_2489,N_2297);
or UO_412 (O_412,N_2363,N_2315);
nor UO_413 (O_413,N_2376,N_2942);
nor UO_414 (O_414,N_2508,N_2048);
nor UO_415 (O_415,N_2221,N_2968);
and UO_416 (O_416,N_2792,N_2712);
or UO_417 (O_417,N_2260,N_2565);
nor UO_418 (O_418,N_2639,N_2227);
and UO_419 (O_419,N_2618,N_2536);
nand UO_420 (O_420,N_2736,N_2670);
and UO_421 (O_421,N_2657,N_2896);
nand UO_422 (O_422,N_2200,N_2979);
nand UO_423 (O_423,N_2095,N_2411);
nand UO_424 (O_424,N_2505,N_2936);
or UO_425 (O_425,N_2306,N_2660);
or UO_426 (O_426,N_2407,N_2892);
or UO_427 (O_427,N_2169,N_2863);
and UO_428 (O_428,N_2609,N_2997);
or UO_429 (O_429,N_2502,N_2812);
or UO_430 (O_430,N_2516,N_2301);
and UO_431 (O_431,N_2506,N_2719);
xor UO_432 (O_432,N_2467,N_2273);
and UO_433 (O_433,N_2218,N_2650);
xor UO_434 (O_434,N_2170,N_2640);
nand UO_435 (O_435,N_2304,N_2581);
or UO_436 (O_436,N_2893,N_2209);
nor UO_437 (O_437,N_2799,N_2125);
and UO_438 (O_438,N_2139,N_2009);
or UO_439 (O_439,N_2706,N_2918);
and UO_440 (O_440,N_2692,N_2130);
and UO_441 (O_441,N_2599,N_2677);
nand UO_442 (O_442,N_2077,N_2724);
nor UO_443 (O_443,N_2228,N_2801);
xnor UO_444 (O_444,N_2973,N_2490);
or UO_445 (O_445,N_2291,N_2441);
nand UO_446 (O_446,N_2603,N_2465);
nor UO_447 (O_447,N_2832,N_2063);
and UO_448 (O_448,N_2102,N_2208);
or UO_449 (O_449,N_2229,N_2978);
nand UO_450 (O_450,N_2344,N_2010);
and UO_451 (O_451,N_2866,N_2949);
nor UO_452 (O_452,N_2206,N_2374);
and UO_453 (O_453,N_2929,N_2856);
xor UO_454 (O_454,N_2875,N_2941);
or UO_455 (O_455,N_2846,N_2858);
and UO_456 (O_456,N_2190,N_2931);
and UO_457 (O_457,N_2105,N_2365);
and UO_458 (O_458,N_2539,N_2755);
or UO_459 (O_459,N_2840,N_2784);
xnor UO_460 (O_460,N_2574,N_2653);
nor UO_461 (O_461,N_2917,N_2466);
nand UO_462 (O_462,N_2479,N_2617);
or UO_463 (O_463,N_2150,N_2020);
nor UO_464 (O_464,N_2876,N_2430);
or UO_465 (O_465,N_2071,N_2904);
nor UO_466 (O_466,N_2770,N_2980);
xnor UO_467 (O_467,N_2568,N_2199);
and UO_468 (O_468,N_2843,N_2478);
nor UO_469 (O_469,N_2733,N_2290);
nor UO_470 (O_470,N_2926,N_2347);
nand UO_471 (O_471,N_2086,N_2316);
or UO_472 (O_472,N_2500,N_2809);
or UO_473 (O_473,N_2275,N_2737);
nand UO_474 (O_474,N_2764,N_2345);
nor UO_475 (O_475,N_2438,N_2066);
nor UO_476 (O_476,N_2212,N_2176);
and UO_477 (O_477,N_2494,N_2591);
nand UO_478 (O_478,N_2957,N_2598);
or UO_479 (O_479,N_2885,N_2760);
xor UO_480 (O_480,N_2517,N_2213);
nor UO_481 (O_481,N_2642,N_2243);
xnor UO_482 (O_482,N_2461,N_2960);
and UO_483 (O_483,N_2024,N_2474);
and UO_484 (O_484,N_2038,N_2322);
and UO_485 (O_485,N_2432,N_2248);
xor UO_486 (O_486,N_2252,N_2682);
or UO_487 (O_487,N_2668,N_2113);
or UO_488 (O_488,N_2433,N_2644);
nand UO_489 (O_489,N_2687,N_2094);
or UO_490 (O_490,N_2134,N_2237);
nand UO_491 (O_491,N_2142,N_2754);
and UO_492 (O_492,N_2000,N_2320);
nor UO_493 (O_493,N_2989,N_2384);
nor UO_494 (O_494,N_2001,N_2092);
and UO_495 (O_495,N_2204,N_2835);
nand UO_496 (O_496,N_2555,N_2477);
nor UO_497 (O_497,N_2710,N_2922);
nor UO_498 (O_498,N_2356,N_2058);
or UO_499 (O_499,N_2485,N_2877);
endmodule