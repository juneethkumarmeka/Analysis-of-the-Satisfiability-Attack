module basic_1000_10000_1500_20_levels_10xor_4(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999;
and U0 (N_0,In_861,In_795);
xor U1 (N_1,In_476,In_460);
and U2 (N_2,In_183,In_105);
or U3 (N_3,In_671,In_805);
nand U4 (N_4,In_243,In_283);
or U5 (N_5,In_330,In_164);
nand U6 (N_6,In_650,In_22);
nand U7 (N_7,In_894,In_913);
nor U8 (N_8,In_548,In_579);
nand U9 (N_9,In_191,In_961);
nor U10 (N_10,In_386,In_552);
nand U11 (N_11,In_29,In_714);
and U12 (N_12,In_116,In_748);
nand U13 (N_13,In_610,In_702);
nand U14 (N_14,In_238,In_37);
or U15 (N_15,In_735,In_267);
or U16 (N_16,In_663,In_690);
nand U17 (N_17,In_763,In_766);
nor U18 (N_18,In_721,In_398);
or U19 (N_19,In_176,In_237);
nor U20 (N_20,In_455,In_179);
xnor U21 (N_21,In_305,In_727);
nor U22 (N_22,In_965,In_438);
nand U23 (N_23,In_377,In_51);
and U24 (N_24,In_797,In_4);
nor U25 (N_25,In_102,In_551);
and U26 (N_26,In_391,In_198);
nand U27 (N_27,In_863,In_24);
or U28 (N_28,In_138,In_311);
nand U29 (N_29,In_847,In_917);
nor U30 (N_30,In_118,In_877);
nand U31 (N_31,In_645,In_779);
nand U32 (N_32,In_354,In_905);
nand U33 (N_33,In_173,In_434);
and U34 (N_34,In_636,In_891);
nor U35 (N_35,In_637,In_49);
nand U36 (N_36,In_135,In_812);
nor U37 (N_37,In_294,In_565);
and U38 (N_38,In_194,In_472);
or U39 (N_39,In_413,In_292);
xnor U40 (N_40,In_642,In_293);
xnor U41 (N_41,In_152,In_127);
xnor U42 (N_42,In_655,In_181);
xor U43 (N_43,In_34,In_31);
nor U44 (N_44,In_983,In_373);
or U45 (N_45,In_252,In_653);
nand U46 (N_46,In_800,In_33);
or U47 (N_47,In_555,In_9);
nand U48 (N_48,In_502,In_92);
nand U49 (N_49,In_69,In_833);
or U50 (N_50,In_55,In_215);
nor U51 (N_51,In_487,In_226);
xor U52 (N_52,In_785,In_873);
xnor U53 (N_53,In_932,In_190);
or U54 (N_54,In_395,In_617);
and U55 (N_55,In_47,In_389);
or U56 (N_56,In_924,In_83);
or U57 (N_57,In_420,In_910);
xor U58 (N_58,In_374,In_335);
and U59 (N_59,In_436,In_888);
nand U60 (N_60,In_204,In_717);
and U61 (N_61,In_115,In_951);
nand U62 (N_62,In_208,In_949);
or U63 (N_63,In_449,In_38);
and U64 (N_64,In_558,In_236);
xnor U65 (N_65,In_782,In_819);
xnor U66 (N_66,In_783,In_295);
nand U67 (N_67,In_255,In_985);
and U68 (N_68,In_998,In_734);
xnor U69 (N_69,In_43,In_697);
nand U70 (N_70,In_789,In_367);
nand U71 (N_71,In_578,In_214);
nand U72 (N_72,In_784,In_160);
or U73 (N_73,In_402,In_992);
xor U74 (N_74,In_131,In_856);
and U75 (N_75,In_545,In_950);
or U76 (N_76,In_284,In_750);
xor U77 (N_77,In_537,In_874);
nor U78 (N_78,In_633,In_234);
and U79 (N_79,In_987,In_870);
nand U80 (N_80,In_346,In_62);
nor U81 (N_81,In_385,In_189);
xor U82 (N_82,In_241,In_435);
nand U83 (N_83,In_375,In_796);
or U84 (N_84,In_128,In_549);
nor U85 (N_85,In_353,In_248);
nand U86 (N_86,In_712,In_614);
or U87 (N_87,In_749,In_121);
xnor U88 (N_88,In_600,In_976);
nand U89 (N_89,In_348,In_729);
or U90 (N_90,In_103,In_325);
nand U91 (N_91,In_569,In_20);
and U92 (N_92,In_495,In_494);
and U93 (N_93,In_559,In_948);
nand U94 (N_94,In_590,In_58);
and U95 (N_95,In_538,In_516);
nand U96 (N_96,In_475,In_153);
and U97 (N_97,In_981,In_591);
and U98 (N_98,In_492,In_171);
nand U99 (N_99,In_309,In_188);
xnor U100 (N_100,In_711,In_817);
or U101 (N_101,In_986,In_124);
or U102 (N_102,In_718,In_521);
xnor U103 (N_103,In_908,In_822);
xor U104 (N_104,In_67,In_527);
and U105 (N_105,In_867,In_461);
or U106 (N_106,In_601,In_792);
nand U107 (N_107,In_694,In_358);
xnor U108 (N_108,In_428,In_235);
nand U109 (N_109,In_496,In_895);
xor U110 (N_110,In_658,In_846);
xnor U111 (N_111,In_919,In_68);
and U112 (N_112,In_643,In_915);
or U113 (N_113,In_363,In_64);
nand U114 (N_114,In_211,In_753);
nor U115 (N_115,In_979,In_141);
nand U116 (N_116,In_927,In_786);
and U117 (N_117,In_306,In_553);
or U118 (N_118,In_710,In_627);
or U119 (N_119,In_594,In_321);
nand U120 (N_120,In_533,In_666);
nand U121 (N_121,In_145,In_299);
or U122 (N_122,In_76,In_317);
or U123 (N_123,In_78,In_212);
and U124 (N_124,In_519,In_349);
nand U125 (N_125,In_225,In_341);
or U126 (N_126,In_931,In_599);
nor U127 (N_127,In_644,In_376);
xor U128 (N_128,In_430,In_952);
or U129 (N_129,In_380,In_586);
or U130 (N_130,In_577,In_607);
or U131 (N_131,In_126,In_246);
xor U132 (N_132,In_480,In_256);
nor U133 (N_133,In_878,In_946);
nor U134 (N_134,In_746,In_427);
nand U135 (N_135,In_429,In_865);
or U136 (N_136,In_674,In_387);
xnor U137 (N_137,In_889,In_447);
nand U138 (N_138,In_532,In_875);
nand U139 (N_139,In_770,In_206);
nand U140 (N_140,In_597,In_265);
xor U141 (N_141,In_871,In_254);
and U142 (N_142,In_862,In_724);
nand U143 (N_143,In_356,In_0);
and U144 (N_144,In_576,In_524);
and U145 (N_145,In_806,In_28);
or U146 (N_146,In_593,In_409);
nand U147 (N_147,In_901,In_32);
nor U148 (N_148,In_980,In_818);
nand U149 (N_149,In_955,In_612);
nand U150 (N_150,In_540,In_315);
and U151 (N_151,In_960,In_944);
xnor U152 (N_152,In_972,In_692);
xor U153 (N_153,In_771,In_454);
xor U154 (N_154,In_536,In_168);
nand U155 (N_155,In_247,In_570);
xnor U156 (N_156,In_675,In_106);
nor U157 (N_157,In_827,In_896);
nand U158 (N_158,In_403,In_323);
or U159 (N_159,In_903,In_898);
nand U160 (N_160,In_959,In_744);
or U161 (N_161,In_529,In_77);
and U162 (N_162,In_528,In_759);
or U163 (N_163,In_186,In_40);
or U164 (N_164,In_362,In_157);
nand U165 (N_165,In_816,In_334);
nand U166 (N_166,In_379,In_406);
nand U167 (N_167,In_720,In_573);
and U168 (N_168,In_661,In_942);
and U169 (N_169,In_921,In_57);
or U170 (N_170,In_835,In_479);
and U171 (N_171,In_703,In_146);
nand U172 (N_172,In_444,In_707);
xor U173 (N_173,In_508,In_264);
and U174 (N_174,In_592,In_556);
and U175 (N_175,In_125,In_332);
xor U176 (N_176,In_880,In_338);
and U177 (N_177,In_716,In_88);
nand U178 (N_178,In_513,In_995);
or U179 (N_179,In_359,In_365);
nand U180 (N_180,In_589,In_90);
and U181 (N_181,In_336,In_500);
or U182 (N_182,In_313,In_993);
xor U183 (N_183,In_240,In_139);
and U184 (N_184,In_518,In_974);
and U185 (N_185,In_756,In_631);
xnor U186 (N_186,In_81,In_616);
or U187 (N_187,In_504,In_776);
nand U188 (N_188,In_858,In_497);
and U189 (N_189,In_218,In_651);
nor U190 (N_190,In_144,In_531);
xnor U191 (N_191,In_273,In_799);
and U192 (N_192,In_301,In_114);
xnor U193 (N_193,In_344,In_973);
nor U194 (N_194,In_509,In_935);
and U195 (N_195,In_854,In_688);
xor U196 (N_196,In_456,In_693);
nand U197 (N_197,In_488,In_250);
and U198 (N_198,In_625,In_458);
nand U199 (N_199,In_794,In_154);
xnor U200 (N_200,In_638,In_731);
xor U201 (N_201,In_316,In_91);
or U202 (N_202,In_30,In_314);
nor U203 (N_203,In_418,In_280);
nand U204 (N_204,In_737,In_382);
nor U205 (N_205,In_680,In_978);
xor U206 (N_206,In_649,In_408);
xnor U207 (N_207,In_535,In_485);
nor U208 (N_208,In_452,In_44);
and U209 (N_209,In_904,In_12);
xor U210 (N_210,In_469,In_684);
or U211 (N_211,In_676,In_654);
or U212 (N_212,In_407,In_704);
and U213 (N_213,In_61,In_249);
and U214 (N_214,In_290,In_554);
or U215 (N_215,In_813,In_665);
xor U216 (N_216,In_659,In_459);
xnor U217 (N_217,In_575,In_130);
nor U218 (N_218,In_132,In_587);
or U219 (N_219,In_6,In_802);
xor U220 (N_220,In_259,In_270);
or U221 (N_221,In_768,In_681);
nand U222 (N_222,In_715,In_804);
xor U223 (N_223,In_210,In_21);
nand U224 (N_224,In_137,In_165);
nor U225 (N_225,In_677,In_393);
nor U226 (N_226,In_736,In_886);
or U227 (N_227,In_517,In_953);
nand U228 (N_228,In_611,In_343);
and U229 (N_229,In_312,In_87);
or U230 (N_230,In_79,In_129);
and U231 (N_231,In_624,In_491);
and U232 (N_232,In_852,In_885);
and U233 (N_233,In_933,In_708);
nor U234 (N_234,In_791,In_123);
nand U235 (N_235,In_781,In_689);
and U236 (N_236,In_269,In_468);
nand U237 (N_237,In_371,In_635);
xor U238 (N_238,In_390,In_628);
nor U239 (N_239,In_902,In_941);
or U240 (N_240,In_322,In_392);
nor U241 (N_241,In_222,In_357);
nor U242 (N_242,In_840,In_440);
and U243 (N_243,In_80,In_988);
xor U244 (N_244,In_738,In_629);
nand U245 (N_245,In_831,In_997);
nor U246 (N_246,In_775,In_178);
or U247 (N_247,In_872,In_845);
nor U248 (N_248,In_741,In_542);
nand U249 (N_249,In_962,In_672);
nor U250 (N_250,In_945,In_347);
nand U251 (N_251,In_414,In_448);
xnor U252 (N_252,In_760,In_85);
nand U253 (N_253,In_350,In_368);
or U254 (N_254,In_41,In_372);
nand U255 (N_255,In_740,In_467);
and U256 (N_256,In_630,In_483);
and U257 (N_257,In_268,In_745);
nand U258 (N_258,In_899,In_975);
nand U259 (N_259,In_310,In_523);
nor U260 (N_260,In_482,In_388);
or U261 (N_261,In_272,In_303);
nor U262 (N_262,In_39,In_148);
or U263 (N_263,In_842,In_260);
and U264 (N_264,In_939,In_698);
and U265 (N_265,In_887,In_892);
or U266 (N_266,In_820,In_620);
nand U267 (N_267,In_404,In_54);
and U268 (N_268,In_405,In_982);
nor U269 (N_269,In_163,In_275);
and U270 (N_270,In_696,In_10);
xnor U271 (N_271,In_477,In_583);
and U272 (N_272,In_767,In_286);
nand U273 (N_273,In_251,In_754);
nor U274 (N_274,In_808,In_977);
nor U275 (N_275,In_568,In_825);
and U276 (N_276,In_327,In_177);
xnor U277 (N_277,In_296,In_691);
nor U278 (N_278,In_522,In_287);
nand U279 (N_279,In_732,In_656);
or U280 (N_280,In_828,In_113);
nor U281 (N_281,In_954,In_462);
nand U282 (N_282,In_416,In_169);
and U283 (N_283,In_196,In_761);
xnor U284 (N_284,In_23,In_70);
xor U285 (N_285,In_897,In_324);
or U286 (N_286,In_423,In_826);
xor U287 (N_287,In_490,In_74);
xor U288 (N_288,In_743,In_911);
or U289 (N_289,In_928,In_832);
xor U290 (N_290,In_857,In_86);
nor U291 (N_291,In_850,In_200);
and U292 (N_292,In_120,In_401);
nor U293 (N_293,In_209,In_709);
nand U294 (N_294,In_733,In_197);
and U295 (N_295,In_907,In_231);
nor U296 (N_296,In_790,In_450);
and U297 (N_297,In_229,In_442);
xor U298 (N_298,In_220,In_342);
xnor U299 (N_299,In_758,In_969);
nor U300 (N_300,In_415,In_580);
nor U301 (N_301,In_609,In_967);
nor U302 (N_302,In_788,In_605);
and U303 (N_303,In_426,In_397);
nor U304 (N_304,In_958,In_89);
xnor U305 (N_305,In_506,In_337);
and U306 (N_306,In_158,In_167);
or U307 (N_307,In_446,In_308);
xor U308 (N_308,In_909,In_999);
or U309 (N_309,In_984,In_632);
or U310 (N_310,In_780,In_17);
nand U311 (N_311,In_762,In_96);
nand U312 (N_312,In_394,In_673);
nor U313 (N_313,In_662,In_352);
and U314 (N_314,In_968,In_101);
nor U315 (N_315,In_505,In_384);
or U316 (N_316,In_574,In_439);
or U317 (N_317,In_608,In_747);
nor U318 (N_318,In_134,In_13);
nand U319 (N_319,In_615,In_203);
or U320 (N_320,In_765,In_934);
or U321 (N_321,In_544,In_278);
xor U322 (N_322,In_550,In_63);
nand U323 (N_323,In_400,In_360);
nor U324 (N_324,In_36,In_59);
or U325 (N_325,In_72,In_53);
nand U326 (N_326,In_572,In_670);
or U327 (N_327,In_228,In_166);
xnor U328 (N_328,In_929,In_143);
xnor U329 (N_329,In_445,In_192);
and U330 (N_330,In_7,In_291);
nor U331 (N_331,In_956,In_668);
nand U332 (N_332,In_752,In_457);
and U333 (N_333,In_253,In_772);
xor U334 (N_334,In_882,In_258);
and U335 (N_335,In_742,In_498);
xnor U336 (N_336,In_626,In_331);
nor U337 (N_337,In_814,In_227);
xor U338 (N_338,In_302,In_660);
or U339 (N_339,In_262,In_232);
nand U340 (N_340,In_151,In_507);
nand U341 (N_341,In_739,In_890);
xor U342 (N_342,In_162,In_701);
nor U343 (N_343,In_15,In_602);
xor U344 (N_344,In_562,In_937);
nor U345 (N_345,In_868,In_184);
or U346 (N_346,In_111,In_582);
or U347 (N_347,In_318,In_824);
nand U348 (N_348,In_340,In_117);
and U349 (N_349,In_839,In_722);
or U350 (N_350,In_396,In_94);
nand U351 (N_351,In_122,In_351);
xor U352 (N_352,In_99,In_185);
nand U353 (N_353,In_838,In_851);
xnor U354 (N_354,In_581,In_412);
or U355 (N_355,In_464,In_916);
nor U356 (N_356,In_48,In_369);
nor U357 (N_357,In_26,In_652);
nor U358 (N_358,In_297,In_634);
nand U359 (N_359,In_841,In_478);
nand U360 (N_360,In_514,In_474);
or U361 (N_361,In_725,In_433);
nand U362 (N_362,In_465,In_530);
xor U363 (N_363,In_619,In_217);
nor U364 (N_364,In_180,In_424);
nand U365 (N_365,In_432,In_525);
and U366 (N_366,In_855,In_526);
and U367 (N_367,In_304,In_864);
or U368 (N_368,In_65,In_906);
or U369 (N_369,In_773,In_471);
nand U370 (N_370,In_859,In_618);
or U371 (N_371,In_104,In_245);
and U372 (N_372,In_383,In_19);
xor U373 (N_373,In_991,In_571);
xor U374 (N_374,In_46,In_281);
nand U375 (N_375,In_35,In_27);
and U376 (N_376,In_947,In_584);
or U377 (N_377,In_489,In_811);
nor U378 (N_378,In_561,In_473);
and U379 (N_379,In_511,In_261);
or U380 (N_380,In_604,In_75);
xnor U381 (N_381,In_142,In_966);
nand U382 (N_382,In_830,In_809);
nand U383 (N_383,In_606,In_879);
nand U384 (N_384,In_801,In_437);
or U385 (N_385,In_567,In_914);
nand U386 (N_386,In_98,In_174);
or U387 (N_387,In_66,In_499);
nand U388 (N_388,In_940,In_774);
and U389 (N_389,In_453,In_5);
and U390 (N_390,In_205,In_598);
xor U391 (N_391,In_187,In_541);
and U392 (N_392,In_853,In_682);
and U393 (N_393,In_777,In_520);
or U394 (N_394,In_943,In_257);
or U395 (N_395,In_501,In_370);
xor U396 (N_396,In_639,In_989);
or U397 (N_397,In_133,In_920);
and U398 (N_398,In_695,In_207);
and U399 (N_399,In_560,In_699);
nand U400 (N_400,In_274,In_421);
or U401 (N_401,In_289,In_730);
nor U402 (N_402,In_221,In_244);
nor U403 (N_403,In_849,In_441);
nand U404 (N_404,In_679,In_647);
or U405 (N_405,In_155,In_723);
or U406 (N_406,In_893,In_233);
or U407 (N_407,In_787,In_71);
xnor U408 (N_408,In_829,In_112);
nand U409 (N_409,In_149,In_484);
nand U410 (N_410,In_93,In_378);
or U411 (N_411,In_613,In_82);
xor U412 (N_412,In_843,In_361);
xor U413 (N_413,In_300,In_18);
or U414 (N_414,In_345,In_242);
nand U415 (N_415,In_411,In_685);
nand U416 (N_416,In_60,In_224);
xnor U417 (N_417,In_109,In_900);
and U418 (N_418,In_486,In_669);
or U419 (N_419,In_640,In_687);
nand U420 (N_420,In_172,In_778);
or U421 (N_421,In_883,In_73);
and U422 (N_422,In_751,In_288);
xor U423 (N_423,In_664,In_451);
and U424 (N_424,In_239,In_564);
xor U425 (N_425,In_333,In_100);
nand U426 (N_426,In_970,In_648);
nor U427 (N_427,In_990,In_355);
nor U428 (N_428,In_912,In_821);
nand U429 (N_429,In_667,In_657);
or U430 (N_430,In_547,In_266);
or U431 (N_431,In_534,In_866);
nor U432 (N_432,In_971,In_175);
nand U433 (N_433,In_503,In_326);
nor U434 (N_434,In_603,In_3);
and U435 (N_435,In_147,In_938);
nand U436 (N_436,In_140,In_546);
and U437 (N_437,In_276,In_84);
or U438 (N_438,In_282,In_470);
nor U439 (N_439,In_622,In_156);
nand U440 (N_440,In_159,In_621);
xor U441 (N_441,In_881,In_339);
and U442 (N_442,In_646,In_431);
nor U443 (N_443,In_56,In_623);
or U444 (N_444,In_161,In_182);
and U445 (N_445,In_810,In_277);
nor U446 (N_446,In_419,In_11);
nand U447 (N_447,In_199,In_563);
xnor U448 (N_448,In_320,In_755);
nand U449 (N_449,In_807,In_25);
nand U450 (N_450,In_193,In_836);
xnor U451 (N_451,In_463,In_793);
or U452 (N_452,In_764,In_923);
nor U453 (N_453,In_757,In_996);
nor U454 (N_454,In_719,In_493);
nor U455 (N_455,In_42,In_700);
nand U456 (N_456,In_769,In_466);
nor U457 (N_457,In_641,In_678);
xor U458 (N_458,In_515,In_230);
nand U459 (N_459,In_512,In_848);
nor U460 (N_460,In_136,In_263);
and U461 (N_461,In_957,In_922);
or U462 (N_462,In_686,In_45);
or U463 (N_463,In_195,In_319);
nand U464 (N_464,In_728,In_285);
and U465 (N_465,In_417,In_844);
nand U466 (N_466,In_97,In_963);
xor U467 (N_467,In_860,In_834);
and U468 (N_468,In_713,In_328);
nor U469 (N_469,In_52,In_837);
nor U470 (N_470,In_50,In_994);
nand U471 (N_471,In_298,In_223);
nor U472 (N_472,In_2,In_307);
nand U473 (N_473,In_399,In_595);
nor U474 (N_474,In_925,In_279);
nand U475 (N_475,In_119,In_930);
and U476 (N_476,In_588,In_683);
or U477 (N_477,In_705,In_481);
nand U478 (N_478,In_110,In_107);
xnor U479 (N_479,In_726,In_557);
nand U480 (N_480,In_706,In_16);
or U481 (N_481,In_815,In_539);
or U482 (N_482,In_443,In_150);
nor U483 (N_483,In_1,In_964);
and U484 (N_484,In_596,In_219);
or U485 (N_485,In_803,In_936);
or U486 (N_486,In_95,In_381);
or U487 (N_487,In_170,In_202);
nand U488 (N_488,In_271,In_329);
or U489 (N_489,In_422,In_926);
or U490 (N_490,In_366,In_869);
xnor U491 (N_491,In_213,In_216);
nor U492 (N_492,In_884,In_823);
and U493 (N_493,In_364,In_410);
nor U494 (N_494,In_425,In_876);
or U495 (N_495,In_510,In_918);
xor U496 (N_496,In_201,In_8);
or U497 (N_497,In_14,In_566);
nor U498 (N_498,In_585,In_798);
nand U499 (N_499,In_543,In_108);
nand U500 (N_500,N_130,N_288);
nand U501 (N_501,N_150,N_100);
nand U502 (N_502,N_359,N_197);
nand U503 (N_503,N_117,N_131);
or U504 (N_504,N_142,N_394);
or U505 (N_505,N_86,N_302);
nor U506 (N_506,N_367,N_257);
nand U507 (N_507,N_106,N_23);
nor U508 (N_508,N_355,N_442);
or U509 (N_509,N_183,N_304);
nor U510 (N_510,N_72,N_381);
nand U511 (N_511,N_167,N_346);
xnor U512 (N_512,N_42,N_209);
or U513 (N_513,N_264,N_454);
or U514 (N_514,N_126,N_401);
and U515 (N_515,N_472,N_398);
nand U516 (N_516,N_119,N_17);
nor U517 (N_517,N_203,N_93);
or U518 (N_518,N_2,N_434);
nand U519 (N_519,N_275,N_244);
and U520 (N_520,N_323,N_411);
and U521 (N_521,N_189,N_280);
xnor U522 (N_522,N_110,N_213);
nand U523 (N_523,N_137,N_307);
xor U524 (N_524,N_335,N_347);
and U525 (N_525,N_223,N_153);
nor U526 (N_526,N_166,N_349);
nor U527 (N_527,N_8,N_309);
xnor U528 (N_528,N_39,N_241);
nand U529 (N_529,N_299,N_460);
nand U530 (N_530,N_206,N_435);
xnor U531 (N_531,N_64,N_360);
nand U532 (N_532,N_320,N_218);
and U533 (N_533,N_379,N_68);
nand U534 (N_534,N_370,N_92);
and U535 (N_535,N_227,N_295);
or U536 (N_536,N_80,N_459);
xor U537 (N_537,N_172,N_176);
xor U538 (N_538,N_233,N_1);
nand U539 (N_539,N_29,N_350);
or U540 (N_540,N_195,N_65);
nor U541 (N_541,N_371,N_466);
nor U542 (N_542,N_276,N_177);
xor U543 (N_543,N_416,N_333);
xnor U544 (N_544,N_358,N_98);
and U545 (N_545,N_338,N_208);
xnor U546 (N_546,N_62,N_180);
or U547 (N_547,N_268,N_407);
or U548 (N_548,N_105,N_285);
nor U549 (N_549,N_271,N_99);
or U550 (N_550,N_238,N_441);
or U551 (N_551,N_373,N_497);
and U552 (N_552,N_90,N_240);
or U553 (N_553,N_365,N_476);
and U554 (N_554,N_118,N_418);
nor U555 (N_555,N_449,N_192);
nand U556 (N_556,N_164,N_428);
xnor U557 (N_557,N_114,N_242);
nand U558 (N_558,N_159,N_0);
xor U559 (N_559,N_125,N_267);
nor U560 (N_560,N_111,N_327);
nor U561 (N_561,N_224,N_234);
or U562 (N_562,N_12,N_392);
nor U563 (N_563,N_190,N_79);
or U564 (N_564,N_220,N_406);
nand U565 (N_565,N_174,N_396);
and U566 (N_566,N_67,N_334);
xnor U567 (N_567,N_48,N_284);
and U568 (N_568,N_60,N_134);
xor U569 (N_569,N_246,N_112);
nand U570 (N_570,N_467,N_141);
nand U571 (N_571,N_361,N_71);
nor U572 (N_572,N_260,N_115);
nor U573 (N_573,N_91,N_292);
nor U574 (N_574,N_353,N_461);
nor U575 (N_575,N_188,N_127);
nand U576 (N_576,N_311,N_84);
and U577 (N_577,N_430,N_486);
xnor U578 (N_578,N_340,N_363);
xor U579 (N_579,N_279,N_265);
nand U580 (N_580,N_254,N_41);
and U581 (N_581,N_103,N_154);
nor U582 (N_582,N_54,N_322);
or U583 (N_583,N_456,N_423);
and U584 (N_584,N_161,N_287);
nand U585 (N_585,N_298,N_282);
xor U586 (N_586,N_286,N_377);
nand U587 (N_587,N_70,N_326);
or U588 (N_588,N_193,N_32);
xor U589 (N_589,N_354,N_494);
nor U590 (N_590,N_24,N_236);
nand U591 (N_591,N_222,N_149);
nand U592 (N_592,N_453,N_101);
nand U593 (N_593,N_471,N_255);
and U594 (N_594,N_290,N_132);
nor U595 (N_595,N_372,N_393);
or U596 (N_596,N_308,N_475);
and U597 (N_597,N_22,N_325);
and U598 (N_598,N_306,N_210);
nand U599 (N_599,N_412,N_13);
and U600 (N_600,N_336,N_4);
or U601 (N_601,N_452,N_305);
or U602 (N_602,N_49,N_143);
nor U603 (N_603,N_490,N_324);
or U604 (N_604,N_7,N_16);
xnor U605 (N_605,N_57,N_201);
nor U606 (N_606,N_185,N_191);
xnor U607 (N_607,N_107,N_179);
or U608 (N_608,N_215,N_169);
or U609 (N_609,N_439,N_249);
nor U610 (N_610,N_283,N_251);
or U611 (N_611,N_151,N_395);
nor U612 (N_612,N_481,N_463);
or U613 (N_613,N_138,N_165);
nor U614 (N_614,N_297,N_53);
nor U615 (N_615,N_319,N_207);
nor U616 (N_616,N_273,N_199);
xnor U617 (N_617,N_194,N_480);
or U618 (N_618,N_383,N_66);
or U619 (N_619,N_450,N_424);
and U620 (N_620,N_30,N_173);
nor U621 (N_621,N_455,N_216);
and U622 (N_622,N_278,N_313);
nand U623 (N_623,N_404,N_45);
or U624 (N_624,N_170,N_77);
or U625 (N_625,N_432,N_33);
xnor U626 (N_626,N_487,N_385);
xnor U627 (N_627,N_378,N_421);
and U628 (N_628,N_496,N_235);
xor U629 (N_629,N_274,N_163);
xnor U630 (N_630,N_196,N_139);
or U631 (N_631,N_499,N_51);
nand U632 (N_632,N_148,N_155);
and U633 (N_633,N_78,N_36);
nor U634 (N_634,N_56,N_146);
and U635 (N_635,N_321,N_205);
xor U636 (N_636,N_243,N_368);
or U637 (N_637,N_156,N_229);
and U638 (N_638,N_427,N_375);
or U639 (N_639,N_133,N_50);
and U640 (N_640,N_25,N_85);
xor U641 (N_641,N_226,N_330);
or U642 (N_642,N_414,N_436);
and U643 (N_643,N_269,N_468);
and U644 (N_644,N_303,N_145);
and U645 (N_645,N_409,N_492);
nor U646 (N_646,N_410,N_445);
nand U647 (N_647,N_178,N_369);
or U648 (N_648,N_47,N_277);
nand U649 (N_649,N_58,N_37);
nor U650 (N_650,N_113,N_458);
nor U651 (N_651,N_415,N_69);
nor U652 (N_652,N_237,N_120);
and U653 (N_653,N_217,N_382);
nand U654 (N_654,N_10,N_402);
nand U655 (N_655,N_491,N_75);
nor U656 (N_656,N_478,N_352);
and U657 (N_657,N_109,N_52);
nor U658 (N_658,N_437,N_187);
and U659 (N_659,N_87,N_348);
nand U660 (N_660,N_433,N_121);
xor U661 (N_661,N_477,N_19);
or U662 (N_662,N_211,N_102);
nor U663 (N_663,N_248,N_88);
nand U664 (N_664,N_293,N_26);
nor U665 (N_665,N_140,N_403);
nor U666 (N_666,N_444,N_417);
and U667 (N_667,N_200,N_182);
nand U668 (N_668,N_11,N_160);
or U669 (N_669,N_252,N_397);
nand U670 (N_670,N_429,N_81);
and U671 (N_671,N_270,N_144);
or U672 (N_672,N_400,N_342);
nor U673 (N_673,N_28,N_259);
xnor U674 (N_674,N_328,N_184);
nor U675 (N_675,N_446,N_6);
xnor U676 (N_676,N_89,N_440);
and U677 (N_677,N_46,N_55);
or U678 (N_678,N_135,N_204);
xor U679 (N_679,N_431,N_425);
and U680 (N_680,N_262,N_232);
xor U681 (N_681,N_95,N_221);
or U682 (N_682,N_74,N_63);
xor U683 (N_683,N_422,N_245);
nand U684 (N_684,N_380,N_408);
nor U685 (N_685,N_364,N_366);
and U686 (N_686,N_443,N_374);
or U687 (N_687,N_59,N_388);
xnor U688 (N_688,N_488,N_448);
xor U689 (N_689,N_464,N_43);
nand U690 (N_690,N_362,N_212);
nor U691 (N_691,N_314,N_474);
or U692 (N_692,N_76,N_301);
nand U693 (N_693,N_123,N_498);
nor U694 (N_694,N_136,N_317);
and U695 (N_695,N_399,N_186);
and U696 (N_696,N_484,N_250);
or U697 (N_697,N_289,N_129);
and U698 (N_698,N_152,N_14);
or U699 (N_699,N_258,N_413);
nor U700 (N_700,N_239,N_35);
nand U701 (N_701,N_344,N_219);
xor U702 (N_702,N_465,N_21);
nor U703 (N_703,N_479,N_281);
xor U704 (N_704,N_9,N_15);
or U705 (N_705,N_116,N_96);
xor U706 (N_706,N_339,N_108);
xnor U707 (N_707,N_473,N_389);
nor U708 (N_708,N_171,N_310);
and U709 (N_709,N_256,N_225);
nor U710 (N_710,N_261,N_20);
nand U711 (N_711,N_247,N_485);
or U712 (N_712,N_122,N_420);
and U713 (N_713,N_266,N_157);
nor U714 (N_714,N_202,N_40);
and U715 (N_715,N_272,N_5);
and U716 (N_716,N_341,N_356);
nand U717 (N_717,N_391,N_315);
nor U718 (N_718,N_316,N_214);
xor U719 (N_719,N_387,N_147);
and U720 (N_720,N_82,N_419);
nand U721 (N_721,N_44,N_168);
and U722 (N_722,N_104,N_253);
and U723 (N_723,N_61,N_128);
and U724 (N_724,N_489,N_34);
nand U725 (N_725,N_493,N_351);
xnor U726 (N_726,N_451,N_300);
and U727 (N_727,N_457,N_175);
and U728 (N_728,N_482,N_345);
nand U729 (N_729,N_230,N_462);
xor U730 (N_730,N_337,N_376);
xnor U731 (N_731,N_405,N_27);
nor U732 (N_732,N_483,N_198);
or U733 (N_733,N_83,N_331);
nor U734 (N_734,N_228,N_296);
nand U735 (N_735,N_469,N_73);
nand U736 (N_736,N_470,N_438);
nand U737 (N_737,N_386,N_231);
or U738 (N_738,N_312,N_94);
or U739 (N_739,N_357,N_3);
and U740 (N_740,N_181,N_291);
nor U741 (N_741,N_158,N_332);
and U742 (N_742,N_18,N_343);
xor U743 (N_743,N_447,N_263);
or U744 (N_744,N_426,N_329);
nand U745 (N_745,N_495,N_384);
nor U746 (N_746,N_162,N_97);
and U747 (N_747,N_38,N_294);
xnor U748 (N_748,N_390,N_31);
or U749 (N_749,N_318,N_124);
nor U750 (N_750,N_359,N_421);
and U751 (N_751,N_213,N_386);
nor U752 (N_752,N_278,N_489);
or U753 (N_753,N_341,N_102);
or U754 (N_754,N_110,N_324);
xnor U755 (N_755,N_8,N_375);
and U756 (N_756,N_346,N_255);
or U757 (N_757,N_90,N_5);
nor U758 (N_758,N_5,N_199);
xor U759 (N_759,N_358,N_398);
and U760 (N_760,N_373,N_296);
nand U761 (N_761,N_253,N_9);
nand U762 (N_762,N_187,N_367);
or U763 (N_763,N_189,N_248);
and U764 (N_764,N_254,N_274);
or U765 (N_765,N_130,N_230);
xor U766 (N_766,N_101,N_185);
or U767 (N_767,N_51,N_209);
and U768 (N_768,N_352,N_21);
and U769 (N_769,N_17,N_410);
and U770 (N_770,N_273,N_425);
or U771 (N_771,N_391,N_208);
or U772 (N_772,N_378,N_276);
or U773 (N_773,N_2,N_108);
or U774 (N_774,N_166,N_324);
or U775 (N_775,N_403,N_202);
xor U776 (N_776,N_201,N_457);
xnor U777 (N_777,N_477,N_297);
nor U778 (N_778,N_478,N_334);
xor U779 (N_779,N_273,N_398);
nor U780 (N_780,N_47,N_488);
nor U781 (N_781,N_10,N_90);
and U782 (N_782,N_296,N_65);
and U783 (N_783,N_156,N_452);
nand U784 (N_784,N_428,N_357);
nor U785 (N_785,N_76,N_44);
nor U786 (N_786,N_498,N_227);
or U787 (N_787,N_3,N_208);
xnor U788 (N_788,N_71,N_267);
xor U789 (N_789,N_237,N_482);
nor U790 (N_790,N_309,N_277);
nand U791 (N_791,N_212,N_39);
nor U792 (N_792,N_13,N_39);
nor U793 (N_793,N_414,N_201);
xor U794 (N_794,N_59,N_417);
nand U795 (N_795,N_193,N_476);
nand U796 (N_796,N_400,N_339);
and U797 (N_797,N_203,N_455);
xor U798 (N_798,N_477,N_401);
nand U799 (N_799,N_219,N_370);
xor U800 (N_800,N_50,N_148);
nand U801 (N_801,N_195,N_235);
or U802 (N_802,N_83,N_43);
and U803 (N_803,N_183,N_93);
and U804 (N_804,N_27,N_80);
and U805 (N_805,N_455,N_445);
xor U806 (N_806,N_467,N_416);
nand U807 (N_807,N_450,N_124);
xnor U808 (N_808,N_348,N_485);
nor U809 (N_809,N_83,N_283);
and U810 (N_810,N_21,N_374);
nor U811 (N_811,N_218,N_116);
or U812 (N_812,N_5,N_374);
and U813 (N_813,N_289,N_301);
nor U814 (N_814,N_309,N_209);
nor U815 (N_815,N_67,N_485);
and U816 (N_816,N_16,N_359);
xnor U817 (N_817,N_461,N_301);
nor U818 (N_818,N_433,N_66);
and U819 (N_819,N_160,N_259);
and U820 (N_820,N_446,N_198);
nand U821 (N_821,N_426,N_165);
or U822 (N_822,N_169,N_449);
nor U823 (N_823,N_203,N_343);
or U824 (N_824,N_404,N_459);
xor U825 (N_825,N_486,N_154);
and U826 (N_826,N_0,N_464);
xnor U827 (N_827,N_195,N_406);
or U828 (N_828,N_402,N_149);
xor U829 (N_829,N_58,N_104);
or U830 (N_830,N_382,N_365);
nand U831 (N_831,N_380,N_379);
and U832 (N_832,N_445,N_103);
nor U833 (N_833,N_489,N_235);
nor U834 (N_834,N_71,N_434);
and U835 (N_835,N_172,N_108);
or U836 (N_836,N_415,N_335);
xor U837 (N_837,N_74,N_496);
nor U838 (N_838,N_311,N_212);
nand U839 (N_839,N_114,N_59);
or U840 (N_840,N_455,N_268);
or U841 (N_841,N_496,N_165);
nand U842 (N_842,N_488,N_495);
and U843 (N_843,N_26,N_333);
nand U844 (N_844,N_219,N_338);
xnor U845 (N_845,N_21,N_347);
and U846 (N_846,N_160,N_452);
and U847 (N_847,N_487,N_337);
nor U848 (N_848,N_260,N_334);
nor U849 (N_849,N_55,N_287);
and U850 (N_850,N_447,N_375);
nand U851 (N_851,N_225,N_249);
nand U852 (N_852,N_189,N_148);
or U853 (N_853,N_283,N_188);
xor U854 (N_854,N_379,N_38);
nand U855 (N_855,N_459,N_490);
nand U856 (N_856,N_399,N_74);
or U857 (N_857,N_255,N_381);
nor U858 (N_858,N_150,N_52);
xor U859 (N_859,N_367,N_357);
nand U860 (N_860,N_157,N_418);
nor U861 (N_861,N_115,N_43);
and U862 (N_862,N_80,N_474);
and U863 (N_863,N_187,N_230);
nor U864 (N_864,N_132,N_378);
nand U865 (N_865,N_408,N_32);
xnor U866 (N_866,N_231,N_175);
nor U867 (N_867,N_179,N_177);
nand U868 (N_868,N_222,N_379);
nor U869 (N_869,N_88,N_326);
nand U870 (N_870,N_45,N_9);
nor U871 (N_871,N_8,N_72);
and U872 (N_872,N_28,N_212);
xnor U873 (N_873,N_427,N_22);
and U874 (N_874,N_407,N_178);
or U875 (N_875,N_247,N_442);
and U876 (N_876,N_225,N_236);
xor U877 (N_877,N_329,N_178);
xor U878 (N_878,N_292,N_177);
nand U879 (N_879,N_276,N_469);
or U880 (N_880,N_280,N_245);
or U881 (N_881,N_486,N_206);
and U882 (N_882,N_78,N_134);
nand U883 (N_883,N_194,N_104);
xnor U884 (N_884,N_186,N_439);
nor U885 (N_885,N_396,N_359);
xnor U886 (N_886,N_396,N_349);
and U887 (N_887,N_17,N_298);
xnor U888 (N_888,N_239,N_288);
or U889 (N_889,N_97,N_19);
and U890 (N_890,N_220,N_285);
nor U891 (N_891,N_455,N_466);
xnor U892 (N_892,N_413,N_380);
nor U893 (N_893,N_39,N_493);
nor U894 (N_894,N_262,N_33);
nor U895 (N_895,N_250,N_166);
nand U896 (N_896,N_251,N_397);
or U897 (N_897,N_370,N_56);
nor U898 (N_898,N_284,N_442);
xnor U899 (N_899,N_394,N_328);
and U900 (N_900,N_442,N_487);
nand U901 (N_901,N_61,N_316);
nand U902 (N_902,N_418,N_64);
nor U903 (N_903,N_404,N_452);
or U904 (N_904,N_436,N_82);
nor U905 (N_905,N_176,N_73);
or U906 (N_906,N_41,N_90);
or U907 (N_907,N_29,N_255);
and U908 (N_908,N_428,N_401);
xnor U909 (N_909,N_425,N_199);
nand U910 (N_910,N_349,N_194);
nor U911 (N_911,N_188,N_265);
nor U912 (N_912,N_103,N_330);
nand U913 (N_913,N_92,N_304);
nand U914 (N_914,N_271,N_165);
xnor U915 (N_915,N_57,N_119);
xor U916 (N_916,N_40,N_455);
nand U917 (N_917,N_162,N_384);
nand U918 (N_918,N_382,N_52);
xor U919 (N_919,N_93,N_254);
and U920 (N_920,N_194,N_206);
nand U921 (N_921,N_228,N_392);
and U922 (N_922,N_474,N_126);
xnor U923 (N_923,N_220,N_187);
and U924 (N_924,N_288,N_389);
or U925 (N_925,N_127,N_116);
nor U926 (N_926,N_451,N_385);
and U927 (N_927,N_443,N_491);
xnor U928 (N_928,N_116,N_12);
xor U929 (N_929,N_156,N_478);
nand U930 (N_930,N_97,N_281);
nand U931 (N_931,N_21,N_467);
nand U932 (N_932,N_154,N_303);
or U933 (N_933,N_50,N_340);
xnor U934 (N_934,N_189,N_312);
xnor U935 (N_935,N_354,N_15);
nand U936 (N_936,N_234,N_223);
or U937 (N_937,N_408,N_364);
xnor U938 (N_938,N_49,N_369);
or U939 (N_939,N_411,N_15);
and U940 (N_940,N_4,N_448);
or U941 (N_941,N_236,N_459);
and U942 (N_942,N_197,N_257);
nand U943 (N_943,N_303,N_164);
and U944 (N_944,N_194,N_190);
nor U945 (N_945,N_218,N_63);
nor U946 (N_946,N_224,N_29);
or U947 (N_947,N_377,N_457);
and U948 (N_948,N_231,N_163);
xor U949 (N_949,N_156,N_6);
nor U950 (N_950,N_262,N_149);
nor U951 (N_951,N_244,N_307);
xnor U952 (N_952,N_319,N_273);
or U953 (N_953,N_452,N_436);
nor U954 (N_954,N_218,N_495);
xor U955 (N_955,N_85,N_290);
nand U956 (N_956,N_387,N_404);
nor U957 (N_957,N_92,N_480);
or U958 (N_958,N_266,N_291);
xnor U959 (N_959,N_204,N_108);
nand U960 (N_960,N_65,N_337);
and U961 (N_961,N_56,N_451);
nand U962 (N_962,N_439,N_333);
nand U963 (N_963,N_449,N_280);
or U964 (N_964,N_18,N_425);
xor U965 (N_965,N_338,N_280);
or U966 (N_966,N_303,N_41);
nor U967 (N_967,N_392,N_104);
or U968 (N_968,N_435,N_459);
xnor U969 (N_969,N_109,N_461);
xor U970 (N_970,N_275,N_417);
xnor U971 (N_971,N_348,N_458);
nor U972 (N_972,N_341,N_274);
or U973 (N_973,N_55,N_406);
xor U974 (N_974,N_110,N_347);
or U975 (N_975,N_163,N_275);
nand U976 (N_976,N_346,N_171);
or U977 (N_977,N_306,N_91);
and U978 (N_978,N_246,N_374);
nor U979 (N_979,N_354,N_418);
nor U980 (N_980,N_263,N_463);
and U981 (N_981,N_114,N_317);
nand U982 (N_982,N_185,N_98);
or U983 (N_983,N_265,N_123);
nand U984 (N_984,N_359,N_434);
nor U985 (N_985,N_304,N_131);
and U986 (N_986,N_408,N_469);
nor U987 (N_987,N_26,N_105);
nor U988 (N_988,N_313,N_18);
nor U989 (N_989,N_432,N_296);
or U990 (N_990,N_321,N_278);
or U991 (N_991,N_124,N_389);
nor U992 (N_992,N_144,N_203);
nand U993 (N_993,N_235,N_179);
and U994 (N_994,N_437,N_424);
xnor U995 (N_995,N_317,N_98);
xor U996 (N_996,N_114,N_360);
nand U997 (N_997,N_355,N_63);
or U998 (N_998,N_252,N_6);
nand U999 (N_999,N_183,N_140);
nor U1000 (N_1000,N_955,N_941);
nand U1001 (N_1001,N_511,N_874);
nand U1002 (N_1002,N_529,N_903);
xnor U1003 (N_1003,N_801,N_725);
or U1004 (N_1004,N_852,N_888);
and U1005 (N_1005,N_840,N_626);
nand U1006 (N_1006,N_567,N_655);
nand U1007 (N_1007,N_897,N_999);
xor U1008 (N_1008,N_792,N_550);
nand U1009 (N_1009,N_571,N_872);
and U1010 (N_1010,N_856,N_798);
or U1011 (N_1011,N_810,N_868);
nand U1012 (N_1012,N_913,N_618);
nor U1013 (N_1013,N_653,N_589);
or U1014 (N_1014,N_946,N_839);
and U1015 (N_1015,N_680,N_758);
and U1016 (N_1016,N_735,N_780);
xor U1017 (N_1017,N_776,N_826);
and U1018 (N_1018,N_960,N_821);
or U1019 (N_1019,N_578,N_790);
nor U1020 (N_1020,N_895,N_564);
nor U1021 (N_1021,N_814,N_817);
and U1022 (N_1022,N_679,N_682);
nand U1023 (N_1023,N_527,N_530);
nand U1024 (N_1024,N_560,N_849);
or U1025 (N_1025,N_835,N_968);
and U1026 (N_1026,N_995,N_741);
nor U1027 (N_1027,N_555,N_642);
and U1028 (N_1028,N_966,N_886);
xnor U1029 (N_1029,N_557,N_635);
and U1030 (N_1030,N_911,N_942);
or U1031 (N_1031,N_640,N_883);
or U1032 (N_1032,N_611,N_787);
xor U1033 (N_1033,N_918,N_534);
nand U1034 (N_1034,N_580,N_851);
xnor U1035 (N_1035,N_882,N_771);
or U1036 (N_1036,N_685,N_985);
xnor U1037 (N_1037,N_768,N_830);
or U1038 (N_1038,N_742,N_535);
xor U1039 (N_1039,N_881,N_816);
or U1040 (N_1040,N_880,N_753);
or U1041 (N_1041,N_850,N_538);
nand U1042 (N_1042,N_879,N_854);
xnor U1043 (N_1043,N_605,N_834);
nand U1044 (N_1044,N_965,N_857);
or U1045 (N_1045,N_583,N_670);
xnor U1046 (N_1046,N_979,N_774);
nand U1047 (N_1047,N_772,N_733);
xnor U1048 (N_1048,N_971,N_623);
xor U1049 (N_1049,N_706,N_590);
nand U1050 (N_1050,N_906,N_683);
and U1051 (N_1051,N_637,N_656);
or U1052 (N_1052,N_820,N_700);
or U1053 (N_1053,N_707,N_908);
xor U1054 (N_1054,N_940,N_657);
xor U1055 (N_1055,N_989,N_639);
xnor U1056 (N_1056,N_812,N_508);
or U1057 (N_1057,N_842,N_689);
xor U1058 (N_1058,N_586,N_982);
xnor U1059 (N_1059,N_907,N_691);
nand U1060 (N_1060,N_565,N_766);
nor U1061 (N_1061,N_576,N_591);
nor U1062 (N_1062,N_953,N_891);
nand U1063 (N_1063,N_582,N_693);
or U1064 (N_1064,N_734,N_935);
nand U1065 (N_1065,N_944,N_889);
nor U1066 (N_1066,N_559,N_617);
xor U1067 (N_1067,N_797,N_896);
or U1068 (N_1068,N_606,N_638);
nand U1069 (N_1069,N_573,N_815);
nor U1070 (N_1070,N_750,N_751);
and U1071 (N_1071,N_947,N_556);
nor U1072 (N_1072,N_673,N_804);
nand U1073 (N_1073,N_848,N_825);
nand U1074 (N_1074,N_831,N_859);
xnor U1075 (N_1075,N_763,N_615);
xor U1076 (N_1076,N_662,N_841);
nand U1077 (N_1077,N_521,N_552);
or U1078 (N_1078,N_975,N_669);
xor U1079 (N_1079,N_684,N_869);
nand U1080 (N_1080,N_516,N_893);
xor U1081 (N_1081,N_870,N_809);
xnor U1082 (N_1082,N_858,N_745);
or U1083 (N_1083,N_844,N_972);
nand U1084 (N_1084,N_647,N_905);
xnor U1085 (N_1085,N_712,N_514);
or U1086 (N_1086,N_788,N_624);
nand U1087 (N_1087,N_900,N_658);
and U1088 (N_1088,N_708,N_926);
nand U1089 (N_1089,N_899,N_740);
and U1090 (N_1090,N_866,N_987);
and U1091 (N_1091,N_661,N_901);
or U1092 (N_1092,N_863,N_813);
nor U1093 (N_1093,N_607,N_961);
nor U1094 (N_1094,N_819,N_528);
and U1095 (N_1095,N_959,N_568);
xor U1096 (N_1096,N_885,N_549);
nand U1097 (N_1097,N_954,N_991);
and U1098 (N_1098,N_577,N_934);
nor U1099 (N_1099,N_631,N_986);
nor U1100 (N_1100,N_919,N_778);
xnor U1101 (N_1101,N_862,N_930);
nor U1102 (N_1102,N_686,N_978);
or U1103 (N_1103,N_633,N_505);
nand U1104 (N_1104,N_915,N_931);
xor U1105 (N_1105,N_558,N_600);
xnor U1106 (N_1106,N_988,N_922);
xor U1107 (N_1107,N_561,N_805);
and U1108 (N_1108,N_646,N_619);
and U1109 (N_1109,N_634,N_553);
xor U1110 (N_1110,N_864,N_981);
or U1111 (N_1111,N_699,N_838);
xor U1112 (N_1112,N_936,N_599);
xor U1113 (N_1113,N_724,N_824);
or U1114 (N_1114,N_546,N_504);
and U1115 (N_1115,N_932,N_672);
and U1116 (N_1116,N_920,N_917);
xor U1117 (N_1117,N_747,N_976);
and U1118 (N_1118,N_594,N_752);
nor U1119 (N_1119,N_519,N_629);
nor U1120 (N_1120,N_543,N_924);
nand U1121 (N_1121,N_613,N_717);
nand U1122 (N_1122,N_645,N_974);
xor U1123 (N_1123,N_769,N_997);
and U1124 (N_1124,N_595,N_873);
and U1125 (N_1125,N_929,N_531);
or U1126 (N_1126,N_608,N_865);
nand U1127 (N_1127,N_588,N_721);
or U1128 (N_1128,N_784,N_566);
xor U1129 (N_1129,N_761,N_690);
nand U1130 (N_1130,N_542,N_861);
xor U1131 (N_1131,N_716,N_783);
nor U1132 (N_1132,N_695,N_912);
nor U1133 (N_1133,N_601,N_811);
and U1134 (N_1134,N_927,N_625);
xnor U1135 (N_1135,N_994,N_938);
xor U1136 (N_1136,N_644,N_948);
nand U1137 (N_1137,N_539,N_630);
nor U1138 (N_1138,N_973,N_536);
or U1139 (N_1139,N_703,N_800);
and U1140 (N_1140,N_894,N_674);
and U1141 (N_1141,N_803,N_525);
or U1142 (N_1142,N_943,N_789);
nor U1143 (N_1143,N_827,N_579);
and U1144 (N_1144,N_990,N_668);
and U1145 (N_1145,N_755,N_781);
xor U1146 (N_1146,N_678,N_620);
or U1147 (N_1147,N_727,N_822);
nor U1148 (N_1148,N_701,N_904);
xnor U1149 (N_1149,N_945,N_828);
nand U1150 (N_1150,N_962,N_748);
or U1151 (N_1151,N_501,N_983);
nand U1152 (N_1152,N_671,N_729);
xor U1153 (N_1153,N_964,N_969);
or U1154 (N_1154,N_833,N_796);
nor U1155 (N_1155,N_709,N_950);
and U1156 (N_1156,N_602,N_933);
or U1157 (N_1157,N_587,N_609);
nor U1158 (N_1158,N_612,N_916);
nand U1159 (N_1159,N_984,N_520);
xor U1160 (N_1160,N_726,N_643);
and U1161 (N_1161,N_537,N_597);
nor U1162 (N_1162,N_795,N_697);
nor U1163 (N_1163,N_570,N_837);
nor U1164 (N_1164,N_547,N_677);
or U1165 (N_1165,N_925,N_939);
and U1166 (N_1166,N_676,N_794);
or U1167 (N_1167,N_736,N_698);
xor U1168 (N_1168,N_584,N_977);
nor U1169 (N_1169,N_749,N_764);
xnor U1170 (N_1170,N_718,N_807);
xor U1171 (N_1171,N_890,N_506);
nor U1172 (N_1172,N_715,N_770);
and U1173 (N_1173,N_808,N_777);
and U1174 (N_1174,N_544,N_694);
or U1175 (N_1175,N_756,N_843);
nand U1176 (N_1176,N_762,N_711);
and U1177 (N_1177,N_738,N_688);
and U1178 (N_1178,N_730,N_949);
or U1179 (N_1179,N_710,N_628);
or U1180 (N_1180,N_887,N_667);
and U1181 (N_1181,N_760,N_902);
nor U1182 (N_1182,N_503,N_754);
and U1183 (N_1183,N_509,N_636);
xnor U1184 (N_1184,N_675,N_829);
nand U1185 (N_1185,N_779,N_993);
and U1186 (N_1186,N_875,N_541);
nor U1187 (N_1187,N_732,N_574);
nor U1188 (N_1188,N_967,N_951);
nand U1189 (N_1189,N_855,N_793);
nand U1190 (N_1190,N_853,N_649);
nor U1191 (N_1191,N_802,N_627);
or U1192 (N_1192,N_791,N_666);
nand U1193 (N_1193,N_540,N_757);
and U1194 (N_1194,N_575,N_512);
nand U1195 (N_1195,N_702,N_782);
or U1196 (N_1196,N_502,N_603);
and U1197 (N_1197,N_923,N_963);
and U1198 (N_1198,N_799,N_598);
xor U1199 (N_1199,N_518,N_775);
nor U1200 (N_1200,N_563,N_737);
xor U1201 (N_1201,N_759,N_692);
or U1202 (N_1202,N_500,N_739);
xnor U1203 (N_1203,N_845,N_818);
or U1204 (N_1204,N_562,N_523);
or U1205 (N_1205,N_722,N_705);
nor U1206 (N_1206,N_632,N_524);
nor U1207 (N_1207,N_921,N_723);
or U1208 (N_1208,N_515,N_714);
and U1209 (N_1209,N_876,N_614);
and U1210 (N_1210,N_720,N_604);
nor U1211 (N_1211,N_687,N_958);
and U1212 (N_1212,N_654,N_998);
nor U1213 (N_1213,N_952,N_719);
nor U1214 (N_1214,N_867,N_847);
or U1215 (N_1215,N_664,N_956);
nor U1216 (N_1216,N_545,N_786);
nand U1217 (N_1217,N_704,N_610);
or U1218 (N_1218,N_892,N_957);
nor U1219 (N_1219,N_832,N_522);
nand U1220 (N_1220,N_909,N_836);
nand U1221 (N_1221,N_871,N_652);
nor U1222 (N_1222,N_898,N_641);
nand U1223 (N_1223,N_713,N_937);
or U1224 (N_1224,N_622,N_696);
nor U1225 (N_1225,N_593,N_970);
nor U1226 (N_1226,N_592,N_659);
nand U1227 (N_1227,N_746,N_914);
and U1228 (N_1228,N_663,N_554);
xor U1229 (N_1229,N_665,N_878);
and U1230 (N_1230,N_910,N_569);
nor U1231 (N_1231,N_581,N_532);
xnor U1232 (N_1232,N_773,N_860);
xnor U1233 (N_1233,N_765,N_996);
and U1234 (N_1234,N_596,N_660);
xnor U1235 (N_1235,N_743,N_650);
and U1236 (N_1236,N_621,N_785);
nand U1237 (N_1237,N_510,N_806);
or U1238 (N_1238,N_681,N_548);
nor U1239 (N_1239,N_507,N_884);
nor U1240 (N_1240,N_992,N_651);
or U1241 (N_1241,N_648,N_767);
nand U1242 (N_1242,N_585,N_846);
nor U1243 (N_1243,N_513,N_728);
or U1244 (N_1244,N_616,N_744);
nand U1245 (N_1245,N_533,N_928);
nand U1246 (N_1246,N_877,N_731);
or U1247 (N_1247,N_823,N_572);
or U1248 (N_1248,N_526,N_980);
or U1249 (N_1249,N_517,N_551);
and U1250 (N_1250,N_807,N_753);
nor U1251 (N_1251,N_556,N_883);
xor U1252 (N_1252,N_925,N_783);
nand U1253 (N_1253,N_630,N_684);
nor U1254 (N_1254,N_567,N_949);
and U1255 (N_1255,N_841,N_759);
nand U1256 (N_1256,N_861,N_990);
nand U1257 (N_1257,N_866,N_942);
nor U1258 (N_1258,N_559,N_919);
xor U1259 (N_1259,N_830,N_751);
nor U1260 (N_1260,N_613,N_818);
nand U1261 (N_1261,N_963,N_991);
nand U1262 (N_1262,N_644,N_951);
and U1263 (N_1263,N_842,N_545);
xor U1264 (N_1264,N_927,N_525);
nand U1265 (N_1265,N_824,N_571);
nand U1266 (N_1266,N_745,N_525);
and U1267 (N_1267,N_925,N_988);
xnor U1268 (N_1268,N_760,N_670);
nand U1269 (N_1269,N_855,N_953);
and U1270 (N_1270,N_554,N_602);
and U1271 (N_1271,N_924,N_692);
xor U1272 (N_1272,N_817,N_546);
or U1273 (N_1273,N_606,N_602);
and U1274 (N_1274,N_679,N_564);
nor U1275 (N_1275,N_566,N_833);
or U1276 (N_1276,N_853,N_579);
or U1277 (N_1277,N_736,N_602);
or U1278 (N_1278,N_861,N_610);
and U1279 (N_1279,N_841,N_799);
or U1280 (N_1280,N_832,N_836);
xor U1281 (N_1281,N_544,N_675);
or U1282 (N_1282,N_543,N_958);
xnor U1283 (N_1283,N_849,N_991);
nand U1284 (N_1284,N_747,N_592);
nand U1285 (N_1285,N_551,N_689);
xor U1286 (N_1286,N_768,N_850);
nor U1287 (N_1287,N_536,N_623);
nor U1288 (N_1288,N_644,N_893);
or U1289 (N_1289,N_945,N_992);
nand U1290 (N_1290,N_654,N_751);
nand U1291 (N_1291,N_604,N_752);
xor U1292 (N_1292,N_936,N_636);
nor U1293 (N_1293,N_903,N_639);
nand U1294 (N_1294,N_747,N_636);
nor U1295 (N_1295,N_769,N_678);
nor U1296 (N_1296,N_682,N_542);
nand U1297 (N_1297,N_795,N_893);
nor U1298 (N_1298,N_683,N_835);
or U1299 (N_1299,N_915,N_608);
nor U1300 (N_1300,N_685,N_876);
or U1301 (N_1301,N_954,N_946);
xor U1302 (N_1302,N_683,N_806);
or U1303 (N_1303,N_758,N_998);
nand U1304 (N_1304,N_762,N_723);
nand U1305 (N_1305,N_924,N_976);
nor U1306 (N_1306,N_943,N_955);
and U1307 (N_1307,N_711,N_782);
and U1308 (N_1308,N_761,N_631);
xnor U1309 (N_1309,N_719,N_789);
or U1310 (N_1310,N_748,N_891);
and U1311 (N_1311,N_900,N_850);
or U1312 (N_1312,N_742,N_681);
nand U1313 (N_1313,N_877,N_932);
nor U1314 (N_1314,N_806,N_556);
nand U1315 (N_1315,N_798,N_793);
or U1316 (N_1316,N_979,N_541);
nor U1317 (N_1317,N_742,N_762);
nor U1318 (N_1318,N_745,N_949);
nand U1319 (N_1319,N_526,N_807);
or U1320 (N_1320,N_567,N_896);
nand U1321 (N_1321,N_567,N_942);
nand U1322 (N_1322,N_727,N_690);
or U1323 (N_1323,N_869,N_533);
nand U1324 (N_1324,N_770,N_971);
nor U1325 (N_1325,N_755,N_714);
and U1326 (N_1326,N_882,N_881);
or U1327 (N_1327,N_839,N_666);
nand U1328 (N_1328,N_931,N_552);
and U1329 (N_1329,N_960,N_816);
or U1330 (N_1330,N_745,N_788);
nand U1331 (N_1331,N_852,N_856);
or U1332 (N_1332,N_574,N_663);
nor U1333 (N_1333,N_878,N_908);
or U1334 (N_1334,N_643,N_651);
or U1335 (N_1335,N_561,N_519);
nand U1336 (N_1336,N_629,N_876);
nand U1337 (N_1337,N_630,N_556);
and U1338 (N_1338,N_603,N_636);
xnor U1339 (N_1339,N_781,N_944);
nand U1340 (N_1340,N_663,N_968);
and U1341 (N_1341,N_568,N_861);
and U1342 (N_1342,N_666,N_746);
nand U1343 (N_1343,N_749,N_517);
xor U1344 (N_1344,N_775,N_938);
nand U1345 (N_1345,N_720,N_566);
nor U1346 (N_1346,N_901,N_527);
and U1347 (N_1347,N_921,N_808);
nor U1348 (N_1348,N_996,N_784);
xnor U1349 (N_1349,N_504,N_943);
or U1350 (N_1350,N_736,N_584);
xor U1351 (N_1351,N_756,N_922);
xnor U1352 (N_1352,N_706,N_651);
and U1353 (N_1353,N_933,N_672);
and U1354 (N_1354,N_649,N_973);
nor U1355 (N_1355,N_836,N_765);
nor U1356 (N_1356,N_690,N_768);
and U1357 (N_1357,N_921,N_710);
or U1358 (N_1358,N_739,N_655);
xor U1359 (N_1359,N_705,N_786);
and U1360 (N_1360,N_534,N_752);
nor U1361 (N_1361,N_847,N_779);
nor U1362 (N_1362,N_890,N_617);
xor U1363 (N_1363,N_523,N_911);
and U1364 (N_1364,N_885,N_803);
nand U1365 (N_1365,N_967,N_750);
nand U1366 (N_1366,N_690,N_862);
nand U1367 (N_1367,N_657,N_891);
nand U1368 (N_1368,N_999,N_901);
nor U1369 (N_1369,N_992,N_633);
xor U1370 (N_1370,N_844,N_573);
and U1371 (N_1371,N_846,N_922);
nand U1372 (N_1372,N_955,N_785);
xnor U1373 (N_1373,N_507,N_815);
xor U1374 (N_1374,N_848,N_724);
nand U1375 (N_1375,N_945,N_757);
or U1376 (N_1376,N_864,N_615);
or U1377 (N_1377,N_940,N_899);
or U1378 (N_1378,N_514,N_593);
or U1379 (N_1379,N_983,N_866);
and U1380 (N_1380,N_534,N_672);
and U1381 (N_1381,N_618,N_794);
and U1382 (N_1382,N_538,N_574);
and U1383 (N_1383,N_717,N_971);
or U1384 (N_1384,N_624,N_873);
xnor U1385 (N_1385,N_849,N_537);
or U1386 (N_1386,N_529,N_800);
nand U1387 (N_1387,N_896,N_917);
nor U1388 (N_1388,N_791,N_690);
nor U1389 (N_1389,N_823,N_552);
xnor U1390 (N_1390,N_595,N_593);
nand U1391 (N_1391,N_521,N_936);
nand U1392 (N_1392,N_610,N_681);
or U1393 (N_1393,N_962,N_524);
nand U1394 (N_1394,N_688,N_573);
nor U1395 (N_1395,N_953,N_787);
xnor U1396 (N_1396,N_795,N_965);
nand U1397 (N_1397,N_896,N_523);
and U1398 (N_1398,N_604,N_743);
nor U1399 (N_1399,N_598,N_973);
xnor U1400 (N_1400,N_875,N_927);
or U1401 (N_1401,N_924,N_865);
or U1402 (N_1402,N_830,N_819);
nand U1403 (N_1403,N_777,N_838);
xor U1404 (N_1404,N_839,N_537);
nor U1405 (N_1405,N_986,N_938);
nand U1406 (N_1406,N_532,N_523);
and U1407 (N_1407,N_866,N_662);
xnor U1408 (N_1408,N_657,N_766);
nand U1409 (N_1409,N_895,N_767);
xnor U1410 (N_1410,N_649,N_815);
nor U1411 (N_1411,N_811,N_863);
nor U1412 (N_1412,N_754,N_864);
nand U1413 (N_1413,N_829,N_741);
nor U1414 (N_1414,N_502,N_895);
xnor U1415 (N_1415,N_858,N_991);
and U1416 (N_1416,N_707,N_685);
xor U1417 (N_1417,N_895,N_593);
and U1418 (N_1418,N_633,N_816);
or U1419 (N_1419,N_671,N_599);
nor U1420 (N_1420,N_523,N_949);
or U1421 (N_1421,N_931,N_705);
nand U1422 (N_1422,N_717,N_857);
xor U1423 (N_1423,N_942,N_654);
nor U1424 (N_1424,N_699,N_716);
or U1425 (N_1425,N_931,N_890);
or U1426 (N_1426,N_724,N_836);
and U1427 (N_1427,N_517,N_776);
and U1428 (N_1428,N_881,N_668);
xnor U1429 (N_1429,N_653,N_525);
or U1430 (N_1430,N_717,N_711);
or U1431 (N_1431,N_841,N_777);
nor U1432 (N_1432,N_850,N_767);
xnor U1433 (N_1433,N_927,N_576);
nor U1434 (N_1434,N_896,N_902);
nor U1435 (N_1435,N_610,N_675);
nand U1436 (N_1436,N_930,N_644);
xor U1437 (N_1437,N_933,N_589);
xor U1438 (N_1438,N_615,N_823);
nand U1439 (N_1439,N_969,N_664);
nand U1440 (N_1440,N_618,N_720);
nor U1441 (N_1441,N_646,N_695);
nor U1442 (N_1442,N_892,N_651);
nand U1443 (N_1443,N_881,N_779);
nor U1444 (N_1444,N_745,N_881);
nor U1445 (N_1445,N_782,N_946);
nor U1446 (N_1446,N_643,N_855);
xnor U1447 (N_1447,N_992,N_527);
and U1448 (N_1448,N_902,N_855);
and U1449 (N_1449,N_821,N_502);
and U1450 (N_1450,N_958,N_515);
nor U1451 (N_1451,N_881,N_896);
xnor U1452 (N_1452,N_639,N_907);
nor U1453 (N_1453,N_557,N_863);
and U1454 (N_1454,N_847,N_740);
nor U1455 (N_1455,N_574,N_869);
or U1456 (N_1456,N_839,N_616);
xor U1457 (N_1457,N_524,N_691);
nand U1458 (N_1458,N_946,N_910);
or U1459 (N_1459,N_630,N_908);
nand U1460 (N_1460,N_875,N_548);
xnor U1461 (N_1461,N_746,N_855);
and U1462 (N_1462,N_886,N_722);
or U1463 (N_1463,N_577,N_823);
and U1464 (N_1464,N_524,N_974);
and U1465 (N_1465,N_694,N_731);
or U1466 (N_1466,N_978,N_617);
nand U1467 (N_1467,N_548,N_520);
nor U1468 (N_1468,N_787,N_587);
nand U1469 (N_1469,N_648,N_661);
nand U1470 (N_1470,N_596,N_520);
or U1471 (N_1471,N_726,N_539);
or U1472 (N_1472,N_940,N_540);
xnor U1473 (N_1473,N_907,N_811);
nand U1474 (N_1474,N_689,N_780);
nor U1475 (N_1475,N_565,N_961);
and U1476 (N_1476,N_895,N_871);
or U1477 (N_1477,N_835,N_777);
nand U1478 (N_1478,N_902,N_933);
xor U1479 (N_1479,N_972,N_897);
xor U1480 (N_1480,N_694,N_545);
and U1481 (N_1481,N_599,N_702);
nor U1482 (N_1482,N_509,N_694);
and U1483 (N_1483,N_504,N_693);
nand U1484 (N_1484,N_743,N_612);
and U1485 (N_1485,N_905,N_550);
xnor U1486 (N_1486,N_584,N_854);
and U1487 (N_1487,N_873,N_833);
xor U1488 (N_1488,N_751,N_808);
and U1489 (N_1489,N_912,N_909);
and U1490 (N_1490,N_561,N_657);
nor U1491 (N_1491,N_648,N_716);
xor U1492 (N_1492,N_738,N_708);
nand U1493 (N_1493,N_801,N_702);
xor U1494 (N_1494,N_761,N_636);
nand U1495 (N_1495,N_782,N_897);
xnor U1496 (N_1496,N_691,N_504);
nand U1497 (N_1497,N_943,N_566);
nand U1498 (N_1498,N_606,N_975);
or U1499 (N_1499,N_990,N_684);
and U1500 (N_1500,N_1271,N_1019);
or U1501 (N_1501,N_1175,N_1146);
xnor U1502 (N_1502,N_1205,N_1290);
xor U1503 (N_1503,N_1497,N_1294);
or U1504 (N_1504,N_1080,N_1253);
or U1505 (N_1505,N_1468,N_1198);
or U1506 (N_1506,N_1001,N_1337);
nor U1507 (N_1507,N_1260,N_1270);
nand U1508 (N_1508,N_1400,N_1144);
xnor U1509 (N_1509,N_1487,N_1318);
xnor U1510 (N_1510,N_1126,N_1339);
and U1511 (N_1511,N_1491,N_1315);
nor U1512 (N_1512,N_1119,N_1121);
nor U1513 (N_1513,N_1051,N_1098);
or U1514 (N_1514,N_1393,N_1344);
and U1515 (N_1515,N_1472,N_1402);
nor U1516 (N_1516,N_1427,N_1350);
xnor U1517 (N_1517,N_1461,N_1475);
and U1518 (N_1518,N_1392,N_1473);
xor U1519 (N_1519,N_1317,N_1432);
or U1520 (N_1520,N_1215,N_1219);
xor U1521 (N_1521,N_1478,N_1267);
or U1522 (N_1522,N_1322,N_1469);
nor U1523 (N_1523,N_1334,N_1272);
or U1524 (N_1524,N_1371,N_1004);
nand U1525 (N_1525,N_1394,N_1380);
nand U1526 (N_1526,N_1189,N_1378);
xnor U1527 (N_1527,N_1025,N_1153);
xor U1528 (N_1528,N_1125,N_1244);
xnor U1529 (N_1529,N_1314,N_1454);
nand U1530 (N_1530,N_1134,N_1470);
xnor U1531 (N_1531,N_1405,N_1381);
nand U1532 (N_1532,N_1423,N_1029);
or U1533 (N_1533,N_1440,N_1073);
and U1534 (N_1534,N_1237,N_1228);
and U1535 (N_1535,N_1036,N_1332);
nor U1536 (N_1536,N_1081,N_1048);
or U1537 (N_1537,N_1164,N_1054);
nor U1538 (N_1538,N_1361,N_1325);
nand U1539 (N_1539,N_1390,N_1068);
xnor U1540 (N_1540,N_1213,N_1488);
nor U1541 (N_1541,N_1217,N_1407);
nor U1542 (N_1542,N_1258,N_1150);
or U1543 (N_1543,N_1462,N_1042);
nor U1544 (N_1544,N_1287,N_1452);
or U1545 (N_1545,N_1474,N_1047);
or U1546 (N_1546,N_1075,N_1159);
nand U1547 (N_1547,N_1338,N_1458);
xnor U1548 (N_1548,N_1301,N_1148);
nor U1549 (N_1549,N_1255,N_1089);
or U1550 (N_1550,N_1070,N_1476);
and U1551 (N_1551,N_1005,N_1037);
and U1552 (N_1552,N_1052,N_1031);
xor U1553 (N_1553,N_1021,N_1082);
nand U1554 (N_1554,N_1499,N_1303);
nor U1555 (N_1555,N_1056,N_1450);
and U1556 (N_1556,N_1254,N_1046);
or U1557 (N_1557,N_1050,N_1349);
and U1558 (N_1558,N_1386,N_1277);
and U1559 (N_1559,N_1252,N_1120);
and U1560 (N_1560,N_1341,N_1142);
xnor U1561 (N_1561,N_1199,N_1094);
and U1562 (N_1562,N_1492,N_1329);
xnor U1563 (N_1563,N_1077,N_1261);
and U1564 (N_1564,N_1279,N_1494);
xnor U1565 (N_1565,N_1248,N_1433);
or U1566 (N_1566,N_1097,N_1323);
and U1567 (N_1567,N_1220,N_1059);
or U1568 (N_1568,N_1284,N_1280);
and U1569 (N_1569,N_1417,N_1099);
nand U1570 (N_1570,N_1293,N_1319);
nor U1571 (N_1571,N_1456,N_1002);
or U1572 (N_1572,N_1058,N_1208);
and U1573 (N_1573,N_1214,N_1291);
nor U1574 (N_1574,N_1145,N_1108);
and U1575 (N_1575,N_1365,N_1235);
and U1576 (N_1576,N_1460,N_1396);
or U1577 (N_1577,N_1328,N_1112);
and U1578 (N_1578,N_1359,N_1116);
and U1579 (N_1579,N_1465,N_1026);
and U1580 (N_1580,N_1347,N_1067);
nand U1581 (N_1581,N_1057,N_1086);
and U1582 (N_1582,N_1201,N_1266);
and U1583 (N_1583,N_1482,N_1195);
nand U1584 (N_1584,N_1012,N_1209);
xnor U1585 (N_1585,N_1246,N_1084);
or U1586 (N_1586,N_1447,N_1128);
nor U1587 (N_1587,N_1348,N_1449);
and U1588 (N_1588,N_1168,N_1188);
nand U1589 (N_1589,N_1178,N_1388);
and U1590 (N_1590,N_1354,N_1045);
and U1591 (N_1591,N_1111,N_1321);
nor U1592 (N_1592,N_1009,N_1180);
and U1593 (N_1593,N_1256,N_1249);
nor U1594 (N_1594,N_1282,N_1300);
and U1595 (N_1595,N_1444,N_1218);
and U1596 (N_1596,N_1434,N_1397);
nand U1597 (N_1597,N_1308,N_1439);
and U1598 (N_1598,N_1040,N_1490);
or U1599 (N_1599,N_1498,N_1181);
nor U1600 (N_1600,N_1281,N_1418);
nand U1601 (N_1601,N_1333,N_1000);
xor U1602 (N_1602,N_1240,N_1053);
nor U1603 (N_1603,N_1395,N_1302);
xnor U1604 (N_1604,N_1273,N_1483);
xor U1605 (N_1605,N_1250,N_1185);
nand U1606 (N_1606,N_1411,N_1191);
nand U1607 (N_1607,N_1151,N_1143);
or U1608 (N_1608,N_1355,N_1165);
nand U1609 (N_1609,N_1182,N_1389);
nand U1610 (N_1610,N_1336,N_1162);
nor U1611 (N_1611,N_1278,N_1018);
xor U1612 (N_1612,N_1342,N_1192);
or U1613 (N_1613,N_1232,N_1442);
and U1614 (N_1614,N_1131,N_1416);
nand U1615 (N_1615,N_1129,N_1179);
nand U1616 (N_1616,N_1072,N_1413);
or U1617 (N_1617,N_1172,N_1312);
or U1618 (N_1618,N_1136,N_1269);
nor U1619 (N_1619,N_1481,N_1352);
nor U1620 (N_1620,N_1231,N_1107);
or U1621 (N_1621,N_1177,N_1197);
xnor U1622 (N_1622,N_1230,N_1095);
nor U1623 (N_1623,N_1010,N_1457);
xnor U1624 (N_1624,N_1257,N_1202);
nor U1625 (N_1625,N_1014,N_1289);
nand U1626 (N_1626,N_1114,N_1087);
or U1627 (N_1627,N_1229,N_1356);
nand U1628 (N_1628,N_1455,N_1043);
nor U1629 (N_1629,N_1376,N_1373);
nand U1630 (N_1630,N_1234,N_1124);
nor U1631 (N_1631,N_1034,N_1425);
nand U1632 (N_1632,N_1268,N_1484);
and U1633 (N_1633,N_1306,N_1101);
nand U1634 (N_1634,N_1083,N_1436);
nand U1635 (N_1635,N_1368,N_1410);
xnor U1636 (N_1636,N_1028,N_1204);
and U1637 (N_1637,N_1216,N_1055);
nand U1638 (N_1638,N_1115,N_1173);
and U1639 (N_1639,N_1309,N_1200);
or U1640 (N_1640,N_1362,N_1438);
xor U1641 (N_1641,N_1013,N_1297);
or U1642 (N_1642,N_1275,N_1313);
nor U1643 (N_1643,N_1123,N_1091);
xor U1644 (N_1644,N_1139,N_1403);
nor U1645 (N_1645,N_1343,N_1135);
nor U1646 (N_1646,N_1307,N_1422);
and U1647 (N_1647,N_1466,N_1154);
or U1648 (N_1648,N_1011,N_1008);
xor U1649 (N_1649,N_1239,N_1259);
nor U1650 (N_1650,N_1316,N_1412);
or U1651 (N_1651,N_1207,N_1074);
nor U1652 (N_1652,N_1221,N_1078);
and U1653 (N_1653,N_1193,N_1076);
xnor U1654 (N_1654,N_1156,N_1263);
or U1655 (N_1655,N_1327,N_1238);
or U1656 (N_1656,N_1069,N_1027);
nand U1657 (N_1657,N_1363,N_1431);
nand U1658 (N_1658,N_1241,N_1190);
and U1659 (N_1659,N_1035,N_1437);
or U1660 (N_1660,N_1443,N_1038);
xnor U1661 (N_1661,N_1104,N_1435);
nor U1662 (N_1662,N_1285,N_1419);
or U1663 (N_1663,N_1226,N_1224);
xor U1664 (N_1664,N_1496,N_1196);
xor U1665 (N_1665,N_1044,N_1464);
xor U1666 (N_1666,N_1007,N_1206);
and U1667 (N_1667,N_1424,N_1030);
xor U1668 (N_1668,N_1369,N_1236);
nor U1669 (N_1669,N_1167,N_1066);
and U1670 (N_1670,N_1299,N_1366);
nor U1671 (N_1671,N_1184,N_1326);
or U1672 (N_1672,N_1064,N_1370);
nand U1673 (N_1673,N_1382,N_1351);
nand U1674 (N_1674,N_1331,N_1033);
and U1675 (N_1675,N_1203,N_1251);
and U1676 (N_1676,N_1305,N_1161);
nor U1677 (N_1677,N_1374,N_1485);
nor U1678 (N_1678,N_1155,N_1233);
xnor U1679 (N_1679,N_1105,N_1049);
or U1680 (N_1680,N_1090,N_1093);
nand U1681 (N_1681,N_1109,N_1428);
and U1682 (N_1682,N_1377,N_1345);
nor U1683 (N_1683,N_1071,N_1157);
xor U1684 (N_1684,N_1140,N_1493);
nor U1685 (N_1685,N_1286,N_1357);
and U1686 (N_1686,N_1262,N_1391);
and U1687 (N_1687,N_1430,N_1292);
xor U1688 (N_1688,N_1360,N_1110);
nor U1689 (N_1689,N_1174,N_1186);
or U1690 (N_1690,N_1210,N_1247);
and U1691 (N_1691,N_1088,N_1212);
nor U1692 (N_1692,N_1222,N_1274);
nor U1693 (N_1693,N_1384,N_1065);
nand U1694 (N_1694,N_1096,N_1409);
or U1695 (N_1695,N_1477,N_1243);
nor U1696 (N_1696,N_1459,N_1296);
nor U1697 (N_1697,N_1364,N_1022);
nand U1698 (N_1698,N_1063,N_1023);
nor U1699 (N_1699,N_1163,N_1152);
nor U1700 (N_1700,N_1324,N_1103);
nand U1701 (N_1701,N_1039,N_1242);
or U1702 (N_1702,N_1379,N_1006);
and U1703 (N_1703,N_1194,N_1429);
xor U1704 (N_1704,N_1137,N_1016);
or U1705 (N_1705,N_1102,N_1024);
nor U1706 (N_1706,N_1445,N_1117);
or U1707 (N_1707,N_1311,N_1062);
xnor U1708 (N_1708,N_1463,N_1169);
xor U1709 (N_1709,N_1404,N_1426);
xor U1710 (N_1710,N_1346,N_1176);
nand U1711 (N_1711,N_1017,N_1138);
xor U1712 (N_1712,N_1288,N_1100);
or U1713 (N_1713,N_1441,N_1495);
nand U1714 (N_1714,N_1118,N_1158);
nand U1715 (N_1715,N_1471,N_1132);
nand U1716 (N_1716,N_1170,N_1320);
xnor U1717 (N_1717,N_1295,N_1406);
nor U1718 (N_1718,N_1171,N_1298);
nor U1719 (N_1719,N_1113,N_1453);
or U1720 (N_1720,N_1304,N_1340);
xor U1721 (N_1721,N_1372,N_1421);
xnor U1722 (N_1722,N_1020,N_1353);
or U1723 (N_1723,N_1467,N_1032);
and U1724 (N_1724,N_1283,N_1264);
or U1725 (N_1725,N_1147,N_1276);
nand U1726 (N_1726,N_1387,N_1130);
xnor U1727 (N_1727,N_1358,N_1160);
xor U1728 (N_1728,N_1489,N_1223);
nor U1729 (N_1729,N_1383,N_1211);
xnor U1730 (N_1730,N_1141,N_1385);
nor U1731 (N_1731,N_1227,N_1448);
nor U1732 (N_1732,N_1085,N_1166);
xnor U1733 (N_1733,N_1401,N_1408);
nand U1734 (N_1734,N_1183,N_1446);
xnor U1735 (N_1735,N_1133,N_1375);
xnor U1736 (N_1736,N_1245,N_1225);
and U1737 (N_1737,N_1061,N_1335);
xor U1738 (N_1738,N_1187,N_1079);
nand U1739 (N_1739,N_1265,N_1003);
xor U1740 (N_1740,N_1420,N_1398);
or U1741 (N_1741,N_1486,N_1015);
or U1742 (N_1742,N_1092,N_1399);
xnor U1743 (N_1743,N_1060,N_1106);
nor U1744 (N_1744,N_1041,N_1451);
or U1745 (N_1745,N_1367,N_1149);
nor U1746 (N_1746,N_1330,N_1479);
nand U1747 (N_1747,N_1127,N_1122);
nand U1748 (N_1748,N_1310,N_1480);
or U1749 (N_1749,N_1415,N_1414);
or U1750 (N_1750,N_1216,N_1186);
or U1751 (N_1751,N_1368,N_1067);
nor U1752 (N_1752,N_1478,N_1166);
and U1753 (N_1753,N_1404,N_1335);
and U1754 (N_1754,N_1172,N_1409);
and U1755 (N_1755,N_1006,N_1329);
nand U1756 (N_1756,N_1291,N_1242);
nand U1757 (N_1757,N_1117,N_1373);
and U1758 (N_1758,N_1468,N_1304);
nand U1759 (N_1759,N_1002,N_1166);
and U1760 (N_1760,N_1322,N_1490);
and U1761 (N_1761,N_1496,N_1219);
nor U1762 (N_1762,N_1403,N_1334);
nor U1763 (N_1763,N_1488,N_1285);
nand U1764 (N_1764,N_1171,N_1251);
and U1765 (N_1765,N_1025,N_1095);
or U1766 (N_1766,N_1146,N_1320);
nand U1767 (N_1767,N_1080,N_1379);
and U1768 (N_1768,N_1084,N_1038);
or U1769 (N_1769,N_1497,N_1264);
and U1770 (N_1770,N_1426,N_1038);
nor U1771 (N_1771,N_1418,N_1324);
xnor U1772 (N_1772,N_1230,N_1171);
or U1773 (N_1773,N_1366,N_1112);
nor U1774 (N_1774,N_1281,N_1139);
xor U1775 (N_1775,N_1379,N_1422);
or U1776 (N_1776,N_1168,N_1032);
nor U1777 (N_1777,N_1144,N_1206);
and U1778 (N_1778,N_1436,N_1052);
nor U1779 (N_1779,N_1434,N_1021);
and U1780 (N_1780,N_1082,N_1271);
nand U1781 (N_1781,N_1494,N_1415);
xnor U1782 (N_1782,N_1415,N_1071);
xor U1783 (N_1783,N_1332,N_1322);
and U1784 (N_1784,N_1280,N_1059);
nor U1785 (N_1785,N_1438,N_1395);
xnor U1786 (N_1786,N_1440,N_1318);
and U1787 (N_1787,N_1125,N_1233);
xnor U1788 (N_1788,N_1227,N_1007);
xnor U1789 (N_1789,N_1012,N_1331);
xnor U1790 (N_1790,N_1314,N_1375);
nand U1791 (N_1791,N_1225,N_1346);
and U1792 (N_1792,N_1298,N_1486);
xnor U1793 (N_1793,N_1147,N_1262);
and U1794 (N_1794,N_1270,N_1301);
nand U1795 (N_1795,N_1097,N_1134);
nor U1796 (N_1796,N_1147,N_1429);
nand U1797 (N_1797,N_1221,N_1453);
nand U1798 (N_1798,N_1236,N_1167);
xnor U1799 (N_1799,N_1202,N_1056);
nand U1800 (N_1800,N_1237,N_1014);
or U1801 (N_1801,N_1126,N_1155);
nor U1802 (N_1802,N_1495,N_1169);
nand U1803 (N_1803,N_1296,N_1264);
or U1804 (N_1804,N_1469,N_1480);
and U1805 (N_1805,N_1362,N_1015);
nand U1806 (N_1806,N_1257,N_1356);
nor U1807 (N_1807,N_1367,N_1071);
or U1808 (N_1808,N_1377,N_1431);
xnor U1809 (N_1809,N_1397,N_1314);
nand U1810 (N_1810,N_1036,N_1297);
xnor U1811 (N_1811,N_1243,N_1294);
and U1812 (N_1812,N_1300,N_1054);
xor U1813 (N_1813,N_1466,N_1284);
and U1814 (N_1814,N_1160,N_1136);
nand U1815 (N_1815,N_1365,N_1199);
nor U1816 (N_1816,N_1262,N_1224);
nor U1817 (N_1817,N_1174,N_1270);
or U1818 (N_1818,N_1406,N_1413);
or U1819 (N_1819,N_1385,N_1381);
xnor U1820 (N_1820,N_1002,N_1393);
or U1821 (N_1821,N_1370,N_1119);
nor U1822 (N_1822,N_1279,N_1356);
or U1823 (N_1823,N_1458,N_1184);
nor U1824 (N_1824,N_1038,N_1346);
nor U1825 (N_1825,N_1435,N_1441);
and U1826 (N_1826,N_1417,N_1351);
or U1827 (N_1827,N_1239,N_1202);
xnor U1828 (N_1828,N_1416,N_1223);
nor U1829 (N_1829,N_1188,N_1446);
nor U1830 (N_1830,N_1324,N_1367);
nand U1831 (N_1831,N_1297,N_1283);
nand U1832 (N_1832,N_1109,N_1217);
or U1833 (N_1833,N_1395,N_1321);
nor U1834 (N_1834,N_1483,N_1118);
and U1835 (N_1835,N_1464,N_1487);
and U1836 (N_1836,N_1330,N_1207);
or U1837 (N_1837,N_1001,N_1367);
nand U1838 (N_1838,N_1354,N_1205);
nand U1839 (N_1839,N_1350,N_1341);
nor U1840 (N_1840,N_1207,N_1383);
and U1841 (N_1841,N_1341,N_1252);
or U1842 (N_1842,N_1233,N_1403);
or U1843 (N_1843,N_1409,N_1405);
nand U1844 (N_1844,N_1217,N_1155);
or U1845 (N_1845,N_1355,N_1051);
and U1846 (N_1846,N_1102,N_1037);
or U1847 (N_1847,N_1158,N_1094);
or U1848 (N_1848,N_1309,N_1261);
or U1849 (N_1849,N_1194,N_1200);
nor U1850 (N_1850,N_1309,N_1419);
and U1851 (N_1851,N_1443,N_1367);
xor U1852 (N_1852,N_1269,N_1131);
xnor U1853 (N_1853,N_1357,N_1394);
or U1854 (N_1854,N_1333,N_1182);
xnor U1855 (N_1855,N_1109,N_1464);
or U1856 (N_1856,N_1276,N_1127);
nand U1857 (N_1857,N_1268,N_1126);
or U1858 (N_1858,N_1127,N_1245);
nand U1859 (N_1859,N_1298,N_1023);
nor U1860 (N_1860,N_1157,N_1316);
nor U1861 (N_1861,N_1093,N_1279);
xnor U1862 (N_1862,N_1414,N_1299);
and U1863 (N_1863,N_1361,N_1114);
and U1864 (N_1864,N_1317,N_1070);
or U1865 (N_1865,N_1343,N_1434);
nor U1866 (N_1866,N_1119,N_1185);
nor U1867 (N_1867,N_1049,N_1363);
or U1868 (N_1868,N_1395,N_1320);
nand U1869 (N_1869,N_1400,N_1185);
nor U1870 (N_1870,N_1418,N_1028);
nor U1871 (N_1871,N_1011,N_1048);
or U1872 (N_1872,N_1440,N_1182);
nor U1873 (N_1873,N_1361,N_1231);
xnor U1874 (N_1874,N_1148,N_1216);
nand U1875 (N_1875,N_1030,N_1407);
nand U1876 (N_1876,N_1266,N_1209);
or U1877 (N_1877,N_1225,N_1103);
nor U1878 (N_1878,N_1178,N_1462);
and U1879 (N_1879,N_1110,N_1414);
or U1880 (N_1880,N_1488,N_1153);
nand U1881 (N_1881,N_1427,N_1318);
nand U1882 (N_1882,N_1117,N_1311);
nor U1883 (N_1883,N_1224,N_1306);
and U1884 (N_1884,N_1361,N_1287);
or U1885 (N_1885,N_1220,N_1381);
or U1886 (N_1886,N_1470,N_1129);
and U1887 (N_1887,N_1434,N_1114);
or U1888 (N_1888,N_1289,N_1453);
and U1889 (N_1889,N_1297,N_1143);
or U1890 (N_1890,N_1357,N_1448);
xnor U1891 (N_1891,N_1272,N_1091);
and U1892 (N_1892,N_1420,N_1052);
xor U1893 (N_1893,N_1415,N_1043);
xnor U1894 (N_1894,N_1461,N_1349);
xor U1895 (N_1895,N_1487,N_1480);
nand U1896 (N_1896,N_1470,N_1150);
and U1897 (N_1897,N_1360,N_1271);
or U1898 (N_1898,N_1383,N_1319);
nand U1899 (N_1899,N_1023,N_1192);
nor U1900 (N_1900,N_1078,N_1038);
nor U1901 (N_1901,N_1158,N_1481);
nand U1902 (N_1902,N_1197,N_1174);
nor U1903 (N_1903,N_1425,N_1431);
xor U1904 (N_1904,N_1418,N_1057);
nand U1905 (N_1905,N_1436,N_1475);
nand U1906 (N_1906,N_1228,N_1355);
or U1907 (N_1907,N_1055,N_1442);
and U1908 (N_1908,N_1002,N_1128);
or U1909 (N_1909,N_1282,N_1467);
nor U1910 (N_1910,N_1254,N_1114);
nor U1911 (N_1911,N_1470,N_1295);
xor U1912 (N_1912,N_1425,N_1499);
xor U1913 (N_1913,N_1198,N_1132);
nand U1914 (N_1914,N_1417,N_1188);
nand U1915 (N_1915,N_1434,N_1079);
nor U1916 (N_1916,N_1435,N_1369);
xnor U1917 (N_1917,N_1070,N_1017);
xor U1918 (N_1918,N_1208,N_1083);
or U1919 (N_1919,N_1056,N_1302);
and U1920 (N_1920,N_1353,N_1058);
nor U1921 (N_1921,N_1039,N_1342);
and U1922 (N_1922,N_1306,N_1420);
xor U1923 (N_1923,N_1174,N_1280);
xor U1924 (N_1924,N_1127,N_1431);
and U1925 (N_1925,N_1284,N_1294);
and U1926 (N_1926,N_1406,N_1085);
nor U1927 (N_1927,N_1077,N_1209);
xor U1928 (N_1928,N_1391,N_1338);
xnor U1929 (N_1929,N_1321,N_1110);
or U1930 (N_1930,N_1285,N_1186);
nor U1931 (N_1931,N_1004,N_1094);
nor U1932 (N_1932,N_1279,N_1393);
or U1933 (N_1933,N_1159,N_1295);
or U1934 (N_1934,N_1178,N_1219);
nand U1935 (N_1935,N_1331,N_1177);
xnor U1936 (N_1936,N_1164,N_1487);
nand U1937 (N_1937,N_1036,N_1333);
nand U1938 (N_1938,N_1249,N_1492);
or U1939 (N_1939,N_1263,N_1419);
nand U1940 (N_1940,N_1022,N_1438);
nor U1941 (N_1941,N_1120,N_1215);
nor U1942 (N_1942,N_1242,N_1116);
or U1943 (N_1943,N_1168,N_1282);
nand U1944 (N_1944,N_1145,N_1241);
nand U1945 (N_1945,N_1217,N_1037);
nor U1946 (N_1946,N_1068,N_1447);
or U1947 (N_1947,N_1367,N_1142);
nand U1948 (N_1948,N_1002,N_1160);
xor U1949 (N_1949,N_1288,N_1295);
or U1950 (N_1950,N_1263,N_1358);
or U1951 (N_1951,N_1308,N_1392);
nor U1952 (N_1952,N_1304,N_1316);
and U1953 (N_1953,N_1469,N_1441);
nand U1954 (N_1954,N_1360,N_1276);
nor U1955 (N_1955,N_1371,N_1078);
or U1956 (N_1956,N_1121,N_1057);
xor U1957 (N_1957,N_1349,N_1272);
nand U1958 (N_1958,N_1451,N_1306);
xnor U1959 (N_1959,N_1103,N_1052);
or U1960 (N_1960,N_1146,N_1214);
nor U1961 (N_1961,N_1018,N_1285);
and U1962 (N_1962,N_1339,N_1489);
nor U1963 (N_1963,N_1152,N_1113);
nor U1964 (N_1964,N_1389,N_1264);
xnor U1965 (N_1965,N_1250,N_1389);
and U1966 (N_1966,N_1165,N_1281);
nor U1967 (N_1967,N_1067,N_1245);
and U1968 (N_1968,N_1090,N_1405);
nand U1969 (N_1969,N_1101,N_1329);
nor U1970 (N_1970,N_1213,N_1424);
or U1971 (N_1971,N_1481,N_1337);
or U1972 (N_1972,N_1499,N_1338);
nand U1973 (N_1973,N_1333,N_1039);
or U1974 (N_1974,N_1427,N_1381);
nand U1975 (N_1975,N_1004,N_1275);
nand U1976 (N_1976,N_1250,N_1340);
or U1977 (N_1977,N_1389,N_1353);
and U1978 (N_1978,N_1271,N_1168);
nor U1979 (N_1979,N_1160,N_1055);
nand U1980 (N_1980,N_1310,N_1362);
and U1981 (N_1981,N_1299,N_1011);
nand U1982 (N_1982,N_1128,N_1198);
nor U1983 (N_1983,N_1358,N_1167);
xnor U1984 (N_1984,N_1027,N_1008);
and U1985 (N_1985,N_1283,N_1019);
xnor U1986 (N_1986,N_1463,N_1167);
xnor U1987 (N_1987,N_1143,N_1223);
or U1988 (N_1988,N_1472,N_1286);
xor U1989 (N_1989,N_1222,N_1192);
nand U1990 (N_1990,N_1486,N_1029);
nor U1991 (N_1991,N_1203,N_1212);
xor U1992 (N_1992,N_1353,N_1126);
and U1993 (N_1993,N_1048,N_1189);
or U1994 (N_1994,N_1426,N_1166);
nor U1995 (N_1995,N_1228,N_1480);
or U1996 (N_1996,N_1130,N_1064);
nor U1997 (N_1997,N_1438,N_1094);
or U1998 (N_1998,N_1447,N_1487);
or U1999 (N_1999,N_1099,N_1309);
xnor U2000 (N_2000,N_1739,N_1672);
nor U2001 (N_2001,N_1743,N_1584);
or U2002 (N_2002,N_1781,N_1643);
nor U2003 (N_2003,N_1725,N_1699);
nor U2004 (N_2004,N_1652,N_1611);
and U2005 (N_2005,N_1581,N_1805);
xnor U2006 (N_2006,N_1825,N_1616);
xnor U2007 (N_2007,N_1697,N_1565);
and U2008 (N_2008,N_1744,N_1789);
xnor U2009 (N_2009,N_1836,N_1729);
nand U2010 (N_2010,N_1635,N_1712);
nand U2011 (N_2011,N_1797,N_1835);
xnor U2012 (N_2012,N_1833,N_1629);
or U2013 (N_2013,N_1579,N_1574);
and U2014 (N_2014,N_1686,N_1976);
and U2015 (N_2015,N_1543,N_1587);
and U2016 (N_2016,N_1909,N_1636);
and U2017 (N_2017,N_1875,N_1950);
xor U2018 (N_2018,N_1904,N_1801);
xor U2019 (N_2019,N_1598,N_1706);
nor U2020 (N_2020,N_1539,N_1834);
xnor U2021 (N_2021,N_1508,N_1595);
or U2022 (N_2022,N_1622,N_1995);
xnor U2023 (N_2023,N_1555,N_1787);
or U2024 (N_2024,N_1972,N_1823);
nand U2025 (N_2025,N_1804,N_1557);
nor U2026 (N_2026,N_1948,N_1917);
nand U2027 (N_2027,N_1958,N_1621);
or U2028 (N_2028,N_1762,N_1504);
xor U2029 (N_2029,N_1988,N_1940);
nor U2030 (N_2030,N_1602,N_1571);
and U2031 (N_2031,N_1883,N_1867);
nor U2032 (N_2032,N_1946,N_1967);
nor U2033 (N_2033,N_1774,N_1855);
nand U2034 (N_2034,N_1898,N_1936);
xor U2035 (N_2035,N_1580,N_1792);
or U2036 (N_2036,N_1600,N_1542);
or U2037 (N_2037,N_1906,N_1740);
and U2038 (N_2038,N_1554,N_1503);
nand U2039 (N_2039,N_1800,N_1943);
and U2040 (N_2040,N_1962,N_1684);
nor U2041 (N_2041,N_1612,N_1530);
nor U2042 (N_2042,N_1859,N_1737);
or U2043 (N_2043,N_1720,N_1960);
or U2044 (N_2044,N_1634,N_1793);
and U2045 (N_2045,N_1751,N_1773);
nand U2046 (N_2046,N_1664,N_1869);
nor U2047 (N_2047,N_1692,N_1517);
nor U2048 (N_2048,N_1933,N_1707);
nor U2049 (N_2049,N_1763,N_1527);
or U2050 (N_2050,N_1551,N_1870);
nor U2051 (N_2051,N_1724,N_1696);
nor U2052 (N_2052,N_1721,N_1726);
nor U2053 (N_2053,N_1914,N_1569);
or U2054 (N_2054,N_1886,N_1644);
nor U2055 (N_2055,N_1837,N_1887);
xor U2056 (N_2056,N_1884,N_1516);
or U2057 (N_2057,N_1889,N_1953);
nor U2058 (N_2058,N_1864,N_1784);
or U2059 (N_2059,N_1528,N_1659);
nor U2060 (N_2060,N_1997,N_1541);
nand U2061 (N_2061,N_1679,N_1657);
nor U2062 (N_2062,N_1925,N_1845);
xor U2063 (N_2063,N_1618,N_1710);
or U2064 (N_2064,N_1691,N_1892);
and U2065 (N_2065,N_1626,N_1844);
xor U2066 (N_2066,N_1601,N_1885);
nand U2067 (N_2067,N_1842,N_1897);
and U2068 (N_2068,N_1808,N_1986);
xor U2069 (N_2069,N_1561,N_1811);
or U2070 (N_2070,N_1782,N_1766);
and U2071 (N_2071,N_1944,N_1695);
and U2072 (N_2072,N_1977,N_1815);
or U2073 (N_2073,N_1814,N_1907);
nor U2074 (N_2074,N_1553,N_1778);
nand U2075 (N_2075,N_1893,N_1592);
xnor U2076 (N_2076,N_1973,N_1521);
or U2077 (N_2077,N_1756,N_1654);
xnor U2078 (N_2078,N_1783,N_1968);
nand U2079 (N_2079,N_1689,N_1798);
nor U2080 (N_2080,N_1704,N_1924);
or U2081 (N_2081,N_1556,N_1594);
nand U2082 (N_2082,N_1531,N_1918);
nand U2083 (N_2083,N_1639,N_1617);
or U2084 (N_2084,N_1529,N_1849);
nand U2085 (N_2085,N_1597,N_1871);
or U2086 (N_2086,N_1980,N_1730);
nand U2087 (N_2087,N_1735,N_1754);
and U2088 (N_2088,N_1812,N_1690);
xor U2089 (N_2089,N_1502,N_1873);
xor U2090 (N_2090,N_1619,N_1938);
or U2091 (N_2091,N_1593,N_1663);
xnor U2092 (N_2092,N_1882,N_1955);
and U2093 (N_2093,N_1670,N_1896);
and U2094 (N_2094,N_1665,N_1645);
or U2095 (N_2095,N_1640,N_1772);
and U2096 (N_2096,N_1714,N_1638);
nand U2097 (N_2097,N_1723,N_1637);
nor U2098 (N_2098,N_1613,N_1518);
nand U2099 (N_2099,N_1526,N_1916);
nand U2100 (N_2100,N_1620,N_1931);
xnor U2101 (N_2101,N_1757,N_1807);
xor U2102 (N_2102,N_1563,N_1777);
or U2103 (N_2103,N_1547,N_1848);
nor U2104 (N_2104,N_1591,N_1866);
xnor U2105 (N_2105,N_1568,N_1996);
nor U2106 (N_2106,N_1559,N_1853);
and U2107 (N_2107,N_1993,N_1850);
or U2108 (N_2108,N_1578,N_1603);
or U2109 (N_2109,N_1770,N_1974);
nand U2110 (N_2110,N_1546,N_1920);
or U2111 (N_2111,N_1749,N_1731);
xnor U2112 (N_2112,N_1919,N_1863);
or U2113 (N_2113,N_1966,N_1874);
or U2114 (N_2114,N_1668,N_1540);
and U2115 (N_2115,N_1820,N_1929);
or U2116 (N_2116,N_1838,N_1912);
or U2117 (N_2117,N_1794,N_1992);
nor U2118 (N_2118,N_1648,N_1915);
xor U2119 (N_2119,N_1562,N_1669);
and U2120 (N_2120,N_1846,N_1544);
xor U2121 (N_2121,N_1750,N_1548);
nor U2122 (N_2122,N_1840,N_1839);
nand U2123 (N_2123,N_1649,N_1716);
nand U2124 (N_2124,N_1558,N_1514);
nand U2125 (N_2125,N_1590,N_1501);
or U2126 (N_2126,N_1956,N_1978);
nor U2127 (N_2127,N_1566,N_1901);
nor U2128 (N_2128,N_1856,N_1513);
nor U2129 (N_2129,N_1718,N_1802);
and U2130 (N_2130,N_1964,N_1709);
xnor U2131 (N_2131,N_1747,N_1876);
nand U2132 (N_2132,N_1570,N_1764);
or U2133 (N_2133,N_1681,N_1656);
xnor U2134 (N_2134,N_1908,N_1816);
nand U2135 (N_2135,N_1606,N_1890);
and U2136 (N_2136,N_1985,N_1810);
or U2137 (N_2137,N_1701,N_1827);
nor U2138 (N_2138,N_1680,N_1758);
and U2139 (N_2139,N_1775,N_1585);
nand U2140 (N_2140,N_1662,N_1868);
nor U2141 (N_2141,N_1965,N_1817);
or U2142 (N_2142,N_1854,N_1700);
xor U2143 (N_2143,N_1608,N_1990);
or U2144 (N_2144,N_1878,N_1567);
nand U2145 (N_2145,N_1831,N_1877);
and U2146 (N_2146,N_1752,N_1545);
nor U2147 (N_2147,N_1650,N_1509);
nor U2148 (N_2148,N_1577,N_1532);
nor U2149 (N_2149,N_1951,N_1771);
nand U2150 (N_2150,N_1549,N_1666);
nand U2151 (N_2151,N_1841,N_1795);
nor U2152 (N_2152,N_1703,N_1922);
or U2153 (N_2153,N_1711,N_1799);
nor U2154 (N_2154,N_1932,N_1623);
nand U2155 (N_2155,N_1755,N_1865);
nand U2156 (N_2156,N_1760,N_1954);
and U2157 (N_2157,N_1660,N_1852);
and U2158 (N_2158,N_1683,N_1941);
xor U2159 (N_2159,N_1687,N_1745);
nand U2160 (N_2160,N_1982,N_1673);
or U2161 (N_2161,N_1949,N_1573);
or U2162 (N_2162,N_1905,N_1675);
nand U2163 (N_2163,N_1520,N_1961);
nor U2164 (N_2164,N_1630,N_1507);
or U2165 (N_2165,N_1589,N_1900);
or U2166 (N_2166,N_1942,N_1525);
xor U2167 (N_2167,N_1632,N_1847);
nor U2168 (N_2168,N_1785,N_1667);
or U2169 (N_2169,N_1881,N_1625);
xnor U2170 (N_2170,N_1694,N_1768);
xnor U2171 (N_2171,N_1661,N_1776);
nand U2172 (N_2172,N_1790,N_1506);
nor U2173 (N_2173,N_1991,N_1819);
nand U2174 (N_2174,N_1605,N_1791);
xnor U2175 (N_2175,N_1926,N_1728);
and U2176 (N_2176,N_1733,N_1767);
nand U2177 (N_2177,N_1983,N_1753);
xor U2178 (N_2178,N_1998,N_1927);
nand U2179 (N_2179,N_1642,N_1537);
nand U2180 (N_2180,N_1921,N_1719);
nor U2181 (N_2181,N_1564,N_1575);
nor U2182 (N_2182,N_1678,N_1769);
nand U2183 (N_2183,N_1832,N_1858);
xnor U2184 (N_2184,N_1533,N_1979);
and U2185 (N_2185,N_1702,N_1693);
nand U2186 (N_2186,N_1633,N_1510);
nor U2187 (N_2187,N_1934,N_1935);
or U2188 (N_2188,N_1627,N_1880);
xor U2189 (N_2189,N_1722,N_1796);
nand U2190 (N_2190,N_1923,N_1913);
nor U2191 (N_2191,N_1538,N_1653);
nand U2192 (N_2192,N_1945,N_1515);
xnor U2193 (N_2193,N_1903,N_1818);
and U2194 (N_2194,N_1788,N_1748);
nand U2195 (N_2195,N_1727,N_1646);
or U2196 (N_2196,N_1872,N_1609);
and U2197 (N_2197,N_1599,N_1851);
nor U2198 (N_2198,N_1959,N_1829);
nand U2199 (N_2199,N_1674,N_1824);
nor U2200 (N_2200,N_1969,N_1582);
nand U2201 (N_2201,N_1713,N_1894);
or U2202 (N_2202,N_1759,N_1975);
nand U2203 (N_2203,N_1821,N_1987);
or U2204 (N_2204,N_1902,N_1780);
nor U2205 (N_2205,N_1522,N_1614);
nor U2206 (N_2206,N_1911,N_1536);
nand U2207 (N_2207,N_1843,N_1523);
nor U2208 (N_2208,N_1765,N_1560);
nand U2209 (N_2209,N_1822,N_1895);
and U2210 (N_2210,N_1550,N_1519);
nor U2211 (N_2211,N_1524,N_1891);
or U2212 (N_2212,N_1809,N_1688);
and U2213 (N_2213,N_1899,N_1939);
nor U2214 (N_2214,N_1761,N_1928);
nand U2215 (N_2215,N_1628,N_1862);
nor U2216 (N_2216,N_1999,N_1708);
nand U2217 (N_2217,N_1604,N_1732);
and U2218 (N_2218,N_1717,N_1607);
nand U2219 (N_2219,N_1742,N_1857);
nand U2220 (N_2220,N_1826,N_1583);
nand U2221 (N_2221,N_1651,N_1511);
and U2222 (N_2222,N_1576,N_1981);
xnor U2223 (N_2223,N_1971,N_1741);
nor U2224 (N_2224,N_1736,N_1641);
xor U2225 (N_2225,N_1952,N_1989);
nand U2226 (N_2226,N_1984,N_1888);
or U2227 (N_2227,N_1947,N_1500);
nand U2228 (N_2228,N_1861,N_1963);
and U2229 (N_2229,N_1615,N_1910);
or U2230 (N_2230,N_1957,N_1930);
nor U2231 (N_2231,N_1596,N_1746);
nor U2232 (N_2232,N_1631,N_1658);
and U2233 (N_2233,N_1715,N_1860);
or U2234 (N_2234,N_1552,N_1813);
nand U2235 (N_2235,N_1677,N_1610);
xnor U2236 (N_2236,N_1655,N_1676);
or U2237 (N_2237,N_1786,N_1534);
or U2238 (N_2238,N_1671,N_1505);
and U2239 (N_2239,N_1572,N_1698);
and U2240 (N_2240,N_1970,N_1588);
nor U2241 (N_2241,N_1586,N_1685);
and U2242 (N_2242,N_1937,N_1738);
xor U2243 (N_2243,N_1806,N_1624);
nor U2244 (N_2244,N_1647,N_1512);
or U2245 (N_2245,N_1803,N_1682);
and U2246 (N_2246,N_1994,N_1879);
xnor U2247 (N_2247,N_1705,N_1830);
or U2248 (N_2248,N_1535,N_1734);
nand U2249 (N_2249,N_1779,N_1828);
nand U2250 (N_2250,N_1916,N_1763);
or U2251 (N_2251,N_1740,N_1859);
nand U2252 (N_2252,N_1928,N_1967);
nand U2253 (N_2253,N_1961,N_1699);
xor U2254 (N_2254,N_1918,N_1645);
and U2255 (N_2255,N_1604,N_1537);
and U2256 (N_2256,N_1577,N_1849);
nand U2257 (N_2257,N_1813,N_1625);
nand U2258 (N_2258,N_1725,N_1676);
xnor U2259 (N_2259,N_1979,N_1945);
and U2260 (N_2260,N_1889,N_1930);
nand U2261 (N_2261,N_1715,N_1833);
and U2262 (N_2262,N_1771,N_1539);
or U2263 (N_2263,N_1914,N_1770);
xor U2264 (N_2264,N_1696,N_1883);
and U2265 (N_2265,N_1945,N_1599);
nor U2266 (N_2266,N_1966,N_1582);
xor U2267 (N_2267,N_1993,N_1871);
xnor U2268 (N_2268,N_1565,N_1835);
nor U2269 (N_2269,N_1948,N_1916);
nand U2270 (N_2270,N_1961,N_1541);
nand U2271 (N_2271,N_1756,N_1895);
or U2272 (N_2272,N_1921,N_1800);
nor U2273 (N_2273,N_1817,N_1591);
or U2274 (N_2274,N_1704,N_1880);
xor U2275 (N_2275,N_1991,N_1623);
nor U2276 (N_2276,N_1970,N_1959);
and U2277 (N_2277,N_1629,N_1678);
nor U2278 (N_2278,N_1824,N_1864);
xnor U2279 (N_2279,N_1741,N_1706);
nor U2280 (N_2280,N_1975,N_1790);
nor U2281 (N_2281,N_1676,N_1589);
and U2282 (N_2282,N_1531,N_1928);
nor U2283 (N_2283,N_1801,N_1639);
nand U2284 (N_2284,N_1819,N_1713);
or U2285 (N_2285,N_1935,N_1835);
and U2286 (N_2286,N_1908,N_1803);
and U2287 (N_2287,N_1900,N_1777);
or U2288 (N_2288,N_1699,N_1636);
or U2289 (N_2289,N_1942,N_1880);
xor U2290 (N_2290,N_1728,N_1771);
or U2291 (N_2291,N_1972,N_1605);
or U2292 (N_2292,N_1627,N_1934);
nand U2293 (N_2293,N_1852,N_1688);
xnor U2294 (N_2294,N_1948,N_1808);
and U2295 (N_2295,N_1610,N_1694);
nand U2296 (N_2296,N_1918,N_1797);
nand U2297 (N_2297,N_1691,N_1710);
xor U2298 (N_2298,N_1651,N_1634);
nand U2299 (N_2299,N_1878,N_1623);
and U2300 (N_2300,N_1694,N_1540);
nor U2301 (N_2301,N_1758,N_1535);
nor U2302 (N_2302,N_1778,N_1813);
nand U2303 (N_2303,N_1943,N_1746);
nor U2304 (N_2304,N_1778,N_1636);
xnor U2305 (N_2305,N_1546,N_1698);
nor U2306 (N_2306,N_1766,N_1896);
nor U2307 (N_2307,N_1805,N_1643);
nand U2308 (N_2308,N_1966,N_1873);
nand U2309 (N_2309,N_1933,N_1892);
nor U2310 (N_2310,N_1719,N_1606);
and U2311 (N_2311,N_1693,N_1665);
nand U2312 (N_2312,N_1981,N_1600);
and U2313 (N_2313,N_1748,N_1735);
or U2314 (N_2314,N_1729,N_1683);
or U2315 (N_2315,N_1650,N_1649);
and U2316 (N_2316,N_1597,N_1839);
nor U2317 (N_2317,N_1539,N_1663);
or U2318 (N_2318,N_1516,N_1847);
nor U2319 (N_2319,N_1967,N_1708);
xnor U2320 (N_2320,N_1508,N_1847);
nand U2321 (N_2321,N_1980,N_1784);
nor U2322 (N_2322,N_1935,N_1531);
xnor U2323 (N_2323,N_1745,N_1610);
nor U2324 (N_2324,N_1944,N_1831);
and U2325 (N_2325,N_1993,N_1778);
and U2326 (N_2326,N_1900,N_1564);
or U2327 (N_2327,N_1946,N_1617);
nor U2328 (N_2328,N_1755,N_1820);
and U2329 (N_2329,N_1925,N_1993);
xor U2330 (N_2330,N_1550,N_1939);
xnor U2331 (N_2331,N_1660,N_1614);
nand U2332 (N_2332,N_1981,N_1974);
or U2333 (N_2333,N_1706,N_1990);
and U2334 (N_2334,N_1952,N_1825);
xor U2335 (N_2335,N_1637,N_1597);
xor U2336 (N_2336,N_1729,N_1951);
or U2337 (N_2337,N_1661,N_1782);
nor U2338 (N_2338,N_1664,N_1931);
or U2339 (N_2339,N_1575,N_1811);
xor U2340 (N_2340,N_1994,N_1527);
and U2341 (N_2341,N_1551,N_1984);
or U2342 (N_2342,N_1527,N_1568);
nor U2343 (N_2343,N_1712,N_1725);
xnor U2344 (N_2344,N_1865,N_1676);
xnor U2345 (N_2345,N_1628,N_1924);
xnor U2346 (N_2346,N_1642,N_1550);
and U2347 (N_2347,N_1867,N_1803);
nor U2348 (N_2348,N_1995,N_1909);
and U2349 (N_2349,N_1620,N_1509);
and U2350 (N_2350,N_1883,N_1690);
and U2351 (N_2351,N_1625,N_1908);
and U2352 (N_2352,N_1619,N_1835);
or U2353 (N_2353,N_1673,N_1771);
or U2354 (N_2354,N_1931,N_1732);
nor U2355 (N_2355,N_1848,N_1641);
and U2356 (N_2356,N_1533,N_1551);
or U2357 (N_2357,N_1763,N_1705);
or U2358 (N_2358,N_1723,N_1923);
nand U2359 (N_2359,N_1966,N_1820);
xor U2360 (N_2360,N_1612,N_1522);
nor U2361 (N_2361,N_1832,N_1838);
and U2362 (N_2362,N_1544,N_1583);
nor U2363 (N_2363,N_1658,N_1614);
or U2364 (N_2364,N_1680,N_1977);
nand U2365 (N_2365,N_1771,N_1908);
nor U2366 (N_2366,N_1573,N_1888);
nand U2367 (N_2367,N_1700,N_1906);
nor U2368 (N_2368,N_1798,N_1532);
and U2369 (N_2369,N_1672,N_1761);
and U2370 (N_2370,N_1834,N_1512);
xor U2371 (N_2371,N_1647,N_1988);
nand U2372 (N_2372,N_1817,N_1681);
or U2373 (N_2373,N_1957,N_1599);
or U2374 (N_2374,N_1960,N_1615);
and U2375 (N_2375,N_1673,N_1840);
nor U2376 (N_2376,N_1860,N_1719);
or U2377 (N_2377,N_1801,N_1897);
or U2378 (N_2378,N_1919,N_1708);
or U2379 (N_2379,N_1616,N_1738);
nor U2380 (N_2380,N_1761,N_1523);
and U2381 (N_2381,N_1837,N_1558);
xor U2382 (N_2382,N_1795,N_1611);
xnor U2383 (N_2383,N_1988,N_1812);
xor U2384 (N_2384,N_1587,N_1668);
nor U2385 (N_2385,N_1771,N_1779);
or U2386 (N_2386,N_1836,N_1851);
and U2387 (N_2387,N_1613,N_1872);
and U2388 (N_2388,N_1646,N_1906);
nor U2389 (N_2389,N_1690,N_1545);
or U2390 (N_2390,N_1649,N_1798);
and U2391 (N_2391,N_1741,N_1738);
and U2392 (N_2392,N_1522,N_1637);
nor U2393 (N_2393,N_1904,N_1821);
nand U2394 (N_2394,N_1557,N_1830);
or U2395 (N_2395,N_1707,N_1773);
nor U2396 (N_2396,N_1660,N_1929);
nand U2397 (N_2397,N_1772,N_1616);
or U2398 (N_2398,N_1539,N_1514);
and U2399 (N_2399,N_1637,N_1770);
nand U2400 (N_2400,N_1682,N_1542);
xor U2401 (N_2401,N_1855,N_1985);
nor U2402 (N_2402,N_1821,N_1901);
nand U2403 (N_2403,N_1837,N_1553);
nand U2404 (N_2404,N_1929,N_1607);
and U2405 (N_2405,N_1578,N_1984);
nand U2406 (N_2406,N_1751,N_1606);
or U2407 (N_2407,N_1556,N_1944);
xor U2408 (N_2408,N_1506,N_1641);
or U2409 (N_2409,N_1791,N_1758);
and U2410 (N_2410,N_1953,N_1721);
or U2411 (N_2411,N_1736,N_1861);
xnor U2412 (N_2412,N_1547,N_1950);
xor U2413 (N_2413,N_1838,N_1580);
or U2414 (N_2414,N_1670,N_1547);
nand U2415 (N_2415,N_1726,N_1962);
and U2416 (N_2416,N_1643,N_1629);
nand U2417 (N_2417,N_1518,N_1950);
or U2418 (N_2418,N_1567,N_1939);
nand U2419 (N_2419,N_1715,N_1542);
or U2420 (N_2420,N_1525,N_1724);
xnor U2421 (N_2421,N_1553,N_1545);
nor U2422 (N_2422,N_1983,N_1747);
nand U2423 (N_2423,N_1963,N_1951);
and U2424 (N_2424,N_1869,N_1866);
nand U2425 (N_2425,N_1569,N_1811);
and U2426 (N_2426,N_1956,N_1750);
nor U2427 (N_2427,N_1732,N_1651);
nand U2428 (N_2428,N_1643,N_1519);
or U2429 (N_2429,N_1828,N_1773);
nand U2430 (N_2430,N_1881,N_1556);
xor U2431 (N_2431,N_1652,N_1640);
xor U2432 (N_2432,N_1986,N_1911);
nand U2433 (N_2433,N_1804,N_1643);
xor U2434 (N_2434,N_1799,N_1816);
nand U2435 (N_2435,N_1506,N_1764);
nand U2436 (N_2436,N_1519,N_1807);
nand U2437 (N_2437,N_1874,N_1648);
xor U2438 (N_2438,N_1921,N_1914);
nand U2439 (N_2439,N_1637,N_1760);
or U2440 (N_2440,N_1660,N_1645);
nor U2441 (N_2441,N_1914,N_1831);
and U2442 (N_2442,N_1973,N_1706);
and U2443 (N_2443,N_1996,N_1773);
and U2444 (N_2444,N_1767,N_1905);
and U2445 (N_2445,N_1502,N_1676);
xnor U2446 (N_2446,N_1747,N_1885);
and U2447 (N_2447,N_1718,N_1897);
or U2448 (N_2448,N_1962,N_1697);
and U2449 (N_2449,N_1902,N_1746);
nor U2450 (N_2450,N_1702,N_1891);
nand U2451 (N_2451,N_1644,N_1839);
xnor U2452 (N_2452,N_1530,N_1576);
nand U2453 (N_2453,N_1942,N_1827);
nor U2454 (N_2454,N_1951,N_1594);
nor U2455 (N_2455,N_1650,N_1606);
nor U2456 (N_2456,N_1782,N_1792);
nor U2457 (N_2457,N_1595,N_1992);
nor U2458 (N_2458,N_1962,N_1883);
or U2459 (N_2459,N_1833,N_1606);
or U2460 (N_2460,N_1768,N_1624);
or U2461 (N_2461,N_1670,N_1740);
and U2462 (N_2462,N_1511,N_1661);
nand U2463 (N_2463,N_1506,N_1955);
xnor U2464 (N_2464,N_1507,N_1929);
xor U2465 (N_2465,N_1629,N_1844);
and U2466 (N_2466,N_1559,N_1851);
and U2467 (N_2467,N_1734,N_1759);
xor U2468 (N_2468,N_1792,N_1629);
or U2469 (N_2469,N_1832,N_1795);
and U2470 (N_2470,N_1793,N_1787);
nand U2471 (N_2471,N_1568,N_1544);
or U2472 (N_2472,N_1655,N_1548);
and U2473 (N_2473,N_1577,N_1653);
and U2474 (N_2474,N_1529,N_1681);
nand U2475 (N_2475,N_1955,N_1723);
and U2476 (N_2476,N_1902,N_1962);
nand U2477 (N_2477,N_1941,N_1981);
nor U2478 (N_2478,N_1696,N_1977);
and U2479 (N_2479,N_1753,N_1634);
and U2480 (N_2480,N_1674,N_1745);
or U2481 (N_2481,N_1959,N_1766);
nor U2482 (N_2482,N_1791,N_1589);
and U2483 (N_2483,N_1500,N_1815);
nor U2484 (N_2484,N_1914,N_1528);
nor U2485 (N_2485,N_1517,N_1880);
xor U2486 (N_2486,N_1554,N_1972);
nor U2487 (N_2487,N_1966,N_1713);
nor U2488 (N_2488,N_1991,N_1979);
xnor U2489 (N_2489,N_1989,N_1588);
xnor U2490 (N_2490,N_1734,N_1546);
and U2491 (N_2491,N_1868,N_1767);
and U2492 (N_2492,N_1752,N_1953);
and U2493 (N_2493,N_1841,N_1740);
and U2494 (N_2494,N_1668,N_1704);
or U2495 (N_2495,N_1864,N_1780);
and U2496 (N_2496,N_1504,N_1580);
or U2497 (N_2497,N_1672,N_1822);
nor U2498 (N_2498,N_1553,N_1527);
or U2499 (N_2499,N_1521,N_1925);
xnor U2500 (N_2500,N_2344,N_2499);
nor U2501 (N_2501,N_2417,N_2158);
and U2502 (N_2502,N_2465,N_2453);
or U2503 (N_2503,N_2123,N_2103);
nor U2504 (N_2504,N_2333,N_2423);
and U2505 (N_2505,N_2494,N_2044);
nor U2506 (N_2506,N_2434,N_2384);
and U2507 (N_2507,N_2173,N_2235);
xnor U2508 (N_2508,N_2051,N_2316);
xnor U2509 (N_2509,N_2137,N_2482);
or U2510 (N_2510,N_2127,N_2356);
and U2511 (N_2511,N_2155,N_2334);
nor U2512 (N_2512,N_2081,N_2397);
nor U2513 (N_2513,N_2476,N_2414);
nor U2514 (N_2514,N_2129,N_2086);
xnor U2515 (N_2515,N_2362,N_2363);
nand U2516 (N_2516,N_2447,N_2041);
and U2517 (N_2517,N_2445,N_2310);
xnor U2518 (N_2518,N_2217,N_2118);
nor U2519 (N_2519,N_2181,N_2105);
and U2520 (N_2520,N_2090,N_2004);
nand U2521 (N_2521,N_2026,N_2413);
nor U2522 (N_2522,N_2210,N_2134);
and U2523 (N_2523,N_2359,N_2467);
or U2524 (N_2524,N_2436,N_2422);
or U2525 (N_2525,N_2109,N_2046);
and U2526 (N_2526,N_2444,N_2163);
xor U2527 (N_2527,N_2115,N_2446);
and U2528 (N_2528,N_2291,N_2021);
or U2529 (N_2529,N_2062,N_2225);
nor U2530 (N_2530,N_2145,N_2393);
or U2531 (N_2531,N_2357,N_2429);
nand U2532 (N_2532,N_2212,N_2076);
xnor U2533 (N_2533,N_2039,N_2289);
or U2534 (N_2534,N_2151,N_2481);
or U2535 (N_2535,N_2084,N_2266);
nor U2536 (N_2536,N_2104,N_2143);
nor U2537 (N_2537,N_2247,N_2202);
or U2538 (N_2538,N_2042,N_2282);
nand U2539 (N_2539,N_2340,N_2029);
nand U2540 (N_2540,N_2207,N_2116);
xnor U2541 (N_2541,N_2443,N_2349);
nor U2542 (N_2542,N_2458,N_2322);
or U2543 (N_2543,N_2464,N_2365);
or U2544 (N_2544,N_2396,N_2477);
nand U2545 (N_2545,N_2036,N_2346);
and U2546 (N_2546,N_2126,N_2187);
nand U2547 (N_2547,N_2161,N_2440);
or U2548 (N_2548,N_2252,N_2017);
nor U2549 (N_2549,N_2050,N_2360);
nand U2550 (N_2550,N_2057,N_2321);
or U2551 (N_2551,N_2468,N_2069);
nor U2552 (N_2552,N_2470,N_2271);
nand U2553 (N_2553,N_2230,N_2475);
xor U2554 (N_2554,N_2408,N_2461);
xnor U2555 (N_2555,N_2338,N_2085);
nor U2556 (N_2556,N_2088,N_2154);
nor U2557 (N_2557,N_2011,N_2337);
and U2558 (N_2558,N_2174,N_2067);
or U2559 (N_2559,N_2001,N_2229);
nor U2560 (N_2560,N_2299,N_2263);
and U2561 (N_2561,N_2493,N_2121);
xnor U2562 (N_2562,N_2361,N_2265);
nor U2563 (N_2563,N_2401,N_2189);
nor U2564 (N_2564,N_2079,N_2025);
nand U2565 (N_2565,N_2111,N_2188);
xnor U2566 (N_2566,N_2466,N_2487);
xnor U2567 (N_2567,N_2166,N_2425);
or U2568 (N_2568,N_2028,N_2370);
xnor U2569 (N_2569,N_2073,N_2192);
xnor U2570 (N_2570,N_2403,N_2351);
xor U2571 (N_2571,N_2296,N_2033);
nand U2572 (N_2572,N_2182,N_2009);
xor U2573 (N_2573,N_2305,N_2054);
xor U2574 (N_2574,N_2018,N_2294);
or U2575 (N_2575,N_2373,N_2135);
or U2576 (N_2576,N_2313,N_2380);
xnor U2577 (N_2577,N_2022,N_2472);
or U2578 (N_2578,N_2378,N_2012);
nor U2579 (N_2579,N_2364,N_2221);
nor U2580 (N_2580,N_2175,N_2257);
nand U2581 (N_2581,N_2233,N_2261);
nor U2582 (N_2582,N_2099,N_2101);
or U2583 (N_2583,N_2259,N_2150);
nand U2584 (N_2584,N_2292,N_2483);
nor U2585 (N_2585,N_2387,N_2335);
nand U2586 (N_2586,N_2249,N_2120);
xnor U2587 (N_2587,N_2048,N_2319);
and U2588 (N_2588,N_2208,N_2255);
xor U2589 (N_2589,N_2285,N_2224);
and U2590 (N_2590,N_2075,N_2382);
and U2591 (N_2591,N_2317,N_2144);
or U2592 (N_2592,N_2110,N_2388);
xnor U2593 (N_2593,N_2002,N_2290);
and U2594 (N_2594,N_2179,N_2352);
nor U2595 (N_2595,N_2049,N_2418);
nand U2596 (N_2596,N_2377,N_2133);
and U2597 (N_2597,N_2180,N_2215);
xnor U2598 (N_2598,N_2139,N_2199);
xnor U2599 (N_2599,N_2368,N_2428);
nor U2600 (N_2600,N_2267,N_2309);
xor U2601 (N_2601,N_2375,N_2183);
or U2602 (N_2602,N_2391,N_2420);
or U2603 (N_2603,N_2456,N_2190);
or U2604 (N_2604,N_2204,N_2213);
or U2605 (N_2605,N_2325,N_2197);
and U2606 (N_2606,N_2131,N_2030);
xnor U2607 (N_2607,N_2201,N_2140);
and U2608 (N_2608,N_2395,N_2411);
nor U2609 (N_2609,N_2035,N_2308);
or U2610 (N_2610,N_2023,N_2037);
nor U2611 (N_2611,N_2089,N_2008);
nor U2612 (N_2612,N_2007,N_2329);
or U2613 (N_2613,N_2096,N_2303);
or U2614 (N_2614,N_2433,N_2191);
nand U2615 (N_2615,N_2078,N_2058);
and U2616 (N_2616,N_2430,N_2047);
nor U2617 (N_2617,N_2122,N_2250);
and U2618 (N_2618,N_2462,N_2353);
xor U2619 (N_2619,N_2124,N_2354);
xnor U2620 (N_2620,N_2318,N_2059);
or U2621 (N_2621,N_2307,N_2093);
nand U2622 (N_2622,N_2358,N_2306);
and U2623 (N_2623,N_2312,N_2248);
nor U2624 (N_2624,N_2372,N_2068);
nand U2625 (N_2625,N_2478,N_2237);
or U2626 (N_2626,N_2284,N_2152);
and U2627 (N_2627,N_2273,N_2060);
nor U2628 (N_2628,N_2167,N_2157);
xnor U2629 (N_2629,N_2106,N_2449);
nor U2630 (N_2630,N_2209,N_2495);
nand U2631 (N_2631,N_2203,N_2366);
nor U2632 (N_2632,N_2473,N_2490);
nand U2633 (N_2633,N_2463,N_2302);
nor U2634 (N_2634,N_2342,N_2184);
nor U2635 (N_2635,N_2256,N_2343);
and U2636 (N_2636,N_2170,N_2112);
and U2637 (N_2637,N_2496,N_2113);
and U2638 (N_2638,N_2064,N_2024);
and U2639 (N_2639,N_2386,N_2206);
or U2640 (N_2640,N_2402,N_2232);
xnor U2641 (N_2641,N_2239,N_2339);
nand U2642 (N_2642,N_2226,N_2485);
nor U2643 (N_2643,N_2066,N_2072);
nand U2644 (N_2644,N_2474,N_2459);
nand U2645 (N_2645,N_2159,N_2092);
nor U2646 (N_2646,N_2277,N_2399);
nor U2647 (N_2647,N_2274,N_2260);
and U2648 (N_2648,N_2400,N_2141);
xnor U2649 (N_2649,N_2063,N_2293);
or U2650 (N_2650,N_2389,N_2435);
nand U2651 (N_2651,N_2003,N_2095);
and U2652 (N_2652,N_2406,N_2398);
and U2653 (N_2653,N_2091,N_2034);
nand U2654 (N_2654,N_2331,N_2176);
xor U2655 (N_2655,N_2350,N_2419);
xor U2656 (N_2656,N_2253,N_2330);
xor U2657 (N_2657,N_2421,N_2214);
and U2658 (N_2658,N_2077,N_2304);
and U2659 (N_2659,N_2489,N_2392);
nand U2660 (N_2660,N_2015,N_2448);
and U2661 (N_2661,N_2246,N_2369);
nand U2662 (N_2662,N_2374,N_2243);
nor U2663 (N_2663,N_2032,N_2000);
nor U2664 (N_2664,N_2149,N_2320);
xor U2665 (N_2665,N_2279,N_2222);
nand U2666 (N_2666,N_2497,N_2245);
nand U2667 (N_2667,N_2052,N_2196);
or U2668 (N_2668,N_2381,N_2227);
or U2669 (N_2669,N_2005,N_2486);
nor U2670 (N_2670,N_2371,N_2231);
nand U2671 (N_2671,N_2480,N_2178);
nand U2672 (N_2672,N_2080,N_2238);
xnor U2673 (N_2673,N_2027,N_2415);
or U2674 (N_2674,N_2390,N_2347);
or U2675 (N_2675,N_2241,N_2488);
nor U2676 (N_2676,N_2244,N_2484);
or U2677 (N_2677,N_2171,N_2138);
or U2678 (N_2678,N_2451,N_2327);
or U2679 (N_2679,N_2288,N_2427);
xnor U2680 (N_2680,N_2177,N_2441);
xor U2681 (N_2681,N_2328,N_2454);
nor U2682 (N_2682,N_2471,N_2114);
or U2683 (N_2683,N_2168,N_2438);
nor U2684 (N_2684,N_2268,N_2376);
or U2685 (N_2685,N_2125,N_2219);
nand U2686 (N_2686,N_2460,N_2045);
nand U2687 (N_2687,N_2269,N_2083);
or U2688 (N_2688,N_2195,N_2275);
or U2689 (N_2689,N_2194,N_2010);
or U2690 (N_2690,N_2070,N_2479);
nand U2691 (N_2691,N_2053,N_2272);
nand U2692 (N_2692,N_2457,N_2348);
and U2693 (N_2693,N_2492,N_2142);
nand U2694 (N_2694,N_2205,N_2450);
and U2695 (N_2695,N_2262,N_2014);
or U2696 (N_2696,N_2102,N_2297);
xor U2697 (N_2697,N_2146,N_2040);
nor U2698 (N_2698,N_2251,N_2065);
nor U2699 (N_2699,N_2276,N_2185);
or U2700 (N_2700,N_2228,N_2281);
nand U2701 (N_2701,N_2038,N_2278);
nand U2702 (N_2702,N_2469,N_2452);
or U2703 (N_2703,N_2006,N_2407);
and U2704 (N_2704,N_2172,N_2431);
and U2705 (N_2705,N_2074,N_2404);
nor U2706 (N_2706,N_2165,N_2162);
nand U2707 (N_2707,N_2383,N_2491);
or U2708 (N_2708,N_2128,N_2198);
or U2709 (N_2709,N_2314,N_2424);
or U2710 (N_2710,N_2218,N_2055);
or U2711 (N_2711,N_2061,N_2132);
or U2712 (N_2712,N_2336,N_2223);
or U2713 (N_2713,N_2020,N_2416);
and U2714 (N_2714,N_2432,N_2286);
or U2715 (N_2715,N_2119,N_2379);
or U2716 (N_2716,N_2410,N_2016);
nor U2717 (N_2717,N_2130,N_2097);
nor U2718 (N_2718,N_2056,N_2148);
or U2719 (N_2719,N_2200,N_2442);
and U2720 (N_2720,N_2169,N_2394);
nor U2721 (N_2721,N_2409,N_2298);
nand U2722 (N_2722,N_2355,N_2098);
nor U2723 (N_2723,N_2280,N_2283);
nand U2724 (N_2724,N_2367,N_2412);
and U2725 (N_2725,N_2071,N_2117);
nand U2726 (N_2726,N_2236,N_2147);
xnor U2727 (N_2727,N_2405,N_2455);
and U2728 (N_2728,N_2254,N_2100);
xor U2729 (N_2729,N_2240,N_2136);
and U2730 (N_2730,N_2295,N_2094);
nor U2731 (N_2731,N_2164,N_2326);
nor U2732 (N_2732,N_2220,N_2270);
or U2733 (N_2733,N_2019,N_2082);
nand U2734 (N_2734,N_2301,N_2216);
and U2735 (N_2735,N_2345,N_2156);
and U2736 (N_2736,N_2323,N_2341);
nand U2737 (N_2737,N_2211,N_2258);
nand U2738 (N_2738,N_2264,N_2031);
and U2739 (N_2739,N_2426,N_2385);
and U2740 (N_2740,N_2439,N_2332);
nand U2741 (N_2741,N_2107,N_2242);
or U2742 (N_2742,N_2153,N_2013);
or U2743 (N_2743,N_2315,N_2108);
xor U2744 (N_2744,N_2287,N_2437);
or U2745 (N_2745,N_2193,N_2498);
or U2746 (N_2746,N_2087,N_2234);
xnor U2747 (N_2747,N_2186,N_2311);
xor U2748 (N_2748,N_2043,N_2300);
xnor U2749 (N_2749,N_2160,N_2324);
and U2750 (N_2750,N_2212,N_2492);
xor U2751 (N_2751,N_2098,N_2125);
or U2752 (N_2752,N_2433,N_2093);
xor U2753 (N_2753,N_2371,N_2223);
and U2754 (N_2754,N_2293,N_2254);
xor U2755 (N_2755,N_2423,N_2087);
and U2756 (N_2756,N_2045,N_2228);
or U2757 (N_2757,N_2198,N_2242);
xor U2758 (N_2758,N_2358,N_2186);
nand U2759 (N_2759,N_2306,N_2075);
nand U2760 (N_2760,N_2041,N_2423);
or U2761 (N_2761,N_2262,N_2439);
and U2762 (N_2762,N_2342,N_2206);
xnor U2763 (N_2763,N_2383,N_2025);
xor U2764 (N_2764,N_2353,N_2461);
xnor U2765 (N_2765,N_2395,N_2200);
xnor U2766 (N_2766,N_2158,N_2489);
and U2767 (N_2767,N_2363,N_2167);
nor U2768 (N_2768,N_2023,N_2403);
or U2769 (N_2769,N_2490,N_2167);
xnor U2770 (N_2770,N_2201,N_2288);
xnor U2771 (N_2771,N_2040,N_2435);
nor U2772 (N_2772,N_2293,N_2104);
nand U2773 (N_2773,N_2135,N_2224);
and U2774 (N_2774,N_2064,N_2475);
and U2775 (N_2775,N_2478,N_2253);
and U2776 (N_2776,N_2349,N_2347);
xnor U2777 (N_2777,N_2399,N_2430);
nor U2778 (N_2778,N_2104,N_2394);
nand U2779 (N_2779,N_2463,N_2143);
nor U2780 (N_2780,N_2292,N_2375);
nor U2781 (N_2781,N_2073,N_2128);
or U2782 (N_2782,N_2088,N_2211);
xor U2783 (N_2783,N_2366,N_2218);
nor U2784 (N_2784,N_2144,N_2251);
nand U2785 (N_2785,N_2494,N_2245);
nand U2786 (N_2786,N_2139,N_2131);
and U2787 (N_2787,N_2112,N_2185);
nand U2788 (N_2788,N_2220,N_2151);
nand U2789 (N_2789,N_2167,N_2122);
or U2790 (N_2790,N_2366,N_2126);
nand U2791 (N_2791,N_2192,N_2486);
and U2792 (N_2792,N_2152,N_2343);
or U2793 (N_2793,N_2342,N_2077);
xnor U2794 (N_2794,N_2498,N_2022);
or U2795 (N_2795,N_2254,N_2487);
nor U2796 (N_2796,N_2283,N_2183);
or U2797 (N_2797,N_2083,N_2490);
and U2798 (N_2798,N_2347,N_2372);
nor U2799 (N_2799,N_2234,N_2040);
nand U2800 (N_2800,N_2218,N_2388);
nand U2801 (N_2801,N_2175,N_2267);
or U2802 (N_2802,N_2250,N_2266);
xnor U2803 (N_2803,N_2040,N_2093);
nor U2804 (N_2804,N_2260,N_2277);
and U2805 (N_2805,N_2314,N_2285);
or U2806 (N_2806,N_2138,N_2179);
nand U2807 (N_2807,N_2236,N_2053);
nand U2808 (N_2808,N_2174,N_2204);
nor U2809 (N_2809,N_2006,N_2041);
or U2810 (N_2810,N_2350,N_2325);
or U2811 (N_2811,N_2279,N_2158);
xor U2812 (N_2812,N_2111,N_2490);
and U2813 (N_2813,N_2462,N_2207);
and U2814 (N_2814,N_2112,N_2320);
and U2815 (N_2815,N_2142,N_2464);
or U2816 (N_2816,N_2194,N_2245);
nand U2817 (N_2817,N_2191,N_2448);
nor U2818 (N_2818,N_2468,N_2295);
xor U2819 (N_2819,N_2052,N_2176);
nor U2820 (N_2820,N_2077,N_2467);
and U2821 (N_2821,N_2475,N_2350);
nand U2822 (N_2822,N_2007,N_2278);
xor U2823 (N_2823,N_2487,N_2460);
nand U2824 (N_2824,N_2272,N_2329);
and U2825 (N_2825,N_2106,N_2397);
or U2826 (N_2826,N_2036,N_2403);
nand U2827 (N_2827,N_2013,N_2269);
nand U2828 (N_2828,N_2379,N_2166);
or U2829 (N_2829,N_2220,N_2211);
nand U2830 (N_2830,N_2390,N_2326);
nand U2831 (N_2831,N_2302,N_2362);
nor U2832 (N_2832,N_2409,N_2471);
nor U2833 (N_2833,N_2295,N_2320);
nand U2834 (N_2834,N_2179,N_2025);
and U2835 (N_2835,N_2232,N_2025);
nor U2836 (N_2836,N_2127,N_2007);
or U2837 (N_2837,N_2164,N_2400);
or U2838 (N_2838,N_2299,N_2435);
or U2839 (N_2839,N_2208,N_2014);
or U2840 (N_2840,N_2380,N_2034);
nand U2841 (N_2841,N_2350,N_2473);
nand U2842 (N_2842,N_2202,N_2104);
nor U2843 (N_2843,N_2017,N_2493);
nand U2844 (N_2844,N_2036,N_2421);
and U2845 (N_2845,N_2430,N_2423);
or U2846 (N_2846,N_2480,N_2123);
nand U2847 (N_2847,N_2496,N_2308);
xor U2848 (N_2848,N_2053,N_2467);
nand U2849 (N_2849,N_2106,N_2359);
nor U2850 (N_2850,N_2140,N_2389);
xnor U2851 (N_2851,N_2059,N_2274);
xnor U2852 (N_2852,N_2081,N_2286);
nor U2853 (N_2853,N_2174,N_2411);
xor U2854 (N_2854,N_2199,N_2248);
or U2855 (N_2855,N_2188,N_2465);
nand U2856 (N_2856,N_2078,N_2295);
xor U2857 (N_2857,N_2351,N_2407);
nand U2858 (N_2858,N_2004,N_2001);
nand U2859 (N_2859,N_2485,N_2483);
nor U2860 (N_2860,N_2428,N_2158);
nor U2861 (N_2861,N_2189,N_2431);
and U2862 (N_2862,N_2062,N_2280);
nor U2863 (N_2863,N_2387,N_2110);
or U2864 (N_2864,N_2391,N_2213);
nor U2865 (N_2865,N_2308,N_2263);
nor U2866 (N_2866,N_2355,N_2498);
or U2867 (N_2867,N_2374,N_2163);
xor U2868 (N_2868,N_2276,N_2308);
nand U2869 (N_2869,N_2035,N_2031);
or U2870 (N_2870,N_2038,N_2330);
nand U2871 (N_2871,N_2313,N_2478);
nor U2872 (N_2872,N_2292,N_2222);
nand U2873 (N_2873,N_2379,N_2326);
nand U2874 (N_2874,N_2341,N_2140);
nand U2875 (N_2875,N_2263,N_2480);
nor U2876 (N_2876,N_2490,N_2197);
and U2877 (N_2877,N_2234,N_2208);
nor U2878 (N_2878,N_2030,N_2090);
and U2879 (N_2879,N_2274,N_2322);
nand U2880 (N_2880,N_2208,N_2085);
nor U2881 (N_2881,N_2322,N_2212);
and U2882 (N_2882,N_2192,N_2419);
nand U2883 (N_2883,N_2265,N_2494);
nor U2884 (N_2884,N_2207,N_2033);
xnor U2885 (N_2885,N_2301,N_2123);
xor U2886 (N_2886,N_2497,N_2060);
nand U2887 (N_2887,N_2499,N_2440);
nand U2888 (N_2888,N_2239,N_2428);
nand U2889 (N_2889,N_2111,N_2081);
xnor U2890 (N_2890,N_2213,N_2453);
or U2891 (N_2891,N_2344,N_2486);
xnor U2892 (N_2892,N_2080,N_2474);
xor U2893 (N_2893,N_2493,N_2085);
xor U2894 (N_2894,N_2116,N_2468);
nor U2895 (N_2895,N_2349,N_2303);
or U2896 (N_2896,N_2437,N_2477);
or U2897 (N_2897,N_2429,N_2393);
xnor U2898 (N_2898,N_2428,N_2232);
and U2899 (N_2899,N_2470,N_2324);
and U2900 (N_2900,N_2465,N_2494);
nand U2901 (N_2901,N_2368,N_2430);
xor U2902 (N_2902,N_2152,N_2491);
and U2903 (N_2903,N_2355,N_2229);
nor U2904 (N_2904,N_2147,N_2055);
nor U2905 (N_2905,N_2466,N_2218);
or U2906 (N_2906,N_2033,N_2066);
and U2907 (N_2907,N_2372,N_2456);
and U2908 (N_2908,N_2309,N_2126);
or U2909 (N_2909,N_2252,N_2161);
nand U2910 (N_2910,N_2210,N_2258);
nand U2911 (N_2911,N_2017,N_2266);
or U2912 (N_2912,N_2182,N_2293);
or U2913 (N_2913,N_2005,N_2469);
or U2914 (N_2914,N_2334,N_2495);
nand U2915 (N_2915,N_2230,N_2416);
nand U2916 (N_2916,N_2261,N_2234);
xnor U2917 (N_2917,N_2073,N_2325);
xor U2918 (N_2918,N_2140,N_2460);
xnor U2919 (N_2919,N_2120,N_2280);
or U2920 (N_2920,N_2002,N_2035);
nand U2921 (N_2921,N_2349,N_2077);
and U2922 (N_2922,N_2103,N_2325);
xnor U2923 (N_2923,N_2270,N_2266);
and U2924 (N_2924,N_2383,N_2086);
or U2925 (N_2925,N_2143,N_2137);
nand U2926 (N_2926,N_2205,N_2053);
or U2927 (N_2927,N_2326,N_2037);
nand U2928 (N_2928,N_2159,N_2062);
nor U2929 (N_2929,N_2248,N_2066);
nand U2930 (N_2930,N_2397,N_2494);
xnor U2931 (N_2931,N_2289,N_2443);
nand U2932 (N_2932,N_2486,N_2075);
xnor U2933 (N_2933,N_2382,N_2414);
nor U2934 (N_2934,N_2240,N_2238);
or U2935 (N_2935,N_2130,N_2133);
nor U2936 (N_2936,N_2477,N_2344);
or U2937 (N_2937,N_2054,N_2483);
nor U2938 (N_2938,N_2301,N_2255);
or U2939 (N_2939,N_2238,N_2361);
and U2940 (N_2940,N_2145,N_2387);
xnor U2941 (N_2941,N_2422,N_2181);
or U2942 (N_2942,N_2046,N_2092);
nand U2943 (N_2943,N_2420,N_2388);
nor U2944 (N_2944,N_2021,N_2180);
and U2945 (N_2945,N_2060,N_2206);
nand U2946 (N_2946,N_2217,N_2133);
nand U2947 (N_2947,N_2080,N_2497);
or U2948 (N_2948,N_2076,N_2456);
nand U2949 (N_2949,N_2498,N_2326);
or U2950 (N_2950,N_2131,N_2390);
xnor U2951 (N_2951,N_2152,N_2115);
xnor U2952 (N_2952,N_2328,N_2352);
nand U2953 (N_2953,N_2106,N_2060);
or U2954 (N_2954,N_2469,N_2003);
xnor U2955 (N_2955,N_2418,N_2313);
nor U2956 (N_2956,N_2468,N_2129);
xor U2957 (N_2957,N_2292,N_2341);
or U2958 (N_2958,N_2108,N_2198);
nor U2959 (N_2959,N_2134,N_2096);
nand U2960 (N_2960,N_2245,N_2221);
or U2961 (N_2961,N_2090,N_2064);
xor U2962 (N_2962,N_2353,N_2364);
and U2963 (N_2963,N_2289,N_2009);
and U2964 (N_2964,N_2331,N_2174);
nand U2965 (N_2965,N_2191,N_2251);
nand U2966 (N_2966,N_2335,N_2449);
nand U2967 (N_2967,N_2005,N_2140);
nand U2968 (N_2968,N_2015,N_2291);
nand U2969 (N_2969,N_2468,N_2435);
nor U2970 (N_2970,N_2190,N_2432);
xor U2971 (N_2971,N_2074,N_2000);
or U2972 (N_2972,N_2431,N_2038);
nor U2973 (N_2973,N_2286,N_2252);
xor U2974 (N_2974,N_2190,N_2117);
and U2975 (N_2975,N_2119,N_2029);
xor U2976 (N_2976,N_2186,N_2470);
or U2977 (N_2977,N_2360,N_2435);
and U2978 (N_2978,N_2465,N_2029);
xnor U2979 (N_2979,N_2047,N_2198);
nand U2980 (N_2980,N_2421,N_2318);
xor U2981 (N_2981,N_2098,N_2394);
and U2982 (N_2982,N_2103,N_2321);
nor U2983 (N_2983,N_2321,N_2054);
and U2984 (N_2984,N_2425,N_2223);
xnor U2985 (N_2985,N_2016,N_2144);
nand U2986 (N_2986,N_2239,N_2119);
xor U2987 (N_2987,N_2403,N_2301);
xnor U2988 (N_2988,N_2467,N_2408);
and U2989 (N_2989,N_2202,N_2313);
xor U2990 (N_2990,N_2229,N_2434);
nor U2991 (N_2991,N_2002,N_2072);
nor U2992 (N_2992,N_2200,N_2343);
and U2993 (N_2993,N_2068,N_2052);
or U2994 (N_2994,N_2478,N_2444);
or U2995 (N_2995,N_2215,N_2076);
xnor U2996 (N_2996,N_2238,N_2330);
xor U2997 (N_2997,N_2275,N_2238);
and U2998 (N_2998,N_2368,N_2350);
xnor U2999 (N_2999,N_2159,N_2410);
xor U3000 (N_3000,N_2740,N_2971);
nor U3001 (N_3001,N_2654,N_2894);
or U3002 (N_3002,N_2653,N_2684);
xor U3003 (N_3003,N_2915,N_2919);
or U3004 (N_3004,N_2949,N_2749);
nand U3005 (N_3005,N_2718,N_2590);
nand U3006 (N_3006,N_2627,N_2720);
xor U3007 (N_3007,N_2735,N_2665);
and U3008 (N_3008,N_2851,N_2522);
and U3009 (N_3009,N_2853,N_2933);
and U3010 (N_3010,N_2931,N_2719);
xnor U3011 (N_3011,N_2578,N_2875);
xor U3012 (N_3012,N_2662,N_2818);
and U3013 (N_3013,N_2605,N_2983);
nor U3014 (N_3014,N_2708,N_2961);
or U3015 (N_3015,N_2682,N_2612);
nor U3016 (N_3016,N_2688,N_2552);
nor U3017 (N_3017,N_2566,N_2955);
nand U3018 (N_3018,N_2643,N_2553);
nand U3019 (N_3019,N_2847,N_2988);
nor U3020 (N_3020,N_2531,N_2633);
nand U3021 (N_3021,N_2539,N_2850);
xnor U3022 (N_3022,N_2524,N_2788);
and U3023 (N_3023,N_2874,N_2517);
and U3024 (N_3024,N_2780,N_2699);
nand U3025 (N_3025,N_2577,N_2791);
nand U3026 (N_3026,N_2856,N_2686);
nor U3027 (N_3027,N_2794,N_2753);
and U3028 (N_3028,N_2506,N_2655);
xnor U3029 (N_3029,N_2816,N_2559);
and U3030 (N_3030,N_2690,N_2835);
xor U3031 (N_3031,N_2798,N_2587);
or U3032 (N_3032,N_2882,N_2770);
nor U3033 (N_3033,N_2683,N_2918);
nand U3034 (N_3034,N_2721,N_2696);
nand U3035 (N_3035,N_2765,N_2639);
xnor U3036 (N_3036,N_2839,N_2928);
nand U3037 (N_3037,N_2990,N_2636);
nand U3038 (N_3038,N_2731,N_2734);
and U3039 (N_3039,N_2622,N_2760);
xnor U3040 (N_3040,N_2940,N_2985);
or U3041 (N_3041,N_2953,N_2693);
or U3042 (N_3042,N_2711,N_2863);
nand U3043 (N_3043,N_2644,N_2806);
nor U3044 (N_3044,N_2664,N_2836);
and U3045 (N_3045,N_2715,N_2695);
nand U3046 (N_3046,N_2634,N_2810);
nor U3047 (N_3047,N_2526,N_2911);
and U3048 (N_3048,N_2595,N_2889);
nand U3049 (N_3049,N_2593,N_2807);
nand U3050 (N_3050,N_2676,N_2594);
nor U3051 (N_3051,N_2642,N_2698);
or U3052 (N_3052,N_2966,N_2814);
or U3053 (N_3053,N_2906,N_2635);
and U3054 (N_3054,N_2541,N_2892);
and U3055 (N_3055,N_2606,N_2581);
nand U3056 (N_3056,N_2588,N_2739);
xnor U3057 (N_3057,N_2782,N_2861);
nor U3058 (N_3058,N_2980,N_2529);
nor U3059 (N_3059,N_2755,N_2631);
or U3060 (N_3060,N_2849,N_2723);
nor U3061 (N_3061,N_2822,N_2573);
or U3062 (N_3062,N_2809,N_2557);
xor U3063 (N_3063,N_2832,N_2535);
xnor U3064 (N_3064,N_2771,N_2989);
xor U3065 (N_3065,N_2674,N_2502);
xor U3066 (N_3066,N_2870,N_2800);
nor U3067 (N_3067,N_2831,N_2925);
or U3068 (N_3068,N_2632,N_2617);
nand U3069 (N_3069,N_2834,N_2991);
or U3070 (N_3070,N_2840,N_2528);
xor U3071 (N_3071,N_2783,N_2886);
xnor U3072 (N_3072,N_2795,N_2694);
nand U3073 (N_3073,N_2689,N_2951);
nor U3074 (N_3074,N_2697,N_2970);
xor U3075 (N_3075,N_2545,N_2930);
xor U3076 (N_3076,N_2844,N_2724);
nand U3077 (N_3077,N_2738,N_2599);
and U3078 (N_3078,N_2984,N_2837);
or U3079 (N_3079,N_2867,N_2544);
nand U3080 (N_3080,N_2910,N_2993);
nand U3081 (N_3081,N_2946,N_2558);
or U3082 (N_3082,N_2941,N_2623);
nor U3083 (N_3083,N_2607,N_2754);
or U3084 (N_3084,N_2859,N_2999);
nor U3085 (N_3085,N_2732,N_2574);
xor U3086 (N_3086,N_2944,N_2895);
nor U3087 (N_3087,N_2979,N_2551);
nor U3088 (N_3088,N_2745,N_2757);
nand U3089 (N_3089,N_2939,N_2790);
nor U3090 (N_3090,N_2714,N_2898);
nand U3091 (N_3091,N_2967,N_2786);
xnor U3092 (N_3092,N_2519,N_2744);
and U3093 (N_3093,N_2878,N_2900);
and U3094 (N_3094,N_2602,N_2527);
or U3095 (N_3095,N_2725,N_2729);
nand U3096 (N_3096,N_2666,N_2704);
and U3097 (N_3097,N_2650,N_2521);
nor U3098 (N_3098,N_2647,N_2703);
and U3099 (N_3099,N_2848,N_2960);
or U3100 (N_3100,N_2625,N_2897);
or U3101 (N_3101,N_2546,N_2669);
and U3102 (N_3102,N_2842,N_2945);
nand U3103 (N_3103,N_2950,N_2920);
and U3104 (N_3104,N_2614,N_2518);
or U3105 (N_3105,N_2767,N_2978);
xnor U3106 (N_3106,N_2962,N_2513);
and U3107 (N_3107,N_2802,N_2808);
xnor U3108 (N_3108,N_2742,N_2883);
and U3109 (N_3109,N_2572,N_2803);
or U3110 (N_3110,N_2997,N_2768);
nor U3111 (N_3111,N_2764,N_2750);
nor U3112 (N_3112,N_2881,N_2514);
xnor U3113 (N_3113,N_2986,N_2620);
nor U3114 (N_3114,N_2854,N_2508);
nor U3115 (N_3115,N_2965,N_2903);
nor U3116 (N_3116,N_2926,N_2880);
nand U3117 (N_3117,N_2779,N_2968);
nand U3118 (N_3118,N_2909,N_2873);
nand U3119 (N_3119,N_2826,N_2678);
nand U3120 (N_3120,N_2793,N_2778);
nand U3121 (N_3121,N_2975,N_2976);
or U3122 (N_3122,N_2943,N_2923);
or U3123 (N_3123,N_2871,N_2741);
and U3124 (N_3124,N_2618,N_2685);
nor U3125 (N_3125,N_2523,N_2667);
nor U3126 (N_3126,N_2532,N_2902);
nand U3127 (N_3127,N_2512,N_2820);
nand U3128 (N_3128,N_2626,N_2656);
xor U3129 (N_3129,N_2759,N_2994);
or U3130 (N_3130,N_2564,N_2860);
and U3131 (N_3131,N_2638,N_2736);
and U3132 (N_3132,N_2710,N_2796);
or U3133 (N_3133,N_2954,N_2872);
and U3134 (N_3134,N_2582,N_2756);
xnor U3135 (N_3135,N_2579,N_2538);
nand U3136 (N_3136,N_2511,N_2821);
or U3137 (N_3137,N_2681,N_2964);
and U3138 (N_3138,N_2751,N_2784);
and U3139 (N_3139,N_2675,N_2733);
nand U3140 (N_3140,N_2973,N_2663);
nand U3141 (N_3141,N_2833,N_2503);
xnor U3142 (N_3142,N_2905,N_2974);
nand U3143 (N_3143,N_2701,N_2864);
nand U3144 (N_3144,N_2628,N_2716);
nor U3145 (N_3145,N_2922,N_2956);
nand U3146 (N_3146,N_2533,N_2937);
or U3147 (N_3147,N_2887,N_2713);
xnor U3148 (N_3148,N_2787,N_2830);
xor U3149 (N_3149,N_2841,N_2672);
xor U3150 (N_3150,N_2624,N_2640);
nand U3151 (N_3151,N_2769,N_2908);
and U3152 (N_3152,N_2547,N_2592);
nand U3153 (N_3153,N_2507,N_2712);
or U3154 (N_3154,N_2589,N_2917);
and U3155 (N_3155,N_2687,N_2890);
nand U3156 (N_3156,N_2657,N_2877);
xnor U3157 (N_3157,N_2537,N_2921);
xor U3158 (N_3158,N_2671,N_2758);
xnor U3159 (N_3159,N_2525,N_2510);
nor U3160 (N_3160,N_2691,N_2648);
nor U3161 (N_3161,N_2829,N_2825);
nand U3162 (N_3162,N_2747,N_2571);
or U3163 (N_3163,N_2661,N_2520);
xnor U3164 (N_3164,N_2865,N_2603);
nand U3165 (N_3165,N_2641,N_2629);
nor U3166 (N_3166,N_2613,N_2575);
nor U3167 (N_3167,N_2550,N_2846);
nor U3168 (N_3168,N_2637,N_2813);
or U3169 (N_3169,N_2598,N_2569);
and U3170 (N_3170,N_2743,N_2823);
nand U3171 (N_3171,N_2660,N_2789);
nand U3172 (N_3172,N_2862,N_2817);
xor U3173 (N_3173,N_2893,N_2540);
and U3174 (N_3174,N_2600,N_2737);
nand U3175 (N_3175,N_2912,N_2580);
xor U3176 (N_3176,N_2611,N_2762);
xnor U3177 (N_3177,N_2935,N_2885);
xnor U3178 (N_3178,N_2815,N_2728);
xor U3179 (N_3179,N_2549,N_2969);
xnor U3180 (N_3180,N_2799,N_2646);
or U3181 (N_3181,N_2709,N_2530);
nor U3182 (N_3182,N_2942,N_2774);
and U3183 (N_3183,N_2869,N_2659);
xnor U3184 (N_3184,N_2958,N_2619);
or U3185 (N_3185,N_2858,N_2500);
and U3186 (N_3186,N_2673,N_2972);
xnor U3187 (N_3187,N_2987,N_2722);
nand U3188 (N_3188,N_2630,N_2584);
nor U3189 (N_3189,N_2649,N_2932);
or U3190 (N_3190,N_2596,N_2568);
and U3191 (N_3191,N_2896,N_2957);
and U3192 (N_3192,N_2838,N_2763);
xnor U3193 (N_3193,N_2777,N_2706);
and U3194 (N_3194,N_2927,N_2766);
and U3195 (N_3195,N_2679,N_2761);
xor U3196 (N_3196,N_2801,N_2608);
nor U3197 (N_3197,N_2616,N_2717);
or U3198 (N_3198,N_2560,N_2509);
nor U3199 (N_3199,N_2785,N_2570);
or U3200 (N_3200,N_2901,N_2651);
and U3201 (N_3201,N_2947,N_2866);
or U3202 (N_3202,N_2585,N_2797);
xor U3203 (N_3203,N_2792,N_2899);
or U3204 (N_3204,N_2907,N_2977);
xor U3205 (N_3205,N_2879,N_2752);
or U3206 (N_3206,N_2852,N_2934);
or U3207 (N_3207,N_2888,N_2998);
or U3208 (N_3208,N_2705,N_2730);
or U3209 (N_3209,N_2548,N_2645);
nor U3210 (N_3210,N_2812,N_2811);
nor U3211 (N_3211,N_2982,N_2515);
xnor U3212 (N_3212,N_2563,N_2772);
nand U3213 (N_3213,N_2924,N_2707);
xor U3214 (N_3214,N_2534,N_2843);
xor U3215 (N_3215,N_2781,N_2501);
or U3216 (N_3216,N_2914,N_2658);
nand U3217 (N_3217,N_2819,N_2504);
nand U3218 (N_3218,N_2562,N_2857);
or U3219 (N_3219,N_2775,N_2604);
nand U3220 (N_3220,N_2543,N_2542);
xor U3221 (N_3221,N_2904,N_2776);
nand U3222 (N_3222,N_2996,N_2609);
nor U3223 (N_3223,N_2702,N_2959);
or U3224 (N_3224,N_2677,N_2748);
or U3225 (N_3225,N_2668,N_2938);
nor U3226 (N_3226,N_2929,N_2692);
nor U3227 (N_3227,N_2597,N_2845);
and U3228 (N_3228,N_2855,N_2948);
nand U3229 (N_3229,N_2913,N_2773);
and U3230 (N_3230,N_2621,N_2827);
and U3231 (N_3231,N_2583,N_2727);
or U3232 (N_3232,N_2554,N_2891);
xor U3233 (N_3233,N_2995,N_2936);
and U3234 (N_3234,N_2876,N_2567);
or U3235 (N_3235,N_2556,N_2615);
xnor U3236 (N_3236,N_2824,N_2670);
nand U3237 (N_3237,N_2981,N_2591);
nor U3238 (N_3238,N_2963,N_2700);
xor U3239 (N_3239,N_2565,N_2726);
nand U3240 (N_3240,N_2586,N_2516);
nor U3241 (N_3241,N_2601,N_2828);
or U3242 (N_3242,N_2868,N_2680);
xor U3243 (N_3243,N_2804,N_2952);
and U3244 (N_3244,N_2561,N_2884);
nand U3245 (N_3245,N_2805,N_2746);
or U3246 (N_3246,N_2916,N_2652);
xnor U3247 (N_3247,N_2992,N_2555);
nand U3248 (N_3248,N_2610,N_2505);
or U3249 (N_3249,N_2536,N_2576);
xor U3250 (N_3250,N_2683,N_2714);
nor U3251 (N_3251,N_2533,N_2930);
nor U3252 (N_3252,N_2629,N_2905);
nand U3253 (N_3253,N_2777,N_2538);
or U3254 (N_3254,N_2860,N_2683);
and U3255 (N_3255,N_2503,N_2934);
xnor U3256 (N_3256,N_2542,N_2944);
nand U3257 (N_3257,N_2626,N_2902);
and U3258 (N_3258,N_2539,N_2675);
xnor U3259 (N_3259,N_2917,N_2748);
and U3260 (N_3260,N_2617,N_2628);
nor U3261 (N_3261,N_2880,N_2555);
or U3262 (N_3262,N_2699,N_2616);
or U3263 (N_3263,N_2654,N_2586);
nand U3264 (N_3264,N_2874,N_2711);
or U3265 (N_3265,N_2823,N_2506);
nor U3266 (N_3266,N_2853,N_2976);
nor U3267 (N_3267,N_2666,N_2658);
xor U3268 (N_3268,N_2706,N_2759);
nor U3269 (N_3269,N_2778,N_2505);
nor U3270 (N_3270,N_2997,N_2922);
nor U3271 (N_3271,N_2508,N_2810);
xnor U3272 (N_3272,N_2517,N_2618);
or U3273 (N_3273,N_2504,N_2772);
xor U3274 (N_3274,N_2943,N_2588);
nor U3275 (N_3275,N_2747,N_2710);
nor U3276 (N_3276,N_2612,N_2520);
and U3277 (N_3277,N_2830,N_2979);
xor U3278 (N_3278,N_2529,N_2614);
and U3279 (N_3279,N_2820,N_2565);
xor U3280 (N_3280,N_2853,N_2543);
or U3281 (N_3281,N_2586,N_2751);
and U3282 (N_3282,N_2946,N_2533);
xnor U3283 (N_3283,N_2617,N_2535);
nor U3284 (N_3284,N_2994,N_2999);
and U3285 (N_3285,N_2647,N_2742);
nor U3286 (N_3286,N_2788,N_2913);
nand U3287 (N_3287,N_2708,N_2722);
xnor U3288 (N_3288,N_2606,N_2815);
and U3289 (N_3289,N_2638,N_2932);
and U3290 (N_3290,N_2899,N_2772);
nor U3291 (N_3291,N_2508,N_2891);
nand U3292 (N_3292,N_2755,N_2533);
and U3293 (N_3293,N_2892,N_2542);
nor U3294 (N_3294,N_2557,N_2774);
nand U3295 (N_3295,N_2655,N_2922);
and U3296 (N_3296,N_2996,N_2768);
or U3297 (N_3297,N_2836,N_2725);
or U3298 (N_3298,N_2798,N_2681);
or U3299 (N_3299,N_2537,N_2556);
xnor U3300 (N_3300,N_2937,N_2978);
and U3301 (N_3301,N_2875,N_2746);
xor U3302 (N_3302,N_2671,N_2797);
nand U3303 (N_3303,N_2515,N_2653);
xnor U3304 (N_3304,N_2588,N_2813);
xnor U3305 (N_3305,N_2948,N_2746);
nand U3306 (N_3306,N_2858,N_2602);
and U3307 (N_3307,N_2920,N_2802);
nand U3308 (N_3308,N_2776,N_2803);
and U3309 (N_3309,N_2845,N_2530);
nand U3310 (N_3310,N_2834,N_2704);
nor U3311 (N_3311,N_2952,N_2681);
and U3312 (N_3312,N_2505,N_2671);
or U3313 (N_3313,N_2802,N_2616);
or U3314 (N_3314,N_2508,N_2941);
nor U3315 (N_3315,N_2594,N_2628);
nor U3316 (N_3316,N_2512,N_2923);
and U3317 (N_3317,N_2774,N_2569);
xor U3318 (N_3318,N_2887,N_2742);
nand U3319 (N_3319,N_2566,N_2561);
nand U3320 (N_3320,N_2721,N_2609);
xor U3321 (N_3321,N_2698,N_2826);
nand U3322 (N_3322,N_2928,N_2915);
xor U3323 (N_3323,N_2658,N_2975);
and U3324 (N_3324,N_2844,N_2511);
or U3325 (N_3325,N_2541,N_2514);
and U3326 (N_3326,N_2578,N_2842);
or U3327 (N_3327,N_2988,N_2925);
or U3328 (N_3328,N_2817,N_2703);
or U3329 (N_3329,N_2506,N_2715);
nand U3330 (N_3330,N_2911,N_2635);
nor U3331 (N_3331,N_2858,N_2928);
or U3332 (N_3332,N_2763,N_2700);
nor U3333 (N_3333,N_2587,N_2654);
or U3334 (N_3334,N_2815,N_2628);
or U3335 (N_3335,N_2536,N_2758);
or U3336 (N_3336,N_2863,N_2816);
nor U3337 (N_3337,N_2858,N_2608);
xor U3338 (N_3338,N_2838,N_2793);
xor U3339 (N_3339,N_2661,N_2952);
xnor U3340 (N_3340,N_2964,N_2917);
nor U3341 (N_3341,N_2661,N_2586);
nand U3342 (N_3342,N_2793,N_2882);
and U3343 (N_3343,N_2699,N_2711);
nand U3344 (N_3344,N_2878,N_2908);
nor U3345 (N_3345,N_2593,N_2696);
xor U3346 (N_3346,N_2642,N_2701);
nand U3347 (N_3347,N_2909,N_2531);
and U3348 (N_3348,N_2916,N_2932);
xnor U3349 (N_3349,N_2938,N_2903);
or U3350 (N_3350,N_2536,N_2560);
nand U3351 (N_3351,N_2778,N_2992);
nor U3352 (N_3352,N_2745,N_2647);
or U3353 (N_3353,N_2507,N_2993);
and U3354 (N_3354,N_2944,N_2881);
and U3355 (N_3355,N_2571,N_2749);
or U3356 (N_3356,N_2503,N_2745);
nor U3357 (N_3357,N_2764,N_2756);
and U3358 (N_3358,N_2527,N_2585);
xor U3359 (N_3359,N_2713,N_2730);
xor U3360 (N_3360,N_2922,N_2844);
or U3361 (N_3361,N_2624,N_2675);
and U3362 (N_3362,N_2630,N_2914);
nand U3363 (N_3363,N_2689,N_2878);
nor U3364 (N_3364,N_2760,N_2915);
xor U3365 (N_3365,N_2899,N_2504);
xnor U3366 (N_3366,N_2847,N_2592);
xor U3367 (N_3367,N_2891,N_2875);
and U3368 (N_3368,N_2580,N_2864);
or U3369 (N_3369,N_2546,N_2588);
xnor U3370 (N_3370,N_2546,N_2748);
nand U3371 (N_3371,N_2847,N_2501);
and U3372 (N_3372,N_2966,N_2851);
and U3373 (N_3373,N_2617,N_2912);
nor U3374 (N_3374,N_2522,N_2810);
and U3375 (N_3375,N_2992,N_2604);
or U3376 (N_3376,N_2694,N_2869);
nor U3377 (N_3377,N_2960,N_2540);
xnor U3378 (N_3378,N_2587,N_2852);
or U3379 (N_3379,N_2840,N_2584);
nor U3380 (N_3380,N_2683,N_2949);
nor U3381 (N_3381,N_2516,N_2627);
nor U3382 (N_3382,N_2692,N_2610);
or U3383 (N_3383,N_2923,N_2639);
and U3384 (N_3384,N_2882,N_2992);
and U3385 (N_3385,N_2811,N_2802);
and U3386 (N_3386,N_2674,N_2836);
xnor U3387 (N_3387,N_2595,N_2860);
xor U3388 (N_3388,N_2578,N_2758);
xnor U3389 (N_3389,N_2789,N_2902);
or U3390 (N_3390,N_2711,N_2931);
or U3391 (N_3391,N_2841,N_2853);
and U3392 (N_3392,N_2602,N_2635);
nand U3393 (N_3393,N_2665,N_2747);
nor U3394 (N_3394,N_2628,N_2549);
and U3395 (N_3395,N_2949,N_2569);
or U3396 (N_3396,N_2754,N_2794);
nor U3397 (N_3397,N_2736,N_2576);
xnor U3398 (N_3398,N_2611,N_2941);
xor U3399 (N_3399,N_2906,N_2590);
nor U3400 (N_3400,N_2579,N_2567);
or U3401 (N_3401,N_2996,N_2614);
and U3402 (N_3402,N_2760,N_2972);
or U3403 (N_3403,N_2593,N_2642);
or U3404 (N_3404,N_2998,N_2765);
and U3405 (N_3405,N_2941,N_2972);
and U3406 (N_3406,N_2745,N_2790);
xnor U3407 (N_3407,N_2541,N_2968);
and U3408 (N_3408,N_2589,N_2948);
nor U3409 (N_3409,N_2585,N_2981);
nand U3410 (N_3410,N_2573,N_2944);
or U3411 (N_3411,N_2900,N_2672);
nand U3412 (N_3412,N_2683,N_2654);
xor U3413 (N_3413,N_2818,N_2890);
and U3414 (N_3414,N_2968,N_2518);
nor U3415 (N_3415,N_2883,N_2706);
nand U3416 (N_3416,N_2923,N_2725);
nand U3417 (N_3417,N_2809,N_2732);
and U3418 (N_3418,N_2905,N_2968);
xnor U3419 (N_3419,N_2884,N_2653);
nand U3420 (N_3420,N_2726,N_2782);
and U3421 (N_3421,N_2675,N_2533);
xor U3422 (N_3422,N_2694,N_2645);
and U3423 (N_3423,N_2543,N_2740);
nand U3424 (N_3424,N_2763,N_2831);
or U3425 (N_3425,N_2834,N_2551);
or U3426 (N_3426,N_2961,N_2678);
xor U3427 (N_3427,N_2708,N_2654);
nand U3428 (N_3428,N_2815,N_2769);
and U3429 (N_3429,N_2517,N_2697);
nor U3430 (N_3430,N_2875,N_2940);
nor U3431 (N_3431,N_2888,N_2605);
nor U3432 (N_3432,N_2622,N_2892);
and U3433 (N_3433,N_2791,N_2949);
or U3434 (N_3434,N_2797,N_2826);
nand U3435 (N_3435,N_2625,N_2781);
nor U3436 (N_3436,N_2560,N_2921);
and U3437 (N_3437,N_2898,N_2678);
nor U3438 (N_3438,N_2653,N_2942);
and U3439 (N_3439,N_2715,N_2789);
nor U3440 (N_3440,N_2769,N_2604);
and U3441 (N_3441,N_2600,N_2869);
nor U3442 (N_3442,N_2827,N_2747);
or U3443 (N_3443,N_2681,N_2715);
nor U3444 (N_3444,N_2520,N_2735);
nor U3445 (N_3445,N_2566,N_2702);
nand U3446 (N_3446,N_2888,N_2726);
nand U3447 (N_3447,N_2975,N_2548);
or U3448 (N_3448,N_2889,N_2695);
xnor U3449 (N_3449,N_2763,N_2508);
or U3450 (N_3450,N_2605,N_2515);
and U3451 (N_3451,N_2741,N_2730);
or U3452 (N_3452,N_2895,N_2654);
or U3453 (N_3453,N_2807,N_2818);
nor U3454 (N_3454,N_2742,N_2598);
nand U3455 (N_3455,N_2950,N_2762);
nor U3456 (N_3456,N_2677,N_2907);
and U3457 (N_3457,N_2633,N_2783);
xor U3458 (N_3458,N_2681,N_2705);
nor U3459 (N_3459,N_2765,N_2547);
nand U3460 (N_3460,N_2856,N_2831);
or U3461 (N_3461,N_2985,N_2528);
nand U3462 (N_3462,N_2997,N_2789);
nor U3463 (N_3463,N_2607,N_2627);
and U3464 (N_3464,N_2619,N_2661);
nor U3465 (N_3465,N_2558,N_2800);
nor U3466 (N_3466,N_2514,N_2977);
nand U3467 (N_3467,N_2690,N_2566);
xnor U3468 (N_3468,N_2785,N_2969);
and U3469 (N_3469,N_2823,N_2826);
nand U3470 (N_3470,N_2585,N_2548);
nand U3471 (N_3471,N_2534,N_2770);
or U3472 (N_3472,N_2973,N_2941);
and U3473 (N_3473,N_2927,N_2563);
or U3474 (N_3474,N_2551,N_2664);
nor U3475 (N_3475,N_2837,N_2948);
nor U3476 (N_3476,N_2599,N_2851);
and U3477 (N_3477,N_2804,N_2904);
nor U3478 (N_3478,N_2525,N_2535);
nor U3479 (N_3479,N_2916,N_2754);
xnor U3480 (N_3480,N_2600,N_2914);
xor U3481 (N_3481,N_2860,N_2713);
xnor U3482 (N_3482,N_2964,N_2816);
and U3483 (N_3483,N_2758,N_2977);
or U3484 (N_3484,N_2658,N_2549);
and U3485 (N_3485,N_2626,N_2736);
and U3486 (N_3486,N_2537,N_2591);
or U3487 (N_3487,N_2847,N_2540);
xor U3488 (N_3488,N_2594,N_2611);
xnor U3489 (N_3489,N_2838,N_2959);
nand U3490 (N_3490,N_2538,N_2762);
xor U3491 (N_3491,N_2759,N_2849);
or U3492 (N_3492,N_2890,N_2829);
and U3493 (N_3493,N_2671,N_2998);
nor U3494 (N_3494,N_2500,N_2681);
and U3495 (N_3495,N_2818,N_2605);
nand U3496 (N_3496,N_2926,N_2808);
and U3497 (N_3497,N_2995,N_2999);
and U3498 (N_3498,N_2953,N_2840);
nand U3499 (N_3499,N_2813,N_2948);
xor U3500 (N_3500,N_3106,N_3482);
or U3501 (N_3501,N_3046,N_3318);
or U3502 (N_3502,N_3494,N_3029);
xor U3503 (N_3503,N_3481,N_3126);
or U3504 (N_3504,N_3406,N_3157);
and U3505 (N_3505,N_3349,N_3411);
and U3506 (N_3506,N_3152,N_3112);
nand U3507 (N_3507,N_3465,N_3372);
nor U3508 (N_3508,N_3258,N_3288);
or U3509 (N_3509,N_3015,N_3385);
xor U3510 (N_3510,N_3345,N_3421);
nand U3511 (N_3511,N_3378,N_3223);
nand U3512 (N_3512,N_3386,N_3480);
and U3513 (N_3513,N_3061,N_3115);
nor U3514 (N_3514,N_3020,N_3243);
or U3515 (N_3515,N_3072,N_3151);
xor U3516 (N_3516,N_3442,N_3292);
or U3517 (N_3517,N_3099,N_3262);
nor U3518 (N_3518,N_3076,N_3323);
xnor U3519 (N_3519,N_3127,N_3149);
nor U3520 (N_3520,N_3159,N_3057);
and U3521 (N_3521,N_3321,N_3108);
nor U3522 (N_3522,N_3395,N_3373);
or U3523 (N_3523,N_3004,N_3211);
nand U3524 (N_3524,N_3478,N_3214);
or U3525 (N_3525,N_3281,N_3059);
or U3526 (N_3526,N_3003,N_3396);
nor U3527 (N_3527,N_3332,N_3013);
nor U3528 (N_3528,N_3233,N_3254);
xnor U3529 (N_3529,N_3484,N_3443);
nor U3530 (N_3530,N_3137,N_3350);
xnor U3531 (N_3531,N_3363,N_3206);
nand U3532 (N_3532,N_3241,N_3371);
nor U3533 (N_3533,N_3186,N_3178);
xnor U3534 (N_3534,N_3416,N_3270);
nand U3535 (N_3535,N_3111,N_3203);
or U3536 (N_3536,N_3040,N_3204);
or U3537 (N_3537,N_3242,N_3148);
nand U3538 (N_3538,N_3287,N_3256);
or U3539 (N_3539,N_3184,N_3437);
nand U3540 (N_3540,N_3239,N_3129);
xnor U3541 (N_3541,N_3294,N_3098);
or U3542 (N_3542,N_3348,N_3354);
and U3543 (N_3543,N_3387,N_3369);
nand U3544 (N_3544,N_3248,N_3028);
xor U3545 (N_3545,N_3268,N_3351);
nor U3546 (N_3546,N_3173,N_3325);
nand U3547 (N_3547,N_3271,N_3140);
xnor U3548 (N_3548,N_3198,N_3289);
nor U3549 (N_3549,N_3295,N_3107);
and U3550 (N_3550,N_3150,N_3327);
or U3551 (N_3551,N_3000,N_3026);
nand U3552 (N_3552,N_3410,N_3341);
nand U3553 (N_3553,N_3272,N_3412);
nor U3554 (N_3554,N_3417,N_3232);
nand U3555 (N_3555,N_3110,N_3430);
xor U3556 (N_3556,N_3449,N_3337);
nand U3557 (N_3557,N_3071,N_3364);
xnor U3558 (N_3558,N_3084,N_3380);
nand U3559 (N_3559,N_3477,N_3425);
nand U3560 (N_3560,N_3130,N_3238);
or U3561 (N_3561,N_3356,N_3212);
nand U3562 (N_3562,N_3264,N_3403);
and U3563 (N_3563,N_3456,N_3224);
or U3564 (N_3564,N_3097,N_3340);
nand U3565 (N_3565,N_3382,N_3170);
and U3566 (N_3566,N_3290,N_3301);
or U3567 (N_3567,N_3060,N_3329);
and U3568 (N_3568,N_3361,N_3434);
and U3569 (N_3569,N_3132,N_3119);
or U3570 (N_3570,N_3083,N_3428);
or U3571 (N_3571,N_3497,N_3285);
nand U3572 (N_3572,N_3078,N_3018);
nor U3573 (N_3573,N_3192,N_3296);
xor U3574 (N_3574,N_3101,N_3463);
and U3575 (N_3575,N_3392,N_3116);
and U3576 (N_3576,N_3236,N_3228);
xor U3577 (N_3577,N_3409,N_3063);
or U3578 (N_3578,N_3488,N_3440);
nor U3579 (N_3579,N_3278,N_3048);
xor U3580 (N_3580,N_3050,N_3429);
and U3581 (N_3581,N_3191,N_3436);
and U3582 (N_3582,N_3094,N_3035);
and U3583 (N_3583,N_3420,N_3310);
or U3584 (N_3584,N_3453,N_3388);
nor U3585 (N_3585,N_3491,N_3069);
nor U3586 (N_3586,N_3259,N_3397);
nor U3587 (N_3587,N_3495,N_3358);
nor U3588 (N_3588,N_3405,N_3165);
nor U3589 (N_3589,N_3041,N_3273);
xnor U3590 (N_3590,N_3324,N_3080);
nor U3591 (N_3591,N_3260,N_3374);
or U3592 (N_3592,N_3042,N_3213);
nand U3593 (N_3593,N_3001,N_3167);
nor U3594 (N_3594,N_3227,N_3008);
nor U3595 (N_3595,N_3304,N_3128);
or U3596 (N_3596,N_3316,N_3118);
or U3597 (N_3597,N_3085,N_3467);
or U3598 (N_3598,N_3024,N_3448);
or U3599 (N_3599,N_3011,N_3355);
or U3600 (N_3600,N_3022,N_3444);
and U3601 (N_3601,N_3333,N_3246);
nand U3602 (N_3602,N_3189,N_3401);
or U3603 (N_3603,N_3188,N_3230);
or U3604 (N_3604,N_3138,N_3210);
or U3605 (N_3605,N_3293,N_3314);
or U3606 (N_3606,N_3122,N_3217);
nand U3607 (N_3607,N_3394,N_3240);
xnor U3608 (N_3608,N_3431,N_3282);
and U3609 (N_3609,N_3313,N_3195);
nor U3610 (N_3610,N_3089,N_3114);
nor U3611 (N_3611,N_3253,N_3439);
nor U3612 (N_3612,N_3353,N_3461);
nand U3613 (N_3613,N_3091,N_3234);
or U3614 (N_3614,N_3124,N_3220);
and U3615 (N_3615,N_3190,N_3245);
and U3616 (N_3616,N_3381,N_3231);
xnor U3617 (N_3617,N_3133,N_3146);
nand U3618 (N_3618,N_3320,N_3215);
and U3619 (N_3619,N_3226,N_3031);
xnor U3620 (N_3620,N_3052,N_3322);
xnor U3621 (N_3621,N_3487,N_3056);
nand U3622 (N_3622,N_3051,N_3162);
and U3623 (N_3623,N_3427,N_3435);
xnor U3624 (N_3624,N_3261,N_3143);
and U3625 (N_3625,N_3187,N_3422);
and U3626 (N_3626,N_3460,N_3081);
or U3627 (N_3627,N_3023,N_3109);
nand U3628 (N_3628,N_3297,N_3441);
xor U3629 (N_3629,N_3413,N_3229);
xor U3630 (N_3630,N_3185,N_3144);
nor U3631 (N_3631,N_3312,N_3275);
nor U3632 (N_3632,N_3183,N_3326);
and U3633 (N_3633,N_3006,N_3362);
nor U3634 (N_3634,N_3389,N_3298);
and U3635 (N_3635,N_3202,N_3047);
nand U3636 (N_3636,N_3486,N_3038);
xor U3637 (N_3637,N_3342,N_3433);
and U3638 (N_3638,N_3193,N_3163);
or U3639 (N_3639,N_3344,N_3168);
xor U3640 (N_3640,N_3266,N_3464);
nand U3641 (N_3641,N_3307,N_3303);
nand U3642 (N_3642,N_3419,N_3036);
nand U3643 (N_3643,N_3113,N_3180);
xor U3644 (N_3644,N_3357,N_3462);
nand U3645 (N_3645,N_3007,N_3045);
xor U3646 (N_3646,N_3249,N_3086);
and U3647 (N_3647,N_3087,N_3336);
nand U3648 (N_3648,N_3483,N_3451);
or U3649 (N_3649,N_3062,N_3100);
nand U3650 (N_3650,N_3221,N_3077);
nand U3651 (N_3651,N_3383,N_3473);
or U3652 (N_3652,N_3402,N_3475);
or U3653 (N_3653,N_3237,N_3068);
nor U3654 (N_3654,N_3175,N_3390);
and U3655 (N_3655,N_3125,N_3088);
xnor U3656 (N_3656,N_3021,N_3141);
or U3657 (N_3657,N_3365,N_3166);
nand U3658 (N_3658,N_3331,N_3017);
nor U3659 (N_3659,N_3257,N_3315);
and U3660 (N_3660,N_3274,N_3010);
and U3661 (N_3661,N_3123,N_3492);
and U3662 (N_3662,N_3019,N_3252);
and U3663 (N_3663,N_3302,N_3103);
nor U3664 (N_3664,N_3445,N_3200);
or U3665 (N_3665,N_3267,N_3432);
xnor U3666 (N_3666,N_3454,N_3067);
nor U3667 (N_3667,N_3330,N_3276);
xnor U3668 (N_3668,N_3309,N_3027);
or U3669 (N_3669,N_3493,N_3219);
and U3670 (N_3670,N_3338,N_3407);
or U3671 (N_3671,N_3147,N_3096);
nand U3672 (N_3672,N_3426,N_3025);
nand U3673 (N_3673,N_3311,N_3197);
nor U3674 (N_3674,N_3093,N_3074);
nor U3675 (N_3675,N_3360,N_3391);
and U3676 (N_3676,N_3370,N_3205);
or U3677 (N_3677,N_3251,N_3247);
nor U3678 (N_3678,N_3044,N_3161);
and U3679 (N_3679,N_3105,N_3033);
nand U3680 (N_3680,N_3194,N_3136);
nand U3681 (N_3681,N_3037,N_3286);
nand U3682 (N_3682,N_3090,N_3255);
or U3683 (N_3683,N_3352,N_3196);
xnor U3684 (N_3684,N_3418,N_3414);
nand U3685 (N_3685,N_3334,N_3457);
and U3686 (N_3686,N_3468,N_3490);
nand U3687 (N_3687,N_3053,N_3277);
nand U3688 (N_3688,N_3176,N_3079);
xnor U3689 (N_3689,N_3469,N_3479);
nand U3690 (N_3690,N_3092,N_3135);
xnor U3691 (N_3691,N_3423,N_3472);
and U3692 (N_3692,N_3154,N_3102);
nor U3693 (N_3693,N_3346,N_3216);
or U3694 (N_3694,N_3030,N_3142);
or U3695 (N_3695,N_3209,N_3299);
nand U3696 (N_3696,N_3156,N_3343);
or U3697 (N_3697,N_3005,N_3174);
or U3698 (N_3698,N_3131,N_3012);
nor U3699 (N_3699,N_3408,N_3250);
nor U3700 (N_3700,N_3009,N_3235);
or U3701 (N_3701,N_3489,N_3179);
xnor U3702 (N_3702,N_3446,N_3308);
nor U3703 (N_3703,N_3158,N_3164);
and U3704 (N_3704,N_3459,N_3496);
nor U3705 (N_3705,N_3328,N_3145);
or U3706 (N_3706,N_3181,N_3485);
nor U3707 (N_3707,N_3455,N_3379);
nor U3708 (N_3708,N_3398,N_3104);
xnor U3709 (N_3709,N_3471,N_3393);
or U3710 (N_3710,N_3384,N_3265);
xnor U3711 (N_3711,N_3377,N_3284);
xor U3712 (N_3712,N_3438,N_3339);
nor U3713 (N_3713,N_3366,N_3034);
nor U3714 (N_3714,N_3347,N_3499);
xnor U3715 (N_3715,N_3317,N_3450);
nor U3716 (N_3716,N_3283,N_3070);
and U3717 (N_3717,N_3016,N_3319);
xor U3718 (N_3718,N_3177,N_3095);
xor U3719 (N_3719,N_3424,N_3280);
nand U3720 (N_3720,N_3153,N_3306);
nor U3721 (N_3721,N_3376,N_3032);
or U3722 (N_3722,N_3014,N_3474);
nand U3723 (N_3723,N_3120,N_3171);
or U3724 (N_3724,N_3160,N_3359);
or U3725 (N_3725,N_3058,N_3367);
xor U3726 (N_3726,N_3415,N_3065);
and U3727 (N_3727,N_3335,N_3208);
nor U3728 (N_3728,N_3375,N_3117);
nor U3729 (N_3729,N_3305,N_3466);
nand U3730 (N_3730,N_3244,N_3055);
or U3731 (N_3731,N_3263,N_3447);
nand U3732 (N_3732,N_3470,N_3182);
nor U3733 (N_3733,N_3225,N_3222);
and U3734 (N_3734,N_3476,N_3172);
nand U3735 (N_3735,N_3400,N_3199);
or U3736 (N_3736,N_3368,N_3155);
or U3737 (N_3737,N_3134,N_3269);
and U3738 (N_3738,N_3066,N_3207);
and U3739 (N_3739,N_3498,N_3291);
xor U3740 (N_3740,N_3399,N_3043);
or U3741 (N_3741,N_3279,N_3201);
or U3742 (N_3742,N_3218,N_3300);
nand U3743 (N_3743,N_3049,N_3054);
and U3744 (N_3744,N_3404,N_3139);
or U3745 (N_3745,N_3075,N_3039);
xnor U3746 (N_3746,N_3082,N_3452);
or U3747 (N_3747,N_3458,N_3073);
or U3748 (N_3748,N_3121,N_3169);
xnor U3749 (N_3749,N_3002,N_3064);
nor U3750 (N_3750,N_3339,N_3490);
xor U3751 (N_3751,N_3372,N_3472);
and U3752 (N_3752,N_3030,N_3049);
xor U3753 (N_3753,N_3194,N_3393);
xnor U3754 (N_3754,N_3339,N_3283);
and U3755 (N_3755,N_3479,N_3451);
nand U3756 (N_3756,N_3114,N_3146);
or U3757 (N_3757,N_3199,N_3034);
xnor U3758 (N_3758,N_3177,N_3232);
or U3759 (N_3759,N_3374,N_3184);
nor U3760 (N_3760,N_3084,N_3135);
nor U3761 (N_3761,N_3064,N_3260);
or U3762 (N_3762,N_3192,N_3287);
xor U3763 (N_3763,N_3219,N_3425);
nand U3764 (N_3764,N_3305,N_3282);
or U3765 (N_3765,N_3001,N_3004);
nand U3766 (N_3766,N_3066,N_3373);
or U3767 (N_3767,N_3180,N_3313);
or U3768 (N_3768,N_3106,N_3002);
xnor U3769 (N_3769,N_3422,N_3294);
nor U3770 (N_3770,N_3392,N_3475);
nand U3771 (N_3771,N_3028,N_3200);
and U3772 (N_3772,N_3234,N_3395);
nor U3773 (N_3773,N_3346,N_3124);
xnor U3774 (N_3774,N_3071,N_3309);
and U3775 (N_3775,N_3126,N_3267);
nand U3776 (N_3776,N_3403,N_3073);
xor U3777 (N_3777,N_3264,N_3251);
xnor U3778 (N_3778,N_3082,N_3026);
or U3779 (N_3779,N_3125,N_3386);
xor U3780 (N_3780,N_3148,N_3388);
or U3781 (N_3781,N_3429,N_3195);
or U3782 (N_3782,N_3114,N_3261);
nor U3783 (N_3783,N_3208,N_3373);
nor U3784 (N_3784,N_3219,N_3090);
and U3785 (N_3785,N_3300,N_3404);
nand U3786 (N_3786,N_3123,N_3409);
nor U3787 (N_3787,N_3477,N_3348);
xor U3788 (N_3788,N_3458,N_3339);
or U3789 (N_3789,N_3385,N_3108);
nand U3790 (N_3790,N_3298,N_3145);
and U3791 (N_3791,N_3389,N_3424);
nor U3792 (N_3792,N_3024,N_3287);
nand U3793 (N_3793,N_3410,N_3100);
and U3794 (N_3794,N_3493,N_3217);
or U3795 (N_3795,N_3321,N_3452);
nor U3796 (N_3796,N_3306,N_3066);
xnor U3797 (N_3797,N_3253,N_3116);
nand U3798 (N_3798,N_3415,N_3443);
xor U3799 (N_3799,N_3092,N_3122);
or U3800 (N_3800,N_3030,N_3435);
nand U3801 (N_3801,N_3113,N_3388);
nor U3802 (N_3802,N_3063,N_3001);
and U3803 (N_3803,N_3412,N_3295);
nor U3804 (N_3804,N_3302,N_3083);
xnor U3805 (N_3805,N_3303,N_3223);
or U3806 (N_3806,N_3065,N_3050);
nand U3807 (N_3807,N_3203,N_3356);
and U3808 (N_3808,N_3185,N_3116);
nand U3809 (N_3809,N_3304,N_3011);
nand U3810 (N_3810,N_3263,N_3432);
nor U3811 (N_3811,N_3246,N_3369);
and U3812 (N_3812,N_3275,N_3077);
and U3813 (N_3813,N_3199,N_3496);
nand U3814 (N_3814,N_3228,N_3023);
and U3815 (N_3815,N_3494,N_3224);
and U3816 (N_3816,N_3192,N_3266);
and U3817 (N_3817,N_3117,N_3351);
xnor U3818 (N_3818,N_3257,N_3111);
nand U3819 (N_3819,N_3180,N_3259);
or U3820 (N_3820,N_3293,N_3484);
nor U3821 (N_3821,N_3122,N_3302);
xnor U3822 (N_3822,N_3203,N_3183);
and U3823 (N_3823,N_3434,N_3333);
nand U3824 (N_3824,N_3192,N_3093);
xor U3825 (N_3825,N_3247,N_3370);
and U3826 (N_3826,N_3224,N_3499);
nor U3827 (N_3827,N_3306,N_3383);
and U3828 (N_3828,N_3330,N_3387);
or U3829 (N_3829,N_3488,N_3439);
and U3830 (N_3830,N_3284,N_3381);
xnor U3831 (N_3831,N_3268,N_3460);
nand U3832 (N_3832,N_3336,N_3148);
xor U3833 (N_3833,N_3366,N_3431);
nor U3834 (N_3834,N_3116,N_3029);
nand U3835 (N_3835,N_3311,N_3464);
or U3836 (N_3836,N_3012,N_3227);
and U3837 (N_3837,N_3496,N_3427);
and U3838 (N_3838,N_3347,N_3307);
xor U3839 (N_3839,N_3073,N_3076);
xnor U3840 (N_3840,N_3362,N_3082);
or U3841 (N_3841,N_3406,N_3015);
nand U3842 (N_3842,N_3304,N_3135);
nand U3843 (N_3843,N_3258,N_3241);
nand U3844 (N_3844,N_3455,N_3000);
xor U3845 (N_3845,N_3483,N_3382);
nor U3846 (N_3846,N_3325,N_3258);
nor U3847 (N_3847,N_3340,N_3079);
nor U3848 (N_3848,N_3127,N_3403);
and U3849 (N_3849,N_3008,N_3461);
xnor U3850 (N_3850,N_3497,N_3110);
or U3851 (N_3851,N_3397,N_3349);
nor U3852 (N_3852,N_3272,N_3397);
or U3853 (N_3853,N_3082,N_3296);
nor U3854 (N_3854,N_3471,N_3400);
or U3855 (N_3855,N_3331,N_3375);
and U3856 (N_3856,N_3190,N_3096);
nand U3857 (N_3857,N_3461,N_3073);
or U3858 (N_3858,N_3321,N_3342);
or U3859 (N_3859,N_3451,N_3307);
nor U3860 (N_3860,N_3437,N_3322);
xor U3861 (N_3861,N_3418,N_3126);
or U3862 (N_3862,N_3139,N_3284);
xnor U3863 (N_3863,N_3366,N_3036);
nor U3864 (N_3864,N_3246,N_3473);
and U3865 (N_3865,N_3472,N_3054);
nand U3866 (N_3866,N_3035,N_3019);
xor U3867 (N_3867,N_3062,N_3073);
or U3868 (N_3868,N_3267,N_3330);
or U3869 (N_3869,N_3052,N_3244);
nand U3870 (N_3870,N_3244,N_3135);
xor U3871 (N_3871,N_3299,N_3261);
or U3872 (N_3872,N_3317,N_3380);
and U3873 (N_3873,N_3442,N_3138);
xnor U3874 (N_3874,N_3419,N_3004);
and U3875 (N_3875,N_3388,N_3217);
or U3876 (N_3876,N_3175,N_3330);
and U3877 (N_3877,N_3008,N_3315);
or U3878 (N_3878,N_3098,N_3066);
xor U3879 (N_3879,N_3021,N_3478);
and U3880 (N_3880,N_3258,N_3176);
nand U3881 (N_3881,N_3095,N_3211);
and U3882 (N_3882,N_3280,N_3420);
xor U3883 (N_3883,N_3039,N_3223);
nand U3884 (N_3884,N_3008,N_3048);
nor U3885 (N_3885,N_3281,N_3352);
xnor U3886 (N_3886,N_3305,N_3081);
nor U3887 (N_3887,N_3296,N_3171);
nand U3888 (N_3888,N_3458,N_3231);
nand U3889 (N_3889,N_3043,N_3006);
nor U3890 (N_3890,N_3106,N_3252);
nand U3891 (N_3891,N_3148,N_3238);
xor U3892 (N_3892,N_3252,N_3138);
or U3893 (N_3893,N_3139,N_3192);
xor U3894 (N_3894,N_3359,N_3103);
and U3895 (N_3895,N_3209,N_3443);
or U3896 (N_3896,N_3220,N_3285);
nand U3897 (N_3897,N_3172,N_3174);
nand U3898 (N_3898,N_3178,N_3326);
xnor U3899 (N_3899,N_3332,N_3217);
nand U3900 (N_3900,N_3397,N_3242);
nor U3901 (N_3901,N_3131,N_3021);
or U3902 (N_3902,N_3363,N_3261);
and U3903 (N_3903,N_3419,N_3247);
xnor U3904 (N_3904,N_3466,N_3221);
and U3905 (N_3905,N_3234,N_3074);
or U3906 (N_3906,N_3342,N_3005);
xnor U3907 (N_3907,N_3295,N_3124);
or U3908 (N_3908,N_3446,N_3018);
and U3909 (N_3909,N_3233,N_3035);
and U3910 (N_3910,N_3272,N_3110);
and U3911 (N_3911,N_3248,N_3363);
nor U3912 (N_3912,N_3385,N_3127);
or U3913 (N_3913,N_3113,N_3056);
and U3914 (N_3914,N_3154,N_3275);
nand U3915 (N_3915,N_3274,N_3080);
or U3916 (N_3916,N_3197,N_3090);
or U3917 (N_3917,N_3493,N_3198);
nor U3918 (N_3918,N_3343,N_3035);
nor U3919 (N_3919,N_3071,N_3493);
xnor U3920 (N_3920,N_3490,N_3472);
nand U3921 (N_3921,N_3373,N_3402);
nor U3922 (N_3922,N_3472,N_3344);
or U3923 (N_3923,N_3235,N_3349);
and U3924 (N_3924,N_3335,N_3402);
nand U3925 (N_3925,N_3086,N_3030);
nor U3926 (N_3926,N_3293,N_3183);
or U3927 (N_3927,N_3443,N_3004);
xnor U3928 (N_3928,N_3283,N_3394);
nor U3929 (N_3929,N_3124,N_3038);
xor U3930 (N_3930,N_3493,N_3458);
nand U3931 (N_3931,N_3288,N_3309);
and U3932 (N_3932,N_3368,N_3191);
xor U3933 (N_3933,N_3304,N_3125);
nand U3934 (N_3934,N_3009,N_3019);
nand U3935 (N_3935,N_3452,N_3425);
or U3936 (N_3936,N_3435,N_3010);
nand U3937 (N_3937,N_3037,N_3464);
and U3938 (N_3938,N_3294,N_3190);
xnor U3939 (N_3939,N_3181,N_3319);
nor U3940 (N_3940,N_3429,N_3357);
xnor U3941 (N_3941,N_3497,N_3492);
nand U3942 (N_3942,N_3356,N_3057);
xnor U3943 (N_3943,N_3368,N_3355);
xnor U3944 (N_3944,N_3279,N_3455);
xor U3945 (N_3945,N_3111,N_3218);
xor U3946 (N_3946,N_3099,N_3078);
xor U3947 (N_3947,N_3366,N_3226);
nand U3948 (N_3948,N_3051,N_3232);
nand U3949 (N_3949,N_3039,N_3470);
nor U3950 (N_3950,N_3022,N_3481);
and U3951 (N_3951,N_3152,N_3418);
nor U3952 (N_3952,N_3484,N_3065);
xor U3953 (N_3953,N_3057,N_3450);
nand U3954 (N_3954,N_3189,N_3492);
and U3955 (N_3955,N_3468,N_3289);
nand U3956 (N_3956,N_3090,N_3439);
or U3957 (N_3957,N_3146,N_3176);
xor U3958 (N_3958,N_3024,N_3328);
and U3959 (N_3959,N_3418,N_3057);
and U3960 (N_3960,N_3219,N_3315);
nor U3961 (N_3961,N_3074,N_3277);
nand U3962 (N_3962,N_3101,N_3042);
and U3963 (N_3963,N_3225,N_3230);
nor U3964 (N_3964,N_3414,N_3300);
nor U3965 (N_3965,N_3373,N_3067);
and U3966 (N_3966,N_3421,N_3454);
xor U3967 (N_3967,N_3217,N_3394);
or U3968 (N_3968,N_3372,N_3041);
nor U3969 (N_3969,N_3499,N_3303);
xor U3970 (N_3970,N_3391,N_3150);
xnor U3971 (N_3971,N_3063,N_3020);
or U3972 (N_3972,N_3410,N_3132);
nand U3973 (N_3973,N_3351,N_3456);
and U3974 (N_3974,N_3061,N_3314);
xor U3975 (N_3975,N_3097,N_3240);
xnor U3976 (N_3976,N_3138,N_3062);
and U3977 (N_3977,N_3074,N_3219);
or U3978 (N_3978,N_3253,N_3192);
xnor U3979 (N_3979,N_3111,N_3245);
nand U3980 (N_3980,N_3196,N_3190);
nor U3981 (N_3981,N_3153,N_3122);
nand U3982 (N_3982,N_3480,N_3332);
nor U3983 (N_3983,N_3302,N_3033);
or U3984 (N_3984,N_3131,N_3461);
or U3985 (N_3985,N_3496,N_3006);
and U3986 (N_3986,N_3300,N_3068);
nor U3987 (N_3987,N_3115,N_3060);
or U3988 (N_3988,N_3045,N_3499);
xnor U3989 (N_3989,N_3401,N_3405);
or U3990 (N_3990,N_3206,N_3074);
nor U3991 (N_3991,N_3013,N_3433);
nand U3992 (N_3992,N_3011,N_3195);
or U3993 (N_3993,N_3027,N_3007);
nand U3994 (N_3994,N_3026,N_3299);
and U3995 (N_3995,N_3093,N_3349);
and U3996 (N_3996,N_3087,N_3332);
nor U3997 (N_3997,N_3378,N_3321);
and U3998 (N_3998,N_3189,N_3388);
nand U3999 (N_3999,N_3341,N_3137);
nand U4000 (N_4000,N_3875,N_3998);
nor U4001 (N_4001,N_3984,N_3709);
or U4002 (N_4002,N_3932,N_3661);
xnor U4003 (N_4003,N_3884,N_3793);
or U4004 (N_4004,N_3936,N_3975);
nand U4005 (N_4005,N_3664,N_3929);
nor U4006 (N_4006,N_3608,N_3504);
nor U4007 (N_4007,N_3509,N_3843);
nand U4008 (N_4008,N_3510,N_3912);
nand U4009 (N_4009,N_3727,N_3581);
nand U4010 (N_4010,N_3853,N_3803);
nor U4011 (N_4011,N_3535,N_3553);
nor U4012 (N_4012,N_3758,N_3696);
or U4013 (N_4013,N_3873,N_3606);
nor U4014 (N_4014,N_3710,N_3980);
or U4015 (N_4015,N_3792,N_3940);
nor U4016 (N_4016,N_3882,N_3533);
or U4017 (N_4017,N_3768,N_3741);
xnor U4018 (N_4018,N_3848,N_3635);
and U4019 (N_4019,N_3777,N_3693);
nand U4020 (N_4020,N_3852,N_3740);
nand U4021 (N_4021,N_3555,N_3755);
nand U4022 (N_4022,N_3500,N_3885);
nor U4023 (N_4023,N_3829,N_3986);
nand U4024 (N_4024,N_3665,N_3917);
xnor U4025 (N_4025,N_3678,N_3840);
nand U4026 (N_4026,N_3810,N_3604);
and U4027 (N_4027,N_3780,N_3673);
or U4028 (N_4028,N_3860,N_3800);
nor U4029 (N_4029,N_3874,N_3839);
xnor U4030 (N_4030,N_3551,N_3545);
or U4031 (N_4031,N_3869,N_3788);
nor U4032 (N_4032,N_3914,N_3719);
or U4033 (N_4033,N_3713,N_3631);
or U4034 (N_4034,N_3592,N_3683);
and U4035 (N_4035,N_3992,N_3970);
or U4036 (N_4036,N_3981,N_3762);
and U4037 (N_4037,N_3522,N_3933);
xor U4038 (N_4038,N_3680,N_3973);
and U4039 (N_4039,N_3819,N_3603);
and U4040 (N_4040,N_3775,N_3989);
and U4041 (N_4041,N_3627,N_3797);
nor U4042 (N_4042,N_3733,N_3677);
or U4043 (N_4043,N_3920,N_3619);
xor U4044 (N_4044,N_3865,N_3764);
and U4045 (N_4045,N_3638,N_3574);
nand U4046 (N_4046,N_3773,N_3960);
nor U4047 (N_4047,N_3612,N_3751);
and U4048 (N_4048,N_3567,N_3763);
or U4049 (N_4049,N_3903,N_3889);
nand U4050 (N_4050,N_3597,N_3937);
or U4051 (N_4051,N_3537,N_3676);
nand U4052 (N_4052,N_3689,N_3939);
nand U4053 (N_4053,N_3894,N_3947);
nor U4054 (N_4054,N_3717,N_3536);
nor U4055 (N_4055,N_3613,N_3811);
and U4056 (N_4056,N_3972,N_3790);
or U4057 (N_4057,N_3923,N_3895);
xor U4058 (N_4058,N_3618,N_3626);
nand U4059 (N_4059,N_3785,N_3691);
or U4060 (N_4060,N_3759,N_3589);
or U4061 (N_4061,N_3783,N_3672);
and U4062 (N_4062,N_3658,N_3890);
nor U4063 (N_4063,N_3897,N_3963);
or U4064 (N_4064,N_3871,N_3556);
nand U4065 (N_4065,N_3909,N_3988);
xnor U4066 (N_4066,N_3594,N_3571);
nand U4067 (N_4067,N_3948,N_3506);
nor U4068 (N_4068,N_3669,N_3760);
xnor U4069 (N_4069,N_3952,N_3904);
or U4070 (N_4070,N_3805,N_3979);
xnor U4071 (N_4071,N_3649,N_3739);
xor U4072 (N_4072,N_3982,N_3667);
xor U4073 (N_4073,N_3930,N_3996);
nor U4074 (N_4074,N_3786,N_3718);
xor U4075 (N_4075,N_3699,N_3644);
or U4076 (N_4076,N_3528,N_3985);
and U4077 (N_4077,N_3624,N_3579);
and U4078 (N_4078,N_3799,N_3549);
nand U4079 (N_4079,N_3744,N_3828);
and U4080 (N_4080,N_3888,N_3637);
and U4081 (N_4081,N_3902,N_3527);
and U4082 (N_4082,N_3891,N_3663);
xor U4083 (N_4083,N_3690,N_3515);
nand U4084 (N_4084,N_3514,N_3507);
or U4085 (N_4085,N_3511,N_3955);
nor U4086 (N_4086,N_3942,N_3765);
xnor U4087 (N_4087,N_3832,N_3841);
xnor U4088 (N_4088,N_3971,N_3812);
or U4089 (N_4089,N_3781,N_3993);
and U4090 (N_4090,N_3610,N_3931);
nand U4091 (N_4091,N_3750,N_3732);
xor U4092 (N_4092,N_3961,N_3916);
nand U4093 (N_4093,N_3628,N_3830);
nor U4094 (N_4094,N_3737,N_3659);
nor U4095 (N_4095,N_3561,N_3962);
nor U4096 (N_4096,N_3681,N_3726);
xor U4097 (N_4097,N_3542,N_3856);
nor U4098 (N_4098,N_3827,N_3734);
xor U4099 (N_4099,N_3602,N_3804);
nor U4100 (N_4100,N_3876,N_3731);
nor U4101 (N_4101,N_3591,N_3629);
or U4102 (N_4102,N_3974,N_3958);
nand U4103 (N_4103,N_3558,N_3508);
nand U4104 (N_4104,N_3587,N_3872);
nor U4105 (N_4105,N_3572,N_3703);
and U4106 (N_4106,N_3994,N_3593);
nand U4107 (N_4107,N_3941,N_3815);
or U4108 (N_4108,N_3531,N_3700);
nand U4109 (N_4109,N_3938,N_3774);
nand U4110 (N_4110,N_3600,N_3798);
or U4111 (N_4111,N_3776,N_3825);
and U4112 (N_4112,N_3576,N_3953);
and U4113 (N_4113,N_3769,N_3701);
or U4114 (N_4114,N_3564,N_3670);
and U4115 (N_4115,N_3950,N_3565);
xnor U4116 (N_4116,N_3820,N_3653);
nand U4117 (N_4117,N_3578,N_3794);
xor U4118 (N_4118,N_3622,N_3879);
nand U4119 (N_4119,N_3711,N_3826);
nand U4120 (N_4120,N_3534,N_3523);
nor U4121 (N_4121,N_3999,N_3599);
nor U4122 (N_4122,N_3706,N_3857);
nand U4123 (N_4123,N_3708,N_3625);
and U4124 (N_4124,N_3684,N_3870);
and U4125 (N_4125,N_3590,N_3822);
nand U4126 (N_4126,N_3559,N_3557);
or U4127 (N_4127,N_3566,N_3813);
or U4128 (N_4128,N_3715,N_3656);
xor U4129 (N_4129,N_3756,N_3648);
nand U4130 (N_4130,N_3789,N_3862);
xor U4131 (N_4131,N_3854,N_3520);
and U4132 (N_4132,N_3687,N_3541);
nor U4133 (N_4133,N_3598,N_3607);
or U4134 (N_4134,N_3913,N_3723);
nand U4135 (N_4135,N_3978,N_3688);
nand U4136 (N_4136,N_3584,N_3666);
or U4137 (N_4137,N_3925,N_3752);
nand U4138 (N_4138,N_3809,N_3521);
xnor U4139 (N_4139,N_3643,N_3646);
and U4140 (N_4140,N_3944,N_3532);
and U4141 (N_4141,N_3632,N_3833);
or U4142 (N_4142,N_3836,N_3802);
nand U4143 (N_4143,N_3991,N_3596);
nand U4144 (N_4144,N_3867,N_3630);
and U4145 (N_4145,N_3801,N_3570);
or U4146 (N_4146,N_3831,N_3838);
and U4147 (N_4147,N_3761,N_3943);
xnor U4148 (N_4148,N_3851,N_3868);
and U4149 (N_4149,N_3617,N_3580);
nand U4150 (N_4150,N_3907,N_3966);
or U4151 (N_4151,N_3512,N_3660);
and U4152 (N_4152,N_3995,N_3787);
nand U4153 (N_4153,N_3766,N_3880);
and U4154 (N_4154,N_3641,N_3883);
and U4155 (N_4155,N_3864,N_3905);
nand U4156 (N_4156,N_3503,N_3725);
or U4157 (N_4157,N_3562,N_3807);
xnor U4158 (N_4158,N_3662,N_3530);
and U4159 (N_4159,N_3910,N_3538);
and U4160 (N_4160,N_3892,N_3863);
or U4161 (N_4161,N_3736,N_3563);
or U4162 (N_4162,N_3539,N_3846);
nand U4163 (N_4163,N_3650,N_3735);
nor U4164 (N_4164,N_3573,N_3749);
xnor U4165 (N_4165,N_3816,N_3771);
xnor U4166 (N_4166,N_3569,N_3784);
nand U4167 (N_4167,N_3518,N_3657);
nand U4168 (N_4168,N_3900,N_3652);
nor U4169 (N_4169,N_3823,N_3834);
and U4170 (N_4170,N_3611,N_3645);
nor U4171 (N_4171,N_3983,N_3621);
and U4172 (N_4172,N_3821,N_3745);
and U4173 (N_4173,N_3906,N_3908);
xnor U4174 (N_4174,N_3837,N_3866);
nand U4175 (N_4175,N_3547,N_3616);
nand U4176 (N_4176,N_3817,N_3921);
nand U4177 (N_4177,N_3550,N_3695);
or U4178 (N_4178,N_3588,N_3540);
and U4179 (N_4179,N_3716,N_3704);
or U4180 (N_4180,N_3634,N_3772);
xor U4181 (N_4181,N_3746,N_3525);
xnor U4182 (N_4182,N_3582,N_3742);
and U4183 (N_4183,N_3965,N_3642);
or U4184 (N_4184,N_3605,N_3881);
and U4185 (N_4185,N_3779,N_3835);
nor U4186 (N_4186,N_3585,N_3791);
xnor U4187 (N_4187,N_3844,N_3918);
or U4188 (N_4188,N_3712,N_3956);
xnor U4189 (N_4189,N_3969,N_3502);
and U4190 (N_4190,N_3639,N_3620);
xnor U4191 (N_4191,N_3721,N_3546);
or U4192 (N_4192,N_3577,N_3796);
or U4193 (N_4193,N_3778,N_3682);
nand U4194 (N_4194,N_3977,N_3850);
nand U4195 (N_4195,N_3782,N_3517);
nor U4196 (N_4196,N_3901,N_3886);
or U4197 (N_4197,N_3859,N_3685);
nor U4198 (N_4198,N_3560,N_3928);
or U4199 (N_4199,N_3738,N_3767);
xnor U4200 (N_4200,N_3548,N_3694);
nand U4201 (N_4201,N_3806,N_3946);
xnor U4202 (N_4202,N_3899,N_3697);
nor U4203 (N_4203,N_3702,N_3858);
or U4204 (N_4204,N_3568,N_3651);
nand U4205 (N_4205,N_3967,N_3516);
nor U4206 (N_4206,N_3926,N_3714);
nor U4207 (N_4207,N_3674,N_3849);
nand U4208 (N_4208,N_3722,N_3935);
nor U4209 (N_4209,N_3698,N_3959);
xor U4210 (N_4210,N_3524,N_3855);
and U4211 (N_4211,N_3583,N_3997);
or U4212 (N_4212,N_3505,N_3519);
nand U4213 (N_4213,N_3949,N_3818);
nor U4214 (N_4214,N_3575,N_3987);
xnor U4215 (N_4215,N_3898,N_3896);
and U4216 (N_4216,N_3808,N_3730);
or U4217 (N_4217,N_3640,N_3877);
or U4218 (N_4218,N_3990,N_3842);
xnor U4219 (N_4219,N_3526,N_3623);
xor U4220 (N_4220,N_3922,N_3747);
or U4221 (N_4221,N_3501,N_3692);
and U4222 (N_4222,N_3945,N_3615);
xnor U4223 (N_4223,N_3911,N_3887);
nand U4224 (N_4224,N_3795,N_3878);
xnor U4225 (N_4225,N_3586,N_3595);
nand U4226 (N_4226,N_3743,N_3705);
and U4227 (N_4227,N_3513,N_3847);
xor U4228 (N_4228,N_3543,N_3636);
and U4229 (N_4229,N_3919,N_3601);
nand U4230 (N_4230,N_3968,N_3927);
nor U4231 (N_4231,N_3893,N_3729);
nand U4232 (N_4232,N_3675,N_3954);
xnor U4233 (N_4233,N_3861,N_3976);
nor U4234 (N_4234,N_3924,N_3679);
or U4235 (N_4235,N_3824,N_3686);
and U4236 (N_4236,N_3770,N_3957);
and U4237 (N_4237,N_3554,N_3934);
nor U4238 (N_4238,N_3647,N_3951);
nor U4239 (N_4239,N_3720,N_3614);
or U4240 (N_4240,N_3814,N_3609);
xnor U4241 (N_4241,N_3728,N_3964);
or U4242 (N_4242,N_3724,N_3754);
nor U4243 (N_4243,N_3671,N_3845);
xnor U4244 (N_4244,N_3668,N_3757);
or U4245 (N_4245,N_3552,N_3655);
nand U4246 (N_4246,N_3529,N_3633);
or U4247 (N_4247,N_3654,N_3544);
or U4248 (N_4248,N_3753,N_3915);
nor U4249 (N_4249,N_3707,N_3748);
and U4250 (N_4250,N_3764,N_3805);
nor U4251 (N_4251,N_3692,N_3666);
nand U4252 (N_4252,N_3976,N_3616);
nand U4253 (N_4253,N_3814,N_3951);
and U4254 (N_4254,N_3933,N_3851);
nor U4255 (N_4255,N_3661,N_3615);
nand U4256 (N_4256,N_3573,N_3798);
xnor U4257 (N_4257,N_3949,N_3564);
xnor U4258 (N_4258,N_3688,N_3804);
and U4259 (N_4259,N_3749,N_3654);
and U4260 (N_4260,N_3624,N_3777);
nor U4261 (N_4261,N_3607,N_3809);
nand U4262 (N_4262,N_3664,N_3883);
nand U4263 (N_4263,N_3848,N_3659);
or U4264 (N_4264,N_3530,N_3567);
nand U4265 (N_4265,N_3773,N_3597);
or U4266 (N_4266,N_3961,N_3871);
or U4267 (N_4267,N_3583,N_3977);
xnor U4268 (N_4268,N_3533,N_3867);
xnor U4269 (N_4269,N_3944,N_3560);
or U4270 (N_4270,N_3649,N_3772);
xor U4271 (N_4271,N_3966,N_3909);
nor U4272 (N_4272,N_3943,N_3795);
nand U4273 (N_4273,N_3705,N_3786);
and U4274 (N_4274,N_3614,N_3812);
xnor U4275 (N_4275,N_3803,N_3552);
nand U4276 (N_4276,N_3967,N_3931);
and U4277 (N_4277,N_3913,N_3676);
nand U4278 (N_4278,N_3588,N_3574);
nor U4279 (N_4279,N_3956,N_3867);
nor U4280 (N_4280,N_3523,N_3980);
nor U4281 (N_4281,N_3522,N_3595);
nand U4282 (N_4282,N_3640,N_3883);
xor U4283 (N_4283,N_3790,N_3524);
nor U4284 (N_4284,N_3804,N_3983);
nor U4285 (N_4285,N_3671,N_3874);
xor U4286 (N_4286,N_3535,N_3893);
xnor U4287 (N_4287,N_3759,N_3649);
or U4288 (N_4288,N_3878,N_3660);
or U4289 (N_4289,N_3616,N_3869);
nor U4290 (N_4290,N_3616,N_3702);
nor U4291 (N_4291,N_3621,N_3562);
nand U4292 (N_4292,N_3689,N_3619);
xor U4293 (N_4293,N_3997,N_3747);
and U4294 (N_4294,N_3650,N_3736);
and U4295 (N_4295,N_3716,N_3889);
nor U4296 (N_4296,N_3675,N_3794);
nor U4297 (N_4297,N_3947,N_3849);
nor U4298 (N_4298,N_3827,N_3861);
or U4299 (N_4299,N_3868,N_3842);
or U4300 (N_4300,N_3702,N_3921);
or U4301 (N_4301,N_3658,N_3528);
or U4302 (N_4302,N_3689,N_3534);
nand U4303 (N_4303,N_3834,N_3901);
and U4304 (N_4304,N_3738,N_3680);
or U4305 (N_4305,N_3923,N_3809);
nand U4306 (N_4306,N_3576,N_3758);
xor U4307 (N_4307,N_3638,N_3868);
nor U4308 (N_4308,N_3959,N_3774);
or U4309 (N_4309,N_3812,N_3532);
nor U4310 (N_4310,N_3521,N_3691);
xnor U4311 (N_4311,N_3527,N_3733);
or U4312 (N_4312,N_3839,N_3746);
and U4313 (N_4313,N_3859,N_3749);
nand U4314 (N_4314,N_3806,N_3859);
nand U4315 (N_4315,N_3866,N_3619);
xor U4316 (N_4316,N_3614,N_3736);
and U4317 (N_4317,N_3509,N_3500);
and U4318 (N_4318,N_3964,N_3610);
nand U4319 (N_4319,N_3846,N_3763);
nand U4320 (N_4320,N_3886,N_3733);
or U4321 (N_4321,N_3730,N_3961);
or U4322 (N_4322,N_3914,N_3648);
nand U4323 (N_4323,N_3525,N_3766);
and U4324 (N_4324,N_3634,N_3974);
and U4325 (N_4325,N_3896,N_3626);
nand U4326 (N_4326,N_3619,N_3950);
or U4327 (N_4327,N_3936,N_3920);
or U4328 (N_4328,N_3788,N_3639);
and U4329 (N_4329,N_3879,N_3760);
nand U4330 (N_4330,N_3511,N_3891);
and U4331 (N_4331,N_3645,N_3845);
or U4332 (N_4332,N_3566,N_3968);
nand U4333 (N_4333,N_3647,N_3953);
nand U4334 (N_4334,N_3622,N_3928);
xnor U4335 (N_4335,N_3976,N_3692);
and U4336 (N_4336,N_3537,N_3953);
and U4337 (N_4337,N_3895,N_3767);
nor U4338 (N_4338,N_3674,N_3517);
nand U4339 (N_4339,N_3953,N_3731);
and U4340 (N_4340,N_3549,N_3701);
nand U4341 (N_4341,N_3770,N_3931);
nand U4342 (N_4342,N_3909,N_3828);
nand U4343 (N_4343,N_3629,N_3867);
and U4344 (N_4344,N_3542,N_3609);
or U4345 (N_4345,N_3672,N_3503);
xnor U4346 (N_4346,N_3544,N_3561);
xor U4347 (N_4347,N_3531,N_3722);
xnor U4348 (N_4348,N_3928,N_3638);
xnor U4349 (N_4349,N_3656,N_3558);
xor U4350 (N_4350,N_3531,N_3872);
xnor U4351 (N_4351,N_3502,N_3966);
xor U4352 (N_4352,N_3526,N_3667);
nor U4353 (N_4353,N_3525,N_3951);
and U4354 (N_4354,N_3784,N_3539);
xnor U4355 (N_4355,N_3810,N_3612);
nand U4356 (N_4356,N_3937,N_3674);
nand U4357 (N_4357,N_3858,N_3608);
and U4358 (N_4358,N_3708,N_3569);
or U4359 (N_4359,N_3698,N_3684);
or U4360 (N_4360,N_3502,N_3791);
nand U4361 (N_4361,N_3657,N_3963);
or U4362 (N_4362,N_3971,N_3924);
nand U4363 (N_4363,N_3850,N_3772);
and U4364 (N_4364,N_3967,N_3789);
and U4365 (N_4365,N_3684,N_3637);
nor U4366 (N_4366,N_3750,N_3528);
xnor U4367 (N_4367,N_3934,N_3942);
or U4368 (N_4368,N_3921,N_3762);
or U4369 (N_4369,N_3999,N_3543);
xor U4370 (N_4370,N_3552,N_3767);
or U4371 (N_4371,N_3659,N_3962);
xnor U4372 (N_4372,N_3826,N_3765);
or U4373 (N_4373,N_3971,N_3846);
or U4374 (N_4374,N_3733,N_3811);
or U4375 (N_4375,N_3550,N_3995);
or U4376 (N_4376,N_3948,N_3808);
xnor U4377 (N_4377,N_3698,N_3739);
or U4378 (N_4378,N_3875,N_3979);
xor U4379 (N_4379,N_3944,N_3522);
nor U4380 (N_4380,N_3956,N_3847);
or U4381 (N_4381,N_3952,N_3702);
or U4382 (N_4382,N_3570,N_3756);
xor U4383 (N_4383,N_3668,N_3533);
nor U4384 (N_4384,N_3540,N_3961);
nand U4385 (N_4385,N_3647,N_3973);
and U4386 (N_4386,N_3594,N_3643);
nor U4387 (N_4387,N_3823,N_3814);
nand U4388 (N_4388,N_3673,N_3769);
and U4389 (N_4389,N_3973,N_3779);
xor U4390 (N_4390,N_3749,N_3780);
and U4391 (N_4391,N_3544,N_3939);
nand U4392 (N_4392,N_3518,N_3750);
nand U4393 (N_4393,N_3500,N_3946);
or U4394 (N_4394,N_3666,N_3703);
xor U4395 (N_4395,N_3594,N_3769);
nor U4396 (N_4396,N_3919,N_3812);
nor U4397 (N_4397,N_3768,N_3690);
xor U4398 (N_4398,N_3960,N_3586);
xnor U4399 (N_4399,N_3934,N_3507);
and U4400 (N_4400,N_3994,N_3854);
nor U4401 (N_4401,N_3906,N_3629);
xor U4402 (N_4402,N_3915,N_3869);
nand U4403 (N_4403,N_3560,N_3852);
xor U4404 (N_4404,N_3747,N_3889);
nand U4405 (N_4405,N_3620,N_3584);
nor U4406 (N_4406,N_3857,N_3932);
nor U4407 (N_4407,N_3908,N_3997);
or U4408 (N_4408,N_3713,N_3892);
nand U4409 (N_4409,N_3837,N_3755);
nand U4410 (N_4410,N_3560,N_3541);
and U4411 (N_4411,N_3513,N_3555);
and U4412 (N_4412,N_3882,N_3696);
xor U4413 (N_4413,N_3902,N_3840);
or U4414 (N_4414,N_3839,N_3767);
nor U4415 (N_4415,N_3606,N_3706);
nand U4416 (N_4416,N_3937,N_3571);
or U4417 (N_4417,N_3696,N_3569);
or U4418 (N_4418,N_3744,N_3949);
or U4419 (N_4419,N_3888,N_3642);
or U4420 (N_4420,N_3833,N_3722);
or U4421 (N_4421,N_3874,N_3709);
nor U4422 (N_4422,N_3788,N_3594);
nand U4423 (N_4423,N_3740,N_3922);
and U4424 (N_4424,N_3925,N_3964);
nor U4425 (N_4425,N_3957,N_3986);
nor U4426 (N_4426,N_3523,N_3872);
nand U4427 (N_4427,N_3504,N_3799);
nor U4428 (N_4428,N_3940,N_3745);
nand U4429 (N_4429,N_3971,N_3519);
nand U4430 (N_4430,N_3730,N_3553);
or U4431 (N_4431,N_3778,N_3541);
nand U4432 (N_4432,N_3773,N_3816);
nor U4433 (N_4433,N_3982,N_3634);
nor U4434 (N_4434,N_3755,N_3686);
nand U4435 (N_4435,N_3951,N_3978);
and U4436 (N_4436,N_3681,N_3831);
nand U4437 (N_4437,N_3809,N_3976);
nand U4438 (N_4438,N_3534,N_3536);
and U4439 (N_4439,N_3702,N_3672);
xor U4440 (N_4440,N_3957,N_3634);
or U4441 (N_4441,N_3984,N_3650);
or U4442 (N_4442,N_3962,N_3750);
nor U4443 (N_4443,N_3751,N_3880);
nand U4444 (N_4444,N_3852,N_3831);
xor U4445 (N_4445,N_3899,N_3889);
nand U4446 (N_4446,N_3507,N_3979);
or U4447 (N_4447,N_3558,N_3511);
xor U4448 (N_4448,N_3614,N_3668);
xnor U4449 (N_4449,N_3969,N_3550);
nand U4450 (N_4450,N_3731,N_3682);
nor U4451 (N_4451,N_3889,N_3524);
or U4452 (N_4452,N_3626,N_3690);
and U4453 (N_4453,N_3894,N_3744);
nor U4454 (N_4454,N_3588,N_3900);
nor U4455 (N_4455,N_3950,N_3926);
nor U4456 (N_4456,N_3814,N_3767);
nor U4457 (N_4457,N_3852,N_3621);
or U4458 (N_4458,N_3593,N_3882);
or U4459 (N_4459,N_3593,N_3744);
and U4460 (N_4460,N_3631,N_3633);
or U4461 (N_4461,N_3539,N_3618);
xnor U4462 (N_4462,N_3556,N_3798);
nand U4463 (N_4463,N_3578,N_3954);
and U4464 (N_4464,N_3840,N_3922);
xor U4465 (N_4465,N_3750,N_3568);
or U4466 (N_4466,N_3708,N_3943);
or U4467 (N_4467,N_3763,N_3808);
xnor U4468 (N_4468,N_3785,N_3960);
or U4469 (N_4469,N_3788,N_3728);
or U4470 (N_4470,N_3782,N_3927);
and U4471 (N_4471,N_3812,N_3945);
nor U4472 (N_4472,N_3907,N_3880);
nor U4473 (N_4473,N_3807,N_3773);
and U4474 (N_4474,N_3688,N_3692);
xor U4475 (N_4475,N_3867,N_3662);
nor U4476 (N_4476,N_3837,N_3706);
and U4477 (N_4477,N_3939,N_3563);
or U4478 (N_4478,N_3522,N_3816);
nand U4479 (N_4479,N_3595,N_3726);
and U4480 (N_4480,N_3893,N_3609);
nand U4481 (N_4481,N_3896,N_3831);
xnor U4482 (N_4482,N_3701,N_3552);
and U4483 (N_4483,N_3833,N_3565);
or U4484 (N_4484,N_3551,N_3691);
nand U4485 (N_4485,N_3992,N_3601);
or U4486 (N_4486,N_3868,N_3527);
and U4487 (N_4487,N_3502,N_3665);
nor U4488 (N_4488,N_3808,N_3503);
xnor U4489 (N_4489,N_3534,N_3854);
and U4490 (N_4490,N_3665,N_3609);
xnor U4491 (N_4491,N_3727,N_3968);
or U4492 (N_4492,N_3578,N_3943);
nor U4493 (N_4493,N_3642,N_3658);
nand U4494 (N_4494,N_3599,N_3786);
xnor U4495 (N_4495,N_3695,N_3902);
nor U4496 (N_4496,N_3695,N_3734);
xor U4497 (N_4497,N_3884,N_3626);
nor U4498 (N_4498,N_3585,N_3763);
nor U4499 (N_4499,N_3807,N_3654);
xor U4500 (N_4500,N_4223,N_4144);
nand U4501 (N_4501,N_4299,N_4078);
nor U4502 (N_4502,N_4374,N_4030);
nor U4503 (N_4503,N_4140,N_4232);
xnor U4504 (N_4504,N_4335,N_4365);
and U4505 (N_4505,N_4449,N_4239);
xnor U4506 (N_4506,N_4105,N_4379);
xor U4507 (N_4507,N_4020,N_4316);
nor U4508 (N_4508,N_4035,N_4005);
xnor U4509 (N_4509,N_4475,N_4034);
nand U4510 (N_4510,N_4019,N_4385);
or U4511 (N_4511,N_4430,N_4151);
nand U4512 (N_4512,N_4132,N_4157);
nand U4513 (N_4513,N_4314,N_4348);
xor U4514 (N_4514,N_4127,N_4126);
and U4515 (N_4515,N_4227,N_4333);
and U4516 (N_4516,N_4468,N_4286);
and U4517 (N_4517,N_4162,N_4395);
or U4518 (N_4518,N_4474,N_4330);
nor U4519 (N_4519,N_4349,N_4000);
xor U4520 (N_4520,N_4325,N_4014);
or U4521 (N_4521,N_4300,N_4022);
nand U4522 (N_4522,N_4161,N_4398);
nand U4523 (N_4523,N_4143,N_4359);
and U4524 (N_4524,N_4495,N_4066);
and U4525 (N_4525,N_4113,N_4252);
nor U4526 (N_4526,N_4195,N_4188);
xor U4527 (N_4527,N_4179,N_4202);
or U4528 (N_4528,N_4448,N_4049);
and U4529 (N_4529,N_4294,N_4094);
nand U4530 (N_4530,N_4269,N_4487);
and U4531 (N_4531,N_4375,N_4290);
nand U4532 (N_4532,N_4399,N_4275);
nor U4533 (N_4533,N_4317,N_4198);
xor U4534 (N_4534,N_4362,N_4021);
and U4535 (N_4535,N_4410,N_4027);
and U4536 (N_4536,N_4381,N_4055);
or U4537 (N_4537,N_4110,N_4007);
and U4538 (N_4538,N_4420,N_4422);
or U4539 (N_4539,N_4102,N_4283);
and U4540 (N_4540,N_4263,N_4409);
xnor U4541 (N_4541,N_4204,N_4150);
nand U4542 (N_4542,N_4208,N_4077);
nand U4543 (N_4543,N_4130,N_4396);
nor U4544 (N_4544,N_4192,N_4224);
and U4545 (N_4545,N_4011,N_4322);
or U4546 (N_4546,N_4218,N_4042);
xnor U4547 (N_4547,N_4366,N_4236);
nor U4548 (N_4548,N_4436,N_4407);
nand U4549 (N_4549,N_4009,N_4016);
or U4550 (N_4550,N_4393,N_4051);
nor U4551 (N_4551,N_4104,N_4092);
xor U4552 (N_4552,N_4197,N_4103);
and U4553 (N_4553,N_4115,N_4018);
or U4554 (N_4554,N_4040,N_4251);
xor U4555 (N_4555,N_4419,N_4068);
and U4556 (N_4556,N_4072,N_4471);
nor U4557 (N_4557,N_4321,N_4203);
and U4558 (N_4558,N_4212,N_4340);
xnor U4559 (N_4559,N_4411,N_4106);
xor U4560 (N_4560,N_4026,N_4033);
xnor U4561 (N_4561,N_4098,N_4280);
xor U4562 (N_4562,N_4477,N_4047);
nand U4563 (N_4563,N_4341,N_4155);
nor U4564 (N_4564,N_4220,N_4160);
and U4565 (N_4565,N_4295,N_4453);
nor U4566 (N_4566,N_4045,N_4258);
xnor U4567 (N_4567,N_4056,N_4063);
and U4568 (N_4568,N_4472,N_4390);
xnor U4569 (N_4569,N_4059,N_4061);
and U4570 (N_4570,N_4323,N_4108);
or U4571 (N_4571,N_4185,N_4264);
nor U4572 (N_4572,N_4326,N_4320);
nor U4573 (N_4573,N_4125,N_4433);
xor U4574 (N_4574,N_4303,N_4214);
nor U4575 (N_4575,N_4431,N_4121);
nor U4576 (N_4576,N_4384,N_4173);
and U4577 (N_4577,N_4165,N_4193);
or U4578 (N_4578,N_4073,N_4378);
and U4579 (N_4579,N_4265,N_4046);
nor U4580 (N_4580,N_4194,N_4332);
nand U4581 (N_4581,N_4081,N_4201);
and U4582 (N_4582,N_4350,N_4071);
and U4583 (N_4583,N_4497,N_4248);
and U4584 (N_4584,N_4039,N_4416);
or U4585 (N_4585,N_4304,N_4250);
nand U4586 (N_4586,N_4156,N_4397);
nand U4587 (N_4587,N_4454,N_4158);
or U4588 (N_4588,N_4228,N_4461);
xor U4589 (N_4589,N_4480,N_4235);
or U4590 (N_4590,N_4344,N_4358);
xor U4591 (N_4591,N_4360,N_4288);
nand U4592 (N_4592,N_4423,N_4270);
and U4593 (N_4593,N_4371,N_4446);
and U4594 (N_4594,N_4476,N_4057);
nand U4595 (N_4595,N_4222,N_4012);
or U4596 (N_4596,N_4498,N_4364);
or U4597 (N_4597,N_4154,N_4319);
xnor U4598 (N_4598,N_4484,N_4262);
nor U4599 (N_4599,N_4435,N_4301);
and U4600 (N_4600,N_4413,N_4470);
nand U4601 (N_4601,N_4003,N_4240);
nor U4602 (N_4602,N_4405,N_4302);
nand U4603 (N_4603,N_4266,N_4353);
nor U4604 (N_4604,N_4052,N_4309);
nor U4605 (N_4605,N_4412,N_4230);
and U4606 (N_4606,N_4207,N_4216);
nor U4607 (N_4607,N_4123,N_4277);
or U4608 (N_4608,N_4013,N_4345);
and U4609 (N_4609,N_4442,N_4452);
nand U4610 (N_4610,N_4006,N_4334);
or U4611 (N_4611,N_4237,N_4255);
nand U4612 (N_4612,N_4174,N_4373);
and U4613 (N_4613,N_4443,N_4135);
and U4614 (N_4614,N_4331,N_4256);
xor U4615 (N_4615,N_4209,N_4354);
nand U4616 (N_4616,N_4168,N_4462);
and U4617 (N_4617,N_4387,N_4440);
and U4618 (N_4618,N_4370,N_4226);
xor U4619 (N_4619,N_4279,N_4141);
and U4620 (N_4620,N_4445,N_4455);
nand U4621 (N_4621,N_4352,N_4170);
nor U4622 (N_4622,N_4196,N_4400);
xor U4623 (N_4623,N_4086,N_4041);
nand U4624 (N_4624,N_4496,N_4029);
xor U4625 (N_4625,N_4129,N_4246);
xor U4626 (N_4626,N_4267,N_4153);
and U4627 (N_4627,N_4437,N_4394);
nand U4628 (N_4628,N_4243,N_4367);
xor U4629 (N_4629,N_4478,N_4176);
nand U4630 (N_4630,N_4089,N_4145);
and U4631 (N_4631,N_4439,N_4008);
xnor U4632 (N_4632,N_4441,N_4479);
or U4633 (N_4633,N_4032,N_4087);
and U4634 (N_4634,N_4101,N_4297);
nor U4635 (N_4635,N_4249,N_4128);
nand U4636 (N_4636,N_4432,N_4493);
xnor U4637 (N_4637,N_4166,N_4434);
and U4638 (N_4638,N_4274,N_4417);
nor U4639 (N_4639,N_4464,N_4306);
or U4640 (N_4640,N_4050,N_4038);
and U4641 (N_4641,N_4282,N_4037);
nor U4642 (N_4642,N_4285,N_4120);
nand U4643 (N_4643,N_4424,N_4025);
and U4644 (N_4644,N_4124,N_4079);
nor U4645 (N_4645,N_4023,N_4109);
nand U4646 (N_4646,N_4402,N_4069);
xnor U4647 (N_4647,N_4408,N_4254);
nor U4648 (N_4648,N_4327,N_4119);
or U4649 (N_4649,N_4138,N_4093);
nand U4650 (N_4650,N_4082,N_4293);
or U4651 (N_4651,N_4229,N_4134);
or U4652 (N_4652,N_4117,N_4311);
xnor U4653 (N_4653,N_4289,N_4190);
nor U4654 (N_4654,N_4356,N_4372);
or U4655 (N_4655,N_4171,N_4191);
nor U4656 (N_4656,N_4483,N_4451);
xor U4657 (N_4657,N_4064,N_4244);
nor U4658 (N_4658,N_4221,N_4276);
nand U4659 (N_4659,N_4465,N_4292);
nand U4660 (N_4660,N_4107,N_4043);
and U4661 (N_4661,N_4088,N_4428);
nor U4662 (N_4662,N_4225,N_4147);
nor U4663 (N_4663,N_4184,N_4458);
nand U4664 (N_4664,N_4217,N_4388);
and U4665 (N_4665,N_4091,N_4096);
and U4666 (N_4666,N_4346,N_4163);
xnor U4667 (N_4667,N_4178,N_4233);
nor U4668 (N_4668,N_4463,N_4142);
and U4669 (N_4669,N_4065,N_4466);
or U4670 (N_4670,N_4404,N_4189);
nor U4671 (N_4671,N_4257,N_4481);
xnor U4672 (N_4672,N_4447,N_4377);
xor U4673 (N_4673,N_4067,N_4485);
and U4674 (N_4674,N_4231,N_4181);
nand U4675 (N_4675,N_4084,N_4376);
nor U4676 (N_4676,N_4048,N_4131);
and U4677 (N_4677,N_4438,N_4467);
nand U4678 (N_4678,N_4425,N_4062);
xor U4679 (N_4679,N_4308,N_4172);
and U4680 (N_4680,N_4186,N_4368);
and U4681 (N_4681,N_4427,N_4004);
or U4682 (N_4682,N_4338,N_4219);
or U4683 (N_4683,N_4152,N_4342);
or U4684 (N_4684,N_4259,N_4296);
xnor U4685 (N_4685,N_4391,N_4313);
and U4686 (N_4686,N_4175,N_4137);
nor U4687 (N_4687,N_4403,N_4253);
nor U4688 (N_4688,N_4099,N_4028);
xnor U4689 (N_4689,N_4305,N_4260);
or U4690 (N_4690,N_4164,N_4183);
nand U4691 (N_4691,N_4261,N_4414);
nand U4692 (N_4692,N_4075,N_4482);
nand U4693 (N_4693,N_4460,N_4247);
nand U4694 (N_4694,N_4001,N_4116);
nand U4695 (N_4695,N_4205,N_4090);
nor U4696 (N_4696,N_4097,N_4347);
and U4697 (N_4697,N_4426,N_4492);
nand U4698 (N_4698,N_4187,N_4118);
xnor U4699 (N_4699,N_4489,N_4083);
xnor U4700 (N_4700,N_4343,N_4281);
or U4701 (N_4701,N_4010,N_4076);
nand U4702 (N_4702,N_4383,N_4074);
nand U4703 (N_4703,N_4486,N_4122);
and U4704 (N_4704,N_4298,N_4241);
nor U4705 (N_4705,N_4429,N_4112);
and U4706 (N_4706,N_4242,N_4339);
xor U4707 (N_4707,N_4380,N_4182);
xnor U4708 (N_4708,N_4114,N_4085);
and U4709 (N_4709,N_4382,N_4100);
and U4710 (N_4710,N_4328,N_4058);
nand U4711 (N_4711,N_4111,N_4324);
nor U4712 (N_4712,N_4284,N_4273);
nand U4713 (N_4713,N_4490,N_4133);
nand U4714 (N_4714,N_4002,N_4315);
and U4715 (N_4715,N_4095,N_4177);
and U4716 (N_4716,N_4271,N_4336);
nor U4717 (N_4717,N_4488,N_4139);
and U4718 (N_4718,N_4357,N_4421);
and U4719 (N_4719,N_4053,N_4238);
or U4720 (N_4720,N_4363,N_4159);
nand U4721 (N_4721,N_4491,N_4310);
xnor U4722 (N_4722,N_4287,N_4200);
nor U4723 (N_4723,N_4469,N_4318);
nand U4724 (N_4724,N_4015,N_4312);
nor U4725 (N_4725,N_4329,N_4169);
or U4726 (N_4726,N_4406,N_4245);
and U4727 (N_4727,N_4024,N_4389);
and U4728 (N_4728,N_4386,N_4494);
xnor U4729 (N_4729,N_4054,N_4211);
nand U4730 (N_4730,N_4361,N_4457);
and U4731 (N_4731,N_4415,N_4017);
and U4732 (N_4732,N_4307,N_4215);
xor U4733 (N_4733,N_4180,N_4148);
and U4734 (N_4734,N_4234,N_4459);
xor U4735 (N_4735,N_4036,N_4450);
and U4736 (N_4736,N_4272,N_4206);
nand U4737 (N_4737,N_4291,N_4060);
or U4738 (N_4738,N_4369,N_4418);
and U4739 (N_4739,N_4136,N_4167);
xnor U4740 (N_4740,N_4337,N_4456);
xor U4741 (N_4741,N_4268,N_4499);
and U4742 (N_4742,N_4044,N_4031);
nand U4743 (N_4743,N_4080,N_4444);
or U4744 (N_4744,N_4146,N_4210);
nand U4745 (N_4745,N_4278,N_4473);
nor U4746 (N_4746,N_4199,N_4070);
or U4747 (N_4747,N_4351,N_4213);
nand U4748 (N_4748,N_4392,N_4355);
or U4749 (N_4749,N_4401,N_4149);
xor U4750 (N_4750,N_4227,N_4377);
nand U4751 (N_4751,N_4342,N_4061);
and U4752 (N_4752,N_4388,N_4448);
and U4753 (N_4753,N_4221,N_4013);
or U4754 (N_4754,N_4341,N_4444);
nor U4755 (N_4755,N_4473,N_4009);
nand U4756 (N_4756,N_4469,N_4355);
xnor U4757 (N_4757,N_4455,N_4197);
nor U4758 (N_4758,N_4384,N_4129);
or U4759 (N_4759,N_4321,N_4246);
xor U4760 (N_4760,N_4371,N_4373);
or U4761 (N_4761,N_4223,N_4338);
xnor U4762 (N_4762,N_4389,N_4328);
or U4763 (N_4763,N_4466,N_4308);
nor U4764 (N_4764,N_4450,N_4057);
nand U4765 (N_4765,N_4269,N_4160);
nand U4766 (N_4766,N_4025,N_4224);
nor U4767 (N_4767,N_4247,N_4444);
nor U4768 (N_4768,N_4482,N_4424);
and U4769 (N_4769,N_4021,N_4225);
and U4770 (N_4770,N_4194,N_4189);
nand U4771 (N_4771,N_4311,N_4211);
xnor U4772 (N_4772,N_4225,N_4436);
nand U4773 (N_4773,N_4218,N_4058);
nand U4774 (N_4774,N_4058,N_4147);
or U4775 (N_4775,N_4322,N_4270);
xor U4776 (N_4776,N_4044,N_4077);
xor U4777 (N_4777,N_4427,N_4343);
and U4778 (N_4778,N_4183,N_4301);
nand U4779 (N_4779,N_4044,N_4221);
or U4780 (N_4780,N_4185,N_4453);
nor U4781 (N_4781,N_4209,N_4364);
nor U4782 (N_4782,N_4365,N_4243);
and U4783 (N_4783,N_4292,N_4149);
nand U4784 (N_4784,N_4413,N_4045);
xnor U4785 (N_4785,N_4243,N_4095);
and U4786 (N_4786,N_4341,N_4064);
or U4787 (N_4787,N_4398,N_4142);
or U4788 (N_4788,N_4047,N_4199);
or U4789 (N_4789,N_4153,N_4107);
nand U4790 (N_4790,N_4201,N_4155);
nor U4791 (N_4791,N_4051,N_4264);
and U4792 (N_4792,N_4464,N_4068);
and U4793 (N_4793,N_4456,N_4148);
or U4794 (N_4794,N_4446,N_4219);
nor U4795 (N_4795,N_4293,N_4219);
or U4796 (N_4796,N_4486,N_4493);
nor U4797 (N_4797,N_4223,N_4016);
xor U4798 (N_4798,N_4289,N_4420);
nand U4799 (N_4799,N_4454,N_4315);
nand U4800 (N_4800,N_4399,N_4371);
or U4801 (N_4801,N_4007,N_4272);
and U4802 (N_4802,N_4435,N_4448);
or U4803 (N_4803,N_4287,N_4230);
nor U4804 (N_4804,N_4381,N_4376);
xnor U4805 (N_4805,N_4390,N_4247);
nor U4806 (N_4806,N_4286,N_4266);
or U4807 (N_4807,N_4025,N_4362);
or U4808 (N_4808,N_4479,N_4141);
xnor U4809 (N_4809,N_4100,N_4400);
nand U4810 (N_4810,N_4191,N_4310);
nand U4811 (N_4811,N_4439,N_4309);
xor U4812 (N_4812,N_4149,N_4057);
xor U4813 (N_4813,N_4426,N_4345);
and U4814 (N_4814,N_4230,N_4257);
and U4815 (N_4815,N_4179,N_4467);
xor U4816 (N_4816,N_4211,N_4419);
nand U4817 (N_4817,N_4410,N_4003);
nand U4818 (N_4818,N_4305,N_4384);
xnor U4819 (N_4819,N_4290,N_4165);
and U4820 (N_4820,N_4194,N_4282);
or U4821 (N_4821,N_4275,N_4499);
xnor U4822 (N_4822,N_4003,N_4218);
xor U4823 (N_4823,N_4242,N_4174);
nand U4824 (N_4824,N_4493,N_4174);
nand U4825 (N_4825,N_4367,N_4021);
and U4826 (N_4826,N_4306,N_4066);
xor U4827 (N_4827,N_4226,N_4189);
xnor U4828 (N_4828,N_4459,N_4145);
nor U4829 (N_4829,N_4371,N_4129);
nand U4830 (N_4830,N_4088,N_4402);
or U4831 (N_4831,N_4144,N_4194);
nor U4832 (N_4832,N_4431,N_4244);
nor U4833 (N_4833,N_4070,N_4003);
and U4834 (N_4834,N_4127,N_4274);
or U4835 (N_4835,N_4334,N_4097);
nor U4836 (N_4836,N_4490,N_4255);
nand U4837 (N_4837,N_4225,N_4111);
or U4838 (N_4838,N_4438,N_4121);
and U4839 (N_4839,N_4352,N_4112);
or U4840 (N_4840,N_4210,N_4080);
nand U4841 (N_4841,N_4286,N_4274);
xnor U4842 (N_4842,N_4010,N_4128);
xnor U4843 (N_4843,N_4373,N_4417);
and U4844 (N_4844,N_4405,N_4103);
and U4845 (N_4845,N_4371,N_4175);
or U4846 (N_4846,N_4062,N_4357);
xor U4847 (N_4847,N_4428,N_4465);
and U4848 (N_4848,N_4151,N_4488);
and U4849 (N_4849,N_4279,N_4153);
nand U4850 (N_4850,N_4191,N_4006);
or U4851 (N_4851,N_4284,N_4445);
and U4852 (N_4852,N_4167,N_4147);
nand U4853 (N_4853,N_4384,N_4445);
nand U4854 (N_4854,N_4447,N_4263);
nand U4855 (N_4855,N_4012,N_4030);
and U4856 (N_4856,N_4004,N_4290);
or U4857 (N_4857,N_4380,N_4029);
nand U4858 (N_4858,N_4495,N_4469);
xor U4859 (N_4859,N_4263,N_4396);
and U4860 (N_4860,N_4483,N_4408);
or U4861 (N_4861,N_4416,N_4359);
or U4862 (N_4862,N_4096,N_4124);
and U4863 (N_4863,N_4030,N_4383);
nor U4864 (N_4864,N_4439,N_4368);
nand U4865 (N_4865,N_4151,N_4410);
nor U4866 (N_4866,N_4339,N_4447);
and U4867 (N_4867,N_4456,N_4235);
nand U4868 (N_4868,N_4026,N_4314);
nor U4869 (N_4869,N_4297,N_4390);
xnor U4870 (N_4870,N_4202,N_4422);
or U4871 (N_4871,N_4054,N_4017);
nor U4872 (N_4872,N_4346,N_4479);
and U4873 (N_4873,N_4063,N_4130);
or U4874 (N_4874,N_4024,N_4204);
nor U4875 (N_4875,N_4491,N_4199);
nand U4876 (N_4876,N_4069,N_4258);
or U4877 (N_4877,N_4065,N_4291);
and U4878 (N_4878,N_4301,N_4046);
nor U4879 (N_4879,N_4291,N_4450);
nor U4880 (N_4880,N_4323,N_4241);
nor U4881 (N_4881,N_4103,N_4090);
or U4882 (N_4882,N_4220,N_4167);
nor U4883 (N_4883,N_4377,N_4254);
xor U4884 (N_4884,N_4427,N_4339);
and U4885 (N_4885,N_4220,N_4481);
and U4886 (N_4886,N_4388,N_4371);
nor U4887 (N_4887,N_4251,N_4044);
nand U4888 (N_4888,N_4318,N_4488);
nand U4889 (N_4889,N_4244,N_4243);
nor U4890 (N_4890,N_4253,N_4260);
nand U4891 (N_4891,N_4406,N_4095);
and U4892 (N_4892,N_4152,N_4195);
nand U4893 (N_4893,N_4203,N_4015);
and U4894 (N_4894,N_4272,N_4303);
or U4895 (N_4895,N_4150,N_4448);
xor U4896 (N_4896,N_4404,N_4241);
nand U4897 (N_4897,N_4159,N_4386);
nor U4898 (N_4898,N_4185,N_4053);
and U4899 (N_4899,N_4194,N_4020);
nor U4900 (N_4900,N_4284,N_4499);
nor U4901 (N_4901,N_4367,N_4164);
xor U4902 (N_4902,N_4306,N_4151);
nand U4903 (N_4903,N_4385,N_4365);
nor U4904 (N_4904,N_4099,N_4065);
nor U4905 (N_4905,N_4471,N_4307);
nor U4906 (N_4906,N_4116,N_4077);
and U4907 (N_4907,N_4084,N_4098);
nor U4908 (N_4908,N_4491,N_4406);
nor U4909 (N_4909,N_4087,N_4365);
xnor U4910 (N_4910,N_4080,N_4199);
nand U4911 (N_4911,N_4318,N_4316);
nor U4912 (N_4912,N_4407,N_4256);
nand U4913 (N_4913,N_4139,N_4228);
and U4914 (N_4914,N_4004,N_4412);
and U4915 (N_4915,N_4338,N_4329);
xor U4916 (N_4916,N_4497,N_4179);
xnor U4917 (N_4917,N_4021,N_4269);
xor U4918 (N_4918,N_4427,N_4263);
or U4919 (N_4919,N_4460,N_4039);
nand U4920 (N_4920,N_4469,N_4239);
nor U4921 (N_4921,N_4096,N_4262);
nor U4922 (N_4922,N_4198,N_4277);
and U4923 (N_4923,N_4013,N_4115);
xnor U4924 (N_4924,N_4490,N_4069);
nor U4925 (N_4925,N_4360,N_4146);
or U4926 (N_4926,N_4240,N_4035);
and U4927 (N_4927,N_4301,N_4254);
xor U4928 (N_4928,N_4433,N_4201);
nand U4929 (N_4929,N_4429,N_4217);
or U4930 (N_4930,N_4438,N_4406);
nand U4931 (N_4931,N_4419,N_4038);
nand U4932 (N_4932,N_4136,N_4296);
and U4933 (N_4933,N_4475,N_4344);
nand U4934 (N_4934,N_4434,N_4436);
nand U4935 (N_4935,N_4221,N_4215);
nand U4936 (N_4936,N_4095,N_4071);
nor U4937 (N_4937,N_4050,N_4348);
nand U4938 (N_4938,N_4442,N_4091);
nor U4939 (N_4939,N_4169,N_4042);
or U4940 (N_4940,N_4137,N_4484);
xor U4941 (N_4941,N_4237,N_4352);
nor U4942 (N_4942,N_4241,N_4441);
nand U4943 (N_4943,N_4084,N_4159);
and U4944 (N_4944,N_4378,N_4409);
xnor U4945 (N_4945,N_4122,N_4313);
nor U4946 (N_4946,N_4128,N_4377);
or U4947 (N_4947,N_4275,N_4237);
nor U4948 (N_4948,N_4102,N_4292);
and U4949 (N_4949,N_4344,N_4065);
nor U4950 (N_4950,N_4393,N_4482);
nand U4951 (N_4951,N_4064,N_4053);
nor U4952 (N_4952,N_4060,N_4497);
nor U4953 (N_4953,N_4031,N_4436);
or U4954 (N_4954,N_4122,N_4389);
or U4955 (N_4955,N_4031,N_4314);
xor U4956 (N_4956,N_4043,N_4042);
nand U4957 (N_4957,N_4475,N_4267);
xnor U4958 (N_4958,N_4129,N_4285);
nand U4959 (N_4959,N_4021,N_4326);
or U4960 (N_4960,N_4114,N_4339);
nor U4961 (N_4961,N_4165,N_4127);
nand U4962 (N_4962,N_4257,N_4039);
nand U4963 (N_4963,N_4366,N_4436);
nor U4964 (N_4964,N_4174,N_4186);
nor U4965 (N_4965,N_4491,N_4188);
or U4966 (N_4966,N_4020,N_4450);
nor U4967 (N_4967,N_4472,N_4477);
nor U4968 (N_4968,N_4218,N_4336);
and U4969 (N_4969,N_4334,N_4081);
or U4970 (N_4970,N_4039,N_4311);
nor U4971 (N_4971,N_4108,N_4065);
nor U4972 (N_4972,N_4179,N_4344);
xnor U4973 (N_4973,N_4367,N_4189);
or U4974 (N_4974,N_4277,N_4304);
nand U4975 (N_4975,N_4090,N_4461);
xor U4976 (N_4976,N_4239,N_4124);
nand U4977 (N_4977,N_4021,N_4426);
and U4978 (N_4978,N_4171,N_4166);
nand U4979 (N_4979,N_4151,N_4162);
nor U4980 (N_4980,N_4458,N_4464);
and U4981 (N_4981,N_4080,N_4408);
or U4982 (N_4982,N_4111,N_4488);
and U4983 (N_4983,N_4474,N_4071);
or U4984 (N_4984,N_4485,N_4130);
nor U4985 (N_4985,N_4312,N_4440);
xor U4986 (N_4986,N_4044,N_4054);
or U4987 (N_4987,N_4025,N_4318);
or U4988 (N_4988,N_4135,N_4122);
xor U4989 (N_4989,N_4057,N_4076);
nor U4990 (N_4990,N_4249,N_4085);
or U4991 (N_4991,N_4389,N_4079);
or U4992 (N_4992,N_4189,N_4358);
nor U4993 (N_4993,N_4332,N_4272);
or U4994 (N_4994,N_4307,N_4230);
nand U4995 (N_4995,N_4407,N_4201);
xor U4996 (N_4996,N_4281,N_4331);
or U4997 (N_4997,N_4273,N_4494);
or U4998 (N_4998,N_4499,N_4377);
nor U4999 (N_4999,N_4338,N_4416);
xor U5000 (N_5000,N_4763,N_4584);
or U5001 (N_5001,N_4708,N_4932);
nand U5002 (N_5002,N_4614,N_4977);
nor U5003 (N_5003,N_4827,N_4762);
or U5004 (N_5004,N_4947,N_4743);
and U5005 (N_5005,N_4590,N_4722);
or U5006 (N_5006,N_4570,N_4839);
xnor U5007 (N_5007,N_4903,N_4557);
nand U5008 (N_5008,N_4600,N_4595);
nand U5009 (N_5009,N_4807,N_4967);
nand U5010 (N_5010,N_4801,N_4703);
nand U5011 (N_5011,N_4976,N_4825);
xnor U5012 (N_5012,N_4921,N_4504);
xor U5013 (N_5013,N_4653,N_4820);
and U5014 (N_5014,N_4935,N_4870);
or U5015 (N_5015,N_4605,N_4723);
or U5016 (N_5016,N_4919,N_4960);
and U5017 (N_5017,N_4786,N_4791);
nand U5018 (N_5018,N_4568,N_4877);
nor U5019 (N_5019,N_4618,N_4757);
nor U5020 (N_5020,N_4929,N_4729);
or U5021 (N_5021,N_4980,N_4580);
and U5022 (N_5022,N_4565,N_4830);
xnor U5023 (N_5023,N_4965,N_4968);
xnor U5024 (N_5024,N_4519,N_4576);
xor U5025 (N_5025,N_4928,N_4783);
or U5026 (N_5026,N_4892,N_4668);
nor U5027 (N_5027,N_4842,N_4750);
xnor U5028 (N_5028,N_4507,N_4710);
xnor U5029 (N_5029,N_4758,N_4661);
nor U5030 (N_5030,N_4663,N_4948);
and U5031 (N_5031,N_4954,N_4598);
xnor U5032 (N_5032,N_4555,N_4901);
nand U5033 (N_5033,N_4690,N_4638);
and U5034 (N_5034,N_4829,N_4966);
or U5035 (N_5035,N_4814,N_4867);
nand U5036 (N_5036,N_4500,N_4567);
or U5037 (N_5037,N_4621,N_4677);
or U5038 (N_5038,N_4608,N_4549);
nor U5039 (N_5039,N_4637,N_4854);
nor U5040 (N_5040,N_4572,N_4607);
nand U5041 (N_5041,N_4551,N_4984);
xor U5042 (N_5042,N_4674,N_4738);
nor U5043 (N_5043,N_4756,N_4950);
or U5044 (N_5044,N_4823,N_4978);
and U5045 (N_5045,N_4896,N_4782);
xnor U5046 (N_5046,N_4724,N_4620);
nand U5047 (N_5047,N_4520,N_4752);
and U5048 (N_5048,N_4933,N_4619);
nor U5049 (N_5049,N_4588,N_4860);
or U5050 (N_5050,N_4720,N_4672);
xnor U5051 (N_5051,N_4794,N_4865);
nand U5052 (N_5052,N_4804,N_4671);
or U5053 (N_5053,N_4694,N_4678);
nor U5054 (N_5054,N_4734,N_4862);
nor U5055 (N_5055,N_4993,N_4546);
or U5056 (N_5056,N_4518,N_4644);
nand U5057 (N_5057,N_4913,N_4868);
or U5058 (N_5058,N_4925,N_4838);
xor U5059 (N_5059,N_4961,N_4628);
or U5060 (N_5060,N_4503,N_4955);
nand U5061 (N_5061,N_4821,N_4699);
nor U5062 (N_5062,N_4527,N_4872);
or U5063 (N_5063,N_4508,N_4983);
and U5064 (N_5064,N_4533,N_4949);
nand U5065 (N_5065,N_4866,N_4602);
or U5066 (N_5066,N_4880,N_4534);
or U5067 (N_5067,N_4806,N_4561);
or U5068 (N_5068,N_4995,N_4874);
nor U5069 (N_5069,N_4957,N_4630);
nand U5070 (N_5070,N_4819,N_4701);
and U5071 (N_5071,N_4936,N_4755);
nand U5072 (N_5072,N_4560,N_4767);
xor U5073 (N_5073,N_4837,N_4959);
xnor U5074 (N_5074,N_4698,N_4573);
or U5075 (N_5075,N_4731,N_4587);
nor U5076 (N_5076,N_4797,N_4943);
or U5077 (N_5077,N_4988,N_4869);
and U5078 (N_5078,N_4861,N_4654);
or U5079 (N_5079,N_4553,N_4737);
nor U5080 (N_5080,N_4716,N_4702);
or U5081 (N_5081,N_4548,N_4624);
xnor U5082 (N_5082,N_4646,N_4905);
nand U5083 (N_5083,N_4847,N_4704);
and U5084 (N_5084,N_4660,N_4617);
nor U5085 (N_5085,N_4652,N_4688);
or U5086 (N_5086,N_4835,N_4656);
xor U5087 (N_5087,N_4956,N_4585);
nor U5088 (N_5088,N_4680,N_4882);
nand U5089 (N_5089,N_4662,N_4958);
and U5090 (N_5090,N_4831,N_4664);
xor U5091 (N_5091,N_4840,N_4712);
xor U5092 (N_5092,N_4515,N_4883);
nor U5093 (N_5093,N_4878,N_4594);
nor U5094 (N_5094,N_4884,N_4769);
or U5095 (N_5095,N_4922,N_4506);
nor U5096 (N_5096,N_4593,N_4923);
nand U5097 (N_5097,N_4639,N_4599);
nand U5098 (N_5098,N_4986,N_4817);
or U5099 (N_5099,N_4626,N_4787);
and U5100 (N_5100,N_4937,N_4962);
nor U5101 (N_5101,N_4693,N_4574);
or U5102 (N_5102,N_4733,N_4981);
nand U5103 (N_5103,N_4773,N_4643);
nand U5104 (N_5104,N_4779,N_4985);
nor U5105 (N_5105,N_4824,N_4537);
nand U5106 (N_5106,N_4930,N_4924);
nand U5107 (N_5107,N_4843,N_4899);
and U5108 (N_5108,N_4864,N_4938);
and U5109 (N_5109,N_4834,N_4577);
or U5110 (N_5110,N_4741,N_4634);
xnor U5111 (N_5111,N_4761,N_4727);
or U5112 (N_5112,N_4625,N_4610);
and U5113 (N_5113,N_4718,N_4717);
nand U5114 (N_5114,N_4517,N_4784);
xor U5115 (N_5115,N_4990,N_4846);
nand U5116 (N_5116,N_4944,N_4902);
or U5117 (N_5117,N_4844,N_4751);
nor U5118 (N_5118,N_4973,N_4927);
xor U5119 (N_5119,N_4633,N_4525);
nand U5120 (N_5120,N_4885,N_4524);
nor U5121 (N_5121,N_4725,N_4915);
and U5122 (N_5122,N_4815,N_4550);
nand U5123 (N_5123,N_4640,N_4857);
nand U5124 (N_5124,N_4541,N_4647);
nand U5125 (N_5125,N_4895,N_4996);
or U5126 (N_5126,N_4645,N_4686);
and U5127 (N_5127,N_4754,N_4858);
nor U5128 (N_5128,N_4891,N_4951);
xor U5129 (N_5129,N_4953,N_4739);
xor U5130 (N_5130,N_4616,N_4730);
xor U5131 (N_5131,N_4681,N_4530);
nor U5132 (N_5132,N_4700,N_4871);
nand U5133 (N_5133,N_4676,N_4648);
and U5134 (N_5134,N_4516,N_4583);
or U5135 (N_5135,N_4531,N_4521);
or U5136 (N_5136,N_4657,N_4735);
nand U5137 (N_5137,N_4532,N_4604);
and U5138 (N_5138,N_4813,N_4900);
and U5139 (N_5139,N_4636,N_4582);
or U5140 (N_5140,N_4765,N_4746);
and U5141 (N_5141,N_4934,N_4649);
nor U5142 (N_5142,N_4513,N_4501);
or U5143 (N_5143,N_4818,N_4622);
xor U5144 (N_5144,N_4575,N_4912);
and U5145 (N_5145,N_4705,N_4796);
or U5146 (N_5146,N_4780,N_4997);
nand U5147 (N_5147,N_4691,N_4970);
xor U5148 (N_5148,N_4775,N_4897);
xnor U5149 (N_5149,N_4788,N_4963);
and U5150 (N_5150,N_4774,N_4706);
xnor U5151 (N_5151,N_4941,N_4766);
nand U5152 (N_5152,N_4719,N_4511);
or U5153 (N_5153,N_4799,N_4563);
nor U5154 (N_5154,N_4523,N_4969);
or U5155 (N_5155,N_4529,N_4514);
nand U5156 (N_5156,N_4918,N_4669);
nand U5157 (N_5157,N_4859,N_4785);
or U5158 (N_5158,N_4856,N_4512);
or U5159 (N_5159,N_4855,N_4790);
nor U5160 (N_5160,N_4655,N_4945);
nor U5161 (N_5161,N_4509,N_4697);
nor U5162 (N_5162,N_4778,N_4726);
and U5163 (N_5163,N_4659,N_4876);
and U5164 (N_5164,N_4836,N_4810);
and U5165 (N_5165,N_4873,N_4881);
xor U5166 (N_5166,N_4526,N_4745);
nor U5167 (N_5167,N_4714,N_4848);
nand U5168 (N_5168,N_4764,N_4771);
and U5169 (N_5169,N_4695,N_4850);
xor U5170 (N_5170,N_4792,N_4740);
and U5171 (N_5171,N_4890,N_4942);
nand U5172 (N_5172,N_4907,N_4502);
and U5173 (N_5173,N_4609,N_4849);
and U5174 (N_5174,N_4554,N_4781);
or U5175 (N_5175,N_4566,N_4545);
and U5176 (N_5176,N_4579,N_4736);
xnor U5177 (N_5177,N_4709,N_4994);
nor U5178 (N_5178,N_4651,N_4972);
and U5179 (N_5179,N_4615,N_4613);
and U5180 (N_5180,N_4558,N_4917);
xnor U5181 (N_5181,N_4991,N_4728);
xnor U5182 (N_5182,N_4887,N_4552);
and U5183 (N_5183,N_4789,N_4931);
nor U5184 (N_5184,N_4713,N_4793);
nand U5185 (N_5185,N_4581,N_4889);
xor U5186 (N_5186,N_4893,N_4603);
or U5187 (N_5187,N_4952,N_4528);
nand U5188 (N_5188,N_4998,N_4635);
and U5189 (N_5189,N_4732,N_4826);
and U5190 (N_5190,N_4845,N_4571);
and U5191 (N_5191,N_4665,N_4536);
nand U5192 (N_5192,N_4888,N_4667);
or U5193 (N_5193,N_4586,N_4592);
or U5194 (N_5194,N_4692,N_4753);
and U5195 (N_5195,N_4658,N_4776);
and U5196 (N_5196,N_4601,N_4627);
and U5197 (N_5197,N_4982,N_4898);
xnor U5198 (N_5198,N_4711,N_4682);
nor U5199 (N_5199,N_4777,N_4538);
xnor U5200 (N_5200,N_4852,N_4744);
nor U5201 (N_5201,N_4800,N_4910);
or U5202 (N_5202,N_4597,N_4591);
nand U5203 (N_5203,N_4908,N_4641);
or U5204 (N_5204,N_4920,N_4642);
xor U5205 (N_5205,N_4559,N_4768);
and U5206 (N_5206,N_4505,N_4612);
xnor U5207 (N_5207,N_4666,N_4770);
nor U5208 (N_5208,N_4675,N_4816);
and U5209 (N_5209,N_4543,N_4911);
or U5210 (N_5210,N_4759,N_4812);
nor U5211 (N_5211,N_4875,N_4886);
or U5212 (N_5212,N_4940,N_4879);
or U5213 (N_5213,N_4802,N_4894);
xnor U5214 (N_5214,N_4822,N_4679);
or U5215 (N_5215,N_4673,N_4670);
and U5216 (N_5216,N_4629,N_4811);
and U5217 (N_5217,N_4828,N_4510);
or U5218 (N_5218,N_4715,N_4544);
nor U5219 (N_5219,N_4999,N_4689);
nor U5220 (N_5220,N_4589,N_4721);
or U5221 (N_5221,N_4522,N_4684);
nand U5222 (N_5222,N_4987,N_4685);
xor U5223 (N_5223,N_4539,N_4904);
nor U5224 (N_5224,N_4749,N_4851);
xnor U5225 (N_5225,N_4803,N_4564);
nand U5226 (N_5226,N_4596,N_4989);
or U5227 (N_5227,N_4798,N_4542);
nand U5228 (N_5228,N_4562,N_4631);
and U5229 (N_5229,N_4650,N_4696);
nor U5230 (N_5230,N_4926,N_4556);
nand U5231 (N_5231,N_4748,N_4914);
nor U5232 (N_5232,N_4916,N_4687);
and U5233 (N_5233,N_4975,N_4853);
nor U5234 (N_5234,N_4611,N_4992);
xnor U5235 (N_5235,N_4578,N_4683);
or U5236 (N_5236,N_4632,N_4742);
nor U5237 (N_5237,N_4841,N_4569);
nor U5238 (N_5238,N_4795,N_4809);
and U5239 (N_5239,N_4808,N_4964);
nor U5240 (N_5240,N_4939,N_4974);
nor U5241 (N_5241,N_4971,N_4772);
nand U5242 (N_5242,N_4833,N_4707);
xor U5243 (N_5243,N_4906,N_4540);
nand U5244 (N_5244,N_4805,N_4606);
xor U5245 (N_5245,N_4747,N_4535);
xnor U5246 (N_5246,N_4832,N_4760);
xor U5247 (N_5247,N_4946,N_4979);
nand U5248 (N_5248,N_4909,N_4623);
and U5249 (N_5249,N_4863,N_4547);
or U5250 (N_5250,N_4544,N_4987);
nor U5251 (N_5251,N_4552,N_4923);
and U5252 (N_5252,N_4554,N_4504);
or U5253 (N_5253,N_4657,N_4898);
nor U5254 (N_5254,N_4932,N_4740);
xor U5255 (N_5255,N_4933,N_4549);
or U5256 (N_5256,N_4782,N_4708);
nor U5257 (N_5257,N_4529,N_4733);
nor U5258 (N_5258,N_4720,N_4540);
and U5259 (N_5259,N_4739,N_4655);
nand U5260 (N_5260,N_4571,N_4534);
and U5261 (N_5261,N_4558,N_4757);
xnor U5262 (N_5262,N_4666,N_4936);
nor U5263 (N_5263,N_4642,N_4935);
xnor U5264 (N_5264,N_4600,N_4552);
nand U5265 (N_5265,N_4736,N_4867);
xor U5266 (N_5266,N_4859,N_4616);
xor U5267 (N_5267,N_4864,N_4734);
xor U5268 (N_5268,N_4600,N_4934);
or U5269 (N_5269,N_4809,N_4652);
and U5270 (N_5270,N_4575,N_4516);
nor U5271 (N_5271,N_4806,N_4552);
xor U5272 (N_5272,N_4772,N_4742);
or U5273 (N_5273,N_4754,N_4948);
nor U5274 (N_5274,N_4549,N_4571);
xnor U5275 (N_5275,N_4899,N_4764);
xor U5276 (N_5276,N_4639,N_4783);
xnor U5277 (N_5277,N_4536,N_4738);
nor U5278 (N_5278,N_4964,N_4767);
nand U5279 (N_5279,N_4543,N_4619);
or U5280 (N_5280,N_4641,N_4936);
xnor U5281 (N_5281,N_4913,N_4826);
or U5282 (N_5282,N_4586,N_4539);
xor U5283 (N_5283,N_4872,N_4620);
and U5284 (N_5284,N_4918,N_4649);
and U5285 (N_5285,N_4816,N_4951);
or U5286 (N_5286,N_4883,N_4739);
or U5287 (N_5287,N_4572,N_4760);
xor U5288 (N_5288,N_4608,N_4644);
nand U5289 (N_5289,N_4926,N_4770);
xor U5290 (N_5290,N_4684,N_4601);
or U5291 (N_5291,N_4586,N_4587);
or U5292 (N_5292,N_4703,N_4836);
or U5293 (N_5293,N_4608,N_4741);
nand U5294 (N_5294,N_4503,N_4946);
xor U5295 (N_5295,N_4725,N_4639);
nor U5296 (N_5296,N_4679,N_4998);
and U5297 (N_5297,N_4557,N_4985);
or U5298 (N_5298,N_4575,N_4627);
nand U5299 (N_5299,N_4834,N_4966);
xor U5300 (N_5300,N_4592,N_4834);
or U5301 (N_5301,N_4788,N_4617);
and U5302 (N_5302,N_4817,N_4910);
or U5303 (N_5303,N_4810,N_4904);
nor U5304 (N_5304,N_4957,N_4980);
xor U5305 (N_5305,N_4864,N_4659);
nor U5306 (N_5306,N_4702,N_4828);
or U5307 (N_5307,N_4855,N_4715);
and U5308 (N_5308,N_4590,N_4833);
nor U5309 (N_5309,N_4687,N_4561);
xor U5310 (N_5310,N_4802,N_4922);
nor U5311 (N_5311,N_4751,N_4993);
and U5312 (N_5312,N_4954,N_4845);
xor U5313 (N_5313,N_4964,N_4925);
or U5314 (N_5314,N_4839,N_4958);
nor U5315 (N_5315,N_4904,N_4943);
nand U5316 (N_5316,N_4935,N_4762);
nor U5317 (N_5317,N_4689,N_4528);
nand U5318 (N_5318,N_4819,N_4559);
or U5319 (N_5319,N_4999,N_4722);
or U5320 (N_5320,N_4791,N_4879);
nand U5321 (N_5321,N_4549,N_4660);
nand U5322 (N_5322,N_4951,N_4958);
nor U5323 (N_5323,N_4788,N_4517);
and U5324 (N_5324,N_4849,N_4607);
xnor U5325 (N_5325,N_4617,N_4920);
xnor U5326 (N_5326,N_4824,N_4837);
nor U5327 (N_5327,N_4785,N_4917);
and U5328 (N_5328,N_4684,N_4774);
nand U5329 (N_5329,N_4672,N_4674);
and U5330 (N_5330,N_4624,N_4601);
nand U5331 (N_5331,N_4808,N_4867);
and U5332 (N_5332,N_4917,N_4654);
nand U5333 (N_5333,N_4968,N_4884);
and U5334 (N_5334,N_4920,N_4949);
xor U5335 (N_5335,N_4855,N_4596);
nand U5336 (N_5336,N_4968,N_4967);
nand U5337 (N_5337,N_4614,N_4924);
xnor U5338 (N_5338,N_4851,N_4782);
and U5339 (N_5339,N_4711,N_4789);
and U5340 (N_5340,N_4822,N_4751);
nand U5341 (N_5341,N_4991,N_4974);
or U5342 (N_5342,N_4928,N_4812);
or U5343 (N_5343,N_4516,N_4905);
nand U5344 (N_5344,N_4848,N_4630);
or U5345 (N_5345,N_4876,N_4809);
xnor U5346 (N_5346,N_4839,N_4528);
and U5347 (N_5347,N_4577,N_4926);
and U5348 (N_5348,N_4809,N_4600);
and U5349 (N_5349,N_4547,N_4524);
xnor U5350 (N_5350,N_4843,N_4842);
or U5351 (N_5351,N_4583,N_4867);
nor U5352 (N_5352,N_4566,N_4959);
xnor U5353 (N_5353,N_4568,N_4555);
and U5354 (N_5354,N_4996,N_4574);
or U5355 (N_5355,N_4792,N_4958);
nand U5356 (N_5356,N_4744,N_4631);
and U5357 (N_5357,N_4634,N_4961);
nor U5358 (N_5358,N_4755,N_4616);
xnor U5359 (N_5359,N_4634,N_4520);
and U5360 (N_5360,N_4792,N_4857);
and U5361 (N_5361,N_4619,N_4700);
xor U5362 (N_5362,N_4881,N_4610);
nand U5363 (N_5363,N_4999,N_4931);
nor U5364 (N_5364,N_4721,N_4530);
nand U5365 (N_5365,N_4666,N_4621);
and U5366 (N_5366,N_4899,N_4883);
or U5367 (N_5367,N_4987,N_4644);
or U5368 (N_5368,N_4570,N_4718);
nor U5369 (N_5369,N_4923,N_4514);
or U5370 (N_5370,N_4566,N_4853);
or U5371 (N_5371,N_4757,N_4643);
nor U5372 (N_5372,N_4715,N_4524);
and U5373 (N_5373,N_4547,N_4658);
or U5374 (N_5374,N_4751,N_4758);
and U5375 (N_5375,N_4857,N_4999);
and U5376 (N_5376,N_4648,N_4927);
nor U5377 (N_5377,N_4689,N_4880);
nand U5378 (N_5378,N_4627,N_4506);
xor U5379 (N_5379,N_4839,N_4564);
or U5380 (N_5380,N_4537,N_4589);
nand U5381 (N_5381,N_4688,N_4773);
nand U5382 (N_5382,N_4579,N_4516);
and U5383 (N_5383,N_4791,N_4537);
xor U5384 (N_5384,N_4537,N_4564);
nor U5385 (N_5385,N_4763,N_4989);
nor U5386 (N_5386,N_4779,N_4726);
nor U5387 (N_5387,N_4713,N_4915);
or U5388 (N_5388,N_4857,N_4572);
xor U5389 (N_5389,N_4539,N_4653);
nor U5390 (N_5390,N_4680,N_4962);
xor U5391 (N_5391,N_4982,N_4642);
nand U5392 (N_5392,N_4955,N_4509);
nor U5393 (N_5393,N_4969,N_4797);
xnor U5394 (N_5394,N_4970,N_4520);
nand U5395 (N_5395,N_4823,N_4986);
xor U5396 (N_5396,N_4762,N_4973);
or U5397 (N_5397,N_4759,N_4951);
nand U5398 (N_5398,N_4577,N_4758);
nand U5399 (N_5399,N_4712,N_4687);
nor U5400 (N_5400,N_4771,N_4920);
xnor U5401 (N_5401,N_4754,N_4598);
or U5402 (N_5402,N_4776,N_4932);
nor U5403 (N_5403,N_4501,N_4699);
and U5404 (N_5404,N_4933,N_4713);
xnor U5405 (N_5405,N_4557,N_4604);
and U5406 (N_5406,N_4867,N_4684);
xnor U5407 (N_5407,N_4941,N_4658);
or U5408 (N_5408,N_4514,N_4879);
xnor U5409 (N_5409,N_4860,N_4871);
or U5410 (N_5410,N_4571,N_4514);
nor U5411 (N_5411,N_4844,N_4569);
and U5412 (N_5412,N_4723,N_4797);
and U5413 (N_5413,N_4885,N_4519);
nor U5414 (N_5414,N_4708,N_4923);
or U5415 (N_5415,N_4855,N_4771);
xnor U5416 (N_5416,N_4700,N_4846);
nor U5417 (N_5417,N_4595,N_4852);
and U5418 (N_5418,N_4803,N_4798);
nor U5419 (N_5419,N_4882,N_4907);
nand U5420 (N_5420,N_4886,N_4792);
nand U5421 (N_5421,N_4960,N_4512);
nor U5422 (N_5422,N_4564,N_4613);
xnor U5423 (N_5423,N_4641,N_4644);
and U5424 (N_5424,N_4688,N_4839);
nor U5425 (N_5425,N_4925,N_4874);
and U5426 (N_5426,N_4856,N_4593);
xor U5427 (N_5427,N_4625,N_4861);
xnor U5428 (N_5428,N_4765,N_4570);
nand U5429 (N_5429,N_4742,N_4802);
nand U5430 (N_5430,N_4513,N_4896);
and U5431 (N_5431,N_4812,N_4938);
and U5432 (N_5432,N_4538,N_4663);
and U5433 (N_5433,N_4940,N_4853);
and U5434 (N_5434,N_4833,N_4545);
xnor U5435 (N_5435,N_4675,N_4998);
nand U5436 (N_5436,N_4945,N_4870);
nor U5437 (N_5437,N_4870,N_4507);
xor U5438 (N_5438,N_4556,N_4616);
xor U5439 (N_5439,N_4777,N_4958);
and U5440 (N_5440,N_4503,N_4696);
or U5441 (N_5441,N_4970,N_4949);
or U5442 (N_5442,N_4714,N_4960);
and U5443 (N_5443,N_4732,N_4873);
nor U5444 (N_5444,N_4754,N_4817);
nor U5445 (N_5445,N_4798,N_4899);
nand U5446 (N_5446,N_4515,N_4601);
and U5447 (N_5447,N_4513,N_4597);
and U5448 (N_5448,N_4809,N_4892);
xor U5449 (N_5449,N_4906,N_4883);
or U5450 (N_5450,N_4641,N_4562);
xnor U5451 (N_5451,N_4767,N_4671);
nand U5452 (N_5452,N_4828,N_4802);
xnor U5453 (N_5453,N_4963,N_4998);
and U5454 (N_5454,N_4812,N_4567);
nand U5455 (N_5455,N_4867,N_4648);
and U5456 (N_5456,N_4773,N_4964);
and U5457 (N_5457,N_4788,N_4959);
or U5458 (N_5458,N_4619,N_4660);
xor U5459 (N_5459,N_4697,N_4619);
xor U5460 (N_5460,N_4866,N_4765);
xor U5461 (N_5461,N_4635,N_4629);
or U5462 (N_5462,N_4778,N_4752);
nand U5463 (N_5463,N_4504,N_4518);
xor U5464 (N_5464,N_4830,N_4685);
xnor U5465 (N_5465,N_4843,N_4713);
nand U5466 (N_5466,N_4602,N_4539);
or U5467 (N_5467,N_4510,N_4710);
nand U5468 (N_5468,N_4557,N_4651);
nand U5469 (N_5469,N_4626,N_4600);
nor U5470 (N_5470,N_4514,N_4925);
nand U5471 (N_5471,N_4870,N_4987);
nor U5472 (N_5472,N_4873,N_4595);
nor U5473 (N_5473,N_4528,N_4663);
xor U5474 (N_5474,N_4547,N_4768);
nor U5475 (N_5475,N_4600,N_4771);
nor U5476 (N_5476,N_4742,N_4965);
nand U5477 (N_5477,N_4637,N_4547);
xnor U5478 (N_5478,N_4669,N_4826);
nor U5479 (N_5479,N_4623,N_4645);
xnor U5480 (N_5480,N_4671,N_4908);
or U5481 (N_5481,N_4690,N_4630);
nand U5482 (N_5482,N_4658,N_4520);
or U5483 (N_5483,N_4697,N_4910);
and U5484 (N_5484,N_4744,N_4824);
nor U5485 (N_5485,N_4700,N_4512);
nor U5486 (N_5486,N_4512,N_4833);
and U5487 (N_5487,N_4693,N_4994);
nand U5488 (N_5488,N_4933,N_4562);
and U5489 (N_5489,N_4984,N_4642);
xnor U5490 (N_5490,N_4639,N_4943);
nor U5491 (N_5491,N_4553,N_4986);
xnor U5492 (N_5492,N_4691,N_4887);
or U5493 (N_5493,N_4706,N_4576);
nor U5494 (N_5494,N_4925,N_4856);
or U5495 (N_5495,N_4849,N_4781);
or U5496 (N_5496,N_4683,N_4745);
and U5497 (N_5497,N_4637,N_4807);
and U5498 (N_5498,N_4670,N_4917);
or U5499 (N_5499,N_4884,N_4921);
or U5500 (N_5500,N_5200,N_5164);
and U5501 (N_5501,N_5397,N_5224);
nand U5502 (N_5502,N_5116,N_5080);
nor U5503 (N_5503,N_5068,N_5411);
or U5504 (N_5504,N_5028,N_5112);
nand U5505 (N_5505,N_5268,N_5439);
nand U5506 (N_5506,N_5421,N_5419);
nand U5507 (N_5507,N_5108,N_5212);
nand U5508 (N_5508,N_5223,N_5194);
nand U5509 (N_5509,N_5216,N_5002);
xnor U5510 (N_5510,N_5050,N_5434);
or U5511 (N_5511,N_5077,N_5408);
or U5512 (N_5512,N_5415,N_5204);
and U5513 (N_5513,N_5320,N_5088);
or U5514 (N_5514,N_5167,N_5140);
nand U5515 (N_5515,N_5329,N_5205);
and U5516 (N_5516,N_5151,N_5255);
nor U5517 (N_5517,N_5136,N_5407);
and U5518 (N_5518,N_5305,N_5250);
xnor U5519 (N_5519,N_5284,N_5190);
and U5520 (N_5520,N_5180,N_5213);
xor U5521 (N_5521,N_5176,N_5263);
and U5522 (N_5522,N_5006,N_5385);
xor U5523 (N_5523,N_5342,N_5131);
and U5524 (N_5524,N_5064,N_5048);
xnor U5525 (N_5525,N_5058,N_5008);
or U5526 (N_5526,N_5490,N_5285);
nand U5527 (N_5527,N_5466,N_5318);
nand U5528 (N_5528,N_5383,N_5471);
nor U5529 (N_5529,N_5307,N_5450);
nand U5530 (N_5530,N_5356,N_5147);
nor U5531 (N_5531,N_5161,N_5470);
or U5532 (N_5532,N_5106,N_5483);
nor U5533 (N_5533,N_5452,N_5481);
nand U5534 (N_5534,N_5267,N_5225);
and U5535 (N_5535,N_5179,N_5257);
or U5536 (N_5536,N_5114,N_5290);
and U5537 (N_5537,N_5403,N_5062);
nor U5538 (N_5538,N_5334,N_5226);
and U5539 (N_5539,N_5326,N_5299);
and U5540 (N_5540,N_5003,N_5322);
and U5541 (N_5541,N_5266,N_5429);
or U5542 (N_5542,N_5245,N_5492);
and U5543 (N_5543,N_5251,N_5443);
xor U5544 (N_5544,N_5377,N_5327);
or U5545 (N_5545,N_5096,N_5005);
or U5546 (N_5546,N_5037,N_5269);
or U5547 (N_5547,N_5402,N_5170);
nand U5548 (N_5548,N_5043,N_5217);
or U5549 (N_5549,N_5332,N_5085);
and U5550 (N_5550,N_5472,N_5172);
and U5551 (N_5551,N_5258,N_5132);
or U5552 (N_5552,N_5289,N_5244);
nor U5553 (N_5553,N_5261,N_5463);
or U5554 (N_5554,N_5484,N_5392);
nor U5555 (N_5555,N_5358,N_5345);
nand U5556 (N_5556,N_5207,N_5338);
and U5557 (N_5557,N_5348,N_5432);
nand U5558 (N_5558,N_5023,N_5174);
or U5559 (N_5559,N_5323,N_5294);
or U5560 (N_5560,N_5034,N_5486);
and U5561 (N_5561,N_5222,N_5365);
or U5562 (N_5562,N_5361,N_5124);
nand U5563 (N_5563,N_5182,N_5337);
xor U5564 (N_5564,N_5030,N_5083);
nor U5565 (N_5565,N_5369,N_5013);
and U5566 (N_5566,N_5293,N_5291);
nor U5567 (N_5567,N_5027,N_5070);
and U5568 (N_5568,N_5395,N_5390);
or U5569 (N_5569,N_5229,N_5409);
and U5570 (N_5570,N_5417,N_5047);
and U5571 (N_5571,N_5309,N_5391);
or U5572 (N_5572,N_5396,N_5275);
nand U5573 (N_5573,N_5456,N_5449);
nor U5574 (N_5574,N_5093,N_5115);
or U5575 (N_5575,N_5234,N_5061);
nor U5576 (N_5576,N_5451,N_5279);
nand U5577 (N_5577,N_5311,N_5335);
xor U5578 (N_5578,N_5160,N_5343);
nand U5579 (N_5579,N_5227,N_5134);
xnor U5580 (N_5580,N_5082,N_5230);
nand U5581 (N_5581,N_5295,N_5152);
xnor U5582 (N_5582,N_5087,N_5032);
and U5583 (N_5583,N_5150,N_5171);
or U5584 (N_5584,N_5435,N_5367);
and U5585 (N_5585,N_5253,N_5324);
or U5586 (N_5586,N_5495,N_5353);
and U5587 (N_5587,N_5328,N_5214);
or U5588 (N_5588,N_5110,N_5181);
xnor U5589 (N_5589,N_5312,N_5125);
nor U5590 (N_5590,N_5482,N_5094);
xnor U5591 (N_5591,N_5420,N_5376);
or U5592 (N_5592,N_5169,N_5412);
xor U5593 (N_5593,N_5394,N_5260);
nor U5594 (N_5594,N_5063,N_5319);
xnor U5595 (N_5595,N_5215,N_5233);
xnor U5596 (N_5596,N_5304,N_5236);
nor U5597 (N_5597,N_5431,N_5056);
or U5598 (N_5598,N_5464,N_5206);
nor U5599 (N_5599,N_5247,N_5398);
and U5600 (N_5600,N_5366,N_5388);
xor U5601 (N_5601,N_5145,N_5264);
or U5602 (N_5602,N_5044,N_5078);
xor U5603 (N_5603,N_5469,N_5441);
nand U5604 (N_5604,N_5098,N_5273);
or U5605 (N_5605,N_5011,N_5118);
or U5606 (N_5606,N_5177,N_5184);
and U5607 (N_5607,N_5404,N_5359);
nand U5608 (N_5608,N_5202,N_5079);
nor U5609 (N_5609,N_5102,N_5186);
or U5610 (N_5610,N_5221,N_5243);
or U5611 (N_5611,N_5235,N_5185);
and U5612 (N_5612,N_5040,N_5086);
and U5613 (N_5613,N_5113,N_5081);
xor U5614 (N_5614,N_5109,N_5026);
and U5615 (N_5615,N_5017,N_5178);
xnor U5616 (N_5616,N_5475,N_5331);
nand U5617 (N_5617,N_5371,N_5288);
or U5618 (N_5618,N_5137,N_5231);
and U5619 (N_5619,N_5209,N_5302);
nor U5620 (N_5620,N_5352,N_5380);
nand U5621 (N_5621,N_5135,N_5406);
and U5622 (N_5622,N_5042,N_5413);
nand U5623 (N_5623,N_5189,N_5347);
and U5624 (N_5624,N_5453,N_5091);
and U5625 (N_5625,N_5424,N_5461);
and U5626 (N_5626,N_5300,N_5423);
nand U5627 (N_5627,N_5467,N_5336);
or U5628 (N_5628,N_5485,N_5220);
xnor U5629 (N_5629,N_5121,N_5089);
nor U5630 (N_5630,N_5045,N_5072);
xnor U5631 (N_5631,N_5046,N_5122);
or U5632 (N_5632,N_5019,N_5198);
nor U5633 (N_5633,N_5433,N_5468);
xnor U5634 (N_5634,N_5281,N_5051);
xor U5635 (N_5635,N_5029,N_5237);
nand U5636 (N_5636,N_5210,N_5148);
nand U5637 (N_5637,N_5095,N_5344);
nand U5638 (N_5638,N_5310,N_5025);
nor U5639 (N_5639,N_5351,N_5022);
or U5640 (N_5640,N_5438,N_5455);
nor U5641 (N_5641,N_5370,N_5084);
nor U5642 (N_5642,N_5159,N_5035);
and U5643 (N_5643,N_5410,N_5036);
and U5644 (N_5644,N_5149,N_5308);
or U5645 (N_5645,N_5041,N_5350);
and U5646 (N_5646,N_5418,N_5049);
nor U5647 (N_5647,N_5071,N_5059);
nand U5648 (N_5648,N_5426,N_5057);
nor U5649 (N_5649,N_5203,N_5448);
xnor U5650 (N_5650,N_5054,N_5117);
nor U5651 (N_5651,N_5065,N_5321);
and U5652 (N_5652,N_5362,N_5066);
nor U5653 (N_5653,N_5239,N_5156);
nand U5654 (N_5654,N_5400,N_5489);
or U5655 (N_5655,N_5382,N_5497);
nor U5656 (N_5656,N_5020,N_5241);
xnor U5657 (N_5657,N_5018,N_5246);
xnor U5658 (N_5658,N_5414,N_5039);
nor U5659 (N_5659,N_5173,N_5364);
and U5660 (N_5660,N_5199,N_5462);
nand U5661 (N_5661,N_5249,N_5422);
xnor U5662 (N_5662,N_5254,N_5007);
or U5663 (N_5663,N_5010,N_5256);
and U5664 (N_5664,N_5447,N_5330);
and U5665 (N_5665,N_5103,N_5073);
nand U5666 (N_5666,N_5265,N_5069);
xor U5667 (N_5667,N_5012,N_5428);
and U5668 (N_5668,N_5168,N_5154);
or U5669 (N_5669,N_5274,N_5128);
nor U5670 (N_5670,N_5287,N_5141);
or U5671 (N_5671,N_5314,N_5496);
or U5672 (N_5672,N_5075,N_5191);
and U5673 (N_5673,N_5104,N_5143);
nor U5674 (N_5674,N_5060,N_5317);
nor U5675 (N_5675,N_5494,N_5357);
and U5676 (N_5676,N_5129,N_5446);
and U5677 (N_5677,N_5126,N_5240);
xnor U5678 (N_5678,N_5242,N_5127);
nor U5679 (N_5679,N_5133,N_5009);
and U5680 (N_5680,N_5457,N_5099);
xnor U5681 (N_5681,N_5120,N_5499);
nor U5682 (N_5682,N_5301,N_5437);
nand U5683 (N_5683,N_5473,N_5272);
and U5684 (N_5684,N_5399,N_5163);
and U5685 (N_5685,N_5092,N_5107);
or U5686 (N_5686,N_5297,N_5155);
xor U5687 (N_5687,N_5487,N_5262);
nand U5688 (N_5688,N_5339,N_5393);
and U5689 (N_5689,N_5175,N_5349);
nand U5690 (N_5690,N_5031,N_5142);
and U5691 (N_5691,N_5074,N_5459);
or U5692 (N_5692,N_5100,N_5401);
nand U5693 (N_5693,N_5478,N_5090);
and U5694 (N_5694,N_5346,N_5021);
xor U5695 (N_5695,N_5123,N_5076);
xnor U5696 (N_5696,N_5296,N_5157);
nor U5697 (N_5697,N_5440,N_5333);
xnor U5698 (N_5698,N_5038,N_5378);
xnor U5699 (N_5699,N_5476,N_5477);
or U5700 (N_5700,N_5183,N_5201);
or U5701 (N_5701,N_5381,N_5219);
and U5702 (N_5702,N_5442,N_5354);
and U5703 (N_5703,N_5427,N_5014);
nand U5704 (N_5704,N_5303,N_5105);
nor U5705 (N_5705,N_5004,N_5416);
nand U5706 (N_5706,N_5144,N_5101);
xnor U5707 (N_5707,N_5444,N_5188);
or U5708 (N_5708,N_5196,N_5460);
nor U5709 (N_5709,N_5491,N_5479);
xor U5710 (N_5710,N_5052,N_5379);
or U5711 (N_5711,N_5368,N_5425);
or U5712 (N_5712,N_5454,N_5248);
and U5713 (N_5713,N_5016,N_5228);
nand U5714 (N_5714,N_5445,N_5197);
nand U5715 (N_5715,N_5341,N_5363);
xor U5716 (N_5716,N_5139,N_5373);
or U5717 (N_5717,N_5292,N_5372);
or U5718 (N_5718,N_5138,N_5192);
nor U5719 (N_5719,N_5286,N_5389);
nor U5720 (N_5720,N_5306,N_5280);
xor U5721 (N_5721,N_5465,N_5387);
and U5722 (N_5722,N_5000,N_5053);
and U5723 (N_5723,N_5430,N_5313);
nor U5724 (N_5724,N_5211,N_5187);
xor U5725 (N_5725,N_5015,N_5375);
xnor U5726 (N_5726,N_5283,N_5193);
nand U5727 (N_5727,N_5374,N_5355);
xnor U5728 (N_5728,N_5158,N_5232);
or U5729 (N_5729,N_5480,N_5316);
xnor U5730 (N_5730,N_5315,N_5119);
nor U5731 (N_5731,N_5153,N_5001);
xnor U5732 (N_5732,N_5282,N_5033);
xnor U5733 (N_5733,N_5298,N_5252);
or U5734 (N_5734,N_5360,N_5493);
or U5735 (N_5735,N_5218,N_5474);
nor U5736 (N_5736,N_5276,N_5340);
nand U5737 (N_5737,N_5195,N_5130);
xnor U5738 (N_5738,N_5498,N_5384);
xor U5739 (N_5739,N_5277,N_5067);
nor U5740 (N_5740,N_5270,N_5238);
and U5741 (N_5741,N_5278,N_5165);
xor U5742 (N_5742,N_5386,N_5111);
nand U5743 (N_5743,N_5325,N_5162);
nand U5744 (N_5744,N_5166,N_5436);
nand U5745 (N_5745,N_5024,N_5488);
nand U5746 (N_5746,N_5259,N_5405);
nand U5747 (N_5747,N_5097,N_5271);
nor U5748 (N_5748,N_5458,N_5146);
nand U5749 (N_5749,N_5055,N_5208);
and U5750 (N_5750,N_5470,N_5315);
and U5751 (N_5751,N_5411,N_5433);
or U5752 (N_5752,N_5299,N_5224);
xor U5753 (N_5753,N_5308,N_5330);
nand U5754 (N_5754,N_5239,N_5297);
and U5755 (N_5755,N_5231,N_5052);
nand U5756 (N_5756,N_5358,N_5377);
nor U5757 (N_5757,N_5419,N_5486);
xnor U5758 (N_5758,N_5427,N_5199);
xnor U5759 (N_5759,N_5003,N_5116);
or U5760 (N_5760,N_5436,N_5215);
or U5761 (N_5761,N_5146,N_5480);
nor U5762 (N_5762,N_5102,N_5324);
and U5763 (N_5763,N_5198,N_5044);
xnor U5764 (N_5764,N_5016,N_5031);
and U5765 (N_5765,N_5235,N_5254);
or U5766 (N_5766,N_5270,N_5109);
nor U5767 (N_5767,N_5128,N_5434);
xor U5768 (N_5768,N_5430,N_5471);
xor U5769 (N_5769,N_5327,N_5410);
or U5770 (N_5770,N_5131,N_5033);
nor U5771 (N_5771,N_5446,N_5119);
xnor U5772 (N_5772,N_5099,N_5024);
nand U5773 (N_5773,N_5477,N_5101);
and U5774 (N_5774,N_5424,N_5033);
nor U5775 (N_5775,N_5182,N_5474);
nor U5776 (N_5776,N_5362,N_5394);
nand U5777 (N_5777,N_5315,N_5342);
nand U5778 (N_5778,N_5093,N_5357);
nand U5779 (N_5779,N_5407,N_5481);
nor U5780 (N_5780,N_5289,N_5272);
and U5781 (N_5781,N_5084,N_5025);
nand U5782 (N_5782,N_5175,N_5133);
nor U5783 (N_5783,N_5000,N_5065);
xor U5784 (N_5784,N_5297,N_5003);
nor U5785 (N_5785,N_5386,N_5233);
nand U5786 (N_5786,N_5334,N_5308);
xor U5787 (N_5787,N_5279,N_5131);
nand U5788 (N_5788,N_5099,N_5359);
and U5789 (N_5789,N_5008,N_5196);
or U5790 (N_5790,N_5395,N_5445);
or U5791 (N_5791,N_5160,N_5282);
xnor U5792 (N_5792,N_5029,N_5308);
nand U5793 (N_5793,N_5354,N_5035);
and U5794 (N_5794,N_5237,N_5010);
or U5795 (N_5795,N_5110,N_5149);
and U5796 (N_5796,N_5059,N_5452);
nor U5797 (N_5797,N_5010,N_5423);
and U5798 (N_5798,N_5033,N_5466);
and U5799 (N_5799,N_5351,N_5031);
xnor U5800 (N_5800,N_5173,N_5181);
nand U5801 (N_5801,N_5203,N_5006);
xnor U5802 (N_5802,N_5183,N_5119);
or U5803 (N_5803,N_5033,N_5008);
nor U5804 (N_5804,N_5232,N_5491);
xnor U5805 (N_5805,N_5389,N_5435);
nand U5806 (N_5806,N_5166,N_5143);
or U5807 (N_5807,N_5379,N_5386);
nor U5808 (N_5808,N_5224,N_5230);
or U5809 (N_5809,N_5461,N_5490);
and U5810 (N_5810,N_5033,N_5065);
or U5811 (N_5811,N_5352,N_5366);
nor U5812 (N_5812,N_5266,N_5411);
and U5813 (N_5813,N_5027,N_5167);
nor U5814 (N_5814,N_5350,N_5187);
and U5815 (N_5815,N_5021,N_5260);
and U5816 (N_5816,N_5086,N_5023);
xnor U5817 (N_5817,N_5302,N_5006);
xnor U5818 (N_5818,N_5415,N_5004);
or U5819 (N_5819,N_5037,N_5376);
nand U5820 (N_5820,N_5156,N_5427);
xnor U5821 (N_5821,N_5213,N_5193);
or U5822 (N_5822,N_5288,N_5025);
and U5823 (N_5823,N_5425,N_5063);
xor U5824 (N_5824,N_5290,N_5392);
nor U5825 (N_5825,N_5040,N_5432);
and U5826 (N_5826,N_5196,N_5152);
nor U5827 (N_5827,N_5492,N_5257);
or U5828 (N_5828,N_5362,N_5072);
or U5829 (N_5829,N_5217,N_5033);
and U5830 (N_5830,N_5329,N_5091);
and U5831 (N_5831,N_5456,N_5156);
nor U5832 (N_5832,N_5393,N_5358);
and U5833 (N_5833,N_5161,N_5008);
or U5834 (N_5834,N_5466,N_5114);
and U5835 (N_5835,N_5074,N_5462);
nand U5836 (N_5836,N_5126,N_5296);
xnor U5837 (N_5837,N_5170,N_5133);
and U5838 (N_5838,N_5238,N_5051);
or U5839 (N_5839,N_5136,N_5231);
and U5840 (N_5840,N_5021,N_5227);
or U5841 (N_5841,N_5088,N_5189);
nand U5842 (N_5842,N_5270,N_5024);
and U5843 (N_5843,N_5139,N_5084);
and U5844 (N_5844,N_5064,N_5491);
or U5845 (N_5845,N_5281,N_5498);
and U5846 (N_5846,N_5415,N_5000);
xnor U5847 (N_5847,N_5118,N_5245);
nor U5848 (N_5848,N_5475,N_5381);
nand U5849 (N_5849,N_5382,N_5347);
or U5850 (N_5850,N_5478,N_5371);
or U5851 (N_5851,N_5490,N_5072);
nor U5852 (N_5852,N_5261,N_5447);
nand U5853 (N_5853,N_5104,N_5253);
nand U5854 (N_5854,N_5202,N_5137);
and U5855 (N_5855,N_5296,N_5430);
nand U5856 (N_5856,N_5110,N_5267);
xnor U5857 (N_5857,N_5417,N_5012);
nand U5858 (N_5858,N_5017,N_5495);
nor U5859 (N_5859,N_5400,N_5155);
xor U5860 (N_5860,N_5292,N_5214);
nor U5861 (N_5861,N_5491,N_5178);
nand U5862 (N_5862,N_5131,N_5312);
or U5863 (N_5863,N_5064,N_5476);
and U5864 (N_5864,N_5260,N_5209);
xnor U5865 (N_5865,N_5054,N_5099);
nor U5866 (N_5866,N_5280,N_5137);
nor U5867 (N_5867,N_5117,N_5187);
nor U5868 (N_5868,N_5328,N_5121);
and U5869 (N_5869,N_5393,N_5466);
xnor U5870 (N_5870,N_5152,N_5393);
xor U5871 (N_5871,N_5423,N_5060);
nor U5872 (N_5872,N_5228,N_5454);
nor U5873 (N_5873,N_5259,N_5009);
nor U5874 (N_5874,N_5291,N_5101);
nand U5875 (N_5875,N_5212,N_5104);
or U5876 (N_5876,N_5078,N_5363);
and U5877 (N_5877,N_5434,N_5227);
or U5878 (N_5878,N_5464,N_5454);
nand U5879 (N_5879,N_5429,N_5316);
xnor U5880 (N_5880,N_5459,N_5368);
xnor U5881 (N_5881,N_5290,N_5314);
nor U5882 (N_5882,N_5154,N_5128);
xor U5883 (N_5883,N_5129,N_5218);
xor U5884 (N_5884,N_5424,N_5203);
or U5885 (N_5885,N_5068,N_5222);
nand U5886 (N_5886,N_5408,N_5350);
xor U5887 (N_5887,N_5387,N_5096);
and U5888 (N_5888,N_5163,N_5455);
xor U5889 (N_5889,N_5047,N_5030);
or U5890 (N_5890,N_5391,N_5294);
and U5891 (N_5891,N_5337,N_5315);
and U5892 (N_5892,N_5306,N_5332);
xor U5893 (N_5893,N_5041,N_5202);
or U5894 (N_5894,N_5231,N_5036);
nor U5895 (N_5895,N_5433,N_5110);
xor U5896 (N_5896,N_5281,N_5381);
or U5897 (N_5897,N_5309,N_5135);
nor U5898 (N_5898,N_5147,N_5447);
nor U5899 (N_5899,N_5266,N_5434);
or U5900 (N_5900,N_5339,N_5008);
nor U5901 (N_5901,N_5263,N_5209);
and U5902 (N_5902,N_5493,N_5455);
nor U5903 (N_5903,N_5310,N_5442);
xnor U5904 (N_5904,N_5055,N_5002);
or U5905 (N_5905,N_5209,N_5355);
or U5906 (N_5906,N_5447,N_5457);
or U5907 (N_5907,N_5013,N_5420);
xnor U5908 (N_5908,N_5222,N_5469);
xor U5909 (N_5909,N_5221,N_5069);
nor U5910 (N_5910,N_5277,N_5187);
nand U5911 (N_5911,N_5056,N_5446);
and U5912 (N_5912,N_5425,N_5259);
and U5913 (N_5913,N_5386,N_5449);
or U5914 (N_5914,N_5363,N_5277);
or U5915 (N_5915,N_5296,N_5082);
nor U5916 (N_5916,N_5031,N_5284);
and U5917 (N_5917,N_5430,N_5218);
nand U5918 (N_5918,N_5130,N_5463);
nand U5919 (N_5919,N_5331,N_5239);
xor U5920 (N_5920,N_5261,N_5199);
nor U5921 (N_5921,N_5176,N_5105);
nor U5922 (N_5922,N_5310,N_5125);
and U5923 (N_5923,N_5042,N_5492);
or U5924 (N_5924,N_5187,N_5336);
and U5925 (N_5925,N_5120,N_5236);
nand U5926 (N_5926,N_5087,N_5487);
xnor U5927 (N_5927,N_5262,N_5175);
and U5928 (N_5928,N_5149,N_5132);
nand U5929 (N_5929,N_5182,N_5301);
xor U5930 (N_5930,N_5246,N_5116);
nand U5931 (N_5931,N_5373,N_5388);
xor U5932 (N_5932,N_5322,N_5400);
xnor U5933 (N_5933,N_5269,N_5499);
and U5934 (N_5934,N_5108,N_5391);
xor U5935 (N_5935,N_5402,N_5450);
or U5936 (N_5936,N_5149,N_5436);
nand U5937 (N_5937,N_5308,N_5449);
xnor U5938 (N_5938,N_5046,N_5269);
or U5939 (N_5939,N_5034,N_5360);
and U5940 (N_5940,N_5101,N_5339);
and U5941 (N_5941,N_5219,N_5359);
nor U5942 (N_5942,N_5311,N_5472);
or U5943 (N_5943,N_5074,N_5198);
nor U5944 (N_5944,N_5007,N_5016);
and U5945 (N_5945,N_5059,N_5488);
and U5946 (N_5946,N_5414,N_5328);
xor U5947 (N_5947,N_5307,N_5074);
or U5948 (N_5948,N_5300,N_5112);
xor U5949 (N_5949,N_5217,N_5034);
and U5950 (N_5950,N_5068,N_5237);
nand U5951 (N_5951,N_5377,N_5348);
or U5952 (N_5952,N_5308,N_5068);
xnor U5953 (N_5953,N_5082,N_5242);
xnor U5954 (N_5954,N_5475,N_5050);
or U5955 (N_5955,N_5007,N_5355);
and U5956 (N_5956,N_5442,N_5128);
or U5957 (N_5957,N_5148,N_5024);
and U5958 (N_5958,N_5252,N_5408);
nand U5959 (N_5959,N_5394,N_5237);
nor U5960 (N_5960,N_5454,N_5041);
or U5961 (N_5961,N_5087,N_5434);
or U5962 (N_5962,N_5185,N_5454);
or U5963 (N_5963,N_5037,N_5308);
and U5964 (N_5964,N_5113,N_5291);
xor U5965 (N_5965,N_5282,N_5185);
xnor U5966 (N_5966,N_5282,N_5275);
xor U5967 (N_5967,N_5192,N_5355);
nor U5968 (N_5968,N_5429,N_5322);
xnor U5969 (N_5969,N_5393,N_5405);
or U5970 (N_5970,N_5062,N_5290);
xnor U5971 (N_5971,N_5354,N_5369);
nand U5972 (N_5972,N_5399,N_5227);
or U5973 (N_5973,N_5439,N_5459);
xnor U5974 (N_5974,N_5116,N_5226);
or U5975 (N_5975,N_5214,N_5156);
or U5976 (N_5976,N_5336,N_5075);
or U5977 (N_5977,N_5446,N_5131);
or U5978 (N_5978,N_5168,N_5356);
or U5979 (N_5979,N_5386,N_5041);
nor U5980 (N_5980,N_5120,N_5275);
xor U5981 (N_5981,N_5445,N_5076);
nand U5982 (N_5982,N_5290,N_5498);
or U5983 (N_5983,N_5188,N_5152);
and U5984 (N_5984,N_5425,N_5497);
or U5985 (N_5985,N_5285,N_5435);
nand U5986 (N_5986,N_5437,N_5090);
nor U5987 (N_5987,N_5273,N_5206);
and U5988 (N_5988,N_5050,N_5181);
and U5989 (N_5989,N_5457,N_5458);
xnor U5990 (N_5990,N_5448,N_5148);
xor U5991 (N_5991,N_5266,N_5358);
and U5992 (N_5992,N_5184,N_5465);
and U5993 (N_5993,N_5151,N_5386);
xnor U5994 (N_5994,N_5430,N_5489);
and U5995 (N_5995,N_5386,N_5005);
xor U5996 (N_5996,N_5007,N_5350);
or U5997 (N_5997,N_5332,N_5182);
or U5998 (N_5998,N_5490,N_5422);
nand U5999 (N_5999,N_5258,N_5026);
nand U6000 (N_6000,N_5967,N_5558);
and U6001 (N_6001,N_5784,N_5753);
and U6002 (N_6002,N_5793,N_5681);
xor U6003 (N_6003,N_5723,N_5976);
xnor U6004 (N_6004,N_5633,N_5996);
and U6005 (N_6005,N_5594,N_5655);
nand U6006 (N_6006,N_5796,N_5981);
or U6007 (N_6007,N_5550,N_5649);
and U6008 (N_6008,N_5787,N_5674);
nand U6009 (N_6009,N_5794,N_5559);
nand U6010 (N_6010,N_5914,N_5581);
and U6011 (N_6011,N_5859,N_5819);
nor U6012 (N_6012,N_5809,N_5945);
nand U6013 (N_6013,N_5907,N_5733);
and U6014 (N_6014,N_5806,N_5864);
or U6015 (N_6015,N_5815,N_5802);
and U6016 (N_6016,N_5818,N_5837);
xor U6017 (N_6017,N_5648,N_5567);
or U6018 (N_6018,N_5952,N_5805);
xnor U6019 (N_6019,N_5552,N_5501);
or U6020 (N_6020,N_5947,N_5946);
nand U6021 (N_6021,N_5507,N_5771);
or U6022 (N_6022,N_5549,N_5894);
and U6023 (N_6023,N_5535,N_5988);
and U6024 (N_6024,N_5767,N_5642);
nand U6025 (N_6025,N_5697,N_5656);
or U6026 (N_6026,N_5643,N_5895);
or U6027 (N_6027,N_5726,N_5635);
or U6028 (N_6028,N_5951,N_5898);
and U6029 (N_6029,N_5950,N_5521);
nand U6030 (N_6030,N_5855,N_5523);
or U6031 (N_6031,N_5561,N_5932);
nand U6032 (N_6032,N_5536,N_5710);
nand U6033 (N_6033,N_5966,N_5740);
xnor U6034 (N_6034,N_5944,N_5694);
and U6035 (N_6035,N_5547,N_5530);
or U6036 (N_6036,N_5730,N_5964);
and U6037 (N_6037,N_5872,N_5798);
or U6038 (N_6038,N_5576,N_5638);
or U6039 (N_6039,N_5686,N_5687);
nand U6040 (N_6040,N_5644,N_5953);
nand U6041 (N_6041,N_5654,N_5678);
nand U6042 (N_6042,N_5579,N_5554);
nor U6043 (N_6043,N_5808,N_5690);
nand U6044 (N_6044,N_5537,N_5508);
or U6045 (N_6045,N_5799,N_5754);
and U6046 (N_6046,N_5738,N_5823);
nand U6047 (N_6047,N_5725,N_5543);
and U6048 (N_6048,N_5931,N_5789);
or U6049 (N_6049,N_5841,N_5857);
xnor U6050 (N_6050,N_5941,N_5689);
nor U6051 (N_6051,N_5908,N_5765);
xor U6052 (N_6052,N_5783,N_5748);
and U6053 (N_6053,N_5997,N_5595);
xor U6054 (N_6054,N_5620,N_5786);
and U6055 (N_6055,N_5705,N_5919);
nand U6056 (N_6056,N_5511,N_5875);
or U6057 (N_6057,N_5943,N_5604);
or U6058 (N_6058,N_5637,N_5848);
nor U6059 (N_6059,N_5890,N_5887);
xor U6060 (N_6060,N_5634,N_5948);
and U6061 (N_6061,N_5827,N_5528);
nor U6062 (N_6062,N_5551,N_5647);
and U6063 (N_6063,N_5957,N_5938);
nand U6064 (N_6064,N_5980,N_5760);
or U6065 (N_6065,N_5704,N_5514);
and U6066 (N_6066,N_5825,N_5830);
and U6067 (N_6067,N_5688,N_5795);
and U6068 (N_6068,N_5517,N_5540);
nor U6069 (N_6069,N_5628,N_5699);
xnor U6070 (N_6070,N_5824,N_5568);
or U6071 (N_6071,N_5846,N_5665);
or U6072 (N_6072,N_5928,N_5901);
or U6073 (N_6073,N_5608,N_5519);
nand U6074 (N_6074,N_5734,N_5987);
nor U6075 (N_6075,N_5813,N_5691);
and U6076 (N_6076,N_5556,N_5924);
and U6077 (N_6077,N_5842,N_5564);
nor U6078 (N_6078,N_5975,N_5539);
or U6079 (N_6079,N_5591,N_5971);
or U6080 (N_6080,N_5548,N_5743);
nor U6081 (N_6081,N_5879,N_5968);
and U6082 (N_6082,N_5553,N_5735);
and U6083 (N_6083,N_5820,N_5852);
xnor U6084 (N_6084,N_5916,N_5792);
nor U6085 (N_6085,N_5807,N_5741);
and U6086 (N_6086,N_5613,N_5700);
nand U6087 (N_6087,N_5949,N_5986);
and U6088 (N_6088,N_5565,N_5719);
and U6089 (N_6089,N_5926,N_5664);
and U6090 (N_6090,N_5758,N_5578);
or U6091 (N_6091,N_5526,N_5718);
nand U6092 (N_6092,N_5563,N_5627);
nand U6093 (N_6093,N_5516,N_5918);
nand U6094 (N_6094,N_5545,N_5600);
or U6095 (N_6095,N_5970,N_5961);
or U6096 (N_6096,N_5675,N_5520);
xor U6097 (N_6097,N_5874,N_5828);
nor U6098 (N_6098,N_5721,N_5869);
nor U6099 (N_6099,N_5587,N_5515);
nand U6100 (N_6100,N_5992,N_5920);
or U6101 (N_6101,N_5751,N_5598);
nand U6102 (N_6102,N_5937,N_5663);
nand U6103 (N_6103,N_5965,N_5821);
nand U6104 (N_6104,N_5892,N_5646);
nor U6105 (N_6105,N_5571,N_5847);
nor U6106 (N_6106,N_5863,N_5685);
or U6107 (N_6107,N_5676,N_5629);
xor U6108 (N_6108,N_5546,N_5666);
and U6109 (N_6109,N_5885,N_5990);
nand U6110 (N_6110,N_5876,N_5624);
and U6111 (N_6111,N_5702,N_5977);
nand U6112 (N_6112,N_5732,N_5707);
or U6113 (N_6113,N_5804,N_5601);
nand U6114 (N_6114,N_5695,N_5590);
or U6115 (N_6115,N_5871,N_5671);
nand U6116 (N_6116,N_5617,N_5762);
xor U6117 (N_6117,N_5673,N_5557);
nor U6118 (N_6118,N_5782,N_5715);
nor U6119 (N_6119,N_5877,N_5840);
and U6120 (N_6120,N_5903,N_5684);
and U6121 (N_6121,N_5929,N_5905);
and U6122 (N_6122,N_5881,N_5683);
and U6123 (N_6123,N_5983,N_5909);
nand U6124 (N_6124,N_5999,N_5641);
or U6125 (N_6125,N_5915,N_5816);
and U6126 (N_6126,N_5770,N_5882);
nand U6127 (N_6127,N_5921,N_5836);
nand U6128 (N_6128,N_5910,N_5614);
nand U6129 (N_6129,N_5845,N_5778);
or U6130 (N_6130,N_5737,N_5593);
nand U6131 (N_6131,N_5995,N_5714);
xnor U6132 (N_6132,N_5503,N_5883);
and U6133 (N_6133,N_5582,N_5693);
nand U6134 (N_6134,N_5619,N_5533);
and U6135 (N_6135,N_5831,N_5978);
xnor U6136 (N_6136,N_5630,N_5925);
nor U6137 (N_6137,N_5911,N_5788);
or U6138 (N_6138,N_5764,N_5658);
nor U6139 (N_6139,N_5870,N_5716);
and U6140 (N_6140,N_5667,N_5973);
nand U6141 (N_6141,N_5761,N_5505);
nor U6142 (N_6142,N_5660,N_5560);
nand U6143 (N_6143,N_5998,N_5574);
nand U6144 (N_6144,N_5592,N_5506);
nor U6145 (N_6145,N_5777,N_5917);
xor U6146 (N_6146,N_5755,N_5886);
nand U6147 (N_6147,N_5891,N_5853);
or U6148 (N_6148,N_5839,N_5680);
xnor U6149 (N_6149,N_5780,N_5766);
or U6150 (N_6150,N_5652,N_5622);
nand U6151 (N_6151,N_5812,N_5527);
nor U6152 (N_6152,N_5888,N_5974);
or U6153 (N_6153,N_5742,N_5989);
nor U6154 (N_6154,N_5960,N_5858);
nand U6155 (N_6155,N_5939,N_5868);
or U6156 (N_6156,N_5657,N_5889);
xnor U6157 (N_6157,N_5832,N_5509);
xor U6158 (N_6158,N_5711,N_5756);
xnor U6159 (N_6159,N_5833,N_5829);
or U6160 (N_6160,N_5724,N_5811);
and U6161 (N_6161,N_5736,N_5631);
nand U6162 (N_6162,N_5729,N_5902);
or U6163 (N_6163,N_5513,N_5822);
xnor U6164 (N_6164,N_5636,N_5942);
or U6165 (N_6165,N_5826,N_5851);
nor U6166 (N_6166,N_5612,N_5835);
nor U6167 (N_6167,N_5585,N_5569);
and U6168 (N_6168,N_5873,N_5679);
and U6169 (N_6169,N_5677,N_5906);
nand U6170 (N_6170,N_5645,N_5956);
nand U6171 (N_6171,N_5541,N_5984);
nor U6172 (N_6172,N_5534,N_5698);
xnor U6173 (N_6173,N_5745,N_5991);
or U6174 (N_6174,N_5632,N_5834);
and U6175 (N_6175,N_5927,N_5522);
nand U6176 (N_6176,N_5602,N_5555);
nor U6177 (N_6177,N_5797,N_5933);
xor U6178 (N_6178,N_5532,N_5512);
nand U6179 (N_6179,N_5640,N_5708);
nand U6180 (N_6180,N_5529,N_5650);
xor U6181 (N_6181,N_5800,N_5623);
or U6182 (N_6182,N_5713,N_5994);
xor U6183 (N_6183,N_5703,N_5790);
nor U6184 (N_6184,N_5959,N_5525);
nor U6185 (N_6185,N_5586,N_5934);
xnor U6186 (N_6186,N_5922,N_5566);
xnor U6187 (N_6187,N_5672,N_5862);
or U6188 (N_6188,N_5803,N_5639);
or U6189 (N_6189,N_5544,N_5781);
xnor U6190 (N_6190,N_5596,N_5954);
nor U6191 (N_6191,N_5731,N_5610);
or U6192 (N_6192,N_5768,N_5930);
xor U6193 (N_6193,N_5969,N_5940);
nand U6194 (N_6194,N_5861,N_5597);
xnor U6195 (N_6195,N_5720,N_5854);
or U6196 (N_6196,N_5860,N_5982);
and U6197 (N_6197,N_5609,N_5878);
nand U6198 (N_6198,N_5884,N_5856);
nand U6199 (N_6199,N_5744,N_5772);
and U6200 (N_6200,N_5570,N_5575);
xor U6201 (N_6201,N_5897,N_5615);
xnor U6202 (N_6202,N_5502,N_5573);
nand U6203 (N_6203,N_5746,N_5993);
xnor U6204 (N_6204,N_5577,N_5662);
nand U6205 (N_6205,N_5696,N_5606);
nor U6206 (N_6206,N_5923,N_5572);
xnor U6207 (N_6207,N_5936,N_5580);
xnor U6208 (N_6208,N_5867,N_5979);
xor U6209 (N_6209,N_5504,N_5801);
nand U6210 (N_6210,N_5599,N_5769);
xor U6211 (N_6211,N_5682,N_5712);
nor U6212 (N_6212,N_5893,N_5935);
nor U6213 (N_6213,N_5912,N_5814);
nand U6214 (N_6214,N_5701,N_5616);
xor U6215 (N_6215,N_5880,N_5651);
xor U6216 (N_6216,N_5817,N_5776);
nor U6217 (N_6217,N_5538,N_5749);
or U6218 (N_6218,N_5618,N_5589);
nor U6219 (N_6219,N_5562,N_5727);
xnor U6220 (N_6220,N_5518,N_5865);
nand U6221 (N_6221,N_5692,N_5785);
nand U6222 (N_6222,N_5670,N_5524);
and U6223 (N_6223,N_5850,N_5625);
xnor U6224 (N_6224,N_5626,N_5611);
or U6225 (N_6225,N_5605,N_5621);
xnor U6226 (N_6226,N_5774,N_5963);
xor U6227 (N_6227,N_5500,N_5913);
or U6228 (N_6228,N_5763,N_5899);
or U6229 (N_6229,N_5728,N_5752);
or U6230 (N_6230,N_5668,N_5773);
xnor U6231 (N_6231,N_5849,N_5588);
or U6232 (N_6232,N_5531,N_5709);
nand U6233 (N_6233,N_5653,N_5722);
xnor U6234 (N_6234,N_5542,N_5779);
and U6235 (N_6235,N_5661,N_5706);
or U6236 (N_6236,N_5985,N_5896);
and U6237 (N_6237,N_5659,N_5603);
nand U6238 (N_6238,N_5747,N_5583);
or U6239 (N_6239,N_5955,N_5510);
nand U6240 (N_6240,N_5739,N_5958);
nand U6241 (N_6241,N_5669,N_5843);
and U6242 (N_6242,N_5838,N_5810);
xor U6243 (N_6243,N_5584,N_5791);
or U6244 (N_6244,N_5775,N_5759);
xnor U6245 (N_6245,N_5717,N_5757);
or U6246 (N_6246,N_5750,N_5972);
nor U6247 (N_6247,N_5900,N_5844);
nand U6248 (N_6248,N_5904,N_5607);
nand U6249 (N_6249,N_5866,N_5962);
and U6250 (N_6250,N_5808,N_5937);
nor U6251 (N_6251,N_5670,N_5616);
xnor U6252 (N_6252,N_5953,N_5894);
nand U6253 (N_6253,N_5665,N_5893);
xnor U6254 (N_6254,N_5838,N_5731);
nand U6255 (N_6255,N_5743,N_5622);
xnor U6256 (N_6256,N_5695,N_5910);
nor U6257 (N_6257,N_5724,N_5526);
nor U6258 (N_6258,N_5742,N_5666);
or U6259 (N_6259,N_5629,N_5669);
nor U6260 (N_6260,N_5612,N_5950);
nand U6261 (N_6261,N_5679,N_5787);
nand U6262 (N_6262,N_5903,N_5879);
xor U6263 (N_6263,N_5943,N_5645);
and U6264 (N_6264,N_5707,N_5597);
and U6265 (N_6265,N_5704,N_5980);
nand U6266 (N_6266,N_5708,N_5786);
xor U6267 (N_6267,N_5844,N_5990);
and U6268 (N_6268,N_5728,N_5886);
nand U6269 (N_6269,N_5727,N_5720);
nand U6270 (N_6270,N_5892,N_5982);
and U6271 (N_6271,N_5736,N_5920);
and U6272 (N_6272,N_5789,N_5717);
nand U6273 (N_6273,N_5571,N_5893);
xor U6274 (N_6274,N_5567,N_5793);
nand U6275 (N_6275,N_5506,N_5842);
nor U6276 (N_6276,N_5873,N_5962);
nor U6277 (N_6277,N_5672,N_5595);
nand U6278 (N_6278,N_5807,N_5932);
nand U6279 (N_6279,N_5650,N_5843);
xnor U6280 (N_6280,N_5693,N_5534);
nor U6281 (N_6281,N_5608,N_5612);
and U6282 (N_6282,N_5883,N_5901);
nor U6283 (N_6283,N_5749,N_5745);
nor U6284 (N_6284,N_5808,N_5727);
or U6285 (N_6285,N_5892,N_5599);
nand U6286 (N_6286,N_5980,N_5776);
xor U6287 (N_6287,N_5820,N_5682);
nand U6288 (N_6288,N_5781,N_5706);
nor U6289 (N_6289,N_5973,N_5516);
nor U6290 (N_6290,N_5639,N_5501);
or U6291 (N_6291,N_5853,N_5897);
xnor U6292 (N_6292,N_5852,N_5653);
or U6293 (N_6293,N_5706,N_5875);
nand U6294 (N_6294,N_5738,N_5894);
and U6295 (N_6295,N_5618,N_5985);
or U6296 (N_6296,N_5860,N_5986);
xnor U6297 (N_6297,N_5695,N_5789);
and U6298 (N_6298,N_5729,N_5841);
nand U6299 (N_6299,N_5795,N_5660);
and U6300 (N_6300,N_5988,N_5993);
and U6301 (N_6301,N_5947,N_5716);
and U6302 (N_6302,N_5726,N_5767);
or U6303 (N_6303,N_5769,N_5836);
xnor U6304 (N_6304,N_5685,N_5648);
or U6305 (N_6305,N_5772,N_5519);
nor U6306 (N_6306,N_5888,N_5507);
xnor U6307 (N_6307,N_5641,N_5653);
nand U6308 (N_6308,N_5709,N_5775);
and U6309 (N_6309,N_5642,N_5587);
nand U6310 (N_6310,N_5538,N_5599);
nand U6311 (N_6311,N_5614,N_5828);
and U6312 (N_6312,N_5934,N_5513);
xnor U6313 (N_6313,N_5700,N_5702);
xor U6314 (N_6314,N_5952,N_5763);
nand U6315 (N_6315,N_5915,N_5532);
nor U6316 (N_6316,N_5724,N_5607);
or U6317 (N_6317,N_5561,N_5619);
nand U6318 (N_6318,N_5563,N_5793);
nor U6319 (N_6319,N_5819,N_5867);
and U6320 (N_6320,N_5520,N_5737);
nand U6321 (N_6321,N_5698,N_5563);
nand U6322 (N_6322,N_5972,N_5538);
xnor U6323 (N_6323,N_5706,N_5811);
and U6324 (N_6324,N_5664,N_5878);
nor U6325 (N_6325,N_5624,N_5588);
or U6326 (N_6326,N_5888,N_5667);
nor U6327 (N_6327,N_5504,N_5894);
and U6328 (N_6328,N_5772,N_5899);
and U6329 (N_6329,N_5519,N_5647);
and U6330 (N_6330,N_5761,N_5775);
and U6331 (N_6331,N_5518,N_5714);
or U6332 (N_6332,N_5752,N_5953);
nand U6333 (N_6333,N_5761,N_5531);
nand U6334 (N_6334,N_5912,N_5588);
or U6335 (N_6335,N_5980,N_5932);
and U6336 (N_6336,N_5897,N_5792);
and U6337 (N_6337,N_5751,N_5543);
nor U6338 (N_6338,N_5941,N_5922);
or U6339 (N_6339,N_5903,N_5973);
or U6340 (N_6340,N_5761,N_5537);
nor U6341 (N_6341,N_5805,N_5672);
and U6342 (N_6342,N_5806,N_5712);
or U6343 (N_6343,N_5522,N_5896);
xor U6344 (N_6344,N_5834,N_5639);
xnor U6345 (N_6345,N_5935,N_5627);
and U6346 (N_6346,N_5639,N_5918);
xnor U6347 (N_6347,N_5963,N_5586);
nor U6348 (N_6348,N_5963,N_5780);
nand U6349 (N_6349,N_5734,N_5796);
nand U6350 (N_6350,N_5998,N_5632);
or U6351 (N_6351,N_5798,N_5804);
and U6352 (N_6352,N_5744,N_5955);
xnor U6353 (N_6353,N_5724,N_5977);
xnor U6354 (N_6354,N_5591,N_5933);
nor U6355 (N_6355,N_5945,N_5562);
xor U6356 (N_6356,N_5797,N_5853);
and U6357 (N_6357,N_5556,N_5522);
or U6358 (N_6358,N_5937,N_5864);
nand U6359 (N_6359,N_5613,N_5761);
xnor U6360 (N_6360,N_5732,N_5972);
xnor U6361 (N_6361,N_5831,N_5973);
xnor U6362 (N_6362,N_5722,N_5960);
nor U6363 (N_6363,N_5561,N_5827);
or U6364 (N_6364,N_5983,N_5945);
nor U6365 (N_6365,N_5721,N_5860);
or U6366 (N_6366,N_5830,N_5668);
xnor U6367 (N_6367,N_5595,N_5701);
nand U6368 (N_6368,N_5846,N_5733);
nor U6369 (N_6369,N_5654,N_5928);
and U6370 (N_6370,N_5635,N_5737);
xnor U6371 (N_6371,N_5533,N_5558);
nor U6372 (N_6372,N_5702,N_5854);
and U6373 (N_6373,N_5515,N_5556);
and U6374 (N_6374,N_5672,N_5757);
nor U6375 (N_6375,N_5512,N_5731);
or U6376 (N_6376,N_5968,N_5663);
and U6377 (N_6377,N_5737,N_5894);
and U6378 (N_6378,N_5671,N_5682);
nor U6379 (N_6379,N_5964,N_5755);
or U6380 (N_6380,N_5679,N_5868);
nor U6381 (N_6381,N_5933,N_5831);
nand U6382 (N_6382,N_5818,N_5854);
or U6383 (N_6383,N_5784,N_5739);
and U6384 (N_6384,N_5930,N_5797);
nand U6385 (N_6385,N_5881,N_5500);
and U6386 (N_6386,N_5726,N_5853);
nand U6387 (N_6387,N_5990,N_5650);
nand U6388 (N_6388,N_5787,N_5896);
nand U6389 (N_6389,N_5562,N_5880);
and U6390 (N_6390,N_5855,N_5880);
nor U6391 (N_6391,N_5732,N_5996);
and U6392 (N_6392,N_5701,N_5608);
or U6393 (N_6393,N_5624,N_5970);
nor U6394 (N_6394,N_5743,N_5818);
nand U6395 (N_6395,N_5966,N_5560);
and U6396 (N_6396,N_5684,N_5502);
nor U6397 (N_6397,N_5766,N_5828);
nor U6398 (N_6398,N_5724,N_5781);
nand U6399 (N_6399,N_5832,N_5679);
nor U6400 (N_6400,N_5814,N_5751);
xor U6401 (N_6401,N_5977,N_5824);
nor U6402 (N_6402,N_5765,N_5786);
nand U6403 (N_6403,N_5821,N_5956);
or U6404 (N_6404,N_5860,N_5738);
nor U6405 (N_6405,N_5568,N_5738);
and U6406 (N_6406,N_5639,N_5853);
xor U6407 (N_6407,N_5830,N_5795);
and U6408 (N_6408,N_5777,N_5821);
and U6409 (N_6409,N_5809,N_5707);
or U6410 (N_6410,N_5844,N_5680);
nor U6411 (N_6411,N_5654,N_5509);
or U6412 (N_6412,N_5776,N_5542);
nand U6413 (N_6413,N_5737,N_5684);
or U6414 (N_6414,N_5816,N_5563);
xor U6415 (N_6415,N_5787,N_5728);
or U6416 (N_6416,N_5742,N_5892);
nand U6417 (N_6417,N_5977,N_5607);
or U6418 (N_6418,N_5602,N_5601);
nor U6419 (N_6419,N_5511,N_5800);
or U6420 (N_6420,N_5751,N_5517);
xor U6421 (N_6421,N_5624,N_5507);
nor U6422 (N_6422,N_5543,N_5711);
or U6423 (N_6423,N_5671,N_5756);
and U6424 (N_6424,N_5767,N_5781);
nand U6425 (N_6425,N_5532,N_5713);
nand U6426 (N_6426,N_5813,N_5992);
xnor U6427 (N_6427,N_5703,N_5565);
xor U6428 (N_6428,N_5560,N_5503);
xnor U6429 (N_6429,N_5572,N_5553);
xor U6430 (N_6430,N_5554,N_5880);
or U6431 (N_6431,N_5539,N_5881);
and U6432 (N_6432,N_5669,N_5758);
and U6433 (N_6433,N_5845,N_5640);
xor U6434 (N_6434,N_5940,N_5726);
nor U6435 (N_6435,N_5655,N_5783);
nor U6436 (N_6436,N_5792,N_5848);
nand U6437 (N_6437,N_5736,N_5588);
xnor U6438 (N_6438,N_5906,N_5765);
and U6439 (N_6439,N_5956,N_5689);
xnor U6440 (N_6440,N_5747,N_5585);
xnor U6441 (N_6441,N_5718,N_5880);
or U6442 (N_6442,N_5806,N_5540);
nor U6443 (N_6443,N_5715,N_5909);
and U6444 (N_6444,N_5652,N_5546);
and U6445 (N_6445,N_5889,N_5735);
nor U6446 (N_6446,N_5973,N_5631);
or U6447 (N_6447,N_5549,N_5590);
nand U6448 (N_6448,N_5513,N_5725);
nand U6449 (N_6449,N_5632,N_5511);
xor U6450 (N_6450,N_5770,N_5897);
nand U6451 (N_6451,N_5518,N_5636);
and U6452 (N_6452,N_5624,N_5657);
or U6453 (N_6453,N_5729,N_5556);
and U6454 (N_6454,N_5726,N_5865);
or U6455 (N_6455,N_5938,N_5950);
and U6456 (N_6456,N_5838,N_5798);
nand U6457 (N_6457,N_5817,N_5815);
nor U6458 (N_6458,N_5958,N_5813);
or U6459 (N_6459,N_5625,N_5904);
and U6460 (N_6460,N_5506,N_5876);
and U6461 (N_6461,N_5831,N_5866);
nor U6462 (N_6462,N_5830,N_5613);
nand U6463 (N_6463,N_5578,N_5643);
nor U6464 (N_6464,N_5970,N_5854);
or U6465 (N_6465,N_5709,N_5764);
and U6466 (N_6466,N_5996,N_5984);
xnor U6467 (N_6467,N_5674,N_5705);
nor U6468 (N_6468,N_5611,N_5660);
or U6469 (N_6469,N_5681,N_5960);
or U6470 (N_6470,N_5742,N_5626);
or U6471 (N_6471,N_5742,N_5532);
nand U6472 (N_6472,N_5969,N_5741);
nand U6473 (N_6473,N_5795,N_5714);
nor U6474 (N_6474,N_5512,N_5830);
xnor U6475 (N_6475,N_5682,N_5641);
nand U6476 (N_6476,N_5820,N_5690);
nor U6477 (N_6477,N_5706,N_5753);
xor U6478 (N_6478,N_5500,N_5877);
nand U6479 (N_6479,N_5834,N_5893);
or U6480 (N_6480,N_5761,N_5867);
xnor U6481 (N_6481,N_5553,N_5652);
xor U6482 (N_6482,N_5736,N_5994);
or U6483 (N_6483,N_5640,N_5916);
nor U6484 (N_6484,N_5994,N_5885);
and U6485 (N_6485,N_5771,N_5589);
nand U6486 (N_6486,N_5886,N_5944);
and U6487 (N_6487,N_5506,N_5500);
nor U6488 (N_6488,N_5784,N_5821);
nor U6489 (N_6489,N_5561,N_5761);
nor U6490 (N_6490,N_5921,N_5696);
xor U6491 (N_6491,N_5974,N_5864);
and U6492 (N_6492,N_5557,N_5723);
nor U6493 (N_6493,N_5880,N_5555);
and U6494 (N_6494,N_5973,N_5889);
nand U6495 (N_6495,N_5972,N_5728);
or U6496 (N_6496,N_5618,N_5725);
and U6497 (N_6497,N_5614,N_5646);
xor U6498 (N_6498,N_5937,N_5994);
nand U6499 (N_6499,N_5539,N_5920);
or U6500 (N_6500,N_6158,N_6153);
or U6501 (N_6501,N_6183,N_6152);
and U6502 (N_6502,N_6292,N_6213);
nor U6503 (N_6503,N_6099,N_6453);
xnor U6504 (N_6504,N_6498,N_6046);
xor U6505 (N_6505,N_6067,N_6148);
nand U6506 (N_6506,N_6492,N_6223);
xnor U6507 (N_6507,N_6442,N_6089);
xnor U6508 (N_6508,N_6035,N_6493);
nor U6509 (N_6509,N_6389,N_6130);
or U6510 (N_6510,N_6120,N_6367);
nand U6511 (N_6511,N_6331,N_6311);
and U6512 (N_6512,N_6450,N_6312);
nand U6513 (N_6513,N_6055,N_6346);
xnor U6514 (N_6514,N_6171,N_6326);
and U6515 (N_6515,N_6418,N_6253);
and U6516 (N_6516,N_6234,N_6071);
or U6517 (N_6517,N_6134,N_6110);
xor U6518 (N_6518,N_6485,N_6323);
or U6519 (N_6519,N_6305,N_6200);
nand U6520 (N_6520,N_6195,N_6207);
and U6521 (N_6521,N_6033,N_6194);
xor U6522 (N_6522,N_6411,N_6202);
or U6523 (N_6523,N_6060,N_6366);
or U6524 (N_6524,N_6063,N_6407);
nand U6525 (N_6525,N_6347,N_6256);
and U6526 (N_6526,N_6027,N_6144);
xor U6527 (N_6527,N_6433,N_6447);
nand U6528 (N_6528,N_6233,N_6106);
or U6529 (N_6529,N_6296,N_6357);
nor U6530 (N_6530,N_6294,N_6477);
nand U6531 (N_6531,N_6359,N_6181);
xor U6532 (N_6532,N_6214,N_6472);
nor U6533 (N_6533,N_6039,N_6102);
nand U6534 (N_6534,N_6275,N_6444);
and U6535 (N_6535,N_6496,N_6182);
nor U6536 (N_6536,N_6461,N_6034);
nand U6537 (N_6537,N_6395,N_6222);
nand U6538 (N_6538,N_6340,N_6180);
nand U6539 (N_6539,N_6306,N_6392);
and U6540 (N_6540,N_6459,N_6156);
nand U6541 (N_6541,N_6057,N_6137);
or U6542 (N_6542,N_6211,N_6119);
nand U6543 (N_6543,N_6210,N_6186);
xor U6544 (N_6544,N_6344,N_6164);
and U6545 (N_6545,N_6351,N_6341);
and U6546 (N_6546,N_6072,N_6486);
and U6547 (N_6547,N_6150,N_6307);
nand U6548 (N_6548,N_6416,N_6017);
nor U6549 (N_6549,N_6278,N_6143);
xor U6550 (N_6550,N_6266,N_6385);
nand U6551 (N_6551,N_6022,N_6258);
or U6552 (N_6552,N_6023,N_6086);
and U6553 (N_6553,N_6008,N_6402);
nand U6554 (N_6554,N_6097,N_6135);
xnor U6555 (N_6555,N_6077,N_6238);
or U6556 (N_6556,N_6269,N_6149);
or U6557 (N_6557,N_6235,N_6428);
nor U6558 (N_6558,N_6073,N_6469);
and U6559 (N_6559,N_6398,N_6004);
and U6560 (N_6560,N_6473,N_6084);
nor U6561 (N_6561,N_6456,N_6165);
nor U6562 (N_6562,N_6147,N_6121);
nor U6563 (N_6563,N_6226,N_6010);
nor U6564 (N_6564,N_6413,N_6203);
and U6565 (N_6565,N_6481,N_6045);
or U6566 (N_6566,N_6262,N_6064);
nand U6567 (N_6567,N_6179,N_6076);
xor U6568 (N_6568,N_6257,N_6132);
xor U6569 (N_6569,N_6362,N_6224);
nand U6570 (N_6570,N_6408,N_6217);
or U6571 (N_6571,N_6128,N_6085);
or U6572 (N_6572,N_6437,N_6454);
xor U6573 (N_6573,N_6264,N_6123);
nand U6574 (N_6574,N_6320,N_6052);
or U6575 (N_6575,N_6284,N_6197);
and U6576 (N_6576,N_6490,N_6024);
and U6577 (N_6577,N_6393,N_6404);
nor U6578 (N_6578,N_6126,N_6087);
nor U6579 (N_6579,N_6487,N_6031);
nand U6580 (N_6580,N_6216,N_6310);
xnor U6581 (N_6581,N_6348,N_6322);
nand U6582 (N_6582,N_6409,N_6139);
and U6583 (N_6583,N_6251,N_6370);
nor U6584 (N_6584,N_6184,N_6475);
xnor U6585 (N_6585,N_6178,N_6199);
xor U6586 (N_6586,N_6001,N_6382);
nand U6587 (N_6587,N_6029,N_6040);
or U6588 (N_6588,N_6096,N_6019);
nor U6589 (N_6589,N_6254,N_6208);
or U6590 (N_6590,N_6044,N_6423);
or U6591 (N_6591,N_6100,N_6173);
and U6592 (N_6592,N_6265,N_6098);
or U6593 (N_6593,N_6279,N_6425);
or U6594 (N_6594,N_6479,N_6056);
xor U6595 (N_6595,N_6113,N_6299);
nor U6596 (N_6596,N_6157,N_6336);
xor U6597 (N_6597,N_6452,N_6474);
nand U6598 (N_6598,N_6274,N_6109);
nor U6599 (N_6599,N_6062,N_6049);
nand U6600 (N_6600,N_6020,N_6298);
xnor U6601 (N_6601,N_6397,N_6295);
nand U6602 (N_6602,N_6094,N_6250);
and U6603 (N_6603,N_6261,N_6212);
and U6604 (N_6604,N_6154,N_6354);
xnor U6605 (N_6605,N_6048,N_6009);
and U6606 (N_6606,N_6494,N_6427);
nor U6607 (N_6607,N_6379,N_6104);
nor U6608 (N_6608,N_6438,N_6328);
nor U6609 (N_6609,N_6188,N_6327);
nand U6610 (N_6610,N_6196,N_6365);
xnor U6611 (N_6611,N_6457,N_6315);
and U6612 (N_6612,N_6304,N_6495);
or U6613 (N_6613,N_6483,N_6293);
or U6614 (N_6614,N_6316,N_6421);
nor U6615 (N_6615,N_6018,N_6015);
and U6616 (N_6616,N_6169,N_6297);
xnor U6617 (N_6617,N_6314,N_6036);
nand U6618 (N_6618,N_6191,N_6026);
and U6619 (N_6619,N_6410,N_6353);
and U6620 (N_6620,N_6415,N_6313);
nand U6621 (N_6621,N_6339,N_6422);
xnor U6622 (N_6622,N_6228,N_6381);
xnor U6623 (N_6623,N_6032,N_6175);
xnor U6624 (N_6624,N_6374,N_6361);
or U6625 (N_6625,N_6277,N_6405);
and U6626 (N_6626,N_6300,N_6230);
nand U6627 (N_6627,N_6038,N_6112);
and U6628 (N_6628,N_6050,N_6364);
nor U6629 (N_6629,N_6333,N_6136);
nor U6630 (N_6630,N_6163,N_6133);
xor U6631 (N_6631,N_6319,N_6282);
and U6632 (N_6632,N_6174,N_6412);
xnor U6633 (N_6633,N_6462,N_6061);
nand U6634 (N_6634,N_6105,N_6047);
xor U6635 (N_6635,N_6243,N_6387);
or U6636 (N_6636,N_6125,N_6006);
xor U6637 (N_6637,N_6070,N_6225);
and U6638 (N_6638,N_6499,N_6236);
nor U6639 (N_6639,N_6122,N_6455);
and U6640 (N_6640,N_6114,N_6219);
and U6641 (N_6641,N_6318,N_6273);
nand U6642 (N_6642,N_6394,N_6435);
nand U6643 (N_6643,N_6041,N_6317);
xor U6644 (N_6644,N_6215,N_6115);
nor U6645 (N_6645,N_6237,N_6414);
or U6646 (N_6646,N_6209,N_6103);
or U6647 (N_6647,N_6082,N_6482);
nor U6648 (N_6648,N_6376,N_6360);
xor U6649 (N_6649,N_6054,N_6193);
nand U6650 (N_6650,N_6218,N_6484);
and U6651 (N_6651,N_6424,N_6170);
xnor U6652 (N_6652,N_6124,N_6281);
nand U6653 (N_6653,N_6140,N_6375);
nand U6654 (N_6654,N_6465,N_6160);
xor U6655 (N_6655,N_6380,N_6467);
nand U6656 (N_6656,N_6016,N_6025);
or U6657 (N_6657,N_6276,N_6349);
nor U6658 (N_6658,N_6489,N_6324);
nand U6659 (N_6659,N_6287,N_6204);
nand U6660 (N_6660,N_6338,N_6068);
xnor U6661 (N_6661,N_6259,N_6343);
nand U6662 (N_6662,N_6372,N_6248);
and U6663 (N_6663,N_6384,N_6246);
or U6664 (N_6664,N_6189,N_6345);
or U6665 (N_6665,N_6131,N_6232);
and U6666 (N_6666,N_6014,N_6166);
or U6667 (N_6667,N_6329,N_6302);
nand U6668 (N_6668,N_6332,N_6005);
and U6669 (N_6669,N_6286,N_6268);
xnor U6670 (N_6670,N_6013,N_6363);
or U6671 (N_6671,N_6075,N_6146);
nand U6672 (N_6672,N_6445,N_6288);
nand U6673 (N_6673,N_6478,N_6187);
or U6674 (N_6674,N_6065,N_6242);
nor U6675 (N_6675,N_6468,N_6406);
nor U6676 (N_6676,N_6373,N_6285);
xor U6677 (N_6677,N_6291,N_6419);
or U6678 (N_6678,N_6289,N_6491);
nor U6679 (N_6679,N_6301,N_6162);
or U6680 (N_6680,N_6352,N_6458);
xnor U6681 (N_6681,N_6466,N_6069);
nor U6682 (N_6682,N_6325,N_6240);
nor U6683 (N_6683,N_6101,N_6272);
xor U6684 (N_6684,N_6396,N_6107);
xnor U6685 (N_6685,N_6043,N_6007);
or U6686 (N_6686,N_6434,N_6358);
xnor U6687 (N_6687,N_6066,N_6190);
nor U6688 (N_6688,N_6000,N_6280);
or U6689 (N_6689,N_6172,N_6127);
nor U6690 (N_6690,N_6111,N_6451);
nand U6691 (N_6691,N_6220,N_6206);
xor U6692 (N_6692,N_6037,N_6334);
and U6693 (N_6693,N_6309,N_6141);
nand U6694 (N_6694,N_6449,N_6429);
or U6695 (N_6695,N_6391,N_6058);
nor U6696 (N_6696,N_6471,N_6371);
xor U6697 (N_6697,N_6108,N_6488);
or U6698 (N_6698,N_6463,N_6403);
xnor U6699 (N_6699,N_6470,N_6439);
and U6700 (N_6700,N_6118,N_6177);
nor U6701 (N_6701,N_6308,N_6093);
or U6702 (N_6702,N_6460,N_6337);
and U6703 (N_6703,N_6247,N_6446);
and U6704 (N_6704,N_6003,N_6092);
and U6705 (N_6705,N_6078,N_6021);
nand U6706 (N_6706,N_6377,N_6443);
and U6707 (N_6707,N_6145,N_6263);
nor U6708 (N_6708,N_6388,N_6356);
or U6709 (N_6709,N_6270,N_6267);
xnor U6710 (N_6710,N_6168,N_6192);
or U6711 (N_6711,N_6244,N_6231);
and U6712 (N_6712,N_6355,N_6350);
nor U6713 (N_6713,N_6383,N_6497);
nand U6714 (N_6714,N_6399,N_6378);
or U6715 (N_6715,N_6129,N_6151);
and U6716 (N_6716,N_6426,N_6117);
and U6717 (N_6717,N_6042,N_6249);
nand U6718 (N_6718,N_6142,N_6330);
nor U6719 (N_6719,N_6205,N_6255);
and U6720 (N_6720,N_6053,N_6079);
nor U6721 (N_6721,N_6167,N_6400);
nand U6722 (N_6722,N_6369,N_6271);
nand U6723 (N_6723,N_6431,N_6260);
and U6724 (N_6724,N_6074,N_6030);
nor U6725 (N_6725,N_6051,N_6390);
or U6726 (N_6726,N_6059,N_6011);
and U6727 (N_6727,N_6221,N_6229);
and U6728 (N_6728,N_6012,N_6028);
or U6729 (N_6729,N_6401,N_6081);
or U6730 (N_6730,N_6335,N_6002);
xor U6731 (N_6731,N_6176,N_6303);
nand U6732 (N_6732,N_6417,N_6283);
and U6733 (N_6733,N_6436,N_6116);
or U6734 (N_6734,N_6159,N_6091);
nor U6735 (N_6735,N_6083,N_6185);
nor U6736 (N_6736,N_6441,N_6321);
xnor U6737 (N_6737,N_6252,N_6245);
nor U6738 (N_6738,N_6155,N_6480);
nor U6739 (N_6739,N_6090,N_6368);
xor U6740 (N_6740,N_6080,N_6239);
and U6741 (N_6741,N_6420,N_6448);
or U6742 (N_6742,N_6095,N_6198);
or U6743 (N_6743,N_6241,N_6088);
xnor U6744 (N_6744,N_6386,N_6440);
nand U6745 (N_6745,N_6432,N_6201);
or U6746 (N_6746,N_6138,N_6227);
nand U6747 (N_6747,N_6342,N_6161);
nor U6748 (N_6748,N_6464,N_6290);
xnor U6749 (N_6749,N_6430,N_6476);
nand U6750 (N_6750,N_6090,N_6250);
xnor U6751 (N_6751,N_6192,N_6313);
nor U6752 (N_6752,N_6495,N_6102);
and U6753 (N_6753,N_6109,N_6499);
or U6754 (N_6754,N_6446,N_6342);
nor U6755 (N_6755,N_6344,N_6161);
nor U6756 (N_6756,N_6239,N_6163);
or U6757 (N_6757,N_6158,N_6472);
or U6758 (N_6758,N_6192,N_6288);
nor U6759 (N_6759,N_6099,N_6114);
nand U6760 (N_6760,N_6141,N_6214);
nand U6761 (N_6761,N_6267,N_6198);
nand U6762 (N_6762,N_6004,N_6240);
or U6763 (N_6763,N_6478,N_6458);
nand U6764 (N_6764,N_6077,N_6271);
or U6765 (N_6765,N_6196,N_6476);
and U6766 (N_6766,N_6193,N_6166);
or U6767 (N_6767,N_6362,N_6227);
xnor U6768 (N_6768,N_6218,N_6248);
xor U6769 (N_6769,N_6396,N_6254);
and U6770 (N_6770,N_6240,N_6473);
and U6771 (N_6771,N_6120,N_6443);
and U6772 (N_6772,N_6492,N_6165);
xnor U6773 (N_6773,N_6208,N_6213);
xnor U6774 (N_6774,N_6491,N_6070);
nand U6775 (N_6775,N_6099,N_6115);
nor U6776 (N_6776,N_6447,N_6371);
nand U6777 (N_6777,N_6438,N_6392);
or U6778 (N_6778,N_6090,N_6032);
nor U6779 (N_6779,N_6140,N_6251);
or U6780 (N_6780,N_6225,N_6006);
or U6781 (N_6781,N_6409,N_6193);
nand U6782 (N_6782,N_6137,N_6251);
or U6783 (N_6783,N_6118,N_6193);
nand U6784 (N_6784,N_6216,N_6146);
or U6785 (N_6785,N_6026,N_6259);
and U6786 (N_6786,N_6268,N_6377);
nand U6787 (N_6787,N_6392,N_6096);
and U6788 (N_6788,N_6117,N_6030);
nand U6789 (N_6789,N_6091,N_6118);
xnor U6790 (N_6790,N_6108,N_6250);
xor U6791 (N_6791,N_6225,N_6257);
nand U6792 (N_6792,N_6162,N_6307);
xor U6793 (N_6793,N_6434,N_6368);
xnor U6794 (N_6794,N_6309,N_6020);
or U6795 (N_6795,N_6470,N_6427);
and U6796 (N_6796,N_6305,N_6431);
xor U6797 (N_6797,N_6244,N_6143);
xnor U6798 (N_6798,N_6053,N_6319);
nor U6799 (N_6799,N_6465,N_6377);
nand U6800 (N_6800,N_6126,N_6033);
or U6801 (N_6801,N_6447,N_6390);
nor U6802 (N_6802,N_6088,N_6422);
xor U6803 (N_6803,N_6095,N_6422);
or U6804 (N_6804,N_6218,N_6427);
nor U6805 (N_6805,N_6155,N_6065);
nor U6806 (N_6806,N_6312,N_6139);
xnor U6807 (N_6807,N_6217,N_6330);
xnor U6808 (N_6808,N_6281,N_6056);
nand U6809 (N_6809,N_6145,N_6464);
xnor U6810 (N_6810,N_6157,N_6475);
or U6811 (N_6811,N_6195,N_6369);
nand U6812 (N_6812,N_6059,N_6143);
and U6813 (N_6813,N_6139,N_6070);
nor U6814 (N_6814,N_6364,N_6416);
and U6815 (N_6815,N_6319,N_6189);
or U6816 (N_6816,N_6224,N_6398);
nor U6817 (N_6817,N_6033,N_6260);
nand U6818 (N_6818,N_6326,N_6228);
xnor U6819 (N_6819,N_6172,N_6087);
or U6820 (N_6820,N_6230,N_6492);
and U6821 (N_6821,N_6444,N_6216);
and U6822 (N_6822,N_6176,N_6197);
nand U6823 (N_6823,N_6060,N_6246);
nand U6824 (N_6824,N_6326,N_6066);
xor U6825 (N_6825,N_6289,N_6411);
and U6826 (N_6826,N_6482,N_6216);
xor U6827 (N_6827,N_6380,N_6426);
and U6828 (N_6828,N_6490,N_6065);
or U6829 (N_6829,N_6087,N_6170);
xnor U6830 (N_6830,N_6152,N_6456);
xor U6831 (N_6831,N_6392,N_6092);
and U6832 (N_6832,N_6102,N_6310);
nor U6833 (N_6833,N_6026,N_6459);
or U6834 (N_6834,N_6370,N_6450);
nor U6835 (N_6835,N_6202,N_6429);
xnor U6836 (N_6836,N_6256,N_6087);
or U6837 (N_6837,N_6484,N_6285);
nand U6838 (N_6838,N_6257,N_6484);
nand U6839 (N_6839,N_6238,N_6010);
nand U6840 (N_6840,N_6241,N_6069);
or U6841 (N_6841,N_6459,N_6251);
and U6842 (N_6842,N_6260,N_6355);
nor U6843 (N_6843,N_6234,N_6440);
nand U6844 (N_6844,N_6264,N_6204);
and U6845 (N_6845,N_6346,N_6112);
nand U6846 (N_6846,N_6107,N_6033);
nor U6847 (N_6847,N_6377,N_6365);
or U6848 (N_6848,N_6373,N_6283);
nand U6849 (N_6849,N_6344,N_6441);
and U6850 (N_6850,N_6219,N_6279);
nor U6851 (N_6851,N_6324,N_6014);
and U6852 (N_6852,N_6173,N_6019);
nand U6853 (N_6853,N_6274,N_6090);
or U6854 (N_6854,N_6480,N_6328);
or U6855 (N_6855,N_6165,N_6080);
or U6856 (N_6856,N_6320,N_6332);
xor U6857 (N_6857,N_6269,N_6264);
or U6858 (N_6858,N_6484,N_6215);
or U6859 (N_6859,N_6032,N_6478);
or U6860 (N_6860,N_6228,N_6255);
or U6861 (N_6861,N_6090,N_6272);
or U6862 (N_6862,N_6375,N_6175);
or U6863 (N_6863,N_6301,N_6025);
or U6864 (N_6864,N_6191,N_6004);
and U6865 (N_6865,N_6380,N_6156);
or U6866 (N_6866,N_6053,N_6155);
and U6867 (N_6867,N_6237,N_6262);
nand U6868 (N_6868,N_6397,N_6334);
and U6869 (N_6869,N_6242,N_6186);
nor U6870 (N_6870,N_6314,N_6247);
or U6871 (N_6871,N_6169,N_6394);
nor U6872 (N_6872,N_6328,N_6253);
and U6873 (N_6873,N_6184,N_6214);
nor U6874 (N_6874,N_6282,N_6499);
nor U6875 (N_6875,N_6064,N_6056);
or U6876 (N_6876,N_6193,N_6242);
and U6877 (N_6877,N_6356,N_6335);
xnor U6878 (N_6878,N_6237,N_6065);
nand U6879 (N_6879,N_6253,N_6151);
nand U6880 (N_6880,N_6355,N_6136);
or U6881 (N_6881,N_6239,N_6418);
or U6882 (N_6882,N_6019,N_6295);
xor U6883 (N_6883,N_6092,N_6245);
or U6884 (N_6884,N_6113,N_6423);
nor U6885 (N_6885,N_6478,N_6274);
nor U6886 (N_6886,N_6354,N_6326);
or U6887 (N_6887,N_6128,N_6206);
or U6888 (N_6888,N_6006,N_6298);
and U6889 (N_6889,N_6038,N_6150);
nand U6890 (N_6890,N_6216,N_6335);
xor U6891 (N_6891,N_6025,N_6425);
or U6892 (N_6892,N_6342,N_6469);
xnor U6893 (N_6893,N_6488,N_6207);
xnor U6894 (N_6894,N_6054,N_6038);
xor U6895 (N_6895,N_6023,N_6172);
nand U6896 (N_6896,N_6312,N_6145);
nand U6897 (N_6897,N_6430,N_6049);
nand U6898 (N_6898,N_6026,N_6272);
or U6899 (N_6899,N_6358,N_6184);
or U6900 (N_6900,N_6374,N_6311);
or U6901 (N_6901,N_6123,N_6112);
nand U6902 (N_6902,N_6291,N_6184);
or U6903 (N_6903,N_6151,N_6220);
nor U6904 (N_6904,N_6417,N_6372);
xnor U6905 (N_6905,N_6269,N_6441);
or U6906 (N_6906,N_6045,N_6444);
xnor U6907 (N_6907,N_6253,N_6142);
nand U6908 (N_6908,N_6396,N_6468);
nor U6909 (N_6909,N_6054,N_6255);
or U6910 (N_6910,N_6135,N_6278);
nor U6911 (N_6911,N_6315,N_6041);
xor U6912 (N_6912,N_6115,N_6380);
nand U6913 (N_6913,N_6261,N_6295);
or U6914 (N_6914,N_6389,N_6036);
xor U6915 (N_6915,N_6158,N_6086);
or U6916 (N_6916,N_6181,N_6328);
and U6917 (N_6917,N_6200,N_6454);
nor U6918 (N_6918,N_6320,N_6245);
nand U6919 (N_6919,N_6457,N_6114);
nand U6920 (N_6920,N_6479,N_6219);
nor U6921 (N_6921,N_6390,N_6346);
nor U6922 (N_6922,N_6400,N_6030);
or U6923 (N_6923,N_6210,N_6117);
xnor U6924 (N_6924,N_6124,N_6358);
nor U6925 (N_6925,N_6051,N_6098);
and U6926 (N_6926,N_6308,N_6094);
nand U6927 (N_6927,N_6058,N_6494);
nor U6928 (N_6928,N_6390,N_6247);
nand U6929 (N_6929,N_6119,N_6192);
nand U6930 (N_6930,N_6451,N_6217);
nor U6931 (N_6931,N_6370,N_6077);
nor U6932 (N_6932,N_6439,N_6227);
and U6933 (N_6933,N_6171,N_6269);
xnor U6934 (N_6934,N_6119,N_6357);
nand U6935 (N_6935,N_6189,N_6378);
or U6936 (N_6936,N_6032,N_6357);
or U6937 (N_6937,N_6234,N_6172);
nor U6938 (N_6938,N_6262,N_6452);
nand U6939 (N_6939,N_6119,N_6436);
nand U6940 (N_6940,N_6162,N_6093);
xor U6941 (N_6941,N_6407,N_6469);
nand U6942 (N_6942,N_6286,N_6321);
or U6943 (N_6943,N_6043,N_6054);
nor U6944 (N_6944,N_6443,N_6337);
xnor U6945 (N_6945,N_6138,N_6460);
nor U6946 (N_6946,N_6424,N_6014);
nor U6947 (N_6947,N_6498,N_6174);
and U6948 (N_6948,N_6398,N_6015);
nor U6949 (N_6949,N_6297,N_6254);
or U6950 (N_6950,N_6149,N_6338);
nand U6951 (N_6951,N_6069,N_6289);
or U6952 (N_6952,N_6463,N_6158);
or U6953 (N_6953,N_6479,N_6326);
nand U6954 (N_6954,N_6404,N_6304);
and U6955 (N_6955,N_6079,N_6398);
or U6956 (N_6956,N_6045,N_6147);
and U6957 (N_6957,N_6454,N_6013);
xor U6958 (N_6958,N_6401,N_6122);
xor U6959 (N_6959,N_6316,N_6130);
nand U6960 (N_6960,N_6317,N_6303);
or U6961 (N_6961,N_6360,N_6089);
or U6962 (N_6962,N_6205,N_6200);
or U6963 (N_6963,N_6268,N_6129);
xor U6964 (N_6964,N_6047,N_6104);
xor U6965 (N_6965,N_6490,N_6423);
nor U6966 (N_6966,N_6478,N_6073);
nand U6967 (N_6967,N_6393,N_6251);
xnor U6968 (N_6968,N_6340,N_6241);
nand U6969 (N_6969,N_6393,N_6220);
or U6970 (N_6970,N_6354,N_6390);
and U6971 (N_6971,N_6137,N_6052);
xnor U6972 (N_6972,N_6372,N_6190);
xor U6973 (N_6973,N_6414,N_6231);
or U6974 (N_6974,N_6240,N_6267);
and U6975 (N_6975,N_6422,N_6011);
xor U6976 (N_6976,N_6091,N_6198);
nor U6977 (N_6977,N_6104,N_6292);
or U6978 (N_6978,N_6472,N_6335);
nand U6979 (N_6979,N_6385,N_6312);
nor U6980 (N_6980,N_6298,N_6281);
xor U6981 (N_6981,N_6455,N_6318);
xnor U6982 (N_6982,N_6047,N_6143);
nand U6983 (N_6983,N_6337,N_6004);
nand U6984 (N_6984,N_6424,N_6088);
and U6985 (N_6985,N_6019,N_6471);
nand U6986 (N_6986,N_6133,N_6146);
xnor U6987 (N_6987,N_6494,N_6330);
and U6988 (N_6988,N_6075,N_6032);
xor U6989 (N_6989,N_6230,N_6088);
nand U6990 (N_6990,N_6432,N_6453);
xnor U6991 (N_6991,N_6236,N_6426);
xnor U6992 (N_6992,N_6272,N_6054);
and U6993 (N_6993,N_6444,N_6239);
and U6994 (N_6994,N_6265,N_6094);
nand U6995 (N_6995,N_6417,N_6162);
nor U6996 (N_6996,N_6253,N_6090);
nor U6997 (N_6997,N_6432,N_6265);
nand U6998 (N_6998,N_6063,N_6440);
or U6999 (N_6999,N_6275,N_6042);
and U7000 (N_7000,N_6652,N_6745);
or U7001 (N_7001,N_6597,N_6547);
and U7002 (N_7002,N_6509,N_6873);
and U7003 (N_7003,N_6684,N_6777);
xnor U7004 (N_7004,N_6616,N_6897);
and U7005 (N_7005,N_6676,N_6655);
nand U7006 (N_7006,N_6571,N_6693);
nor U7007 (N_7007,N_6635,N_6596);
xnor U7008 (N_7008,N_6633,N_6771);
nor U7009 (N_7009,N_6669,N_6586);
xor U7010 (N_7010,N_6766,N_6550);
and U7011 (N_7011,N_6713,N_6931);
xnor U7012 (N_7012,N_6627,N_6945);
or U7013 (N_7013,N_6634,N_6820);
or U7014 (N_7014,N_6724,N_6532);
nand U7015 (N_7015,N_6716,N_6804);
nor U7016 (N_7016,N_6651,N_6666);
xor U7017 (N_7017,N_6695,N_6670);
and U7018 (N_7018,N_6915,N_6859);
nor U7019 (N_7019,N_6902,N_6846);
nor U7020 (N_7020,N_6889,N_6769);
xnor U7021 (N_7021,N_6842,N_6872);
nor U7022 (N_7022,N_6883,N_6743);
and U7023 (N_7023,N_6639,N_6973);
nor U7024 (N_7024,N_6779,N_6994);
and U7025 (N_7025,N_6988,N_6910);
and U7026 (N_7026,N_6563,N_6912);
nand U7027 (N_7027,N_6914,N_6824);
nor U7028 (N_7028,N_6870,N_6643);
xnor U7029 (N_7029,N_6538,N_6558);
xor U7030 (N_7030,N_6932,N_6511);
nor U7031 (N_7031,N_6933,N_6927);
nand U7032 (N_7032,N_6867,N_6857);
or U7033 (N_7033,N_6710,N_6986);
and U7034 (N_7034,N_6928,N_6683);
nor U7035 (N_7035,N_6949,N_6637);
nor U7036 (N_7036,N_6853,N_6561);
and U7037 (N_7037,N_6908,N_6685);
nor U7038 (N_7038,N_6767,N_6874);
xnor U7039 (N_7039,N_6696,N_6956);
or U7040 (N_7040,N_6798,N_6725);
and U7041 (N_7041,N_6658,N_6972);
or U7042 (N_7042,N_6821,N_6880);
and U7043 (N_7043,N_6899,N_6649);
nand U7044 (N_7044,N_6922,N_6833);
nand U7045 (N_7045,N_6791,N_6521);
nor U7046 (N_7046,N_6794,N_6930);
xnor U7047 (N_7047,N_6541,N_6885);
and U7048 (N_7048,N_6925,N_6587);
or U7049 (N_7049,N_6730,N_6506);
xnor U7050 (N_7050,N_6985,N_6705);
xnor U7051 (N_7051,N_6628,N_6584);
nand U7052 (N_7052,N_6917,N_6524);
or U7053 (N_7053,N_6989,N_6665);
nand U7054 (N_7054,N_6540,N_6965);
or U7055 (N_7055,N_6592,N_6756);
xor U7056 (N_7056,N_6687,N_6508);
or U7057 (N_7057,N_6784,N_6507);
nand U7058 (N_7058,N_6613,N_6739);
xnor U7059 (N_7059,N_6717,N_6752);
xnor U7060 (N_7060,N_6572,N_6722);
xnor U7061 (N_7061,N_6523,N_6653);
or U7062 (N_7062,N_6667,N_6823);
xnor U7063 (N_7063,N_6625,N_6975);
nand U7064 (N_7064,N_6736,N_6799);
nor U7065 (N_7065,N_6602,N_6951);
nand U7066 (N_7066,N_6900,N_6935);
xor U7067 (N_7067,N_6882,N_6701);
nor U7068 (N_7068,N_6734,N_6677);
and U7069 (N_7069,N_6887,N_6732);
and U7070 (N_7070,N_6761,N_6786);
nand U7071 (N_7071,N_6689,N_6575);
or U7072 (N_7072,N_6668,N_6517);
and U7073 (N_7073,N_6773,N_6817);
and U7074 (N_7074,N_6615,N_6694);
nand U7075 (N_7075,N_6618,N_6849);
nand U7076 (N_7076,N_6591,N_6603);
xnor U7077 (N_7077,N_6714,N_6648);
nand U7078 (N_7078,N_6795,N_6848);
nor U7079 (N_7079,N_6623,N_6569);
nand U7080 (N_7080,N_6647,N_6692);
nand U7081 (N_7081,N_6827,N_6865);
or U7082 (N_7082,N_6715,N_6758);
nor U7083 (N_7083,N_6774,N_6789);
or U7084 (N_7084,N_6838,N_6557);
or U7085 (N_7085,N_6898,N_6860);
or U7086 (N_7086,N_6936,N_6918);
xnor U7087 (N_7087,N_6564,N_6967);
or U7088 (N_7088,N_6548,N_6620);
or U7089 (N_7089,N_6680,N_6772);
or U7090 (N_7090,N_6529,N_6905);
nand U7091 (N_7091,N_6686,N_6500);
or U7092 (N_7092,N_6578,N_6585);
or U7093 (N_7093,N_6921,N_6530);
or U7094 (N_7094,N_6744,N_6733);
or U7095 (N_7095,N_6505,N_6886);
xnor U7096 (N_7096,N_6929,N_6958);
nand U7097 (N_7097,N_6545,N_6626);
or U7098 (N_7098,N_6796,N_6818);
nand U7099 (N_7099,N_6963,N_6681);
xnor U7100 (N_7100,N_6978,N_6518);
nor U7101 (N_7101,N_6600,N_6519);
or U7102 (N_7102,N_6711,N_6810);
nor U7103 (N_7103,N_6590,N_6565);
nand U7104 (N_7104,N_6504,N_6837);
nand U7105 (N_7105,N_6974,N_6803);
xor U7106 (N_7106,N_6982,N_6559);
or U7107 (N_7107,N_6993,N_6619);
nor U7108 (N_7108,N_6863,N_6574);
nand U7109 (N_7109,N_6924,N_6934);
xor U7110 (N_7110,N_6757,N_6845);
nand U7111 (N_7111,N_6811,N_6806);
or U7112 (N_7112,N_6990,N_6727);
nand U7113 (N_7113,N_6778,N_6913);
and U7114 (N_7114,N_6536,N_6866);
nand U7115 (N_7115,N_6690,N_6721);
or U7116 (N_7116,N_6879,N_6871);
nand U7117 (N_7117,N_6851,N_6642);
nand U7118 (N_7118,N_6904,N_6788);
xnor U7119 (N_7119,N_6555,N_6709);
and U7120 (N_7120,N_6875,N_6916);
nand U7121 (N_7121,N_6992,N_6790);
nor U7122 (N_7122,N_6737,N_6957);
xnor U7123 (N_7123,N_6944,N_6976);
xor U7124 (N_7124,N_6723,N_6601);
and U7125 (N_7125,N_6691,N_6549);
nand U7126 (N_7126,N_6868,N_6567);
xor U7127 (N_7127,N_6780,N_6661);
nor U7128 (N_7128,N_6775,N_6969);
nand U7129 (N_7129,N_6970,N_6759);
xor U7130 (N_7130,N_6594,N_6862);
and U7131 (N_7131,N_6726,N_6527);
or U7132 (N_7132,N_6729,N_6828);
or U7133 (N_7133,N_6593,N_6891);
xor U7134 (N_7134,N_6749,N_6844);
or U7135 (N_7135,N_6942,N_6983);
xor U7136 (N_7136,N_6996,N_6835);
nand U7137 (N_7137,N_6675,N_6840);
nand U7138 (N_7138,N_6706,N_6740);
or U7139 (N_7139,N_6528,N_6770);
and U7140 (N_7140,N_6582,N_6566);
nor U7141 (N_7141,N_6588,N_6673);
xor U7142 (N_7142,N_6702,N_6955);
or U7143 (N_7143,N_6819,N_6869);
nand U7144 (N_7144,N_6698,N_6577);
xnor U7145 (N_7145,N_6608,N_6920);
nor U7146 (N_7146,N_6854,N_6632);
nor U7147 (N_7147,N_6662,N_6700);
nand U7148 (N_7148,N_6834,N_6896);
xor U7149 (N_7149,N_6741,N_6570);
nor U7150 (N_7150,N_6510,N_6946);
xor U7151 (N_7151,N_6544,N_6881);
and U7152 (N_7152,N_6947,N_6793);
nor U7153 (N_7153,N_6631,N_6814);
xor U7154 (N_7154,N_6843,N_6551);
nor U7155 (N_7155,N_6878,N_6977);
nand U7156 (N_7156,N_6901,N_6589);
nor U7157 (N_7157,N_6813,N_6964);
or U7158 (N_7158,N_6979,N_6808);
nand U7159 (N_7159,N_6830,N_6501);
and U7160 (N_7160,N_6512,N_6611);
xor U7161 (N_7161,N_6783,N_6839);
nand U7162 (N_7162,N_6847,N_6877);
xnor U7163 (N_7163,N_6797,N_6852);
xor U7164 (N_7164,N_6580,N_6535);
nor U7165 (N_7165,N_6579,N_6952);
xor U7166 (N_7166,N_6809,N_6903);
and U7167 (N_7167,N_6624,N_6938);
xnor U7168 (N_7168,N_6629,N_6640);
and U7169 (N_7169,N_6776,N_6768);
nand U7170 (N_7170,N_6966,N_6531);
xnor U7171 (N_7171,N_6815,N_6525);
nand U7172 (N_7172,N_6858,N_6672);
or U7173 (N_7173,N_6971,N_6950);
xor U7174 (N_7174,N_6699,N_6503);
and U7175 (N_7175,N_6607,N_6650);
and U7176 (N_7176,N_6678,N_6754);
or U7177 (N_7177,N_6622,N_6641);
and U7178 (N_7178,N_6841,N_6760);
and U7179 (N_7179,N_6812,N_6763);
xor U7180 (N_7180,N_6805,N_6553);
or U7181 (N_7181,N_6907,N_6537);
nor U7182 (N_7182,N_6671,N_6543);
and U7183 (N_7183,N_6679,N_6660);
xor U7184 (N_7184,N_6638,N_6836);
and U7185 (N_7185,N_6961,N_6906);
or U7186 (N_7186,N_6998,N_6831);
nor U7187 (N_7187,N_6522,N_6636);
nor U7188 (N_7188,N_6984,N_6703);
nand U7189 (N_7189,N_6939,N_6573);
nor U7190 (N_7190,N_6822,N_6539);
nand U7191 (N_7191,N_6612,N_6892);
nor U7192 (N_7192,N_6552,N_6514);
nand U7193 (N_7193,N_6765,N_6782);
xor U7194 (N_7194,N_6610,N_6542);
nor U7195 (N_7195,N_6962,N_6911);
or U7196 (N_7196,N_6785,N_6595);
and U7197 (N_7197,N_6832,N_6747);
and U7198 (N_7198,N_6981,N_6598);
or U7199 (N_7199,N_6850,N_6750);
nor U7200 (N_7200,N_6720,N_6630);
nand U7201 (N_7201,N_6893,N_6856);
and U7202 (N_7202,N_6787,N_6513);
nand U7203 (N_7203,N_6968,N_6583);
and U7204 (N_7204,N_6940,N_6712);
or U7205 (N_7205,N_6581,N_6718);
nor U7206 (N_7206,N_6864,N_6534);
or U7207 (N_7207,N_6959,N_6943);
or U7208 (N_7208,N_6825,N_6707);
and U7209 (N_7209,N_6895,N_6576);
xor U7210 (N_7210,N_6645,N_6919);
and U7211 (N_7211,N_6688,N_6755);
xor U7212 (N_7212,N_6909,N_6807);
and U7213 (N_7213,N_6560,N_6654);
and U7214 (N_7214,N_6997,N_6515);
and U7215 (N_7215,N_6704,N_6753);
nand U7216 (N_7216,N_6748,N_6991);
nor U7217 (N_7217,N_6533,N_6738);
and U7218 (N_7218,N_6708,N_6656);
or U7219 (N_7219,N_6599,N_6604);
nor U7220 (N_7220,N_6742,N_6953);
xor U7221 (N_7221,N_6960,N_6876);
and U7222 (N_7222,N_6617,N_6802);
and U7223 (N_7223,N_6888,N_6697);
and U7224 (N_7224,N_6516,N_6948);
or U7225 (N_7225,N_6657,N_6562);
and U7226 (N_7226,N_6751,N_6800);
xor U7227 (N_7227,N_6664,N_6999);
or U7228 (N_7228,N_6568,N_6926);
or U7229 (N_7229,N_6923,N_6526);
or U7230 (N_7230,N_6605,N_6735);
xor U7231 (N_7231,N_6556,N_6987);
nand U7232 (N_7232,N_6674,N_6663);
and U7233 (N_7233,N_6609,N_6621);
xnor U7234 (N_7234,N_6861,N_6980);
xnor U7235 (N_7235,N_6659,N_6646);
nor U7236 (N_7236,N_6719,N_6995);
xor U7237 (N_7237,N_6731,N_6781);
xor U7238 (N_7238,N_6614,N_6554);
and U7239 (N_7239,N_6829,N_6746);
nor U7240 (N_7240,N_6890,N_6682);
and U7241 (N_7241,N_6937,N_6728);
nor U7242 (N_7242,N_6855,N_6826);
nand U7243 (N_7243,N_6894,N_6884);
nand U7244 (N_7244,N_6954,N_6801);
or U7245 (N_7245,N_6764,N_6941);
nand U7246 (N_7246,N_6792,N_6762);
nor U7247 (N_7247,N_6520,N_6546);
or U7248 (N_7248,N_6606,N_6644);
nor U7249 (N_7249,N_6502,N_6816);
nand U7250 (N_7250,N_6905,N_6980);
nand U7251 (N_7251,N_6885,N_6884);
nand U7252 (N_7252,N_6875,N_6862);
nand U7253 (N_7253,N_6810,N_6958);
nor U7254 (N_7254,N_6857,N_6789);
and U7255 (N_7255,N_6852,N_6677);
or U7256 (N_7256,N_6544,N_6593);
xor U7257 (N_7257,N_6557,N_6643);
nor U7258 (N_7258,N_6592,N_6816);
nor U7259 (N_7259,N_6737,N_6749);
nand U7260 (N_7260,N_6512,N_6613);
nor U7261 (N_7261,N_6550,N_6540);
xnor U7262 (N_7262,N_6639,N_6516);
and U7263 (N_7263,N_6599,N_6779);
xor U7264 (N_7264,N_6680,N_6551);
nand U7265 (N_7265,N_6953,N_6652);
nor U7266 (N_7266,N_6712,N_6559);
nor U7267 (N_7267,N_6974,N_6734);
nor U7268 (N_7268,N_6618,N_6576);
or U7269 (N_7269,N_6662,N_6785);
or U7270 (N_7270,N_6614,N_6621);
and U7271 (N_7271,N_6888,N_6757);
nand U7272 (N_7272,N_6950,N_6998);
nor U7273 (N_7273,N_6507,N_6509);
nor U7274 (N_7274,N_6907,N_6731);
xor U7275 (N_7275,N_6680,N_6741);
or U7276 (N_7276,N_6638,N_6769);
nor U7277 (N_7277,N_6522,N_6756);
xor U7278 (N_7278,N_6909,N_6790);
and U7279 (N_7279,N_6853,N_6733);
nand U7280 (N_7280,N_6955,N_6758);
nor U7281 (N_7281,N_6502,N_6615);
and U7282 (N_7282,N_6650,N_6507);
nor U7283 (N_7283,N_6731,N_6583);
nor U7284 (N_7284,N_6829,N_6589);
nand U7285 (N_7285,N_6956,N_6753);
and U7286 (N_7286,N_6825,N_6505);
or U7287 (N_7287,N_6617,N_6604);
or U7288 (N_7288,N_6534,N_6874);
nor U7289 (N_7289,N_6841,N_6717);
nor U7290 (N_7290,N_6608,N_6765);
nor U7291 (N_7291,N_6999,N_6814);
nor U7292 (N_7292,N_6773,N_6655);
nor U7293 (N_7293,N_6815,N_6857);
nor U7294 (N_7294,N_6790,N_6530);
xnor U7295 (N_7295,N_6735,N_6625);
nand U7296 (N_7296,N_6762,N_6528);
or U7297 (N_7297,N_6720,N_6811);
nor U7298 (N_7298,N_6500,N_6870);
nand U7299 (N_7299,N_6774,N_6721);
and U7300 (N_7300,N_6694,N_6536);
nor U7301 (N_7301,N_6553,N_6695);
and U7302 (N_7302,N_6646,N_6817);
nor U7303 (N_7303,N_6712,N_6605);
xnor U7304 (N_7304,N_6661,N_6880);
nand U7305 (N_7305,N_6713,N_6803);
nand U7306 (N_7306,N_6976,N_6700);
or U7307 (N_7307,N_6513,N_6529);
nor U7308 (N_7308,N_6701,N_6847);
or U7309 (N_7309,N_6802,N_6615);
xor U7310 (N_7310,N_6503,N_6701);
and U7311 (N_7311,N_6617,N_6878);
and U7312 (N_7312,N_6505,N_6755);
xor U7313 (N_7313,N_6705,N_6581);
or U7314 (N_7314,N_6659,N_6996);
or U7315 (N_7315,N_6986,N_6658);
nand U7316 (N_7316,N_6959,N_6830);
xor U7317 (N_7317,N_6789,N_6731);
and U7318 (N_7318,N_6794,N_6641);
nor U7319 (N_7319,N_6856,N_6811);
and U7320 (N_7320,N_6539,N_6983);
nor U7321 (N_7321,N_6648,N_6878);
or U7322 (N_7322,N_6808,N_6619);
and U7323 (N_7323,N_6856,N_6616);
nor U7324 (N_7324,N_6933,N_6939);
nand U7325 (N_7325,N_6591,N_6509);
nand U7326 (N_7326,N_6716,N_6641);
and U7327 (N_7327,N_6908,N_6586);
nand U7328 (N_7328,N_6975,N_6927);
or U7329 (N_7329,N_6505,N_6939);
xnor U7330 (N_7330,N_6777,N_6550);
nand U7331 (N_7331,N_6672,N_6726);
nand U7332 (N_7332,N_6905,N_6970);
and U7333 (N_7333,N_6885,N_6825);
xor U7334 (N_7334,N_6613,N_6788);
xor U7335 (N_7335,N_6936,N_6959);
or U7336 (N_7336,N_6866,N_6540);
xor U7337 (N_7337,N_6894,N_6518);
nand U7338 (N_7338,N_6520,N_6648);
or U7339 (N_7339,N_6803,N_6929);
and U7340 (N_7340,N_6618,N_6822);
and U7341 (N_7341,N_6734,N_6815);
or U7342 (N_7342,N_6723,N_6991);
nand U7343 (N_7343,N_6530,N_6751);
xnor U7344 (N_7344,N_6592,N_6722);
and U7345 (N_7345,N_6694,N_6692);
xor U7346 (N_7346,N_6721,N_6757);
xor U7347 (N_7347,N_6636,N_6994);
and U7348 (N_7348,N_6999,N_6712);
nor U7349 (N_7349,N_6888,N_6501);
xor U7350 (N_7350,N_6752,N_6919);
or U7351 (N_7351,N_6797,N_6551);
xor U7352 (N_7352,N_6618,N_6579);
nor U7353 (N_7353,N_6933,N_6545);
or U7354 (N_7354,N_6606,N_6746);
and U7355 (N_7355,N_6724,N_6951);
nor U7356 (N_7356,N_6732,N_6685);
and U7357 (N_7357,N_6853,N_6959);
xor U7358 (N_7358,N_6965,N_6565);
xnor U7359 (N_7359,N_6509,N_6922);
xor U7360 (N_7360,N_6823,N_6971);
nor U7361 (N_7361,N_6667,N_6953);
or U7362 (N_7362,N_6570,N_6730);
or U7363 (N_7363,N_6606,N_6514);
and U7364 (N_7364,N_6674,N_6946);
nor U7365 (N_7365,N_6501,N_6657);
nand U7366 (N_7366,N_6770,N_6753);
nand U7367 (N_7367,N_6697,N_6872);
xnor U7368 (N_7368,N_6939,N_6926);
and U7369 (N_7369,N_6899,N_6673);
xor U7370 (N_7370,N_6579,N_6592);
nor U7371 (N_7371,N_6865,N_6602);
and U7372 (N_7372,N_6727,N_6565);
nand U7373 (N_7373,N_6751,N_6890);
and U7374 (N_7374,N_6741,N_6862);
and U7375 (N_7375,N_6525,N_6857);
nand U7376 (N_7376,N_6703,N_6549);
xor U7377 (N_7377,N_6923,N_6632);
or U7378 (N_7378,N_6671,N_6986);
and U7379 (N_7379,N_6920,N_6944);
or U7380 (N_7380,N_6931,N_6786);
or U7381 (N_7381,N_6745,N_6604);
nand U7382 (N_7382,N_6853,N_6724);
or U7383 (N_7383,N_6670,N_6806);
xnor U7384 (N_7384,N_6608,N_6529);
or U7385 (N_7385,N_6662,N_6947);
xnor U7386 (N_7386,N_6523,N_6840);
nand U7387 (N_7387,N_6805,N_6781);
or U7388 (N_7388,N_6672,N_6579);
or U7389 (N_7389,N_6872,N_6631);
or U7390 (N_7390,N_6768,N_6904);
nand U7391 (N_7391,N_6819,N_6840);
xor U7392 (N_7392,N_6593,N_6668);
or U7393 (N_7393,N_6864,N_6902);
nor U7394 (N_7394,N_6716,N_6633);
or U7395 (N_7395,N_6899,N_6730);
xor U7396 (N_7396,N_6530,N_6966);
and U7397 (N_7397,N_6972,N_6758);
or U7398 (N_7398,N_6943,N_6572);
or U7399 (N_7399,N_6820,N_6552);
and U7400 (N_7400,N_6760,N_6537);
or U7401 (N_7401,N_6991,N_6767);
or U7402 (N_7402,N_6860,N_6837);
and U7403 (N_7403,N_6733,N_6933);
or U7404 (N_7404,N_6827,N_6831);
or U7405 (N_7405,N_6589,N_6813);
and U7406 (N_7406,N_6844,N_6955);
or U7407 (N_7407,N_6773,N_6926);
nor U7408 (N_7408,N_6744,N_6687);
and U7409 (N_7409,N_6756,N_6719);
nor U7410 (N_7410,N_6992,N_6591);
and U7411 (N_7411,N_6974,N_6613);
xor U7412 (N_7412,N_6671,N_6746);
nor U7413 (N_7413,N_6976,N_6612);
or U7414 (N_7414,N_6653,N_6587);
and U7415 (N_7415,N_6561,N_6879);
or U7416 (N_7416,N_6663,N_6759);
nor U7417 (N_7417,N_6971,N_6764);
nor U7418 (N_7418,N_6577,N_6645);
nand U7419 (N_7419,N_6535,N_6636);
nand U7420 (N_7420,N_6960,N_6504);
xnor U7421 (N_7421,N_6665,N_6819);
or U7422 (N_7422,N_6547,N_6788);
nand U7423 (N_7423,N_6814,N_6601);
nand U7424 (N_7424,N_6853,N_6591);
nand U7425 (N_7425,N_6747,N_6566);
nand U7426 (N_7426,N_6604,N_6531);
or U7427 (N_7427,N_6739,N_6719);
nand U7428 (N_7428,N_6777,N_6932);
and U7429 (N_7429,N_6684,N_6886);
or U7430 (N_7430,N_6592,N_6726);
nand U7431 (N_7431,N_6906,N_6950);
xor U7432 (N_7432,N_6898,N_6543);
nor U7433 (N_7433,N_6648,N_6825);
nor U7434 (N_7434,N_6805,N_6984);
or U7435 (N_7435,N_6801,N_6735);
nand U7436 (N_7436,N_6733,N_6719);
nor U7437 (N_7437,N_6700,N_6622);
or U7438 (N_7438,N_6794,N_6868);
nand U7439 (N_7439,N_6750,N_6825);
and U7440 (N_7440,N_6873,N_6906);
and U7441 (N_7441,N_6588,N_6531);
nor U7442 (N_7442,N_6506,N_6968);
nor U7443 (N_7443,N_6595,N_6879);
xnor U7444 (N_7444,N_6830,N_6949);
nor U7445 (N_7445,N_6583,N_6885);
xnor U7446 (N_7446,N_6531,N_6704);
nor U7447 (N_7447,N_6560,N_6690);
and U7448 (N_7448,N_6791,N_6688);
and U7449 (N_7449,N_6539,N_6598);
or U7450 (N_7450,N_6691,N_6763);
nand U7451 (N_7451,N_6997,N_6666);
or U7452 (N_7452,N_6751,N_6741);
xor U7453 (N_7453,N_6652,N_6654);
nand U7454 (N_7454,N_6792,N_6906);
nor U7455 (N_7455,N_6742,N_6754);
nand U7456 (N_7456,N_6635,N_6602);
nand U7457 (N_7457,N_6518,N_6797);
nand U7458 (N_7458,N_6799,N_6698);
and U7459 (N_7459,N_6831,N_6870);
nand U7460 (N_7460,N_6801,N_6951);
xnor U7461 (N_7461,N_6581,N_6655);
or U7462 (N_7462,N_6796,N_6812);
nand U7463 (N_7463,N_6739,N_6962);
xor U7464 (N_7464,N_6568,N_6596);
and U7465 (N_7465,N_6673,N_6657);
nor U7466 (N_7466,N_6559,N_6512);
nand U7467 (N_7467,N_6806,N_6910);
nand U7468 (N_7468,N_6786,N_6795);
and U7469 (N_7469,N_6692,N_6758);
and U7470 (N_7470,N_6570,N_6934);
or U7471 (N_7471,N_6841,N_6699);
xnor U7472 (N_7472,N_6877,N_6984);
xnor U7473 (N_7473,N_6876,N_6858);
nand U7474 (N_7474,N_6927,N_6971);
or U7475 (N_7475,N_6621,N_6863);
and U7476 (N_7476,N_6804,N_6736);
nand U7477 (N_7477,N_6627,N_6546);
xnor U7478 (N_7478,N_6889,N_6717);
xor U7479 (N_7479,N_6964,N_6886);
nand U7480 (N_7480,N_6586,N_6859);
or U7481 (N_7481,N_6522,N_6926);
xor U7482 (N_7482,N_6745,N_6686);
and U7483 (N_7483,N_6561,N_6666);
or U7484 (N_7484,N_6582,N_6827);
xor U7485 (N_7485,N_6724,N_6698);
or U7486 (N_7486,N_6557,N_6907);
and U7487 (N_7487,N_6552,N_6635);
or U7488 (N_7488,N_6686,N_6939);
nand U7489 (N_7489,N_6580,N_6608);
or U7490 (N_7490,N_6770,N_6552);
or U7491 (N_7491,N_6601,N_6702);
nor U7492 (N_7492,N_6810,N_6719);
nand U7493 (N_7493,N_6891,N_6984);
or U7494 (N_7494,N_6573,N_6549);
xor U7495 (N_7495,N_6563,N_6543);
or U7496 (N_7496,N_6599,N_6682);
and U7497 (N_7497,N_6669,N_6761);
nor U7498 (N_7498,N_6724,N_6797);
or U7499 (N_7499,N_6729,N_6946);
xnor U7500 (N_7500,N_7458,N_7466);
xnor U7501 (N_7501,N_7419,N_7344);
nor U7502 (N_7502,N_7151,N_7492);
nand U7503 (N_7503,N_7482,N_7444);
xor U7504 (N_7504,N_7379,N_7368);
and U7505 (N_7505,N_7037,N_7446);
nand U7506 (N_7506,N_7480,N_7290);
and U7507 (N_7507,N_7380,N_7157);
nand U7508 (N_7508,N_7386,N_7360);
nand U7509 (N_7509,N_7412,N_7439);
nor U7510 (N_7510,N_7213,N_7226);
xnor U7511 (N_7511,N_7479,N_7276);
nor U7512 (N_7512,N_7023,N_7041);
or U7513 (N_7513,N_7417,N_7388);
nand U7514 (N_7514,N_7264,N_7060);
nand U7515 (N_7515,N_7159,N_7073);
and U7516 (N_7516,N_7189,N_7399);
or U7517 (N_7517,N_7208,N_7232);
and U7518 (N_7518,N_7281,N_7071);
nor U7519 (N_7519,N_7366,N_7053);
or U7520 (N_7520,N_7364,N_7470);
xor U7521 (N_7521,N_7358,N_7147);
or U7522 (N_7522,N_7080,N_7477);
and U7523 (N_7523,N_7097,N_7429);
xnor U7524 (N_7524,N_7187,N_7322);
and U7525 (N_7525,N_7017,N_7178);
nand U7526 (N_7526,N_7355,N_7059);
xor U7527 (N_7527,N_7155,N_7202);
and U7528 (N_7528,N_7445,N_7292);
nand U7529 (N_7529,N_7451,N_7047);
nor U7530 (N_7530,N_7294,N_7449);
nor U7531 (N_7531,N_7204,N_7486);
xnor U7532 (N_7532,N_7141,N_7282);
nand U7533 (N_7533,N_7374,N_7296);
nor U7534 (N_7534,N_7148,N_7117);
xor U7535 (N_7535,N_7179,N_7332);
and U7536 (N_7536,N_7400,N_7257);
nor U7537 (N_7537,N_7267,N_7197);
nor U7538 (N_7538,N_7311,N_7370);
or U7539 (N_7539,N_7464,N_7215);
xor U7540 (N_7540,N_7490,N_7090);
and U7541 (N_7541,N_7127,N_7002);
and U7542 (N_7542,N_7062,N_7418);
xnor U7543 (N_7543,N_7167,N_7277);
and U7544 (N_7544,N_7485,N_7044);
or U7545 (N_7545,N_7089,N_7307);
nand U7546 (N_7546,N_7401,N_7042);
or U7547 (N_7547,N_7103,N_7180);
nand U7548 (N_7548,N_7182,N_7009);
nor U7549 (N_7549,N_7415,N_7468);
and U7550 (N_7550,N_7383,N_7373);
and U7551 (N_7551,N_7420,N_7057);
nor U7552 (N_7552,N_7132,N_7454);
nor U7553 (N_7553,N_7392,N_7312);
xor U7554 (N_7554,N_7483,N_7450);
xor U7555 (N_7555,N_7069,N_7183);
or U7556 (N_7556,N_7195,N_7173);
and U7557 (N_7557,N_7496,N_7046);
nand U7558 (N_7558,N_7299,N_7020);
nand U7559 (N_7559,N_7193,N_7194);
nand U7560 (N_7560,N_7237,N_7301);
nor U7561 (N_7561,N_7138,N_7121);
and U7562 (N_7562,N_7150,N_7135);
or U7563 (N_7563,N_7295,N_7263);
and U7564 (N_7564,N_7251,N_7235);
nor U7565 (N_7565,N_7261,N_7376);
nor U7566 (N_7566,N_7222,N_7385);
xor U7567 (N_7567,N_7199,N_7184);
xor U7568 (N_7568,N_7395,N_7457);
or U7569 (N_7569,N_7109,N_7064);
or U7570 (N_7570,N_7402,N_7221);
nand U7571 (N_7571,N_7153,N_7421);
nor U7572 (N_7572,N_7461,N_7433);
nand U7573 (N_7573,N_7072,N_7349);
and U7574 (N_7574,N_7164,N_7128);
nand U7575 (N_7575,N_7414,N_7129);
nand U7576 (N_7576,N_7315,N_7130);
and U7577 (N_7577,N_7345,N_7122);
or U7578 (N_7578,N_7317,N_7170);
nor U7579 (N_7579,N_7165,N_7493);
or U7580 (N_7580,N_7359,N_7156);
xnor U7581 (N_7581,N_7387,N_7448);
xor U7582 (N_7582,N_7110,N_7453);
xnor U7583 (N_7583,N_7365,N_7049);
nand U7584 (N_7584,N_7298,N_7306);
xor U7585 (N_7585,N_7242,N_7275);
and U7586 (N_7586,N_7131,N_7196);
nand U7587 (N_7587,N_7061,N_7323);
nand U7588 (N_7588,N_7216,N_7015);
nor U7589 (N_7589,N_7025,N_7287);
or U7590 (N_7590,N_7106,N_7269);
or U7591 (N_7591,N_7394,N_7176);
or U7592 (N_7592,N_7120,N_7337);
and U7593 (N_7593,N_7036,N_7363);
nand U7594 (N_7594,N_7190,N_7459);
and U7595 (N_7595,N_7227,N_7123);
nor U7596 (N_7596,N_7030,N_7168);
nand U7597 (N_7597,N_7104,N_7174);
nor U7598 (N_7598,N_7207,N_7443);
xnor U7599 (N_7599,N_7024,N_7175);
nor U7600 (N_7600,N_7438,N_7022);
xor U7601 (N_7601,N_7166,N_7003);
and U7602 (N_7602,N_7491,N_7381);
xnor U7603 (N_7603,N_7067,N_7247);
and U7604 (N_7604,N_7239,N_7331);
and U7605 (N_7605,N_7126,N_7043);
and U7606 (N_7606,N_7115,N_7158);
nor U7607 (N_7607,N_7473,N_7181);
and U7608 (N_7608,N_7101,N_7350);
or U7609 (N_7609,N_7074,N_7352);
xor U7610 (N_7610,N_7372,N_7346);
and U7611 (N_7611,N_7076,N_7498);
or U7612 (N_7612,N_7338,N_7302);
xnor U7613 (N_7613,N_7185,N_7078);
xor U7614 (N_7614,N_7432,N_7413);
xor U7615 (N_7615,N_7001,N_7487);
nand U7616 (N_7616,N_7140,N_7068);
xnor U7617 (N_7617,N_7038,N_7431);
and U7618 (N_7618,N_7427,N_7478);
xor U7619 (N_7619,N_7212,N_7118);
nor U7620 (N_7620,N_7082,N_7006);
nand U7621 (N_7621,N_7441,N_7308);
xor U7622 (N_7622,N_7342,N_7469);
or U7623 (N_7623,N_7303,N_7304);
nor U7624 (N_7624,N_7476,N_7467);
nor U7625 (N_7625,N_7495,N_7447);
and U7626 (N_7626,N_7268,N_7404);
nand U7627 (N_7627,N_7206,N_7143);
nor U7628 (N_7628,N_7333,N_7192);
or U7629 (N_7629,N_7029,N_7499);
xor U7630 (N_7630,N_7011,N_7018);
or U7631 (N_7631,N_7188,N_7318);
nor U7632 (N_7632,N_7007,N_7066);
xnor U7633 (N_7633,N_7111,N_7055);
nand U7634 (N_7634,N_7391,N_7050);
nor U7635 (N_7635,N_7091,N_7489);
or U7636 (N_7636,N_7475,N_7063);
xnor U7637 (N_7637,N_7133,N_7356);
xnor U7638 (N_7638,N_7330,N_7334);
nand U7639 (N_7639,N_7035,N_7077);
and U7640 (N_7640,N_7305,N_7396);
nor U7641 (N_7641,N_7309,N_7497);
nand U7642 (N_7642,N_7172,N_7326);
and U7643 (N_7643,N_7357,N_7005);
or U7644 (N_7644,N_7327,N_7134);
nor U7645 (N_7645,N_7260,N_7398);
and U7646 (N_7646,N_7389,N_7280);
nor U7647 (N_7647,N_7136,N_7142);
nand U7648 (N_7648,N_7341,N_7058);
nor U7649 (N_7649,N_7085,N_7440);
xnor U7650 (N_7650,N_7285,N_7377);
nor U7651 (N_7651,N_7086,N_7384);
and U7652 (N_7652,N_7152,N_7336);
xor U7653 (N_7653,N_7019,N_7435);
nor U7654 (N_7654,N_7075,N_7408);
or U7655 (N_7655,N_7297,N_7228);
or U7656 (N_7656,N_7014,N_7070);
or U7657 (N_7657,N_7171,N_7096);
xnor U7658 (N_7658,N_7314,N_7016);
or U7659 (N_7659,N_7256,N_7218);
xnor U7660 (N_7660,N_7230,N_7324);
xnor U7661 (N_7661,N_7219,N_7186);
and U7662 (N_7662,N_7291,N_7065);
xnor U7663 (N_7663,N_7273,N_7390);
nand U7664 (N_7664,N_7032,N_7393);
nor U7665 (N_7665,N_7236,N_7021);
or U7666 (N_7666,N_7351,N_7255);
nand U7667 (N_7667,N_7004,N_7116);
nor U7668 (N_7668,N_7146,N_7220);
and U7669 (N_7669,N_7200,N_7300);
and U7670 (N_7670,N_7428,N_7371);
nor U7671 (N_7671,N_7040,N_7270);
nand U7672 (N_7672,N_7249,N_7272);
and U7673 (N_7673,N_7409,N_7259);
or U7674 (N_7674,N_7154,N_7229);
or U7675 (N_7675,N_7378,N_7026);
or U7676 (N_7676,N_7284,N_7462);
xor U7677 (N_7677,N_7163,N_7161);
xor U7678 (N_7678,N_7137,N_7405);
nand U7679 (N_7679,N_7092,N_7205);
or U7680 (N_7680,N_7083,N_7052);
or U7681 (N_7681,N_7149,N_7362);
nor U7682 (N_7682,N_7426,N_7369);
nor U7683 (N_7683,N_7382,N_7430);
or U7684 (N_7684,N_7162,N_7340);
xor U7685 (N_7685,N_7217,N_7416);
and U7686 (N_7686,N_7367,N_7225);
or U7687 (N_7687,N_7406,N_7248);
nor U7688 (N_7688,N_7198,N_7279);
or U7689 (N_7689,N_7442,N_7160);
nor U7690 (N_7690,N_7093,N_7319);
and U7691 (N_7691,N_7481,N_7099);
and U7692 (N_7692,N_7045,N_7262);
xor U7693 (N_7693,N_7425,N_7000);
or U7694 (N_7694,N_7100,N_7139);
nand U7695 (N_7695,N_7201,N_7328);
or U7696 (N_7696,N_7098,N_7114);
or U7697 (N_7697,N_7471,N_7286);
nor U7698 (N_7698,N_7246,N_7320);
or U7699 (N_7699,N_7124,N_7094);
and U7700 (N_7700,N_7339,N_7112);
and U7701 (N_7701,N_7087,N_7210);
xor U7702 (N_7702,N_7316,N_7233);
and U7703 (N_7703,N_7240,N_7424);
and U7704 (N_7704,N_7231,N_7031);
and U7705 (N_7705,N_7484,N_7403);
xor U7706 (N_7706,N_7271,N_7488);
and U7707 (N_7707,N_7119,N_7455);
xnor U7708 (N_7708,N_7245,N_7335);
nor U7709 (N_7709,N_7108,N_7238);
nand U7710 (N_7710,N_7293,N_7353);
and U7711 (N_7711,N_7107,N_7407);
or U7712 (N_7712,N_7283,N_7494);
or U7713 (N_7713,N_7437,N_7051);
nand U7714 (N_7714,N_7278,N_7191);
xor U7715 (N_7715,N_7177,N_7211);
or U7716 (N_7716,N_7258,N_7243);
nor U7717 (N_7717,N_7265,N_7474);
or U7718 (N_7718,N_7234,N_7423);
and U7719 (N_7719,N_7169,N_7463);
nand U7720 (N_7720,N_7144,N_7375);
or U7721 (N_7721,N_7102,N_7347);
or U7722 (N_7722,N_7081,N_7224);
or U7723 (N_7723,N_7241,N_7266);
and U7724 (N_7724,N_7244,N_7214);
nand U7725 (N_7725,N_7113,N_7033);
and U7726 (N_7726,N_7310,N_7145);
nor U7727 (N_7727,N_7329,N_7008);
nor U7728 (N_7728,N_7288,N_7223);
or U7729 (N_7729,N_7125,N_7289);
or U7730 (N_7730,N_7436,N_7456);
and U7731 (N_7731,N_7079,N_7252);
and U7732 (N_7732,N_7010,N_7472);
and U7733 (N_7733,N_7250,N_7410);
nand U7734 (N_7734,N_7397,N_7034);
nor U7735 (N_7735,N_7354,N_7422);
xnor U7736 (N_7736,N_7434,N_7321);
or U7737 (N_7737,N_7012,N_7105);
xor U7738 (N_7738,N_7411,N_7039);
xor U7739 (N_7739,N_7343,N_7313);
nor U7740 (N_7740,N_7348,N_7460);
nand U7741 (N_7741,N_7452,N_7088);
or U7742 (N_7742,N_7209,N_7013);
nand U7743 (N_7743,N_7325,N_7048);
nand U7744 (N_7744,N_7054,N_7095);
or U7745 (N_7745,N_7027,N_7361);
and U7746 (N_7746,N_7084,N_7028);
xor U7747 (N_7747,N_7056,N_7203);
and U7748 (N_7748,N_7465,N_7253);
and U7749 (N_7749,N_7274,N_7254);
nor U7750 (N_7750,N_7461,N_7024);
and U7751 (N_7751,N_7465,N_7045);
nand U7752 (N_7752,N_7387,N_7124);
nand U7753 (N_7753,N_7095,N_7290);
and U7754 (N_7754,N_7492,N_7275);
nand U7755 (N_7755,N_7306,N_7069);
or U7756 (N_7756,N_7306,N_7477);
and U7757 (N_7757,N_7187,N_7446);
or U7758 (N_7758,N_7486,N_7334);
nor U7759 (N_7759,N_7411,N_7461);
nor U7760 (N_7760,N_7433,N_7249);
or U7761 (N_7761,N_7267,N_7167);
nand U7762 (N_7762,N_7096,N_7128);
and U7763 (N_7763,N_7010,N_7116);
and U7764 (N_7764,N_7446,N_7003);
nor U7765 (N_7765,N_7133,N_7184);
nand U7766 (N_7766,N_7215,N_7267);
nor U7767 (N_7767,N_7367,N_7178);
nor U7768 (N_7768,N_7414,N_7239);
and U7769 (N_7769,N_7048,N_7125);
xor U7770 (N_7770,N_7185,N_7165);
and U7771 (N_7771,N_7017,N_7316);
nor U7772 (N_7772,N_7016,N_7330);
xnor U7773 (N_7773,N_7382,N_7289);
nor U7774 (N_7774,N_7250,N_7306);
nand U7775 (N_7775,N_7259,N_7250);
nand U7776 (N_7776,N_7004,N_7250);
nor U7777 (N_7777,N_7078,N_7083);
nand U7778 (N_7778,N_7304,N_7237);
nor U7779 (N_7779,N_7016,N_7387);
or U7780 (N_7780,N_7158,N_7080);
nand U7781 (N_7781,N_7063,N_7429);
or U7782 (N_7782,N_7045,N_7183);
nor U7783 (N_7783,N_7358,N_7079);
xnor U7784 (N_7784,N_7325,N_7198);
nor U7785 (N_7785,N_7232,N_7268);
nand U7786 (N_7786,N_7383,N_7408);
nand U7787 (N_7787,N_7098,N_7269);
xor U7788 (N_7788,N_7343,N_7433);
and U7789 (N_7789,N_7073,N_7377);
or U7790 (N_7790,N_7092,N_7095);
nor U7791 (N_7791,N_7160,N_7338);
nor U7792 (N_7792,N_7376,N_7126);
nor U7793 (N_7793,N_7284,N_7162);
xor U7794 (N_7794,N_7350,N_7274);
xnor U7795 (N_7795,N_7194,N_7054);
xor U7796 (N_7796,N_7312,N_7230);
nand U7797 (N_7797,N_7193,N_7176);
or U7798 (N_7798,N_7420,N_7167);
or U7799 (N_7799,N_7373,N_7274);
or U7800 (N_7800,N_7301,N_7459);
and U7801 (N_7801,N_7369,N_7204);
nor U7802 (N_7802,N_7187,N_7319);
or U7803 (N_7803,N_7150,N_7272);
or U7804 (N_7804,N_7134,N_7399);
and U7805 (N_7805,N_7489,N_7263);
nor U7806 (N_7806,N_7478,N_7368);
or U7807 (N_7807,N_7493,N_7232);
xor U7808 (N_7808,N_7439,N_7198);
or U7809 (N_7809,N_7245,N_7426);
or U7810 (N_7810,N_7079,N_7322);
or U7811 (N_7811,N_7070,N_7441);
or U7812 (N_7812,N_7011,N_7109);
nor U7813 (N_7813,N_7443,N_7216);
nor U7814 (N_7814,N_7336,N_7227);
xor U7815 (N_7815,N_7282,N_7220);
and U7816 (N_7816,N_7335,N_7018);
and U7817 (N_7817,N_7325,N_7489);
nor U7818 (N_7818,N_7256,N_7208);
nor U7819 (N_7819,N_7133,N_7255);
nor U7820 (N_7820,N_7418,N_7271);
or U7821 (N_7821,N_7249,N_7087);
or U7822 (N_7822,N_7120,N_7335);
nor U7823 (N_7823,N_7106,N_7356);
xor U7824 (N_7824,N_7115,N_7159);
nor U7825 (N_7825,N_7467,N_7322);
nor U7826 (N_7826,N_7374,N_7077);
or U7827 (N_7827,N_7347,N_7359);
and U7828 (N_7828,N_7038,N_7030);
or U7829 (N_7829,N_7483,N_7389);
xnor U7830 (N_7830,N_7414,N_7016);
or U7831 (N_7831,N_7483,N_7125);
or U7832 (N_7832,N_7183,N_7105);
and U7833 (N_7833,N_7168,N_7487);
nand U7834 (N_7834,N_7259,N_7463);
nor U7835 (N_7835,N_7020,N_7480);
or U7836 (N_7836,N_7362,N_7256);
xor U7837 (N_7837,N_7015,N_7041);
nor U7838 (N_7838,N_7274,N_7213);
and U7839 (N_7839,N_7383,N_7224);
and U7840 (N_7840,N_7318,N_7099);
or U7841 (N_7841,N_7190,N_7251);
and U7842 (N_7842,N_7282,N_7194);
or U7843 (N_7843,N_7392,N_7042);
nor U7844 (N_7844,N_7212,N_7417);
nor U7845 (N_7845,N_7402,N_7085);
and U7846 (N_7846,N_7027,N_7399);
and U7847 (N_7847,N_7313,N_7463);
nor U7848 (N_7848,N_7015,N_7126);
or U7849 (N_7849,N_7334,N_7003);
or U7850 (N_7850,N_7239,N_7272);
nand U7851 (N_7851,N_7421,N_7047);
nor U7852 (N_7852,N_7493,N_7003);
nand U7853 (N_7853,N_7264,N_7000);
or U7854 (N_7854,N_7041,N_7218);
nand U7855 (N_7855,N_7188,N_7238);
nand U7856 (N_7856,N_7346,N_7198);
and U7857 (N_7857,N_7055,N_7189);
and U7858 (N_7858,N_7276,N_7227);
or U7859 (N_7859,N_7004,N_7453);
xor U7860 (N_7860,N_7266,N_7357);
nand U7861 (N_7861,N_7031,N_7334);
nand U7862 (N_7862,N_7121,N_7271);
and U7863 (N_7863,N_7391,N_7059);
nand U7864 (N_7864,N_7466,N_7095);
and U7865 (N_7865,N_7221,N_7120);
or U7866 (N_7866,N_7114,N_7408);
or U7867 (N_7867,N_7328,N_7006);
and U7868 (N_7868,N_7498,N_7462);
nor U7869 (N_7869,N_7173,N_7073);
and U7870 (N_7870,N_7044,N_7098);
nand U7871 (N_7871,N_7046,N_7284);
nand U7872 (N_7872,N_7266,N_7268);
nand U7873 (N_7873,N_7209,N_7126);
nand U7874 (N_7874,N_7284,N_7089);
xnor U7875 (N_7875,N_7494,N_7259);
nor U7876 (N_7876,N_7035,N_7369);
nor U7877 (N_7877,N_7487,N_7488);
xor U7878 (N_7878,N_7380,N_7349);
nor U7879 (N_7879,N_7038,N_7482);
and U7880 (N_7880,N_7017,N_7487);
nor U7881 (N_7881,N_7023,N_7002);
xor U7882 (N_7882,N_7363,N_7429);
nand U7883 (N_7883,N_7310,N_7000);
and U7884 (N_7884,N_7126,N_7330);
xor U7885 (N_7885,N_7321,N_7415);
or U7886 (N_7886,N_7012,N_7310);
nand U7887 (N_7887,N_7108,N_7268);
nand U7888 (N_7888,N_7102,N_7350);
or U7889 (N_7889,N_7384,N_7202);
and U7890 (N_7890,N_7493,N_7027);
nor U7891 (N_7891,N_7427,N_7239);
nor U7892 (N_7892,N_7270,N_7071);
nand U7893 (N_7893,N_7298,N_7216);
nand U7894 (N_7894,N_7219,N_7463);
and U7895 (N_7895,N_7010,N_7202);
and U7896 (N_7896,N_7179,N_7347);
or U7897 (N_7897,N_7240,N_7206);
nor U7898 (N_7898,N_7330,N_7380);
xnor U7899 (N_7899,N_7023,N_7110);
nand U7900 (N_7900,N_7465,N_7032);
nand U7901 (N_7901,N_7419,N_7430);
xor U7902 (N_7902,N_7132,N_7036);
xnor U7903 (N_7903,N_7294,N_7267);
xor U7904 (N_7904,N_7030,N_7307);
xnor U7905 (N_7905,N_7406,N_7367);
nor U7906 (N_7906,N_7452,N_7254);
and U7907 (N_7907,N_7461,N_7237);
nor U7908 (N_7908,N_7285,N_7398);
xnor U7909 (N_7909,N_7377,N_7061);
xnor U7910 (N_7910,N_7226,N_7023);
nand U7911 (N_7911,N_7173,N_7232);
xnor U7912 (N_7912,N_7085,N_7012);
xor U7913 (N_7913,N_7457,N_7109);
nand U7914 (N_7914,N_7382,N_7221);
or U7915 (N_7915,N_7489,N_7033);
nor U7916 (N_7916,N_7361,N_7001);
or U7917 (N_7917,N_7106,N_7226);
xnor U7918 (N_7918,N_7128,N_7004);
or U7919 (N_7919,N_7379,N_7138);
or U7920 (N_7920,N_7451,N_7195);
nor U7921 (N_7921,N_7215,N_7422);
or U7922 (N_7922,N_7484,N_7273);
and U7923 (N_7923,N_7301,N_7070);
xor U7924 (N_7924,N_7375,N_7344);
nor U7925 (N_7925,N_7153,N_7434);
xor U7926 (N_7926,N_7254,N_7156);
xor U7927 (N_7927,N_7212,N_7327);
xor U7928 (N_7928,N_7254,N_7066);
and U7929 (N_7929,N_7257,N_7081);
nor U7930 (N_7930,N_7073,N_7425);
xor U7931 (N_7931,N_7495,N_7163);
xor U7932 (N_7932,N_7317,N_7365);
nor U7933 (N_7933,N_7262,N_7036);
nand U7934 (N_7934,N_7454,N_7252);
nand U7935 (N_7935,N_7432,N_7077);
or U7936 (N_7936,N_7384,N_7256);
and U7937 (N_7937,N_7367,N_7045);
or U7938 (N_7938,N_7181,N_7009);
or U7939 (N_7939,N_7413,N_7018);
nand U7940 (N_7940,N_7283,N_7268);
nand U7941 (N_7941,N_7147,N_7330);
or U7942 (N_7942,N_7251,N_7160);
nor U7943 (N_7943,N_7011,N_7007);
or U7944 (N_7944,N_7238,N_7359);
nor U7945 (N_7945,N_7179,N_7107);
nor U7946 (N_7946,N_7196,N_7009);
and U7947 (N_7947,N_7444,N_7300);
and U7948 (N_7948,N_7181,N_7220);
and U7949 (N_7949,N_7459,N_7381);
nand U7950 (N_7950,N_7085,N_7487);
nand U7951 (N_7951,N_7370,N_7333);
nand U7952 (N_7952,N_7378,N_7328);
xnor U7953 (N_7953,N_7212,N_7497);
nor U7954 (N_7954,N_7478,N_7075);
nor U7955 (N_7955,N_7164,N_7447);
and U7956 (N_7956,N_7344,N_7320);
or U7957 (N_7957,N_7356,N_7193);
nor U7958 (N_7958,N_7064,N_7263);
or U7959 (N_7959,N_7229,N_7069);
and U7960 (N_7960,N_7271,N_7457);
nor U7961 (N_7961,N_7438,N_7016);
or U7962 (N_7962,N_7403,N_7071);
and U7963 (N_7963,N_7029,N_7463);
nand U7964 (N_7964,N_7228,N_7356);
and U7965 (N_7965,N_7130,N_7149);
nor U7966 (N_7966,N_7445,N_7270);
nor U7967 (N_7967,N_7276,N_7191);
nand U7968 (N_7968,N_7414,N_7427);
and U7969 (N_7969,N_7303,N_7326);
and U7970 (N_7970,N_7319,N_7065);
or U7971 (N_7971,N_7465,N_7219);
nor U7972 (N_7972,N_7069,N_7178);
xor U7973 (N_7973,N_7469,N_7201);
nor U7974 (N_7974,N_7343,N_7318);
nand U7975 (N_7975,N_7285,N_7354);
xor U7976 (N_7976,N_7362,N_7282);
or U7977 (N_7977,N_7362,N_7411);
and U7978 (N_7978,N_7368,N_7232);
or U7979 (N_7979,N_7000,N_7216);
xnor U7980 (N_7980,N_7378,N_7392);
xnor U7981 (N_7981,N_7086,N_7408);
xnor U7982 (N_7982,N_7249,N_7165);
xor U7983 (N_7983,N_7350,N_7134);
nand U7984 (N_7984,N_7006,N_7034);
or U7985 (N_7985,N_7070,N_7068);
or U7986 (N_7986,N_7049,N_7172);
or U7987 (N_7987,N_7029,N_7008);
nand U7988 (N_7988,N_7387,N_7214);
nand U7989 (N_7989,N_7426,N_7163);
and U7990 (N_7990,N_7139,N_7199);
xnor U7991 (N_7991,N_7231,N_7486);
nand U7992 (N_7992,N_7010,N_7486);
and U7993 (N_7993,N_7498,N_7061);
xnor U7994 (N_7994,N_7220,N_7163);
nand U7995 (N_7995,N_7192,N_7456);
or U7996 (N_7996,N_7417,N_7163);
and U7997 (N_7997,N_7482,N_7387);
nand U7998 (N_7998,N_7005,N_7073);
and U7999 (N_7999,N_7485,N_7231);
nor U8000 (N_8000,N_7565,N_7626);
xnor U8001 (N_8001,N_7514,N_7775);
xnor U8002 (N_8002,N_7559,N_7687);
and U8003 (N_8003,N_7892,N_7958);
xnor U8004 (N_8004,N_7532,N_7543);
xnor U8005 (N_8005,N_7686,N_7880);
or U8006 (N_8006,N_7818,N_7595);
nor U8007 (N_8007,N_7506,N_7799);
and U8008 (N_8008,N_7986,N_7743);
xnor U8009 (N_8009,N_7871,N_7710);
nand U8010 (N_8010,N_7918,N_7522);
and U8011 (N_8011,N_7531,N_7689);
xnor U8012 (N_8012,N_7549,N_7624);
xnor U8013 (N_8013,N_7648,N_7682);
nor U8014 (N_8014,N_7589,N_7823);
xnor U8015 (N_8015,N_7608,N_7616);
and U8016 (N_8016,N_7784,N_7936);
and U8017 (N_8017,N_7778,N_7951);
xor U8018 (N_8018,N_7696,N_7852);
or U8019 (N_8019,N_7859,N_7867);
nand U8020 (N_8020,N_7874,N_7932);
nand U8021 (N_8021,N_7917,N_7903);
and U8022 (N_8022,N_7947,N_7795);
and U8023 (N_8023,N_7929,N_7792);
nand U8024 (N_8024,N_7647,N_7649);
and U8025 (N_8025,N_7965,N_7629);
xnor U8026 (N_8026,N_7598,N_7521);
xnor U8027 (N_8027,N_7864,N_7612);
and U8028 (N_8028,N_7806,N_7617);
and U8029 (N_8029,N_7691,N_7828);
xnor U8030 (N_8030,N_7955,N_7935);
nand U8031 (N_8031,N_7734,N_7782);
nand U8032 (N_8032,N_7976,N_7953);
and U8033 (N_8033,N_7827,N_7961);
nand U8034 (N_8034,N_7798,N_7633);
nor U8035 (N_8035,N_7848,N_7754);
nor U8036 (N_8036,N_7893,N_7911);
and U8037 (N_8037,N_7540,N_7830);
nand U8038 (N_8038,N_7943,N_7855);
nor U8039 (N_8039,N_7685,N_7980);
nor U8040 (N_8040,N_7739,N_7501);
nor U8041 (N_8041,N_7677,N_7923);
or U8042 (N_8042,N_7785,N_7846);
nor U8043 (N_8043,N_7789,N_7581);
xor U8044 (N_8044,N_7679,N_7749);
nor U8045 (N_8045,N_7946,N_7535);
nand U8046 (N_8046,N_7908,N_7721);
and U8047 (N_8047,N_7740,N_7518);
nand U8048 (N_8048,N_7611,N_7551);
and U8049 (N_8049,N_7809,N_7578);
xor U8050 (N_8050,N_7653,N_7610);
nor U8051 (N_8051,N_7523,N_7954);
and U8052 (N_8052,N_7618,N_7674);
nor U8053 (N_8053,N_7991,N_7796);
nor U8054 (N_8054,N_7952,N_7534);
nand U8055 (N_8055,N_7845,N_7662);
xnor U8056 (N_8056,N_7762,N_7969);
or U8057 (N_8057,N_7832,N_7652);
and U8058 (N_8058,N_7605,N_7547);
nor U8059 (N_8059,N_7994,N_7715);
xor U8060 (N_8060,N_7949,N_7901);
xor U8061 (N_8061,N_7810,N_7684);
nand U8062 (N_8062,N_7841,N_7517);
xor U8063 (N_8063,N_7770,N_7794);
or U8064 (N_8064,N_7621,N_7930);
and U8065 (N_8065,N_7704,N_7613);
nand U8066 (N_8066,N_7902,N_7819);
or U8067 (N_8067,N_7977,N_7519);
or U8068 (N_8068,N_7698,N_7676);
xnor U8069 (N_8069,N_7758,N_7881);
xor U8070 (N_8070,N_7764,N_7590);
nand U8071 (N_8071,N_7886,N_7574);
nand U8072 (N_8072,N_7926,N_7971);
nand U8073 (N_8073,N_7808,N_7709);
xor U8074 (N_8074,N_7887,N_7722);
xnor U8075 (N_8075,N_7931,N_7509);
and U8076 (N_8076,N_7592,N_7718);
or U8077 (N_8077,N_7694,N_7913);
xnor U8078 (N_8078,N_7587,N_7548);
nor U8079 (N_8079,N_7620,N_7642);
and U8080 (N_8080,N_7673,N_7640);
and U8081 (N_8081,N_7757,N_7964);
or U8082 (N_8082,N_7561,N_7688);
xnor U8083 (N_8083,N_7525,N_7868);
or U8084 (N_8084,N_7815,N_7856);
or U8085 (N_8085,N_7787,N_7727);
nor U8086 (N_8086,N_7860,N_7761);
or U8087 (N_8087,N_7714,N_7631);
or U8088 (N_8088,N_7777,N_7712);
nand U8089 (N_8089,N_7672,N_7670);
nand U8090 (N_8090,N_7550,N_7767);
xnor U8091 (N_8091,N_7713,N_7570);
xor U8092 (N_8092,N_7733,N_7656);
nor U8093 (N_8093,N_7847,N_7566);
nand U8094 (N_8094,N_7584,N_7690);
nand U8095 (N_8095,N_7527,N_7728);
nand U8096 (N_8096,N_7599,N_7512);
xnor U8097 (N_8097,N_7801,N_7800);
and U8098 (N_8098,N_7650,N_7663);
and U8099 (N_8099,N_7602,N_7862);
and U8100 (N_8100,N_7884,N_7507);
nor U8101 (N_8101,N_7934,N_7813);
or U8102 (N_8102,N_7836,N_7972);
or U8103 (N_8103,N_7513,N_7904);
xor U8104 (N_8104,N_7744,N_7779);
xnor U8105 (N_8105,N_7555,N_7863);
and U8106 (N_8106,N_7962,N_7563);
or U8107 (N_8107,N_7707,N_7987);
nand U8108 (N_8108,N_7791,N_7600);
nor U8109 (N_8109,N_7924,N_7760);
or U8110 (N_8110,N_7948,N_7582);
or U8111 (N_8111,N_7984,N_7771);
nor U8112 (N_8112,N_7556,N_7831);
or U8113 (N_8113,N_7637,N_7838);
nand U8114 (N_8114,N_7788,N_7735);
nand U8115 (N_8115,N_7865,N_7752);
nor U8116 (N_8116,N_7857,N_7664);
and U8117 (N_8117,N_7639,N_7692);
xor U8118 (N_8118,N_7843,N_7607);
and U8119 (N_8119,N_7866,N_7719);
nor U8120 (N_8120,N_7996,N_7768);
and U8121 (N_8121,N_7805,N_7928);
xnor U8122 (N_8122,N_7835,N_7585);
or U8123 (N_8123,N_7909,N_7897);
nor U8124 (N_8124,N_7981,N_7746);
and U8125 (N_8125,N_7655,N_7572);
nor U8126 (N_8126,N_7644,N_7729);
nand U8127 (N_8127,N_7554,N_7993);
or U8128 (N_8128,N_7877,N_7957);
or U8129 (N_8129,N_7837,N_7628);
and U8130 (N_8130,N_7940,N_7938);
nor U8131 (N_8131,N_7573,N_7705);
xnor U8132 (N_8132,N_7944,N_7678);
and U8133 (N_8133,N_7973,N_7533);
and U8134 (N_8134,N_7680,N_7671);
or U8135 (N_8135,N_7623,N_7668);
or U8136 (N_8136,N_7583,N_7557);
or U8137 (N_8137,N_7515,N_7634);
nand U8138 (N_8138,N_7769,N_7569);
nand U8139 (N_8139,N_7726,N_7576);
xnor U8140 (N_8140,N_7790,N_7919);
nor U8141 (N_8141,N_7748,N_7500);
nor U8142 (N_8142,N_7807,N_7888);
or U8143 (N_8143,N_7822,N_7502);
nand U8144 (N_8144,N_7783,N_7907);
xnor U8145 (N_8145,N_7833,N_7520);
xnor U8146 (N_8146,N_7669,N_7898);
xor U8147 (N_8147,N_7516,N_7627);
or U8148 (N_8148,N_7596,N_7594);
xnor U8149 (N_8149,N_7839,N_7606);
nand U8150 (N_8150,N_7890,N_7979);
nor U8151 (N_8151,N_7895,N_7651);
or U8152 (N_8152,N_7916,N_7829);
or U8153 (N_8153,N_7701,N_7503);
nor U8154 (N_8154,N_7797,N_7537);
nor U8155 (N_8155,N_7699,N_7879);
nand U8156 (N_8156,N_7854,N_7568);
and U8157 (N_8157,N_7586,N_7635);
or U8158 (N_8158,N_7660,N_7723);
nand U8159 (N_8159,N_7840,N_7530);
and U8160 (N_8160,N_7505,N_7869);
nor U8161 (N_8161,N_7542,N_7661);
and U8162 (N_8162,N_7541,N_7910);
nand U8163 (N_8163,N_7885,N_7774);
or U8164 (N_8164,N_7646,N_7636);
nand U8165 (N_8165,N_7967,N_7816);
and U8166 (N_8166,N_7745,N_7683);
nor U8167 (N_8167,N_7804,N_7659);
xor U8168 (N_8168,N_7853,N_7510);
xor U8169 (N_8169,N_7968,N_7759);
or U8170 (N_8170,N_7703,N_7755);
nor U8171 (N_8171,N_7997,N_7876);
and U8172 (N_8172,N_7825,N_7803);
and U8173 (N_8173,N_7614,N_7643);
nand U8174 (N_8174,N_7658,N_7738);
nand U8175 (N_8175,N_7546,N_7702);
xnor U8176 (N_8176,N_7905,N_7978);
and U8177 (N_8177,N_7942,N_7939);
nand U8178 (N_8178,N_7882,N_7922);
or U8179 (N_8179,N_7850,N_7878);
and U8180 (N_8180,N_7750,N_7988);
nor U8181 (N_8181,N_7921,N_7657);
xor U8182 (N_8182,N_7700,N_7553);
or U8183 (N_8183,N_7511,N_7870);
or U8184 (N_8184,N_7894,N_7579);
or U8185 (N_8185,N_7970,N_7708);
and U8186 (N_8186,N_7544,N_7737);
or U8187 (N_8187,N_7889,N_7725);
xor U8188 (N_8188,N_7645,N_7802);
and U8189 (N_8189,N_7912,N_7619);
nor U8190 (N_8190,N_7577,N_7529);
nor U8191 (N_8191,N_7667,N_7925);
nand U8192 (N_8192,N_7593,N_7834);
nand U8193 (N_8193,N_7766,N_7588);
nor U8194 (N_8194,N_7772,N_7844);
xor U8195 (N_8195,N_7504,N_7601);
nand U8196 (N_8196,N_7851,N_7604);
and U8197 (N_8197,N_7820,N_7883);
nand U8198 (N_8198,N_7591,N_7781);
and U8199 (N_8199,N_7695,N_7539);
nor U8200 (N_8200,N_7985,N_7567);
and U8201 (N_8201,N_7983,N_7975);
or U8202 (N_8202,N_7927,N_7950);
or U8203 (N_8203,N_7575,N_7524);
xnor U8204 (N_8204,N_7697,N_7960);
nand U8205 (N_8205,N_7625,N_7990);
and U8206 (N_8206,N_7641,N_7811);
xnor U8207 (N_8207,N_7861,N_7681);
or U8208 (N_8208,N_7793,N_7724);
xnor U8209 (N_8209,N_7742,N_7992);
nor U8210 (N_8210,N_7609,N_7941);
nor U8211 (N_8211,N_7900,N_7817);
and U8212 (N_8212,N_7933,N_7873);
or U8213 (N_8213,N_7536,N_7824);
xnor U8214 (N_8214,N_7716,N_7693);
and U8215 (N_8215,N_7622,N_7736);
or U8216 (N_8216,N_7508,N_7821);
and U8217 (N_8217,N_7763,N_7632);
xnor U8218 (N_8218,N_7751,N_7914);
nand U8219 (N_8219,N_7891,N_7776);
xnor U8220 (N_8220,N_7753,N_7571);
or U8221 (N_8221,N_7666,N_7920);
nor U8222 (N_8222,N_7731,N_7741);
or U8223 (N_8223,N_7717,N_7937);
xnor U8224 (N_8224,N_7526,N_7603);
nand U8225 (N_8225,N_7773,N_7558);
and U8226 (N_8226,N_7654,N_7786);
nand U8227 (N_8227,N_7959,N_7597);
nor U8228 (N_8228,N_7720,N_7999);
nand U8229 (N_8229,N_7899,N_7906);
and U8230 (N_8230,N_7765,N_7812);
nand U8231 (N_8231,N_7956,N_7747);
and U8232 (N_8232,N_7552,N_7963);
nor U8233 (N_8233,N_7732,N_7982);
nand U8234 (N_8234,N_7638,N_7528);
and U8235 (N_8235,N_7615,N_7989);
nor U8236 (N_8236,N_7826,N_7730);
nand U8237 (N_8237,N_7562,N_7974);
xor U8238 (N_8238,N_7756,N_7538);
nor U8239 (N_8239,N_7711,N_7780);
xnor U8240 (N_8240,N_7545,N_7945);
nor U8241 (N_8241,N_7966,N_7665);
xnor U8242 (N_8242,N_7858,N_7814);
nand U8243 (N_8243,N_7896,N_7849);
nand U8244 (N_8244,N_7706,N_7872);
xnor U8245 (N_8245,N_7564,N_7998);
nand U8246 (N_8246,N_7915,N_7875);
and U8247 (N_8247,N_7995,N_7630);
nand U8248 (N_8248,N_7580,N_7842);
nor U8249 (N_8249,N_7560,N_7675);
xnor U8250 (N_8250,N_7849,N_7682);
or U8251 (N_8251,N_7991,N_7580);
nor U8252 (N_8252,N_7772,N_7631);
nand U8253 (N_8253,N_7509,N_7584);
nand U8254 (N_8254,N_7710,N_7540);
xor U8255 (N_8255,N_7984,N_7892);
nand U8256 (N_8256,N_7779,N_7986);
xor U8257 (N_8257,N_7863,N_7648);
and U8258 (N_8258,N_7828,N_7835);
nor U8259 (N_8259,N_7870,N_7876);
xnor U8260 (N_8260,N_7922,N_7600);
and U8261 (N_8261,N_7844,N_7516);
nand U8262 (N_8262,N_7990,N_7941);
xnor U8263 (N_8263,N_7844,N_7984);
or U8264 (N_8264,N_7613,N_7632);
nor U8265 (N_8265,N_7913,N_7923);
nor U8266 (N_8266,N_7609,N_7506);
and U8267 (N_8267,N_7867,N_7717);
nand U8268 (N_8268,N_7539,N_7698);
nor U8269 (N_8269,N_7839,N_7713);
and U8270 (N_8270,N_7758,N_7837);
xnor U8271 (N_8271,N_7642,N_7998);
nand U8272 (N_8272,N_7661,N_7958);
xnor U8273 (N_8273,N_7944,N_7948);
xnor U8274 (N_8274,N_7940,N_7535);
xor U8275 (N_8275,N_7739,N_7957);
xor U8276 (N_8276,N_7992,N_7736);
or U8277 (N_8277,N_7698,N_7835);
and U8278 (N_8278,N_7962,N_7983);
and U8279 (N_8279,N_7723,N_7708);
nor U8280 (N_8280,N_7578,N_7789);
and U8281 (N_8281,N_7910,N_7949);
or U8282 (N_8282,N_7628,N_7626);
nor U8283 (N_8283,N_7526,N_7869);
nand U8284 (N_8284,N_7758,N_7715);
xnor U8285 (N_8285,N_7846,N_7943);
or U8286 (N_8286,N_7896,N_7764);
nor U8287 (N_8287,N_7506,N_7514);
nor U8288 (N_8288,N_7756,N_7967);
nor U8289 (N_8289,N_7688,N_7822);
nor U8290 (N_8290,N_7760,N_7737);
nand U8291 (N_8291,N_7706,N_7566);
nor U8292 (N_8292,N_7604,N_7731);
nor U8293 (N_8293,N_7846,N_7818);
and U8294 (N_8294,N_7553,N_7650);
nand U8295 (N_8295,N_7547,N_7763);
and U8296 (N_8296,N_7929,N_7800);
or U8297 (N_8297,N_7512,N_7981);
xnor U8298 (N_8298,N_7688,N_7618);
xor U8299 (N_8299,N_7664,N_7902);
or U8300 (N_8300,N_7877,N_7544);
and U8301 (N_8301,N_7618,N_7847);
or U8302 (N_8302,N_7655,N_7635);
nand U8303 (N_8303,N_7800,N_7589);
nand U8304 (N_8304,N_7959,N_7950);
or U8305 (N_8305,N_7854,N_7839);
xnor U8306 (N_8306,N_7699,N_7920);
or U8307 (N_8307,N_7776,N_7535);
or U8308 (N_8308,N_7986,N_7937);
or U8309 (N_8309,N_7788,N_7510);
xor U8310 (N_8310,N_7581,N_7829);
or U8311 (N_8311,N_7862,N_7535);
or U8312 (N_8312,N_7884,N_7861);
nor U8313 (N_8313,N_7574,N_7749);
nand U8314 (N_8314,N_7507,N_7898);
nand U8315 (N_8315,N_7621,N_7948);
or U8316 (N_8316,N_7724,N_7633);
or U8317 (N_8317,N_7707,N_7864);
or U8318 (N_8318,N_7745,N_7895);
nor U8319 (N_8319,N_7630,N_7697);
nand U8320 (N_8320,N_7731,N_7885);
or U8321 (N_8321,N_7949,N_7858);
and U8322 (N_8322,N_7635,N_7900);
nor U8323 (N_8323,N_7594,N_7723);
and U8324 (N_8324,N_7686,N_7738);
xnor U8325 (N_8325,N_7690,N_7678);
and U8326 (N_8326,N_7601,N_7778);
nor U8327 (N_8327,N_7948,N_7743);
nor U8328 (N_8328,N_7865,N_7630);
or U8329 (N_8329,N_7833,N_7581);
nor U8330 (N_8330,N_7666,N_7758);
or U8331 (N_8331,N_7552,N_7786);
or U8332 (N_8332,N_7938,N_7945);
nor U8333 (N_8333,N_7646,N_7786);
xor U8334 (N_8334,N_7800,N_7653);
and U8335 (N_8335,N_7879,N_7565);
and U8336 (N_8336,N_7935,N_7766);
xnor U8337 (N_8337,N_7977,N_7751);
nor U8338 (N_8338,N_7768,N_7612);
nor U8339 (N_8339,N_7632,N_7890);
nand U8340 (N_8340,N_7753,N_7955);
or U8341 (N_8341,N_7847,N_7504);
nor U8342 (N_8342,N_7557,N_7712);
and U8343 (N_8343,N_7780,N_7662);
xnor U8344 (N_8344,N_7644,N_7826);
or U8345 (N_8345,N_7521,N_7803);
and U8346 (N_8346,N_7856,N_7792);
or U8347 (N_8347,N_7892,N_7930);
and U8348 (N_8348,N_7842,N_7737);
xnor U8349 (N_8349,N_7918,N_7604);
nor U8350 (N_8350,N_7679,N_7805);
nand U8351 (N_8351,N_7961,N_7927);
or U8352 (N_8352,N_7586,N_7684);
and U8353 (N_8353,N_7606,N_7747);
or U8354 (N_8354,N_7755,N_7934);
xor U8355 (N_8355,N_7539,N_7918);
xnor U8356 (N_8356,N_7821,N_7608);
nor U8357 (N_8357,N_7772,N_7833);
and U8358 (N_8358,N_7693,N_7890);
nand U8359 (N_8359,N_7860,N_7960);
xor U8360 (N_8360,N_7778,N_7731);
nand U8361 (N_8361,N_7643,N_7574);
nor U8362 (N_8362,N_7554,N_7921);
nor U8363 (N_8363,N_7998,N_7582);
and U8364 (N_8364,N_7564,N_7928);
or U8365 (N_8365,N_7732,N_7971);
and U8366 (N_8366,N_7725,N_7799);
and U8367 (N_8367,N_7879,N_7979);
xor U8368 (N_8368,N_7563,N_7502);
nand U8369 (N_8369,N_7634,N_7503);
xor U8370 (N_8370,N_7934,N_7883);
nand U8371 (N_8371,N_7803,N_7962);
and U8372 (N_8372,N_7626,N_7782);
nand U8373 (N_8373,N_7759,N_7716);
and U8374 (N_8374,N_7561,N_7749);
or U8375 (N_8375,N_7989,N_7901);
and U8376 (N_8376,N_7990,N_7888);
xor U8377 (N_8377,N_7633,N_7875);
and U8378 (N_8378,N_7953,N_7511);
nand U8379 (N_8379,N_7916,N_7929);
or U8380 (N_8380,N_7984,N_7961);
or U8381 (N_8381,N_7759,N_7794);
or U8382 (N_8382,N_7822,N_7821);
xor U8383 (N_8383,N_7686,N_7901);
nor U8384 (N_8384,N_7906,N_7653);
nor U8385 (N_8385,N_7865,N_7863);
nand U8386 (N_8386,N_7524,N_7772);
and U8387 (N_8387,N_7651,N_7928);
nor U8388 (N_8388,N_7905,N_7628);
and U8389 (N_8389,N_7973,N_7702);
or U8390 (N_8390,N_7913,N_7699);
nor U8391 (N_8391,N_7980,N_7665);
or U8392 (N_8392,N_7926,N_7718);
nand U8393 (N_8393,N_7700,N_7647);
nor U8394 (N_8394,N_7902,N_7878);
nor U8395 (N_8395,N_7620,N_7575);
nor U8396 (N_8396,N_7741,N_7775);
xnor U8397 (N_8397,N_7782,N_7993);
nand U8398 (N_8398,N_7507,N_7606);
or U8399 (N_8399,N_7901,N_7775);
nand U8400 (N_8400,N_7664,N_7748);
nor U8401 (N_8401,N_7577,N_7986);
xor U8402 (N_8402,N_7881,N_7998);
or U8403 (N_8403,N_7968,N_7650);
nand U8404 (N_8404,N_7869,N_7551);
nand U8405 (N_8405,N_7654,N_7939);
nor U8406 (N_8406,N_7920,N_7616);
nor U8407 (N_8407,N_7569,N_7750);
nand U8408 (N_8408,N_7931,N_7854);
nor U8409 (N_8409,N_7862,N_7848);
nand U8410 (N_8410,N_7957,N_7637);
nor U8411 (N_8411,N_7940,N_7591);
or U8412 (N_8412,N_7714,N_7935);
nor U8413 (N_8413,N_7600,N_7797);
or U8414 (N_8414,N_7807,N_7688);
nor U8415 (N_8415,N_7661,N_7590);
and U8416 (N_8416,N_7839,N_7905);
nand U8417 (N_8417,N_7647,N_7943);
or U8418 (N_8418,N_7758,N_7511);
nor U8419 (N_8419,N_7559,N_7802);
nand U8420 (N_8420,N_7577,N_7556);
xnor U8421 (N_8421,N_7953,N_7968);
xor U8422 (N_8422,N_7931,N_7534);
and U8423 (N_8423,N_7573,N_7738);
nand U8424 (N_8424,N_7869,N_7537);
xnor U8425 (N_8425,N_7729,N_7945);
nor U8426 (N_8426,N_7892,N_7781);
nand U8427 (N_8427,N_7690,N_7601);
or U8428 (N_8428,N_7538,N_7615);
nand U8429 (N_8429,N_7885,N_7506);
nand U8430 (N_8430,N_7746,N_7679);
xor U8431 (N_8431,N_7543,N_7923);
nor U8432 (N_8432,N_7709,N_7760);
or U8433 (N_8433,N_7760,N_7735);
or U8434 (N_8434,N_7559,N_7882);
nor U8435 (N_8435,N_7559,N_7864);
and U8436 (N_8436,N_7566,N_7878);
nor U8437 (N_8437,N_7781,N_7803);
nor U8438 (N_8438,N_7926,N_7741);
xnor U8439 (N_8439,N_7562,N_7886);
and U8440 (N_8440,N_7947,N_7561);
nor U8441 (N_8441,N_7586,N_7993);
xor U8442 (N_8442,N_7615,N_7828);
and U8443 (N_8443,N_7512,N_7623);
or U8444 (N_8444,N_7535,N_7931);
xor U8445 (N_8445,N_7600,N_7831);
xnor U8446 (N_8446,N_7661,N_7783);
nand U8447 (N_8447,N_7711,N_7958);
xnor U8448 (N_8448,N_7557,N_7574);
or U8449 (N_8449,N_7915,N_7636);
nand U8450 (N_8450,N_7852,N_7693);
nand U8451 (N_8451,N_7687,N_7572);
and U8452 (N_8452,N_7713,N_7969);
and U8453 (N_8453,N_7621,N_7534);
or U8454 (N_8454,N_7746,N_7919);
and U8455 (N_8455,N_7561,N_7678);
or U8456 (N_8456,N_7559,N_7974);
nor U8457 (N_8457,N_7768,N_7959);
nand U8458 (N_8458,N_7930,N_7532);
nand U8459 (N_8459,N_7767,N_7835);
or U8460 (N_8460,N_7869,N_7804);
or U8461 (N_8461,N_7762,N_7813);
xnor U8462 (N_8462,N_7663,N_7706);
nor U8463 (N_8463,N_7656,N_7705);
or U8464 (N_8464,N_7955,N_7983);
and U8465 (N_8465,N_7578,N_7983);
nand U8466 (N_8466,N_7987,N_7797);
nor U8467 (N_8467,N_7582,N_7721);
xor U8468 (N_8468,N_7537,N_7861);
nand U8469 (N_8469,N_7574,N_7815);
nand U8470 (N_8470,N_7889,N_7555);
xnor U8471 (N_8471,N_7794,N_7678);
or U8472 (N_8472,N_7641,N_7580);
xor U8473 (N_8473,N_7760,N_7652);
and U8474 (N_8474,N_7929,N_7837);
and U8475 (N_8475,N_7828,N_7933);
and U8476 (N_8476,N_7736,N_7956);
and U8477 (N_8477,N_7820,N_7723);
or U8478 (N_8478,N_7898,N_7591);
and U8479 (N_8479,N_7675,N_7978);
nand U8480 (N_8480,N_7871,N_7799);
and U8481 (N_8481,N_7667,N_7888);
or U8482 (N_8482,N_7829,N_7623);
or U8483 (N_8483,N_7906,N_7913);
nand U8484 (N_8484,N_7556,N_7593);
and U8485 (N_8485,N_7727,N_7615);
and U8486 (N_8486,N_7742,N_7980);
and U8487 (N_8487,N_7810,N_7879);
or U8488 (N_8488,N_7574,N_7773);
and U8489 (N_8489,N_7698,N_7791);
xnor U8490 (N_8490,N_7604,N_7966);
or U8491 (N_8491,N_7615,N_7922);
nor U8492 (N_8492,N_7855,N_7517);
or U8493 (N_8493,N_7777,N_7573);
nand U8494 (N_8494,N_7701,N_7980);
nand U8495 (N_8495,N_7923,N_7827);
xnor U8496 (N_8496,N_7939,N_7675);
xor U8497 (N_8497,N_7513,N_7654);
and U8498 (N_8498,N_7778,N_7554);
nor U8499 (N_8499,N_7944,N_7583);
nand U8500 (N_8500,N_8300,N_8388);
nand U8501 (N_8501,N_8231,N_8368);
nand U8502 (N_8502,N_8022,N_8271);
or U8503 (N_8503,N_8083,N_8427);
nor U8504 (N_8504,N_8445,N_8342);
or U8505 (N_8505,N_8493,N_8356);
nor U8506 (N_8506,N_8030,N_8399);
nor U8507 (N_8507,N_8261,N_8216);
nor U8508 (N_8508,N_8260,N_8277);
nand U8509 (N_8509,N_8064,N_8471);
nor U8510 (N_8510,N_8447,N_8486);
or U8511 (N_8511,N_8332,N_8213);
nand U8512 (N_8512,N_8351,N_8166);
nor U8513 (N_8513,N_8264,N_8115);
nand U8514 (N_8514,N_8498,N_8311);
or U8515 (N_8515,N_8331,N_8034);
nand U8516 (N_8516,N_8262,N_8473);
nor U8517 (N_8517,N_8167,N_8379);
and U8518 (N_8518,N_8048,N_8164);
xnor U8519 (N_8519,N_8067,N_8403);
xnor U8520 (N_8520,N_8198,N_8093);
nor U8521 (N_8521,N_8484,N_8131);
nand U8522 (N_8522,N_8393,N_8138);
or U8523 (N_8523,N_8060,N_8318);
or U8524 (N_8524,N_8135,N_8426);
or U8525 (N_8525,N_8220,N_8481);
and U8526 (N_8526,N_8172,N_8469);
and U8527 (N_8527,N_8415,N_8100);
or U8528 (N_8528,N_8329,N_8401);
nand U8529 (N_8529,N_8487,N_8425);
nor U8530 (N_8530,N_8025,N_8299);
nor U8531 (N_8531,N_8459,N_8126);
nor U8532 (N_8532,N_8363,N_8139);
nor U8533 (N_8533,N_8346,N_8273);
nand U8534 (N_8534,N_8463,N_8149);
nor U8535 (N_8535,N_8389,N_8298);
and U8536 (N_8536,N_8244,N_8287);
nor U8537 (N_8537,N_8091,N_8122);
xnor U8538 (N_8538,N_8250,N_8457);
and U8539 (N_8539,N_8171,N_8058);
xor U8540 (N_8540,N_8012,N_8482);
and U8541 (N_8541,N_8191,N_8321);
nor U8542 (N_8542,N_8499,N_8162);
and U8543 (N_8543,N_8263,N_8188);
nor U8544 (N_8544,N_8328,N_8002);
xnor U8545 (N_8545,N_8113,N_8327);
xor U8546 (N_8546,N_8392,N_8380);
nand U8547 (N_8547,N_8458,N_8047);
xor U8548 (N_8548,N_8108,N_8404);
xnor U8549 (N_8549,N_8312,N_8133);
xor U8550 (N_8550,N_8341,N_8151);
xor U8551 (N_8551,N_8015,N_8170);
and U8552 (N_8552,N_8288,N_8344);
or U8553 (N_8553,N_8410,N_8168);
nor U8554 (N_8554,N_8465,N_8041);
nor U8555 (N_8555,N_8116,N_8395);
nand U8556 (N_8556,N_8295,N_8021);
nor U8557 (N_8557,N_8136,N_8468);
nor U8558 (N_8558,N_8079,N_8381);
nand U8559 (N_8559,N_8339,N_8086);
nand U8560 (N_8560,N_8307,N_8477);
xnor U8561 (N_8561,N_8396,N_8435);
or U8562 (N_8562,N_8306,N_8485);
xnor U8563 (N_8563,N_8259,N_8452);
xor U8564 (N_8564,N_8189,N_8117);
xnor U8565 (N_8565,N_8422,N_8109);
or U8566 (N_8566,N_8227,N_8107);
nand U8567 (N_8567,N_8206,N_8219);
or U8568 (N_8568,N_8038,N_8150);
and U8569 (N_8569,N_8205,N_8101);
or U8570 (N_8570,N_8418,N_8456);
xnor U8571 (N_8571,N_8013,N_8185);
nand U8572 (N_8572,N_8431,N_8102);
nand U8573 (N_8573,N_8143,N_8472);
and U8574 (N_8574,N_8195,N_8444);
nand U8575 (N_8575,N_8240,N_8155);
nand U8576 (N_8576,N_8005,N_8297);
nand U8577 (N_8577,N_8334,N_8095);
or U8578 (N_8578,N_8003,N_8496);
nor U8579 (N_8579,N_8176,N_8467);
and U8580 (N_8580,N_8454,N_8152);
or U8581 (N_8581,N_8296,N_8258);
nand U8582 (N_8582,N_8436,N_8180);
and U8583 (N_8583,N_8008,N_8066);
or U8584 (N_8584,N_8040,N_8330);
and U8585 (N_8585,N_8081,N_8209);
xnor U8586 (N_8586,N_8073,N_8480);
nand U8587 (N_8587,N_8045,N_8232);
nor U8588 (N_8588,N_8382,N_8080);
and U8589 (N_8589,N_8269,N_8178);
or U8590 (N_8590,N_8223,N_8397);
nor U8591 (N_8591,N_8196,N_8438);
xor U8592 (N_8592,N_8280,N_8127);
nand U8593 (N_8593,N_8129,N_8224);
and U8594 (N_8594,N_8084,N_8007);
nor U8595 (N_8595,N_8023,N_8462);
and U8596 (N_8596,N_8001,N_8247);
and U8597 (N_8597,N_8183,N_8310);
or U8598 (N_8598,N_8061,N_8144);
nor U8599 (N_8599,N_8432,N_8384);
and U8600 (N_8600,N_8451,N_8376);
nor U8601 (N_8601,N_8055,N_8278);
xnor U8602 (N_8602,N_8281,N_8377);
nand U8603 (N_8603,N_8215,N_8423);
nor U8604 (N_8604,N_8450,N_8386);
or U8605 (N_8605,N_8305,N_8257);
xnor U8606 (N_8606,N_8338,N_8494);
nor U8607 (N_8607,N_8375,N_8214);
or U8608 (N_8608,N_8320,N_8068);
nor U8609 (N_8609,N_8347,N_8199);
xor U8610 (N_8610,N_8071,N_8076);
nor U8611 (N_8611,N_8365,N_8190);
and U8612 (N_8612,N_8405,N_8235);
or U8613 (N_8613,N_8229,N_8114);
or U8614 (N_8614,N_8218,N_8163);
xnor U8615 (N_8615,N_8367,N_8208);
and U8616 (N_8616,N_8430,N_8433);
or U8617 (N_8617,N_8411,N_8085);
nor U8618 (N_8618,N_8286,N_8488);
and U8619 (N_8619,N_8192,N_8317);
nand U8620 (N_8620,N_8130,N_8239);
or U8621 (N_8621,N_8019,N_8359);
xnor U8622 (N_8622,N_8051,N_8408);
xor U8623 (N_8623,N_8323,N_8077);
or U8624 (N_8624,N_8302,N_8345);
nand U8625 (N_8625,N_8104,N_8029);
or U8626 (N_8626,N_8470,N_8251);
or U8627 (N_8627,N_8406,N_8125);
or U8628 (N_8628,N_8236,N_8274);
or U8629 (N_8629,N_8413,N_8285);
nor U8630 (N_8630,N_8440,N_8439);
xor U8631 (N_8631,N_8070,N_8234);
and U8632 (N_8632,N_8291,N_8265);
nor U8633 (N_8633,N_8146,N_8242);
or U8634 (N_8634,N_8420,N_8398);
or U8635 (N_8635,N_8187,N_8355);
and U8636 (N_8636,N_8200,N_8004);
or U8637 (N_8637,N_8449,N_8090);
xnor U8638 (N_8638,N_8429,N_8326);
nand U8639 (N_8639,N_8282,N_8464);
nor U8640 (N_8640,N_8042,N_8460);
nor U8641 (N_8641,N_8243,N_8497);
and U8642 (N_8642,N_8092,N_8194);
xnor U8643 (N_8643,N_8407,N_8476);
and U8644 (N_8644,N_8197,N_8358);
nor U8645 (N_8645,N_8222,N_8461);
nand U8646 (N_8646,N_8279,N_8063);
xnor U8647 (N_8647,N_8304,N_8391);
nor U8648 (N_8648,N_8052,N_8303);
and U8649 (N_8649,N_8360,N_8315);
xor U8650 (N_8650,N_8402,N_8373);
nor U8651 (N_8651,N_8255,N_8186);
nand U8652 (N_8652,N_8106,N_8096);
and U8653 (N_8653,N_8169,N_8142);
or U8654 (N_8654,N_8453,N_8414);
xor U8655 (N_8655,N_8443,N_8174);
xnor U8656 (N_8656,N_8412,N_8221);
nand U8657 (N_8657,N_8230,N_8324);
or U8658 (N_8658,N_8201,N_8211);
nand U8659 (N_8659,N_8446,N_8020);
xnor U8660 (N_8660,N_8348,N_8018);
xor U8661 (N_8661,N_8204,N_8448);
and U8662 (N_8662,N_8409,N_8434);
xor U8663 (N_8663,N_8120,N_8417);
or U8664 (N_8664,N_8010,N_8483);
xor U8665 (N_8665,N_8158,N_8253);
nand U8666 (N_8666,N_8322,N_8094);
xnor U8667 (N_8667,N_8340,N_8027);
nor U8668 (N_8668,N_8437,N_8137);
xor U8669 (N_8669,N_8350,N_8028);
nor U8670 (N_8670,N_8256,N_8241);
nand U8671 (N_8671,N_8110,N_8087);
xnor U8672 (N_8672,N_8193,N_8237);
nand U8673 (N_8673,N_8147,N_8011);
or U8674 (N_8674,N_8228,N_8466);
nor U8675 (N_8675,N_8016,N_8387);
or U8676 (N_8676,N_8428,N_8378);
and U8677 (N_8677,N_8366,N_8225);
and U8678 (N_8678,N_8354,N_8075);
or U8679 (N_8679,N_8290,N_8372);
xor U8680 (N_8680,N_8078,N_8475);
xnor U8681 (N_8681,N_8270,N_8049);
xnor U8682 (N_8682,N_8140,N_8046);
or U8683 (N_8683,N_8000,N_8054);
or U8684 (N_8684,N_8154,N_8069);
nand U8685 (N_8685,N_8314,N_8026);
xnor U8686 (N_8686,N_8124,N_8289);
nand U8687 (N_8687,N_8062,N_8336);
nor U8688 (N_8688,N_8442,N_8371);
xnor U8689 (N_8689,N_8495,N_8161);
nor U8690 (N_8690,N_8394,N_8141);
xnor U8691 (N_8691,N_8337,N_8249);
nand U8692 (N_8692,N_8173,N_8050);
or U8693 (N_8693,N_8006,N_8292);
and U8694 (N_8694,N_8179,N_8043);
and U8695 (N_8695,N_8478,N_8313);
and U8696 (N_8696,N_8268,N_8309);
nor U8697 (N_8697,N_8370,N_8238);
nor U8698 (N_8698,N_8059,N_8316);
nor U8699 (N_8699,N_8132,N_8293);
and U8700 (N_8700,N_8400,N_8088);
nand U8701 (N_8701,N_8056,N_8390);
nor U8702 (N_8702,N_8121,N_8333);
nor U8703 (N_8703,N_8284,N_8217);
nor U8704 (N_8704,N_8072,N_8416);
or U8705 (N_8705,N_8479,N_8089);
nor U8706 (N_8706,N_8160,N_8009);
xor U8707 (N_8707,N_8357,N_8252);
nor U8708 (N_8708,N_8031,N_8202);
xnor U8709 (N_8709,N_8369,N_8474);
and U8710 (N_8710,N_8057,N_8421);
nor U8711 (N_8711,N_8103,N_8308);
nor U8712 (N_8712,N_8039,N_8112);
and U8713 (N_8713,N_8082,N_8226);
or U8714 (N_8714,N_8153,N_8343);
nand U8715 (N_8715,N_8419,N_8032);
nor U8716 (N_8716,N_8156,N_8492);
nand U8717 (N_8717,N_8207,N_8233);
nor U8718 (N_8718,N_8159,N_8212);
nor U8719 (N_8719,N_8035,N_8148);
and U8720 (N_8720,N_8053,N_8033);
and U8721 (N_8721,N_8119,N_8036);
nand U8722 (N_8722,N_8325,N_8455);
xor U8723 (N_8723,N_8165,N_8489);
and U8724 (N_8724,N_8017,N_8276);
xor U8725 (N_8725,N_8203,N_8105);
or U8726 (N_8726,N_8099,N_8097);
nor U8727 (N_8727,N_8272,N_8210);
or U8728 (N_8728,N_8024,N_8044);
or U8729 (N_8729,N_8361,N_8245);
nand U8730 (N_8730,N_8145,N_8267);
or U8731 (N_8731,N_8074,N_8275);
or U8732 (N_8732,N_8177,N_8065);
and U8733 (N_8733,N_8128,N_8184);
xor U8734 (N_8734,N_8374,N_8491);
nand U8735 (N_8735,N_8294,N_8349);
xor U8736 (N_8736,N_8118,N_8248);
or U8737 (N_8737,N_8181,N_8424);
xor U8738 (N_8738,N_8037,N_8385);
and U8739 (N_8739,N_8362,N_8014);
nand U8740 (N_8740,N_8335,N_8182);
or U8741 (N_8741,N_8352,N_8098);
nand U8742 (N_8742,N_8319,N_8283);
nor U8743 (N_8743,N_8123,N_8134);
nand U8744 (N_8744,N_8301,N_8175);
or U8745 (N_8745,N_8157,N_8353);
and U8746 (N_8746,N_8364,N_8441);
nor U8747 (N_8747,N_8266,N_8490);
nor U8748 (N_8748,N_8254,N_8111);
and U8749 (N_8749,N_8383,N_8246);
nand U8750 (N_8750,N_8350,N_8237);
nand U8751 (N_8751,N_8400,N_8135);
and U8752 (N_8752,N_8256,N_8201);
xnor U8753 (N_8753,N_8491,N_8265);
nor U8754 (N_8754,N_8261,N_8068);
or U8755 (N_8755,N_8040,N_8052);
nand U8756 (N_8756,N_8250,N_8106);
nand U8757 (N_8757,N_8178,N_8453);
nor U8758 (N_8758,N_8043,N_8419);
xnor U8759 (N_8759,N_8301,N_8416);
xnor U8760 (N_8760,N_8208,N_8113);
nor U8761 (N_8761,N_8025,N_8407);
xor U8762 (N_8762,N_8134,N_8316);
or U8763 (N_8763,N_8066,N_8121);
nor U8764 (N_8764,N_8175,N_8309);
xnor U8765 (N_8765,N_8122,N_8203);
or U8766 (N_8766,N_8396,N_8227);
xor U8767 (N_8767,N_8424,N_8472);
nor U8768 (N_8768,N_8048,N_8427);
nor U8769 (N_8769,N_8452,N_8033);
nor U8770 (N_8770,N_8310,N_8447);
nand U8771 (N_8771,N_8049,N_8222);
xnor U8772 (N_8772,N_8332,N_8032);
xnor U8773 (N_8773,N_8087,N_8159);
nand U8774 (N_8774,N_8100,N_8106);
nor U8775 (N_8775,N_8338,N_8348);
nor U8776 (N_8776,N_8442,N_8319);
and U8777 (N_8777,N_8057,N_8193);
or U8778 (N_8778,N_8111,N_8164);
xnor U8779 (N_8779,N_8033,N_8359);
xnor U8780 (N_8780,N_8448,N_8341);
or U8781 (N_8781,N_8278,N_8469);
or U8782 (N_8782,N_8107,N_8208);
and U8783 (N_8783,N_8023,N_8011);
or U8784 (N_8784,N_8344,N_8289);
nand U8785 (N_8785,N_8051,N_8399);
nand U8786 (N_8786,N_8302,N_8185);
or U8787 (N_8787,N_8051,N_8106);
nor U8788 (N_8788,N_8142,N_8120);
nor U8789 (N_8789,N_8276,N_8216);
or U8790 (N_8790,N_8345,N_8293);
or U8791 (N_8791,N_8023,N_8169);
or U8792 (N_8792,N_8241,N_8074);
xor U8793 (N_8793,N_8192,N_8203);
and U8794 (N_8794,N_8272,N_8384);
nor U8795 (N_8795,N_8263,N_8418);
or U8796 (N_8796,N_8120,N_8380);
xor U8797 (N_8797,N_8042,N_8396);
nand U8798 (N_8798,N_8061,N_8160);
nand U8799 (N_8799,N_8356,N_8236);
or U8800 (N_8800,N_8402,N_8249);
and U8801 (N_8801,N_8329,N_8146);
nand U8802 (N_8802,N_8065,N_8248);
nor U8803 (N_8803,N_8460,N_8341);
xnor U8804 (N_8804,N_8207,N_8198);
xnor U8805 (N_8805,N_8109,N_8098);
or U8806 (N_8806,N_8481,N_8328);
or U8807 (N_8807,N_8486,N_8339);
nand U8808 (N_8808,N_8090,N_8004);
and U8809 (N_8809,N_8025,N_8026);
nor U8810 (N_8810,N_8261,N_8228);
or U8811 (N_8811,N_8067,N_8349);
xnor U8812 (N_8812,N_8307,N_8482);
and U8813 (N_8813,N_8394,N_8017);
xor U8814 (N_8814,N_8262,N_8238);
or U8815 (N_8815,N_8033,N_8338);
xor U8816 (N_8816,N_8161,N_8364);
xor U8817 (N_8817,N_8000,N_8377);
nor U8818 (N_8818,N_8355,N_8274);
and U8819 (N_8819,N_8197,N_8150);
xnor U8820 (N_8820,N_8252,N_8099);
nand U8821 (N_8821,N_8232,N_8004);
and U8822 (N_8822,N_8000,N_8046);
and U8823 (N_8823,N_8004,N_8177);
and U8824 (N_8824,N_8323,N_8326);
or U8825 (N_8825,N_8182,N_8065);
nand U8826 (N_8826,N_8221,N_8066);
nand U8827 (N_8827,N_8390,N_8204);
nor U8828 (N_8828,N_8294,N_8499);
and U8829 (N_8829,N_8485,N_8496);
xnor U8830 (N_8830,N_8153,N_8421);
and U8831 (N_8831,N_8120,N_8076);
xor U8832 (N_8832,N_8316,N_8196);
nor U8833 (N_8833,N_8139,N_8085);
nand U8834 (N_8834,N_8060,N_8110);
or U8835 (N_8835,N_8218,N_8235);
nand U8836 (N_8836,N_8145,N_8106);
xnor U8837 (N_8837,N_8429,N_8028);
xnor U8838 (N_8838,N_8019,N_8444);
xnor U8839 (N_8839,N_8223,N_8035);
or U8840 (N_8840,N_8019,N_8343);
xor U8841 (N_8841,N_8295,N_8230);
xnor U8842 (N_8842,N_8256,N_8279);
or U8843 (N_8843,N_8019,N_8426);
or U8844 (N_8844,N_8298,N_8006);
and U8845 (N_8845,N_8472,N_8304);
or U8846 (N_8846,N_8222,N_8425);
and U8847 (N_8847,N_8031,N_8495);
xor U8848 (N_8848,N_8240,N_8137);
nor U8849 (N_8849,N_8242,N_8248);
nor U8850 (N_8850,N_8164,N_8133);
nor U8851 (N_8851,N_8073,N_8251);
nor U8852 (N_8852,N_8204,N_8432);
and U8853 (N_8853,N_8495,N_8481);
or U8854 (N_8854,N_8499,N_8092);
xnor U8855 (N_8855,N_8205,N_8028);
xor U8856 (N_8856,N_8026,N_8061);
nand U8857 (N_8857,N_8292,N_8266);
nand U8858 (N_8858,N_8001,N_8495);
xor U8859 (N_8859,N_8212,N_8177);
xnor U8860 (N_8860,N_8418,N_8029);
xor U8861 (N_8861,N_8090,N_8493);
nand U8862 (N_8862,N_8450,N_8206);
nand U8863 (N_8863,N_8262,N_8495);
xor U8864 (N_8864,N_8144,N_8416);
or U8865 (N_8865,N_8204,N_8208);
nand U8866 (N_8866,N_8356,N_8165);
nor U8867 (N_8867,N_8038,N_8023);
nor U8868 (N_8868,N_8072,N_8461);
xnor U8869 (N_8869,N_8446,N_8382);
or U8870 (N_8870,N_8077,N_8446);
or U8871 (N_8871,N_8191,N_8076);
xor U8872 (N_8872,N_8041,N_8053);
nor U8873 (N_8873,N_8259,N_8078);
nand U8874 (N_8874,N_8119,N_8272);
xor U8875 (N_8875,N_8444,N_8135);
or U8876 (N_8876,N_8175,N_8294);
nand U8877 (N_8877,N_8279,N_8198);
nor U8878 (N_8878,N_8086,N_8202);
or U8879 (N_8879,N_8297,N_8062);
or U8880 (N_8880,N_8461,N_8048);
and U8881 (N_8881,N_8207,N_8403);
nor U8882 (N_8882,N_8039,N_8035);
nand U8883 (N_8883,N_8084,N_8447);
nand U8884 (N_8884,N_8304,N_8465);
and U8885 (N_8885,N_8376,N_8383);
and U8886 (N_8886,N_8308,N_8422);
nand U8887 (N_8887,N_8210,N_8039);
or U8888 (N_8888,N_8259,N_8059);
xor U8889 (N_8889,N_8472,N_8216);
nand U8890 (N_8890,N_8166,N_8137);
xnor U8891 (N_8891,N_8190,N_8329);
xnor U8892 (N_8892,N_8336,N_8396);
nor U8893 (N_8893,N_8117,N_8102);
xnor U8894 (N_8894,N_8454,N_8442);
and U8895 (N_8895,N_8370,N_8007);
nor U8896 (N_8896,N_8209,N_8321);
or U8897 (N_8897,N_8067,N_8300);
nand U8898 (N_8898,N_8423,N_8426);
nor U8899 (N_8899,N_8125,N_8175);
xor U8900 (N_8900,N_8067,N_8082);
nand U8901 (N_8901,N_8103,N_8181);
nand U8902 (N_8902,N_8261,N_8323);
and U8903 (N_8903,N_8231,N_8235);
or U8904 (N_8904,N_8028,N_8111);
or U8905 (N_8905,N_8351,N_8010);
and U8906 (N_8906,N_8475,N_8351);
xor U8907 (N_8907,N_8181,N_8374);
nor U8908 (N_8908,N_8433,N_8392);
nor U8909 (N_8909,N_8412,N_8298);
and U8910 (N_8910,N_8288,N_8272);
nand U8911 (N_8911,N_8240,N_8399);
nor U8912 (N_8912,N_8005,N_8172);
xnor U8913 (N_8913,N_8036,N_8217);
and U8914 (N_8914,N_8452,N_8042);
nand U8915 (N_8915,N_8456,N_8126);
xor U8916 (N_8916,N_8410,N_8065);
or U8917 (N_8917,N_8447,N_8452);
xnor U8918 (N_8918,N_8383,N_8105);
nand U8919 (N_8919,N_8413,N_8458);
nand U8920 (N_8920,N_8111,N_8115);
and U8921 (N_8921,N_8157,N_8008);
or U8922 (N_8922,N_8212,N_8045);
nor U8923 (N_8923,N_8076,N_8457);
and U8924 (N_8924,N_8245,N_8330);
and U8925 (N_8925,N_8033,N_8214);
xnor U8926 (N_8926,N_8051,N_8497);
xor U8927 (N_8927,N_8359,N_8340);
nor U8928 (N_8928,N_8385,N_8437);
nand U8929 (N_8929,N_8487,N_8126);
and U8930 (N_8930,N_8227,N_8452);
xor U8931 (N_8931,N_8178,N_8078);
nand U8932 (N_8932,N_8280,N_8369);
nor U8933 (N_8933,N_8423,N_8163);
xor U8934 (N_8934,N_8172,N_8301);
xor U8935 (N_8935,N_8135,N_8191);
xor U8936 (N_8936,N_8451,N_8052);
and U8937 (N_8937,N_8223,N_8295);
or U8938 (N_8938,N_8252,N_8003);
nand U8939 (N_8939,N_8045,N_8380);
nand U8940 (N_8940,N_8216,N_8245);
and U8941 (N_8941,N_8335,N_8056);
xnor U8942 (N_8942,N_8326,N_8450);
or U8943 (N_8943,N_8460,N_8464);
nand U8944 (N_8944,N_8332,N_8241);
xor U8945 (N_8945,N_8174,N_8390);
nor U8946 (N_8946,N_8354,N_8108);
nor U8947 (N_8947,N_8062,N_8038);
nor U8948 (N_8948,N_8093,N_8444);
nor U8949 (N_8949,N_8210,N_8160);
or U8950 (N_8950,N_8276,N_8035);
and U8951 (N_8951,N_8004,N_8093);
and U8952 (N_8952,N_8248,N_8359);
or U8953 (N_8953,N_8185,N_8183);
nor U8954 (N_8954,N_8367,N_8317);
or U8955 (N_8955,N_8207,N_8121);
or U8956 (N_8956,N_8243,N_8063);
nor U8957 (N_8957,N_8128,N_8271);
nand U8958 (N_8958,N_8393,N_8126);
and U8959 (N_8959,N_8475,N_8146);
nor U8960 (N_8960,N_8208,N_8062);
xor U8961 (N_8961,N_8227,N_8285);
nor U8962 (N_8962,N_8361,N_8018);
xnor U8963 (N_8963,N_8028,N_8256);
or U8964 (N_8964,N_8322,N_8428);
xnor U8965 (N_8965,N_8207,N_8320);
xnor U8966 (N_8966,N_8108,N_8202);
nand U8967 (N_8967,N_8329,N_8319);
nand U8968 (N_8968,N_8307,N_8274);
xor U8969 (N_8969,N_8226,N_8072);
or U8970 (N_8970,N_8190,N_8141);
or U8971 (N_8971,N_8025,N_8121);
or U8972 (N_8972,N_8448,N_8168);
nand U8973 (N_8973,N_8111,N_8305);
nand U8974 (N_8974,N_8064,N_8468);
nand U8975 (N_8975,N_8195,N_8451);
nor U8976 (N_8976,N_8255,N_8466);
or U8977 (N_8977,N_8082,N_8393);
or U8978 (N_8978,N_8201,N_8245);
nor U8979 (N_8979,N_8221,N_8012);
and U8980 (N_8980,N_8162,N_8026);
or U8981 (N_8981,N_8020,N_8199);
nor U8982 (N_8982,N_8316,N_8122);
nor U8983 (N_8983,N_8248,N_8058);
or U8984 (N_8984,N_8307,N_8102);
nand U8985 (N_8985,N_8246,N_8225);
or U8986 (N_8986,N_8334,N_8094);
nor U8987 (N_8987,N_8169,N_8313);
and U8988 (N_8988,N_8359,N_8175);
xnor U8989 (N_8989,N_8313,N_8397);
nor U8990 (N_8990,N_8406,N_8393);
nor U8991 (N_8991,N_8081,N_8417);
or U8992 (N_8992,N_8259,N_8273);
and U8993 (N_8993,N_8427,N_8231);
or U8994 (N_8994,N_8024,N_8164);
and U8995 (N_8995,N_8188,N_8349);
nor U8996 (N_8996,N_8136,N_8444);
and U8997 (N_8997,N_8314,N_8051);
or U8998 (N_8998,N_8332,N_8242);
xor U8999 (N_8999,N_8056,N_8401);
and U9000 (N_9000,N_8628,N_8650);
and U9001 (N_9001,N_8899,N_8838);
nand U9002 (N_9002,N_8626,N_8710);
and U9003 (N_9003,N_8961,N_8658);
xor U9004 (N_9004,N_8613,N_8602);
nor U9005 (N_9005,N_8890,N_8592);
or U9006 (N_9006,N_8660,N_8641);
nand U9007 (N_9007,N_8597,N_8981);
nor U9008 (N_9008,N_8885,N_8500);
xnor U9009 (N_9009,N_8969,N_8913);
and U9010 (N_9010,N_8857,N_8737);
xor U9011 (N_9011,N_8783,N_8933);
nand U9012 (N_9012,N_8798,N_8587);
and U9013 (N_9013,N_8951,N_8740);
or U9014 (N_9014,N_8720,N_8861);
xor U9015 (N_9015,N_8774,N_8880);
or U9016 (N_9016,N_8950,N_8759);
xor U9017 (N_9017,N_8754,N_8580);
or U9018 (N_9018,N_8905,N_8591);
nand U9019 (N_9019,N_8860,N_8878);
and U9020 (N_9020,N_8538,N_8635);
nand U9021 (N_9021,N_8788,N_8785);
and U9022 (N_9022,N_8634,N_8937);
nor U9023 (N_9023,N_8687,N_8505);
or U9024 (N_9024,N_8945,N_8817);
or U9025 (N_9025,N_8990,N_8565);
or U9026 (N_9026,N_8742,N_8988);
nand U9027 (N_9027,N_8823,N_8517);
or U9028 (N_9028,N_8924,N_8590);
and U9029 (N_9029,N_8713,N_8734);
xor U9030 (N_9030,N_8866,N_8735);
nand U9031 (N_9031,N_8901,N_8779);
and U9032 (N_9032,N_8839,N_8822);
or U9033 (N_9033,N_8697,N_8661);
xnor U9034 (N_9034,N_8757,N_8728);
xor U9035 (N_9035,N_8653,N_8691);
nor U9036 (N_9036,N_8993,N_8884);
nor U9037 (N_9037,N_8649,N_8944);
xnor U9038 (N_9038,N_8741,N_8549);
and U9039 (N_9039,N_8518,N_8540);
nand U9040 (N_9040,N_8999,N_8576);
and U9041 (N_9041,N_8927,N_8585);
xnor U9042 (N_9042,N_8868,N_8664);
and U9043 (N_9043,N_8980,N_8876);
xnor U9044 (N_9044,N_8732,N_8572);
nor U9045 (N_9045,N_8813,N_8651);
nor U9046 (N_9046,N_8588,N_8815);
or U9047 (N_9047,N_8692,N_8543);
or U9048 (N_9048,N_8546,N_8812);
nor U9049 (N_9049,N_8504,N_8535);
and U9050 (N_9050,N_8683,N_8765);
and U9051 (N_9051,N_8555,N_8943);
xnor U9052 (N_9052,N_8654,N_8589);
xor U9053 (N_9053,N_8881,N_8851);
nand U9054 (N_9054,N_8624,N_8704);
nor U9055 (N_9055,N_8766,N_8618);
xor U9056 (N_9056,N_8917,N_8608);
or U9057 (N_9057,N_8938,N_8696);
nor U9058 (N_9058,N_8841,N_8837);
or U9059 (N_9059,N_8743,N_8909);
nor U9060 (N_9060,N_8832,N_8559);
xor U9061 (N_9061,N_8579,N_8510);
xnor U9062 (N_9062,N_8786,N_8932);
nand U9063 (N_9063,N_8915,N_8895);
or U9064 (N_9064,N_8719,N_8723);
and U9065 (N_9065,N_8948,N_8685);
or U9066 (N_9066,N_8949,N_8994);
and U9067 (N_9067,N_8528,N_8897);
nand U9068 (N_9068,N_8514,N_8553);
and U9069 (N_9069,N_8908,N_8930);
nand U9070 (N_9070,N_8984,N_8600);
xnor U9071 (N_9071,N_8607,N_8573);
nand U9072 (N_9072,N_8936,N_8724);
or U9073 (N_9073,N_8680,N_8964);
or U9074 (N_9074,N_8639,N_8974);
or U9075 (N_9075,N_8700,N_8879);
nor U9076 (N_9076,N_8914,N_8819);
nand U9077 (N_9077,N_8756,N_8609);
xor U9078 (N_9078,N_8693,N_8893);
nand U9079 (N_9079,N_8707,N_8566);
xor U9080 (N_9080,N_8793,N_8637);
nor U9081 (N_9081,N_8581,N_8954);
and U9082 (N_9082,N_8663,N_8862);
or U9083 (N_9083,N_8770,N_8665);
nor U9084 (N_9084,N_8548,N_8656);
xnor U9085 (N_9085,N_8906,N_8955);
or U9086 (N_9086,N_8567,N_8551);
and U9087 (N_9087,N_8575,N_8630);
nand U9088 (N_9088,N_8708,N_8633);
nor U9089 (N_9089,N_8542,N_8869);
nor U9090 (N_9090,N_8978,N_8956);
nor U9091 (N_9091,N_8667,N_8939);
and U9092 (N_9092,N_8789,N_8775);
nand U9093 (N_9093,N_8865,N_8596);
and U9094 (N_9094,N_8797,N_8795);
xor U9095 (N_9095,N_8947,N_8843);
nor U9096 (N_9096,N_8807,N_8733);
xor U9097 (N_9097,N_8574,N_8648);
nand U9098 (N_9098,N_8725,N_8811);
or U9099 (N_9099,N_8946,N_8856);
or U9100 (N_9100,N_8896,N_8529);
nor U9101 (N_9101,N_8532,N_8738);
nor U9102 (N_9102,N_8531,N_8750);
nand U9103 (N_9103,N_8818,N_8689);
nor U9104 (N_9104,N_8631,N_8805);
and U9105 (N_9105,N_8809,N_8644);
or U9106 (N_9106,N_8627,N_8989);
and U9107 (N_9107,N_8796,N_8836);
xnor U9108 (N_9108,N_8802,N_8957);
nand U9109 (N_9109,N_8903,N_8831);
nand U9110 (N_9110,N_8564,N_8935);
or U9111 (N_9111,N_8702,N_8621);
and U9112 (N_9112,N_8675,N_8894);
and U9113 (N_9113,N_8547,N_8749);
nor U9114 (N_9114,N_8617,N_8959);
xor U9115 (N_9115,N_8717,N_8698);
nand U9116 (N_9116,N_8530,N_8769);
nor U9117 (N_9117,N_8888,N_8763);
or U9118 (N_9118,N_8558,N_8828);
and U9119 (N_9119,N_8671,N_8715);
nor U9120 (N_9120,N_8554,N_8577);
xor U9121 (N_9121,N_8891,N_8777);
xor U9122 (N_9122,N_8799,N_8810);
nor U9123 (N_9123,N_8636,N_8673);
nand U9124 (N_9124,N_8858,N_8960);
nand U9125 (N_9125,N_8545,N_8983);
and U9126 (N_9126,N_8681,N_8527);
and U9127 (N_9127,N_8595,N_8875);
xnor U9128 (N_9128,N_8982,N_8830);
and U9129 (N_9129,N_8722,N_8995);
or U9130 (N_9130,N_8712,N_8760);
or U9131 (N_9131,N_8787,N_8803);
nor U9132 (N_9132,N_8721,N_8847);
and U9133 (N_9133,N_8882,N_8963);
and U9134 (N_9134,N_8781,N_8910);
nor U9135 (N_9135,N_8561,N_8729);
or U9136 (N_9136,N_8773,N_8782);
xnor U9137 (N_9137,N_8764,N_8525);
nor U9138 (N_9138,N_8537,N_8611);
xnor U9139 (N_9139,N_8699,N_8557);
and U9140 (N_9140,N_8752,N_8616);
nor U9141 (N_9141,N_8973,N_8652);
xor U9142 (N_9142,N_8835,N_8736);
nand U9143 (N_9143,N_8790,N_8987);
xor U9144 (N_9144,N_8643,N_8968);
xnor U9145 (N_9145,N_8544,N_8501);
xnor U9146 (N_9146,N_8709,N_8521);
xor U9147 (N_9147,N_8916,N_8670);
nor U9148 (N_9148,N_8829,N_8872);
xor U9149 (N_9149,N_8694,N_8791);
nor U9150 (N_9150,N_8755,N_8747);
or U9151 (N_9151,N_8646,N_8934);
or U9152 (N_9152,N_8522,N_8864);
nor U9153 (N_9153,N_8503,N_8674);
nand U9154 (N_9154,N_8761,N_8604);
nor U9155 (N_9155,N_8966,N_8889);
nor U9156 (N_9156,N_8682,N_8727);
and U9157 (N_9157,N_8679,N_8688);
nor U9158 (N_9158,N_8971,N_8762);
xnor U9159 (N_9159,N_8768,N_8739);
or U9160 (N_9160,N_8640,N_8840);
nand U9161 (N_9161,N_8985,N_8509);
or U9162 (N_9162,N_8911,N_8827);
nand U9163 (N_9163,N_8506,N_8584);
and U9164 (N_9164,N_8582,N_8931);
nand U9165 (N_9165,N_8877,N_8751);
xnor U9166 (N_9166,N_8918,N_8842);
xnor U9167 (N_9167,N_8767,N_8508);
or U9168 (N_9168,N_8677,N_8612);
nor U9169 (N_9169,N_8672,N_8539);
xor U9170 (N_9170,N_8863,N_8655);
xnor U9171 (N_9171,N_8867,N_8808);
and U9172 (N_9172,N_8571,N_8668);
and U9173 (N_9173,N_8855,N_8512);
xnor U9174 (N_9174,N_8870,N_8887);
nor U9175 (N_9175,N_8556,N_8645);
and U9176 (N_9176,N_8620,N_8873);
nor U9177 (N_9177,N_8686,N_8507);
or U9178 (N_9178,N_8526,N_8519);
nor U9179 (N_9179,N_8684,N_8629);
xnor U9180 (N_9180,N_8524,N_8996);
or U9181 (N_9181,N_8701,N_8923);
or U9182 (N_9182,N_8711,N_8744);
or U9183 (N_9183,N_8705,N_8922);
nand U9184 (N_9184,N_8718,N_8886);
or U9185 (N_9185,N_8730,N_8850);
nand U9186 (N_9186,N_8515,N_8758);
and U9187 (N_9187,N_8902,N_8970);
nor U9188 (N_9188,N_8776,N_8562);
nor U9189 (N_9189,N_8599,N_8849);
nor U9190 (N_9190,N_8550,N_8520);
xnor U9191 (N_9191,N_8659,N_8965);
nor U9192 (N_9192,N_8975,N_8568);
or U9193 (N_9193,N_8778,N_8513);
or U9194 (N_9194,N_8666,N_8991);
and U9195 (N_9195,N_8845,N_8714);
and U9196 (N_9196,N_8610,N_8986);
xnor U9197 (N_9197,N_8690,N_8941);
or U9198 (N_9198,N_8800,N_8825);
and U9199 (N_9199,N_8919,N_8912);
xor U9200 (N_9200,N_8892,N_8598);
and U9201 (N_9201,N_8560,N_8642);
or U9202 (N_9202,N_8523,N_8962);
nand U9203 (N_9203,N_8594,N_8748);
or U9204 (N_9204,N_8615,N_8859);
nor U9205 (N_9205,N_8806,N_8907);
or U9206 (N_9206,N_8784,N_8929);
nor U9207 (N_9207,N_8801,N_8716);
nand U9208 (N_9208,N_8638,N_8623);
nand U9209 (N_9209,N_8940,N_8552);
or U9210 (N_9210,N_8904,N_8852);
xnor U9211 (N_9211,N_8921,N_8824);
and U9212 (N_9212,N_8669,N_8511);
xnor U9213 (N_9213,N_8920,N_8854);
xor U9214 (N_9214,N_8992,N_8534);
nand U9215 (N_9215,N_8972,N_8977);
and U9216 (N_9216,N_8619,N_8998);
or U9217 (N_9217,N_8578,N_8731);
and U9218 (N_9218,N_8593,N_8953);
nand U9219 (N_9219,N_8772,N_8533);
or U9220 (N_9220,N_8647,N_8952);
or U9221 (N_9221,N_8586,N_8726);
nor U9222 (N_9222,N_8898,N_8820);
or U9223 (N_9223,N_8834,N_8583);
nand U9224 (N_9224,N_8853,N_8883);
or U9225 (N_9225,N_8703,N_8605);
nand U9226 (N_9226,N_8536,N_8846);
or U9227 (N_9227,N_8614,N_8676);
nand U9228 (N_9228,N_8745,N_8826);
nor U9229 (N_9229,N_8871,N_8874);
and U9230 (N_9230,N_8606,N_8844);
or U9231 (N_9231,N_8780,N_8746);
nand U9232 (N_9232,N_8502,N_8804);
nand U9233 (N_9233,N_8814,N_8569);
nand U9234 (N_9234,N_8816,N_8833);
or U9235 (N_9235,N_8541,N_8792);
nor U9236 (N_9236,N_8570,N_8928);
or U9237 (N_9237,N_8625,N_8657);
xnor U9238 (N_9238,N_8925,N_8753);
nor U9239 (N_9239,N_8603,N_8967);
nand U9240 (N_9240,N_8958,N_8662);
nand U9241 (N_9241,N_8622,N_8926);
or U9242 (N_9242,N_8794,N_8601);
xor U9243 (N_9243,N_8942,N_8516);
or U9244 (N_9244,N_8563,N_8997);
or U9245 (N_9245,N_8976,N_8900);
nor U9246 (N_9246,N_8678,N_8632);
or U9247 (N_9247,N_8848,N_8771);
nor U9248 (N_9248,N_8706,N_8695);
xnor U9249 (N_9249,N_8979,N_8821);
or U9250 (N_9250,N_8599,N_8907);
or U9251 (N_9251,N_8932,N_8739);
or U9252 (N_9252,N_8583,N_8762);
and U9253 (N_9253,N_8684,N_8920);
or U9254 (N_9254,N_8604,N_8717);
nor U9255 (N_9255,N_8806,N_8689);
and U9256 (N_9256,N_8670,N_8982);
or U9257 (N_9257,N_8996,N_8568);
xnor U9258 (N_9258,N_8582,N_8764);
or U9259 (N_9259,N_8870,N_8578);
and U9260 (N_9260,N_8618,N_8554);
xnor U9261 (N_9261,N_8822,N_8642);
and U9262 (N_9262,N_8835,N_8656);
nand U9263 (N_9263,N_8957,N_8756);
xnor U9264 (N_9264,N_8563,N_8651);
and U9265 (N_9265,N_8548,N_8798);
xnor U9266 (N_9266,N_8967,N_8587);
and U9267 (N_9267,N_8990,N_8538);
and U9268 (N_9268,N_8926,N_8577);
nor U9269 (N_9269,N_8754,N_8766);
or U9270 (N_9270,N_8800,N_8754);
nand U9271 (N_9271,N_8888,N_8766);
or U9272 (N_9272,N_8985,N_8849);
or U9273 (N_9273,N_8901,N_8964);
nand U9274 (N_9274,N_8949,N_8890);
nor U9275 (N_9275,N_8738,N_8869);
nand U9276 (N_9276,N_8611,N_8555);
nand U9277 (N_9277,N_8799,N_8988);
nand U9278 (N_9278,N_8707,N_8792);
and U9279 (N_9279,N_8821,N_8518);
or U9280 (N_9280,N_8780,N_8946);
or U9281 (N_9281,N_8601,N_8777);
nand U9282 (N_9282,N_8969,N_8723);
nor U9283 (N_9283,N_8767,N_8573);
and U9284 (N_9284,N_8925,N_8778);
nand U9285 (N_9285,N_8840,N_8930);
xor U9286 (N_9286,N_8743,N_8628);
xor U9287 (N_9287,N_8655,N_8682);
and U9288 (N_9288,N_8847,N_8517);
or U9289 (N_9289,N_8977,N_8568);
or U9290 (N_9290,N_8548,N_8573);
nand U9291 (N_9291,N_8740,N_8865);
nand U9292 (N_9292,N_8504,N_8686);
nand U9293 (N_9293,N_8839,N_8816);
and U9294 (N_9294,N_8958,N_8700);
or U9295 (N_9295,N_8784,N_8774);
nand U9296 (N_9296,N_8911,N_8552);
nor U9297 (N_9297,N_8733,N_8732);
nand U9298 (N_9298,N_8796,N_8789);
xnor U9299 (N_9299,N_8631,N_8538);
nand U9300 (N_9300,N_8797,N_8851);
xnor U9301 (N_9301,N_8612,N_8889);
nor U9302 (N_9302,N_8867,N_8801);
or U9303 (N_9303,N_8777,N_8918);
and U9304 (N_9304,N_8938,N_8709);
nand U9305 (N_9305,N_8828,N_8768);
and U9306 (N_9306,N_8623,N_8812);
xor U9307 (N_9307,N_8642,N_8775);
xnor U9308 (N_9308,N_8504,N_8874);
or U9309 (N_9309,N_8906,N_8811);
nand U9310 (N_9310,N_8782,N_8503);
and U9311 (N_9311,N_8680,N_8717);
or U9312 (N_9312,N_8869,N_8927);
xor U9313 (N_9313,N_8537,N_8927);
and U9314 (N_9314,N_8618,N_8616);
or U9315 (N_9315,N_8713,N_8607);
xor U9316 (N_9316,N_8596,N_8676);
and U9317 (N_9317,N_8590,N_8857);
xnor U9318 (N_9318,N_8546,N_8738);
nor U9319 (N_9319,N_8573,N_8876);
nand U9320 (N_9320,N_8833,N_8743);
xnor U9321 (N_9321,N_8775,N_8735);
or U9322 (N_9322,N_8528,N_8899);
xor U9323 (N_9323,N_8811,N_8624);
nor U9324 (N_9324,N_8616,N_8802);
nand U9325 (N_9325,N_8500,N_8981);
nor U9326 (N_9326,N_8590,N_8758);
and U9327 (N_9327,N_8669,N_8872);
or U9328 (N_9328,N_8788,N_8907);
or U9329 (N_9329,N_8970,N_8651);
and U9330 (N_9330,N_8940,N_8636);
nand U9331 (N_9331,N_8807,N_8991);
nand U9332 (N_9332,N_8693,N_8790);
or U9333 (N_9333,N_8950,N_8902);
and U9334 (N_9334,N_8610,N_8740);
nand U9335 (N_9335,N_8644,N_8616);
xor U9336 (N_9336,N_8700,N_8793);
nor U9337 (N_9337,N_8789,N_8577);
and U9338 (N_9338,N_8765,N_8852);
nand U9339 (N_9339,N_8859,N_8569);
nor U9340 (N_9340,N_8771,N_8625);
nor U9341 (N_9341,N_8828,N_8603);
nor U9342 (N_9342,N_8865,N_8631);
nor U9343 (N_9343,N_8997,N_8550);
and U9344 (N_9344,N_8908,N_8901);
nor U9345 (N_9345,N_8762,N_8798);
and U9346 (N_9346,N_8753,N_8999);
nor U9347 (N_9347,N_8631,N_8582);
xor U9348 (N_9348,N_8728,N_8531);
nand U9349 (N_9349,N_8924,N_8888);
and U9350 (N_9350,N_8941,N_8664);
nor U9351 (N_9351,N_8643,N_8558);
xor U9352 (N_9352,N_8543,N_8913);
nor U9353 (N_9353,N_8766,N_8610);
xor U9354 (N_9354,N_8790,N_8704);
nor U9355 (N_9355,N_8540,N_8763);
nand U9356 (N_9356,N_8755,N_8923);
nor U9357 (N_9357,N_8796,N_8825);
nand U9358 (N_9358,N_8605,N_8763);
xor U9359 (N_9359,N_8782,N_8575);
and U9360 (N_9360,N_8883,N_8821);
or U9361 (N_9361,N_8851,N_8763);
and U9362 (N_9362,N_8762,N_8748);
and U9363 (N_9363,N_8644,N_8510);
and U9364 (N_9364,N_8991,N_8770);
or U9365 (N_9365,N_8967,N_8785);
nand U9366 (N_9366,N_8564,N_8907);
and U9367 (N_9367,N_8737,N_8946);
nor U9368 (N_9368,N_8916,N_8519);
and U9369 (N_9369,N_8806,N_8696);
and U9370 (N_9370,N_8947,N_8547);
or U9371 (N_9371,N_8660,N_8838);
and U9372 (N_9372,N_8811,N_8657);
nor U9373 (N_9373,N_8649,N_8811);
and U9374 (N_9374,N_8894,N_8591);
and U9375 (N_9375,N_8510,N_8552);
xor U9376 (N_9376,N_8684,N_8829);
or U9377 (N_9377,N_8634,N_8991);
and U9378 (N_9378,N_8916,N_8683);
xor U9379 (N_9379,N_8728,N_8905);
nor U9380 (N_9380,N_8784,N_8945);
nor U9381 (N_9381,N_8662,N_8758);
nand U9382 (N_9382,N_8532,N_8809);
xnor U9383 (N_9383,N_8905,N_8549);
and U9384 (N_9384,N_8774,N_8903);
nor U9385 (N_9385,N_8557,N_8685);
xnor U9386 (N_9386,N_8862,N_8954);
nor U9387 (N_9387,N_8716,N_8804);
or U9388 (N_9388,N_8740,N_8597);
nor U9389 (N_9389,N_8616,N_8823);
nor U9390 (N_9390,N_8886,N_8830);
xnor U9391 (N_9391,N_8862,N_8632);
nand U9392 (N_9392,N_8904,N_8683);
xor U9393 (N_9393,N_8632,N_8641);
nor U9394 (N_9394,N_8544,N_8831);
or U9395 (N_9395,N_8601,N_8630);
xor U9396 (N_9396,N_8512,N_8524);
and U9397 (N_9397,N_8611,N_8927);
nand U9398 (N_9398,N_8982,N_8587);
nor U9399 (N_9399,N_8852,N_8682);
nand U9400 (N_9400,N_8637,N_8579);
xnor U9401 (N_9401,N_8731,N_8882);
nand U9402 (N_9402,N_8975,N_8740);
and U9403 (N_9403,N_8688,N_8630);
nand U9404 (N_9404,N_8629,N_8776);
and U9405 (N_9405,N_8615,N_8848);
and U9406 (N_9406,N_8535,N_8522);
and U9407 (N_9407,N_8679,N_8643);
nor U9408 (N_9408,N_8753,N_8880);
or U9409 (N_9409,N_8845,N_8962);
and U9410 (N_9410,N_8809,N_8813);
and U9411 (N_9411,N_8609,N_8507);
nand U9412 (N_9412,N_8755,N_8507);
or U9413 (N_9413,N_8924,N_8592);
nor U9414 (N_9414,N_8503,N_8646);
nand U9415 (N_9415,N_8962,N_8865);
xor U9416 (N_9416,N_8797,N_8802);
or U9417 (N_9417,N_8639,N_8638);
and U9418 (N_9418,N_8964,N_8903);
xor U9419 (N_9419,N_8848,N_8712);
nand U9420 (N_9420,N_8670,N_8693);
xnor U9421 (N_9421,N_8761,N_8884);
xnor U9422 (N_9422,N_8594,N_8583);
nor U9423 (N_9423,N_8943,N_8540);
nand U9424 (N_9424,N_8790,N_8972);
xor U9425 (N_9425,N_8916,N_8524);
xor U9426 (N_9426,N_8707,N_8659);
or U9427 (N_9427,N_8520,N_8985);
nand U9428 (N_9428,N_8855,N_8636);
nand U9429 (N_9429,N_8765,N_8755);
xor U9430 (N_9430,N_8751,N_8519);
xnor U9431 (N_9431,N_8905,N_8615);
nor U9432 (N_9432,N_8883,N_8513);
xnor U9433 (N_9433,N_8888,N_8742);
or U9434 (N_9434,N_8617,N_8710);
nor U9435 (N_9435,N_8983,N_8850);
nand U9436 (N_9436,N_8897,N_8988);
and U9437 (N_9437,N_8976,N_8860);
and U9438 (N_9438,N_8791,N_8589);
or U9439 (N_9439,N_8588,N_8675);
or U9440 (N_9440,N_8832,N_8531);
and U9441 (N_9441,N_8824,N_8662);
xnor U9442 (N_9442,N_8938,N_8537);
or U9443 (N_9443,N_8638,N_8657);
nor U9444 (N_9444,N_8841,N_8672);
nand U9445 (N_9445,N_8664,N_8535);
and U9446 (N_9446,N_8665,N_8575);
nand U9447 (N_9447,N_8553,N_8871);
or U9448 (N_9448,N_8857,N_8796);
or U9449 (N_9449,N_8657,N_8689);
or U9450 (N_9450,N_8807,N_8680);
or U9451 (N_9451,N_8943,N_8582);
nand U9452 (N_9452,N_8904,N_8886);
xnor U9453 (N_9453,N_8810,N_8871);
and U9454 (N_9454,N_8970,N_8953);
nand U9455 (N_9455,N_8916,N_8940);
and U9456 (N_9456,N_8670,N_8806);
and U9457 (N_9457,N_8975,N_8532);
nand U9458 (N_9458,N_8760,N_8663);
nand U9459 (N_9459,N_8776,N_8823);
nand U9460 (N_9460,N_8528,N_8781);
and U9461 (N_9461,N_8832,N_8761);
and U9462 (N_9462,N_8870,N_8502);
xnor U9463 (N_9463,N_8706,N_8930);
nand U9464 (N_9464,N_8650,N_8747);
nor U9465 (N_9465,N_8801,N_8924);
nand U9466 (N_9466,N_8920,N_8923);
xor U9467 (N_9467,N_8650,N_8602);
xor U9468 (N_9468,N_8552,N_8946);
nor U9469 (N_9469,N_8677,N_8693);
nand U9470 (N_9470,N_8909,N_8934);
xor U9471 (N_9471,N_8555,N_8661);
nor U9472 (N_9472,N_8570,N_8999);
xnor U9473 (N_9473,N_8973,N_8843);
or U9474 (N_9474,N_8614,N_8796);
nand U9475 (N_9475,N_8523,N_8598);
xnor U9476 (N_9476,N_8702,N_8812);
or U9477 (N_9477,N_8902,N_8664);
nor U9478 (N_9478,N_8823,N_8683);
nor U9479 (N_9479,N_8690,N_8615);
and U9480 (N_9480,N_8579,N_8593);
xor U9481 (N_9481,N_8592,N_8942);
and U9482 (N_9482,N_8841,N_8644);
xor U9483 (N_9483,N_8757,N_8706);
and U9484 (N_9484,N_8727,N_8645);
and U9485 (N_9485,N_8846,N_8749);
or U9486 (N_9486,N_8972,N_8898);
nand U9487 (N_9487,N_8905,N_8909);
nand U9488 (N_9488,N_8723,N_8895);
or U9489 (N_9489,N_8503,N_8886);
nand U9490 (N_9490,N_8758,N_8979);
nor U9491 (N_9491,N_8841,N_8859);
or U9492 (N_9492,N_8609,N_8579);
and U9493 (N_9493,N_8708,N_8779);
or U9494 (N_9494,N_8949,N_8523);
and U9495 (N_9495,N_8561,N_8549);
or U9496 (N_9496,N_8760,N_8734);
or U9497 (N_9497,N_8741,N_8990);
nor U9498 (N_9498,N_8792,N_8939);
or U9499 (N_9499,N_8800,N_8655);
and U9500 (N_9500,N_9406,N_9013);
nand U9501 (N_9501,N_9209,N_9242);
nand U9502 (N_9502,N_9398,N_9129);
or U9503 (N_9503,N_9054,N_9462);
and U9504 (N_9504,N_9315,N_9121);
nor U9505 (N_9505,N_9080,N_9337);
nor U9506 (N_9506,N_9473,N_9085);
xor U9507 (N_9507,N_9015,N_9296);
and U9508 (N_9508,N_9231,N_9482);
and U9509 (N_9509,N_9317,N_9050);
nand U9510 (N_9510,N_9366,N_9396);
nor U9511 (N_9511,N_9443,N_9078);
and U9512 (N_9512,N_9048,N_9359);
or U9513 (N_9513,N_9348,N_9476);
and U9514 (N_9514,N_9238,N_9498);
xor U9515 (N_9515,N_9141,N_9388);
nor U9516 (N_9516,N_9481,N_9103);
and U9517 (N_9517,N_9469,N_9172);
xnor U9518 (N_9518,N_9225,N_9002);
or U9519 (N_9519,N_9422,N_9424);
and U9520 (N_9520,N_9435,N_9160);
nand U9521 (N_9521,N_9258,N_9007);
or U9522 (N_9522,N_9148,N_9426);
or U9523 (N_9523,N_9440,N_9003);
nand U9524 (N_9524,N_9299,N_9470);
and U9525 (N_9525,N_9061,N_9226);
xnor U9526 (N_9526,N_9474,N_9267);
nor U9527 (N_9527,N_9253,N_9360);
nand U9528 (N_9528,N_9112,N_9136);
xnor U9529 (N_9529,N_9222,N_9450);
xor U9530 (N_9530,N_9218,N_9309);
xor U9531 (N_9531,N_9252,N_9384);
or U9532 (N_9532,N_9284,N_9488);
nor U9533 (N_9533,N_9330,N_9117);
xor U9534 (N_9534,N_9104,N_9133);
and U9535 (N_9535,N_9162,N_9320);
nand U9536 (N_9536,N_9207,N_9261);
and U9537 (N_9537,N_9182,N_9107);
nor U9538 (N_9538,N_9217,N_9467);
xnor U9539 (N_9539,N_9028,N_9194);
nor U9540 (N_9540,N_9039,N_9446);
nor U9541 (N_9541,N_9322,N_9154);
nor U9542 (N_9542,N_9466,N_9239);
nor U9543 (N_9543,N_9205,N_9200);
nor U9544 (N_9544,N_9010,N_9202);
nor U9545 (N_9545,N_9419,N_9185);
xor U9546 (N_9546,N_9113,N_9233);
or U9547 (N_9547,N_9389,N_9471);
nand U9548 (N_9548,N_9275,N_9211);
nand U9549 (N_9549,N_9127,N_9004);
nand U9550 (N_9550,N_9180,N_9092);
nand U9551 (N_9551,N_9352,N_9118);
or U9552 (N_9552,N_9232,N_9087);
nand U9553 (N_9553,N_9431,N_9228);
and U9554 (N_9554,N_9430,N_9340);
xnor U9555 (N_9555,N_9140,N_9489);
xor U9556 (N_9556,N_9070,N_9386);
nor U9557 (N_9557,N_9434,N_9313);
nor U9558 (N_9558,N_9206,N_9302);
or U9559 (N_9559,N_9365,N_9270);
xor U9560 (N_9560,N_9197,N_9081);
or U9561 (N_9561,N_9318,N_9123);
and U9562 (N_9562,N_9094,N_9373);
xor U9563 (N_9563,N_9150,N_9495);
nand U9564 (N_9564,N_9060,N_9427);
and U9565 (N_9565,N_9083,N_9001);
nand U9566 (N_9566,N_9369,N_9246);
nor U9567 (N_9567,N_9012,N_9041);
nor U9568 (N_9568,N_9375,N_9266);
nand U9569 (N_9569,N_9114,N_9043);
and U9570 (N_9570,N_9237,N_9086);
xnor U9571 (N_9571,N_9240,N_9046);
and U9572 (N_9572,N_9174,N_9491);
or U9573 (N_9573,N_9382,N_9063);
xnor U9574 (N_9574,N_9091,N_9444);
and U9575 (N_9575,N_9356,N_9165);
and U9576 (N_9576,N_9478,N_9090);
nor U9577 (N_9577,N_9387,N_9203);
nand U9578 (N_9578,N_9137,N_9390);
and U9579 (N_9579,N_9135,N_9288);
and U9580 (N_9580,N_9184,N_9310);
xnor U9581 (N_9581,N_9022,N_9327);
and U9582 (N_9582,N_9040,N_9014);
xor U9583 (N_9583,N_9105,N_9181);
or U9584 (N_9584,N_9357,N_9000);
and U9585 (N_9585,N_9490,N_9006);
xor U9586 (N_9586,N_9005,N_9188);
nor U9587 (N_9587,N_9319,N_9407);
or U9588 (N_9588,N_9273,N_9345);
or U9589 (N_9589,N_9169,N_9416);
nand U9590 (N_9590,N_9370,N_9096);
and U9591 (N_9591,N_9032,N_9143);
nor U9592 (N_9592,N_9280,N_9047);
and U9593 (N_9593,N_9147,N_9251);
nand U9594 (N_9594,N_9248,N_9343);
nor U9595 (N_9595,N_9351,N_9264);
and U9596 (N_9596,N_9037,N_9074);
or U9597 (N_9597,N_9304,N_9215);
nand U9598 (N_9598,N_9452,N_9088);
or U9599 (N_9599,N_9325,N_9418);
xor U9600 (N_9600,N_9229,N_9475);
nor U9601 (N_9601,N_9179,N_9290);
nand U9602 (N_9602,N_9176,N_9276);
xor U9603 (N_9603,N_9234,N_9372);
xor U9604 (N_9604,N_9018,N_9235);
nor U9605 (N_9605,N_9106,N_9159);
nand U9606 (N_9606,N_9463,N_9338);
and U9607 (N_9607,N_9448,N_9298);
and U9608 (N_9608,N_9358,N_9021);
xnor U9609 (N_9609,N_9198,N_9336);
nand U9610 (N_9610,N_9259,N_9282);
nor U9611 (N_9611,N_9368,N_9189);
nor U9612 (N_9612,N_9067,N_9055);
nand U9613 (N_9613,N_9029,N_9151);
nand U9614 (N_9614,N_9454,N_9451);
and U9615 (N_9615,N_9401,N_9163);
nor U9616 (N_9616,N_9052,N_9378);
and U9617 (N_9617,N_9016,N_9095);
nor U9618 (N_9618,N_9305,N_9171);
xnor U9619 (N_9619,N_9271,N_9472);
nand U9620 (N_9620,N_9036,N_9414);
nand U9621 (N_9621,N_9494,N_9377);
xnor U9622 (N_9622,N_9277,N_9301);
xnor U9623 (N_9623,N_9241,N_9058);
nand U9624 (N_9624,N_9221,N_9256);
nor U9625 (N_9625,N_9486,N_9392);
nor U9626 (N_9626,N_9109,N_9316);
and U9627 (N_9627,N_9349,N_9247);
nor U9628 (N_9628,N_9220,N_9287);
nor U9629 (N_9629,N_9030,N_9069);
nand U9630 (N_9630,N_9193,N_9099);
nor U9631 (N_9631,N_9487,N_9158);
or U9632 (N_9632,N_9272,N_9230);
xor U9633 (N_9633,N_9329,N_9308);
xor U9634 (N_9634,N_9260,N_9149);
xnor U9635 (N_9635,N_9265,N_9101);
nand U9636 (N_9636,N_9332,N_9363);
or U9637 (N_9637,N_9017,N_9364);
xnor U9638 (N_9638,N_9497,N_9461);
or U9639 (N_9639,N_9412,N_9411);
nor U9640 (N_9640,N_9208,N_9057);
or U9641 (N_9641,N_9307,N_9331);
nand U9642 (N_9642,N_9409,N_9051);
nand U9643 (N_9643,N_9145,N_9279);
or U9644 (N_9644,N_9072,N_9367);
or U9645 (N_9645,N_9263,N_9300);
or U9646 (N_9646,N_9291,N_9084);
and U9647 (N_9647,N_9404,N_9219);
or U9648 (N_9648,N_9460,N_9415);
nor U9649 (N_9649,N_9457,N_9479);
and U9650 (N_9650,N_9429,N_9334);
xor U9651 (N_9651,N_9496,N_9045);
or U9652 (N_9652,N_9168,N_9283);
or U9653 (N_9653,N_9468,N_9437);
and U9654 (N_9654,N_9152,N_9326);
xor U9655 (N_9655,N_9328,N_9066);
and U9656 (N_9656,N_9341,N_9269);
nand U9657 (N_9657,N_9441,N_9285);
xnor U9658 (N_9658,N_9402,N_9480);
and U9659 (N_9659,N_9019,N_9049);
or U9660 (N_9660,N_9499,N_9177);
xnor U9661 (N_9661,N_9224,N_9038);
and U9662 (N_9662,N_9216,N_9214);
or U9663 (N_9663,N_9199,N_9442);
or U9664 (N_9664,N_9314,N_9459);
nor U9665 (N_9665,N_9410,N_9347);
or U9666 (N_9666,N_9161,N_9312);
xor U9667 (N_9667,N_9191,N_9223);
or U9668 (N_9668,N_9025,N_9120);
nor U9669 (N_9669,N_9183,N_9399);
nor U9670 (N_9670,N_9195,N_9131);
xnor U9671 (N_9671,N_9009,N_9027);
or U9672 (N_9672,N_9056,N_9115);
xor U9673 (N_9673,N_9249,N_9178);
nor U9674 (N_9674,N_9423,N_9380);
xnor U9675 (N_9675,N_9201,N_9295);
xnor U9676 (N_9676,N_9255,N_9428);
nor U9677 (N_9677,N_9024,N_9465);
and U9678 (N_9678,N_9125,N_9068);
or U9679 (N_9679,N_9439,N_9034);
or U9680 (N_9680,N_9035,N_9134);
or U9681 (N_9681,N_9484,N_9031);
nand U9682 (N_9682,N_9243,N_9436);
and U9683 (N_9683,N_9033,N_9371);
nor U9684 (N_9684,N_9190,N_9236);
nand U9685 (N_9685,N_9303,N_9065);
or U9686 (N_9686,N_9408,N_9458);
or U9687 (N_9687,N_9293,N_9286);
nor U9688 (N_9688,N_9342,N_9438);
nand U9689 (N_9689,N_9391,N_9324);
nor U9690 (N_9690,N_9173,N_9130);
or U9691 (N_9691,N_9076,N_9254);
xnor U9692 (N_9692,N_9355,N_9071);
nand U9693 (N_9693,N_9346,N_9379);
nand U9694 (N_9694,N_9268,N_9432);
and U9695 (N_9695,N_9311,N_9420);
and U9696 (N_9696,N_9245,N_9167);
nand U9697 (N_9697,N_9108,N_9455);
or U9698 (N_9698,N_9155,N_9492);
xnor U9699 (N_9699,N_9353,N_9212);
or U9700 (N_9700,N_9425,N_9383);
nand U9701 (N_9701,N_9321,N_9111);
nor U9702 (N_9702,N_9144,N_9153);
and U9703 (N_9703,N_9456,N_9323);
xor U9704 (N_9704,N_9175,N_9164);
and U9705 (N_9705,N_9403,N_9306);
and U9706 (N_9706,N_9292,N_9400);
nor U9707 (N_9707,N_9257,N_9335);
xor U9708 (N_9708,N_9376,N_9297);
or U9709 (N_9709,N_9350,N_9294);
and U9710 (N_9710,N_9381,N_9413);
or U9711 (N_9711,N_9250,N_9082);
and U9712 (N_9712,N_9187,N_9344);
nor U9713 (N_9713,N_9166,N_9170);
and U9714 (N_9714,N_9333,N_9075);
and U9715 (N_9715,N_9433,N_9008);
or U9716 (N_9716,N_9042,N_9062);
xor U9717 (N_9717,N_9281,N_9122);
nor U9718 (N_9718,N_9210,N_9339);
xor U9719 (N_9719,N_9102,N_9077);
or U9720 (N_9720,N_9278,N_9362);
xnor U9721 (N_9721,N_9100,N_9110);
xor U9722 (N_9722,N_9126,N_9093);
nor U9723 (N_9723,N_9089,N_9445);
xor U9724 (N_9724,N_9011,N_9196);
nand U9725 (N_9725,N_9139,N_9204);
and U9726 (N_9726,N_9213,N_9274);
xor U9727 (N_9727,N_9397,N_9421);
and U9728 (N_9728,N_9374,N_9447);
or U9729 (N_9729,N_9142,N_9156);
nand U9730 (N_9730,N_9289,N_9186);
xor U9731 (N_9731,N_9385,N_9405);
and U9732 (N_9732,N_9262,N_9079);
and U9733 (N_9733,N_9354,N_9157);
or U9734 (N_9734,N_9192,N_9485);
nor U9735 (N_9735,N_9395,N_9146);
xnor U9736 (N_9736,N_9449,N_9119);
and U9737 (N_9737,N_9124,N_9044);
xnor U9738 (N_9738,N_9464,N_9138);
or U9739 (N_9739,N_9059,N_9026);
nand U9740 (N_9740,N_9097,N_9020);
nor U9741 (N_9741,N_9132,N_9417);
xor U9742 (N_9742,N_9483,N_9023);
or U9743 (N_9743,N_9453,N_9477);
nand U9744 (N_9744,N_9116,N_9073);
xnor U9745 (N_9745,N_9053,N_9244);
nor U9746 (N_9746,N_9361,N_9393);
or U9747 (N_9747,N_9098,N_9493);
xor U9748 (N_9748,N_9128,N_9394);
nor U9749 (N_9749,N_9227,N_9064);
nand U9750 (N_9750,N_9341,N_9228);
and U9751 (N_9751,N_9170,N_9495);
nand U9752 (N_9752,N_9279,N_9170);
nor U9753 (N_9753,N_9060,N_9042);
or U9754 (N_9754,N_9463,N_9001);
nand U9755 (N_9755,N_9059,N_9135);
xnor U9756 (N_9756,N_9189,N_9449);
and U9757 (N_9757,N_9296,N_9177);
or U9758 (N_9758,N_9431,N_9135);
nor U9759 (N_9759,N_9207,N_9375);
nor U9760 (N_9760,N_9341,N_9140);
and U9761 (N_9761,N_9411,N_9159);
nand U9762 (N_9762,N_9174,N_9421);
and U9763 (N_9763,N_9090,N_9072);
nand U9764 (N_9764,N_9151,N_9394);
xnor U9765 (N_9765,N_9024,N_9363);
xor U9766 (N_9766,N_9362,N_9183);
nor U9767 (N_9767,N_9126,N_9174);
or U9768 (N_9768,N_9499,N_9049);
and U9769 (N_9769,N_9097,N_9481);
and U9770 (N_9770,N_9203,N_9157);
nand U9771 (N_9771,N_9145,N_9324);
xnor U9772 (N_9772,N_9297,N_9379);
or U9773 (N_9773,N_9210,N_9310);
nand U9774 (N_9774,N_9076,N_9222);
nor U9775 (N_9775,N_9096,N_9151);
or U9776 (N_9776,N_9490,N_9162);
nor U9777 (N_9777,N_9077,N_9017);
nand U9778 (N_9778,N_9140,N_9069);
and U9779 (N_9779,N_9048,N_9483);
nor U9780 (N_9780,N_9041,N_9350);
or U9781 (N_9781,N_9178,N_9397);
nand U9782 (N_9782,N_9479,N_9466);
xor U9783 (N_9783,N_9230,N_9465);
nand U9784 (N_9784,N_9171,N_9302);
xor U9785 (N_9785,N_9484,N_9180);
or U9786 (N_9786,N_9262,N_9139);
nor U9787 (N_9787,N_9003,N_9001);
and U9788 (N_9788,N_9310,N_9423);
xnor U9789 (N_9789,N_9301,N_9153);
or U9790 (N_9790,N_9469,N_9227);
nand U9791 (N_9791,N_9083,N_9214);
xor U9792 (N_9792,N_9370,N_9359);
xor U9793 (N_9793,N_9045,N_9409);
or U9794 (N_9794,N_9255,N_9449);
xor U9795 (N_9795,N_9197,N_9215);
or U9796 (N_9796,N_9440,N_9193);
nand U9797 (N_9797,N_9462,N_9263);
nor U9798 (N_9798,N_9201,N_9488);
or U9799 (N_9799,N_9304,N_9242);
and U9800 (N_9800,N_9199,N_9274);
nor U9801 (N_9801,N_9028,N_9296);
xnor U9802 (N_9802,N_9269,N_9230);
and U9803 (N_9803,N_9074,N_9132);
xnor U9804 (N_9804,N_9280,N_9087);
nor U9805 (N_9805,N_9315,N_9415);
and U9806 (N_9806,N_9339,N_9037);
nor U9807 (N_9807,N_9419,N_9080);
nor U9808 (N_9808,N_9473,N_9285);
nor U9809 (N_9809,N_9056,N_9014);
nor U9810 (N_9810,N_9404,N_9159);
or U9811 (N_9811,N_9403,N_9272);
xor U9812 (N_9812,N_9253,N_9218);
nor U9813 (N_9813,N_9367,N_9067);
and U9814 (N_9814,N_9344,N_9102);
nor U9815 (N_9815,N_9225,N_9422);
nor U9816 (N_9816,N_9351,N_9267);
nor U9817 (N_9817,N_9000,N_9316);
nand U9818 (N_9818,N_9204,N_9000);
and U9819 (N_9819,N_9305,N_9005);
nor U9820 (N_9820,N_9347,N_9083);
and U9821 (N_9821,N_9487,N_9219);
xnor U9822 (N_9822,N_9223,N_9037);
or U9823 (N_9823,N_9196,N_9093);
or U9824 (N_9824,N_9127,N_9468);
and U9825 (N_9825,N_9036,N_9180);
xor U9826 (N_9826,N_9269,N_9310);
nand U9827 (N_9827,N_9162,N_9475);
xor U9828 (N_9828,N_9436,N_9249);
and U9829 (N_9829,N_9363,N_9012);
xnor U9830 (N_9830,N_9364,N_9285);
and U9831 (N_9831,N_9095,N_9226);
or U9832 (N_9832,N_9404,N_9033);
nand U9833 (N_9833,N_9363,N_9329);
xor U9834 (N_9834,N_9045,N_9012);
and U9835 (N_9835,N_9400,N_9319);
nor U9836 (N_9836,N_9419,N_9047);
and U9837 (N_9837,N_9177,N_9089);
nand U9838 (N_9838,N_9253,N_9493);
nor U9839 (N_9839,N_9044,N_9133);
and U9840 (N_9840,N_9195,N_9221);
nor U9841 (N_9841,N_9357,N_9180);
xor U9842 (N_9842,N_9468,N_9394);
or U9843 (N_9843,N_9241,N_9062);
nand U9844 (N_9844,N_9220,N_9257);
and U9845 (N_9845,N_9234,N_9473);
xnor U9846 (N_9846,N_9329,N_9333);
nand U9847 (N_9847,N_9179,N_9005);
and U9848 (N_9848,N_9462,N_9439);
nand U9849 (N_9849,N_9360,N_9230);
nand U9850 (N_9850,N_9346,N_9222);
or U9851 (N_9851,N_9434,N_9089);
xor U9852 (N_9852,N_9308,N_9434);
xnor U9853 (N_9853,N_9402,N_9354);
or U9854 (N_9854,N_9370,N_9405);
nand U9855 (N_9855,N_9362,N_9491);
xnor U9856 (N_9856,N_9030,N_9303);
xor U9857 (N_9857,N_9121,N_9112);
xnor U9858 (N_9858,N_9437,N_9446);
xnor U9859 (N_9859,N_9017,N_9454);
nor U9860 (N_9860,N_9452,N_9472);
nand U9861 (N_9861,N_9087,N_9402);
nor U9862 (N_9862,N_9446,N_9426);
and U9863 (N_9863,N_9315,N_9077);
nor U9864 (N_9864,N_9234,N_9394);
nor U9865 (N_9865,N_9380,N_9348);
and U9866 (N_9866,N_9135,N_9151);
xnor U9867 (N_9867,N_9381,N_9437);
or U9868 (N_9868,N_9063,N_9491);
or U9869 (N_9869,N_9315,N_9336);
and U9870 (N_9870,N_9249,N_9420);
nor U9871 (N_9871,N_9192,N_9307);
and U9872 (N_9872,N_9126,N_9306);
nor U9873 (N_9873,N_9407,N_9402);
or U9874 (N_9874,N_9295,N_9411);
nor U9875 (N_9875,N_9318,N_9250);
nor U9876 (N_9876,N_9336,N_9065);
xor U9877 (N_9877,N_9130,N_9351);
nor U9878 (N_9878,N_9039,N_9225);
nor U9879 (N_9879,N_9196,N_9294);
or U9880 (N_9880,N_9241,N_9289);
and U9881 (N_9881,N_9087,N_9494);
nand U9882 (N_9882,N_9033,N_9138);
and U9883 (N_9883,N_9071,N_9019);
nand U9884 (N_9884,N_9104,N_9355);
xnor U9885 (N_9885,N_9032,N_9157);
and U9886 (N_9886,N_9483,N_9392);
xor U9887 (N_9887,N_9290,N_9314);
or U9888 (N_9888,N_9258,N_9411);
and U9889 (N_9889,N_9437,N_9187);
xor U9890 (N_9890,N_9072,N_9172);
and U9891 (N_9891,N_9338,N_9308);
nor U9892 (N_9892,N_9181,N_9445);
nor U9893 (N_9893,N_9101,N_9373);
and U9894 (N_9894,N_9438,N_9351);
nand U9895 (N_9895,N_9212,N_9222);
xor U9896 (N_9896,N_9068,N_9434);
nand U9897 (N_9897,N_9269,N_9189);
or U9898 (N_9898,N_9180,N_9179);
or U9899 (N_9899,N_9436,N_9164);
xor U9900 (N_9900,N_9197,N_9086);
nor U9901 (N_9901,N_9479,N_9117);
and U9902 (N_9902,N_9350,N_9413);
nand U9903 (N_9903,N_9016,N_9022);
and U9904 (N_9904,N_9101,N_9222);
nor U9905 (N_9905,N_9044,N_9276);
nor U9906 (N_9906,N_9358,N_9012);
xnor U9907 (N_9907,N_9381,N_9161);
xnor U9908 (N_9908,N_9272,N_9325);
and U9909 (N_9909,N_9287,N_9462);
and U9910 (N_9910,N_9386,N_9345);
and U9911 (N_9911,N_9291,N_9365);
xor U9912 (N_9912,N_9180,N_9132);
or U9913 (N_9913,N_9464,N_9228);
xor U9914 (N_9914,N_9175,N_9320);
xor U9915 (N_9915,N_9105,N_9459);
xnor U9916 (N_9916,N_9190,N_9029);
or U9917 (N_9917,N_9106,N_9386);
xnor U9918 (N_9918,N_9084,N_9365);
or U9919 (N_9919,N_9004,N_9477);
nand U9920 (N_9920,N_9356,N_9487);
xor U9921 (N_9921,N_9497,N_9436);
nor U9922 (N_9922,N_9164,N_9272);
and U9923 (N_9923,N_9063,N_9233);
nor U9924 (N_9924,N_9314,N_9108);
and U9925 (N_9925,N_9063,N_9164);
and U9926 (N_9926,N_9055,N_9407);
and U9927 (N_9927,N_9160,N_9222);
nand U9928 (N_9928,N_9091,N_9005);
or U9929 (N_9929,N_9155,N_9438);
and U9930 (N_9930,N_9005,N_9147);
and U9931 (N_9931,N_9303,N_9140);
or U9932 (N_9932,N_9413,N_9310);
nor U9933 (N_9933,N_9032,N_9218);
or U9934 (N_9934,N_9191,N_9099);
nand U9935 (N_9935,N_9282,N_9088);
and U9936 (N_9936,N_9342,N_9220);
nor U9937 (N_9937,N_9416,N_9239);
nor U9938 (N_9938,N_9118,N_9268);
xor U9939 (N_9939,N_9328,N_9194);
xor U9940 (N_9940,N_9232,N_9432);
and U9941 (N_9941,N_9433,N_9259);
or U9942 (N_9942,N_9371,N_9171);
nand U9943 (N_9943,N_9042,N_9367);
xor U9944 (N_9944,N_9373,N_9068);
nor U9945 (N_9945,N_9013,N_9443);
xor U9946 (N_9946,N_9064,N_9229);
nor U9947 (N_9947,N_9300,N_9363);
nor U9948 (N_9948,N_9406,N_9392);
xor U9949 (N_9949,N_9026,N_9244);
or U9950 (N_9950,N_9299,N_9359);
or U9951 (N_9951,N_9334,N_9296);
nor U9952 (N_9952,N_9162,N_9398);
xnor U9953 (N_9953,N_9409,N_9482);
or U9954 (N_9954,N_9426,N_9233);
nor U9955 (N_9955,N_9291,N_9349);
and U9956 (N_9956,N_9155,N_9015);
nand U9957 (N_9957,N_9371,N_9117);
xor U9958 (N_9958,N_9022,N_9454);
or U9959 (N_9959,N_9478,N_9094);
nand U9960 (N_9960,N_9444,N_9112);
xnor U9961 (N_9961,N_9135,N_9001);
nand U9962 (N_9962,N_9218,N_9439);
and U9963 (N_9963,N_9331,N_9012);
nor U9964 (N_9964,N_9273,N_9344);
or U9965 (N_9965,N_9168,N_9025);
nor U9966 (N_9966,N_9342,N_9335);
nand U9967 (N_9967,N_9499,N_9285);
and U9968 (N_9968,N_9252,N_9055);
nor U9969 (N_9969,N_9015,N_9346);
nor U9970 (N_9970,N_9477,N_9350);
nand U9971 (N_9971,N_9392,N_9154);
nor U9972 (N_9972,N_9379,N_9255);
nor U9973 (N_9973,N_9074,N_9485);
or U9974 (N_9974,N_9028,N_9236);
nand U9975 (N_9975,N_9429,N_9016);
nand U9976 (N_9976,N_9068,N_9414);
and U9977 (N_9977,N_9365,N_9034);
and U9978 (N_9978,N_9054,N_9324);
or U9979 (N_9979,N_9373,N_9474);
or U9980 (N_9980,N_9039,N_9227);
xor U9981 (N_9981,N_9225,N_9008);
xor U9982 (N_9982,N_9298,N_9499);
and U9983 (N_9983,N_9247,N_9167);
and U9984 (N_9984,N_9288,N_9342);
xnor U9985 (N_9985,N_9129,N_9460);
or U9986 (N_9986,N_9246,N_9121);
or U9987 (N_9987,N_9259,N_9087);
nand U9988 (N_9988,N_9038,N_9014);
or U9989 (N_9989,N_9394,N_9018);
nor U9990 (N_9990,N_9319,N_9443);
xnor U9991 (N_9991,N_9103,N_9051);
xnor U9992 (N_9992,N_9251,N_9450);
xnor U9993 (N_9993,N_9491,N_9059);
or U9994 (N_9994,N_9025,N_9059);
nand U9995 (N_9995,N_9204,N_9010);
and U9996 (N_9996,N_9143,N_9337);
nand U9997 (N_9997,N_9185,N_9107);
nor U9998 (N_9998,N_9435,N_9380);
xnor U9999 (N_9999,N_9099,N_9117);
or UO_0 (O_0,N_9598,N_9959);
nor UO_1 (O_1,N_9907,N_9679);
nand UO_2 (O_2,N_9800,N_9678);
nor UO_3 (O_3,N_9542,N_9975);
and UO_4 (O_4,N_9763,N_9563);
nor UO_5 (O_5,N_9577,N_9881);
nor UO_6 (O_6,N_9627,N_9568);
or UO_7 (O_7,N_9602,N_9761);
nor UO_8 (O_8,N_9701,N_9523);
or UO_9 (O_9,N_9788,N_9847);
or UO_10 (O_10,N_9873,N_9978);
or UO_11 (O_11,N_9738,N_9795);
and UO_12 (O_12,N_9977,N_9583);
nor UO_13 (O_13,N_9629,N_9833);
nor UO_14 (O_14,N_9700,N_9768);
nand UO_15 (O_15,N_9826,N_9698);
nor UO_16 (O_16,N_9606,N_9658);
or UO_17 (O_17,N_9500,N_9814);
and UO_18 (O_18,N_9965,N_9643);
or UO_19 (O_19,N_9601,N_9612);
and UO_20 (O_20,N_9920,N_9727);
xnor UO_21 (O_21,N_9773,N_9995);
nor UO_22 (O_22,N_9515,N_9501);
nand UO_23 (O_23,N_9840,N_9807);
or UO_24 (O_24,N_9575,N_9589);
and UO_25 (O_25,N_9597,N_9869);
and UO_26 (O_26,N_9534,N_9675);
xnor UO_27 (O_27,N_9518,N_9691);
and UO_28 (O_28,N_9699,N_9633);
nor UO_29 (O_29,N_9586,N_9513);
and UO_30 (O_30,N_9981,N_9536);
xor UO_31 (O_31,N_9646,N_9935);
xor UO_32 (O_32,N_9966,N_9637);
or UO_33 (O_33,N_9539,N_9685);
nand UO_34 (O_34,N_9593,N_9968);
nand UO_35 (O_35,N_9852,N_9744);
or UO_36 (O_36,N_9745,N_9916);
and UO_37 (O_37,N_9882,N_9546);
nor UO_38 (O_38,N_9532,N_9838);
or UO_39 (O_39,N_9922,N_9724);
xnor UO_40 (O_40,N_9541,N_9723);
xnor UO_41 (O_41,N_9799,N_9780);
nand UO_42 (O_42,N_9998,N_9816);
and UO_43 (O_43,N_9704,N_9789);
xnor UO_44 (O_44,N_9991,N_9710);
or UO_45 (O_45,N_9645,N_9504);
and UO_46 (O_46,N_9734,N_9828);
or UO_47 (O_47,N_9638,N_9730);
nor UO_48 (O_48,N_9844,N_9621);
nor UO_49 (O_49,N_9617,N_9867);
xnor UO_50 (O_50,N_9615,N_9819);
and UO_51 (O_51,N_9599,N_9692);
nand UO_52 (O_52,N_9958,N_9930);
or UO_53 (O_53,N_9857,N_9798);
or UO_54 (O_54,N_9535,N_9822);
nand UO_55 (O_55,N_9879,N_9951);
nor UO_56 (O_56,N_9683,N_9905);
and UO_57 (O_57,N_9506,N_9717);
nor UO_58 (O_58,N_9581,N_9817);
nand UO_59 (O_59,N_9859,N_9558);
nand UO_60 (O_60,N_9676,N_9642);
and UO_61 (O_61,N_9861,N_9823);
or UO_62 (O_62,N_9886,N_9618);
nor UO_63 (O_63,N_9524,N_9839);
nand UO_64 (O_64,N_9554,N_9936);
and UO_65 (O_65,N_9845,N_9543);
and UO_66 (O_66,N_9754,N_9674);
nor UO_67 (O_67,N_9806,N_9737);
nor UO_68 (O_68,N_9555,N_9655);
xnor UO_69 (O_69,N_9887,N_9703);
and UO_70 (O_70,N_9830,N_9739);
and UO_71 (O_71,N_9640,N_9862);
and UO_72 (O_72,N_9808,N_9897);
and UO_73 (O_73,N_9585,N_9866);
or UO_74 (O_74,N_9749,N_9853);
and UO_75 (O_75,N_9711,N_9996);
or UO_76 (O_76,N_9588,N_9697);
or UO_77 (O_77,N_9979,N_9782);
or UO_78 (O_78,N_9664,N_9502);
or UO_79 (O_79,N_9911,N_9596);
nand UO_80 (O_80,N_9970,N_9791);
nand UO_81 (O_81,N_9982,N_9986);
nor UO_82 (O_82,N_9553,N_9707);
nor UO_83 (O_83,N_9573,N_9760);
nor UO_84 (O_84,N_9537,N_9915);
or UO_85 (O_85,N_9651,N_9579);
nand UO_86 (O_86,N_9630,N_9824);
xor UO_87 (O_87,N_9669,N_9976);
nand UO_88 (O_88,N_9639,N_9559);
and UO_89 (O_89,N_9894,N_9946);
and UO_90 (O_90,N_9993,N_9530);
nand UO_91 (O_91,N_9973,N_9756);
and UO_92 (O_92,N_9706,N_9628);
nor UO_93 (O_93,N_9681,N_9731);
xor UO_94 (O_94,N_9927,N_9941);
or UO_95 (O_95,N_9516,N_9777);
or UO_96 (O_96,N_9810,N_9925);
xnor UO_97 (O_97,N_9784,N_9942);
nor UO_98 (O_98,N_9713,N_9752);
nor UO_99 (O_99,N_9693,N_9619);
nand UO_100 (O_100,N_9963,N_9868);
and UO_101 (O_101,N_9871,N_9770);
and UO_102 (O_102,N_9665,N_9906);
and UO_103 (O_103,N_9755,N_9758);
and UO_104 (O_104,N_9885,N_9902);
nand UO_105 (O_105,N_9688,N_9514);
nand UO_106 (O_106,N_9635,N_9801);
and UO_107 (O_107,N_9549,N_9551);
xnor UO_108 (O_108,N_9714,N_9631);
nand UO_109 (O_109,N_9552,N_9953);
nand UO_110 (O_110,N_9748,N_9570);
and UO_111 (O_111,N_9964,N_9636);
nor UO_112 (O_112,N_9736,N_9608);
or UO_113 (O_113,N_9985,N_9781);
and UO_114 (O_114,N_9997,N_9815);
nand UO_115 (O_115,N_9662,N_9827);
and UO_116 (O_116,N_9896,N_9945);
nor UO_117 (O_117,N_9876,N_9569);
or UO_118 (O_118,N_9743,N_9939);
nand UO_119 (O_119,N_9813,N_9811);
xnor UO_120 (O_120,N_9891,N_9609);
nand UO_121 (O_121,N_9863,N_9910);
xor UO_122 (O_122,N_9783,N_9929);
nand UO_123 (O_123,N_9955,N_9895);
nor UO_124 (O_124,N_9820,N_9695);
nor UO_125 (O_125,N_9557,N_9931);
nor UO_126 (O_126,N_9888,N_9898);
and UO_127 (O_127,N_9509,N_9948);
xor UO_128 (O_128,N_9903,N_9874);
and UO_129 (O_129,N_9846,N_9538);
or UO_130 (O_130,N_9767,N_9666);
or UO_131 (O_131,N_9503,N_9521);
xor UO_132 (O_132,N_9528,N_9550);
and UO_133 (O_133,N_9605,N_9769);
xnor UO_134 (O_134,N_9864,N_9992);
or UO_135 (O_135,N_9582,N_9607);
xnor UO_136 (O_136,N_9893,N_9989);
or UO_137 (O_137,N_9843,N_9620);
nand UO_138 (O_138,N_9900,N_9590);
nor UO_139 (O_139,N_9829,N_9591);
and UO_140 (O_140,N_9511,N_9746);
xnor UO_141 (O_141,N_9994,N_9841);
or UO_142 (O_142,N_9741,N_9682);
or UO_143 (O_143,N_9933,N_9860);
and UO_144 (O_144,N_9821,N_9574);
xor UO_145 (O_145,N_9614,N_9956);
nor UO_146 (O_146,N_9786,N_9842);
or UO_147 (O_147,N_9519,N_9556);
and UO_148 (O_148,N_9694,N_9547);
nor UO_149 (O_149,N_9753,N_9854);
xor UO_150 (O_150,N_9880,N_9856);
or UO_151 (O_151,N_9751,N_9580);
nor UO_152 (O_152,N_9778,N_9878);
and UO_153 (O_153,N_9677,N_9671);
or UO_154 (O_154,N_9600,N_9571);
nand UO_155 (O_155,N_9926,N_9766);
and UO_156 (O_156,N_9949,N_9604);
nand UO_157 (O_157,N_9572,N_9947);
nor UO_158 (O_158,N_9520,N_9690);
or UO_159 (O_159,N_9790,N_9765);
and UO_160 (O_160,N_9625,N_9718);
and UO_161 (O_161,N_9603,N_9937);
nand UO_162 (O_162,N_9984,N_9566);
nand UO_163 (O_163,N_9648,N_9702);
nor UO_164 (O_164,N_9708,N_9952);
or UO_165 (O_165,N_9923,N_9709);
nor UO_166 (O_166,N_9527,N_9510);
xnor UO_167 (O_167,N_9884,N_9892);
or UO_168 (O_168,N_9657,N_9507);
xnor UO_169 (O_169,N_9687,N_9774);
and UO_170 (O_170,N_9670,N_9576);
xnor UO_171 (O_171,N_9747,N_9735);
nand UO_172 (O_172,N_9680,N_9684);
or UO_173 (O_173,N_9632,N_9792);
and UO_174 (O_174,N_9890,N_9613);
xnor UO_175 (O_175,N_9668,N_9624);
and UO_176 (O_176,N_9517,N_9720);
and UO_177 (O_177,N_9961,N_9587);
or UO_178 (O_178,N_9921,N_9851);
nand UO_179 (O_179,N_9661,N_9850);
and UO_180 (O_180,N_9940,N_9913);
nand UO_181 (O_181,N_9875,N_9831);
nand UO_182 (O_182,N_9653,N_9525);
xor UO_183 (O_183,N_9721,N_9794);
xnor UO_184 (O_184,N_9872,N_9729);
nor UO_185 (O_185,N_9865,N_9899);
nand UO_186 (O_186,N_9610,N_9855);
and UO_187 (O_187,N_9889,N_9972);
or UO_188 (O_188,N_9787,N_9740);
nand UO_189 (O_189,N_9932,N_9505);
nor UO_190 (O_190,N_9650,N_9595);
or UO_191 (O_191,N_9522,N_9967);
xnor UO_192 (O_192,N_9987,N_9649);
nand UO_193 (O_193,N_9712,N_9512);
nand UO_194 (O_194,N_9689,N_9641);
and UO_195 (O_195,N_9759,N_9834);
and UO_196 (O_196,N_9531,N_9943);
or UO_197 (O_197,N_9654,N_9848);
nand UO_198 (O_198,N_9849,N_9934);
nor UO_199 (O_199,N_9835,N_9918);
or UO_200 (O_200,N_9914,N_9944);
nor UO_201 (O_201,N_9858,N_9924);
xnor UO_202 (O_202,N_9797,N_9622);
and UO_203 (O_203,N_9673,N_9950);
xnor UO_204 (O_204,N_9954,N_9647);
nor UO_205 (O_205,N_9545,N_9544);
or UO_206 (O_206,N_9508,N_9726);
xnor UO_207 (O_207,N_9732,N_9974);
nor UO_208 (O_208,N_9971,N_9686);
and UO_209 (O_209,N_9832,N_9812);
nor UO_210 (O_210,N_9796,N_9526);
nand UO_211 (O_211,N_9771,N_9870);
nor UO_212 (O_212,N_9805,N_9990);
xnor UO_213 (O_213,N_9750,N_9928);
and UO_214 (O_214,N_9663,N_9779);
nor UO_215 (O_215,N_9656,N_9623);
xnor UO_216 (O_216,N_9764,N_9567);
xnor UO_217 (O_217,N_9909,N_9584);
nor UO_218 (O_218,N_9659,N_9616);
nand UO_219 (O_219,N_9626,N_9728);
and UO_220 (O_220,N_9938,N_9917);
xnor UO_221 (O_221,N_9548,N_9592);
nand UO_222 (O_222,N_9705,N_9912);
nor UO_223 (O_223,N_9804,N_9776);
xnor UO_224 (O_224,N_9672,N_9561);
nand UO_225 (O_225,N_9660,N_9634);
nor UO_226 (O_226,N_9565,N_9652);
nor UO_227 (O_227,N_9696,N_9733);
nand UO_228 (O_228,N_9901,N_9809);
and UO_229 (O_229,N_9594,N_9962);
nand UO_230 (O_230,N_9611,N_9540);
nor UO_231 (O_231,N_9919,N_9980);
xor UO_232 (O_232,N_9757,N_9722);
and UO_233 (O_233,N_9742,N_9715);
xor UO_234 (O_234,N_9825,N_9560);
xor UO_235 (O_235,N_9877,N_9969);
nand UO_236 (O_236,N_9564,N_9772);
or UO_237 (O_237,N_9988,N_9802);
nor UO_238 (O_238,N_9667,N_9725);
and UO_239 (O_239,N_9803,N_9883);
xnor UO_240 (O_240,N_9644,N_9818);
xnor UO_241 (O_241,N_9762,N_9904);
and UO_242 (O_242,N_9529,N_9562);
nand UO_243 (O_243,N_9578,N_9957);
and UO_244 (O_244,N_9775,N_9837);
xor UO_245 (O_245,N_9983,N_9908);
nand UO_246 (O_246,N_9960,N_9719);
nand UO_247 (O_247,N_9793,N_9785);
xor UO_248 (O_248,N_9716,N_9999);
nand UO_249 (O_249,N_9836,N_9533);
and UO_250 (O_250,N_9608,N_9713);
nor UO_251 (O_251,N_9731,N_9842);
or UO_252 (O_252,N_9992,N_9684);
and UO_253 (O_253,N_9837,N_9868);
xnor UO_254 (O_254,N_9699,N_9984);
or UO_255 (O_255,N_9847,N_9961);
nor UO_256 (O_256,N_9681,N_9899);
or UO_257 (O_257,N_9639,N_9974);
and UO_258 (O_258,N_9897,N_9510);
and UO_259 (O_259,N_9823,N_9597);
nor UO_260 (O_260,N_9648,N_9507);
or UO_261 (O_261,N_9764,N_9601);
or UO_262 (O_262,N_9776,N_9947);
nor UO_263 (O_263,N_9903,N_9511);
nand UO_264 (O_264,N_9924,N_9591);
and UO_265 (O_265,N_9887,N_9524);
nand UO_266 (O_266,N_9806,N_9634);
or UO_267 (O_267,N_9865,N_9965);
nor UO_268 (O_268,N_9832,N_9822);
nand UO_269 (O_269,N_9820,N_9598);
nor UO_270 (O_270,N_9505,N_9548);
or UO_271 (O_271,N_9797,N_9828);
xor UO_272 (O_272,N_9814,N_9926);
nor UO_273 (O_273,N_9696,N_9888);
nor UO_274 (O_274,N_9691,N_9508);
or UO_275 (O_275,N_9844,N_9551);
or UO_276 (O_276,N_9729,N_9998);
and UO_277 (O_277,N_9749,N_9612);
and UO_278 (O_278,N_9577,N_9615);
xor UO_279 (O_279,N_9820,N_9857);
nand UO_280 (O_280,N_9728,N_9939);
or UO_281 (O_281,N_9986,N_9834);
nor UO_282 (O_282,N_9892,N_9868);
nor UO_283 (O_283,N_9836,N_9933);
and UO_284 (O_284,N_9750,N_9543);
and UO_285 (O_285,N_9627,N_9657);
nor UO_286 (O_286,N_9879,N_9674);
nor UO_287 (O_287,N_9597,N_9588);
nand UO_288 (O_288,N_9962,N_9518);
and UO_289 (O_289,N_9903,N_9940);
and UO_290 (O_290,N_9962,N_9990);
nor UO_291 (O_291,N_9789,N_9696);
nor UO_292 (O_292,N_9852,N_9502);
nand UO_293 (O_293,N_9888,N_9637);
nor UO_294 (O_294,N_9816,N_9551);
xor UO_295 (O_295,N_9544,N_9638);
or UO_296 (O_296,N_9617,N_9866);
nand UO_297 (O_297,N_9626,N_9768);
nand UO_298 (O_298,N_9676,N_9645);
and UO_299 (O_299,N_9978,N_9759);
nor UO_300 (O_300,N_9982,N_9980);
nor UO_301 (O_301,N_9769,N_9888);
nand UO_302 (O_302,N_9553,N_9907);
nand UO_303 (O_303,N_9898,N_9829);
and UO_304 (O_304,N_9792,N_9978);
nor UO_305 (O_305,N_9502,N_9913);
nand UO_306 (O_306,N_9866,N_9516);
xor UO_307 (O_307,N_9974,N_9936);
nand UO_308 (O_308,N_9736,N_9710);
or UO_309 (O_309,N_9671,N_9891);
or UO_310 (O_310,N_9501,N_9659);
nand UO_311 (O_311,N_9961,N_9644);
xnor UO_312 (O_312,N_9802,N_9627);
nor UO_313 (O_313,N_9608,N_9882);
nor UO_314 (O_314,N_9804,N_9981);
xor UO_315 (O_315,N_9849,N_9992);
nand UO_316 (O_316,N_9937,N_9901);
or UO_317 (O_317,N_9892,N_9930);
nand UO_318 (O_318,N_9570,N_9862);
and UO_319 (O_319,N_9768,N_9814);
nand UO_320 (O_320,N_9529,N_9856);
and UO_321 (O_321,N_9897,N_9634);
nor UO_322 (O_322,N_9899,N_9567);
and UO_323 (O_323,N_9951,N_9516);
nor UO_324 (O_324,N_9608,N_9743);
and UO_325 (O_325,N_9849,N_9936);
and UO_326 (O_326,N_9673,N_9585);
and UO_327 (O_327,N_9541,N_9737);
or UO_328 (O_328,N_9598,N_9728);
or UO_329 (O_329,N_9979,N_9846);
nand UO_330 (O_330,N_9511,N_9663);
or UO_331 (O_331,N_9875,N_9824);
and UO_332 (O_332,N_9858,N_9551);
nor UO_333 (O_333,N_9835,N_9538);
nand UO_334 (O_334,N_9621,N_9885);
nand UO_335 (O_335,N_9974,N_9834);
nor UO_336 (O_336,N_9996,N_9937);
nor UO_337 (O_337,N_9719,N_9503);
xor UO_338 (O_338,N_9933,N_9764);
and UO_339 (O_339,N_9525,N_9527);
nor UO_340 (O_340,N_9949,N_9620);
nor UO_341 (O_341,N_9895,N_9657);
and UO_342 (O_342,N_9828,N_9532);
nor UO_343 (O_343,N_9506,N_9669);
nor UO_344 (O_344,N_9678,N_9594);
nor UO_345 (O_345,N_9841,N_9549);
or UO_346 (O_346,N_9902,N_9981);
nor UO_347 (O_347,N_9930,N_9624);
or UO_348 (O_348,N_9722,N_9789);
nor UO_349 (O_349,N_9923,N_9950);
and UO_350 (O_350,N_9587,N_9774);
nor UO_351 (O_351,N_9938,N_9541);
nand UO_352 (O_352,N_9575,N_9993);
nor UO_353 (O_353,N_9704,N_9637);
nor UO_354 (O_354,N_9623,N_9570);
or UO_355 (O_355,N_9606,N_9785);
nand UO_356 (O_356,N_9719,N_9765);
and UO_357 (O_357,N_9554,N_9611);
and UO_358 (O_358,N_9536,N_9839);
nand UO_359 (O_359,N_9875,N_9775);
nand UO_360 (O_360,N_9665,N_9913);
xor UO_361 (O_361,N_9857,N_9689);
nor UO_362 (O_362,N_9996,N_9890);
and UO_363 (O_363,N_9629,N_9834);
and UO_364 (O_364,N_9629,N_9520);
or UO_365 (O_365,N_9755,N_9999);
nor UO_366 (O_366,N_9546,N_9769);
nor UO_367 (O_367,N_9748,N_9721);
nor UO_368 (O_368,N_9902,N_9953);
xnor UO_369 (O_369,N_9826,N_9876);
and UO_370 (O_370,N_9881,N_9806);
xnor UO_371 (O_371,N_9552,N_9743);
nand UO_372 (O_372,N_9648,N_9638);
and UO_373 (O_373,N_9769,N_9970);
nand UO_374 (O_374,N_9507,N_9505);
or UO_375 (O_375,N_9553,N_9719);
and UO_376 (O_376,N_9638,N_9598);
xor UO_377 (O_377,N_9521,N_9742);
nand UO_378 (O_378,N_9963,N_9579);
nor UO_379 (O_379,N_9951,N_9992);
nand UO_380 (O_380,N_9665,N_9639);
and UO_381 (O_381,N_9515,N_9885);
and UO_382 (O_382,N_9582,N_9917);
or UO_383 (O_383,N_9537,N_9716);
or UO_384 (O_384,N_9944,N_9689);
nand UO_385 (O_385,N_9611,N_9575);
xor UO_386 (O_386,N_9841,N_9530);
or UO_387 (O_387,N_9922,N_9738);
nor UO_388 (O_388,N_9789,N_9969);
or UO_389 (O_389,N_9854,N_9950);
xor UO_390 (O_390,N_9958,N_9637);
or UO_391 (O_391,N_9900,N_9977);
or UO_392 (O_392,N_9674,N_9669);
xor UO_393 (O_393,N_9864,N_9691);
or UO_394 (O_394,N_9843,N_9556);
nor UO_395 (O_395,N_9675,N_9954);
nor UO_396 (O_396,N_9861,N_9654);
xor UO_397 (O_397,N_9519,N_9977);
or UO_398 (O_398,N_9800,N_9671);
nor UO_399 (O_399,N_9993,N_9686);
xor UO_400 (O_400,N_9929,N_9845);
xor UO_401 (O_401,N_9522,N_9624);
xnor UO_402 (O_402,N_9754,N_9695);
or UO_403 (O_403,N_9940,N_9744);
and UO_404 (O_404,N_9885,N_9715);
or UO_405 (O_405,N_9663,N_9587);
nor UO_406 (O_406,N_9698,N_9829);
and UO_407 (O_407,N_9714,N_9855);
and UO_408 (O_408,N_9700,N_9843);
and UO_409 (O_409,N_9922,N_9592);
nand UO_410 (O_410,N_9531,N_9549);
nor UO_411 (O_411,N_9639,N_9585);
xnor UO_412 (O_412,N_9639,N_9529);
or UO_413 (O_413,N_9752,N_9604);
or UO_414 (O_414,N_9734,N_9622);
nand UO_415 (O_415,N_9992,N_9617);
nor UO_416 (O_416,N_9561,N_9866);
and UO_417 (O_417,N_9689,N_9673);
nor UO_418 (O_418,N_9801,N_9833);
xnor UO_419 (O_419,N_9643,N_9728);
xor UO_420 (O_420,N_9585,N_9522);
nand UO_421 (O_421,N_9759,N_9733);
xnor UO_422 (O_422,N_9879,N_9786);
xnor UO_423 (O_423,N_9534,N_9772);
and UO_424 (O_424,N_9524,N_9951);
and UO_425 (O_425,N_9728,N_9757);
and UO_426 (O_426,N_9764,N_9613);
nand UO_427 (O_427,N_9598,N_9697);
xor UO_428 (O_428,N_9563,N_9701);
and UO_429 (O_429,N_9674,N_9963);
xnor UO_430 (O_430,N_9625,N_9876);
and UO_431 (O_431,N_9589,N_9641);
or UO_432 (O_432,N_9794,N_9689);
or UO_433 (O_433,N_9729,N_9945);
xnor UO_434 (O_434,N_9824,N_9542);
xnor UO_435 (O_435,N_9945,N_9981);
nor UO_436 (O_436,N_9958,N_9952);
and UO_437 (O_437,N_9710,N_9832);
xor UO_438 (O_438,N_9911,N_9948);
and UO_439 (O_439,N_9749,N_9628);
nor UO_440 (O_440,N_9880,N_9755);
or UO_441 (O_441,N_9600,N_9994);
or UO_442 (O_442,N_9569,N_9736);
nand UO_443 (O_443,N_9626,N_9733);
nor UO_444 (O_444,N_9540,N_9731);
nor UO_445 (O_445,N_9980,N_9788);
xnor UO_446 (O_446,N_9980,N_9658);
xor UO_447 (O_447,N_9583,N_9710);
nand UO_448 (O_448,N_9748,N_9509);
xnor UO_449 (O_449,N_9624,N_9909);
nor UO_450 (O_450,N_9575,N_9892);
or UO_451 (O_451,N_9898,N_9879);
nor UO_452 (O_452,N_9918,N_9851);
nand UO_453 (O_453,N_9693,N_9894);
nand UO_454 (O_454,N_9896,N_9819);
xor UO_455 (O_455,N_9662,N_9696);
nand UO_456 (O_456,N_9698,N_9995);
xor UO_457 (O_457,N_9659,N_9945);
or UO_458 (O_458,N_9872,N_9608);
and UO_459 (O_459,N_9858,N_9550);
nand UO_460 (O_460,N_9642,N_9743);
xor UO_461 (O_461,N_9558,N_9586);
and UO_462 (O_462,N_9752,N_9557);
xnor UO_463 (O_463,N_9579,N_9992);
or UO_464 (O_464,N_9914,N_9702);
nor UO_465 (O_465,N_9940,N_9736);
nand UO_466 (O_466,N_9743,N_9710);
nand UO_467 (O_467,N_9509,N_9925);
nor UO_468 (O_468,N_9816,N_9578);
and UO_469 (O_469,N_9921,N_9579);
nor UO_470 (O_470,N_9841,N_9879);
or UO_471 (O_471,N_9977,N_9582);
and UO_472 (O_472,N_9827,N_9518);
nand UO_473 (O_473,N_9870,N_9814);
nor UO_474 (O_474,N_9913,N_9699);
nor UO_475 (O_475,N_9947,N_9876);
and UO_476 (O_476,N_9720,N_9754);
and UO_477 (O_477,N_9686,N_9565);
or UO_478 (O_478,N_9601,N_9857);
nand UO_479 (O_479,N_9743,N_9987);
nor UO_480 (O_480,N_9531,N_9992);
xnor UO_481 (O_481,N_9933,N_9627);
or UO_482 (O_482,N_9864,N_9815);
or UO_483 (O_483,N_9992,N_9506);
nor UO_484 (O_484,N_9719,N_9602);
nor UO_485 (O_485,N_9885,N_9787);
nand UO_486 (O_486,N_9692,N_9540);
nand UO_487 (O_487,N_9704,N_9701);
nand UO_488 (O_488,N_9524,N_9867);
xor UO_489 (O_489,N_9946,N_9570);
nand UO_490 (O_490,N_9722,N_9835);
nor UO_491 (O_491,N_9874,N_9747);
and UO_492 (O_492,N_9555,N_9919);
nor UO_493 (O_493,N_9756,N_9680);
and UO_494 (O_494,N_9913,N_9832);
nor UO_495 (O_495,N_9805,N_9891);
or UO_496 (O_496,N_9872,N_9859);
xor UO_497 (O_497,N_9937,N_9846);
xor UO_498 (O_498,N_9959,N_9538);
nor UO_499 (O_499,N_9653,N_9763);
xor UO_500 (O_500,N_9715,N_9989);
and UO_501 (O_501,N_9927,N_9687);
nand UO_502 (O_502,N_9912,N_9679);
xor UO_503 (O_503,N_9915,N_9740);
xnor UO_504 (O_504,N_9946,N_9723);
nor UO_505 (O_505,N_9927,N_9724);
or UO_506 (O_506,N_9559,N_9840);
or UO_507 (O_507,N_9663,N_9865);
xnor UO_508 (O_508,N_9572,N_9500);
and UO_509 (O_509,N_9767,N_9805);
nand UO_510 (O_510,N_9503,N_9596);
and UO_511 (O_511,N_9658,N_9635);
nor UO_512 (O_512,N_9747,N_9632);
xor UO_513 (O_513,N_9890,N_9822);
nor UO_514 (O_514,N_9612,N_9785);
nand UO_515 (O_515,N_9781,N_9638);
nand UO_516 (O_516,N_9846,N_9557);
nand UO_517 (O_517,N_9582,N_9974);
xor UO_518 (O_518,N_9718,N_9639);
or UO_519 (O_519,N_9932,N_9768);
nor UO_520 (O_520,N_9703,N_9982);
nand UO_521 (O_521,N_9638,N_9880);
xnor UO_522 (O_522,N_9838,N_9657);
nand UO_523 (O_523,N_9905,N_9882);
or UO_524 (O_524,N_9558,N_9697);
nor UO_525 (O_525,N_9502,N_9689);
nand UO_526 (O_526,N_9919,N_9892);
or UO_527 (O_527,N_9613,N_9802);
nor UO_528 (O_528,N_9997,N_9820);
xnor UO_529 (O_529,N_9831,N_9806);
nor UO_530 (O_530,N_9761,N_9899);
and UO_531 (O_531,N_9708,N_9881);
nand UO_532 (O_532,N_9986,N_9823);
or UO_533 (O_533,N_9639,N_9754);
nand UO_534 (O_534,N_9618,N_9570);
and UO_535 (O_535,N_9642,N_9922);
nand UO_536 (O_536,N_9922,N_9546);
xor UO_537 (O_537,N_9988,N_9969);
and UO_538 (O_538,N_9549,N_9739);
xor UO_539 (O_539,N_9739,N_9631);
and UO_540 (O_540,N_9993,N_9721);
or UO_541 (O_541,N_9697,N_9536);
nand UO_542 (O_542,N_9961,N_9978);
nor UO_543 (O_543,N_9732,N_9784);
and UO_544 (O_544,N_9959,N_9923);
and UO_545 (O_545,N_9837,N_9653);
and UO_546 (O_546,N_9883,N_9785);
or UO_547 (O_547,N_9562,N_9502);
nor UO_548 (O_548,N_9990,N_9874);
nor UO_549 (O_549,N_9997,N_9837);
or UO_550 (O_550,N_9733,N_9794);
or UO_551 (O_551,N_9928,N_9660);
or UO_552 (O_552,N_9897,N_9678);
nand UO_553 (O_553,N_9955,N_9558);
and UO_554 (O_554,N_9540,N_9971);
and UO_555 (O_555,N_9987,N_9994);
nand UO_556 (O_556,N_9594,N_9842);
or UO_557 (O_557,N_9679,N_9880);
nand UO_558 (O_558,N_9754,N_9774);
or UO_559 (O_559,N_9848,N_9564);
nand UO_560 (O_560,N_9831,N_9805);
nand UO_561 (O_561,N_9715,N_9639);
and UO_562 (O_562,N_9801,N_9573);
nor UO_563 (O_563,N_9713,N_9517);
xnor UO_564 (O_564,N_9536,N_9780);
or UO_565 (O_565,N_9591,N_9813);
or UO_566 (O_566,N_9559,N_9680);
nand UO_567 (O_567,N_9808,N_9746);
nor UO_568 (O_568,N_9653,N_9862);
xnor UO_569 (O_569,N_9802,N_9805);
and UO_570 (O_570,N_9900,N_9649);
and UO_571 (O_571,N_9735,N_9602);
nand UO_572 (O_572,N_9766,N_9687);
nand UO_573 (O_573,N_9716,N_9530);
or UO_574 (O_574,N_9661,N_9880);
nand UO_575 (O_575,N_9997,N_9506);
nor UO_576 (O_576,N_9759,N_9546);
xnor UO_577 (O_577,N_9516,N_9869);
nand UO_578 (O_578,N_9757,N_9655);
xor UO_579 (O_579,N_9529,N_9772);
nor UO_580 (O_580,N_9963,N_9982);
nand UO_581 (O_581,N_9573,N_9891);
or UO_582 (O_582,N_9998,N_9683);
xor UO_583 (O_583,N_9807,N_9704);
xor UO_584 (O_584,N_9655,N_9660);
xor UO_585 (O_585,N_9757,N_9764);
nand UO_586 (O_586,N_9873,N_9703);
and UO_587 (O_587,N_9630,N_9969);
or UO_588 (O_588,N_9739,N_9719);
nand UO_589 (O_589,N_9630,N_9535);
and UO_590 (O_590,N_9667,N_9742);
and UO_591 (O_591,N_9916,N_9570);
xor UO_592 (O_592,N_9568,N_9767);
nor UO_593 (O_593,N_9601,N_9944);
and UO_594 (O_594,N_9947,N_9767);
nor UO_595 (O_595,N_9867,N_9933);
nor UO_596 (O_596,N_9981,N_9775);
and UO_597 (O_597,N_9868,N_9820);
and UO_598 (O_598,N_9855,N_9659);
xor UO_599 (O_599,N_9784,N_9821);
nand UO_600 (O_600,N_9868,N_9513);
nand UO_601 (O_601,N_9868,N_9914);
nand UO_602 (O_602,N_9586,N_9589);
nand UO_603 (O_603,N_9760,N_9611);
xor UO_604 (O_604,N_9872,N_9712);
and UO_605 (O_605,N_9927,N_9778);
and UO_606 (O_606,N_9740,N_9978);
and UO_607 (O_607,N_9808,N_9701);
xnor UO_608 (O_608,N_9523,N_9867);
or UO_609 (O_609,N_9611,N_9866);
nor UO_610 (O_610,N_9865,N_9908);
nor UO_611 (O_611,N_9660,N_9672);
xor UO_612 (O_612,N_9730,N_9649);
xor UO_613 (O_613,N_9976,N_9851);
nand UO_614 (O_614,N_9701,N_9765);
and UO_615 (O_615,N_9987,N_9713);
and UO_616 (O_616,N_9545,N_9693);
or UO_617 (O_617,N_9573,N_9876);
or UO_618 (O_618,N_9960,N_9533);
nor UO_619 (O_619,N_9619,N_9898);
or UO_620 (O_620,N_9816,N_9599);
nand UO_621 (O_621,N_9806,N_9745);
nor UO_622 (O_622,N_9520,N_9819);
and UO_623 (O_623,N_9536,N_9521);
xor UO_624 (O_624,N_9570,N_9788);
nand UO_625 (O_625,N_9858,N_9797);
xnor UO_626 (O_626,N_9877,N_9554);
xor UO_627 (O_627,N_9970,N_9600);
nand UO_628 (O_628,N_9812,N_9901);
nor UO_629 (O_629,N_9762,N_9676);
and UO_630 (O_630,N_9633,N_9855);
nand UO_631 (O_631,N_9686,N_9778);
xnor UO_632 (O_632,N_9649,N_9669);
or UO_633 (O_633,N_9519,N_9617);
xor UO_634 (O_634,N_9642,N_9508);
xor UO_635 (O_635,N_9700,N_9665);
or UO_636 (O_636,N_9996,N_9860);
and UO_637 (O_637,N_9618,N_9550);
nand UO_638 (O_638,N_9599,N_9759);
nor UO_639 (O_639,N_9639,N_9693);
xnor UO_640 (O_640,N_9686,N_9840);
nor UO_641 (O_641,N_9845,N_9591);
xnor UO_642 (O_642,N_9951,N_9746);
nand UO_643 (O_643,N_9855,N_9666);
or UO_644 (O_644,N_9909,N_9982);
xnor UO_645 (O_645,N_9827,N_9713);
and UO_646 (O_646,N_9871,N_9728);
and UO_647 (O_647,N_9869,N_9757);
nor UO_648 (O_648,N_9912,N_9816);
or UO_649 (O_649,N_9502,N_9557);
xor UO_650 (O_650,N_9704,N_9871);
or UO_651 (O_651,N_9848,N_9614);
xor UO_652 (O_652,N_9685,N_9750);
nand UO_653 (O_653,N_9900,N_9709);
and UO_654 (O_654,N_9932,N_9900);
xnor UO_655 (O_655,N_9507,N_9865);
or UO_656 (O_656,N_9726,N_9641);
nand UO_657 (O_657,N_9790,N_9809);
nand UO_658 (O_658,N_9718,N_9829);
nor UO_659 (O_659,N_9732,N_9623);
nand UO_660 (O_660,N_9972,N_9803);
nand UO_661 (O_661,N_9799,N_9985);
xnor UO_662 (O_662,N_9978,N_9555);
nor UO_663 (O_663,N_9797,N_9887);
xnor UO_664 (O_664,N_9872,N_9998);
xor UO_665 (O_665,N_9938,N_9616);
nand UO_666 (O_666,N_9782,N_9645);
or UO_667 (O_667,N_9602,N_9971);
xnor UO_668 (O_668,N_9562,N_9552);
and UO_669 (O_669,N_9599,N_9847);
and UO_670 (O_670,N_9935,N_9706);
or UO_671 (O_671,N_9807,N_9969);
nor UO_672 (O_672,N_9662,N_9519);
nand UO_673 (O_673,N_9786,N_9911);
or UO_674 (O_674,N_9854,N_9699);
nor UO_675 (O_675,N_9782,N_9719);
xor UO_676 (O_676,N_9906,N_9639);
nand UO_677 (O_677,N_9749,N_9588);
and UO_678 (O_678,N_9539,N_9720);
nor UO_679 (O_679,N_9525,N_9876);
nor UO_680 (O_680,N_9667,N_9914);
or UO_681 (O_681,N_9982,N_9833);
xnor UO_682 (O_682,N_9582,N_9623);
xor UO_683 (O_683,N_9568,N_9547);
nand UO_684 (O_684,N_9987,N_9636);
or UO_685 (O_685,N_9877,N_9973);
nor UO_686 (O_686,N_9891,N_9874);
and UO_687 (O_687,N_9980,N_9949);
and UO_688 (O_688,N_9942,N_9705);
or UO_689 (O_689,N_9868,N_9857);
and UO_690 (O_690,N_9581,N_9641);
or UO_691 (O_691,N_9552,N_9542);
xnor UO_692 (O_692,N_9854,N_9835);
nor UO_693 (O_693,N_9895,N_9589);
nor UO_694 (O_694,N_9852,N_9831);
xor UO_695 (O_695,N_9525,N_9858);
xnor UO_696 (O_696,N_9576,N_9963);
nor UO_697 (O_697,N_9594,N_9685);
nand UO_698 (O_698,N_9532,N_9989);
and UO_699 (O_699,N_9725,N_9693);
or UO_700 (O_700,N_9614,N_9967);
nand UO_701 (O_701,N_9577,N_9983);
xor UO_702 (O_702,N_9643,N_9544);
nor UO_703 (O_703,N_9828,N_9591);
and UO_704 (O_704,N_9998,N_9533);
nor UO_705 (O_705,N_9538,N_9787);
or UO_706 (O_706,N_9909,N_9596);
nor UO_707 (O_707,N_9637,N_9782);
or UO_708 (O_708,N_9540,N_9941);
nor UO_709 (O_709,N_9560,N_9568);
or UO_710 (O_710,N_9795,N_9574);
or UO_711 (O_711,N_9816,N_9695);
and UO_712 (O_712,N_9533,N_9823);
nand UO_713 (O_713,N_9767,N_9920);
and UO_714 (O_714,N_9568,N_9815);
nor UO_715 (O_715,N_9514,N_9554);
nor UO_716 (O_716,N_9878,N_9851);
and UO_717 (O_717,N_9626,N_9684);
nor UO_718 (O_718,N_9824,N_9650);
nor UO_719 (O_719,N_9817,N_9764);
or UO_720 (O_720,N_9670,N_9694);
nor UO_721 (O_721,N_9947,N_9983);
nor UO_722 (O_722,N_9732,N_9892);
and UO_723 (O_723,N_9679,N_9741);
or UO_724 (O_724,N_9546,N_9651);
xnor UO_725 (O_725,N_9829,N_9508);
nand UO_726 (O_726,N_9989,N_9958);
or UO_727 (O_727,N_9984,N_9579);
nand UO_728 (O_728,N_9785,N_9859);
and UO_729 (O_729,N_9607,N_9848);
or UO_730 (O_730,N_9695,N_9860);
nor UO_731 (O_731,N_9686,N_9793);
nor UO_732 (O_732,N_9741,N_9948);
nor UO_733 (O_733,N_9823,N_9632);
or UO_734 (O_734,N_9755,N_9899);
xnor UO_735 (O_735,N_9549,N_9816);
and UO_736 (O_736,N_9801,N_9941);
xor UO_737 (O_737,N_9995,N_9949);
or UO_738 (O_738,N_9721,N_9798);
nand UO_739 (O_739,N_9982,N_9609);
or UO_740 (O_740,N_9732,N_9593);
and UO_741 (O_741,N_9688,N_9609);
or UO_742 (O_742,N_9896,N_9737);
and UO_743 (O_743,N_9843,N_9909);
or UO_744 (O_744,N_9862,N_9687);
or UO_745 (O_745,N_9998,N_9791);
and UO_746 (O_746,N_9642,N_9937);
or UO_747 (O_747,N_9690,N_9874);
or UO_748 (O_748,N_9535,N_9776);
or UO_749 (O_749,N_9525,N_9879);
nor UO_750 (O_750,N_9992,N_9556);
nor UO_751 (O_751,N_9971,N_9728);
or UO_752 (O_752,N_9582,N_9542);
nand UO_753 (O_753,N_9854,N_9749);
nand UO_754 (O_754,N_9819,N_9949);
and UO_755 (O_755,N_9514,N_9788);
nand UO_756 (O_756,N_9608,N_9798);
xor UO_757 (O_757,N_9806,N_9975);
xnor UO_758 (O_758,N_9735,N_9930);
or UO_759 (O_759,N_9627,N_9899);
or UO_760 (O_760,N_9695,N_9601);
xor UO_761 (O_761,N_9799,N_9984);
xnor UO_762 (O_762,N_9798,N_9752);
nand UO_763 (O_763,N_9804,N_9886);
nor UO_764 (O_764,N_9629,N_9873);
or UO_765 (O_765,N_9645,N_9742);
nor UO_766 (O_766,N_9754,N_9514);
and UO_767 (O_767,N_9710,N_9915);
nand UO_768 (O_768,N_9562,N_9659);
nand UO_769 (O_769,N_9648,N_9598);
nand UO_770 (O_770,N_9703,N_9699);
xnor UO_771 (O_771,N_9770,N_9995);
and UO_772 (O_772,N_9693,N_9967);
or UO_773 (O_773,N_9660,N_9614);
nand UO_774 (O_774,N_9755,N_9869);
nor UO_775 (O_775,N_9548,N_9785);
xnor UO_776 (O_776,N_9819,N_9510);
xnor UO_777 (O_777,N_9706,N_9602);
xor UO_778 (O_778,N_9992,N_9722);
nand UO_779 (O_779,N_9968,N_9872);
and UO_780 (O_780,N_9790,N_9670);
xnor UO_781 (O_781,N_9936,N_9874);
or UO_782 (O_782,N_9572,N_9786);
and UO_783 (O_783,N_9693,N_9621);
nor UO_784 (O_784,N_9731,N_9699);
nor UO_785 (O_785,N_9516,N_9610);
and UO_786 (O_786,N_9656,N_9558);
and UO_787 (O_787,N_9584,N_9561);
nor UO_788 (O_788,N_9837,N_9761);
nand UO_789 (O_789,N_9785,N_9866);
nand UO_790 (O_790,N_9610,N_9910);
or UO_791 (O_791,N_9503,N_9923);
or UO_792 (O_792,N_9824,N_9580);
or UO_793 (O_793,N_9773,N_9913);
xor UO_794 (O_794,N_9771,N_9640);
or UO_795 (O_795,N_9962,N_9535);
xnor UO_796 (O_796,N_9929,N_9643);
and UO_797 (O_797,N_9623,N_9966);
xnor UO_798 (O_798,N_9939,N_9770);
or UO_799 (O_799,N_9848,N_9791);
xor UO_800 (O_800,N_9666,N_9894);
and UO_801 (O_801,N_9657,N_9617);
xnor UO_802 (O_802,N_9865,N_9577);
nor UO_803 (O_803,N_9846,N_9712);
or UO_804 (O_804,N_9926,N_9691);
nor UO_805 (O_805,N_9907,N_9539);
and UO_806 (O_806,N_9972,N_9967);
nand UO_807 (O_807,N_9589,N_9763);
nor UO_808 (O_808,N_9825,N_9646);
nand UO_809 (O_809,N_9675,N_9725);
xor UO_810 (O_810,N_9997,N_9733);
nor UO_811 (O_811,N_9814,N_9730);
xnor UO_812 (O_812,N_9560,N_9814);
or UO_813 (O_813,N_9802,N_9609);
nor UO_814 (O_814,N_9821,N_9616);
or UO_815 (O_815,N_9588,N_9552);
or UO_816 (O_816,N_9732,N_9572);
nor UO_817 (O_817,N_9652,N_9668);
nor UO_818 (O_818,N_9685,N_9963);
nor UO_819 (O_819,N_9527,N_9893);
and UO_820 (O_820,N_9772,N_9721);
nand UO_821 (O_821,N_9809,N_9505);
and UO_822 (O_822,N_9630,N_9514);
nor UO_823 (O_823,N_9886,N_9690);
and UO_824 (O_824,N_9843,N_9925);
xnor UO_825 (O_825,N_9734,N_9515);
or UO_826 (O_826,N_9886,N_9542);
nand UO_827 (O_827,N_9688,N_9668);
or UO_828 (O_828,N_9503,N_9616);
or UO_829 (O_829,N_9871,N_9733);
xor UO_830 (O_830,N_9697,N_9505);
nand UO_831 (O_831,N_9788,N_9819);
or UO_832 (O_832,N_9536,N_9875);
and UO_833 (O_833,N_9881,N_9673);
and UO_834 (O_834,N_9815,N_9985);
xnor UO_835 (O_835,N_9969,N_9542);
nor UO_836 (O_836,N_9653,N_9859);
nand UO_837 (O_837,N_9905,N_9928);
or UO_838 (O_838,N_9670,N_9905);
or UO_839 (O_839,N_9985,N_9603);
nor UO_840 (O_840,N_9623,N_9987);
or UO_841 (O_841,N_9693,N_9525);
nand UO_842 (O_842,N_9559,N_9668);
nor UO_843 (O_843,N_9933,N_9932);
xnor UO_844 (O_844,N_9732,N_9688);
and UO_845 (O_845,N_9854,N_9533);
or UO_846 (O_846,N_9636,N_9820);
nor UO_847 (O_847,N_9730,N_9517);
nor UO_848 (O_848,N_9670,N_9738);
xor UO_849 (O_849,N_9991,N_9920);
or UO_850 (O_850,N_9579,N_9660);
nand UO_851 (O_851,N_9756,N_9916);
nand UO_852 (O_852,N_9641,N_9585);
and UO_853 (O_853,N_9907,N_9507);
or UO_854 (O_854,N_9529,N_9536);
xnor UO_855 (O_855,N_9796,N_9979);
and UO_856 (O_856,N_9646,N_9552);
nor UO_857 (O_857,N_9871,N_9718);
or UO_858 (O_858,N_9984,N_9996);
nor UO_859 (O_859,N_9989,N_9851);
or UO_860 (O_860,N_9856,N_9733);
nand UO_861 (O_861,N_9513,N_9754);
nor UO_862 (O_862,N_9990,N_9956);
or UO_863 (O_863,N_9869,N_9533);
nor UO_864 (O_864,N_9522,N_9810);
and UO_865 (O_865,N_9940,N_9740);
or UO_866 (O_866,N_9714,N_9770);
nor UO_867 (O_867,N_9941,N_9565);
and UO_868 (O_868,N_9618,N_9589);
xor UO_869 (O_869,N_9777,N_9530);
xor UO_870 (O_870,N_9643,N_9742);
nand UO_871 (O_871,N_9952,N_9505);
xnor UO_872 (O_872,N_9538,N_9593);
xor UO_873 (O_873,N_9752,N_9767);
nand UO_874 (O_874,N_9966,N_9569);
nand UO_875 (O_875,N_9794,N_9642);
or UO_876 (O_876,N_9706,N_9818);
and UO_877 (O_877,N_9921,N_9501);
nand UO_878 (O_878,N_9903,N_9649);
or UO_879 (O_879,N_9563,N_9971);
and UO_880 (O_880,N_9588,N_9779);
nand UO_881 (O_881,N_9964,N_9553);
or UO_882 (O_882,N_9859,N_9670);
nor UO_883 (O_883,N_9768,N_9868);
nor UO_884 (O_884,N_9547,N_9510);
xor UO_885 (O_885,N_9846,N_9649);
nand UO_886 (O_886,N_9946,N_9586);
or UO_887 (O_887,N_9631,N_9735);
and UO_888 (O_888,N_9552,N_9998);
or UO_889 (O_889,N_9795,N_9695);
xnor UO_890 (O_890,N_9596,N_9869);
and UO_891 (O_891,N_9724,N_9597);
nor UO_892 (O_892,N_9987,N_9539);
nor UO_893 (O_893,N_9752,N_9651);
and UO_894 (O_894,N_9828,N_9889);
and UO_895 (O_895,N_9962,N_9972);
xor UO_896 (O_896,N_9947,N_9749);
nand UO_897 (O_897,N_9721,N_9527);
nor UO_898 (O_898,N_9950,N_9521);
or UO_899 (O_899,N_9572,N_9913);
nand UO_900 (O_900,N_9791,N_9777);
nor UO_901 (O_901,N_9870,N_9789);
xnor UO_902 (O_902,N_9995,N_9669);
nor UO_903 (O_903,N_9778,N_9765);
nor UO_904 (O_904,N_9504,N_9886);
and UO_905 (O_905,N_9653,N_9795);
xor UO_906 (O_906,N_9779,N_9627);
nand UO_907 (O_907,N_9511,N_9718);
nor UO_908 (O_908,N_9511,N_9540);
or UO_909 (O_909,N_9685,N_9998);
or UO_910 (O_910,N_9753,N_9648);
xor UO_911 (O_911,N_9997,N_9816);
or UO_912 (O_912,N_9528,N_9548);
and UO_913 (O_913,N_9639,N_9838);
xnor UO_914 (O_914,N_9617,N_9826);
nand UO_915 (O_915,N_9781,N_9648);
nand UO_916 (O_916,N_9831,N_9827);
xor UO_917 (O_917,N_9957,N_9974);
nor UO_918 (O_918,N_9943,N_9608);
nor UO_919 (O_919,N_9989,N_9754);
nor UO_920 (O_920,N_9620,N_9548);
and UO_921 (O_921,N_9518,N_9613);
or UO_922 (O_922,N_9977,N_9858);
nor UO_923 (O_923,N_9937,N_9787);
xnor UO_924 (O_924,N_9680,N_9813);
and UO_925 (O_925,N_9746,N_9955);
xnor UO_926 (O_926,N_9542,N_9658);
and UO_927 (O_927,N_9670,N_9974);
nand UO_928 (O_928,N_9786,N_9978);
nand UO_929 (O_929,N_9686,N_9871);
xnor UO_930 (O_930,N_9606,N_9967);
nor UO_931 (O_931,N_9742,N_9593);
and UO_932 (O_932,N_9969,N_9794);
xnor UO_933 (O_933,N_9899,N_9532);
nor UO_934 (O_934,N_9636,N_9815);
or UO_935 (O_935,N_9601,N_9600);
or UO_936 (O_936,N_9963,N_9619);
nand UO_937 (O_937,N_9955,N_9773);
xor UO_938 (O_938,N_9799,N_9923);
nand UO_939 (O_939,N_9753,N_9730);
nor UO_940 (O_940,N_9775,N_9652);
nand UO_941 (O_941,N_9618,N_9745);
or UO_942 (O_942,N_9682,N_9722);
xor UO_943 (O_943,N_9629,N_9871);
or UO_944 (O_944,N_9849,N_9614);
xor UO_945 (O_945,N_9636,N_9643);
nor UO_946 (O_946,N_9647,N_9909);
xor UO_947 (O_947,N_9660,N_9746);
and UO_948 (O_948,N_9616,N_9722);
nor UO_949 (O_949,N_9872,N_9691);
xor UO_950 (O_950,N_9586,N_9744);
nor UO_951 (O_951,N_9958,N_9685);
and UO_952 (O_952,N_9967,N_9588);
nand UO_953 (O_953,N_9998,N_9592);
and UO_954 (O_954,N_9603,N_9503);
nand UO_955 (O_955,N_9807,N_9695);
nand UO_956 (O_956,N_9784,N_9626);
nand UO_957 (O_957,N_9966,N_9880);
nand UO_958 (O_958,N_9776,N_9989);
and UO_959 (O_959,N_9956,N_9686);
or UO_960 (O_960,N_9701,N_9815);
nor UO_961 (O_961,N_9789,N_9660);
nor UO_962 (O_962,N_9795,N_9524);
nor UO_963 (O_963,N_9575,N_9539);
nand UO_964 (O_964,N_9876,N_9592);
nand UO_965 (O_965,N_9949,N_9582);
nand UO_966 (O_966,N_9510,N_9600);
or UO_967 (O_967,N_9654,N_9840);
nand UO_968 (O_968,N_9643,N_9867);
xnor UO_969 (O_969,N_9909,N_9598);
xor UO_970 (O_970,N_9531,N_9944);
nand UO_971 (O_971,N_9995,N_9935);
nand UO_972 (O_972,N_9589,N_9952);
and UO_973 (O_973,N_9580,N_9623);
and UO_974 (O_974,N_9812,N_9658);
or UO_975 (O_975,N_9673,N_9674);
xnor UO_976 (O_976,N_9503,N_9846);
and UO_977 (O_977,N_9821,N_9892);
or UO_978 (O_978,N_9797,N_9802);
xnor UO_979 (O_979,N_9852,N_9745);
and UO_980 (O_980,N_9613,N_9505);
xor UO_981 (O_981,N_9812,N_9847);
xnor UO_982 (O_982,N_9811,N_9659);
or UO_983 (O_983,N_9964,N_9658);
xnor UO_984 (O_984,N_9905,N_9782);
or UO_985 (O_985,N_9883,N_9867);
xor UO_986 (O_986,N_9753,N_9954);
or UO_987 (O_987,N_9693,N_9569);
nand UO_988 (O_988,N_9729,N_9513);
or UO_989 (O_989,N_9706,N_9921);
and UO_990 (O_990,N_9910,N_9748);
nand UO_991 (O_991,N_9981,N_9518);
or UO_992 (O_992,N_9933,N_9806);
or UO_993 (O_993,N_9678,N_9908);
nor UO_994 (O_994,N_9881,N_9677);
or UO_995 (O_995,N_9569,N_9855);
and UO_996 (O_996,N_9586,N_9761);
and UO_997 (O_997,N_9542,N_9909);
and UO_998 (O_998,N_9943,N_9973);
xnor UO_999 (O_999,N_9610,N_9825);
nor UO_1000 (O_1000,N_9621,N_9589);
and UO_1001 (O_1001,N_9760,N_9528);
and UO_1002 (O_1002,N_9951,N_9855);
nor UO_1003 (O_1003,N_9842,N_9945);
nand UO_1004 (O_1004,N_9695,N_9712);
and UO_1005 (O_1005,N_9614,N_9738);
and UO_1006 (O_1006,N_9560,N_9577);
nor UO_1007 (O_1007,N_9732,N_9695);
and UO_1008 (O_1008,N_9900,N_9612);
and UO_1009 (O_1009,N_9545,N_9607);
and UO_1010 (O_1010,N_9806,N_9743);
and UO_1011 (O_1011,N_9632,N_9786);
or UO_1012 (O_1012,N_9545,N_9836);
or UO_1013 (O_1013,N_9807,N_9863);
nor UO_1014 (O_1014,N_9823,N_9752);
and UO_1015 (O_1015,N_9999,N_9522);
or UO_1016 (O_1016,N_9513,N_9650);
or UO_1017 (O_1017,N_9811,N_9625);
xor UO_1018 (O_1018,N_9963,N_9625);
nand UO_1019 (O_1019,N_9976,N_9714);
and UO_1020 (O_1020,N_9561,N_9948);
xor UO_1021 (O_1021,N_9881,N_9604);
and UO_1022 (O_1022,N_9619,N_9570);
xor UO_1023 (O_1023,N_9568,N_9693);
nor UO_1024 (O_1024,N_9825,N_9844);
nor UO_1025 (O_1025,N_9867,N_9664);
and UO_1026 (O_1026,N_9836,N_9766);
or UO_1027 (O_1027,N_9572,N_9979);
or UO_1028 (O_1028,N_9720,N_9736);
nor UO_1029 (O_1029,N_9525,N_9628);
nand UO_1030 (O_1030,N_9692,N_9546);
nor UO_1031 (O_1031,N_9557,N_9754);
and UO_1032 (O_1032,N_9877,N_9897);
and UO_1033 (O_1033,N_9543,N_9953);
nor UO_1034 (O_1034,N_9578,N_9772);
or UO_1035 (O_1035,N_9744,N_9904);
or UO_1036 (O_1036,N_9501,N_9806);
or UO_1037 (O_1037,N_9954,N_9618);
nor UO_1038 (O_1038,N_9820,N_9825);
or UO_1039 (O_1039,N_9521,N_9728);
nor UO_1040 (O_1040,N_9898,N_9526);
or UO_1041 (O_1041,N_9805,N_9616);
and UO_1042 (O_1042,N_9591,N_9507);
nand UO_1043 (O_1043,N_9596,N_9939);
or UO_1044 (O_1044,N_9869,N_9805);
xor UO_1045 (O_1045,N_9976,N_9502);
nand UO_1046 (O_1046,N_9624,N_9538);
xnor UO_1047 (O_1047,N_9941,N_9584);
nor UO_1048 (O_1048,N_9531,N_9995);
xor UO_1049 (O_1049,N_9852,N_9636);
nand UO_1050 (O_1050,N_9549,N_9893);
and UO_1051 (O_1051,N_9945,N_9551);
xnor UO_1052 (O_1052,N_9721,N_9582);
xnor UO_1053 (O_1053,N_9972,N_9798);
or UO_1054 (O_1054,N_9819,N_9791);
and UO_1055 (O_1055,N_9903,N_9908);
nand UO_1056 (O_1056,N_9905,N_9733);
nand UO_1057 (O_1057,N_9686,N_9746);
xor UO_1058 (O_1058,N_9790,N_9951);
nor UO_1059 (O_1059,N_9671,N_9947);
nor UO_1060 (O_1060,N_9966,N_9669);
or UO_1061 (O_1061,N_9768,N_9820);
nand UO_1062 (O_1062,N_9608,N_9620);
nand UO_1063 (O_1063,N_9918,N_9737);
and UO_1064 (O_1064,N_9957,N_9889);
nor UO_1065 (O_1065,N_9728,N_9930);
nor UO_1066 (O_1066,N_9674,N_9647);
nor UO_1067 (O_1067,N_9505,N_9855);
nand UO_1068 (O_1068,N_9733,N_9580);
xor UO_1069 (O_1069,N_9560,N_9711);
nand UO_1070 (O_1070,N_9583,N_9837);
and UO_1071 (O_1071,N_9874,N_9529);
xor UO_1072 (O_1072,N_9643,N_9878);
nand UO_1073 (O_1073,N_9885,N_9534);
or UO_1074 (O_1074,N_9754,N_9897);
nand UO_1075 (O_1075,N_9832,N_9808);
or UO_1076 (O_1076,N_9579,N_9657);
nor UO_1077 (O_1077,N_9560,N_9871);
nor UO_1078 (O_1078,N_9702,N_9991);
or UO_1079 (O_1079,N_9826,N_9597);
and UO_1080 (O_1080,N_9760,N_9536);
or UO_1081 (O_1081,N_9557,N_9906);
nor UO_1082 (O_1082,N_9612,N_9663);
xnor UO_1083 (O_1083,N_9657,N_9962);
or UO_1084 (O_1084,N_9616,N_9935);
nand UO_1085 (O_1085,N_9523,N_9511);
nor UO_1086 (O_1086,N_9975,N_9692);
xor UO_1087 (O_1087,N_9946,N_9799);
nand UO_1088 (O_1088,N_9881,N_9655);
nor UO_1089 (O_1089,N_9875,N_9873);
nor UO_1090 (O_1090,N_9965,N_9789);
nand UO_1091 (O_1091,N_9869,N_9631);
nand UO_1092 (O_1092,N_9929,N_9890);
nand UO_1093 (O_1093,N_9972,N_9551);
nor UO_1094 (O_1094,N_9632,N_9921);
xnor UO_1095 (O_1095,N_9928,N_9841);
and UO_1096 (O_1096,N_9746,N_9983);
xor UO_1097 (O_1097,N_9580,N_9709);
and UO_1098 (O_1098,N_9509,N_9814);
xnor UO_1099 (O_1099,N_9731,N_9583);
or UO_1100 (O_1100,N_9562,N_9892);
xnor UO_1101 (O_1101,N_9574,N_9826);
nand UO_1102 (O_1102,N_9904,N_9653);
nor UO_1103 (O_1103,N_9808,N_9850);
xnor UO_1104 (O_1104,N_9790,N_9643);
xor UO_1105 (O_1105,N_9640,N_9741);
or UO_1106 (O_1106,N_9880,N_9625);
or UO_1107 (O_1107,N_9535,N_9586);
xnor UO_1108 (O_1108,N_9691,N_9689);
or UO_1109 (O_1109,N_9813,N_9984);
xor UO_1110 (O_1110,N_9640,N_9752);
and UO_1111 (O_1111,N_9632,N_9906);
xnor UO_1112 (O_1112,N_9952,N_9858);
nor UO_1113 (O_1113,N_9637,N_9983);
nor UO_1114 (O_1114,N_9719,N_9939);
and UO_1115 (O_1115,N_9806,N_9976);
nor UO_1116 (O_1116,N_9764,N_9880);
or UO_1117 (O_1117,N_9947,N_9887);
xnor UO_1118 (O_1118,N_9898,N_9744);
and UO_1119 (O_1119,N_9807,N_9943);
and UO_1120 (O_1120,N_9663,N_9746);
nand UO_1121 (O_1121,N_9576,N_9597);
nor UO_1122 (O_1122,N_9677,N_9513);
xnor UO_1123 (O_1123,N_9906,N_9870);
nand UO_1124 (O_1124,N_9989,N_9578);
nand UO_1125 (O_1125,N_9913,N_9521);
or UO_1126 (O_1126,N_9737,N_9633);
nand UO_1127 (O_1127,N_9910,N_9859);
or UO_1128 (O_1128,N_9814,N_9724);
nor UO_1129 (O_1129,N_9749,N_9622);
nand UO_1130 (O_1130,N_9858,N_9722);
nor UO_1131 (O_1131,N_9892,N_9828);
or UO_1132 (O_1132,N_9679,N_9651);
or UO_1133 (O_1133,N_9757,N_9930);
or UO_1134 (O_1134,N_9809,N_9858);
xnor UO_1135 (O_1135,N_9518,N_9702);
xor UO_1136 (O_1136,N_9851,N_9874);
nor UO_1137 (O_1137,N_9904,N_9834);
nor UO_1138 (O_1138,N_9726,N_9595);
nor UO_1139 (O_1139,N_9636,N_9632);
and UO_1140 (O_1140,N_9840,N_9770);
nor UO_1141 (O_1141,N_9591,N_9571);
xor UO_1142 (O_1142,N_9767,N_9780);
nor UO_1143 (O_1143,N_9639,N_9842);
nand UO_1144 (O_1144,N_9794,N_9773);
or UO_1145 (O_1145,N_9699,N_9621);
nor UO_1146 (O_1146,N_9619,N_9896);
or UO_1147 (O_1147,N_9690,N_9912);
and UO_1148 (O_1148,N_9980,N_9977);
xnor UO_1149 (O_1149,N_9923,N_9979);
and UO_1150 (O_1150,N_9582,N_9594);
nor UO_1151 (O_1151,N_9896,N_9736);
nor UO_1152 (O_1152,N_9746,N_9834);
nand UO_1153 (O_1153,N_9859,N_9856);
nand UO_1154 (O_1154,N_9780,N_9540);
nor UO_1155 (O_1155,N_9849,N_9878);
nand UO_1156 (O_1156,N_9990,N_9918);
xnor UO_1157 (O_1157,N_9524,N_9743);
and UO_1158 (O_1158,N_9668,N_9978);
and UO_1159 (O_1159,N_9572,N_9584);
nand UO_1160 (O_1160,N_9791,N_9968);
nand UO_1161 (O_1161,N_9967,N_9998);
and UO_1162 (O_1162,N_9675,N_9844);
or UO_1163 (O_1163,N_9753,N_9990);
nor UO_1164 (O_1164,N_9757,N_9974);
and UO_1165 (O_1165,N_9919,N_9913);
and UO_1166 (O_1166,N_9576,N_9980);
and UO_1167 (O_1167,N_9944,N_9849);
and UO_1168 (O_1168,N_9705,N_9636);
and UO_1169 (O_1169,N_9522,N_9651);
nand UO_1170 (O_1170,N_9660,N_9719);
xor UO_1171 (O_1171,N_9960,N_9593);
xor UO_1172 (O_1172,N_9581,N_9546);
and UO_1173 (O_1173,N_9949,N_9758);
nand UO_1174 (O_1174,N_9748,N_9884);
or UO_1175 (O_1175,N_9834,N_9503);
or UO_1176 (O_1176,N_9930,N_9545);
xnor UO_1177 (O_1177,N_9578,N_9680);
and UO_1178 (O_1178,N_9512,N_9570);
xor UO_1179 (O_1179,N_9885,N_9666);
xnor UO_1180 (O_1180,N_9881,N_9632);
nand UO_1181 (O_1181,N_9906,N_9708);
xnor UO_1182 (O_1182,N_9857,N_9815);
nor UO_1183 (O_1183,N_9543,N_9614);
nand UO_1184 (O_1184,N_9642,N_9650);
xor UO_1185 (O_1185,N_9760,N_9619);
and UO_1186 (O_1186,N_9938,N_9837);
and UO_1187 (O_1187,N_9549,N_9959);
xnor UO_1188 (O_1188,N_9665,N_9977);
or UO_1189 (O_1189,N_9550,N_9804);
nand UO_1190 (O_1190,N_9719,N_9941);
or UO_1191 (O_1191,N_9575,N_9927);
xor UO_1192 (O_1192,N_9964,N_9991);
nor UO_1193 (O_1193,N_9576,N_9629);
or UO_1194 (O_1194,N_9940,N_9902);
nand UO_1195 (O_1195,N_9681,N_9613);
nand UO_1196 (O_1196,N_9940,N_9531);
and UO_1197 (O_1197,N_9936,N_9823);
and UO_1198 (O_1198,N_9514,N_9868);
xor UO_1199 (O_1199,N_9923,N_9727);
nand UO_1200 (O_1200,N_9795,N_9826);
or UO_1201 (O_1201,N_9519,N_9708);
and UO_1202 (O_1202,N_9774,N_9640);
xnor UO_1203 (O_1203,N_9893,N_9642);
or UO_1204 (O_1204,N_9690,N_9894);
or UO_1205 (O_1205,N_9692,N_9903);
or UO_1206 (O_1206,N_9703,N_9990);
nor UO_1207 (O_1207,N_9580,N_9878);
xor UO_1208 (O_1208,N_9576,N_9999);
xor UO_1209 (O_1209,N_9984,N_9657);
nor UO_1210 (O_1210,N_9827,N_9758);
xor UO_1211 (O_1211,N_9548,N_9579);
and UO_1212 (O_1212,N_9801,N_9795);
xor UO_1213 (O_1213,N_9527,N_9762);
nand UO_1214 (O_1214,N_9811,N_9943);
xnor UO_1215 (O_1215,N_9525,N_9826);
xor UO_1216 (O_1216,N_9810,N_9748);
nand UO_1217 (O_1217,N_9551,N_9631);
nor UO_1218 (O_1218,N_9577,N_9950);
and UO_1219 (O_1219,N_9561,N_9994);
or UO_1220 (O_1220,N_9630,N_9865);
nor UO_1221 (O_1221,N_9785,N_9928);
nor UO_1222 (O_1222,N_9981,N_9918);
nor UO_1223 (O_1223,N_9617,N_9719);
and UO_1224 (O_1224,N_9777,N_9584);
nor UO_1225 (O_1225,N_9663,N_9512);
or UO_1226 (O_1226,N_9850,N_9821);
nor UO_1227 (O_1227,N_9934,N_9520);
and UO_1228 (O_1228,N_9993,N_9906);
nor UO_1229 (O_1229,N_9511,N_9737);
or UO_1230 (O_1230,N_9866,N_9598);
xor UO_1231 (O_1231,N_9662,N_9939);
or UO_1232 (O_1232,N_9847,N_9523);
nand UO_1233 (O_1233,N_9517,N_9816);
and UO_1234 (O_1234,N_9556,N_9849);
nand UO_1235 (O_1235,N_9930,N_9704);
xor UO_1236 (O_1236,N_9955,N_9572);
nor UO_1237 (O_1237,N_9520,N_9527);
nor UO_1238 (O_1238,N_9598,N_9927);
or UO_1239 (O_1239,N_9791,N_9990);
nor UO_1240 (O_1240,N_9524,N_9633);
nor UO_1241 (O_1241,N_9637,N_9838);
or UO_1242 (O_1242,N_9517,N_9960);
xor UO_1243 (O_1243,N_9773,N_9736);
nor UO_1244 (O_1244,N_9592,N_9605);
xnor UO_1245 (O_1245,N_9895,N_9695);
and UO_1246 (O_1246,N_9938,N_9832);
xor UO_1247 (O_1247,N_9560,N_9638);
nand UO_1248 (O_1248,N_9927,N_9591);
xnor UO_1249 (O_1249,N_9992,N_9644);
or UO_1250 (O_1250,N_9566,N_9767);
nand UO_1251 (O_1251,N_9993,N_9540);
and UO_1252 (O_1252,N_9831,N_9596);
and UO_1253 (O_1253,N_9548,N_9512);
nand UO_1254 (O_1254,N_9943,N_9695);
or UO_1255 (O_1255,N_9805,N_9721);
xor UO_1256 (O_1256,N_9615,N_9935);
or UO_1257 (O_1257,N_9797,N_9553);
nand UO_1258 (O_1258,N_9601,N_9864);
xnor UO_1259 (O_1259,N_9637,N_9540);
nor UO_1260 (O_1260,N_9623,N_9661);
nor UO_1261 (O_1261,N_9917,N_9797);
nand UO_1262 (O_1262,N_9711,N_9818);
xor UO_1263 (O_1263,N_9872,N_9542);
or UO_1264 (O_1264,N_9915,N_9840);
or UO_1265 (O_1265,N_9709,N_9565);
or UO_1266 (O_1266,N_9743,N_9614);
or UO_1267 (O_1267,N_9699,N_9630);
nor UO_1268 (O_1268,N_9976,N_9505);
xor UO_1269 (O_1269,N_9524,N_9899);
nand UO_1270 (O_1270,N_9833,N_9605);
xor UO_1271 (O_1271,N_9998,N_9502);
or UO_1272 (O_1272,N_9531,N_9900);
xor UO_1273 (O_1273,N_9684,N_9556);
and UO_1274 (O_1274,N_9951,N_9798);
or UO_1275 (O_1275,N_9715,N_9726);
or UO_1276 (O_1276,N_9952,N_9654);
and UO_1277 (O_1277,N_9999,N_9656);
or UO_1278 (O_1278,N_9513,N_9906);
xor UO_1279 (O_1279,N_9603,N_9941);
xor UO_1280 (O_1280,N_9875,N_9651);
and UO_1281 (O_1281,N_9953,N_9507);
nand UO_1282 (O_1282,N_9527,N_9974);
and UO_1283 (O_1283,N_9552,N_9664);
and UO_1284 (O_1284,N_9888,N_9995);
nor UO_1285 (O_1285,N_9604,N_9669);
xor UO_1286 (O_1286,N_9916,N_9982);
nand UO_1287 (O_1287,N_9501,N_9526);
nand UO_1288 (O_1288,N_9784,N_9913);
and UO_1289 (O_1289,N_9896,N_9560);
nor UO_1290 (O_1290,N_9987,N_9692);
xnor UO_1291 (O_1291,N_9738,N_9842);
nand UO_1292 (O_1292,N_9681,N_9723);
nand UO_1293 (O_1293,N_9593,N_9879);
nand UO_1294 (O_1294,N_9819,N_9580);
nand UO_1295 (O_1295,N_9962,N_9758);
nand UO_1296 (O_1296,N_9970,N_9991);
xnor UO_1297 (O_1297,N_9526,N_9757);
or UO_1298 (O_1298,N_9991,N_9688);
or UO_1299 (O_1299,N_9983,N_9897);
nand UO_1300 (O_1300,N_9578,N_9922);
nand UO_1301 (O_1301,N_9555,N_9611);
nand UO_1302 (O_1302,N_9534,N_9972);
nand UO_1303 (O_1303,N_9771,N_9724);
nand UO_1304 (O_1304,N_9531,N_9641);
nor UO_1305 (O_1305,N_9848,N_9599);
or UO_1306 (O_1306,N_9524,N_9990);
nand UO_1307 (O_1307,N_9557,N_9792);
xnor UO_1308 (O_1308,N_9588,N_9712);
or UO_1309 (O_1309,N_9676,N_9500);
nand UO_1310 (O_1310,N_9975,N_9553);
nand UO_1311 (O_1311,N_9824,N_9800);
nand UO_1312 (O_1312,N_9686,N_9928);
or UO_1313 (O_1313,N_9713,N_9882);
or UO_1314 (O_1314,N_9816,N_9960);
nand UO_1315 (O_1315,N_9523,N_9684);
xor UO_1316 (O_1316,N_9654,N_9749);
nand UO_1317 (O_1317,N_9637,N_9645);
xnor UO_1318 (O_1318,N_9546,N_9580);
or UO_1319 (O_1319,N_9784,N_9535);
nor UO_1320 (O_1320,N_9993,N_9784);
and UO_1321 (O_1321,N_9970,N_9691);
nor UO_1322 (O_1322,N_9931,N_9731);
nor UO_1323 (O_1323,N_9863,N_9533);
and UO_1324 (O_1324,N_9700,N_9601);
nor UO_1325 (O_1325,N_9911,N_9689);
and UO_1326 (O_1326,N_9554,N_9810);
and UO_1327 (O_1327,N_9818,N_9546);
or UO_1328 (O_1328,N_9604,N_9960);
nor UO_1329 (O_1329,N_9577,N_9664);
nor UO_1330 (O_1330,N_9778,N_9541);
nand UO_1331 (O_1331,N_9720,N_9953);
and UO_1332 (O_1332,N_9804,N_9575);
nor UO_1333 (O_1333,N_9958,N_9556);
or UO_1334 (O_1334,N_9994,N_9659);
nor UO_1335 (O_1335,N_9769,N_9643);
nand UO_1336 (O_1336,N_9563,N_9658);
or UO_1337 (O_1337,N_9686,N_9930);
and UO_1338 (O_1338,N_9986,N_9688);
or UO_1339 (O_1339,N_9658,N_9794);
or UO_1340 (O_1340,N_9838,N_9902);
nand UO_1341 (O_1341,N_9519,N_9503);
or UO_1342 (O_1342,N_9573,N_9955);
or UO_1343 (O_1343,N_9539,N_9696);
nand UO_1344 (O_1344,N_9926,N_9807);
nor UO_1345 (O_1345,N_9955,N_9833);
and UO_1346 (O_1346,N_9874,N_9606);
nand UO_1347 (O_1347,N_9531,N_9517);
nor UO_1348 (O_1348,N_9880,N_9687);
nand UO_1349 (O_1349,N_9727,N_9507);
nand UO_1350 (O_1350,N_9739,N_9525);
and UO_1351 (O_1351,N_9512,N_9773);
and UO_1352 (O_1352,N_9541,N_9834);
and UO_1353 (O_1353,N_9723,N_9971);
xnor UO_1354 (O_1354,N_9999,N_9521);
and UO_1355 (O_1355,N_9547,N_9807);
xnor UO_1356 (O_1356,N_9936,N_9660);
and UO_1357 (O_1357,N_9720,N_9807);
nor UO_1358 (O_1358,N_9503,N_9938);
nand UO_1359 (O_1359,N_9835,N_9922);
nor UO_1360 (O_1360,N_9547,N_9509);
xnor UO_1361 (O_1361,N_9655,N_9980);
or UO_1362 (O_1362,N_9736,N_9741);
or UO_1363 (O_1363,N_9726,N_9658);
xor UO_1364 (O_1364,N_9919,N_9772);
xor UO_1365 (O_1365,N_9950,N_9506);
nand UO_1366 (O_1366,N_9908,N_9904);
and UO_1367 (O_1367,N_9504,N_9517);
or UO_1368 (O_1368,N_9955,N_9634);
and UO_1369 (O_1369,N_9711,N_9694);
nor UO_1370 (O_1370,N_9605,N_9682);
or UO_1371 (O_1371,N_9565,N_9942);
or UO_1372 (O_1372,N_9510,N_9618);
and UO_1373 (O_1373,N_9547,N_9532);
and UO_1374 (O_1374,N_9694,N_9831);
and UO_1375 (O_1375,N_9762,N_9750);
nand UO_1376 (O_1376,N_9841,N_9845);
xor UO_1377 (O_1377,N_9958,N_9751);
xor UO_1378 (O_1378,N_9642,N_9936);
xnor UO_1379 (O_1379,N_9749,N_9589);
or UO_1380 (O_1380,N_9698,N_9963);
nand UO_1381 (O_1381,N_9736,N_9687);
nand UO_1382 (O_1382,N_9990,N_9512);
or UO_1383 (O_1383,N_9814,N_9722);
nand UO_1384 (O_1384,N_9560,N_9705);
nand UO_1385 (O_1385,N_9597,N_9906);
nor UO_1386 (O_1386,N_9508,N_9621);
or UO_1387 (O_1387,N_9781,N_9546);
or UO_1388 (O_1388,N_9689,N_9550);
nand UO_1389 (O_1389,N_9725,N_9635);
nor UO_1390 (O_1390,N_9554,N_9857);
nand UO_1391 (O_1391,N_9735,N_9640);
or UO_1392 (O_1392,N_9539,N_9762);
nand UO_1393 (O_1393,N_9569,N_9686);
nor UO_1394 (O_1394,N_9757,N_9927);
and UO_1395 (O_1395,N_9934,N_9551);
and UO_1396 (O_1396,N_9860,N_9998);
nor UO_1397 (O_1397,N_9827,N_9973);
or UO_1398 (O_1398,N_9547,N_9538);
and UO_1399 (O_1399,N_9807,N_9613);
and UO_1400 (O_1400,N_9786,N_9687);
and UO_1401 (O_1401,N_9656,N_9745);
nor UO_1402 (O_1402,N_9909,N_9791);
and UO_1403 (O_1403,N_9984,N_9812);
xnor UO_1404 (O_1404,N_9761,N_9857);
xor UO_1405 (O_1405,N_9628,N_9952);
nand UO_1406 (O_1406,N_9579,N_9723);
and UO_1407 (O_1407,N_9996,N_9777);
nor UO_1408 (O_1408,N_9732,N_9556);
nor UO_1409 (O_1409,N_9660,N_9525);
xor UO_1410 (O_1410,N_9758,N_9933);
or UO_1411 (O_1411,N_9562,N_9645);
and UO_1412 (O_1412,N_9580,N_9997);
and UO_1413 (O_1413,N_9716,N_9964);
and UO_1414 (O_1414,N_9522,N_9792);
or UO_1415 (O_1415,N_9671,N_9579);
nor UO_1416 (O_1416,N_9571,N_9550);
or UO_1417 (O_1417,N_9853,N_9748);
nand UO_1418 (O_1418,N_9776,N_9583);
nand UO_1419 (O_1419,N_9580,N_9860);
xnor UO_1420 (O_1420,N_9924,N_9855);
nand UO_1421 (O_1421,N_9829,N_9702);
nor UO_1422 (O_1422,N_9672,N_9541);
nor UO_1423 (O_1423,N_9554,N_9875);
or UO_1424 (O_1424,N_9927,N_9923);
xor UO_1425 (O_1425,N_9730,N_9642);
nand UO_1426 (O_1426,N_9872,N_9547);
and UO_1427 (O_1427,N_9683,N_9755);
nand UO_1428 (O_1428,N_9931,N_9953);
xnor UO_1429 (O_1429,N_9517,N_9651);
nor UO_1430 (O_1430,N_9978,N_9776);
or UO_1431 (O_1431,N_9845,N_9523);
nand UO_1432 (O_1432,N_9645,N_9819);
nor UO_1433 (O_1433,N_9635,N_9637);
nor UO_1434 (O_1434,N_9800,N_9740);
xnor UO_1435 (O_1435,N_9706,N_9755);
xor UO_1436 (O_1436,N_9608,N_9978);
or UO_1437 (O_1437,N_9981,N_9550);
xnor UO_1438 (O_1438,N_9668,N_9546);
or UO_1439 (O_1439,N_9699,N_9756);
nand UO_1440 (O_1440,N_9872,N_9821);
and UO_1441 (O_1441,N_9604,N_9552);
and UO_1442 (O_1442,N_9730,N_9515);
nor UO_1443 (O_1443,N_9845,N_9952);
nor UO_1444 (O_1444,N_9530,N_9592);
nor UO_1445 (O_1445,N_9505,N_9913);
or UO_1446 (O_1446,N_9990,N_9522);
nand UO_1447 (O_1447,N_9527,N_9587);
or UO_1448 (O_1448,N_9841,N_9834);
nor UO_1449 (O_1449,N_9795,N_9622);
and UO_1450 (O_1450,N_9966,N_9825);
nor UO_1451 (O_1451,N_9802,N_9885);
nand UO_1452 (O_1452,N_9718,N_9721);
nand UO_1453 (O_1453,N_9814,N_9599);
and UO_1454 (O_1454,N_9639,N_9948);
nand UO_1455 (O_1455,N_9826,N_9753);
nand UO_1456 (O_1456,N_9585,N_9557);
nor UO_1457 (O_1457,N_9810,N_9869);
and UO_1458 (O_1458,N_9650,N_9605);
xnor UO_1459 (O_1459,N_9522,N_9769);
nand UO_1460 (O_1460,N_9943,N_9705);
or UO_1461 (O_1461,N_9754,N_9549);
nand UO_1462 (O_1462,N_9832,N_9511);
xnor UO_1463 (O_1463,N_9629,N_9859);
or UO_1464 (O_1464,N_9800,N_9607);
nor UO_1465 (O_1465,N_9892,N_9936);
nor UO_1466 (O_1466,N_9991,N_9517);
xnor UO_1467 (O_1467,N_9860,N_9890);
nor UO_1468 (O_1468,N_9990,N_9875);
nand UO_1469 (O_1469,N_9500,N_9968);
nand UO_1470 (O_1470,N_9818,N_9802);
xor UO_1471 (O_1471,N_9641,N_9579);
nor UO_1472 (O_1472,N_9563,N_9586);
nand UO_1473 (O_1473,N_9815,N_9600);
nand UO_1474 (O_1474,N_9862,N_9928);
nand UO_1475 (O_1475,N_9553,N_9667);
xor UO_1476 (O_1476,N_9675,N_9797);
or UO_1477 (O_1477,N_9604,N_9666);
and UO_1478 (O_1478,N_9815,N_9621);
or UO_1479 (O_1479,N_9589,N_9572);
xor UO_1480 (O_1480,N_9649,N_9635);
nand UO_1481 (O_1481,N_9594,N_9977);
xnor UO_1482 (O_1482,N_9918,N_9763);
and UO_1483 (O_1483,N_9777,N_9889);
xnor UO_1484 (O_1484,N_9714,N_9597);
and UO_1485 (O_1485,N_9834,N_9783);
nor UO_1486 (O_1486,N_9945,N_9937);
nor UO_1487 (O_1487,N_9581,N_9993);
and UO_1488 (O_1488,N_9594,N_9876);
nor UO_1489 (O_1489,N_9884,N_9573);
nand UO_1490 (O_1490,N_9662,N_9929);
xor UO_1491 (O_1491,N_9800,N_9928);
nor UO_1492 (O_1492,N_9558,N_9536);
and UO_1493 (O_1493,N_9644,N_9979);
and UO_1494 (O_1494,N_9881,N_9605);
and UO_1495 (O_1495,N_9644,N_9762);
nand UO_1496 (O_1496,N_9895,N_9906);
nor UO_1497 (O_1497,N_9914,N_9836);
nor UO_1498 (O_1498,N_9852,N_9529);
or UO_1499 (O_1499,N_9777,N_9705);
endmodule