module basic_1000_10000_1500_20_levels_2xor_2(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999;
nor U0 (N_0,In_50,In_221);
or U1 (N_1,In_808,In_832);
and U2 (N_2,In_799,In_260);
or U3 (N_3,In_560,In_711);
nand U4 (N_4,In_175,In_914);
or U5 (N_5,In_98,In_220);
nand U6 (N_6,In_358,In_860);
or U7 (N_7,In_971,In_74);
nor U8 (N_8,In_253,In_844);
and U9 (N_9,In_536,In_399);
or U10 (N_10,In_198,In_369);
and U11 (N_11,In_575,In_847);
nand U12 (N_12,In_161,In_514);
xor U13 (N_13,In_697,In_783);
and U14 (N_14,In_73,In_280);
nand U15 (N_15,In_194,In_292);
nor U16 (N_16,In_972,In_347);
and U17 (N_17,In_484,In_945);
nor U18 (N_18,In_479,In_499);
or U19 (N_19,In_123,In_275);
or U20 (N_20,In_142,In_355);
nor U21 (N_21,In_254,In_295);
and U22 (N_22,In_871,In_249);
nand U23 (N_23,In_384,In_821);
nand U24 (N_24,In_563,In_430);
and U25 (N_25,In_931,In_215);
or U26 (N_26,In_473,In_163);
nand U27 (N_27,In_731,In_354);
nand U28 (N_28,In_174,In_265);
xor U29 (N_29,In_848,In_995);
or U30 (N_30,In_24,In_680);
nor U31 (N_31,In_736,In_495);
nor U32 (N_32,In_827,In_489);
nand U33 (N_33,In_330,In_466);
and U34 (N_34,In_624,In_77);
nor U35 (N_35,In_264,In_956);
and U36 (N_36,In_283,In_468);
xnor U37 (N_37,In_587,In_35);
and U38 (N_38,In_471,In_781);
nand U39 (N_39,In_531,In_81);
or U40 (N_40,In_78,In_303);
nand U41 (N_41,In_352,In_1);
nand U42 (N_42,In_792,In_704);
and U43 (N_43,In_884,In_107);
and U44 (N_44,In_177,In_322);
nand U45 (N_45,In_753,In_338);
nand U46 (N_46,In_869,In_777);
nor U47 (N_47,In_565,In_447);
nand U48 (N_48,In_502,In_544);
and U49 (N_49,In_239,In_444);
and U50 (N_50,In_814,In_651);
nand U51 (N_51,In_452,In_41);
and U52 (N_52,In_294,In_729);
xnor U53 (N_53,In_831,In_888);
and U54 (N_54,In_771,In_515);
nand U55 (N_55,In_698,In_682);
nor U56 (N_56,In_877,In_183);
nor U57 (N_57,In_569,In_719);
nor U58 (N_58,In_402,In_478);
or U59 (N_59,In_897,In_291);
xor U60 (N_60,In_141,In_297);
nand U61 (N_61,In_806,In_703);
or U62 (N_62,In_820,In_327);
nor U63 (N_63,In_333,In_969);
nor U64 (N_64,In_755,In_258);
or U65 (N_65,In_532,In_638);
or U66 (N_66,In_613,In_159);
or U67 (N_67,In_597,In_273);
and U68 (N_68,In_342,In_760);
nand U69 (N_69,In_718,In_454);
or U70 (N_70,In_158,In_930);
nor U71 (N_71,In_51,In_817);
xnor U72 (N_72,In_964,In_193);
nor U73 (N_73,In_679,In_615);
nand U74 (N_74,In_356,In_100);
nand U75 (N_75,In_395,In_812);
and U76 (N_76,In_708,In_789);
nand U77 (N_77,In_106,In_86);
nand U78 (N_78,In_405,In_689);
nor U79 (N_79,In_534,In_735);
and U80 (N_80,In_385,In_951);
nand U81 (N_81,In_893,In_339);
nand U82 (N_82,In_379,In_111);
nand U83 (N_83,In_721,In_5);
and U84 (N_84,In_334,In_92);
nand U85 (N_85,In_132,In_419);
nor U86 (N_86,In_448,In_632);
nor U87 (N_87,In_881,In_400);
and U88 (N_88,In_629,In_293);
nand U89 (N_89,In_285,In_653);
xnor U90 (N_90,In_568,In_64);
or U91 (N_91,In_887,In_125);
nor U92 (N_92,In_391,In_701);
nand U93 (N_93,In_166,In_612);
nor U94 (N_94,In_657,In_620);
nand U95 (N_95,In_313,In_171);
nand U96 (N_96,In_747,In_553);
or U97 (N_97,In_639,In_407);
or U98 (N_98,In_938,In_700);
nor U99 (N_99,In_255,In_925);
nor U100 (N_100,In_117,In_187);
or U101 (N_101,In_909,In_833);
nor U102 (N_102,In_943,In_242);
nor U103 (N_103,In_192,In_97);
and U104 (N_104,In_59,In_683);
or U105 (N_105,In_501,In_199);
nor U106 (N_106,In_218,In_717);
or U107 (N_107,In_602,In_907);
nand U108 (N_108,In_2,In_247);
nor U109 (N_109,In_415,In_101);
nand U110 (N_110,In_904,In_486);
or U111 (N_111,In_427,In_761);
nor U112 (N_112,In_655,In_425);
nand U113 (N_113,In_169,In_866);
nor U114 (N_114,In_900,In_139);
or U115 (N_115,In_661,In_337);
xor U116 (N_116,In_750,In_883);
nand U117 (N_117,In_197,In_482);
and U118 (N_118,In_195,In_234);
nand U119 (N_119,In_189,In_593);
or U120 (N_120,In_541,In_367);
or U121 (N_121,In_397,In_380);
nand U122 (N_122,In_941,In_607);
nand U123 (N_123,In_540,In_66);
or U124 (N_124,In_965,In_228);
nand U125 (N_125,In_115,In_674);
nand U126 (N_126,In_572,In_745);
and U127 (N_127,In_456,In_811);
or U128 (N_128,In_326,In_362);
nand U129 (N_129,In_867,In_702);
nor U130 (N_130,In_967,In_937);
nand U131 (N_131,In_80,In_667);
nor U132 (N_132,In_574,In_598);
nand U133 (N_133,In_609,In_469);
nand U134 (N_134,In_923,In_852);
nand U135 (N_135,In_374,In_759);
nand U136 (N_136,In_76,In_691);
nor U137 (N_137,In_627,In_672);
or U138 (N_138,In_329,In_591);
nor U139 (N_139,In_105,In_987);
nor U140 (N_140,In_626,In_270);
or U141 (N_141,In_699,In_3);
nand U142 (N_142,In_918,In_188);
and U143 (N_143,In_126,In_858);
nand U144 (N_144,In_782,In_984);
and U145 (N_145,In_710,In_850);
and U146 (N_146,In_446,In_91);
nor U147 (N_147,In_252,In_770);
and U148 (N_148,In_631,In_670);
or U149 (N_149,In_418,In_509);
nand U150 (N_150,In_842,In_716);
nor U151 (N_151,In_511,In_480);
and U152 (N_152,In_17,In_746);
nand U153 (N_153,In_768,In_20);
nor U154 (N_154,In_343,In_641);
or U155 (N_155,In_288,In_325);
xor U156 (N_156,In_185,In_955);
and U157 (N_157,In_633,In_944);
or U158 (N_158,In_10,In_491);
nor U159 (N_159,In_774,In_723);
nand U160 (N_160,In_70,In_611);
and U161 (N_161,In_26,In_411);
nand U162 (N_162,In_776,In_829);
nor U163 (N_163,In_894,In_304);
and U164 (N_164,In_131,In_772);
xor U165 (N_165,In_335,In_530);
and U166 (N_166,In_421,In_919);
and U167 (N_167,In_201,In_619);
or U168 (N_168,In_147,In_44);
nand U169 (N_169,In_580,In_826);
nand U170 (N_170,In_960,In_251);
or U171 (N_171,In_998,In_715);
and U172 (N_172,In_975,In_173);
nand U173 (N_173,In_88,In_610);
or U174 (N_174,In_289,In_27);
nor U175 (N_175,In_18,In_233);
and U176 (N_176,In_500,In_835);
nor U177 (N_177,In_140,In_879);
nor U178 (N_178,In_259,In_567);
nand U179 (N_179,In_706,In_589);
and U180 (N_180,In_310,In_604);
or U181 (N_181,In_460,In_566);
nand U182 (N_182,In_982,In_642);
or U183 (N_183,In_301,In_219);
or U184 (N_184,In_94,In_467);
nor U185 (N_185,In_980,In_529);
and U186 (N_186,In_578,In_526);
nor U187 (N_187,In_459,In_836);
nor U188 (N_188,In_726,In_796);
nand U189 (N_189,In_896,In_451);
nor U190 (N_190,In_744,In_913);
nand U191 (N_191,In_905,In_660);
nor U192 (N_192,In_241,In_742);
or U193 (N_193,In_124,In_316);
nor U194 (N_194,In_784,In_29);
nor U195 (N_195,In_788,In_924);
and U196 (N_196,In_45,In_227);
nand U197 (N_197,In_681,In_992);
and U198 (N_198,In_908,In_226);
nand U199 (N_199,In_84,In_794);
or U200 (N_200,In_396,In_722);
nor U201 (N_201,In_331,In_705);
nor U202 (N_202,In_517,In_961);
xnor U203 (N_203,In_733,In_190);
xnor U204 (N_204,In_538,In_49);
nand U205 (N_205,In_780,In_802);
nand U206 (N_206,In_42,In_637);
nor U207 (N_207,In_217,In_312);
nor U208 (N_208,In_96,In_581);
and U209 (N_209,In_263,In_378);
and U210 (N_210,In_245,In_898);
or U211 (N_211,In_947,In_351);
or U212 (N_212,In_795,In_516);
or U213 (N_213,In_953,In_790);
nor U214 (N_214,In_562,In_773);
nor U215 (N_215,In_693,In_52);
nand U216 (N_216,In_599,In_696);
nand U217 (N_217,In_184,In_548);
xor U218 (N_218,In_109,In_144);
nand U219 (N_219,In_63,In_841);
nand U220 (N_220,In_90,In_886);
nand U221 (N_221,In_431,In_861);
nor U222 (N_222,In_122,In_320);
nor U223 (N_223,In_546,In_623);
nand U224 (N_224,In_487,In_170);
or U225 (N_225,In_481,In_819);
and U226 (N_226,In_590,In_475);
or U227 (N_227,In_791,In_628);
nand U228 (N_228,In_856,In_207);
and U229 (N_229,In_527,In_954);
and U230 (N_230,In_970,In_377);
nand U231 (N_231,In_853,In_864);
and U232 (N_232,In_146,In_839);
or U233 (N_233,In_53,In_506);
and U234 (N_234,In_749,In_855);
nor U235 (N_235,In_424,In_143);
nor U236 (N_236,In_68,In_981);
xnor U237 (N_237,In_859,In_976);
xor U238 (N_238,In_818,In_991);
nand U239 (N_239,In_116,In_155);
and U240 (N_240,In_640,In_151);
nor U241 (N_241,In_804,In_82);
nand U242 (N_242,In_916,In_55);
nand U243 (N_243,In_205,In_934);
nand U244 (N_244,In_878,In_19);
or U245 (N_245,In_110,In_461);
and U246 (N_246,In_556,In_603);
or U247 (N_247,In_420,In_994);
nor U248 (N_248,In_974,In_805);
and U249 (N_249,In_360,In_618);
nand U250 (N_250,In_318,In_868);
or U251 (N_251,In_150,In_307);
nor U252 (N_252,In_462,In_305);
nand U253 (N_253,In_644,In_47);
nand U254 (N_254,In_436,In_872);
and U255 (N_255,In_959,In_349);
nand U256 (N_256,In_838,In_413);
and U257 (N_257,In_57,In_72);
or U258 (N_258,In_39,In_341);
and U259 (N_259,In_714,In_738);
nand U260 (N_260,In_102,In_204);
and U261 (N_261,In_528,In_373);
and U262 (N_262,In_211,In_523);
and U263 (N_263,In_936,In_551);
and U264 (N_264,In_649,In_137);
and U265 (N_265,In_634,In_825);
nor U266 (N_266,In_282,In_157);
or U267 (N_267,In_389,In_267);
or U268 (N_268,In_135,In_752);
nand U269 (N_269,In_366,In_686);
or U270 (N_270,In_164,In_748);
nand U271 (N_271,In_659,In_963);
or U272 (N_272,In_727,In_793);
or U273 (N_273,In_12,In_375);
nor U274 (N_274,In_685,In_797);
or U275 (N_275,In_906,In_206);
nor U276 (N_276,In_200,In_21);
nand U277 (N_277,In_33,In_62);
nand U278 (N_278,In_939,In_845);
and U279 (N_279,In_261,In_350);
nor U280 (N_280,In_596,In_186);
nand U281 (N_281,In_977,In_635);
or U282 (N_282,In_180,In_892);
nor U283 (N_283,In_690,In_988);
nor U284 (N_284,In_741,In_669);
or U285 (N_285,In_160,In_594);
nor U286 (N_286,In_915,In_584);
nor U287 (N_287,In_743,In_483);
and U288 (N_288,In_429,In_688);
and U289 (N_289,In_223,In_554);
and U290 (N_290,In_668,In_296);
or U291 (N_291,In_966,In_321);
and U292 (N_292,In_309,In_724);
or U293 (N_293,In_570,In_406);
nand U294 (N_294,In_231,In_404);
or U295 (N_295,In_940,In_388);
nand U296 (N_296,In_208,In_889);
and U297 (N_297,In_588,In_266);
or U298 (N_298,In_248,In_778);
nor U299 (N_299,In_903,In_393);
and U300 (N_300,In_364,In_525);
nand U301 (N_301,In_910,In_558);
nand U302 (N_302,In_559,In_435);
nor U303 (N_303,In_809,In_497);
nand U304 (N_304,In_785,In_300);
or U305 (N_305,In_465,In_537);
nor U306 (N_306,In_48,In_917);
or U307 (N_307,In_9,In_764);
xor U308 (N_308,In_32,In_621);
and U309 (N_309,In_348,In_154);
nor U310 (N_310,In_663,In_692);
and U311 (N_311,In_93,In_948);
nor U312 (N_312,In_87,In_127);
nand U313 (N_313,In_636,In_95);
and U314 (N_314,In_216,In_687);
and U315 (N_315,In_196,In_758);
or U316 (N_316,In_46,In_958);
or U317 (N_317,In_911,In_875);
nand U318 (N_318,In_803,In_646);
or U319 (N_319,In_237,In_6);
nand U320 (N_320,In_608,In_815);
or U321 (N_321,In_614,In_665);
nand U322 (N_322,In_235,In_457);
and U323 (N_323,In_230,In_181);
nor U324 (N_324,In_561,In_571);
and U325 (N_325,In_153,In_176);
nor U326 (N_326,In_824,In_214);
or U327 (N_327,In_165,In_455);
and U328 (N_328,In_973,In_268);
or U329 (N_329,In_576,In_328);
nand U330 (N_330,In_394,In_108);
nand U331 (N_331,In_156,In_863);
and U332 (N_332,In_440,In_524);
nor U333 (N_333,In_800,In_392);
nand U334 (N_334,In_645,In_13);
or U335 (N_335,In_210,In_315);
and U336 (N_336,In_134,In_450);
nor U337 (N_337,In_786,In_408);
or U338 (N_338,In_573,In_225);
nor U339 (N_339,In_23,In_762);
and U340 (N_340,In_43,In_775);
nand U341 (N_341,In_503,In_376);
or U342 (N_342,In_922,In_179);
nor U343 (N_343,In_178,In_324);
nand U344 (N_344,In_119,In_658);
and U345 (N_345,In_191,In_854);
nand U346 (N_346,In_549,In_85);
xnor U347 (N_347,In_895,In_891);
or U348 (N_348,In_485,In_209);
or U349 (N_349,In_99,In_224);
nor U350 (N_350,In_993,In_946);
and U351 (N_351,In_458,In_387);
nor U352 (N_352,In_279,In_314);
nand U353 (N_353,In_383,In_779);
nor U354 (N_354,In_290,In_422);
nand U355 (N_355,In_999,In_65);
nand U356 (N_356,In_577,In_488);
and U357 (N_357,In_508,In_595);
nor U358 (N_358,In_353,In_694);
xor U359 (N_359,In_601,In_932);
xnor U360 (N_360,In_823,In_662);
and U361 (N_361,In_656,In_882);
nor U362 (N_362,In_535,In_521);
nor U363 (N_363,In_510,In_433);
nand U364 (N_364,In_464,In_432);
and U365 (N_365,In_308,In_920);
nand U366 (N_366,In_250,In_287);
and U367 (N_367,In_606,In_807);
or U368 (N_368,In_370,In_363);
and U369 (N_369,In_345,In_121);
and U370 (N_370,In_732,In_512);
nand U371 (N_371,In_410,In_162);
or U372 (N_372,In_707,In_767);
nand U373 (N_373,In_401,In_822);
nand U374 (N_374,In_298,In_311);
nand U375 (N_375,In_149,In_582);
nand U376 (N_376,In_985,In_0);
xor U377 (N_377,In_262,In_996);
or U378 (N_378,In_31,In_625);
nor U379 (N_379,In_403,In_751);
and U380 (N_380,In_368,In_713);
nand U381 (N_381,In_921,In_890);
or U382 (N_382,In_552,In_678);
nor U383 (N_383,In_720,In_677);
and U384 (N_384,In_880,In_89);
nor U385 (N_385,In_272,In_494);
nand U386 (N_386,In_118,In_409);
and U387 (N_387,In_622,In_453);
nor U388 (N_388,In_129,In_650);
and U389 (N_389,In_332,In_664);
and U390 (N_390,In_145,In_935);
and U391 (N_391,In_498,In_167);
and U392 (N_392,In_490,In_968);
nand U393 (N_393,In_676,In_357);
or U394 (N_394,In_256,In_439);
nand U395 (N_395,In_182,In_801);
and U396 (N_396,In_361,In_238);
or U397 (N_397,In_885,In_257);
or U398 (N_398,In_952,In_417);
or U399 (N_399,In_426,In_7);
nor U400 (N_400,In_695,In_605);
and U401 (N_401,In_477,In_507);
nand U402 (N_402,In_843,In_128);
or U403 (N_403,In_445,In_929);
and U404 (N_404,In_386,In_928);
or U405 (N_405,In_876,In_269);
nor U406 (N_406,In_449,In_986);
and U407 (N_407,In_274,In_840);
nor U408 (N_408,In_412,In_104);
xnor U409 (N_409,In_550,In_505);
or U410 (N_410,In_133,In_438);
nor U411 (N_411,In_236,In_203);
nand U412 (N_412,In_202,In_319);
nand U413 (N_413,In_754,In_120);
and U414 (N_414,In_654,In_666);
nand U415 (N_415,In_933,In_281);
nand U416 (N_416,In_585,In_229);
and U417 (N_417,In_152,In_730);
nor U418 (N_418,In_849,In_712);
nand U419 (N_419,In_583,In_284);
and U420 (N_420,In_671,In_302);
nor U421 (N_421,In_390,In_130);
nor U422 (N_422,In_504,In_949);
xnor U423 (N_423,In_851,In_901);
nand U424 (N_424,In_564,In_617);
nand U425 (N_425,In_15,In_492);
or U426 (N_426,In_912,In_37);
and U427 (N_427,In_513,In_58);
or U428 (N_428,In_979,In_4);
nand U429 (N_429,In_398,In_728);
and U430 (N_430,In_336,In_846);
and U431 (N_431,In_428,In_865);
nor U432 (N_432,In_616,In_519);
xnor U433 (N_433,In_114,In_71);
nand U434 (N_434,In_243,In_103);
and U435 (N_435,In_543,In_962);
nand U436 (N_436,In_725,In_278);
nand U437 (N_437,In_600,In_8);
or U438 (N_438,In_763,In_11);
or U439 (N_439,In_518,In_830);
and U440 (N_440,In_942,In_34);
and U441 (N_441,In_899,In_212);
and U442 (N_442,In_56,In_816);
or U443 (N_443,In_359,In_28);
or U444 (N_444,In_902,In_522);
xnor U445 (N_445,In_276,In_113);
and U446 (N_446,In_244,In_22);
nand U447 (N_447,In_926,In_927);
nor U448 (N_448,In_734,In_739);
or U449 (N_449,In_168,In_246);
nor U450 (N_450,In_54,In_539);
and U451 (N_451,In_957,In_533);
nand U452 (N_452,In_75,In_810);
nor U453 (N_453,In_240,In_470);
or U454 (N_454,In_989,In_557);
nor U455 (N_455,In_766,In_474);
nor U456 (N_456,In_813,In_769);
nand U457 (N_457,In_40,In_340);
or U458 (N_458,In_673,In_675);
or U459 (N_459,In_441,In_870);
and U460 (N_460,In_647,In_496);
and U461 (N_461,In_547,In_472);
nor U462 (N_462,In_873,In_67);
nor U463 (N_463,In_950,In_434);
and U464 (N_464,In_30,In_148);
or U465 (N_465,In_382,In_643);
or U466 (N_466,In_317,In_38);
nand U467 (N_467,In_765,In_542);
and U468 (N_468,In_787,In_323);
and U469 (N_469,In_592,In_112);
or U470 (N_470,In_443,In_586);
nor U471 (N_471,In_463,In_493);
or U472 (N_472,In_442,In_83);
or U473 (N_473,In_416,In_16);
and U474 (N_474,In_346,In_61);
nor U475 (N_475,In_737,In_306);
and U476 (N_476,In_286,In_277);
nor U477 (N_477,In_648,In_740);
nand U478 (N_478,In_213,In_983);
nand U479 (N_479,In_857,In_372);
nand U480 (N_480,In_136,In_14);
or U481 (N_481,In_60,In_299);
nor U482 (N_482,In_997,In_25);
and U483 (N_483,In_138,In_232);
nand U484 (N_484,In_990,In_371);
and U485 (N_485,In_684,In_545);
or U486 (N_486,In_555,In_172);
nand U487 (N_487,In_271,In_579);
and U488 (N_488,In_874,In_798);
and U489 (N_489,In_978,In_834);
or U490 (N_490,In_520,In_828);
and U491 (N_491,In_630,In_79);
and U492 (N_492,In_414,In_652);
or U493 (N_493,In_709,In_36);
nand U494 (N_494,In_344,In_381);
nand U495 (N_495,In_757,In_437);
or U496 (N_496,In_69,In_756);
nand U497 (N_497,In_476,In_862);
xnor U498 (N_498,In_837,In_423);
and U499 (N_499,In_222,In_365);
nand U500 (N_500,N_448,N_29);
or U501 (N_501,N_151,N_98);
nor U502 (N_502,N_10,N_325);
nor U503 (N_503,N_335,N_281);
and U504 (N_504,N_252,N_407);
nor U505 (N_505,N_282,N_232);
nand U506 (N_506,N_78,N_422);
or U507 (N_507,N_189,N_50);
or U508 (N_508,N_376,N_226);
nor U509 (N_509,N_323,N_87);
nor U510 (N_510,N_466,N_334);
nand U511 (N_511,N_75,N_249);
and U512 (N_512,N_479,N_165);
xor U513 (N_513,N_289,N_357);
nor U514 (N_514,N_305,N_264);
or U515 (N_515,N_168,N_431);
nor U516 (N_516,N_337,N_438);
or U517 (N_517,N_480,N_33);
or U518 (N_518,N_248,N_359);
nand U519 (N_519,N_457,N_172);
or U520 (N_520,N_6,N_313);
or U521 (N_521,N_434,N_76);
and U522 (N_522,N_403,N_452);
nand U523 (N_523,N_352,N_474);
nor U524 (N_524,N_51,N_208);
nor U525 (N_525,N_294,N_327);
nor U526 (N_526,N_418,N_231);
and U527 (N_527,N_336,N_306);
nand U528 (N_528,N_175,N_136);
nand U529 (N_529,N_284,N_303);
nor U530 (N_530,N_21,N_495);
or U531 (N_531,N_94,N_242);
or U532 (N_532,N_465,N_401);
and U533 (N_533,N_52,N_421);
and U534 (N_534,N_430,N_370);
nor U535 (N_535,N_372,N_30);
or U536 (N_536,N_131,N_103);
nor U537 (N_537,N_406,N_222);
xor U538 (N_538,N_490,N_395);
or U539 (N_539,N_214,N_298);
nor U540 (N_540,N_258,N_144);
nand U541 (N_541,N_365,N_227);
nand U542 (N_542,N_229,N_114);
or U543 (N_543,N_130,N_183);
nor U544 (N_544,N_2,N_170);
or U545 (N_545,N_262,N_476);
and U546 (N_546,N_410,N_106);
and U547 (N_547,N_110,N_148);
nor U548 (N_548,N_246,N_485);
or U549 (N_549,N_216,N_13);
nor U550 (N_550,N_290,N_363);
or U551 (N_551,N_489,N_177);
or U552 (N_552,N_55,N_54);
or U553 (N_553,N_269,N_204);
or U554 (N_554,N_125,N_414);
or U555 (N_555,N_176,N_219);
or U556 (N_556,N_478,N_20);
nand U557 (N_557,N_169,N_424);
nor U558 (N_558,N_429,N_455);
nor U559 (N_559,N_192,N_350);
and U560 (N_560,N_161,N_321);
nor U561 (N_561,N_201,N_283);
nor U562 (N_562,N_446,N_74);
or U563 (N_563,N_251,N_35);
or U564 (N_564,N_259,N_80);
nor U565 (N_565,N_211,N_0);
nand U566 (N_566,N_362,N_358);
xor U567 (N_567,N_42,N_18);
nor U568 (N_568,N_253,N_326);
and U569 (N_569,N_400,N_330);
nor U570 (N_570,N_353,N_344);
nor U571 (N_571,N_3,N_271);
nor U572 (N_572,N_188,N_387);
nand U573 (N_573,N_311,N_193);
nor U574 (N_574,N_63,N_237);
and U575 (N_575,N_482,N_364);
and U576 (N_576,N_300,N_408);
and U577 (N_577,N_27,N_36);
nor U578 (N_578,N_8,N_383);
and U579 (N_579,N_276,N_375);
or U580 (N_580,N_447,N_243);
nor U581 (N_581,N_159,N_149);
or U582 (N_582,N_469,N_77);
and U583 (N_583,N_164,N_32);
nand U584 (N_584,N_142,N_435);
nand U585 (N_585,N_411,N_171);
and U586 (N_586,N_346,N_312);
or U587 (N_587,N_113,N_109);
or U588 (N_588,N_166,N_292);
or U589 (N_589,N_184,N_461);
or U590 (N_590,N_467,N_484);
nor U591 (N_591,N_349,N_266);
nand U592 (N_592,N_121,N_296);
xor U593 (N_593,N_156,N_389);
nand U594 (N_594,N_318,N_450);
and U595 (N_595,N_128,N_45);
nor U596 (N_596,N_380,N_118);
or U597 (N_597,N_157,N_49);
nor U598 (N_598,N_138,N_56);
and U599 (N_599,N_409,N_268);
and U600 (N_600,N_5,N_162);
nand U601 (N_601,N_320,N_388);
nand U602 (N_602,N_198,N_210);
nor U603 (N_603,N_57,N_16);
or U604 (N_604,N_417,N_345);
and U605 (N_605,N_1,N_101);
nand U606 (N_606,N_412,N_302);
or U607 (N_607,N_65,N_378);
nor U608 (N_608,N_355,N_356);
nand U609 (N_609,N_37,N_493);
nor U610 (N_610,N_270,N_93);
and U611 (N_611,N_58,N_212);
nor U612 (N_612,N_487,N_293);
or U613 (N_613,N_333,N_158);
or U614 (N_614,N_471,N_154);
and U615 (N_615,N_316,N_497);
or U616 (N_616,N_426,N_133);
nand U617 (N_617,N_89,N_381);
nand U618 (N_618,N_100,N_153);
nor U619 (N_619,N_404,N_126);
nand U620 (N_620,N_69,N_197);
and U621 (N_621,N_245,N_265);
nand U622 (N_622,N_397,N_419);
or U623 (N_623,N_129,N_343);
xor U624 (N_624,N_41,N_234);
nor U625 (N_625,N_483,N_339);
nand U626 (N_626,N_230,N_44);
nand U627 (N_627,N_119,N_40);
nand U628 (N_628,N_132,N_235);
and U629 (N_629,N_205,N_371);
nor U630 (N_630,N_239,N_348);
and U631 (N_631,N_286,N_396);
nand U632 (N_632,N_143,N_39);
nand U633 (N_633,N_472,N_297);
or U634 (N_634,N_97,N_64);
and U635 (N_635,N_67,N_202);
and U636 (N_636,N_117,N_386);
or U637 (N_637,N_458,N_111);
or U638 (N_638,N_31,N_445);
nand U639 (N_639,N_468,N_360);
or U640 (N_640,N_152,N_307);
or U641 (N_641,N_374,N_477);
nand U642 (N_642,N_317,N_280);
nor U643 (N_643,N_427,N_108);
and U644 (N_644,N_92,N_498);
or U645 (N_645,N_213,N_134);
or U646 (N_646,N_444,N_393);
or U647 (N_647,N_60,N_390);
nor U648 (N_648,N_81,N_66);
nor U649 (N_649,N_274,N_104);
or U650 (N_650,N_25,N_53);
and U651 (N_651,N_377,N_279);
and U652 (N_652,N_443,N_382);
or U653 (N_653,N_361,N_432);
nor U654 (N_654,N_309,N_272);
nand U655 (N_655,N_217,N_491);
nor U656 (N_656,N_405,N_34);
and U657 (N_657,N_373,N_451);
xnor U658 (N_658,N_43,N_181);
nor U659 (N_659,N_199,N_299);
and U660 (N_660,N_285,N_494);
nand U661 (N_661,N_354,N_225);
nor U662 (N_662,N_191,N_90);
or U663 (N_663,N_23,N_185);
nand U664 (N_664,N_102,N_449);
nor U665 (N_665,N_62,N_72);
nand U666 (N_666,N_241,N_220);
nor U667 (N_667,N_398,N_347);
or U668 (N_668,N_70,N_112);
and U669 (N_669,N_462,N_261);
or U670 (N_670,N_394,N_203);
or U671 (N_671,N_24,N_442);
xor U672 (N_672,N_250,N_460);
xor U673 (N_673,N_470,N_291);
and U674 (N_674,N_79,N_392);
and U675 (N_675,N_137,N_123);
nor U676 (N_676,N_145,N_86);
nor U677 (N_677,N_304,N_486);
or U678 (N_678,N_182,N_423);
nand U679 (N_679,N_47,N_464);
and U680 (N_680,N_351,N_174);
nand U681 (N_681,N_329,N_140);
nand U682 (N_682,N_319,N_341);
or U683 (N_683,N_221,N_496);
nand U684 (N_684,N_116,N_322);
xor U685 (N_685,N_207,N_420);
nor U686 (N_686,N_278,N_186);
nand U687 (N_687,N_218,N_11);
or U688 (N_688,N_328,N_187);
nor U689 (N_689,N_425,N_342);
nor U690 (N_690,N_499,N_84);
nor U691 (N_691,N_332,N_15);
nand U692 (N_692,N_88,N_135);
or U693 (N_693,N_155,N_436);
nand U694 (N_694,N_415,N_340);
or U695 (N_695,N_275,N_238);
or U696 (N_696,N_4,N_331);
and U697 (N_697,N_301,N_295);
nand U698 (N_698,N_247,N_463);
or U699 (N_699,N_399,N_96);
nand U700 (N_700,N_173,N_141);
and U701 (N_701,N_223,N_456);
and U702 (N_702,N_273,N_475);
and U703 (N_703,N_38,N_209);
nand U704 (N_704,N_59,N_163);
or U705 (N_705,N_26,N_146);
or U706 (N_706,N_402,N_194);
or U707 (N_707,N_139,N_7);
or U708 (N_708,N_83,N_481);
and U709 (N_709,N_190,N_260);
nand U710 (N_710,N_473,N_179);
nor U711 (N_711,N_308,N_180);
nand U712 (N_712,N_196,N_367);
nor U713 (N_713,N_256,N_385);
and U714 (N_714,N_206,N_384);
and U715 (N_715,N_9,N_195);
and U716 (N_716,N_107,N_488);
nor U717 (N_717,N_228,N_46);
or U718 (N_718,N_277,N_105);
nand U719 (N_719,N_254,N_91);
or U720 (N_720,N_459,N_122);
and U721 (N_721,N_22,N_437);
nor U722 (N_722,N_17,N_310);
or U723 (N_723,N_366,N_127);
nor U724 (N_724,N_492,N_267);
or U725 (N_725,N_120,N_288);
nor U726 (N_726,N_233,N_236);
nand U727 (N_727,N_224,N_95);
nand U728 (N_728,N_453,N_379);
nand U729 (N_729,N_315,N_12);
and U730 (N_730,N_255,N_73);
nand U731 (N_731,N_440,N_150);
nand U732 (N_732,N_240,N_28);
nor U733 (N_733,N_257,N_48);
nand U734 (N_734,N_433,N_82);
and U735 (N_735,N_416,N_338);
nand U736 (N_736,N_19,N_314);
and U737 (N_737,N_85,N_147);
or U738 (N_738,N_454,N_160);
and U739 (N_739,N_391,N_287);
or U740 (N_740,N_368,N_215);
and U741 (N_741,N_124,N_244);
nand U742 (N_742,N_115,N_439);
nand U743 (N_743,N_263,N_68);
nand U744 (N_744,N_167,N_14);
nor U745 (N_745,N_324,N_369);
or U746 (N_746,N_61,N_200);
nand U747 (N_747,N_99,N_71);
xnor U748 (N_748,N_428,N_441);
nand U749 (N_749,N_413,N_178);
or U750 (N_750,N_208,N_158);
and U751 (N_751,N_410,N_307);
nand U752 (N_752,N_393,N_196);
or U753 (N_753,N_403,N_224);
or U754 (N_754,N_280,N_403);
nand U755 (N_755,N_143,N_190);
nand U756 (N_756,N_59,N_264);
and U757 (N_757,N_107,N_21);
or U758 (N_758,N_446,N_496);
nor U759 (N_759,N_386,N_166);
nand U760 (N_760,N_149,N_160);
or U761 (N_761,N_276,N_70);
and U762 (N_762,N_229,N_204);
nand U763 (N_763,N_441,N_454);
and U764 (N_764,N_186,N_184);
nor U765 (N_765,N_5,N_202);
or U766 (N_766,N_486,N_147);
and U767 (N_767,N_177,N_352);
nand U768 (N_768,N_490,N_230);
nand U769 (N_769,N_127,N_431);
or U770 (N_770,N_208,N_495);
or U771 (N_771,N_246,N_476);
and U772 (N_772,N_417,N_246);
nand U773 (N_773,N_266,N_393);
and U774 (N_774,N_281,N_164);
and U775 (N_775,N_443,N_15);
nand U776 (N_776,N_267,N_352);
nand U777 (N_777,N_75,N_425);
nand U778 (N_778,N_450,N_355);
or U779 (N_779,N_360,N_211);
nand U780 (N_780,N_125,N_266);
nor U781 (N_781,N_443,N_417);
nor U782 (N_782,N_0,N_303);
nand U783 (N_783,N_121,N_383);
nor U784 (N_784,N_133,N_237);
or U785 (N_785,N_334,N_108);
and U786 (N_786,N_425,N_245);
nand U787 (N_787,N_79,N_460);
nand U788 (N_788,N_185,N_468);
nor U789 (N_789,N_138,N_455);
and U790 (N_790,N_165,N_120);
or U791 (N_791,N_9,N_391);
nor U792 (N_792,N_338,N_395);
and U793 (N_793,N_403,N_211);
nand U794 (N_794,N_116,N_264);
nand U795 (N_795,N_75,N_44);
xor U796 (N_796,N_119,N_397);
or U797 (N_797,N_389,N_179);
nor U798 (N_798,N_160,N_190);
xor U799 (N_799,N_412,N_75);
or U800 (N_800,N_371,N_28);
and U801 (N_801,N_102,N_357);
and U802 (N_802,N_22,N_162);
or U803 (N_803,N_173,N_197);
or U804 (N_804,N_230,N_211);
and U805 (N_805,N_463,N_89);
nor U806 (N_806,N_198,N_333);
nor U807 (N_807,N_95,N_126);
nor U808 (N_808,N_108,N_351);
and U809 (N_809,N_310,N_55);
or U810 (N_810,N_318,N_238);
nor U811 (N_811,N_421,N_53);
and U812 (N_812,N_345,N_462);
nand U813 (N_813,N_333,N_489);
or U814 (N_814,N_469,N_420);
xnor U815 (N_815,N_460,N_46);
or U816 (N_816,N_380,N_322);
nand U817 (N_817,N_87,N_380);
or U818 (N_818,N_387,N_374);
or U819 (N_819,N_351,N_379);
nand U820 (N_820,N_351,N_382);
and U821 (N_821,N_371,N_320);
and U822 (N_822,N_252,N_108);
and U823 (N_823,N_215,N_140);
nor U824 (N_824,N_101,N_371);
or U825 (N_825,N_124,N_213);
nand U826 (N_826,N_189,N_88);
or U827 (N_827,N_140,N_391);
nor U828 (N_828,N_58,N_365);
or U829 (N_829,N_374,N_51);
xnor U830 (N_830,N_258,N_351);
or U831 (N_831,N_54,N_118);
and U832 (N_832,N_342,N_63);
and U833 (N_833,N_49,N_239);
and U834 (N_834,N_269,N_253);
or U835 (N_835,N_180,N_227);
and U836 (N_836,N_91,N_67);
or U837 (N_837,N_173,N_230);
nand U838 (N_838,N_383,N_397);
and U839 (N_839,N_390,N_95);
nor U840 (N_840,N_8,N_260);
nand U841 (N_841,N_344,N_429);
nor U842 (N_842,N_154,N_137);
nor U843 (N_843,N_495,N_439);
xor U844 (N_844,N_420,N_363);
and U845 (N_845,N_225,N_448);
nand U846 (N_846,N_456,N_230);
or U847 (N_847,N_489,N_16);
or U848 (N_848,N_84,N_49);
nand U849 (N_849,N_463,N_230);
and U850 (N_850,N_356,N_76);
and U851 (N_851,N_116,N_338);
and U852 (N_852,N_384,N_359);
nor U853 (N_853,N_348,N_393);
nand U854 (N_854,N_186,N_376);
and U855 (N_855,N_237,N_440);
nand U856 (N_856,N_321,N_186);
nor U857 (N_857,N_251,N_163);
and U858 (N_858,N_6,N_328);
or U859 (N_859,N_470,N_40);
and U860 (N_860,N_407,N_116);
and U861 (N_861,N_184,N_79);
and U862 (N_862,N_85,N_278);
and U863 (N_863,N_40,N_494);
nor U864 (N_864,N_144,N_63);
nand U865 (N_865,N_449,N_7);
and U866 (N_866,N_357,N_86);
xor U867 (N_867,N_121,N_281);
or U868 (N_868,N_35,N_341);
and U869 (N_869,N_129,N_331);
and U870 (N_870,N_233,N_181);
and U871 (N_871,N_119,N_90);
and U872 (N_872,N_178,N_446);
nor U873 (N_873,N_430,N_26);
or U874 (N_874,N_474,N_392);
and U875 (N_875,N_60,N_243);
nor U876 (N_876,N_381,N_411);
and U877 (N_877,N_120,N_97);
or U878 (N_878,N_498,N_206);
nand U879 (N_879,N_48,N_180);
nand U880 (N_880,N_249,N_410);
nor U881 (N_881,N_320,N_118);
nor U882 (N_882,N_9,N_143);
or U883 (N_883,N_298,N_354);
nor U884 (N_884,N_318,N_433);
nor U885 (N_885,N_94,N_378);
nor U886 (N_886,N_453,N_459);
or U887 (N_887,N_20,N_90);
nand U888 (N_888,N_236,N_419);
or U889 (N_889,N_319,N_144);
or U890 (N_890,N_235,N_284);
nand U891 (N_891,N_76,N_137);
nand U892 (N_892,N_189,N_421);
nor U893 (N_893,N_89,N_212);
and U894 (N_894,N_442,N_55);
nand U895 (N_895,N_483,N_388);
and U896 (N_896,N_455,N_335);
and U897 (N_897,N_341,N_367);
or U898 (N_898,N_432,N_111);
nor U899 (N_899,N_198,N_417);
nor U900 (N_900,N_232,N_415);
nand U901 (N_901,N_324,N_498);
nand U902 (N_902,N_40,N_22);
and U903 (N_903,N_138,N_189);
nand U904 (N_904,N_499,N_468);
nand U905 (N_905,N_252,N_294);
or U906 (N_906,N_116,N_275);
nand U907 (N_907,N_248,N_286);
nor U908 (N_908,N_210,N_119);
or U909 (N_909,N_80,N_3);
and U910 (N_910,N_464,N_180);
nor U911 (N_911,N_351,N_243);
and U912 (N_912,N_247,N_349);
nand U913 (N_913,N_466,N_135);
or U914 (N_914,N_425,N_114);
or U915 (N_915,N_182,N_190);
nand U916 (N_916,N_403,N_262);
nand U917 (N_917,N_402,N_148);
or U918 (N_918,N_334,N_422);
nand U919 (N_919,N_153,N_62);
or U920 (N_920,N_67,N_361);
or U921 (N_921,N_403,N_12);
and U922 (N_922,N_20,N_381);
or U923 (N_923,N_228,N_184);
or U924 (N_924,N_63,N_436);
or U925 (N_925,N_362,N_55);
or U926 (N_926,N_5,N_477);
or U927 (N_927,N_468,N_166);
nand U928 (N_928,N_481,N_141);
nor U929 (N_929,N_377,N_214);
nand U930 (N_930,N_400,N_368);
nor U931 (N_931,N_375,N_443);
or U932 (N_932,N_404,N_320);
and U933 (N_933,N_432,N_288);
and U934 (N_934,N_307,N_398);
nor U935 (N_935,N_479,N_156);
nand U936 (N_936,N_209,N_284);
or U937 (N_937,N_314,N_492);
nand U938 (N_938,N_363,N_432);
nand U939 (N_939,N_473,N_15);
nor U940 (N_940,N_403,N_450);
or U941 (N_941,N_331,N_170);
nand U942 (N_942,N_368,N_145);
or U943 (N_943,N_429,N_362);
nand U944 (N_944,N_9,N_297);
or U945 (N_945,N_484,N_290);
nor U946 (N_946,N_425,N_367);
nor U947 (N_947,N_280,N_110);
nor U948 (N_948,N_239,N_250);
and U949 (N_949,N_164,N_86);
or U950 (N_950,N_319,N_243);
nand U951 (N_951,N_166,N_491);
nand U952 (N_952,N_445,N_0);
or U953 (N_953,N_239,N_186);
and U954 (N_954,N_436,N_407);
or U955 (N_955,N_124,N_360);
nand U956 (N_956,N_336,N_457);
nand U957 (N_957,N_222,N_28);
and U958 (N_958,N_286,N_304);
nor U959 (N_959,N_438,N_287);
or U960 (N_960,N_343,N_365);
and U961 (N_961,N_125,N_154);
or U962 (N_962,N_0,N_122);
nor U963 (N_963,N_35,N_343);
and U964 (N_964,N_1,N_472);
or U965 (N_965,N_256,N_31);
nand U966 (N_966,N_261,N_120);
and U967 (N_967,N_431,N_246);
and U968 (N_968,N_433,N_130);
xnor U969 (N_969,N_66,N_159);
and U970 (N_970,N_357,N_43);
nor U971 (N_971,N_373,N_489);
or U972 (N_972,N_495,N_291);
and U973 (N_973,N_61,N_186);
and U974 (N_974,N_390,N_96);
and U975 (N_975,N_50,N_212);
nor U976 (N_976,N_306,N_259);
or U977 (N_977,N_211,N_6);
and U978 (N_978,N_85,N_157);
nand U979 (N_979,N_455,N_74);
and U980 (N_980,N_155,N_17);
and U981 (N_981,N_314,N_283);
or U982 (N_982,N_251,N_383);
and U983 (N_983,N_249,N_357);
or U984 (N_984,N_336,N_346);
nand U985 (N_985,N_465,N_436);
or U986 (N_986,N_252,N_0);
nor U987 (N_987,N_64,N_451);
and U988 (N_988,N_211,N_229);
nand U989 (N_989,N_273,N_235);
nor U990 (N_990,N_456,N_256);
or U991 (N_991,N_170,N_229);
and U992 (N_992,N_287,N_477);
nor U993 (N_993,N_282,N_260);
xor U994 (N_994,N_177,N_472);
and U995 (N_995,N_93,N_356);
and U996 (N_996,N_301,N_139);
nand U997 (N_997,N_482,N_199);
nor U998 (N_998,N_484,N_283);
nand U999 (N_999,N_68,N_81);
xnor U1000 (N_1000,N_956,N_608);
nor U1001 (N_1001,N_706,N_880);
nor U1002 (N_1002,N_762,N_787);
or U1003 (N_1003,N_599,N_737);
or U1004 (N_1004,N_555,N_980);
nor U1005 (N_1005,N_856,N_840);
or U1006 (N_1006,N_894,N_752);
nand U1007 (N_1007,N_807,N_930);
and U1008 (N_1008,N_895,N_575);
or U1009 (N_1009,N_615,N_512);
xor U1010 (N_1010,N_743,N_636);
nand U1011 (N_1011,N_943,N_872);
or U1012 (N_1012,N_750,N_982);
nand U1013 (N_1013,N_988,N_538);
nor U1014 (N_1014,N_848,N_852);
nor U1015 (N_1015,N_849,N_885);
or U1016 (N_1016,N_686,N_514);
nand U1017 (N_1017,N_991,N_830);
and U1018 (N_1018,N_677,N_594);
xor U1019 (N_1019,N_923,N_975);
nand U1020 (N_1020,N_713,N_716);
nand U1021 (N_1021,N_959,N_875);
or U1022 (N_1022,N_727,N_712);
nand U1023 (N_1023,N_629,N_847);
nand U1024 (N_1024,N_561,N_623);
nor U1025 (N_1025,N_996,N_540);
or U1026 (N_1026,N_524,N_928);
or U1027 (N_1027,N_945,N_919);
nand U1028 (N_1028,N_854,N_559);
nor U1029 (N_1029,N_839,N_770);
xor U1030 (N_1030,N_841,N_700);
and U1031 (N_1031,N_614,N_981);
nor U1032 (N_1032,N_544,N_808);
nand U1033 (N_1033,N_979,N_970);
or U1034 (N_1034,N_595,N_501);
or U1035 (N_1035,N_523,N_925);
and U1036 (N_1036,N_796,N_661);
nand U1037 (N_1037,N_844,N_744);
and U1038 (N_1038,N_778,N_936);
or U1039 (N_1039,N_725,N_905);
or U1040 (N_1040,N_568,N_721);
nor U1041 (N_1041,N_672,N_652);
or U1042 (N_1042,N_971,N_817);
and U1043 (N_1043,N_962,N_863);
or U1044 (N_1044,N_904,N_711);
and U1045 (N_1045,N_803,N_909);
and U1046 (N_1046,N_763,N_972);
nand U1047 (N_1047,N_583,N_658);
nor U1048 (N_1048,N_992,N_676);
or U1049 (N_1049,N_751,N_809);
or U1050 (N_1050,N_704,N_550);
nor U1051 (N_1051,N_968,N_864);
nand U1052 (N_1052,N_703,N_588);
and U1053 (N_1053,N_838,N_877);
nor U1054 (N_1054,N_579,N_797);
nand U1055 (N_1055,N_846,N_696);
nor U1056 (N_1056,N_545,N_735);
nor U1057 (N_1057,N_690,N_776);
nand U1058 (N_1058,N_539,N_795);
or U1059 (N_1059,N_630,N_589);
and U1060 (N_1060,N_612,N_714);
nand U1061 (N_1061,N_887,N_946);
nand U1062 (N_1062,N_566,N_871);
or U1063 (N_1063,N_800,N_571);
or U1064 (N_1064,N_698,N_632);
and U1065 (N_1065,N_834,N_574);
and U1066 (N_1066,N_502,N_705);
and U1067 (N_1067,N_537,N_974);
or U1068 (N_1068,N_689,N_753);
nor U1069 (N_1069,N_774,N_964);
or U1070 (N_1070,N_606,N_912);
nand U1071 (N_1071,N_784,N_929);
nor U1072 (N_1072,N_626,N_892);
and U1073 (N_1073,N_679,N_738);
nor U1074 (N_1074,N_810,N_908);
or U1075 (N_1075,N_673,N_733);
and U1076 (N_1076,N_990,N_769);
or U1077 (N_1077,N_886,N_605);
or U1078 (N_1078,N_879,N_611);
nor U1079 (N_1079,N_995,N_596);
nor U1080 (N_1080,N_598,N_754);
xnor U1081 (N_1081,N_940,N_997);
and U1082 (N_1082,N_791,N_881);
or U1083 (N_1083,N_508,N_527);
xnor U1084 (N_1084,N_569,N_782);
and U1085 (N_1085,N_897,N_667);
nor U1086 (N_1086,N_899,N_507);
nand U1087 (N_1087,N_767,N_647);
nor U1088 (N_1088,N_720,N_771);
nand U1089 (N_1089,N_789,N_531);
nor U1090 (N_1090,N_656,N_828);
or U1091 (N_1091,N_509,N_586);
nand U1092 (N_1092,N_640,N_966);
nand U1093 (N_1093,N_688,N_958);
or U1094 (N_1094,N_913,N_792);
nor U1095 (N_1095,N_578,N_824);
or U1096 (N_1096,N_581,N_639);
xnor U1097 (N_1097,N_858,N_627);
xor U1098 (N_1098,N_503,N_907);
nor U1099 (N_1099,N_708,N_532);
and U1100 (N_1100,N_746,N_624);
and U1101 (N_1101,N_518,N_917);
or U1102 (N_1102,N_622,N_857);
and U1103 (N_1103,N_937,N_593);
nor U1104 (N_1104,N_790,N_853);
nand U1105 (N_1105,N_671,N_699);
and U1106 (N_1106,N_822,N_950);
or U1107 (N_1107,N_691,N_765);
nand U1108 (N_1108,N_944,N_761);
nor U1109 (N_1109,N_873,N_906);
nand U1110 (N_1110,N_963,N_707);
xnor U1111 (N_1111,N_793,N_893);
or U1112 (N_1112,N_883,N_903);
nand U1113 (N_1113,N_576,N_734);
nand U1114 (N_1114,N_526,N_603);
nand U1115 (N_1115,N_868,N_773);
nand U1116 (N_1116,N_642,N_911);
nor U1117 (N_1117,N_842,N_645);
nand U1118 (N_1118,N_729,N_674);
nand U1119 (N_1119,N_573,N_604);
nand U1120 (N_1120,N_556,N_920);
nor U1121 (N_1121,N_833,N_684);
nand U1122 (N_1122,N_914,N_542);
nand U1123 (N_1123,N_548,N_815);
nand U1124 (N_1124,N_748,N_506);
nand U1125 (N_1125,N_553,N_558);
nand U1126 (N_1126,N_916,N_653);
or U1127 (N_1127,N_513,N_643);
and U1128 (N_1128,N_620,N_654);
or U1129 (N_1129,N_898,N_775);
or U1130 (N_1130,N_938,N_866);
or U1131 (N_1131,N_695,N_924);
nor U1132 (N_1132,N_889,N_987);
nand U1133 (N_1133,N_567,N_682);
or U1134 (N_1134,N_625,N_888);
nor U1135 (N_1135,N_777,N_665);
and U1136 (N_1136,N_819,N_739);
nand U1137 (N_1137,N_504,N_836);
nor U1138 (N_1138,N_572,N_741);
or U1139 (N_1139,N_510,N_517);
or U1140 (N_1140,N_546,N_867);
or U1141 (N_1141,N_685,N_601);
or U1142 (N_1142,N_998,N_927);
nand U1143 (N_1143,N_683,N_804);
nor U1144 (N_1144,N_760,N_516);
nor U1145 (N_1145,N_755,N_780);
nor U1146 (N_1146,N_657,N_939);
nor U1147 (N_1147,N_663,N_994);
and U1148 (N_1148,N_882,N_697);
nand U1149 (N_1149,N_650,N_747);
or U1150 (N_1150,N_591,N_613);
nor U1151 (N_1151,N_659,N_745);
and U1152 (N_1152,N_814,N_635);
or U1153 (N_1153,N_687,N_560);
and U1154 (N_1154,N_977,N_818);
or U1155 (N_1155,N_715,N_655);
nand U1156 (N_1156,N_641,N_597);
or U1157 (N_1157,N_669,N_931);
or U1158 (N_1158,N_802,N_781);
and U1159 (N_1159,N_621,N_986);
or U1160 (N_1160,N_736,N_855);
nand U1161 (N_1161,N_918,N_816);
or U1162 (N_1162,N_835,N_884);
or U1163 (N_1163,N_851,N_609);
or U1164 (N_1164,N_701,N_876);
nor U1165 (N_1165,N_617,N_993);
nand U1166 (N_1166,N_585,N_941);
nand U1167 (N_1167,N_528,N_772);
nand U1168 (N_1168,N_520,N_577);
or U1169 (N_1169,N_779,N_798);
or U1170 (N_1170,N_536,N_662);
or U1171 (N_1171,N_860,N_702);
nand U1172 (N_1172,N_717,N_519);
or U1173 (N_1173,N_580,N_511);
nor U1174 (N_1174,N_607,N_983);
or U1175 (N_1175,N_633,N_610);
and U1176 (N_1176,N_718,N_955);
and U1177 (N_1177,N_709,N_949);
nand U1178 (N_1178,N_587,N_600);
nor U1179 (N_1179,N_722,N_649);
nor U1180 (N_1180,N_890,N_813);
nor U1181 (N_1181,N_823,N_989);
and U1182 (N_1182,N_680,N_935);
or U1183 (N_1183,N_845,N_843);
nand U1184 (N_1184,N_878,N_551);
nor U1185 (N_1185,N_953,N_869);
nor U1186 (N_1186,N_829,N_758);
and U1187 (N_1187,N_783,N_694);
or U1188 (N_1188,N_731,N_616);
nand U1189 (N_1189,N_522,N_666);
nor U1190 (N_1190,N_644,N_646);
or U1191 (N_1191,N_535,N_582);
nand U1192 (N_1192,N_957,N_757);
and U1193 (N_1193,N_831,N_692);
and U1194 (N_1194,N_821,N_901);
or U1195 (N_1195,N_759,N_564);
and U1196 (N_1196,N_805,N_984);
nor U1197 (N_1197,N_948,N_965);
nand U1198 (N_1198,N_732,N_549);
nor U1199 (N_1199,N_710,N_521);
or U1200 (N_1200,N_541,N_788);
or U1201 (N_1201,N_826,N_547);
and U1202 (N_1202,N_861,N_832);
or U1203 (N_1203,N_926,N_954);
nand U1204 (N_1204,N_942,N_563);
or U1205 (N_1205,N_634,N_602);
or U1206 (N_1206,N_742,N_921);
or U1207 (N_1207,N_500,N_862);
nand U1208 (N_1208,N_670,N_664);
nand U1209 (N_1209,N_973,N_902);
nand U1210 (N_1210,N_801,N_764);
nor U1211 (N_1211,N_969,N_505);
or U1212 (N_1212,N_529,N_756);
nor U1213 (N_1213,N_554,N_557);
nor U1214 (N_1214,N_515,N_749);
or U1215 (N_1215,N_719,N_806);
and U1216 (N_1216,N_900,N_590);
nor U1217 (N_1217,N_976,N_530);
and U1218 (N_1218,N_799,N_668);
nand U1219 (N_1219,N_874,N_896);
nand U1220 (N_1220,N_961,N_811);
or U1221 (N_1221,N_865,N_785);
and U1222 (N_1222,N_915,N_570);
nor U1223 (N_1223,N_543,N_681);
nor U1224 (N_1224,N_533,N_628);
or U1225 (N_1225,N_525,N_794);
and U1226 (N_1226,N_870,N_837);
nor U1227 (N_1227,N_565,N_786);
nor U1228 (N_1228,N_978,N_951);
or U1229 (N_1229,N_985,N_934);
and U1230 (N_1230,N_932,N_820);
and U1231 (N_1231,N_651,N_825);
nor U1232 (N_1232,N_859,N_584);
nor U1233 (N_1233,N_728,N_922);
nor U1234 (N_1234,N_726,N_960);
nand U1235 (N_1235,N_952,N_933);
and U1236 (N_1236,N_891,N_693);
or U1237 (N_1237,N_812,N_910);
nand U1238 (N_1238,N_619,N_827);
or U1239 (N_1239,N_740,N_631);
nand U1240 (N_1240,N_967,N_552);
nand U1241 (N_1241,N_947,N_730);
nor U1242 (N_1242,N_562,N_768);
nand U1243 (N_1243,N_648,N_618);
or U1244 (N_1244,N_660,N_850);
nor U1245 (N_1245,N_637,N_724);
nand U1246 (N_1246,N_766,N_675);
nand U1247 (N_1247,N_678,N_534);
or U1248 (N_1248,N_638,N_999);
nor U1249 (N_1249,N_723,N_592);
and U1250 (N_1250,N_609,N_809);
nand U1251 (N_1251,N_711,N_564);
nand U1252 (N_1252,N_979,N_643);
nor U1253 (N_1253,N_706,N_694);
nand U1254 (N_1254,N_888,N_652);
nor U1255 (N_1255,N_966,N_941);
nor U1256 (N_1256,N_905,N_787);
nor U1257 (N_1257,N_976,N_811);
and U1258 (N_1258,N_981,N_538);
and U1259 (N_1259,N_965,N_580);
or U1260 (N_1260,N_553,N_632);
or U1261 (N_1261,N_588,N_889);
xnor U1262 (N_1262,N_648,N_995);
nor U1263 (N_1263,N_527,N_982);
nand U1264 (N_1264,N_592,N_790);
nand U1265 (N_1265,N_652,N_682);
and U1266 (N_1266,N_757,N_947);
nor U1267 (N_1267,N_848,N_598);
and U1268 (N_1268,N_916,N_773);
nand U1269 (N_1269,N_817,N_827);
or U1270 (N_1270,N_607,N_862);
nand U1271 (N_1271,N_974,N_806);
nor U1272 (N_1272,N_919,N_839);
nand U1273 (N_1273,N_576,N_699);
or U1274 (N_1274,N_750,N_701);
nor U1275 (N_1275,N_568,N_801);
nand U1276 (N_1276,N_814,N_610);
nor U1277 (N_1277,N_554,N_809);
or U1278 (N_1278,N_858,N_747);
and U1279 (N_1279,N_533,N_666);
nor U1280 (N_1280,N_595,N_974);
nor U1281 (N_1281,N_840,N_987);
or U1282 (N_1282,N_568,N_744);
or U1283 (N_1283,N_923,N_757);
nand U1284 (N_1284,N_839,N_920);
or U1285 (N_1285,N_722,N_527);
nor U1286 (N_1286,N_722,N_511);
nor U1287 (N_1287,N_742,N_708);
or U1288 (N_1288,N_773,N_794);
and U1289 (N_1289,N_652,N_503);
and U1290 (N_1290,N_527,N_639);
nor U1291 (N_1291,N_810,N_725);
nor U1292 (N_1292,N_800,N_540);
and U1293 (N_1293,N_753,N_836);
nor U1294 (N_1294,N_975,N_516);
or U1295 (N_1295,N_738,N_681);
nand U1296 (N_1296,N_563,N_575);
and U1297 (N_1297,N_933,N_793);
and U1298 (N_1298,N_916,N_611);
nor U1299 (N_1299,N_842,N_649);
nor U1300 (N_1300,N_701,N_597);
and U1301 (N_1301,N_935,N_899);
nand U1302 (N_1302,N_616,N_596);
nor U1303 (N_1303,N_662,N_642);
nand U1304 (N_1304,N_842,N_651);
nor U1305 (N_1305,N_716,N_703);
and U1306 (N_1306,N_624,N_686);
and U1307 (N_1307,N_980,N_603);
nor U1308 (N_1308,N_992,N_767);
nand U1309 (N_1309,N_634,N_873);
xor U1310 (N_1310,N_783,N_534);
or U1311 (N_1311,N_646,N_564);
or U1312 (N_1312,N_572,N_658);
and U1313 (N_1313,N_520,N_867);
or U1314 (N_1314,N_825,N_876);
nor U1315 (N_1315,N_512,N_957);
xnor U1316 (N_1316,N_591,N_766);
nand U1317 (N_1317,N_919,N_918);
and U1318 (N_1318,N_652,N_829);
or U1319 (N_1319,N_515,N_733);
and U1320 (N_1320,N_745,N_931);
and U1321 (N_1321,N_607,N_854);
and U1322 (N_1322,N_758,N_927);
nand U1323 (N_1323,N_765,N_757);
or U1324 (N_1324,N_913,N_911);
or U1325 (N_1325,N_677,N_509);
and U1326 (N_1326,N_624,N_984);
nand U1327 (N_1327,N_858,N_899);
nand U1328 (N_1328,N_611,N_563);
nor U1329 (N_1329,N_809,N_511);
nor U1330 (N_1330,N_921,N_600);
and U1331 (N_1331,N_734,N_546);
or U1332 (N_1332,N_600,N_937);
nand U1333 (N_1333,N_676,N_860);
nor U1334 (N_1334,N_862,N_825);
nor U1335 (N_1335,N_915,N_828);
nor U1336 (N_1336,N_527,N_885);
and U1337 (N_1337,N_904,N_573);
or U1338 (N_1338,N_910,N_717);
nand U1339 (N_1339,N_733,N_556);
and U1340 (N_1340,N_605,N_789);
or U1341 (N_1341,N_896,N_990);
and U1342 (N_1342,N_575,N_875);
nor U1343 (N_1343,N_711,N_842);
and U1344 (N_1344,N_632,N_923);
and U1345 (N_1345,N_969,N_904);
or U1346 (N_1346,N_601,N_688);
and U1347 (N_1347,N_971,N_991);
nor U1348 (N_1348,N_542,N_960);
nand U1349 (N_1349,N_819,N_815);
or U1350 (N_1350,N_723,N_839);
nor U1351 (N_1351,N_601,N_801);
nor U1352 (N_1352,N_794,N_915);
and U1353 (N_1353,N_581,N_902);
or U1354 (N_1354,N_980,N_885);
nand U1355 (N_1355,N_604,N_685);
nand U1356 (N_1356,N_552,N_512);
or U1357 (N_1357,N_743,N_976);
nand U1358 (N_1358,N_740,N_911);
nand U1359 (N_1359,N_636,N_672);
and U1360 (N_1360,N_571,N_694);
nand U1361 (N_1361,N_751,N_652);
or U1362 (N_1362,N_644,N_592);
nand U1363 (N_1363,N_967,N_559);
or U1364 (N_1364,N_956,N_930);
nor U1365 (N_1365,N_550,N_887);
xor U1366 (N_1366,N_903,N_562);
nand U1367 (N_1367,N_661,N_699);
nor U1368 (N_1368,N_787,N_504);
or U1369 (N_1369,N_504,N_861);
nor U1370 (N_1370,N_972,N_907);
or U1371 (N_1371,N_790,N_604);
nor U1372 (N_1372,N_854,N_683);
and U1373 (N_1373,N_812,N_921);
or U1374 (N_1374,N_778,N_634);
or U1375 (N_1375,N_998,N_556);
xor U1376 (N_1376,N_637,N_828);
or U1377 (N_1377,N_889,N_674);
nor U1378 (N_1378,N_593,N_573);
or U1379 (N_1379,N_618,N_890);
and U1380 (N_1380,N_920,N_540);
or U1381 (N_1381,N_669,N_930);
nor U1382 (N_1382,N_570,N_533);
nor U1383 (N_1383,N_506,N_746);
or U1384 (N_1384,N_740,N_866);
nand U1385 (N_1385,N_665,N_516);
nor U1386 (N_1386,N_751,N_708);
nand U1387 (N_1387,N_882,N_514);
or U1388 (N_1388,N_657,N_960);
nor U1389 (N_1389,N_735,N_947);
xnor U1390 (N_1390,N_966,N_511);
nor U1391 (N_1391,N_844,N_901);
or U1392 (N_1392,N_607,N_608);
or U1393 (N_1393,N_562,N_783);
nand U1394 (N_1394,N_713,N_820);
nor U1395 (N_1395,N_606,N_805);
nand U1396 (N_1396,N_626,N_761);
or U1397 (N_1397,N_572,N_655);
nand U1398 (N_1398,N_596,N_529);
and U1399 (N_1399,N_990,N_814);
or U1400 (N_1400,N_927,N_878);
nor U1401 (N_1401,N_813,N_752);
nor U1402 (N_1402,N_502,N_678);
nor U1403 (N_1403,N_669,N_912);
and U1404 (N_1404,N_685,N_933);
or U1405 (N_1405,N_862,N_695);
or U1406 (N_1406,N_876,N_607);
nor U1407 (N_1407,N_512,N_804);
nand U1408 (N_1408,N_786,N_723);
nor U1409 (N_1409,N_794,N_654);
and U1410 (N_1410,N_622,N_885);
nand U1411 (N_1411,N_566,N_805);
nand U1412 (N_1412,N_932,N_878);
nand U1413 (N_1413,N_852,N_517);
nand U1414 (N_1414,N_859,N_720);
and U1415 (N_1415,N_618,N_636);
nand U1416 (N_1416,N_866,N_655);
or U1417 (N_1417,N_860,N_552);
xor U1418 (N_1418,N_657,N_975);
xor U1419 (N_1419,N_509,N_934);
nor U1420 (N_1420,N_618,N_614);
nand U1421 (N_1421,N_948,N_656);
or U1422 (N_1422,N_860,N_839);
nor U1423 (N_1423,N_824,N_571);
and U1424 (N_1424,N_568,N_745);
and U1425 (N_1425,N_975,N_728);
and U1426 (N_1426,N_983,N_552);
nand U1427 (N_1427,N_658,N_764);
nor U1428 (N_1428,N_835,N_656);
or U1429 (N_1429,N_847,N_916);
nor U1430 (N_1430,N_851,N_651);
nor U1431 (N_1431,N_928,N_975);
nor U1432 (N_1432,N_726,N_734);
nor U1433 (N_1433,N_936,N_662);
or U1434 (N_1434,N_935,N_715);
or U1435 (N_1435,N_581,N_575);
nand U1436 (N_1436,N_904,N_886);
or U1437 (N_1437,N_778,N_602);
nor U1438 (N_1438,N_966,N_655);
and U1439 (N_1439,N_739,N_701);
nand U1440 (N_1440,N_701,N_543);
and U1441 (N_1441,N_826,N_950);
and U1442 (N_1442,N_694,N_954);
nor U1443 (N_1443,N_580,N_928);
nand U1444 (N_1444,N_706,N_594);
and U1445 (N_1445,N_906,N_637);
nand U1446 (N_1446,N_697,N_537);
and U1447 (N_1447,N_722,N_711);
nor U1448 (N_1448,N_755,N_591);
or U1449 (N_1449,N_623,N_819);
and U1450 (N_1450,N_870,N_748);
nor U1451 (N_1451,N_771,N_511);
nand U1452 (N_1452,N_687,N_723);
or U1453 (N_1453,N_687,N_604);
nand U1454 (N_1454,N_825,N_739);
and U1455 (N_1455,N_668,N_695);
nor U1456 (N_1456,N_929,N_736);
nor U1457 (N_1457,N_533,N_921);
or U1458 (N_1458,N_538,N_946);
and U1459 (N_1459,N_540,N_738);
and U1460 (N_1460,N_995,N_542);
or U1461 (N_1461,N_699,N_692);
nand U1462 (N_1462,N_547,N_843);
or U1463 (N_1463,N_529,N_590);
and U1464 (N_1464,N_545,N_994);
nand U1465 (N_1465,N_638,N_796);
nand U1466 (N_1466,N_755,N_714);
and U1467 (N_1467,N_595,N_848);
nand U1468 (N_1468,N_863,N_650);
xnor U1469 (N_1469,N_799,N_765);
or U1470 (N_1470,N_517,N_888);
nand U1471 (N_1471,N_837,N_674);
nand U1472 (N_1472,N_862,N_975);
and U1473 (N_1473,N_894,N_927);
nor U1474 (N_1474,N_841,N_958);
nor U1475 (N_1475,N_919,N_772);
and U1476 (N_1476,N_949,N_733);
nor U1477 (N_1477,N_591,N_749);
or U1478 (N_1478,N_754,N_607);
nor U1479 (N_1479,N_655,N_574);
or U1480 (N_1480,N_840,N_728);
nand U1481 (N_1481,N_538,N_768);
or U1482 (N_1482,N_631,N_775);
nor U1483 (N_1483,N_523,N_555);
and U1484 (N_1484,N_654,N_993);
nand U1485 (N_1485,N_870,N_620);
nand U1486 (N_1486,N_554,N_902);
nand U1487 (N_1487,N_885,N_997);
or U1488 (N_1488,N_700,N_647);
nand U1489 (N_1489,N_631,N_820);
nor U1490 (N_1490,N_980,N_534);
and U1491 (N_1491,N_607,N_618);
and U1492 (N_1492,N_954,N_896);
or U1493 (N_1493,N_525,N_624);
nor U1494 (N_1494,N_511,N_817);
nand U1495 (N_1495,N_815,N_818);
nand U1496 (N_1496,N_612,N_782);
and U1497 (N_1497,N_801,N_966);
xnor U1498 (N_1498,N_975,N_808);
or U1499 (N_1499,N_872,N_715);
or U1500 (N_1500,N_1059,N_1493);
nand U1501 (N_1501,N_1464,N_1311);
nand U1502 (N_1502,N_1370,N_1488);
nor U1503 (N_1503,N_1112,N_1271);
and U1504 (N_1504,N_1149,N_1000);
and U1505 (N_1505,N_1086,N_1301);
nand U1506 (N_1506,N_1003,N_1489);
nor U1507 (N_1507,N_1126,N_1344);
nand U1508 (N_1508,N_1241,N_1165);
nor U1509 (N_1509,N_1440,N_1342);
xnor U1510 (N_1510,N_1247,N_1103);
nor U1511 (N_1511,N_1083,N_1025);
nor U1512 (N_1512,N_1033,N_1049);
and U1513 (N_1513,N_1379,N_1145);
nor U1514 (N_1514,N_1360,N_1334);
or U1515 (N_1515,N_1436,N_1220);
and U1516 (N_1516,N_1016,N_1499);
nand U1517 (N_1517,N_1321,N_1391);
nand U1518 (N_1518,N_1261,N_1434);
nand U1519 (N_1519,N_1482,N_1082);
nor U1520 (N_1520,N_1067,N_1189);
and U1521 (N_1521,N_1209,N_1029);
nand U1522 (N_1522,N_1309,N_1166);
nor U1523 (N_1523,N_1208,N_1120);
or U1524 (N_1524,N_1286,N_1280);
and U1525 (N_1525,N_1007,N_1066);
or U1526 (N_1526,N_1069,N_1054);
nand U1527 (N_1527,N_1310,N_1032);
nor U1528 (N_1528,N_1131,N_1398);
or U1529 (N_1529,N_1390,N_1161);
and U1530 (N_1530,N_1384,N_1143);
and U1531 (N_1531,N_1432,N_1445);
or U1532 (N_1532,N_1352,N_1496);
or U1533 (N_1533,N_1117,N_1195);
nand U1534 (N_1534,N_1463,N_1410);
or U1535 (N_1535,N_1084,N_1290);
and U1536 (N_1536,N_1037,N_1315);
xnor U1537 (N_1537,N_1106,N_1147);
xnor U1538 (N_1538,N_1284,N_1018);
or U1539 (N_1539,N_1475,N_1369);
nor U1540 (N_1540,N_1402,N_1154);
or U1541 (N_1541,N_1134,N_1444);
nor U1542 (N_1542,N_1420,N_1047);
nand U1543 (N_1543,N_1164,N_1468);
nand U1544 (N_1544,N_1326,N_1486);
nand U1545 (N_1545,N_1275,N_1171);
nand U1546 (N_1546,N_1413,N_1480);
nand U1547 (N_1547,N_1130,N_1108);
nand U1548 (N_1548,N_1462,N_1122);
nor U1549 (N_1549,N_1495,N_1196);
nor U1550 (N_1550,N_1257,N_1385);
and U1551 (N_1551,N_1021,N_1023);
and U1552 (N_1552,N_1438,N_1074);
and U1553 (N_1553,N_1065,N_1456);
xnor U1554 (N_1554,N_1393,N_1332);
or U1555 (N_1555,N_1291,N_1467);
nand U1556 (N_1556,N_1098,N_1242);
or U1557 (N_1557,N_1300,N_1197);
or U1558 (N_1558,N_1124,N_1179);
nand U1559 (N_1559,N_1478,N_1279);
nor U1560 (N_1560,N_1494,N_1399);
and U1561 (N_1561,N_1357,N_1135);
and U1562 (N_1562,N_1061,N_1203);
nor U1563 (N_1563,N_1243,N_1210);
nand U1564 (N_1564,N_1153,N_1036);
or U1565 (N_1565,N_1019,N_1157);
nor U1566 (N_1566,N_1027,N_1328);
or U1567 (N_1567,N_1417,N_1090);
nand U1568 (N_1568,N_1050,N_1364);
nor U1569 (N_1569,N_1115,N_1471);
or U1570 (N_1570,N_1362,N_1485);
or U1571 (N_1571,N_1324,N_1176);
and U1572 (N_1572,N_1312,N_1233);
or U1573 (N_1573,N_1336,N_1389);
nor U1574 (N_1574,N_1017,N_1407);
and U1575 (N_1575,N_1356,N_1093);
nand U1576 (N_1576,N_1296,N_1162);
or U1577 (N_1577,N_1015,N_1237);
or U1578 (N_1578,N_1193,N_1238);
and U1579 (N_1579,N_1483,N_1221);
xnor U1580 (N_1580,N_1139,N_1278);
or U1581 (N_1581,N_1219,N_1451);
and U1582 (N_1582,N_1313,N_1425);
nand U1583 (N_1583,N_1298,N_1064);
nand U1584 (N_1584,N_1335,N_1151);
nand U1585 (N_1585,N_1454,N_1028);
nand U1586 (N_1586,N_1405,N_1097);
nor U1587 (N_1587,N_1381,N_1319);
nor U1588 (N_1588,N_1186,N_1116);
and U1589 (N_1589,N_1392,N_1226);
nand U1590 (N_1590,N_1258,N_1387);
nand U1591 (N_1591,N_1129,N_1394);
nand U1592 (N_1592,N_1026,N_1079);
or U1593 (N_1593,N_1285,N_1492);
or U1594 (N_1594,N_1232,N_1331);
and U1595 (N_1595,N_1373,N_1272);
or U1596 (N_1596,N_1293,N_1401);
nand U1597 (N_1597,N_1371,N_1188);
or U1598 (N_1598,N_1100,N_1452);
nor U1599 (N_1599,N_1148,N_1449);
or U1600 (N_1600,N_1138,N_1376);
or U1601 (N_1601,N_1046,N_1395);
nand U1602 (N_1602,N_1076,N_1170);
and U1603 (N_1603,N_1002,N_1031);
or U1604 (N_1604,N_1366,N_1424);
xor U1605 (N_1605,N_1088,N_1141);
and U1606 (N_1606,N_1472,N_1294);
and U1607 (N_1607,N_1338,N_1078);
and U1608 (N_1608,N_1206,N_1118);
or U1609 (N_1609,N_1034,N_1288);
or U1610 (N_1610,N_1248,N_1253);
nor U1611 (N_1611,N_1024,N_1109);
and U1612 (N_1612,N_1256,N_1137);
and U1613 (N_1613,N_1460,N_1001);
or U1614 (N_1614,N_1412,N_1419);
nor U1615 (N_1615,N_1234,N_1068);
and U1616 (N_1616,N_1222,N_1388);
nand U1617 (N_1617,N_1156,N_1457);
nand U1618 (N_1618,N_1330,N_1128);
nand U1619 (N_1619,N_1265,N_1406);
and U1620 (N_1620,N_1022,N_1400);
or U1621 (N_1621,N_1229,N_1358);
nand U1622 (N_1622,N_1178,N_1051);
and U1623 (N_1623,N_1240,N_1180);
nor U1624 (N_1624,N_1262,N_1063);
and U1625 (N_1625,N_1397,N_1194);
nand U1626 (N_1626,N_1473,N_1142);
and U1627 (N_1627,N_1453,N_1487);
nor U1628 (N_1628,N_1416,N_1250);
and U1629 (N_1629,N_1055,N_1191);
xor U1630 (N_1630,N_1200,N_1132);
or U1631 (N_1631,N_1375,N_1236);
nand U1632 (N_1632,N_1378,N_1269);
nand U1633 (N_1633,N_1089,N_1254);
nor U1634 (N_1634,N_1304,N_1428);
and U1635 (N_1635,N_1249,N_1213);
nor U1636 (N_1636,N_1461,N_1427);
or U1637 (N_1637,N_1008,N_1423);
or U1638 (N_1638,N_1094,N_1484);
nor U1639 (N_1639,N_1035,N_1295);
nor U1640 (N_1640,N_1264,N_1174);
or U1641 (N_1641,N_1167,N_1274);
nand U1642 (N_1642,N_1333,N_1266);
nand U1643 (N_1643,N_1433,N_1377);
or U1644 (N_1644,N_1190,N_1058);
nand U1645 (N_1645,N_1421,N_1204);
or U1646 (N_1646,N_1173,N_1125);
nor U1647 (N_1647,N_1458,N_1133);
and U1648 (N_1648,N_1070,N_1317);
nand U1649 (N_1649,N_1255,N_1207);
and U1650 (N_1650,N_1012,N_1404);
nand U1651 (N_1651,N_1305,N_1211);
nand U1652 (N_1652,N_1408,N_1235);
and U1653 (N_1653,N_1155,N_1341);
nor U1654 (N_1654,N_1396,N_1177);
and U1655 (N_1655,N_1490,N_1431);
nand U1656 (N_1656,N_1276,N_1123);
or U1657 (N_1657,N_1119,N_1216);
nor U1658 (N_1658,N_1214,N_1011);
nor U1659 (N_1659,N_1355,N_1048);
nand U1660 (N_1660,N_1056,N_1323);
nor U1661 (N_1661,N_1231,N_1325);
nand U1662 (N_1662,N_1481,N_1013);
or U1663 (N_1663,N_1185,N_1497);
or U1664 (N_1664,N_1107,N_1443);
and U1665 (N_1665,N_1367,N_1320);
nor U1666 (N_1666,N_1192,N_1072);
or U1667 (N_1667,N_1184,N_1447);
nand U1668 (N_1668,N_1096,N_1459);
and U1669 (N_1669,N_1303,N_1057);
nand U1670 (N_1670,N_1201,N_1225);
or U1671 (N_1671,N_1337,N_1409);
and U1672 (N_1672,N_1380,N_1297);
nand U1673 (N_1673,N_1365,N_1168);
and U1674 (N_1674,N_1439,N_1175);
nor U1675 (N_1675,N_1113,N_1127);
and U1676 (N_1676,N_1227,N_1415);
nand U1677 (N_1677,N_1040,N_1136);
and U1678 (N_1678,N_1349,N_1469);
and U1679 (N_1679,N_1474,N_1363);
nand U1680 (N_1680,N_1004,N_1246);
and U1681 (N_1681,N_1429,N_1006);
and U1682 (N_1682,N_1435,N_1160);
nor U1683 (N_1683,N_1307,N_1060);
or U1684 (N_1684,N_1466,N_1308);
nor U1685 (N_1685,N_1010,N_1260);
and U1686 (N_1686,N_1202,N_1092);
nand U1687 (N_1687,N_1306,N_1411);
nor U1688 (N_1688,N_1150,N_1350);
nand U1689 (N_1689,N_1374,N_1347);
nor U1690 (N_1690,N_1169,N_1386);
nand U1691 (N_1691,N_1181,N_1403);
nand U1692 (N_1692,N_1111,N_1302);
and U1693 (N_1693,N_1414,N_1372);
and U1694 (N_1694,N_1073,N_1224);
and U1695 (N_1695,N_1277,N_1292);
and U1696 (N_1696,N_1081,N_1045);
or U1697 (N_1697,N_1267,N_1442);
or U1698 (N_1698,N_1418,N_1259);
and U1699 (N_1699,N_1144,N_1251);
nor U1700 (N_1700,N_1140,N_1041);
and U1701 (N_1701,N_1270,N_1102);
nand U1702 (N_1702,N_1263,N_1455);
or U1703 (N_1703,N_1382,N_1368);
nand U1704 (N_1704,N_1239,N_1316);
xnor U1705 (N_1705,N_1062,N_1479);
nor U1706 (N_1706,N_1268,N_1446);
or U1707 (N_1707,N_1470,N_1014);
or U1708 (N_1708,N_1182,N_1383);
and U1709 (N_1709,N_1020,N_1230);
or U1710 (N_1710,N_1289,N_1318);
nor U1711 (N_1711,N_1353,N_1044);
or U1712 (N_1712,N_1085,N_1282);
and U1713 (N_1713,N_1287,N_1223);
or U1714 (N_1714,N_1101,N_1354);
nor U1715 (N_1715,N_1450,N_1077);
nand U1716 (N_1716,N_1110,N_1422);
or U1717 (N_1717,N_1075,N_1329);
and U1718 (N_1718,N_1465,N_1105);
or U1719 (N_1719,N_1114,N_1498);
nor U1720 (N_1720,N_1053,N_1322);
nand U1721 (N_1721,N_1281,N_1245);
nor U1722 (N_1722,N_1043,N_1361);
nor U1723 (N_1723,N_1158,N_1327);
and U1724 (N_1724,N_1215,N_1351);
or U1725 (N_1725,N_1039,N_1430);
or U1726 (N_1726,N_1205,N_1345);
and U1727 (N_1727,N_1009,N_1042);
nor U1728 (N_1728,N_1071,N_1340);
nor U1729 (N_1729,N_1491,N_1163);
nor U1730 (N_1730,N_1477,N_1198);
nand U1731 (N_1731,N_1228,N_1080);
and U1732 (N_1732,N_1437,N_1091);
nor U1733 (N_1733,N_1348,N_1159);
or U1734 (N_1734,N_1087,N_1172);
or U1735 (N_1735,N_1273,N_1218);
nand U1736 (N_1736,N_1252,N_1244);
nand U1737 (N_1737,N_1212,N_1448);
or U1738 (N_1738,N_1187,N_1030);
nand U1739 (N_1739,N_1299,N_1199);
nor U1740 (N_1740,N_1441,N_1359);
nand U1741 (N_1741,N_1152,N_1476);
nand U1742 (N_1742,N_1038,N_1339);
nand U1743 (N_1743,N_1099,N_1121);
or U1744 (N_1744,N_1217,N_1146);
or U1745 (N_1745,N_1095,N_1343);
and U1746 (N_1746,N_1426,N_1183);
and U1747 (N_1747,N_1104,N_1314);
and U1748 (N_1748,N_1346,N_1052);
nand U1749 (N_1749,N_1005,N_1283);
nand U1750 (N_1750,N_1028,N_1275);
or U1751 (N_1751,N_1353,N_1180);
and U1752 (N_1752,N_1266,N_1340);
nand U1753 (N_1753,N_1072,N_1038);
nor U1754 (N_1754,N_1031,N_1047);
nand U1755 (N_1755,N_1284,N_1275);
and U1756 (N_1756,N_1480,N_1079);
and U1757 (N_1757,N_1348,N_1432);
nor U1758 (N_1758,N_1211,N_1198);
and U1759 (N_1759,N_1248,N_1496);
and U1760 (N_1760,N_1328,N_1389);
nand U1761 (N_1761,N_1015,N_1410);
or U1762 (N_1762,N_1469,N_1493);
or U1763 (N_1763,N_1057,N_1113);
and U1764 (N_1764,N_1465,N_1357);
and U1765 (N_1765,N_1140,N_1157);
nor U1766 (N_1766,N_1494,N_1037);
nor U1767 (N_1767,N_1328,N_1104);
nand U1768 (N_1768,N_1145,N_1263);
or U1769 (N_1769,N_1086,N_1397);
nor U1770 (N_1770,N_1354,N_1020);
nor U1771 (N_1771,N_1477,N_1086);
or U1772 (N_1772,N_1015,N_1487);
nor U1773 (N_1773,N_1027,N_1287);
nor U1774 (N_1774,N_1167,N_1082);
nand U1775 (N_1775,N_1455,N_1448);
nor U1776 (N_1776,N_1334,N_1441);
or U1777 (N_1777,N_1079,N_1277);
or U1778 (N_1778,N_1002,N_1064);
or U1779 (N_1779,N_1172,N_1046);
nor U1780 (N_1780,N_1498,N_1038);
and U1781 (N_1781,N_1100,N_1341);
nor U1782 (N_1782,N_1330,N_1118);
nor U1783 (N_1783,N_1337,N_1098);
nor U1784 (N_1784,N_1295,N_1101);
and U1785 (N_1785,N_1408,N_1293);
xnor U1786 (N_1786,N_1014,N_1007);
and U1787 (N_1787,N_1395,N_1094);
or U1788 (N_1788,N_1016,N_1298);
nor U1789 (N_1789,N_1048,N_1452);
or U1790 (N_1790,N_1308,N_1393);
nand U1791 (N_1791,N_1047,N_1341);
or U1792 (N_1792,N_1366,N_1298);
and U1793 (N_1793,N_1157,N_1458);
and U1794 (N_1794,N_1069,N_1356);
nand U1795 (N_1795,N_1085,N_1095);
or U1796 (N_1796,N_1289,N_1317);
or U1797 (N_1797,N_1444,N_1412);
nand U1798 (N_1798,N_1447,N_1481);
or U1799 (N_1799,N_1158,N_1450);
nor U1800 (N_1800,N_1340,N_1171);
or U1801 (N_1801,N_1284,N_1413);
nor U1802 (N_1802,N_1026,N_1203);
or U1803 (N_1803,N_1194,N_1188);
and U1804 (N_1804,N_1329,N_1095);
or U1805 (N_1805,N_1466,N_1447);
nand U1806 (N_1806,N_1280,N_1353);
nor U1807 (N_1807,N_1344,N_1009);
nor U1808 (N_1808,N_1287,N_1265);
or U1809 (N_1809,N_1135,N_1010);
or U1810 (N_1810,N_1126,N_1347);
nor U1811 (N_1811,N_1369,N_1242);
or U1812 (N_1812,N_1251,N_1063);
nand U1813 (N_1813,N_1097,N_1267);
or U1814 (N_1814,N_1191,N_1440);
nor U1815 (N_1815,N_1400,N_1472);
nand U1816 (N_1816,N_1271,N_1119);
and U1817 (N_1817,N_1091,N_1389);
nor U1818 (N_1818,N_1214,N_1156);
nor U1819 (N_1819,N_1451,N_1151);
or U1820 (N_1820,N_1061,N_1105);
nand U1821 (N_1821,N_1476,N_1209);
and U1822 (N_1822,N_1216,N_1318);
nand U1823 (N_1823,N_1220,N_1006);
xor U1824 (N_1824,N_1319,N_1255);
nand U1825 (N_1825,N_1234,N_1496);
or U1826 (N_1826,N_1492,N_1346);
and U1827 (N_1827,N_1463,N_1425);
nand U1828 (N_1828,N_1402,N_1033);
nor U1829 (N_1829,N_1401,N_1284);
nand U1830 (N_1830,N_1267,N_1303);
nand U1831 (N_1831,N_1365,N_1140);
and U1832 (N_1832,N_1299,N_1014);
or U1833 (N_1833,N_1238,N_1317);
nor U1834 (N_1834,N_1004,N_1468);
nand U1835 (N_1835,N_1416,N_1285);
nand U1836 (N_1836,N_1234,N_1173);
or U1837 (N_1837,N_1383,N_1229);
nor U1838 (N_1838,N_1080,N_1483);
xnor U1839 (N_1839,N_1481,N_1109);
or U1840 (N_1840,N_1375,N_1271);
or U1841 (N_1841,N_1188,N_1450);
nand U1842 (N_1842,N_1492,N_1491);
nor U1843 (N_1843,N_1155,N_1068);
and U1844 (N_1844,N_1311,N_1391);
and U1845 (N_1845,N_1000,N_1296);
nand U1846 (N_1846,N_1152,N_1230);
and U1847 (N_1847,N_1077,N_1185);
and U1848 (N_1848,N_1280,N_1135);
or U1849 (N_1849,N_1339,N_1428);
nand U1850 (N_1850,N_1128,N_1221);
nand U1851 (N_1851,N_1305,N_1088);
xor U1852 (N_1852,N_1174,N_1496);
xor U1853 (N_1853,N_1352,N_1309);
and U1854 (N_1854,N_1410,N_1180);
and U1855 (N_1855,N_1482,N_1355);
or U1856 (N_1856,N_1375,N_1341);
and U1857 (N_1857,N_1411,N_1124);
and U1858 (N_1858,N_1357,N_1381);
nor U1859 (N_1859,N_1339,N_1496);
and U1860 (N_1860,N_1226,N_1372);
and U1861 (N_1861,N_1046,N_1420);
or U1862 (N_1862,N_1271,N_1175);
nor U1863 (N_1863,N_1133,N_1327);
and U1864 (N_1864,N_1071,N_1205);
or U1865 (N_1865,N_1025,N_1041);
nor U1866 (N_1866,N_1189,N_1203);
or U1867 (N_1867,N_1437,N_1308);
nor U1868 (N_1868,N_1007,N_1082);
nor U1869 (N_1869,N_1107,N_1456);
or U1870 (N_1870,N_1161,N_1072);
and U1871 (N_1871,N_1497,N_1488);
and U1872 (N_1872,N_1091,N_1036);
nor U1873 (N_1873,N_1051,N_1036);
nor U1874 (N_1874,N_1298,N_1100);
and U1875 (N_1875,N_1202,N_1319);
nand U1876 (N_1876,N_1461,N_1271);
or U1877 (N_1877,N_1499,N_1186);
and U1878 (N_1878,N_1238,N_1131);
nand U1879 (N_1879,N_1065,N_1308);
or U1880 (N_1880,N_1242,N_1446);
and U1881 (N_1881,N_1058,N_1007);
or U1882 (N_1882,N_1152,N_1434);
nor U1883 (N_1883,N_1334,N_1072);
nand U1884 (N_1884,N_1253,N_1183);
nor U1885 (N_1885,N_1001,N_1357);
xnor U1886 (N_1886,N_1229,N_1334);
nor U1887 (N_1887,N_1185,N_1153);
nor U1888 (N_1888,N_1335,N_1342);
or U1889 (N_1889,N_1086,N_1249);
nor U1890 (N_1890,N_1388,N_1409);
nor U1891 (N_1891,N_1122,N_1078);
nand U1892 (N_1892,N_1177,N_1071);
or U1893 (N_1893,N_1073,N_1110);
and U1894 (N_1894,N_1497,N_1034);
and U1895 (N_1895,N_1448,N_1492);
or U1896 (N_1896,N_1488,N_1126);
and U1897 (N_1897,N_1468,N_1034);
nor U1898 (N_1898,N_1299,N_1275);
and U1899 (N_1899,N_1494,N_1484);
nor U1900 (N_1900,N_1434,N_1279);
or U1901 (N_1901,N_1338,N_1166);
nand U1902 (N_1902,N_1228,N_1255);
or U1903 (N_1903,N_1307,N_1105);
nand U1904 (N_1904,N_1021,N_1121);
and U1905 (N_1905,N_1268,N_1328);
nor U1906 (N_1906,N_1441,N_1254);
nand U1907 (N_1907,N_1469,N_1352);
nand U1908 (N_1908,N_1267,N_1405);
or U1909 (N_1909,N_1407,N_1058);
nor U1910 (N_1910,N_1049,N_1034);
or U1911 (N_1911,N_1360,N_1279);
xnor U1912 (N_1912,N_1181,N_1179);
or U1913 (N_1913,N_1309,N_1265);
nand U1914 (N_1914,N_1384,N_1015);
or U1915 (N_1915,N_1230,N_1180);
nand U1916 (N_1916,N_1210,N_1107);
nand U1917 (N_1917,N_1053,N_1131);
nand U1918 (N_1918,N_1264,N_1468);
and U1919 (N_1919,N_1452,N_1273);
and U1920 (N_1920,N_1038,N_1329);
or U1921 (N_1921,N_1476,N_1327);
nor U1922 (N_1922,N_1275,N_1251);
xnor U1923 (N_1923,N_1248,N_1401);
nor U1924 (N_1924,N_1387,N_1264);
nand U1925 (N_1925,N_1067,N_1257);
and U1926 (N_1926,N_1137,N_1324);
or U1927 (N_1927,N_1167,N_1091);
and U1928 (N_1928,N_1145,N_1370);
and U1929 (N_1929,N_1304,N_1492);
nand U1930 (N_1930,N_1013,N_1486);
nor U1931 (N_1931,N_1124,N_1171);
nor U1932 (N_1932,N_1374,N_1132);
nor U1933 (N_1933,N_1146,N_1134);
and U1934 (N_1934,N_1192,N_1080);
nand U1935 (N_1935,N_1090,N_1276);
and U1936 (N_1936,N_1268,N_1074);
or U1937 (N_1937,N_1171,N_1364);
nor U1938 (N_1938,N_1268,N_1184);
xor U1939 (N_1939,N_1120,N_1110);
nand U1940 (N_1940,N_1222,N_1111);
nand U1941 (N_1941,N_1256,N_1013);
and U1942 (N_1942,N_1387,N_1123);
or U1943 (N_1943,N_1399,N_1274);
and U1944 (N_1944,N_1494,N_1188);
and U1945 (N_1945,N_1394,N_1221);
and U1946 (N_1946,N_1088,N_1258);
or U1947 (N_1947,N_1498,N_1371);
nor U1948 (N_1948,N_1038,N_1416);
nand U1949 (N_1949,N_1199,N_1112);
nor U1950 (N_1950,N_1264,N_1046);
nand U1951 (N_1951,N_1257,N_1121);
nor U1952 (N_1952,N_1047,N_1157);
nor U1953 (N_1953,N_1300,N_1268);
nand U1954 (N_1954,N_1439,N_1449);
nor U1955 (N_1955,N_1201,N_1137);
and U1956 (N_1956,N_1004,N_1358);
or U1957 (N_1957,N_1109,N_1341);
and U1958 (N_1958,N_1374,N_1489);
nand U1959 (N_1959,N_1123,N_1040);
nand U1960 (N_1960,N_1145,N_1219);
and U1961 (N_1961,N_1078,N_1351);
nand U1962 (N_1962,N_1395,N_1467);
nor U1963 (N_1963,N_1346,N_1015);
and U1964 (N_1964,N_1478,N_1204);
xnor U1965 (N_1965,N_1015,N_1351);
nand U1966 (N_1966,N_1400,N_1247);
and U1967 (N_1967,N_1138,N_1063);
or U1968 (N_1968,N_1463,N_1246);
nor U1969 (N_1969,N_1115,N_1319);
or U1970 (N_1970,N_1069,N_1346);
and U1971 (N_1971,N_1050,N_1084);
or U1972 (N_1972,N_1433,N_1350);
and U1973 (N_1973,N_1313,N_1030);
or U1974 (N_1974,N_1334,N_1128);
nor U1975 (N_1975,N_1218,N_1240);
nand U1976 (N_1976,N_1360,N_1061);
nor U1977 (N_1977,N_1274,N_1189);
nor U1978 (N_1978,N_1412,N_1004);
and U1979 (N_1979,N_1039,N_1142);
nor U1980 (N_1980,N_1221,N_1433);
nand U1981 (N_1981,N_1438,N_1303);
or U1982 (N_1982,N_1425,N_1136);
or U1983 (N_1983,N_1260,N_1080);
xnor U1984 (N_1984,N_1266,N_1382);
or U1985 (N_1985,N_1041,N_1466);
or U1986 (N_1986,N_1116,N_1415);
xnor U1987 (N_1987,N_1013,N_1119);
xor U1988 (N_1988,N_1481,N_1312);
nand U1989 (N_1989,N_1068,N_1081);
nor U1990 (N_1990,N_1290,N_1192);
nand U1991 (N_1991,N_1231,N_1135);
nand U1992 (N_1992,N_1384,N_1239);
or U1993 (N_1993,N_1473,N_1145);
and U1994 (N_1994,N_1374,N_1249);
nor U1995 (N_1995,N_1061,N_1123);
or U1996 (N_1996,N_1039,N_1181);
and U1997 (N_1997,N_1064,N_1496);
or U1998 (N_1998,N_1102,N_1421);
or U1999 (N_1999,N_1415,N_1407);
nand U2000 (N_2000,N_1707,N_1561);
nand U2001 (N_2001,N_1997,N_1821);
and U2002 (N_2002,N_1625,N_1600);
or U2003 (N_2003,N_1884,N_1987);
nor U2004 (N_2004,N_1623,N_1601);
or U2005 (N_2005,N_1603,N_1781);
nand U2006 (N_2006,N_1942,N_1655);
and U2007 (N_2007,N_1618,N_1830);
or U2008 (N_2008,N_1742,N_1629);
or U2009 (N_2009,N_1509,N_1699);
nand U2010 (N_2010,N_1851,N_1980);
or U2011 (N_2011,N_1711,N_1572);
and U2012 (N_2012,N_1864,N_1900);
nor U2013 (N_2013,N_1822,N_1801);
or U2014 (N_2014,N_1974,N_1986);
nor U2015 (N_2015,N_1857,N_1598);
nand U2016 (N_2016,N_1798,N_1510);
nand U2017 (N_2017,N_1962,N_1688);
or U2018 (N_2018,N_1813,N_1779);
xnor U2019 (N_2019,N_1535,N_1511);
nand U2020 (N_2020,N_1671,N_1916);
nand U2021 (N_2021,N_1966,N_1639);
nand U2022 (N_2022,N_1907,N_1663);
nand U2023 (N_2023,N_1861,N_1836);
or U2024 (N_2024,N_1754,N_1691);
and U2025 (N_2025,N_1724,N_1532);
or U2026 (N_2026,N_1853,N_1810);
nor U2027 (N_2027,N_1709,N_1784);
nor U2028 (N_2028,N_1874,N_1825);
and U2029 (N_2029,N_1653,N_1721);
nor U2030 (N_2030,N_1506,N_1552);
or U2031 (N_2031,N_1934,N_1744);
or U2032 (N_2032,N_1938,N_1776);
nand U2033 (N_2033,N_1602,N_1689);
xor U2034 (N_2034,N_1797,N_1880);
nand U2035 (N_2035,N_1673,N_1740);
or U2036 (N_2036,N_1722,N_1675);
or U2037 (N_2037,N_1659,N_1568);
and U2038 (N_2038,N_1581,N_1931);
nand U2039 (N_2039,N_1878,N_1679);
or U2040 (N_2040,N_1895,N_1984);
nor U2041 (N_2041,N_1956,N_1988);
and U2042 (N_2042,N_1854,N_1534);
and U2043 (N_2043,N_1838,N_1971);
or U2044 (N_2044,N_1745,N_1786);
nand U2045 (N_2045,N_1865,N_1860);
and U2046 (N_2046,N_1644,N_1614);
nor U2047 (N_2047,N_1573,N_1904);
nand U2048 (N_2048,N_1730,N_1547);
nand U2049 (N_2049,N_1785,N_1719);
nor U2050 (N_2050,N_1993,N_1763);
nor U2051 (N_2051,N_1915,N_1991);
and U2052 (N_2052,N_1893,N_1804);
or U2053 (N_2053,N_1589,N_1564);
nor U2054 (N_2054,N_1762,N_1608);
nand U2055 (N_2055,N_1769,N_1992);
and U2056 (N_2056,N_1520,N_1536);
or U2057 (N_2057,N_1518,N_1823);
or U2058 (N_2058,N_1908,N_1641);
nor U2059 (N_2059,N_1866,N_1901);
or U2060 (N_2060,N_1698,N_1947);
nor U2061 (N_2061,N_1648,N_1695);
and U2062 (N_2062,N_1682,N_1761);
nand U2063 (N_2063,N_1670,N_1972);
and U2064 (N_2064,N_1898,N_1835);
and U2065 (N_2065,N_1543,N_1728);
or U2066 (N_2066,N_1579,N_1959);
nor U2067 (N_2067,N_1549,N_1846);
or U2068 (N_2068,N_1867,N_1584);
or U2069 (N_2069,N_1945,N_1593);
nand U2070 (N_2070,N_1727,N_1583);
nand U2071 (N_2071,N_1604,N_1850);
or U2072 (N_2072,N_1713,N_1967);
and U2073 (N_2073,N_1569,N_1859);
or U2074 (N_2074,N_1516,N_1737);
and U2075 (N_2075,N_1676,N_1734);
or U2076 (N_2076,N_1687,N_1530);
and U2077 (N_2077,N_1531,N_1729);
nand U2078 (N_2078,N_1862,N_1886);
nor U2079 (N_2079,N_1523,N_1831);
and U2080 (N_2080,N_1818,N_1940);
and U2081 (N_2081,N_1505,N_1750);
or U2082 (N_2082,N_1844,N_1599);
or U2083 (N_2083,N_1672,N_1944);
nor U2084 (N_2084,N_1774,N_1811);
and U2085 (N_2085,N_1977,N_1789);
nand U2086 (N_2086,N_1758,N_1826);
or U2087 (N_2087,N_1650,N_1999);
nor U2088 (N_2088,N_1560,N_1732);
or U2089 (N_2089,N_1925,N_1527);
nand U2090 (N_2090,N_1649,N_1773);
or U2091 (N_2091,N_1747,N_1712);
nand U2092 (N_2092,N_1611,N_1808);
nor U2093 (N_2093,N_1665,N_1620);
or U2094 (N_2094,N_1897,N_1749);
or U2095 (N_2095,N_1819,N_1802);
nand U2096 (N_2096,N_1871,N_1660);
or U2097 (N_2097,N_1680,N_1705);
nand U2098 (N_2098,N_1922,N_1906);
nand U2099 (N_2099,N_1877,N_1664);
nor U2100 (N_2100,N_1591,N_1949);
and U2101 (N_2101,N_1782,N_1697);
and U2102 (N_2102,N_1950,N_1545);
or U2103 (N_2103,N_1894,N_1519);
or U2104 (N_2104,N_1610,N_1587);
nand U2105 (N_2105,N_1780,N_1958);
and U2106 (N_2106,N_1500,N_1556);
and U2107 (N_2107,N_1626,N_1981);
nand U2108 (N_2108,N_1704,N_1631);
nor U2109 (N_2109,N_1766,N_1787);
or U2110 (N_2110,N_1803,N_1996);
nand U2111 (N_2111,N_1507,N_1985);
and U2112 (N_2112,N_1582,N_1903);
nand U2113 (N_2113,N_1829,N_1933);
nor U2114 (N_2114,N_1968,N_1989);
and U2115 (N_2115,N_1768,N_1508);
nor U2116 (N_2116,N_1863,N_1788);
nor U2117 (N_2117,N_1794,N_1647);
nand U2118 (N_2118,N_1674,N_1632);
nand U2119 (N_2119,N_1553,N_1638);
nor U2120 (N_2120,N_1615,N_1735);
or U2121 (N_2121,N_1733,N_1783);
xnor U2122 (N_2122,N_1834,N_1590);
nor U2123 (N_2123,N_1953,N_1725);
nor U2124 (N_2124,N_1684,N_1678);
nor U2125 (N_2125,N_1890,N_1912);
nor U2126 (N_2126,N_1995,N_1909);
and U2127 (N_2127,N_1990,N_1771);
and U2128 (N_2128,N_1640,N_1832);
nand U2129 (N_2129,N_1605,N_1833);
nand U2130 (N_2130,N_1855,N_1517);
nor U2131 (N_2131,N_1720,N_1979);
nand U2132 (N_2132,N_1645,N_1924);
nand U2133 (N_2133,N_1970,N_1827);
nor U2134 (N_2134,N_1752,N_1816);
nor U2135 (N_2135,N_1919,N_1790);
or U2136 (N_2136,N_1914,N_1976);
nand U2137 (N_2137,N_1946,N_1576);
and U2138 (N_2138,N_1723,N_1791);
or U2139 (N_2139,N_1716,N_1566);
or U2140 (N_2140,N_1800,N_1551);
nor U2141 (N_2141,N_1570,N_1805);
nand U2142 (N_2142,N_1760,N_1926);
or U2143 (N_2143,N_1841,N_1902);
nor U2144 (N_2144,N_1957,N_1753);
nor U2145 (N_2145,N_1539,N_1501);
and U2146 (N_2146,N_1875,N_1913);
and U2147 (N_2147,N_1872,N_1693);
or U2148 (N_2148,N_1613,N_1726);
and U2149 (N_2149,N_1537,N_1708);
and U2150 (N_2150,N_1792,N_1627);
nor U2151 (N_2151,N_1636,N_1522);
xor U2152 (N_2152,N_1883,N_1619);
nor U2153 (N_2153,N_1548,N_1559);
nand U2154 (N_2154,N_1755,N_1888);
nor U2155 (N_2155,N_1954,N_1935);
nor U2156 (N_2156,N_1738,N_1929);
or U2157 (N_2157,N_1637,N_1597);
nand U2158 (N_2158,N_1557,N_1594);
nor U2159 (N_2159,N_1960,N_1911);
nand U2160 (N_2160,N_1892,N_1681);
and U2161 (N_2161,N_1550,N_1964);
nand U2162 (N_2162,N_1828,N_1651);
and U2163 (N_2163,N_1936,N_1899);
or U2164 (N_2164,N_1703,N_1658);
nor U2165 (N_2165,N_1567,N_1630);
xor U2166 (N_2166,N_1905,N_1796);
and U2167 (N_2167,N_1809,N_1624);
nand U2168 (N_2168,N_1994,N_1503);
or U2169 (N_2169,N_1667,N_1715);
or U2170 (N_2170,N_1927,N_1939);
nor U2171 (N_2171,N_1952,N_1617);
nand U2172 (N_2172,N_1702,N_1876);
xor U2173 (N_2173,N_1662,N_1778);
nor U2174 (N_2174,N_1812,N_1669);
or U2175 (N_2175,N_1546,N_1526);
nand U2176 (N_2176,N_1982,N_1643);
or U2177 (N_2177,N_1542,N_1858);
nand U2178 (N_2178,N_1686,N_1628);
or U2179 (N_2179,N_1683,N_1574);
nor U2180 (N_2180,N_1706,N_1575);
nand U2181 (N_2181,N_1748,N_1529);
nor U2182 (N_2182,N_1504,N_1588);
nor U2183 (N_2183,N_1856,N_1592);
or U2184 (N_2184,N_1634,N_1983);
nor U2185 (N_2185,N_1917,N_1918);
or U2186 (N_2186,N_1596,N_1652);
nand U2187 (N_2187,N_1973,N_1746);
nand U2188 (N_2188,N_1932,N_1795);
nand U2189 (N_2189,N_1852,N_1558);
nor U2190 (N_2190,N_1538,N_1881);
nor U2191 (N_2191,N_1873,N_1694);
nor U2192 (N_2192,N_1837,N_1941);
nor U2193 (N_2193,N_1879,N_1642);
or U2194 (N_2194,N_1621,N_1661);
and U2195 (N_2195,N_1514,N_1889);
or U2196 (N_2196,N_1580,N_1765);
or U2197 (N_2197,N_1690,N_1585);
xnor U2198 (N_2198,N_1717,N_1612);
xnor U2199 (N_2199,N_1814,N_1622);
or U2200 (N_2200,N_1743,N_1777);
nand U2201 (N_2201,N_1891,N_1616);
nor U2202 (N_2202,N_1843,N_1839);
or U2203 (N_2203,N_1607,N_1930);
xor U2204 (N_2204,N_1820,N_1562);
and U2205 (N_2205,N_1513,N_1824);
nand U2206 (N_2206,N_1512,N_1606);
and U2207 (N_2207,N_1767,N_1975);
nand U2208 (N_2208,N_1710,N_1882);
or U2209 (N_2209,N_1969,N_1541);
or U2210 (N_2210,N_1544,N_1961);
and U2211 (N_2211,N_1928,N_1978);
nor U2212 (N_2212,N_1577,N_1515);
nor U2213 (N_2213,N_1571,N_1700);
and U2214 (N_2214,N_1955,N_1696);
nand U2215 (N_2215,N_1840,N_1646);
and U2216 (N_2216,N_1920,N_1937);
or U2217 (N_2217,N_1668,N_1868);
nand U2218 (N_2218,N_1799,N_1502);
and U2219 (N_2219,N_1759,N_1870);
nor U2220 (N_2220,N_1718,N_1817);
or U2221 (N_2221,N_1815,N_1714);
and U2222 (N_2222,N_1923,N_1739);
and U2223 (N_2223,N_1951,N_1578);
nor U2224 (N_2224,N_1666,N_1887);
nand U2225 (N_2225,N_1586,N_1731);
or U2226 (N_2226,N_1595,N_1775);
nand U2227 (N_2227,N_1965,N_1524);
nor U2228 (N_2228,N_1896,N_1842);
or U2229 (N_2229,N_1756,N_1793);
xor U2230 (N_2230,N_1869,N_1998);
or U2231 (N_2231,N_1751,N_1807);
nor U2232 (N_2232,N_1741,N_1885);
nor U2233 (N_2233,N_1757,N_1847);
nand U2234 (N_2234,N_1635,N_1770);
nand U2235 (N_2235,N_1701,N_1533);
nand U2236 (N_2236,N_1736,N_1806);
and U2237 (N_2237,N_1921,N_1657);
nor U2238 (N_2238,N_1963,N_1565);
nor U2239 (N_2239,N_1656,N_1609);
or U2240 (N_2240,N_1910,N_1540);
and U2241 (N_2241,N_1555,N_1685);
or U2242 (N_2242,N_1948,N_1848);
or U2243 (N_2243,N_1525,N_1772);
nand U2244 (N_2244,N_1845,N_1849);
and U2245 (N_2245,N_1554,N_1692);
or U2246 (N_2246,N_1521,N_1528);
and U2247 (N_2247,N_1633,N_1677);
nor U2248 (N_2248,N_1563,N_1764);
or U2249 (N_2249,N_1943,N_1654);
or U2250 (N_2250,N_1823,N_1801);
and U2251 (N_2251,N_1901,N_1769);
or U2252 (N_2252,N_1898,N_1770);
nand U2253 (N_2253,N_1656,N_1607);
xor U2254 (N_2254,N_1584,N_1808);
nor U2255 (N_2255,N_1790,N_1544);
and U2256 (N_2256,N_1545,N_1526);
nor U2257 (N_2257,N_1910,N_1827);
or U2258 (N_2258,N_1821,N_1893);
nor U2259 (N_2259,N_1867,N_1750);
xnor U2260 (N_2260,N_1956,N_1648);
nand U2261 (N_2261,N_1952,N_1633);
and U2262 (N_2262,N_1965,N_1904);
nor U2263 (N_2263,N_1523,N_1570);
or U2264 (N_2264,N_1808,N_1975);
nor U2265 (N_2265,N_1525,N_1622);
nand U2266 (N_2266,N_1720,N_1970);
and U2267 (N_2267,N_1948,N_1899);
nor U2268 (N_2268,N_1680,N_1682);
or U2269 (N_2269,N_1511,N_1905);
or U2270 (N_2270,N_1836,N_1803);
or U2271 (N_2271,N_1982,N_1852);
nand U2272 (N_2272,N_1792,N_1973);
nor U2273 (N_2273,N_1658,N_1943);
and U2274 (N_2274,N_1505,N_1855);
nand U2275 (N_2275,N_1678,N_1899);
nor U2276 (N_2276,N_1883,N_1956);
nor U2277 (N_2277,N_1871,N_1663);
nor U2278 (N_2278,N_1928,N_1899);
nor U2279 (N_2279,N_1642,N_1711);
and U2280 (N_2280,N_1806,N_1899);
nand U2281 (N_2281,N_1621,N_1574);
nand U2282 (N_2282,N_1851,N_1979);
nand U2283 (N_2283,N_1613,N_1780);
and U2284 (N_2284,N_1718,N_1634);
and U2285 (N_2285,N_1561,N_1858);
and U2286 (N_2286,N_1848,N_1771);
nor U2287 (N_2287,N_1937,N_1934);
nor U2288 (N_2288,N_1922,N_1554);
or U2289 (N_2289,N_1890,N_1571);
nor U2290 (N_2290,N_1986,N_1669);
and U2291 (N_2291,N_1861,N_1966);
or U2292 (N_2292,N_1734,N_1950);
and U2293 (N_2293,N_1505,N_1721);
xnor U2294 (N_2294,N_1772,N_1696);
or U2295 (N_2295,N_1855,N_1867);
and U2296 (N_2296,N_1705,N_1834);
nor U2297 (N_2297,N_1805,N_1591);
nor U2298 (N_2298,N_1933,N_1849);
or U2299 (N_2299,N_1663,N_1595);
nand U2300 (N_2300,N_1852,N_1962);
or U2301 (N_2301,N_1807,N_1542);
nor U2302 (N_2302,N_1930,N_1981);
or U2303 (N_2303,N_1701,N_1882);
or U2304 (N_2304,N_1722,N_1636);
nor U2305 (N_2305,N_1669,N_1910);
or U2306 (N_2306,N_1737,N_1758);
and U2307 (N_2307,N_1981,N_1933);
nor U2308 (N_2308,N_1522,N_1594);
or U2309 (N_2309,N_1684,N_1616);
nor U2310 (N_2310,N_1735,N_1850);
or U2311 (N_2311,N_1758,N_1676);
and U2312 (N_2312,N_1541,N_1899);
nor U2313 (N_2313,N_1825,N_1882);
and U2314 (N_2314,N_1907,N_1906);
nor U2315 (N_2315,N_1863,N_1599);
or U2316 (N_2316,N_1625,N_1794);
and U2317 (N_2317,N_1778,N_1963);
or U2318 (N_2318,N_1626,N_1767);
or U2319 (N_2319,N_1930,N_1950);
and U2320 (N_2320,N_1515,N_1684);
nand U2321 (N_2321,N_1514,N_1899);
or U2322 (N_2322,N_1708,N_1935);
and U2323 (N_2323,N_1941,N_1572);
nor U2324 (N_2324,N_1707,N_1786);
or U2325 (N_2325,N_1928,N_1669);
or U2326 (N_2326,N_1590,N_1514);
or U2327 (N_2327,N_1559,N_1919);
nor U2328 (N_2328,N_1540,N_1763);
nor U2329 (N_2329,N_1850,N_1946);
nor U2330 (N_2330,N_1826,N_1594);
and U2331 (N_2331,N_1615,N_1743);
nand U2332 (N_2332,N_1716,N_1970);
and U2333 (N_2333,N_1783,N_1738);
and U2334 (N_2334,N_1700,N_1691);
and U2335 (N_2335,N_1843,N_1832);
and U2336 (N_2336,N_1984,N_1997);
and U2337 (N_2337,N_1905,N_1862);
and U2338 (N_2338,N_1841,N_1730);
and U2339 (N_2339,N_1615,N_1722);
nand U2340 (N_2340,N_1636,N_1823);
nor U2341 (N_2341,N_1859,N_1698);
and U2342 (N_2342,N_1549,N_1916);
or U2343 (N_2343,N_1528,N_1783);
or U2344 (N_2344,N_1561,N_1672);
and U2345 (N_2345,N_1707,N_1770);
nor U2346 (N_2346,N_1575,N_1692);
nand U2347 (N_2347,N_1991,N_1827);
or U2348 (N_2348,N_1640,N_1944);
nor U2349 (N_2349,N_1646,N_1531);
xnor U2350 (N_2350,N_1789,N_1808);
nor U2351 (N_2351,N_1974,N_1752);
nor U2352 (N_2352,N_1963,N_1683);
nand U2353 (N_2353,N_1657,N_1932);
nor U2354 (N_2354,N_1716,N_1759);
nand U2355 (N_2355,N_1540,N_1890);
and U2356 (N_2356,N_1684,N_1634);
nor U2357 (N_2357,N_1905,N_1704);
and U2358 (N_2358,N_1635,N_1643);
nand U2359 (N_2359,N_1672,N_1965);
or U2360 (N_2360,N_1608,N_1703);
nor U2361 (N_2361,N_1650,N_1914);
and U2362 (N_2362,N_1642,N_1772);
nand U2363 (N_2363,N_1691,N_1939);
and U2364 (N_2364,N_1930,N_1629);
or U2365 (N_2365,N_1960,N_1924);
or U2366 (N_2366,N_1693,N_1662);
nand U2367 (N_2367,N_1776,N_1802);
and U2368 (N_2368,N_1690,N_1807);
nor U2369 (N_2369,N_1971,N_1832);
or U2370 (N_2370,N_1861,N_1598);
nor U2371 (N_2371,N_1885,N_1860);
and U2372 (N_2372,N_1505,N_1723);
and U2373 (N_2373,N_1896,N_1651);
nand U2374 (N_2374,N_1742,N_1739);
nor U2375 (N_2375,N_1899,N_1556);
nand U2376 (N_2376,N_1834,N_1916);
nor U2377 (N_2377,N_1973,N_1955);
or U2378 (N_2378,N_1893,N_1708);
nor U2379 (N_2379,N_1970,N_1921);
and U2380 (N_2380,N_1711,N_1835);
nor U2381 (N_2381,N_1696,N_1767);
nand U2382 (N_2382,N_1561,N_1598);
xor U2383 (N_2383,N_1924,N_1811);
nand U2384 (N_2384,N_1692,N_1585);
and U2385 (N_2385,N_1890,N_1739);
xnor U2386 (N_2386,N_1765,N_1813);
nand U2387 (N_2387,N_1761,N_1966);
nand U2388 (N_2388,N_1728,N_1811);
nor U2389 (N_2389,N_1839,N_1636);
nand U2390 (N_2390,N_1547,N_1728);
and U2391 (N_2391,N_1776,N_1892);
xnor U2392 (N_2392,N_1841,N_1927);
nand U2393 (N_2393,N_1817,N_1696);
and U2394 (N_2394,N_1808,N_1616);
nor U2395 (N_2395,N_1992,N_1965);
or U2396 (N_2396,N_1922,N_1680);
and U2397 (N_2397,N_1872,N_1905);
and U2398 (N_2398,N_1751,N_1937);
and U2399 (N_2399,N_1692,N_1807);
and U2400 (N_2400,N_1656,N_1677);
or U2401 (N_2401,N_1619,N_1938);
nand U2402 (N_2402,N_1878,N_1755);
nand U2403 (N_2403,N_1623,N_1816);
and U2404 (N_2404,N_1700,N_1719);
and U2405 (N_2405,N_1982,N_1682);
nor U2406 (N_2406,N_1612,N_1833);
and U2407 (N_2407,N_1771,N_1805);
nand U2408 (N_2408,N_1995,N_1942);
or U2409 (N_2409,N_1656,N_1529);
nor U2410 (N_2410,N_1760,N_1919);
nor U2411 (N_2411,N_1883,N_1547);
nor U2412 (N_2412,N_1709,N_1515);
or U2413 (N_2413,N_1711,N_1734);
nand U2414 (N_2414,N_1778,N_1762);
and U2415 (N_2415,N_1864,N_1603);
or U2416 (N_2416,N_1513,N_1569);
nor U2417 (N_2417,N_1826,N_1602);
and U2418 (N_2418,N_1992,N_1856);
and U2419 (N_2419,N_1746,N_1803);
nand U2420 (N_2420,N_1674,N_1550);
nor U2421 (N_2421,N_1567,N_1585);
nand U2422 (N_2422,N_1951,N_1759);
nor U2423 (N_2423,N_1890,N_1913);
nand U2424 (N_2424,N_1949,N_1820);
nor U2425 (N_2425,N_1549,N_1709);
or U2426 (N_2426,N_1531,N_1556);
nand U2427 (N_2427,N_1824,N_1784);
or U2428 (N_2428,N_1583,N_1673);
xor U2429 (N_2429,N_1696,N_1916);
nor U2430 (N_2430,N_1902,N_1927);
xnor U2431 (N_2431,N_1889,N_1620);
nor U2432 (N_2432,N_1968,N_1727);
nand U2433 (N_2433,N_1589,N_1903);
nor U2434 (N_2434,N_1899,N_1673);
nand U2435 (N_2435,N_1525,N_1593);
or U2436 (N_2436,N_1684,N_1901);
nand U2437 (N_2437,N_1749,N_1951);
xnor U2438 (N_2438,N_1643,N_1784);
xor U2439 (N_2439,N_1590,N_1958);
nor U2440 (N_2440,N_1719,N_1706);
nand U2441 (N_2441,N_1673,N_1772);
or U2442 (N_2442,N_1724,N_1940);
nor U2443 (N_2443,N_1740,N_1674);
or U2444 (N_2444,N_1597,N_1661);
xor U2445 (N_2445,N_1895,N_1790);
or U2446 (N_2446,N_1705,N_1544);
nor U2447 (N_2447,N_1665,N_1942);
nor U2448 (N_2448,N_1917,N_1642);
and U2449 (N_2449,N_1739,N_1882);
or U2450 (N_2450,N_1833,N_1554);
and U2451 (N_2451,N_1556,N_1694);
nand U2452 (N_2452,N_1559,N_1909);
and U2453 (N_2453,N_1522,N_1754);
and U2454 (N_2454,N_1831,N_1599);
nand U2455 (N_2455,N_1576,N_1977);
nand U2456 (N_2456,N_1766,N_1685);
or U2457 (N_2457,N_1540,N_1804);
and U2458 (N_2458,N_1584,N_1991);
and U2459 (N_2459,N_1544,N_1519);
nand U2460 (N_2460,N_1700,N_1635);
and U2461 (N_2461,N_1658,N_1898);
nor U2462 (N_2462,N_1992,N_1980);
nand U2463 (N_2463,N_1516,N_1813);
or U2464 (N_2464,N_1776,N_1923);
and U2465 (N_2465,N_1765,N_1836);
nand U2466 (N_2466,N_1532,N_1742);
nor U2467 (N_2467,N_1799,N_1859);
nand U2468 (N_2468,N_1656,N_1824);
or U2469 (N_2469,N_1560,N_1792);
nand U2470 (N_2470,N_1978,N_1773);
nand U2471 (N_2471,N_1661,N_1773);
and U2472 (N_2472,N_1638,N_1585);
nand U2473 (N_2473,N_1849,N_1561);
and U2474 (N_2474,N_1969,N_1926);
and U2475 (N_2475,N_1636,N_1602);
or U2476 (N_2476,N_1714,N_1742);
and U2477 (N_2477,N_1860,N_1892);
nand U2478 (N_2478,N_1924,N_1773);
nor U2479 (N_2479,N_1750,N_1890);
nand U2480 (N_2480,N_1709,N_1579);
or U2481 (N_2481,N_1574,N_1560);
or U2482 (N_2482,N_1693,N_1878);
or U2483 (N_2483,N_1697,N_1706);
and U2484 (N_2484,N_1850,N_1780);
nor U2485 (N_2485,N_1677,N_1702);
nor U2486 (N_2486,N_1884,N_1934);
nand U2487 (N_2487,N_1563,N_1592);
nand U2488 (N_2488,N_1814,N_1679);
nor U2489 (N_2489,N_1720,N_1955);
nand U2490 (N_2490,N_1976,N_1936);
nand U2491 (N_2491,N_1682,N_1570);
xor U2492 (N_2492,N_1991,N_1592);
and U2493 (N_2493,N_1686,N_1837);
nor U2494 (N_2494,N_1653,N_1553);
or U2495 (N_2495,N_1962,N_1855);
or U2496 (N_2496,N_1778,N_1980);
or U2497 (N_2497,N_1986,N_1976);
nand U2498 (N_2498,N_1844,N_1509);
nor U2499 (N_2499,N_1689,N_1744);
nor U2500 (N_2500,N_2492,N_2163);
nor U2501 (N_2501,N_2319,N_2318);
and U2502 (N_2502,N_2149,N_2044);
and U2503 (N_2503,N_2379,N_2038);
nand U2504 (N_2504,N_2205,N_2181);
nor U2505 (N_2505,N_2306,N_2226);
nand U2506 (N_2506,N_2258,N_2328);
nand U2507 (N_2507,N_2015,N_2183);
nand U2508 (N_2508,N_2124,N_2081);
nand U2509 (N_2509,N_2065,N_2176);
nor U2510 (N_2510,N_2166,N_2434);
nor U2511 (N_2511,N_2324,N_2240);
nor U2512 (N_2512,N_2252,N_2236);
or U2513 (N_2513,N_2125,N_2112);
nor U2514 (N_2514,N_2043,N_2141);
and U2515 (N_2515,N_2344,N_2000);
nor U2516 (N_2516,N_2440,N_2169);
nor U2517 (N_2517,N_2211,N_2210);
or U2518 (N_2518,N_2018,N_2131);
or U2519 (N_2519,N_2419,N_2208);
and U2520 (N_2520,N_2099,N_2050);
or U2521 (N_2521,N_2161,N_2375);
nand U2522 (N_2522,N_2489,N_2037);
and U2523 (N_2523,N_2334,N_2468);
nand U2524 (N_2524,N_2005,N_2311);
nand U2525 (N_2525,N_2416,N_2317);
nand U2526 (N_2526,N_2310,N_2373);
and U2527 (N_2527,N_2076,N_2261);
or U2528 (N_2528,N_2403,N_2188);
nand U2529 (N_2529,N_2206,N_2360);
and U2530 (N_2530,N_2077,N_2260);
nand U2531 (N_2531,N_2048,N_2248);
nand U2532 (N_2532,N_2243,N_2481);
nor U2533 (N_2533,N_2085,N_2233);
nand U2534 (N_2534,N_2136,N_2106);
nor U2535 (N_2535,N_2402,N_2122);
nand U2536 (N_2536,N_2443,N_2144);
and U2537 (N_2537,N_2337,N_2105);
nand U2538 (N_2538,N_2285,N_2126);
nor U2539 (N_2539,N_2145,N_2057);
or U2540 (N_2540,N_2182,N_2263);
nor U2541 (N_2541,N_2372,N_2142);
or U2542 (N_2542,N_2284,N_2457);
nand U2543 (N_2543,N_2363,N_2305);
nor U2544 (N_2544,N_2436,N_2409);
nor U2545 (N_2545,N_2472,N_2341);
and U2546 (N_2546,N_2414,N_2231);
or U2547 (N_2547,N_2281,N_2437);
or U2548 (N_2548,N_2115,N_2449);
or U2549 (N_2549,N_2474,N_2079);
and U2550 (N_2550,N_2304,N_2390);
or U2551 (N_2551,N_2499,N_2199);
and U2552 (N_2552,N_2446,N_2488);
nor U2553 (N_2553,N_2367,N_2086);
and U2554 (N_2554,N_2060,N_2279);
nor U2555 (N_2555,N_2430,N_2030);
nor U2556 (N_2556,N_2498,N_2275);
or U2557 (N_2557,N_2072,N_2022);
xnor U2558 (N_2558,N_2271,N_2359);
or U2559 (N_2559,N_2246,N_2389);
nand U2560 (N_2560,N_2251,N_2380);
nand U2561 (N_2561,N_2160,N_2046);
nand U2562 (N_2562,N_2027,N_2358);
nor U2563 (N_2563,N_2450,N_2392);
and U2564 (N_2564,N_2068,N_2399);
and U2565 (N_2565,N_2137,N_2454);
nor U2566 (N_2566,N_2249,N_2150);
or U2567 (N_2567,N_2152,N_2484);
or U2568 (N_2568,N_2354,N_2276);
or U2569 (N_2569,N_2335,N_2026);
and U2570 (N_2570,N_2098,N_2415);
and U2571 (N_2571,N_2384,N_2366);
nand U2572 (N_2572,N_2218,N_2111);
or U2573 (N_2573,N_2227,N_2331);
or U2574 (N_2574,N_2041,N_2445);
and U2575 (N_2575,N_2217,N_2178);
nor U2576 (N_2576,N_2165,N_2194);
nand U2577 (N_2577,N_2146,N_2003);
and U2578 (N_2578,N_2019,N_2247);
nor U2579 (N_2579,N_2397,N_2496);
or U2580 (N_2580,N_2395,N_2408);
and U2581 (N_2581,N_2300,N_2349);
nor U2582 (N_2582,N_2332,N_2297);
or U2583 (N_2583,N_2173,N_2369);
nand U2584 (N_2584,N_2083,N_2412);
nand U2585 (N_2585,N_2090,N_2376);
or U2586 (N_2586,N_2021,N_2035);
nor U2587 (N_2587,N_2130,N_2031);
xor U2588 (N_2588,N_2033,N_2394);
and U2589 (N_2589,N_2338,N_2177);
nand U2590 (N_2590,N_2386,N_2119);
nand U2591 (N_2591,N_2185,N_2002);
nand U2592 (N_2592,N_2237,N_2042);
nand U2593 (N_2593,N_2429,N_2257);
nor U2594 (N_2594,N_2269,N_2134);
and U2595 (N_2595,N_2428,N_2348);
nand U2596 (N_2596,N_2476,N_2036);
nand U2597 (N_2597,N_2073,N_2097);
or U2598 (N_2598,N_2063,N_2104);
or U2599 (N_2599,N_2064,N_2158);
nand U2600 (N_2600,N_2460,N_2259);
or U2601 (N_2601,N_2241,N_2336);
nor U2602 (N_2602,N_2479,N_2325);
xor U2603 (N_2603,N_2361,N_2345);
or U2604 (N_2604,N_2148,N_2171);
or U2605 (N_2605,N_2316,N_2202);
nand U2606 (N_2606,N_2093,N_2215);
or U2607 (N_2607,N_2262,N_2495);
nand U2608 (N_2608,N_2467,N_2333);
nand U2609 (N_2609,N_2006,N_2406);
and U2610 (N_2610,N_2447,N_2278);
nand U2611 (N_2611,N_2087,N_2024);
nor U2612 (N_2612,N_2453,N_2143);
or U2613 (N_2613,N_2293,N_2029);
xnor U2614 (N_2614,N_2268,N_2422);
nor U2615 (N_2615,N_2225,N_2286);
nor U2616 (N_2616,N_2425,N_2228);
or U2617 (N_2617,N_2491,N_2478);
xor U2618 (N_2618,N_2008,N_2187);
or U2619 (N_2619,N_2209,N_2439);
or U2620 (N_2620,N_2308,N_2290);
or U2621 (N_2621,N_2277,N_2220);
nand U2622 (N_2622,N_2051,N_2121);
or U2623 (N_2623,N_2448,N_2102);
nor U2624 (N_2624,N_2313,N_2184);
nor U2625 (N_2625,N_2192,N_2497);
and U2626 (N_2626,N_2364,N_2047);
nor U2627 (N_2627,N_2393,N_2109);
nand U2628 (N_2628,N_2292,N_2078);
nand U2629 (N_2629,N_2074,N_2438);
nand U2630 (N_2630,N_2471,N_2168);
and U2631 (N_2631,N_2101,N_2426);
and U2632 (N_2632,N_2195,N_2309);
nor U2633 (N_2633,N_2315,N_2113);
nand U2634 (N_2634,N_2061,N_2039);
and U2635 (N_2635,N_2424,N_2396);
xor U2636 (N_2636,N_2155,N_2291);
nor U2637 (N_2637,N_2193,N_2283);
nor U2638 (N_2638,N_2069,N_2433);
nand U2639 (N_2639,N_2219,N_2374);
and U2640 (N_2640,N_2307,N_2080);
nand U2641 (N_2641,N_2295,N_2462);
nor U2642 (N_2642,N_2351,N_2049);
or U2643 (N_2643,N_2296,N_2157);
nand U2644 (N_2644,N_2287,N_2055);
or U2645 (N_2645,N_2298,N_2270);
xor U2646 (N_2646,N_2110,N_2387);
or U2647 (N_2647,N_2197,N_2028);
and U2648 (N_2648,N_2016,N_2362);
or U2649 (N_2649,N_2458,N_2203);
or U2650 (N_2650,N_2013,N_2274);
or U2651 (N_2651,N_2045,N_2343);
or U2652 (N_2652,N_2388,N_2329);
and U2653 (N_2653,N_2242,N_2421);
nand U2654 (N_2654,N_2245,N_2084);
nand U2655 (N_2655,N_2222,N_2264);
nand U2656 (N_2656,N_2123,N_2273);
nand U2657 (N_2657,N_2138,N_2365);
and U2658 (N_2658,N_2214,N_2383);
nor U2659 (N_2659,N_2179,N_2321);
and U2660 (N_2660,N_2229,N_2339);
nand U2661 (N_2661,N_2265,N_2133);
or U2662 (N_2662,N_2014,N_2302);
nand U2663 (N_2663,N_2120,N_2032);
and U2664 (N_2664,N_2054,N_2355);
nor U2665 (N_2665,N_2007,N_2303);
or U2666 (N_2666,N_2127,N_2282);
nor U2667 (N_2667,N_2432,N_2175);
or U2668 (N_2668,N_2483,N_2480);
and U2669 (N_2669,N_2196,N_2012);
or U2670 (N_2670,N_2156,N_2340);
and U2671 (N_2671,N_2100,N_2463);
nor U2672 (N_2672,N_2299,N_2404);
nand U2673 (N_2673,N_2075,N_2289);
nand U2674 (N_2674,N_2473,N_2067);
nand U2675 (N_2675,N_2312,N_2400);
nand U2676 (N_2676,N_2062,N_2417);
nand U2677 (N_2677,N_2056,N_2004);
nor U2678 (N_2678,N_2301,N_2180);
nor U2679 (N_2679,N_2410,N_2370);
nand U2680 (N_2680,N_2162,N_2239);
nand U2681 (N_2681,N_2353,N_2159);
or U2682 (N_2682,N_2451,N_2132);
nand U2683 (N_2683,N_2431,N_2377);
nor U2684 (N_2684,N_2350,N_2459);
nor U2685 (N_2685,N_2427,N_2413);
or U2686 (N_2686,N_2342,N_2401);
or U2687 (N_2687,N_2470,N_2129);
or U2688 (N_2688,N_2174,N_2223);
nor U2689 (N_2689,N_2423,N_2052);
nand U2690 (N_2690,N_2053,N_2189);
or U2691 (N_2691,N_2025,N_2234);
and U2692 (N_2692,N_2235,N_2385);
nor U2693 (N_2693,N_2088,N_2001);
nor U2694 (N_2694,N_2151,N_2294);
and U2695 (N_2695,N_2266,N_2494);
or U2696 (N_2696,N_2322,N_2103);
or U2697 (N_2697,N_2153,N_2116);
or U2698 (N_2698,N_2200,N_2172);
nor U2699 (N_2699,N_2346,N_2186);
nor U2700 (N_2700,N_2154,N_2238);
nand U2701 (N_2701,N_2461,N_2357);
nand U2702 (N_2702,N_2444,N_2095);
and U2703 (N_2703,N_2230,N_2212);
or U2704 (N_2704,N_2010,N_2070);
and U2705 (N_2705,N_2108,N_2190);
or U2706 (N_2706,N_2096,N_2250);
and U2707 (N_2707,N_2140,N_2255);
or U2708 (N_2708,N_2118,N_2020);
nor U2709 (N_2709,N_2213,N_2487);
nor U2710 (N_2710,N_2452,N_2356);
nor U2711 (N_2711,N_2464,N_2280);
or U2712 (N_2712,N_2330,N_2378);
nor U2713 (N_2713,N_2139,N_2201);
and U2714 (N_2714,N_2147,N_2232);
nand U2715 (N_2715,N_2320,N_2058);
or U2716 (N_2716,N_2204,N_2164);
nand U2717 (N_2717,N_2023,N_2288);
and U2718 (N_2718,N_2371,N_2107);
or U2719 (N_2719,N_2009,N_2254);
nand U2720 (N_2720,N_2405,N_2191);
nor U2721 (N_2721,N_2216,N_2092);
and U2722 (N_2722,N_2314,N_2482);
nor U2723 (N_2723,N_2368,N_2059);
nand U2724 (N_2724,N_2253,N_2490);
nand U2725 (N_2725,N_2381,N_2198);
nand U2726 (N_2726,N_2267,N_2011);
and U2727 (N_2727,N_2411,N_2034);
nor U2728 (N_2728,N_2128,N_2221);
xor U2729 (N_2729,N_2117,N_2135);
or U2730 (N_2730,N_2347,N_2477);
and U2731 (N_2731,N_2066,N_2082);
and U2732 (N_2732,N_2224,N_2493);
xor U2733 (N_2733,N_2486,N_2407);
or U2734 (N_2734,N_2469,N_2040);
nor U2735 (N_2735,N_2244,N_2091);
or U2736 (N_2736,N_2089,N_2465);
nand U2737 (N_2737,N_2456,N_2398);
and U2738 (N_2738,N_2170,N_2094);
or U2739 (N_2739,N_2466,N_2441);
nor U2740 (N_2740,N_2382,N_2017);
and U2741 (N_2741,N_2327,N_2391);
nor U2742 (N_2742,N_2435,N_2326);
nand U2743 (N_2743,N_2442,N_2256);
or U2744 (N_2744,N_2323,N_2207);
or U2745 (N_2745,N_2485,N_2167);
xor U2746 (N_2746,N_2455,N_2272);
or U2747 (N_2747,N_2352,N_2114);
nor U2748 (N_2748,N_2071,N_2418);
nor U2749 (N_2749,N_2420,N_2475);
nand U2750 (N_2750,N_2488,N_2462);
nand U2751 (N_2751,N_2294,N_2321);
nand U2752 (N_2752,N_2161,N_2175);
nand U2753 (N_2753,N_2358,N_2386);
or U2754 (N_2754,N_2010,N_2242);
and U2755 (N_2755,N_2007,N_2284);
nand U2756 (N_2756,N_2347,N_2331);
and U2757 (N_2757,N_2179,N_2177);
and U2758 (N_2758,N_2057,N_2403);
or U2759 (N_2759,N_2407,N_2374);
nand U2760 (N_2760,N_2391,N_2494);
nor U2761 (N_2761,N_2123,N_2280);
and U2762 (N_2762,N_2434,N_2364);
nor U2763 (N_2763,N_2417,N_2026);
nor U2764 (N_2764,N_2298,N_2312);
or U2765 (N_2765,N_2053,N_2412);
nor U2766 (N_2766,N_2166,N_2180);
or U2767 (N_2767,N_2262,N_2273);
nor U2768 (N_2768,N_2104,N_2490);
nor U2769 (N_2769,N_2210,N_2150);
and U2770 (N_2770,N_2099,N_2407);
and U2771 (N_2771,N_2424,N_2282);
or U2772 (N_2772,N_2113,N_2322);
nor U2773 (N_2773,N_2207,N_2494);
and U2774 (N_2774,N_2174,N_2145);
nand U2775 (N_2775,N_2133,N_2059);
nand U2776 (N_2776,N_2431,N_2221);
nand U2777 (N_2777,N_2174,N_2379);
nor U2778 (N_2778,N_2125,N_2213);
or U2779 (N_2779,N_2361,N_2145);
or U2780 (N_2780,N_2405,N_2466);
nor U2781 (N_2781,N_2017,N_2296);
and U2782 (N_2782,N_2301,N_2030);
nand U2783 (N_2783,N_2325,N_2054);
and U2784 (N_2784,N_2041,N_2349);
nand U2785 (N_2785,N_2017,N_2073);
or U2786 (N_2786,N_2373,N_2220);
and U2787 (N_2787,N_2407,N_2242);
nand U2788 (N_2788,N_2190,N_2444);
nor U2789 (N_2789,N_2453,N_2035);
nor U2790 (N_2790,N_2467,N_2103);
or U2791 (N_2791,N_2261,N_2456);
or U2792 (N_2792,N_2426,N_2151);
xnor U2793 (N_2793,N_2402,N_2245);
and U2794 (N_2794,N_2088,N_2424);
or U2795 (N_2795,N_2063,N_2190);
or U2796 (N_2796,N_2372,N_2085);
nand U2797 (N_2797,N_2280,N_2330);
and U2798 (N_2798,N_2214,N_2290);
or U2799 (N_2799,N_2490,N_2130);
nand U2800 (N_2800,N_2451,N_2458);
and U2801 (N_2801,N_2340,N_2365);
or U2802 (N_2802,N_2162,N_2212);
or U2803 (N_2803,N_2002,N_2123);
or U2804 (N_2804,N_2459,N_2362);
nor U2805 (N_2805,N_2307,N_2055);
nor U2806 (N_2806,N_2157,N_2449);
nand U2807 (N_2807,N_2247,N_2034);
or U2808 (N_2808,N_2170,N_2360);
nand U2809 (N_2809,N_2255,N_2468);
and U2810 (N_2810,N_2317,N_2478);
or U2811 (N_2811,N_2383,N_2096);
nor U2812 (N_2812,N_2167,N_2202);
or U2813 (N_2813,N_2057,N_2269);
nand U2814 (N_2814,N_2498,N_2157);
or U2815 (N_2815,N_2228,N_2316);
or U2816 (N_2816,N_2447,N_2045);
and U2817 (N_2817,N_2301,N_2254);
and U2818 (N_2818,N_2313,N_2435);
nand U2819 (N_2819,N_2085,N_2195);
and U2820 (N_2820,N_2008,N_2139);
and U2821 (N_2821,N_2221,N_2114);
and U2822 (N_2822,N_2085,N_2018);
nand U2823 (N_2823,N_2364,N_2208);
and U2824 (N_2824,N_2342,N_2109);
nor U2825 (N_2825,N_2047,N_2337);
and U2826 (N_2826,N_2234,N_2294);
and U2827 (N_2827,N_2054,N_2405);
nand U2828 (N_2828,N_2398,N_2315);
or U2829 (N_2829,N_2393,N_2465);
nand U2830 (N_2830,N_2000,N_2444);
or U2831 (N_2831,N_2258,N_2231);
or U2832 (N_2832,N_2311,N_2069);
or U2833 (N_2833,N_2229,N_2037);
or U2834 (N_2834,N_2344,N_2303);
nand U2835 (N_2835,N_2124,N_2429);
and U2836 (N_2836,N_2437,N_2444);
nand U2837 (N_2837,N_2467,N_2252);
or U2838 (N_2838,N_2283,N_2042);
or U2839 (N_2839,N_2232,N_2242);
nand U2840 (N_2840,N_2160,N_2327);
nand U2841 (N_2841,N_2217,N_2456);
and U2842 (N_2842,N_2302,N_2371);
nand U2843 (N_2843,N_2074,N_2280);
nand U2844 (N_2844,N_2294,N_2254);
nand U2845 (N_2845,N_2370,N_2036);
nor U2846 (N_2846,N_2085,N_2377);
nand U2847 (N_2847,N_2481,N_2147);
and U2848 (N_2848,N_2266,N_2289);
and U2849 (N_2849,N_2128,N_2407);
and U2850 (N_2850,N_2110,N_2211);
and U2851 (N_2851,N_2306,N_2390);
nand U2852 (N_2852,N_2365,N_2390);
or U2853 (N_2853,N_2042,N_2479);
and U2854 (N_2854,N_2471,N_2180);
or U2855 (N_2855,N_2379,N_2184);
nor U2856 (N_2856,N_2360,N_2338);
or U2857 (N_2857,N_2006,N_2135);
or U2858 (N_2858,N_2149,N_2302);
nor U2859 (N_2859,N_2061,N_2210);
and U2860 (N_2860,N_2468,N_2406);
and U2861 (N_2861,N_2044,N_2287);
nor U2862 (N_2862,N_2231,N_2492);
nand U2863 (N_2863,N_2288,N_2465);
or U2864 (N_2864,N_2312,N_2429);
nand U2865 (N_2865,N_2227,N_2264);
and U2866 (N_2866,N_2188,N_2397);
or U2867 (N_2867,N_2296,N_2338);
nor U2868 (N_2868,N_2294,N_2490);
and U2869 (N_2869,N_2340,N_2188);
nor U2870 (N_2870,N_2180,N_2293);
or U2871 (N_2871,N_2464,N_2094);
or U2872 (N_2872,N_2336,N_2265);
nor U2873 (N_2873,N_2224,N_2294);
or U2874 (N_2874,N_2398,N_2158);
nor U2875 (N_2875,N_2201,N_2460);
and U2876 (N_2876,N_2390,N_2355);
and U2877 (N_2877,N_2484,N_2238);
nand U2878 (N_2878,N_2452,N_2447);
nand U2879 (N_2879,N_2320,N_2469);
nor U2880 (N_2880,N_2459,N_2455);
nor U2881 (N_2881,N_2009,N_2191);
or U2882 (N_2882,N_2336,N_2032);
nor U2883 (N_2883,N_2250,N_2008);
or U2884 (N_2884,N_2082,N_2078);
nor U2885 (N_2885,N_2380,N_2227);
and U2886 (N_2886,N_2049,N_2407);
nand U2887 (N_2887,N_2421,N_2029);
nor U2888 (N_2888,N_2446,N_2267);
nand U2889 (N_2889,N_2184,N_2021);
and U2890 (N_2890,N_2340,N_2064);
and U2891 (N_2891,N_2356,N_2211);
and U2892 (N_2892,N_2254,N_2242);
and U2893 (N_2893,N_2166,N_2002);
and U2894 (N_2894,N_2366,N_2400);
and U2895 (N_2895,N_2409,N_2433);
nand U2896 (N_2896,N_2481,N_2128);
and U2897 (N_2897,N_2251,N_2021);
and U2898 (N_2898,N_2313,N_2247);
and U2899 (N_2899,N_2300,N_2113);
nand U2900 (N_2900,N_2460,N_2488);
and U2901 (N_2901,N_2479,N_2455);
nand U2902 (N_2902,N_2343,N_2059);
and U2903 (N_2903,N_2470,N_2040);
and U2904 (N_2904,N_2069,N_2499);
and U2905 (N_2905,N_2156,N_2224);
nand U2906 (N_2906,N_2012,N_2146);
and U2907 (N_2907,N_2185,N_2412);
and U2908 (N_2908,N_2021,N_2075);
and U2909 (N_2909,N_2381,N_2440);
nand U2910 (N_2910,N_2170,N_2070);
nor U2911 (N_2911,N_2062,N_2053);
or U2912 (N_2912,N_2179,N_2044);
nor U2913 (N_2913,N_2460,N_2497);
nand U2914 (N_2914,N_2257,N_2034);
nand U2915 (N_2915,N_2140,N_2370);
or U2916 (N_2916,N_2181,N_2499);
nor U2917 (N_2917,N_2067,N_2459);
and U2918 (N_2918,N_2348,N_2038);
and U2919 (N_2919,N_2348,N_2093);
or U2920 (N_2920,N_2050,N_2010);
and U2921 (N_2921,N_2029,N_2381);
or U2922 (N_2922,N_2344,N_2272);
xnor U2923 (N_2923,N_2345,N_2133);
or U2924 (N_2924,N_2375,N_2300);
nand U2925 (N_2925,N_2487,N_2439);
nor U2926 (N_2926,N_2214,N_2357);
nand U2927 (N_2927,N_2088,N_2326);
nand U2928 (N_2928,N_2119,N_2338);
nand U2929 (N_2929,N_2127,N_2168);
nand U2930 (N_2930,N_2224,N_2201);
nand U2931 (N_2931,N_2334,N_2456);
nand U2932 (N_2932,N_2436,N_2213);
nor U2933 (N_2933,N_2416,N_2467);
and U2934 (N_2934,N_2101,N_2226);
nor U2935 (N_2935,N_2025,N_2493);
xor U2936 (N_2936,N_2327,N_2401);
nor U2937 (N_2937,N_2070,N_2128);
nand U2938 (N_2938,N_2073,N_2120);
nor U2939 (N_2939,N_2328,N_2387);
or U2940 (N_2940,N_2493,N_2180);
nand U2941 (N_2941,N_2335,N_2058);
or U2942 (N_2942,N_2442,N_2288);
nor U2943 (N_2943,N_2348,N_2260);
nand U2944 (N_2944,N_2479,N_2122);
nand U2945 (N_2945,N_2489,N_2099);
or U2946 (N_2946,N_2469,N_2066);
or U2947 (N_2947,N_2031,N_2025);
and U2948 (N_2948,N_2260,N_2264);
nor U2949 (N_2949,N_2461,N_2286);
and U2950 (N_2950,N_2168,N_2061);
nand U2951 (N_2951,N_2492,N_2414);
and U2952 (N_2952,N_2091,N_2311);
xnor U2953 (N_2953,N_2355,N_2112);
nand U2954 (N_2954,N_2426,N_2352);
nand U2955 (N_2955,N_2388,N_2381);
nand U2956 (N_2956,N_2026,N_2455);
nor U2957 (N_2957,N_2227,N_2014);
nor U2958 (N_2958,N_2440,N_2425);
xnor U2959 (N_2959,N_2018,N_2390);
and U2960 (N_2960,N_2032,N_2389);
nor U2961 (N_2961,N_2032,N_2133);
nand U2962 (N_2962,N_2275,N_2041);
and U2963 (N_2963,N_2361,N_2146);
nor U2964 (N_2964,N_2317,N_2193);
and U2965 (N_2965,N_2287,N_2136);
or U2966 (N_2966,N_2194,N_2364);
and U2967 (N_2967,N_2256,N_2285);
and U2968 (N_2968,N_2324,N_2304);
nand U2969 (N_2969,N_2065,N_2450);
or U2970 (N_2970,N_2154,N_2418);
and U2971 (N_2971,N_2193,N_2498);
or U2972 (N_2972,N_2062,N_2120);
nand U2973 (N_2973,N_2153,N_2306);
or U2974 (N_2974,N_2268,N_2343);
and U2975 (N_2975,N_2302,N_2108);
and U2976 (N_2976,N_2434,N_2350);
or U2977 (N_2977,N_2478,N_2345);
nand U2978 (N_2978,N_2422,N_2359);
and U2979 (N_2979,N_2347,N_2315);
nor U2980 (N_2980,N_2131,N_2359);
and U2981 (N_2981,N_2374,N_2211);
or U2982 (N_2982,N_2024,N_2417);
nand U2983 (N_2983,N_2208,N_2448);
or U2984 (N_2984,N_2419,N_2471);
nor U2985 (N_2985,N_2289,N_2207);
and U2986 (N_2986,N_2221,N_2373);
and U2987 (N_2987,N_2117,N_2418);
nand U2988 (N_2988,N_2283,N_2372);
nand U2989 (N_2989,N_2401,N_2185);
or U2990 (N_2990,N_2438,N_2061);
and U2991 (N_2991,N_2335,N_2485);
nand U2992 (N_2992,N_2184,N_2129);
or U2993 (N_2993,N_2037,N_2107);
and U2994 (N_2994,N_2205,N_2345);
and U2995 (N_2995,N_2244,N_2095);
nand U2996 (N_2996,N_2383,N_2201);
nor U2997 (N_2997,N_2381,N_2032);
nor U2998 (N_2998,N_2051,N_2300);
or U2999 (N_2999,N_2118,N_2054);
nor U3000 (N_3000,N_2835,N_2887);
nor U3001 (N_3001,N_2995,N_2939);
and U3002 (N_3002,N_2719,N_2631);
nand U3003 (N_3003,N_2564,N_2985);
nor U3004 (N_3004,N_2685,N_2531);
nand U3005 (N_3005,N_2851,N_2525);
nor U3006 (N_3006,N_2524,N_2867);
nand U3007 (N_3007,N_2506,N_2670);
and U3008 (N_3008,N_2639,N_2892);
nor U3009 (N_3009,N_2736,N_2658);
or U3010 (N_3010,N_2630,N_2712);
nand U3011 (N_3011,N_2881,N_2842);
nand U3012 (N_3012,N_2581,N_2812);
or U3013 (N_3013,N_2928,N_2923);
or U3014 (N_3014,N_2596,N_2759);
and U3015 (N_3015,N_2694,N_2772);
or U3016 (N_3016,N_2529,N_2954);
nand U3017 (N_3017,N_2882,N_2557);
or U3018 (N_3018,N_2864,N_2782);
nor U3019 (N_3019,N_2763,N_2755);
and U3020 (N_3020,N_2587,N_2921);
and U3021 (N_3021,N_2951,N_2507);
nand U3022 (N_3022,N_2542,N_2547);
nor U3023 (N_3023,N_2827,N_2967);
nand U3024 (N_3024,N_2559,N_2811);
and U3025 (N_3025,N_2614,N_2555);
or U3026 (N_3026,N_2808,N_2901);
nor U3027 (N_3027,N_2570,N_2907);
nand U3028 (N_3028,N_2909,N_2643);
and U3029 (N_3029,N_2737,N_2747);
nor U3030 (N_3030,N_2624,N_2538);
nor U3031 (N_3031,N_2863,N_2699);
nor U3032 (N_3032,N_2980,N_2688);
nor U3033 (N_3033,N_2611,N_2689);
nor U3034 (N_3034,N_2974,N_2945);
and U3035 (N_3035,N_2791,N_2682);
or U3036 (N_3036,N_2522,N_2979);
nand U3037 (N_3037,N_2621,N_2528);
or U3038 (N_3038,N_2937,N_2815);
nor U3039 (N_3039,N_2911,N_2599);
nand U3040 (N_3040,N_2641,N_2511);
and U3041 (N_3041,N_2657,N_2577);
nor U3042 (N_3042,N_2710,N_2698);
and U3043 (N_3043,N_2852,N_2584);
nand U3044 (N_3044,N_2833,N_2927);
and U3045 (N_3045,N_2595,N_2801);
nand U3046 (N_3046,N_2561,N_2874);
nor U3047 (N_3047,N_2647,N_2947);
nand U3048 (N_3048,N_2862,N_2848);
nand U3049 (N_3049,N_2563,N_2935);
nor U3050 (N_3050,N_2588,N_2975);
and U3051 (N_3051,N_2798,N_2743);
and U3052 (N_3052,N_2741,N_2948);
nor U3053 (N_3053,N_2725,N_2600);
nor U3054 (N_3054,N_2854,N_2970);
nor U3055 (N_3055,N_2777,N_2664);
or U3056 (N_3056,N_2706,N_2604);
nor U3057 (N_3057,N_2780,N_2805);
nand U3058 (N_3058,N_2635,N_2950);
and U3059 (N_3059,N_2671,N_2943);
nand U3060 (N_3060,N_2558,N_2625);
and U3061 (N_3061,N_2649,N_2873);
xnor U3062 (N_3062,N_2830,N_2758);
and U3063 (N_3063,N_2819,N_2549);
and U3064 (N_3064,N_2952,N_2748);
and U3065 (N_3065,N_2971,N_2983);
nor U3066 (N_3066,N_2836,N_2728);
and U3067 (N_3067,N_2821,N_2783);
nand U3068 (N_3068,N_2556,N_2716);
nor U3069 (N_3069,N_2990,N_2606);
nor U3070 (N_3070,N_2828,N_2590);
and U3071 (N_3071,N_2615,N_2638);
and U3072 (N_3072,N_2769,N_2825);
nor U3073 (N_3073,N_2857,N_2778);
and U3074 (N_3074,N_2695,N_2964);
nor U3075 (N_3075,N_2543,N_2930);
and U3076 (N_3076,N_2724,N_2510);
nand U3077 (N_3077,N_2905,N_2788);
nand U3078 (N_3078,N_2541,N_2884);
nor U3079 (N_3079,N_2966,N_2997);
nor U3080 (N_3080,N_2775,N_2608);
nor U3081 (N_3081,N_2767,N_2749);
and U3082 (N_3082,N_2917,N_2687);
nor U3083 (N_3083,N_2790,N_2727);
or U3084 (N_3084,N_2899,N_2554);
or U3085 (N_3085,N_2508,N_2855);
nor U3086 (N_3086,N_2505,N_2626);
nand U3087 (N_3087,N_2871,N_2802);
or U3088 (N_3088,N_2700,N_2822);
and U3089 (N_3089,N_2679,N_2770);
nand U3090 (N_3090,N_2771,N_2675);
nand U3091 (N_3091,N_2886,N_2677);
or U3092 (N_3092,N_2942,N_2589);
and U3093 (N_3093,N_2681,N_2612);
nor U3094 (N_3094,N_2580,N_2651);
nor U3095 (N_3095,N_2504,N_2940);
nand U3096 (N_3096,N_2585,N_2969);
nor U3097 (N_3097,N_2953,N_2718);
nand U3098 (N_3098,N_2645,N_2768);
and U3099 (N_3099,N_2539,N_2934);
and U3100 (N_3100,N_2594,N_2797);
and U3101 (N_3101,N_2617,N_2846);
and U3102 (N_3102,N_2824,N_2931);
nor U3103 (N_3103,N_2799,N_2691);
nand U3104 (N_3104,N_2922,N_2839);
nor U3105 (N_3105,N_2779,N_2904);
and U3106 (N_3106,N_2762,N_2894);
or U3107 (N_3107,N_2629,N_2655);
xnor U3108 (N_3108,N_2800,N_2784);
and U3109 (N_3109,N_2684,N_2620);
and U3110 (N_3110,N_2929,N_2571);
and U3111 (N_3111,N_2832,N_2517);
nor U3112 (N_3112,N_2591,N_2959);
and U3113 (N_3113,N_2750,N_2793);
nand U3114 (N_3114,N_2602,N_2903);
or U3115 (N_3115,N_2733,N_2744);
and U3116 (N_3116,N_2692,N_2708);
nor U3117 (N_3117,N_2521,N_2721);
and U3118 (N_3118,N_2659,N_2993);
and U3119 (N_3119,N_2740,N_2515);
nand U3120 (N_3120,N_2807,N_2958);
nand U3121 (N_3121,N_2598,N_2877);
or U3122 (N_3122,N_2636,N_2876);
or U3123 (N_3123,N_2502,N_2526);
nor U3124 (N_3124,N_2787,N_2984);
xor U3125 (N_3125,N_2880,N_2560);
nor U3126 (N_3126,N_2723,N_2709);
or U3127 (N_3127,N_2715,N_2583);
or U3128 (N_3128,N_2567,N_2856);
or U3129 (N_3129,N_2656,N_2616);
or U3130 (N_3130,N_2789,N_2582);
nand U3131 (N_3131,N_2713,N_2916);
nor U3132 (N_3132,N_2633,N_2720);
nor U3133 (N_3133,N_2760,N_2924);
or U3134 (N_3134,N_2757,N_2912);
nand U3135 (N_3135,N_2756,N_2513);
nand U3136 (N_3136,N_2965,N_2796);
nor U3137 (N_3137,N_2761,N_2628);
and U3138 (N_3138,N_2902,N_2705);
xnor U3139 (N_3139,N_2622,N_2870);
or U3140 (N_3140,N_2861,N_2509);
xor U3141 (N_3141,N_2996,N_2673);
or U3142 (N_3142,N_2774,N_2910);
and U3143 (N_3143,N_2663,N_2512);
nand U3144 (N_3144,N_2500,N_2652);
nor U3145 (N_3145,N_2878,N_2860);
nor U3146 (N_3146,N_2586,N_2773);
nor U3147 (N_3147,N_2781,N_2785);
nor U3148 (N_3148,N_2764,N_2674);
nor U3149 (N_3149,N_2534,N_2562);
or U3150 (N_3150,N_2976,N_2890);
nand U3151 (N_3151,N_2932,N_2661);
or U3152 (N_3152,N_2820,N_2941);
nand U3153 (N_3153,N_2955,N_2765);
nor U3154 (N_3154,N_2806,N_2804);
or U3155 (N_3155,N_2667,N_2690);
or U3156 (N_3156,N_2944,N_2566);
nor U3157 (N_3157,N_2883,N_2746);
nor U3158 (N_3158,N_2516,N_2742);
nor U3159 (N_3159,N_2546,N_2988);
nand U3160 (N_3160,N_2838,N_2915);
or U3161 (N_3161,N_2540,N_2888);
and U3162 (N_3162,N_2869,N_2841);
nor U3163 (N_3163,N_2738,N_2704);
nand U3164 (N_3164,N_2726,N_2813);
and U3165 (N_3165,N_2607,N_2623);
nor U3166 (N_3166,N_2837,N_2662);
or U3167 (N_3167,N_2532,N_2933);
nor U3168 (N_3168,N_2578,N_2696);
nor U3169 (N_3169,N_2537,N_2654);
nor U3170 (N_3170,N_2613,N_2722);
nand U3171 (N_3171,N_2730,N_2994);
or U3172 (N_3172,N_2701,N_2527);
and U3173 (N_3173,N_2752,N_2579);
or U3174 (N_3174,N_2794,N_2568);
and U3175 (N_3175,N_2575,N_2702);
and U3176 (N_3176,N_2850,N_2735);
and U3177 (N_3177,N_2918,N_2981);
nand U3178 (N_3178,N_2593,N_2866);
nor U3179 (N_3179,N_2550,N_2786);
nor U3180 (N_3180,N_2703,N_2792);
and U3181 (N_3181,N_2938,N_2501);
and U3182 (N_3182,N_2987,N_2919);
nand U3183 (N_3183,N_2810,N_2977);
nand U3184 (N_3184,N_2574,N_2648);
nand U3185 (N_3185,N_2572,N_2900);
and U3186 (N_3186,N_2551,N_2666);
or U3187 (N_3187,N_2520,N_2503);
nand U3188 (N_3188,N_2989,N_2686);
or U3189 (N_3189,N_2669,N_2707);
nor U3190 (N_3190,N_2518,N_2535);
and U3191 (N_3191,N_2889,N_2961);
nand U3192 (N_3192,N_2978,N_2717);
nor U3193 (N_3193,N_2803,N_2729);
and U3194 (N_3194,N_2795,N_2597);
and U3195 (N_3195,N_2847,N_2817);
or U3196 (N_3196,N_2968,N_2816);
nand U3197 (N_3197,N_2553,N_2766);
or U3198 (N_3198,N_2678,N_2859);
nor U3199 (N_3199,N_2734,N_2920);
nand U3200 (N_3200,N_2893,N_2896);
nor U3201 (N_3201,N_2936,N_2569);
nor U3202 (N_3202,N_2642,N_2872);
and U3203 (N_3203,N_2697,N_2680);
and U3204 (N_3204,N_2676,N_2897);
and U3205 (N_3205,N_2868,N_2530);
nor U3206 (N_3206,N_2627,N_2865);
nand U3207 (N_3207,N_2536,N_2637);
nand U3208 (N_3208,N_2834,N_2545);
nor U3209 (N_3209,N_2831,N_2573);
nor U3210 (N_3210,N_2660,N_2925);
and U3211 (N_3211,N_2845,N_2853);
nand U3212 (N_3212,N_2818,N_2653);
nor U3213 (N_3213,N_2998,N_2946);
and U3214 (N_3214,N_2672,N_2895);
and U3215 (N_3215,N_2731,N_2523);
nand U3216 (N_3216,N_2960,N_2849);
and U3217 (N_3217,N_2809,N_2814);
and U3218 (N_3218,N_2514,N_2844);
nand U3219 (N_3219,N_2732,N_2533);
nand U3220 (N_3220,N_2739,N_2972);
nor U3221 (N_3221,N_2962,N_2576);
nand U3222 (N_3222,N_2665,N_2693);
nand U3223 (N_3223,N_2683,N_2605);
nand U3224 (N_3224,N_2823,N_2949);
xnor U3225 (N_3225,N_2829,N_2544);
and U3226 (N_3226,N_2618,N_2906);
nor U3227 (N_3227,N_2875,N_2634);
nor U3228 (N_3228,N_2603,N_2552);
nor U3229 (N_3229,N_2986,N_2898);
nand U3230 (N_3230,N_2963,N_2632);
nor U3231 (N_3231,N_2711,N_2519);
and U3232 (N_3232,N_2914,N_2991);
nand U3233 (N_3233,N_2957,N_2601);
nand U3234 (N_3234,N_2982,N_2714);
nand U3235 (N_3235,N_2565,N_2644);
and U3236 (N_3236,N_2646,N_2826);
or U3237 (N_3237,N_2592,N_2913);
or U3238 (N_3238,N_2609,N_2753);
xor U3239 (N_3239,N_2776,N_2891);
and U3240 (N_3240,N_2999,N_2956);
nand U3241 (N_3241,N_2885,N_2754);
xnor U3242 (N_3242,N_2610,N_2640);
nand U3243 (N_3243,N_2548,N_2843);
nor U3244 (N_3244,N_2619,N_2751);
nor U3245 (N_3245,N_2668,N_2650);
or U3246 (N_3246,N_2908,N_2926);
or U3247 (N_3247,N_2879,N_2745);
or U3248 (N_3248,N_2858,N_2973);
and U3249 (N_3249,N_2992,N_2840);
nor U3250 (N_3250,N_2890,N_2752);
or U3251 (N_3251,N_2824,N_2562);
or U3252 (N_3252,N_2661,N_2946);
nand U3253 (N_3253,N_2515,N_2594);
and U3254 (N_3254,N_2602,N_2761);
or U3255 (N_3255,N_2582,N_2710);
nand U3256 (N_3256,N_2696,N_2635);
and U3257 (N_3257,N_2739,N_2967);
and U3258 (N_3258,N_2974,N_2663);
and U3259 (N_3259,N_2903,N_2979);
or U3260 (N_3260,N_2616,N_2576);
or U3261 (N_3261,N_2826,N_2818);
nand U3262 (N_3262,N_2557,N_2692);
or U3263 (N_3263,N_2852,N_2727);
or U3264 (N_3264,N_2981,N_2938);
nand U3265 (N_3265,N_2574,N_2862);
or U3266 (N_3266,N_2847,N_2897);
nand U3267 (N_3267,N_2636,N_2731);
xnor U3268 (N_3268,N_2923,N_2572);
or U3269 (N_3269,N_2601,N_2863);
nor U3270 (N_3270,N_2523,N_2889);
nor U3271 (N_3271,N_2612,N_2601);
and U3272 (N_3272,N_2538,N_2802);
or U3273 (N_3273,N_2701,N_2986);
nand U3274 (N_3274,N_2731,N_2503);
and U3275 (N_3275,N_2528,N_2712);
xor U3276 (N_3276,N_2920,N_2757);
xnor U3277 (N_3277,N_2648,N_2604);
or U3278 (N_3278,N_2780,N_2559);
and U3279 (N_3279,N_2622,N_2979);
or U3280 (N_3280,N_2721,N_2979);
nand U3281 (N_3281,N_2974,N_2859);
nor U3282 (N_3282,N_2520,N_2528);
nand U3283 (N_3283,N_2924,N_2723);
and U3284 (N_3284,N_2818,N_2909);
nor U3285 (N_3285,N_2893,N_2824);
nand U3286 (N_3286,N_2609,N_2767);
or U3287 (N_3287,N_2698,N_2868);
or U3288 (N_3288,N_2807,N_2604);
nand U3289 (N_3289,N_2777,N_2634);
nand U3290 (N_3290,N_2712,N_2670);
and U3291 (N_3291,N_2808,N_2935);
and U3292 (N_3292,N_2586,N_2724);
nand U3293 (N_3293,N_2835,N_2955);
or U3294 (N_3294,N_2763,N_2622);
and U3295 (N_3295,N_2527,N_2756);
and U3296 (N_3296,N_2898,N_2595);
or U3297 (N_3297,N_2953,N_2508);
and U3298 (N_3298,N_2734,N_2603);
or U3299 (N_3299,N_2910,N_2624);
or U3300 (N_3300,N_2947,N_2811);
nor U3301 (N_3301,N_2586,N_2672);
and U3302 (N_3302,N_2781,N_2680);
nand U3303 (N_3303,N_2655,N_2509);
and U3304 (N_3304,N_2984,N_2591);
nor U3305 (N_3305,N_2570,N_2879);
or U3306 (N_3306,N_2588,N_2613);
nand U3307 (N_3307,N_2966,N_2641);
and U3308 (N_3308,N_2733,N_2865);
or U3309 (N_3309,N_2556,N_2968);
and U3310 (N_3310,N_2742,N_2668);
and U3311 (N_3311,N_2763,N_2841);
nor U3312 (N_3312,N_2539,N_2565);
or U3313 (N_3313,N_2687,N_2722);
or U3314 (N_3314,N_2854,N_2550);
nand U3315 (N_3315,N_2803,N_2884);
nand U3316 (N_3316,N_2657,N_2987);
nand U3317 (N_3317,N_2852,N_2598);
and U3318 (N_3318,N_2735,N_2868);
nand U3319 (N_3319,N_2680,N_2570);
and U3320 (N_3320,N_2592,N_2533);
and U3321 (N_3321,N_2722,N_2818);
nor U3322 (N_3322,N_2512,N_2777);
nor U3323 (N_3323,N_2680,N_2862);
and U3324 (N_3324,N_2891,N_2786);
nand U3325 (N_3325,N_2566,N_2715);
nand U3326 (N_3326,N_2919,N_2560);
nand U3327 (N_3327,N_2947,N_2532);
and U3328 (N_3328,N_2661,N_2958);
nor U3329 (N_3329,N_2646,N_2992);
nor U3330 (N_3330,N_2630,N_2624);
or U3331 (N_3331,N_2640,N_2643);
or U3332 (N_3332,N_2776,N_2811);
or U3333 (N_3333,N_2896,N_2638);
nor U3334 (N_3334,N_2758,N_2764);
nand U3335 (N_3335,N_2613,N_2639);
nor U3336 (N_3336,N_2929,N_2983);
and U3337 (N_3337,N_2805,N_2853);
nand U3338 (N_3338,N_2752,N_2592);
nand U3339 (N_3339,N_2756,N_2954);
and U3340 (N_3340,N_2728,N_2802);
or U3341 (N_3341,N_2699,N_2661);
nand U3342 (N_3342,N_2545,N_2636);
and U3343 (N_3343,N_2639,N_2587);
nor U3344 (N_3344,N_2545,N_2745);
or U3345 (N_3345,N_2525,N_2501);
nor U3346 (N_3346,N_2956,N_2963);
or U3347 (N_3347,N_2994,N_2639);
or U3348 (N_3348,N_2760,N_2603);
nor U3349 (N_3349,N_2998,N_2606);
nand U3350 (N_3350,N_2853,N_2949);
and U3351 (N_3351,N_2803,N_2954);
nor U3352 (N_3352,N_2688,N_2917);
nand U3353 (N_3353,N_2817,N_2691);
and U3354 (N_3354,N_2943,N_2617);
nor U3355 (N_3355,N_2684,N_2985);
nor U3356 (N_3356,N_2711,N_2959);
and U3357 (N_3357,N_2972,N_2804);
or U3358 (N_3358,N_2819,N_2856);
nand U3359 (N_3359,N_2542,N_2594);
or U3360 (N_3360,N_2860,N_2803);
nor U3361 (N_3361,N_2740,N_2640);
nand U3362 (N_3362,N_2623,N_2998);
nor U3363 (N_3363,N_2576,N_2968);
and U3364 (N_3364,N_2951,N_2681);
or U3365 (N_3365,N_2577,N_2593);
xor U3366 (N_3366,N_2655,N_2742);
nand U3367 (N_3367,N_2850,N_2671);
nor U3368 (N_3368,N_2584,N_2755);
or U3369 (N_3369,N_2742,N_2608);
nand U3370 (N_3370,N_2800,N_2961);
or U3371 (N_3371,N_2780,N_2522);
nand U3372 (N_3372,N_2835,N_2622);
nor U3373 (N_3373,N_2939,N_2614);
and U3374 (N_3374,N_2993,N_2976);
nand U3375 (N_3375,N_2527,N_2618);
and U3376 (N_3376,N_2789,N_2854);
nor U3377 (N_3377,N_2727,N_2935);
or U3378 (N_3378,N_2782,N_2798);
nor U3379 (N_3379,N_2935,N_2604);
or U3380 (N_3380,N_2999,N_2678);
or U3381 (N_3381,N_2782,N_2922);
nor U3382 (N_3382,N_2824,N_2706);
or U3383 (N_3383,N_2799,N_2670);
or U3384 (N_3384,N_2730,N_2999);
nor U3385 (N_3385,N_2883,N_2817);
nor U3386 (N_3386,N_2791,N_2992);
nand U3387 (N_3387,N_2714,N_2923);
nor U3388 (N_3388,N_2881,N_2685);
nand U3389 (N_3389,N_2916,N_2721);
or U3390 (N_3390,N_2789,N_2989);
nor U3391 (N_3391,N_2508,N_2720);
and U3392 (N_3392,N_2964,N_2981);
and U3393 (N_3393,N_2600,N_2618);
and U3394 (N_3394,N_2747,N_2652);
and U3395 (N_3395,N_2963,N_2805);
nand U3396 (N_3396,N_2604,N_2906);
nand U3397 (N_3397,N_2723,N_2919);
and U3398 (N_3398,N_2822,N_2667);
nand U3399 (N_3399,N_2594,N_2698);
nor U3400 (N_3400,N_2857,N_2776);
nor U3401 (N_3401,N_2722,N_2583);
nor U3402 (N_3402,N_2703,N_2520);
and U3403 (N_3403,N_2947,N_2535);
nor U3404 (N_3404,N_2823,N_2912);
and U3405 (N_3405,N_2827,N_2888);
nor U3406 (N_3406,N_2884,N_2825);
and U3407 (N_3407,N_2624,N_2718);
and U3408 (N_3408,N_2545,N_2662);
and U3409 (N_3409,N_2592,N_2685);
or U3410 (N_3410,N_2990,N_2505);
nor U3411 (N_3411,N_2891,N_2841);
and U3412 (N_3412,N_2568,N_2831);
nand U3413 (N_3413,N_2895,N_2984);
or U3414 (N_3414,N_2957,N_2706);
and U3415 (N_3415,N_2750,N_2723);
nor U3416 (N_3416,N_2555,N_2810);
nor U3417 (N_3417,N_2501,N_2889);
nand U3418 (N_3418,N_2607,N_2978);
nand U3419 (N_3419,N_2558,N_2686);
and U3420 (N_3420,N_2820,N_2566);
nor U3421 (N_3421,N_2643,N_2780);
or U3422 (N_3422,N_2500,N_2922);
nand U3423 (N_3423,N_2908,N_2649);
or U3424 (N_3424,N_2988,N_2575);
and U3425 (N_3425,N_2927,N_2806);
nand U3426 (N_3426,N_2947,N_2910);
nor U3427 (N_3427,N_2639,N_2729);
and U3428 (N_3428,N_2619,N_2587);
and U3429 (N_3429,N_2780,N_2563);
or U3430 (N_3430,N_2635,N_2612);
or U3431 (N_3431,N_2657,N_2681);
and U3432 (N_3432,N_2721,N_2978);
nand U3433 (N_3433,N_2733,N_2835);
or U3434 (N_3434,N_2911,N_2571);
nor U3435 (N_3435,N_2691,N_2704);
nand U3436 (N_3436,N_2620,N_2550);
nor U3437 (N_3437,N_2596,N_2507);
xor U3438 (N_3438,N_2709,N_2953);
and U3439 (N_3439,N_2671,N_2754);
nand U3440 (N_3440,N_2700,N_2711);
and U3441 (N_3441,N_2830,N_2800);
nor U3442 (N_3442,N_2663,N_2507);
xor U3443 (N_3443,N_2950,N_2561);
or U3444 (N_3444,N_2983,N_2755);
or U3445 (N_3445,N_2542,N_2911);
nor U3446 (N_3446,N_2500,N_2901);
or U3447 (N_3447,N_2550,N_2856);
or U3448 (N_3448,N_2502,N_2879);
and U3449 (N_3449,N_2601,N_2627);
and U3450 (N_3450,N_2688,N_2634);
nand U3451 (N_3451,N_2874,N_2530);
and U3452 (N_3452,N_2562,N_2890);
or U3453 (N_3453,N_2735,N_2709);
or U3454 (N_3454,N_2657,N_2958);
or U3455 (N_3455,N_2513,N_2581);
nand U3456 (N_3456,N_2592,N_2660);
nand U3457 (N_3457,N_2951,N_2909);
nor U3458 (N_3458,N_2545,N_2953);
and U3459 (N_3459,N_2819,N_2875);
nor U3460 (N_3460,N_2566,N_2852);
nor U3461 (N_3461,N_2664,N_2672);
or U3462 (N_3462,N_2816,N_2929);
and U3463 (N_3463,N_2501,N_2786);
and U3464 (N_3464,N_2779,N_2710);
or U3465 (N_3465,N_2832,N_2653);
nor U3466 (N_3466,N_2797,N_2974);
or U3467 (N_3467,N_2694,N_2911);
or U3468 (N_3468,N_2597,N_2730);
nand U3469 (N_3469,N_2559,N_2722);
or U3470 (N_3470,N_2914,N_2668);
and U3471 (N_3471,N_2829,N_2518);
and U3472 (N_3472,N_2822,N_2799);
nor U3473 (N_3473,N_2771,N_2598);
or U3474 (N_3474,N_2863,N_2778);
or U3475 (N_3475,N_2937,N_2603);
nor U3476 (N_3476,N_2690,N_2947);
nand U3477 (N_3477,N_2668,N_2800);
or U3478 (N_3478,N_2941,N_2672);
nor U3479 (N_3479,N_2720,N_2763);
or U3480 (N_3480,N_2915,N_2936);
or U3481 (N_3481,N_2805,N_2854);
and U3482 (N_3482,N_2634,N_2969);
xor U3483 (N_3483,N_2991,N_2759);
nor U3484 (N_3484,N_2833,N_2673);
nor U3485 (N_3485,N_2787,N_2812);
nand U3486 (N_3486,N_2781,N_2834);
xor U3487 (N_3487,N_2747,N_2660);
nand U3488 (N_3488,N_2926,N_2674);
nand U3489 (N_3489,N_2920,N_2834);
nand U3490 (N_3490,N_2811,N_2815);
nand U3491 (N_3491,N_2549,N_2514);
or U3492 (N_3492,N_2825,N_2881);
and U3493 (N_3493,N_2744,N_2516);
nand U3494 (N_3494,N_2841,N_2567);
nand U3495 (N_3495,N_2688,N_2752);
nor U3496 (N_3496,N_2558,N_2539);
nor U3497 (N_3497,N_2976,N_2560);
xnor U3498 (N_3498,N_2754,N_2559);
nand U3499 (N_3499,N_2949,N_2513);
and U3500 (N_3500,N_3195,N_3141);
and U3501 (N_3501,N_3377,N_3152);
and U3502 (N_3502,N_3113,N_3043);
or U3503 (N_3503,N_3037,N_3083);
or U3504 (N_3504,N_3451,N_3349);
and U3505 (N_3505,N_3351,N_3208);
nand U3506 (N_3506,N_3173,N_3347);
nor U3507 (N_3507,N_3375,N_3134);
nor U3508 (N_3508,N_3327,N_3336);
or U3509 (N_3509,N_3243,N_3312);
nor U3510 (N_3510,N_3096,N_3398);
or U3511 (N_3511,N_3416,N_3474);
nand U3512 (N_3512,N_3034,N_3009);
or U3513 (N_3513,N_3486,N_3198);
nor U3514 (N_3514,N_3216,N_3240);
nand U3515 (N_3515,N_3437,N_3420);
and U3516 (N_3516,N_3103,N_3084);
or U3517 (N_3517,N_3039,N_3245);
or U3518 (N_3518,N_3030,N_3180);
nor U3519 (N_3519,N_3058,N_3361);
or U3520 (N_3520,N_3256,N_3135);
or U3521 (N_3521,N_3406,N_3476);
or U3522 (N_3522,N_3425,N_3226);
nand U3523 (N_3523,N_3203,N_3271);
xor U3524 (N_3524,N_3223,N_3032);
and U3525 (N_3525,N_3081,N_3296);
or U3526 (N_3526,N_3333,N_3162);
nand U3527 (N_3527,N_3005,N_3038);
xor U3528 (N_3528,N_3066,N_3370);
and U3529 (N_3529,N_3069,N_3379);
nand U3530 (N_3530,N_3497,N_3063);
nand U3531 (N_3531,N_3130,N_3329);
nor U3532 (N_3532,N_3093,N_3491);
nor U3533 (N_3533,N_3239,N_3443);
or U3534 (N_3534,N_3111,N_3316);
nand U3535 (N_3535,N_3222,N_3232);
nor U3536 (N_3536,N_3214,N_3348);
and U3537 (N_3537,N_3026,N_3138);
or U3538 (N_3538,N_3405,N_3384);
nor U3539 (N_3539,N_3422,N_3429);
and U3540 (N_3540,N_3234,N_3300);
nand U3541 (N_3541,N_3006,N_3164);
and U3542 (N_3542,N_3448,N_3190);
and U3543 (N_3543,N_3188,N_3343);
nand U3544 (N_3544,N_3498,N_3309);
or U3545 (N_3545,N_3447,N_3261);
and U3546 (N_3546,N_3494,N_3206);
nand U3547 (N_3547,N_3260,N_3335);
nor U3548 (N_3548,N_3272,N_3076);
nand U3549 (N_3549,N_3374,N_3266);
nor U3550 (N_3550,N_3295,N_3358);
nor U3551 (N_3551,N_3326,N_3465);
and U3552 (N_3552,N_3044,N_3231);
or U3553 (N_3553,N_3079,N_3059);
nand U3554 (N_3554,N_3145,N_3082);
and U3555 (N_3555,N_3244,N_3072);
nor U3556 (N_3556,N_3022,N_3142);
or U3557 (N_3557,N_3487,N_3159);
or U3558 (N_3558,N_3464,N_3478);
nor U3559 (N_3559,N_3047,N_3191);
nor U3560 (N_3560,N_3495,N_3391);
or U3561 (N_3561,N_3105,N_3403);
xnor U3562 (N_3562,N_3182,N_3467);
or U3563 (N_3563,N_3408,N_3383);
nand U3564 (N_3564,N_3115,N_3049);
or U3565 (N_3565,N_3284,N_3364);
or U3566 (N_3566,N_3036,N_3041);
or U3567 (N_3567,N_3492,N_3373);
nor U3568 (N_3568,N_3479,N_3359);
or U3569 (N_3569,N_3340,N_3259);
or U3570 (N_3570,N_3366,N_3046);
or U3571 (N_3571,N_3227,N_3167);
or U3572 (N_3572,N_3303,N_3482);
or U3573 (N_3573,N_3118,N_3166);
nor U3574 (N_3574,N_3413,N_3017);
or U3575 (N_3575,N_3453,N_3278);
and U3576 (N_3576,N_3215,N_3251);
nand U3577 (N_3577,N_3354,N_3293);
nand U3578 (N_3578,N_3485,N_3014);
xor U3579 (N_3579,N_3472,N_3169);
and U3580 (N_3580,N_3407,N_3207);
and U3581 (N_3581,N_3378,N_3094);
xnor U3582 (N_3582,N_3337,N_3064);
and U3583 (N_3583,N_3427,N_3099);
and U3584 (N_3584,N_3328,N_3107);
or U3585 (N_3585,N_3102,N_3496);
nor U3586 (N_3586,N_3025,N_3357);
or U3587 (N_3587,N_3291,N_3139);
and U3588 (N_3588,N_3362,N_3010);
and U3589 (N_3589,N_3268,N_3225);
nor U3590 (N_3590,N_3133,N_3459);
and U3591 (N_3591,N_3089,N_3339);
nand U3592 (N_3592,N_3050,N_3338);
or U3593 (N_3593,N_3299,N_3153);
and U3594 (N_3594,N_3477,N_3365);
nand U3595 (N_3595,N_3192,N_3000);
nand U3596 (N_3596,N_3051,N_3092);
nor U3597 (N_3597,N_3247,N_3021);
nor U3598 (N_3598,N_3062,N_3288);
nand U3599 (N_3599,N_3428,N_3202);
and U3600 (N_3600,N_3053,N_3273);
nor U3601 (N_3601,N_3419,N_3220);
or U3602 (N_3602,N_3380,N_3270);
nand U3603 (N_3603,N_3252,N_3306);
or U3604 (N_3604,N_3040,N_3011);
nor U3605 (N_3605,N_3114,N_3219);
nand U3606 (N_3606,N_3445,N_3031);
or U3607 (N_3607,N_3235,N_3196);
or U3608 (N_3608,N_3004,N_3404);
nor U3609 (N_3609,N_3442,N_3151);
or U3610 (N_3610,N_3087,N_3304);
nor U3611 (N_3611,N_3356,N_3438);
nor U3612 (N_3612,N_3330,N_3471);
nor U3613 (N_3613,N_3056,N_3488);
nand U3614 (N_3614,N_3174,N_3015);
nand U3615 (N_3615,N_3088,N_3386);
and U3616 (N_3616,N_3137,N_3075);
nand U3617 (N_3617,N_3241,N_3301);
and U3618 (N_3618,N_3098,N_3262);
nand U3619 (N_3619,N_3289,N_3435);
nor U3620 (N_3620,N_3267,N_3455);
xor U3621 (N_3621,N_3450,N_3057);
nand U3622 (N_3622,N_3108,N_3382);
or U3623 (N_3623,N_3394,N_3345);
or U3624 (N_3624,N_3283,N_3163);
nor U3625 (N_3625,N_3400,N_3124);
xor U3626 (N_3626,N_3183,N_3157);
nor U3627 (N_3627,N_3481,N_3129);
and U3628 (N_3628,N_3003,N_3433);
and U3629 (N_3629,N_3067,N_3449);
nand U3630 (N_3630,N_3144,N_3468);
or U3631 (N_3631,N_3396,N_3237);
nor U3632 (N_3632,N_3155,N_3028);
nand U3633 (N_3633,N_3172,N_3194);
nor U3634 (N_3634,N_3233,N_3424);
nor U3635 (N_3635,N_3368,N_3305);
nand U3636 (N_3636,N_3297,N_3242);
and U3637 (N_3637,N_3061,N_3332);
nor U3638 (N_3638,N_3432,N_3170);
nand U3639 (N_3639,N_3265,N_3324);
nor U3640 (N_3640,N_3444,N_3292);
nor U3641 (N_3641,N_3321,N_3315);
nand U3642 (N_3642,N_3228,N_3276);
nand U3643 (N_3643,N_3008,N_3436);
nand U3644 (N_3644,N_3140,N_3310);
and U3645 (N_3645,N_3136,N_3371);
nand U3646 (N_3646,N_3409,N_3027);
and U3647 (N_3647,N_3381,N_3213);
nor U3648 (N_3648,N_3250,N_3277);
xor U3649 (N_3649,N_3311,N_3385);
and U3650 (N_3650,N_3020,N_3372);
or U3651 (N_3651,N_3176,N_3001);
or U3652 (N_3652,N_3344,N_3073);
or U3653 (N_3653,N_3007,N_3209);
nor U3654 (N_3654,N_3439,N_3313);
or U3655 (N_3655,N_3186,N_3068);
and U3656 (N_3656,N_3274,N_3168);
or U3657 (N_3657,N_3418,N_3493);
or U3658 (N_3658,N_3002,N_3205);
or U3659 (N_3659,N_3473,N_3426);
nor U3660 (N_3660,N_3045,N_3249);
or U3661 (N_3661,N_3285,N_3258);
or U3662 (N_3662,N_3290,N_3128);
nor U3663 (N_3663,N_3150,N_3042);
or U3664 (N_3664,N_3352,N_3126);
xor U3665 (N_3665,N_3320,N_3121);
and U3666 (N_3666,N_3175,N_3238);
or U3667 (N_3667,N_3298,N_3117);
nor U3668 (N_3668,N_3302,N_3211);
nand U3669 (N_3669,N_3248,N_3221);
nand U3670 (N_3670,N_3390,N_3360);
nor U3671 (N_3671,N_3012,N_3458);
and U3672 (N_3672,N_3112,N_3154);
nand U3673 (N_3673,N_3331,N_3414);
nand U3674 (N_3674,N_3189,N_3342);
or U3675 (N_3675,N_3016,N_3116);
nand U3676 (N_3676,N_3127,N_3171);
or U3677 (N_3677,N_3412,N_3054);
and U3678 (N_3678,N_3125,N_3457);
nand U3679 (N_3679,N_3019,N_3080);
or U3680 (N_3680,N_3160,N_3224);
and U3681 (N_3681,N_3454,N_3078);
nor U3682 (N_3682,N_3218,N_3165);
nand U3683 (N_3683,N_3314,N_3389);
and U3684 (N_3684,N_3148,N_3065);
or U3685 (N_3685,N_3392,N_3264);
nor U3686 (N_3686,N_3395,N_3091);
nand U3687 (N_3687,N_3119,N_3388);
and U3688 (N_3688,N_3446,N_3033);
nor U3689 (N_3689,N_3466,N_3499);
nor U3690 (N_3690,N_3376,N_3095);
and U3691 (N_3691,N_3401,N_3411);
nor U3692 (N_3692,N_3178,N_3325);
and U3693 (N_3693,N_3122,N_3319);
and U3694 (N_3694,N_3109,N_3210);
or U3695 (N_3695,N_3090,N_3280);
and U3696 (N_3696,N_3353,N_3484);
and U3697 (N_3697,N_3212,N_3048);
nor U3698 (N_3698,N_3257,N_3201);
nand U3699 (N_3699,N_3200,N_3023);
nand U3700 (N_3700,N_3060,N_3156);
and U3701 (N_3701,N_3462,N_3294);
and U3702 (N_3702,N_3483,N_3161);
nor U3703 (N_3703,N_3070,N_3052);
and U3704 (N_3704,N_3204,N_3110);
or U3705 (N_3705,N_3393,N_3480);
nand U3706 (N_3706,N_3246,N_3255);
or U3707 (N_3707,N_3441,N_3131);
and U3708 (N_3708,N_3410,N_3399);
nor U3709 (N_3709,N_3236,N_3440);
and U3710 (N_3710,N_3197,N_3149);
nand U3711 (N_3711,N_3490,N_3269);
and U3712 (N_3712,N_3281,N_3434);
and U3713 (N_3713,N_3355,N_3229);
nor U3714 (N_3714,N_3463,N_3158);
nor U3715 (N_3715,N_3217,N_3077);
nor U3716 (N_3716,N_3199,N_3035);
and U3717 (N_3717,N_3132,N_3275);
nand U3718 (N_3718,N_3317,N_3489);
nand U3719 (N_3719,N_3363,N_3120);
and U3720 (N_3720,N_3254,N_3421);
and U3721 (N_3721,N_3179,N_3085);
or U3722 (N_3722,N_3086,N_3460);
nand U3723 (N_3723,N_3475,N_3318);
and U3724 (N_3724,N_3101,N_3263);
and U3725 (N_3725,N_3230,N_3193);
and U3726 (N_3726,N_3024,N_3074);
nand U3727 (N_3727,N_3308,N_3431);
and U3728 (N_3728,N_3071,N_3417);
nand U3729 (N_3729,N_3415,N_3423);
or U3730 (N_3730,N_3286,N_3307);
nand U3731 (N_3731,N_3123,N_3369);
nor U3732 (N_3732,N_3253,N_3461);
xor U3733 (N_3733,N_3177,N_3147);
nand U3734 (N_3734,N_3367,N_3323);
nor U3735 (N_3735,N_3430,N_3106);
nor U3736 (N_3736,N_3013,N_3187);
nand U3737 (N_3737,N_3387,N_3029);
nor U3738 (N_3738,N_3181,N_3018);
nand U3739 (N_3739,N_3341,N_3402);
nor U3740 (N_3740,N_3184,N_3279);
or U3741 (N_3741,N_3146,N_3334);
xor U3742 (N_3742,N_3470,N_3143);
nor U3743 (N_3743,N_3104,N_3100);
or U3744 (N_3744,N_3322,N_3452);
and U3745 (N_3745,N_3097,N_3456);
or U3746 (N_3746,N_3469,N_3185);
nand U3747 (N_3747,N_3397,N_3287);
nor U3748 (N_3748,N_3055,N_3282);
nor U3749 (N_3749,N_3346,N_3350);
and U3750 (N_3750,N_3455,N_3224);
nor U3751 (N_3751,N_3116,N_3279);
or U3752 (N_3752,N_3340,N_3344);
or U3753 (N_3753,N_3025,N_3186);
nand U3754 (N_3754,N_3149,N_3321);
nand U3755 (N_3755,N_3124,N_3379);
or U3756 (N_3756,N_3447,N_3313);
nor U3757 (N_3757,N_3343,N_3186);
nand U3758 (N_3758,N_3284,N_3324);
nand U3759 (N_3759,N_3255,N_3245);
nor U3760 (N_3760,N_3145,N_3308);
nor U3761 (N_3761,N_3420,N_3419);
and U3762 (N_3762,N_3105,N_3492);
and U3763 (N_3763,N_3367,N_3178);
and U3764 (N_3764,N_3274,N_3049);
nand U3765 (N_3765,N_3451,N_3132);
nor U3766 (N_3766,N_3415,N_3010);
xnor U3767 (N_3767,N_3295,N_3184);
and U3768 (N_3768,N_3033,N_3319);
nor U3769 (N_3769,N_3264,N_3027);
or U3770 (N_3770,N_3086,N_3152);
nor U3771 (N_3771,N_3223,N_3259);
and U3772 (N_3772,N_3128,N_3242);
or U3773 (N_3773,N_3096,N_3214);
or U3774 (N_3774,N_3357,N_3296);
nand U3775 (N_3775,N_3073,N_3441);
nand U3776 (N_3776,N_3429,N_3057);
nand U3777 (N_3777,N_3453,N_3132);
and U3778 (N_3778,N_3478,N_3210);
nand U3779 (N_3779,N_3036,N_3345);
xor U3780 (N_3780,N_3135,N_3174);
nor U3781 (N_3781,N_3268,N_3341);
or U3782 (N_3782,N_3246,N_3459);
and U3783 (N_3783,N_3269,N_3196);
nor U3784 (N_3784,N_3248,N_3080);
nand U3785 (N_3785,N_3492,N_3308);
nor U3786 (N_3786,N_3491,N_3299);
nor U3787 (N_3787,N_3081,N_3252);
nand U3788 (N_3788,N_3047,N_3443);
nor U3789 (N_3789,N_3166,N_3064);
xor U3790 (N_3790,N_3243,N_3475);
and U3791 (N_3791,N_3474,N_3044);
nand U3792 (N_3792,N_3073,N_3010);
or U3793 (N_3793,N_3021,N_3336);
nor U3794 (N_3794,N_3343,N_3463);
nor U3795 (N_3795,N_3498,N_3489);
or U3796 (N_3796,N_3108,N_3063);
nor U3797 (N_3797,N_3271,N_3014);
nor U3798 (N_3798,N_3351,N_3447);
xor U3799 (N_3799,N_3391,N_3434);
nand U3800 (N_3800,N_3443,N_3127);
nor U3801 (N_3801,N_3269,N_3337);
nor U3802 (N_3802,N_3499,N_3104);
nand U3803 (N_3803,N_3328,N_3305);
and U3804 (N_3804,N_3410,N_3457);
and U3805 (N_3805,N_3190,N_3398);
nand U3806 (N_3806,N_3213,N_3032);
nand U3807 (N_3807,N_3296,N_3426);
or U3808 (N_3808,N_3483,N_3295);
or U3809 (N_3809,N_3461,N_3194);
nand U3810 (N_3810,N_3193,N_3173);
and U3811 (N_3811,N_3306,N_3434);
and U3812 (N_3812,N_3232,N_3484);
or U3813 (N_3813,N_3160,N_3388);
or U3814 (N_3814,N_3124,N_3283);
xor U3815 (N_3815,N_3491,N_3227);
nor U3816 (N_3816,N_3198,N_3048);
and U3817 (N_3817,N_3204,N_3157);
or U3818 (N_3818,N_3137,N_3143);
nor U3819 (N_3819,N_3020,N_3292);
and U3820 (N_3820,N_3286,N_3048);
nand U3821 (N_3821,N_3251,N_3024);
nand U3822 (N_3822,N_3222,N_3465);
nand U3823 (N_3823,N_3248,N_3278);
nor U3824 (N_3824,N_3447,N_3241);
nand U3825 (N_3825,N_3487,N_3209);
nand U3826 (N_3826,N_3425,N_3406);
or U3827 (N_3827,N_3195,N_3418);
and U3828 (N_3828,N_3382,N_3254);
nand U3829 (N_3829,N_3392,N_3149);
nor U3830 (N_3830,N_3409,N_3384);
nand U3831 (N_3831,N_3137,N_3081);
nor U3832 (N_3832,N_3416,N_3242);
or U3833 (N_3833,N_3207,N_3477);
and U3834 (N_3834,N_3447,N_3018);
and U3835 (N_3835,N_3321,N_3048);
nand U3836 (N_3836,N_3473,N_3131);
nand U3837 (N_3837,N_3083,N_3051);
or U3838 (N_3838,N_3175,N_3252);
and U3839 (N_3839,N_3253,N_3056);
and U3840 (N_3840,N_3324,N_3158);
or U3841 (N_3841,N_3278,N_3449);
or U3842 (N_3842,N_3298,N_3096);
or U3843 (N_3843,N_3489,N_3269);
or U3844 (N_3844,N_3461,N_3243);
nand U3845 (N_3845,N_3205,N_3057);
xnor U3846 (N_3846,N_3296,N_3018);
and U3847 (N_3847,N_3433,N_3279);
xor U3848 (N_3848,N_3459,N_3252);
and U3849 (N_3849,N_3426,N_3325);
nand U3850 (N_3850,N_3413,N_3262);
nand U3851 (N_3851,N_3295,N_3084);
nand U3852 (N_3852,N_3417,N_3189);
or U3853 (N_3853,N_3431,N_3000);
and U3854 (N_3854,N_3233,N_3473);
xnor U3855 (N_3855,N_3349,N_3048);
nand U3856 (N_3856,N_3424,N_3025);
and U3857 (N_3857,N_3309,N_3311);
nor U3858 (N_3858,N_3342,N_3411);
and U3859 (N_3859,N_3482,N_3353);
nor U3860 (N_3860,N_3465,N_3400);
nor U3861 (N_3861,N_3005,N_3022);
nand U3862 (N_3862,N_3156,N_3378);
nand U3863 (N_3863,N_3191,N_3107);
nor U3864 (N_3864,N_3395,N_3499);
and U3865 (N_3865,N_3202,N_3485);
nand U3866 (N_3866,N_3489,N_3397);
and U3867 (N_3867,N_3300,N_3304);
nor U3868 (N_3868,N_3239,N_3096);
nor U3869 (N_3869,N_3378,N_3335);
and U3870 (N_3870,N_3464,N_3495);
nor U3871 (N_3871,N_3001,N_3151);
or U3872 (N_3872,N_3157,N_3129);
nand U3873 (N_3873,N_3180,N_3047);
or U3874 (N_3874,N_3003,N_3035);
or U3875 (N_3875,N_3045,N_3370);
nand U3876 (N_3876,N_3051,N_3424);
and U3877 (N_3877,N_3206,N_3219);
or U3878 (N_3878,N_3219,N_3167);
and U3879 (N_3879,N_3245,N_3463);
nor U3880 (N_3880,N_3376,N_3429);
nor U3881 (N_3881,N_3350,N_3391);
and U3882 (N_3882,N_3047,N_3030);
nand U3883 (N_3883,N_3293,N_3443);
nor U3884 (N_3884,N_3072,N_3110);
nor U3885 (N_3885,N_3393,N_3105);
and U3886 (N_3886,N_3030,N_3219);
or U3887 (N_3887,N_3429,N_3346);
nor U3888 (N_3888,N_3326,N_3006);
nor U3889 (N_3889,N_3290,N_3480);
nor U3890 (N_3890,N_3082,N_3391);
nand U3891 (N_3891,N_3455,N_3436);
and U3892 (N_3892,N_3135,N_3018);
nand U3893 (N_3893,N_3127,N_3244);
or U3894 (N_3894,N_3305,N_3273);
nor U3895 (N_3895,N_3001,N_3084);
nand U3896 (N_3896,N_3431,N_3088);
and U3897 (N_3897,N_3182,N_3006);
and U3898 (N_3898,N_3482,N_3182);
or U3899 (N_3899,N_3100,N_3497);
nor U3900 (N_3900,N_3079,N_3463);
nor U3901 (N_3901,N_3045,N_3083);
and U3902 (N_3902,N_3259,N_3272);
or U3903 (N_3903,N_3448,N_3072);
nand U3904 (N_3904,N_3100,N_3369);
nor U3905 (N_3905,N_3372,N_3499);
nor U3906 (N_3906,N_3415,N_3472);
xnor U3907 (N_3907,N_3313,N_3209);
nand U3908 (N_3908,N_3140,N_3016);
and U3909 (N_3909,N_3291,N_3116);
and U3910 (N_3910,N_3124,N_3418);
nand U3911 (N_3911,N_3044,N_3101);
or U3912 (N_3912,N_3419,N_3046);
or U3913 (N_3913,N_3276,N_3347);
nand U3914 (N_3914,N_3217,N_3155);
and U3915 (N_3915,N_3425,N_3071);
nor U3916 (N_3916,N_3329,N_3360);
nand U3917 (N_3917,N_3466,N_3389);
or U3918 (N_3918,N_3433,N_3139);
nor U3919 (N_3919,N_3396,N_3319);
and U3920 (N_3920,N_3449,N_3012);
nor U3921 (N_3921,N_3193,N_3298);
and U3922 (N_3922,N_3353,N_3135);
and U3923 (N_3923,N_3033,N_3368);
or U3924 (N_3924,N_3444,N_3216);
and U3925 (N_3925,N_3480,N_3241);
or U3926 (N_3926,N_3295,N_3102);
nor U3927 (N_3927,N_3178,N_3436);
nand U3928 (N_3928,N_3358,N_3221);
nand U3929 (N_3929,N_3337,N_3413);
nor U3930 (N_3930,N_3081,N_3185);
nand U3931 (N_3931,N_3415,N_3198);
or U3932 (N_3932,N_3018,N_3331);
nand U3933 (N_3933,N_3216,N_3380);
nand U3934 (N_3934,N_3184,N_3262);
nor U3935 (N_3935,N_3297,N_3326);
or U3936 (N_3936,N_3278,N_3000);
nor U3937 (N_3937,N_3129,N_3423);
nor U3938 (N_3938,N_3352,N_3328);
or U3939 (N_3939,N_3409,N_3198);
or U3940 (N_3940,N_3293,N_3346);
or U3941 (N_3941,N_3095,N_3446);
nand U3942 (N_3942,N_3005,N_3357);
or U3943 (N_3943,N_3375,N_3495);
and U3944 (N_3944,N_3483,N_3187);
nand U3945 (N_3945,N_3326,N_3332);
or U3946 (N_3946,N_3070,N_3229);
nand U3947 (N_3947,N_3398,N_3472);
nand U3948 (N_3948,N_3447,N_3077);
and U3949 (N_3949,N_3389,N_3483);
or U3950 (N_3950,N_3171,N_3499);
nor U3951 (N_3951,N_3198,N_3078);
and U3952 (N_3952,N_3309,N_3322);
or U3953 (N_3953,N_3469,N_3334);
and U3954 (N_3954,N_3001,N_3431);
nor U3955 (N_3955,N_3147,N_3216);
nor U3956 (N_3956,N_3489,N_3008);
or U3957 (N_3957,N_3417,N_3376);
nor U3958 (N_3958,N_3489,N_3038);
or U3959 (N_3959,N_3463,N_3280);
or U3960 (N_3960,N_3209,N_3307);
and U3961 (N_3961,N_3118,N_3003);
nor U3962 (N_3962,N_3192,N_3453);
nand U3963 (N_3963,N_3333,N_3334);
and U3964 (N_3964,N_3404,N_3251);
and U3965 (N_3965,N_3490,N_3218);
nand U3966 (N_3966,N_3273,N_3031);
nand U3967 (N_3967,N_3383,N_3211);
or U3968 (N_3968,N_3429,N_3328);
nor U3969 (N_3969,N_3109,N_3202);
nand U3970 (N_3970,N_3330,N_3464);
nor U3971 (N_3971,N_3368,N_3379);
nor U3972 (N_3972,N_3281,N_3437);
nand U3973 (N_3973,N_3155,N_3479);
nor U3974 (N_3974,N_3053,N_3045);
and U3975 (N_3975,N_3099,N_3487);
nor U3976 (N_3976,N_3494,N_3375);
nor U3977 (N_3977,N_3005,N_3105);
and U3978 (N_3978,N_3359,N_3361);
nand U3979 (N_3979,N_3066,N_3040);
nor U3980 (N_3980,N_3172,N_3088);
and U3981 (N_3981,N_3205,N_3160);
or U3982 (N_3982,N_3148,N_3293);
or U3983 (N_3983,N_3307,N_3244);
and U3984 (N_3984,N_3495,N_3439);
and U3985 (N_3985,N_3277,N_3425);
nor U3986 (N_3986,N_3273,N_3167);
nand U3987 (N_3987,N_3032,N_3308);
and U3988 (N_3988,N_3474,N_3237);
nor U3989 (N_3989,N_3357,N_3069);
nor U3990 (N_3990,N_3074,N_3310);
xor U3991 (N_3991,N_3060,N_3436);
nand U3992 (N_3992,N_3339,N_3399);
and U3993 (N_3993,N_3106,N_3027);
nor U3994 (N_3994,N_3028,N_3476);
and U3995 (N_3995,N_3427,N_3017);
nand U3996 (N_3996,N_3196,N_3142);
or U3997 (N_3997,N_3146,N_3276);
and U3998 (N_3998,N_3441,N_3252);
and U3999 (N_3999,N_3083,N_3035);
nand U4000 (N_4000,N_3723,N_3990);
nor U4001 (N_4001,N_3794,N_3917);
xnor U4002 (N_4002,N_3666,N_3968);
or U4003 (N_4003,N_3928,N_3791);
or U4004 (N_4004,N_3809,N_3697);
nand U4005 (N_4005,N_3537,N_3500);
xor U4006 (N_4006,N_3911,N_3650);
xnor U4007 (N_4007,N_3895,N_3737);
or U4008 (N_4008,N_3565,N_3715);
or U4009 (N_4009,N_3852,N_3975);
xnor U4010 (N_4010,N_3614,N_3627);
or U4011 (N_4011,N_3628,N_3644);
xnor U4012 (N_4012,N_3717,N_3600);
and U4013 (N_4013,N_3949,N_3766);
or U4014 (N_4014,N_3958,N_3813);
nor U4015 (N_4015,N_3573,N_3687);
or U4016 (N_4016,N_3743,N_3775);
or U4017 (N_4017,N_3703,N_3673);
nand U4018 (N_4018,N_3563,N_3993);
or U4019 (N_4019,N_3726,N_3626);
nand U4020 (N_4020,N_3521,N_3718);
nor U4021 (N_4021,N_3839,N_3690);
or U4022 (N_4022,N_3732,N_3876);
nor U4023 (N_4023,N_3858,N_3857);
nor U4024 (N_4024,N_3591,N_3517);
nor U4025 (N_4025,N_3724,N_3598);
nor U4026 (N_4026,N_3580,N_3662);
nand U4027 (N_4027,N_3643,N_3587);
nand U4028 (N_4028,N_3962,N_3758);
and U4029 (N_4029,N_3701,N_3884);
nand U4030 (N_4030,N_3522,N_3868);
or U4031 (N_4031,N_3647,N_3889);
nand U4032 (N_4032,N_3906,N_3608);
and U4033 (N_4033,N_3745,N_3923);
and U4034 (N_4034,N_3931,N_3530);
nor U4035 (N_4035,N_3552,N_3657);
or U4036 (N_4036,N_3756,N_3865);
nor U4037 (N_4037,N_3551,N_3998);
or U4038 (N_4038,N_3991,N_3538);
nor U4039 (N_4039,N_3654,N_3955);
nor U4040 (N_4040,N_3784,N_3945);
or U4041 (N_4041,N_3524,N_3547);
xor U4042 (N_4042,N_3900,N_3891);
nor U4043 (N_4043,N_3705,N_3610);
nand U4044 (N_4044,N_3944,N_3790);
and U4045 (N_4045,N_3820,N_3841);
nor U4046 (N_4046,N_3992,N_3795);
or U4047 (N_4047,N_3965,N_3748);
and U4048 (N_4048,N_3523,N_3698);
and U4049 (N_4049,N_3943,N_3631);
nor U4050 (N_4050,N_3902,N_3555);
nor U4051 (N_4051,N_3772,N_3974);
nor U4052 (N_4052,N_3875,N_3957);
nand U4053 (N_4053,N_3898,N_3616);
xor U4054 (N_4054,N_3503,N_3568);
or U4055 (N_4055,N_3533,N_3874);
or U4056 (N_4056,N_3822,N_3576);
or U4057 (N_4057,N_3562,N_3802);
or U4058 (N_4058,N_3678,N_3672);
or U4059 (N_4059,N_3680,N_3633);
and U4060 (N_4060,N_3693,N_3824);
or U4061 (N_4061,N_3663,N_3785);
and U4062 (N_4062,N_3682,N_3935);
nand U4063 (N_4063,N_3601,N_3982);
and U4064 (N_4064,N_3954,N_3632);
nor U4065 (N_4065,N_3719,N_3752);
or U4066 (N_4066,N_3544,N_3916);
nor U4067 (N_4067,N_3527,N_3816);
nor U4068 (N_4068,N_3854,N_3656);
nor U4069 (N_4069,N_3599,N_3606);
nor U4070 (N_4070,N_3769,N_3787);
nor U4071 (N_4071,N_3881,N_3782);
nand U4072 (N_4072,N_3634,N_3560);
and U4073 (N_4073,N_3519,N_3995);
and U4074 (N_4074,N_3776,N_3780);
nor U4075 (N_4075,N_3762,N_3940);
nand U4076 (N_4076,N_3984,N_3799);
nand U4077 (N_4077,N_3988,N_3863);
nand U4078 (N_4078,N_3735,N_3566);
and U4079 (N_4079,N_3542,N_3751);
and U4080 (N_4080,N_3921,N_3938);
nand U4081 (N_4081,N_3897,N_3676);
nor U4082 (N_4082,N_3515,N_3578);
or U4083 (N_4083,N_3828,N_3589);
or U4084 (N_4084,N_3936,N_3624);
and U4085 (N_4085,N_3727,N_3856);
and U4086 (N_4086,N_3511,N_3877);
or U4087 (N_4087,N_3952,N_3689);
or U4088 (N_4088,N_3843,N_3840);
or U4089 (N_4089,N_3826,N_3759);
nand U4090 (N_4090,N_3878,N_3959);
nand U4091 (N_4091,N_3996,N_3509);
and U4092 (N_4092,N_3770,N_3512);
and U4093 (N_4093,N_3557,N_3640);
or U4094 (N_4094,N_3947,N_3831);
nor U4095 (N_4095,N_3683,N_3611);
nand U4096 (N_4096,N_3778,N_3948);
and U4097 (N_4097,N_3811,N_3963);
and U4098 (N_4098,N_3603,N_3651);
nand U4099 (N_4099,N_3773,N_3939);
nand U4100 (N_4100,N_3604,N_3629);
nand U4101 (N_4101,N_3887,N_3716);
and U4102 (N_4102,N_3847,N_3883);
nand U4103 (N_4103,N_3504,N_3708);
nand U4104 (N_4104,N_3907,N_3637);
nand U4105 (N_4105,N_3607,N_3746);
nand U4106 (N_4106,N_3692,N_3969);
and U4107 (N_4107,N_3671,N_3583);
and U4108 (N_4108,N_3951,N_3910);
nor U4109 (N_4109,N_3804,N_3966);
or U4110 (N_4110,N_3920,N_3691);
nor U4111 (N_4111,N_3722,N_3832);
nand U4112 (N_4112,N_3837,N_3882);
nand U4113 (N_4113,N_3567,N_3674);
or U4114 (N_4114,N_3501,N_3505);
or U4115 (N_4115,N_3873,N_3605);
and U4116 (N_4116,N_3888,N_3588);
and U4117 (N_4117,N_3893,N_3846);
and U4118 (N_4118,N_3710,N_3908);
and U4119 (N_4119,N_3648,N_3972);
nor U4120 (N_4120,N_3658,N_3688);
and U4121 (N_4121,N_3646,N_3535);
and U4122 (N_4122,N_3638,N_3914);
nand U4123 (N_4123,N_3767,N_3903);
and U4124 (N_4124,N_3994,N_3808);
nor U4125 (N_4125,N_3618,N_3559);
and U4126 (N_4126,N_3801,N_3595);
and U4127 (N_4127,N_3602,N_3684);
nor U4128 (N_4128,N_3792,N_3980);
nor U4129 (N_4129,N_3899,N_3681);
and U4130 (N_4130,N_3890,N_3845);
xnor U4131 (N_4131,N_3532,N_3866);
and U4132 (N_4132,N_3669,N_3570);
or U4133 (N_4133,N_3927,N_3979);
nand U4134 (N_4134,N_3549,N_3805);
nor U4135 (N_4135,N_3871,N_3575);
or U4136 (N_4136,N_3649,N_3668);
and U4137 (N_4137,N_3971,N_3729);
nor U4138 (N_4138,N_3976,N_3981);
nor U4139 (N_4139,N_3529,N_3685);
and U4140 (N_4140,N_3937,N_3803);
nand U4141 (N_4141,N_3825,N_3918);
or U4142 (N_4142,N_3569,N_3777);
nand U4143 (N_4143,N_3926,N_3812);
nor U4144 (N_4144,N_3997,N_3941);
nor U4145 (N_4145,N_3985,N_3741);
nand U4146 (N_4146,N_3836,N_3571);
or U4147 (N_4147,N_3919,N_3929);
nand U4148 (N_4148,N_3860,N_3516);
nand U4149 (N_4149,N_3950,N_3556);
and U4150 (N_4150,N_3564,N_3531);
and U4151 (N_4151,N_3536,N_3879);
and U4152 (N_4152,N_3545,N_3933);
and U4153 (N_4153,N_3786,N_3763);
or U4154 (N_4154,N_3789,N_3946);
nor U4155 (N_4155,N_3783,N_3848);
and U4156 (N_4156,N_3768,N_3528);
nand U4157 (N_4157,N_3834,N_3582);
nand U4158 (N_4158,N_3645,N_3740);
nand U4159 (N_4159,N_3728,N_3593);
xnor U4160 (N_4160,N_3967,N_3700);
nor U4161 (N_4161,N_3525,N_3842);
or U4162 (N_4162,N_3986,N_3818);
and U4163 (N_4163,N_3987,N_3541);
nand U4164 (N_4164,N_3696,N_3749);
nand U4165 (N_4165,N_3757,N_3619);
or U4166 (N_4166,N_3546,N_3750);
nor U4167 (N_4167,N_3586,N_3709);
xnor U4168 (N_4168,N_3543,N_3655);
nor U4169 (N_4169,N_3925,N_3507);
or U4170 (N_4170,N_3844,N_3869);
or U4171 (N_4171,N_3999,N_3686);
and U4172 (N_4172,N_3742,N_3872);
nor U4173 (N_4173,N_3807,N_3679);
nand U4174 (N_4174,N_3815,N_3510);
and U4175 (N_4175,N_3913,N_3721);
and U4176 (N_4176,N_3880,N_3514);
nor U4177 (N_4177,N_3659,N_3983);
and U4178 (N_4178,N_3930,N_3725);
or U4179 (N_4179,N_3922,N_3901);
nor U4180 (N_4180,N_3553,N_3753);
and U4181 (N_4181,N_3830,N_3706);
nand U4182 (N_4182,N_3506,N_3579);
nor U4183 (N_4183,N_3660,N_3594);
or U4184 (N_4184,N_3934,N_3764);
nor U4185 (N_4185,N_3704,N_3635);
nor U4186 (N_4186,N_3886,N_3885);
and U4187 (N_4187,N_3652,N_3771);
and U4188 (N_4188,N_3639,N_3636);
and U4189 (N_4189,N_3924,N_3964);
or U4190 (N_4190,N_3806,N_3932);
or U4191 (N_4191,N_3733,N_3829);
or U4192 (N_4192,N_3850,N_3796);
nand U4193 (N_4193,N_3621,N_3833);
nand U4194 (N_4194,N_3960,N_3730);
or U4195 (N_4195,N_3518,N_3581);
nand U4196 (N_4196,N_3779,N_3675);
and U4197 (N_4197,N_3862,N_3953);
or U4198 (N_4198,N_3909,N_3814);
nand U4199 (N_4199,N_3592,N_3774);
nor U4200 (N_4200,N_3713,N_3653);
nand U4201 (N_4201,N_3574,N_3912);
nand U4202 (N_4202,N_3609,N_3590);
nor U4203 (N_4203,N_3699,N_3670);
nand U4204 (N_4204,N_3738,N_3539);
nor U4205 (N_4205,N_3861,N_3597);
nand U4206 (N_4206,N_3620,N_3534);
and U4207 (N_4207,N_3502,N_3838);
nor U4208 (N_4208,N_3548,N_3550);
or U4209 (N_4209,N_3513,N_3904);
nor U4210 (N_4210,N_3744,N_3665);
or U4211 (N_4211,N_3747,N_3625);
nor U4212 (N_4212,N_3970,N_3894);
or U4213 (N_4213,N_3859,N_3855);
nand U4214 (N_4214,N_3765,N_3661);
nand U4215 (N_4215,N_3720,N_3642);
nand U4216 (N_4216,N_3617,N_3819);
nor U4217 (N_4217,N_3827,N_3711);
or U4218 (N_4218,N_3942,N_3558);
nor U4219 (N_4219,N_3540,N_3892);
or U4220 (N_4220,N_3797,N_3781);
nand U4221 (N_4221,N_3615,N_3630);
nand U4222 (N_4222,N_3977,N_3961);
xor U4223 (N_4223,N_3712,N_3835);
and U4224 (N_4224,N_3508,N_3612);
xnor U4225 (N_4225,N_3956,N_3915);
nor U4226 (N_4226,N_3520,N_3755);
nand U4227 (N_4227,N_3973,N_3739);
nand U4228 (N_4228,N_3577,N_3526);
nand U4229 (N_4229,N_3851,N_3702);
nand U4230 (N_4230,N_3905,N_3623);
nand U4231 (N_4231,N_3867,N_3798);
or U4232 (N_4232,N_3572,N_3793);
nand U4233 (N_4233,N_3989,N_3596);
and U4234 (N_4234,N_3561,N_3695);
nand U4235 (N_4235,N_3788,N_3760);
or U4236 (N_4236,N_3734,N_3584);
or U4237 (N_4237,N_3667,N_3853);
and U4238 (N_4238,N_3736,N_3896);
nand U4239 (N_4239,N_3677,N_3641);
and U4240 (N_4240,N_3707,N_3694);
nand U4241 (N_4241,N_3622,N_3870);
nor U4242 (N_4242,N_3761,N_3864);
xor U4243 (N_4243,N_3978,N_3731);
nor U4244 (N_4244,N_3800,N_3849);
and U4245 (N_4245,N_3714,N_3613);
nand U4246 (N_4246,N_3821,N_3810);
nand U4247 (N_4247,N_3664,N_3754);
nor U4248 (N_4248,N_3817,N_3554);
nor U4249 (N_4249,N_3823,N_3585);
and U4250 (N_4250,N_3567,N_3645);
or U4251 (N_4251,N_3710,N_3528);
xnor U4252 (N_4252,N_3998,N_3661);
nand U4253 (N_4253,N_3869,N_3896);
nor U4254 (N_4254,N_3893,N_3588);
nand U4255 (N_4255,N_3662,N_3948);
or U4256 (N_4256,N_3718,N_3838);
and U4257 (N_4257,N_3828,N_3719);
or U4258 (N_4258,N_3731,N_3544);
or U4259 (N_4259,N_3703,N_3806);
nor U4260 (N_4260,N_3647,N_3734);
or U4261 (N_4261,N_3626,N_3791);
nand U4262 (N_4262,N_3873,N_3522);
nand U4263 (N_4263,N_3888,N_3741);
nor U4264 (N_4264,N_3924,N_3898);
nand U4265 (N_4265,N_3556,N_3580);
nor U4266 (N_4266,N_3775,N_3938);
or U4267 (N_4267,N_3945,N_3793);
nand U4268 (N_4268,N_3605,N_3792);
and U4269 (N_4269,N_3837,N_3775);
or U4270 (N_4270,N_3863,N_3903);
or U4271 (N_4271,N_3798,N_3942);
nand U4272 (N_4272,N_3847,N_3699);
nand U4273 (N_4273,N_3597,N_3752);
nand U4274 (N_4274,N_3932,N_3922);
nor U4275 (N_4275,N_3897,N_3668);
and U4276 (N_4276,N_3680,N_3921);
nor U4277 (N_4277,N_3510,N_3659);
nor U4278 (N_4278,N_3668,N_3701);
nor U4279 (N_4279,N_3876,N_3668);
nand U4280 (N_4280,N_3811,N_3564);
and U4281 (N_4281,N_3694,N_3763);
or U4282 (N_4282,N_3754,N_3770);
nor U4283 (N_4283,N_3978,N_3730);
or U4284 (N_4284,N_3991,N_3836);
and U4285 (N_4285,N_3841,N_3502);
or U4286 (N_4286,N_3702,N_3500);
nand U4287 (N_4287,N_3949,N_3951);
or U4288 (N_4288,N_3879,N_3706);
or U4289 (N_4289,N_3924,N_3534);
or U4290 (N_4290,N_3916,N_3501);
or U4291 (N_4291,N_3510,N_3786);
nand U4292 (N_4292,N_3837,N_3718);
xnor U4293 (N_4293,N_3858,N_3850);
or U4294 (N_4294,N_3527,N_3746);
nand U4295 (N_4295,N_3958,N_3747);
or U4296 (N_4296,N_3693,N_3780);
or U4297 (N_4297,N_3806,N_3710);
or U4298 (N_4298,N_3790,N_3814);
and U4299 (N_4299,N_3708,N_3744);
nor U4300 (N_4300,N_3825,N_3824);
and U4301 (N_4301,N_3702,N_3956);
nand U4302 (N_4302,N_3608,N_3541);
nor U4303 (N_4303,N_3579,N_3791);
and U4304 (N_4304,N_3862,N_3693);
nand U4305 (N_4305,N_3749,N_3556);
nor U4306 (N_4306,N_3713,N_3838);
or U4307 (N_4307,N_3964,N_3865);
nand U4308 (N_4308,N_3877,N_3827);
nand U4309 (N_4309,N_3675,N_3746);
or U4310 (N_4310,N_3863,N_3860);
or U4311 (N_4311,N_3928,N_3807);
xor U4312 (N_4312,N_3624,N_3699);
nor U4313 (N_4313,N_3517,N_3859);
nand U4314 (N_4314,N_3636,N_3510);
nor U4315 (N_4315,N_3903,N_3748);
nand U4316 (N_4316,N_3532,N_3741);
nor U4317 (N_4317,N_3934,N_3696);
nand U4318 (N_4318,N_3757,N_3809);
nor U4319 (N_4319,N_3805,N_3956);
or U4320 (N_4320,N_3779,N_3556);
nand U4321 (N_4321,N_3925,N_3550);
and U4322 (N_4322,N_3711,N_3653);
nor U4323 (N_4323,N_3910,N_3774);
and U4324 (N_4324,N_3581,N_3531);
nand U4325 (N_4325,N_3636,N_3734);
nor U4326 (N_4326,N_3523,N_3669);
or U4327 (N_4327,N_3938,N_3846);
nor U4328 (N_4328,N_3700,N_3723);
nand U4329 (N_4329,N_3637,N_3665);
nor U4330 (N_4330,N_3846,N_3664);
or U4331 (N_4331,N_3711,N_3684);
and U4332 (N_4332,N_3525,N_3515);
and U4333 (N_4333,N_3714,N_3805);
nor U4334 (N_4334,N_3703,N_3894);
or U4335 (N_4335,N_3779,N_3897);
and U4336 (N_4336,N_3535,N_3780);
nand U4337 (N_4337,N_3695,N_3554);
and U4338 (N_4338,N_3625,N_3610);
nand U4339 (N_4339,N_3592,N_3525);
nor U4340 (N_4340,N_3817,N_3822);
and U4341 (N_4341,N_3635,N_3802);
and U4342 (N_4342,N_3519,N_3739);
and U4343 (N_4343,N_3997,N_3539);
nor U4344 (N_4344,N_3674,N_3985);
or U4345 (N_4345,N_3975,N_3835);
and U4346 (N_4346,N_3943,N_3608);
nand U4347 (N_4347,N_3767,N_3935);
xor U4348 (N_4348,N_3648,N_3652);
and U4349 (N_4349,N_3859,N_3953);
nand U4350 (N_4350,N_3668,N_3690);
or U4351 (N_4351,N_3630,N_3792);
and U4352 (N_4352,N_3712,N_3764);
nor U4353 (N_4353,N_3871,N_3932);
nand U4354 (N_4354,N_3632,N_3717);
nor U4355 (N_4355,N_3590,N_3884);
nand U4356 (N_4356,N_3981,N_3745);
or U4357 (N_4357,N_3522,N_3689);
or U4358 (N_4358,N_3846,N_3827);
nor U4359 (N_4359,N_3941,N_3751);
nand U4360 (N_4360,N_3767,N_3843);
nor U4361 (N_4361,N_3847,N_3988);
or U4362 (N_4362,N_3760,N_3875);
nand U4363 (N_4363,N_3572,N_3556);
or U4364 (N_4364,N_3715,N_3975);
nand U4365 (N_4365,N_3662,N_3934);
and U4366 (N_4366,N_3939,N_3682);
nor U4367 (N_4367,N_3501,N_3511);
nor U4368 (N_4368,N_3973,N_3868);
or U4369 (N_4369,N_3683,N_3866);
nor U4370 (N_4370,N_3644,N_3580);
or U4371 (N_4371,N_3529,N_3932);
and U4372 (N_4372,N_3843,N_3982);
and U4373 (N_4373,N_3745,N_3600);
or U4374 (N_4374,N_3626,N_3766);
and U4375 (N_4375,N_3947,N_3596);
nand U4376 (N_4376,N_3899,N_3504);
nand U4377 (N_4377,N_3561,N_3605);
or U4378 (N_4378,N_3635,N_3785);
nand U4379 (N_4379,N_3957,N_3853);
nand U4380 (N_4380,N_3847,N_3806);
nor U4381 (N_4381,N_3539,N_3943);
and U4382 (N_4382,N_3505,N_3886);
or U4383 (N_4383,N_3666,N_3776);
nor U4384 (N_4384,N_3891,N_3844);
nand U4385 (N_4385,N_3579,N_3600);
nand U4386 (N_4386,N_3671,N_3534);
nand U4387 (N_4387,N_3815,N_3640);
nor U4388 (N_4388,N_3731,N_3983);
nor U4389 (N_4389,N_3791,N_3535);
and U4390 (N_4390,N_3640,N_3694);
nor U4391 (N_4391,N_3931,N_3704);
xor U4392 (N_4392,N_3517,N_3764);
nor U4393 (N_4393,N_3538,N_3783);
and U4394 (N_4394,N_3685,N_3643);
nand U4395 (N_4395,N_3845,N_3818);
or U4396 (N_4396,N_3518,N_3795);
and U4397 (N_4397,N_3540,N_3919);
nand U4398 (N_4398,N_3725,N_3816);
and U4399 (N_4399,N_3766,N_3710);
nand U4400 (N_4400,N_3514,N_3673);
or U4401 (N_4401,N_3999,N_3850);
and U4402 (N_4402,N_3575,N_3860);
or U4403 (N_4403,N_3991,N_3618);
or U4404 (N_4404,N_3837,N_3729);
and U4405 (N_4405,N_3983,N_3660);
and U4406 (N_4406,N_3695,N_3915);
and U4407 (N_4407,N_3898,N_3793);
and U4408 (N_4408,N_3695,N_3553);
nand U4409 (N_4409,N_3996,N_3714);
and U4410 (N_4410,N_3666,N_3813);
or U4411 (N_4411,N_3782,N_3522);
nor U4412 (N_4412,N_3581,N_3932);
and U4413 (N_4413,N_3833,N_3594);
or U4414 (N_4414,N_3774,N_3969);
nor U4415 (N_4415,N_3782,N_3601);
nor U4416 (N_4416,N_3540,N_3605);
and U4417 (N_4417,N_3503,N_3701);
nor U4418 (N_4418,N_3646,N_3878);
or U4419 (N_4419,N_3819,N_3697);
or U4420 (N_4420,N_3542,N_3814);
and U4421 (N_4421,N_3799,N_3968);
nand U4422 (N_4422,N_3810,N_3650);
nor U4423 (N_4423,N_3808,N_3874);
nand U4424 (N_4424,N_3981,N_3669);
or U4425 (N_4425,N_3980,N_3890);
or U4426 (N_4426,N_3547,N_3532);
or U4427 (N_4427,N_3510,N_3696);
and U4428 (N_4428,N_3642,N_3874);
nand U4429 (N_4429,N_3521,N_3885);
or U4430 (N_4430,N_3594,N_3930);
nand U4431 (N_4431,N_3715,N_3759);
nand U4432 (N_4432,N_3630,N_3881);
nor U4433 (N_4433,N_3767,N_3602);
xnor U4434 (N_4434,N_3520,N_3854);
nand U4435 (N_4435,N_3886,N_3534);
nand U4436 (N_4436,N_3756,N_3810);
or U4437 (N_4437,N_3891,N_3751);
or U4438 (N_4438,N_3829,N_3822);
or U4439 (N_4439,N_3749,N_3821);
nor U4440 (N_4440,N_3646,N_3520);
nor U4441 (N_4441,N_3866,N_3654);
xnor U4442 (N_4442,N_3655,N_3701);
and U4443 (N_4443,N_3679,N_3952);
or U4444 (N_4444,N_3724,N_3690);
or U4445 (N_4445,N_3577,N_3949);
and U4446 (N_4446,N_3732,N_3775);
and U4447 (N_4447,N_3568,N_3611);
nand U4448 (N_4448,N_3967,N_3897);
and U4449 (N_4449,N_3548,N_3916);
or U4450 (N_4450,N_3966,N_3838);
nand U4451 (N_4451,N_3720,N_3975);
and U4452 (N_4452,N_3754,N_3760);
and U4453 (N_4453,N_3890,N_3630);
nand U4454 (N_4454,N_3683,N_3501);
nand U4455 (N_4455,N_3922,N_3575);
and U4456 (N_4456,N_3959,N_3619);
nand U4457 (N_4457,N_3936,N_3932);
nor U4458 (N_4458,N_3900,N_3579);
and U4459 (N_4459,N_3937,N_3541);
and U4460 (N_4460,N_3519,N_3850);
nor U4461 (N_4461,N_3792,N_3836);
or U4462 (N_4462,N_3565,N_3769);
nor U4463 (N_4463,N_3995,N_3855);
nor U4464 (N_4464,N_3938,N_3551);
and U4465 (N_4465,N_3572,N_3979);
nand U4466 (N_4466,N_3515,N_3902);
nand U4467 (N_4467,N_3567,N_3536);
nor U4468 (N_4468,N_3764,N_3715);
or U4469 (N_4469,N_3640,N_3700);
nor U4470 (N_4470,N_3737,N_3713);
and U4471 (N_4471,N_3912,N_3665);
and U4472 (N_4472,N_3669,N_3531);
and U4473 (N_4473,N_3736,N_3988);
nor U4474 (N_4474,N_3825,N_3624);
nand U4475 (N_4475,N_3921,N_3619);
xor U4476 (N_4476,N_3551,N_3514);
nor U4477 (N_4477,N_3974,N_3950);
and U4478 (N_4478,N_3655,N_3878);
nor U4479 (N_4479,N_3646,N_3868);
and U4480 (N_4480,N_3549,N_3871);
nor U4481 (N_4481,N_3916,N_3863);
nor U4482 (N_4482,N_3723,N_3760);
nor U4483 (N_4483,N_3584,N_3783);
or U4484 (N_4484,N_3968,N_3938);
and U4485 (N_4485,N_3605,N_3646);
nor U4486 (N_4486,N_3545,N_3681);
or U4487 (N_4487,N_3790,N_3734);
nand U4488 (N_4488,N_3542,N_3738);
nor U4489 (N_4489,N_3579,N_3882);
or U4490 (N_4490,N_3579,N_3828);
or U4491 (N_4491,N_3517,N_3830);
or U4492 (N_4492,N_3897,N_3742);
and U4493 (N_4493,N_3575,N_3643);
nand U4494 (N_4494,N_3973,N_3907);
and U4495 (N_4495,N_3799,N_3879);
or U4496 (N_4496,N_3728,N_3782);
nor U4497 (N_4497,N_3616,N_3768);
nor U4498 (N_4498,N_3786,N_3757);
nor U4499 (N_4499,N_3885,N_3684);
nand U4500 (N_4500,N_4128,N_4235);
xnor U4501 (N_4501,N_4246,N_4448);
or U4502 (N_4502,N_4006,N_4017);
nor U4503 (N_4503,N_4323,N_4094);
nand U4504 (N_4504,N_4170,N_4333);
nand U4505 (N_4505,N_4185,N_4048);
nand U4506 (N_4506,N_4462,N_4434);
and U4507 (N_4507,N_4282,N_4463);
and U4508 (N_4508,N_4020,N_4401);
nand U4509 (N_4509,N_4150,N_4126);
or U4510 (N_4510,N_4445,N_4438);
and U4511 (N_4511,N_4091,N_4305);
nand U4512 (N_4512,N_4073,N_4441);
or U4513 (N_4513,N_4104,N_4076);
nor U4514 (N_4514,N_4168,N_4457);
and U4515 (N_4515,N_4470,N_4349);
nand U4516 (N_4516,N_4249,N_4204);
nor U4517 (N_4517,N_4269,N_4310);
nor U4518 (N_4518,N_4248,N_4217);
nand U4519 (N_4519,N_4133,N_4139);
or U4520 (N_4520,N_4381,N_4487);
nor U4521 (N_4521,N_4315,N_4374);
or U4522 (N_4522,N_4491,N_4407);
or U4523 (N_4523,N_4067,N_4052);
and U4524 (N_4524,N_4149,N_4499);
and U4525 (N_4525,N_4300,N_4069);
nor U4526 (N_4526,N_4353,N_4112);
nor U4527 (N_4527,N_4225,N_4182);
nand U4528 (N_4528,N_4007,N_4041);
or U4529 (N_4529,N_4483,N_4125);
nor U4530 (N_4530,N_4306,N_4253);
nor U4531 (N_4531,N_4346,N_4026);
and U4532 (N_4532,N_4180,N_4453);
nand U4533 (N_4533,N_4016,N_4392);
and U4534 (N_4534,N_4454,N_4271);
nor U4535 (N_4535,N_4070,N_4080);
and U4536 (N_4536,N_4172,N_4406);
nor U4537 (N_4537,N_4378,N_4409);
nand U4538 (N_4538,N_4242,N_4433);
and U4539 (N_4539,N_4130,N_4356);
or U4540 (N_4540,N_4321,N_4264);
nand U4541 (N_4541,N_4232,N_4102);
and U4542 (N_4542,N_4311,N_4276);
or U4543 (N_4543,N_4473,N_4288);
xnor U4544 (N_4544,N_4215,N_4456);
or U4545 (N_4545,N_4372,N_4044);
and U4546 (N_4546,N_4286,N_4089);
nor U4547 (N_4547,N_4440,N_4029);
and U4548 (N_4548,N_4093,N_4335);
and U4549 (N_4549,N_4416,N_4493);
nand U4550 (N_4550,N_4195,N_4365);
or U4551 (N_4551,N_4354,N_4152);
nor U4552 (N_4552,N_4121,N_4027);
nand U4553 (N_4553,N_4414,N_4480);
or U4554 (N_4554,N_4135,N_4368);
nand U4555 (N_4555,N_4380,N_4050);
and U4556 (N_4556,N_4083,N_4108);
or U4557 (N_4557,N_4032,N_4210);
nand U4558 (N_4558,N_4071,N_4422);
or U4559 (N_4559,N_4161,N_4064);
and U4560 (N_4560,N_4051,N_4008);
nor U4561 (N_4561,N_4224,N_4239);
nor U4562 (N_4562,N_4371,N_4498);
nor U4563 (N_4563,N_4436,N_4338);
nor U4564 (N_4564,N_4400,N_4452);
and U4565 (N_4565,N_4489,N_4360);
and U4566 (N_4566,N_4347,N_4166);
and U4567 (N_4567,N_4298,N_4199);
or U4568 (N_4568,N_4013,N_4458);
nand U4569 (N_4569,N_4496,N_4223);
and U4570 (N_4570,N_4009,N_4326);
nand U4571 (N_4571,N_4475,N_4163);
nor U4572 (N_4572,N_4355,N_4218);
or U4573 (N_4573,N_4294,N_4318);
xor U4574 (N_4574,N_4230,N_4134);
and U4575 (N_4575,N_4228,N_4226);
nand U4576 (N_4576,N_4053,N_4086);
or U4577 (N_4577,N_4307,N_4184);
or U4578 (N_4578,N_4181,N_4390);
and U4579 (N_4579,N_4319,N_4472);
or U4580 (N_4580,N_4369,N_4330);
and U4581 (N_4581,N_4328,N_4268);
nor U4582 (N_4582,N_4046,N_4238);
nor U4583 (N_4583,N_4256,N_4297);
nand U4584 (N_4584,N_4469,N_4003);
nor U4585 (N_4585,N_4122,N_4019);
and U4586 (N_4586,N_4274,N_4272);
and U4587 (N_4587,N_4279,N_4159);
and U4588 (N_4588,N_4012,N_4043);
and U4589 (N_4589,N_4100,N_4148);
nor U4590 (N_4590,N_4485,N_4474);
nor U4591 (N_4591,N_4343,N_4258);
nor U4592 (N_4592,N_4363,N_4156);
nor U4593 (N_4593,N_4442,N_4190);
and U4594 (N_4594,N_4299,N_4107);
nand U4595 (N_4595,N_4429,N_4421);
or U4596 (N_4596,N_4478,N_4432);
nor U4597 (N_4597,N_4477,N_4082);
nor U4598 (N_4598,N_4088,N_4036);
nand U4599 (N_4599,N_4464,N_4110);
nor U4600 (N_4600,N_4492,N_4124);
nor U4601 (N_4601,N_4476,N_4236);
nand U4602 (N_4602,N_4361,N_4424);
and U4603 (N_4603,N_4111,N_4096);
or U4604 (N_4604,N_4320,N_4285);
and U4605 (N_4605,N_4280,N_4337);
and U4606 (N_4606,N_4245,N_4397);
and U4607 (N_4607,N_4038,N_4404);
or U4608 (N_4608,N_4157,N_4266);
and U4609 (N_4609,N_4193,N_4063);
nor U4610 (N_4610,N_4413,N_4000);
nor U4611 (N_4611,N_4281,N_4379);
or U4612 (N_4612,N_4077,N_4175);
nor U4613 (N_4613,N_4097,N_4367);
nor U4614 (N_4614,N_4127,N_4004);
and U4615 (N_4615,N_4153,N_4220);
or U4616 (N_4616,N_4309,N_4261);
and U4617 (N_4617,N_4444,N_4056);
nand U4618 (N_4618,N_4376,N_4028);
and U4619 (N_4619,N_4254,N_4115);
nor U4620 (N_4620,N_4047,N_4132);
nand U4621 (N_4621,N_4138,N_4092);
and U4622 (N_4622,N_4099,N_4141);
nand U4623 (N_4623,N_4058,N_4395);
nand U4624 (N_4624,N_4428,N_4339);
nor U4625 (N_4625,N_4450,N_4085);
or U4626 (N_4626,N_4278,N_4183);
nor U4627 (N_4627,N_4265,N_4074);
and U4628 (N_4628,N_4364,N_4290);
and U4629 (N_4629,N_4382,N_4439);
nor U4630 (N_4630,N_4259,N_4101);
and U4631 (N_4631,N_4113,N_4437);
and U4632 (N_4632,N_4081,N_4200);
and U4633 (N_4633,N_4250,N_4143);
nand U4634 (N_4634,N_4191,N_4405);
nand U4635 (N_4635,N_4431,N_4035);
nor U4636 (N_4636,N_4178,N_4398);
xor U4637 (N_4637,N_4396,N_4332);
nand U4638 (N_4638,N_4207,N_4357);
or U4639 (N_4639,N_4331,N_4103);
and U4640 (N_4640,N_4005,N_4211);
nand U4641 (N_4641,N_4375,N_4119);
nand U4642 (N_4642,N_4196,N_4147);
nand U4643 (N_4643,N_4075,N_4336);
and U4644 (N_4644,N_4468,N_4062);
nand U4645 (N_4645,N_4205,N_4065);
and U4646 (N_4646,N_4233,N_4388);
and U4647 (N_4647,N_4022,N_4061);
nand U4648 (N_4648,N_4169,N_4350);
nand U4649 (N_4649,N_4260,N_4146);
or U4650 (N_4650,N_4284,N_4244);
or U4651 (N_4651,N_4384,N_4277);
and U4652 (N_4652,N_4192,N_4295);
nand U4653 (N_4653,N_4471,N_4197);
and U4654 (N_4654,N_4031,N_4348);
or U4655 (N_4655,N_4171,N_4385);
and U4656 (N_4656,N_4010,N_4131);
and U4657 (N_4657,N_4068,N_4136);
and U4658 (N_4658,N_4234,N_4455);
nor U4659 (N_4659,N_4137,N_4394);
nor U4660 (N_4660,N_4467,N_4351);
or U4661 (N_4661,N_4340,N_4173);
or U4662 (N_4662,N_4317,N_4212);
or U4663 (N_4663,N_4316,N_4072);
and U4664 (N_4664,N_4011,N_4176);
nand U4665 (N_4665,N_4313,N_4229);
nor U4666 (N_4666,N_4079,N_4144);
or U4667 (N_4667,N_4255,N_4186);
and U4668 (N_4668,N_4344,N_4116);
and U4669 (N_4669,N_4021,N_4118);
or U4670 (N_4670,N_4449,N_4377);
nor U4671 (N_4671,N_4057,N_4145);
and U4672 (N_4672,N_4014,N_4042);
nand U4673 (N_4673,N_4423,N_4084);
and U4674 (N_4674,N_4302,N_4055);
nor U4675 (N_4675,N_4345,N_4158);
and U4676 (N_4676,N_4015,N_4213);
or U4677 (N_4677,N_4494,N_4420);
or U4678 (N_4678,N_4293,N_4154);
nor U4679 (N_4679,N_4322,N_4222);
nand U4680 (N_4680,N_4402,N_4263);
and U4681 (N_4681,N_4201,N_4461);
nor U4682 (N_4682,N_4443,N_4209);
and U4683 (N_4683,N_4002,N_4202);
and U4684 (N_4684,N_4106,N_4488);
and U4685 (N_4685,N_4358,N_4039);
and U4686 (N_4686,N_4451,N_4273);
nor U4687 (N_4687,N_4425,N_4227);
or U4688 (N_4688,N_4366,N_4018);
nor U4689 (N_4689,N_4179,N_4417);
and U4690 (N_4690,N_4329,N_4426);
nand U4691 (N_4691,N_4419,N_4095);
nand U4692 (N_4692,N_4023,N_4090);
nor U4693 (N_4693,N_4120,N_4447);
and U4694 (N_4694,N_4030,N_4412);
xor U4695 (N_4695,N_4334,N_4486);
nand U4696 (N_4696,N_4164,N_4495);
or U4697 (N_4697,N_4466,N_4078);
nor U4698 (N_4698,N_4460,N_4165);
and U4699 (N_4699,N_4114,N_4386);
nand U4700 (N_4700,N_4275,N_4098);
nand U4701 (N_4701,N_4240,N_4399);
nor U4702 (N_4702,N_4117,N_4459);
or U4703 (N_4703,N_4303,N_4267);
nand U4704 (N_4704,N_4109,N_4446);
and U4705 (N_4705,N_4024,N_4237);
nand U4706 (N_4706,N_4308,N_4287);
nand U4707 (N_4707,N_4054,N_4252);
xor U4708 (N_4708,N_4325,N_4408);
nor U4709 (N_4709,N_4324,N_4291);
nand U4710 (N_4710,N_4087,N_4403);
or U4711 (N_4711,N_4155,N_4411);
nor U4712 (N_4712,N_4435,N_4283);
nand U4713 (N_4713,N_4479,N_4247);
nand U4714 (N_4714,N_4040,N_4481);
or U4715 (N_4715,N_4418,N_4262);
nor U4716 (N_4716,N_4241,N_4389);
or U4717 (N_4717,N_4177,N_4140);
nand U4718 (N_4718,N_4314,N_4289);
and U4719 (N_4719,N_4216,N_4362);
xnor U4720 (N_4720,N_4025,N_4214);
and U4721 (N_4721,N_4188,N_4341);
nor U4722 (N_4722,N_4312,N_4045);
nor U4723 (N_4723,N_4251,N_4490);
nand U4724 (N_4724,N_4066,N_4465);
nand U4725 (N_4725,N_4203,N_4387);
nor U4726 (N_4726,N_4304,N_4198);
or U4727 (N_4727,N_4033,N_4393);
nor U4728 (N_4728,N_4129,N_4243);
nor U4729 (N_4729,N_4373,N_4342);
and U4730 (N_4730,N_4160,N_4370);
nand U4731 (N_4731,N_4151,N_4059);
nor U4732 (N_4732,N_4231,N_4105);
and U4733 (N_4733,N_4219,N_4167);
and U4734 (N_4734,N_4194,N_4301);
nor U4735 (N_4735,N_4391,N_4162);
nor U4736 (N_4736,N_4206,N_4257);
nor U4737 (N_4737,N_4327,N_4034);
nand U4738 (N_4738,N_4189,N_4484);
nor U4739 (N_4739,N_4415,N_4292);
and U4740 (N_4740,N_4296,N_4383);
nand U4741 (N_4741,N_4270,N_4427);
nand U4742 (N_4742,N_4187,N_4430);
nand U4743 (N_4743,N_4359,N_4123);
or U4744 (N_4744,N_4037,N_4049);
and U4745 (N_4745,N_4001,N_4142);
and U4746 (N_4746,N_4060,N_4352);
or U4747 (N_4747,N_4497,N_4174);
or U4748 (N_4748,N_4208,N_4221);
or U4749 (N_4749,N_4410,N_4482);
or U4750 (N_4750,N_4252,N_4374);
nor U4751 (N_4751,N_4313,N_4462);
nor U4752 (N_4752,N_4359,N_4093);
nand U4753 (N_4753,N_4496,N_4041);
or U4754 (N_4754,N_4247,N_4120);
nand U4755 (N_4755,N_4458,N_4392);
nand U4756 (N_4756,N_4167,N_4273);
nor U4757 (N_4757,N_4191,N_4083);
and U4758 (N_4758,N_4242,N_4019);
and U4759 (N_4759,N_4391,N_4436);
nand U4760 (N_4760,N_4247,N_4446);
and U4761 (N_4761,N_4065,N_4200);
nand U4762 (N_4762,N_4232,N_4094);
and U4763 (N_4763,N_4328,N_4267);
or U4764 (N_4764,N_4320,N_4125);
nor U4765 (N_4765,N_4021,N_4375);
and U4766 (N_4766,N_4494,N_4330);
or U4767 (N_4767,N_4197,N_4092);
or U4768 (N_4768,N_4048,N_4333);
nor U4769 (N_4769,N_4350,N_4486);
or U4770 (N_4770,N_4229,N_4322);
nor U4771 (N_4771,N_4122,N_4458);
and U4772 (N_4772,N_4203,N_4386);
nand U4773 (N_4773,N_4024,N_4072);
and U4774 (N_4774,N_4006,N_4387);
and U4775 (N_4775,N_4336,N_4464);
or U4776 (N_4776,N_4049,N_4178);
nand U4777 (N_4777,N_4356,N_4431);
nand U4778 (N_4778,N_4302,N_4190);
or U4779 (N_4779,N_4321,N_4161);
and U4780 (N_4780,N_4050,N_4298);
nor U4781 (N_4781,N_4454,N_4035);
or U4782 (N_4782,N_4249,N_4270);
nor U4783 (N_4783,N_4285,N_4453);
nand U4784 (N_4784,N_4040,N_4104);
nand U4785 (N_4785,N_4040,N_4322);
and U4786 (N_4786,N_4491,N_4309);
nand U4787 (N_4787,N_4257,N_4046);
nor U4788 (N_4788,N_4187,N_4350);
and U4789 (N_4789,N_4493,N_4285);
or U4790 (N_4790,N_4275,N_4120);
nor U4791 (N_4791,N_4043,N_4117);
nand U4792 (N_4792,N_4212,N_4120);
nand U4793 (N_4793,N_4254,N_4445);
and U4794 (N_4794,N_4321,N_4282);
or U4795 (N_4795,N_4401,N_4206);
or U4796 (N_4796,N_4322,N_4328);
nor U4797 (N_4797,N_4025,N_4390);
nand U4798 (N_4798,N_4240,N_4438);
or U4799 (N_4799,N_4345,N_4383);
nor U4800 (N_4800,N_4021,N_4247);
or U4801 (N_4801,N_4415,N_4051);
nor U4802 (N_4802,N_4080,N_4485);
nor U4803 (N_4803,N_4217,N_4030);
nand U4804 (N_4804,N_4330,N_4232);
xor U4805 (N_4805,N_4309,N_4116);
and U4806 (N_4806,N_4148,N_4231);
and U4807 (N_4807,N_4181,N_4473);
or U4808 (N_4808,N_4202,N_4311);
xnor U4809 (N_4809,N_4028,N_4018);
or U4810 (N_4810,N_4322,N_4493);
or U4811 (N_4811,N_4431,N_4383);
and U4812 (N_4812,N_4184,N_4169);
or U4813 (N_4813,N_4425,N_4450);
nor U4814 (N_4814,N_4359,N_4429);
nand U4815 (N_4815,N_4424,N_4093);
nand U4816 (N_4816,N_4126,N_4435);
and U4817 (N_4817,N_4249,N_4387);
nor U4818 (N_4818,N_4380,N_4416);
or U4819 (N_4819,N_4136,N_4066);
or U4820 (N_4820,N_4390,N_4083);
nor U4821 (N_4821,N_4274,N_4130);
or U4822 (N_4822,N_4074,N_4348);
nor U4823 (N_4823,N_4031,N_4213);
nand U4824 (N_4824,N_4166,N_4476);
nor U4825 (N_4825,N_4070,N_4337);
nor U4826 (N_4826,N_4022,N_4296);
and U4827 (N_4827,N_4284,N_4421);
nor U4828 (N_4828,N_4209,N_4393);
nor U4829 (N_4829,N_4070,N_4379);
nand U4830 (N_4830,N_4336,N_4104);
and U4831 (N_4831,N_4044,N_4162);
nand U4832 (N_4832,N_4323,N_4318);
or U4833 (N_4833,N_4226,N_4286);
nor U4834 (N_4834,N_4460,N_4175);
and U4835 (N_4835,N_4365,N_4037);
nor U4836 (N_4836,N_4455,N_4055);
nor U4837 (N_4837,N_4185,N_4175);
or U4838 (N_4838,N_4246,N_4245);
or U4839 (N_4839,N_4220,N_4389);
and U4840 (N_4840,N_4310,N_4134);
nor U4841 (N_4841,N_4118,N_4482);
or U4842 (N_4842,N_4422,N_4015);
nand U4843 (N_4843,N_4318,N_4023);
or U4844 (N_4844,N_4289,N_4317);
nand U4845 (N_4845,N_4077,N_4078);
and U4846 (N_4846,N_4451,N_4160);
nand U4847 (N_4847,N_4488,N_4218);
nand U4848 (N_4848,N_4053,N_4471);
or U4849 (N_4849,N_4465,N_4173);
and U4850 (N_4850,N_4376,N_4254);
or U4851 (N_4851,N_4456,N_4274);
nand U4852 (N_4852,N_4015,N_4244);
and U4853 (N_4853,N_4147,N_4343);
or U4854 (N_4854,N_4211,N_4185);
nand U4855 (N_4855,N_4468,N_4249);
nand U4856 (N_4856,N_4451,N_4353);
or U4857 (N_4857,N_4361,N_4452);
xor U4858 (N_4858,N_4192,N_4079);
nor U4859 (N_4859,N_4336,N_4183);
or U4860 (N_4860,N_4203,N_4105);
xor U4861 (N_4861,N_4239,N_4359);
nor U4862 (N_4862,N_4201,N_4023);
nor U4863 (N_4863,N_4220,N_4091);
nand U4864 (N_4864,N_4195,N_4201);
or U4865 (N_4865,N_4256,N_4220);
and U4866 (N_4866,N_4279,N_4021);
nand U4867 (N_4867,N_4341,N_4064);
nand U4868 (N_4868,N_4040,N_4144);
or U4869 (N_4869,N_4433,N_4454);
nor U4870 (N_4870,N_4226,N_4155);
nand U4871 (N_4871,N_4202,N_4371);
nand U4872 (N_4872,N_4194,N_4003);
or U4873 (N_4873,N_4288,N_4277);
nand U4874 (N_4874,N_4045,N_4454);
or U4875 (N_4875,N_4196,N_4284);
nand U4876 (N_4876,N_4067,N_4328);
nor U4877 (N_4877,N_4125,N_4118);
or U4878 (N_4878,N_4010,N_4370);
and U4879 (N_4879,N_4339,N_4395);
or U4880 (N_4880,N_4418,N_4358);
or U4881 (N_4881,N_4180,N_4178);
nand U4882 (N_4882,N_4468,N_4211);
nor U4883 (N_4883,N_4363,N_4112);
nor U4884 (N_4884,N_4135,N_4403);
nand U4885 (N_4885,N_4423,N_4078);
or U4886 (N_4886,N_4380,N_4127);
or U4887 (N_4887,N_4107,N_4324);
or U4888 (N_4888,N_4384,N_4198);
nor U4889 (N_4889,N_4145,N_4264);
nor U4890 (N_4890,N_4453,N_4056);
nand U4891 (N_4891,N_4288,N_4068);
nor U4892 (N_4892,N_4151,N_4491);
or U4893 (N_4893,N_4033,N_4400);
or U4894 (N_4894,N_4072,N_4331);
and U4895 (N_4895,N_4234,N_4084);
and U4896 (N_4896,N_4015,N_4464);
nand U4897 (N_4897,N_4003,N_4337);
nor U4898 (N_4898,N_4150,N_4281);
nand U4899 (N_4899,N_4074,N_4444);
or U4900 (N_4900,N_4268,N_4253);
or U4901 (N_4901,N_4410,N_4478);
nand U4902 (N_4902,N_4075,N_4034);
and U4903 (N_4903,N_4089,N_4084);
nand U4904 (N_4904,N_4242,N_4275);
nor U4905 (N_4905,N_4161,N_4111);
nor U4906 (N_4906,N_4261,N_4270);
nand U4907 (N_4907,N_4399,N_4455);
nand U4908 (N_4908,N_4448,N_4015);
and U4909 (N_4909,N_4486,N_4093);
and U4910 (N_4910,N_4412,N_4094);
nor U4911 (N_4911,N_4451,N_4209);
or U4912 (N_4912,N_4267,N_4154);
nand U4913 (N_4913,N_4272,N_4479);
nand U4914 (N_4914,N_4084,N_4476);
nand U4915 (N_4915,N_4220,N_4217);
nand U4916 (N_4916,N_4108,N_4041);
or U4917 (N_4917,N_4163,N_4138);
or U4918 (N_4918,N_4203,N_4098);
or U4919 (N_4919,N_4250,N_4156);
and U4920 (N_4920,N_4161,N_4143);
or U4921 (N_4921,N_4339,N_4474);
and U4922 (N_4922,N_4087,N_4485);
or U4923 (N_4923,N_4322,N_4022);
or U4924 (N_4924,N_4269,N_4353);
nand U4925 (N_4925,N_4321,N_4444);
or U4926 (N_4926,N_4195,N_4471);
nor U4927 (N_4927,N_4160,N_4470);
or U4928 (N_4928,N_4118,N_4137);
nor U4929 (N_4929,N_4457,N_4065);
or U4930 (N_4930,N_4404,N_4040);
and U4931 (N_4931,N_4145,N_4138);
nor U4932 (N_4932,N_4215,N_4177);
or U4933 (N_4933,N_4465,N_4401);
or U4934 (N_4934,N_4299,N_4127);
and U4935 (N_4935,N_4174,N_4381);
nand U4936 (N_4936,N_4402,N_4269);
or U4937 (N_4937,N_4031,N_4054);
and U4938 (N_4938,N_4396,N_4415);
nand U4939 (N_4939,N_4258,N_4354);
or U4940 (N_4940,N_4053,N_4120);
xor U4941 (N_4941,N_4283,N_4100);
nand U4942 (N_4942,N_4093,N_4328);
or U4943 (N_4943,N_4196,N_4168);
and U4944 (N_4944,N_4255,N_4371);
xnor U4945 (N_4945,N_4391,N_4318);
nand U4946 (N_4946,N_4390,N_4439);
nand U4947 (N_4947,N_4156,N_4270);
or U4948 (N_4948,N_4156,N_4373);
nand U4949 (N_4949,N_4369,N_4025);
nand U4950 (N_4950,N_4404,N_4415);
nand U4951 (N_4951,N_4357,N_4442);
nand U4952 (N_4952,N_4459,N_4222);
and U4953 (N_4953,N_4452,N_4097);
or U4954 (N_4954,N_4459,N_4482);
or U4955 (N_4955,N_4446,N_4205);
nor U4956 (N_4956,N_4264,N_4032);
nor U4957 (N_4957,N_4268,N_4402);
or U4958 (N_4958,N_4045,N_4433);
or U4959 (N_4959,N_4427,N_4485);
nor U4960 (N_4960,N_4472,N_4312);
nor U4961 (N_4961,N_4114,N_4408);
or U4962 (N_4962,N_4298,N_4111);
nand U4963 (N_4963,N_4250,N_4000);
nand U4964 (N_4964,N_4147,N_4076);
nor U4965 (N_4965,N_4005,N_4039);
nand U4966 (N_4966,N_4003,N_4489);
nor U4967 (N_4967,N_4306,N_4027);
nor U4968 (N_4968,N_4191,N_4464);
or U4969 (N_4969,N_4199,N_4313);
and U4970 (N_4970,N_4074,N_4126);
nand U4971 (N_4971,N_4002,N_4103);
nor U4972 (N_4972,N_4194,N_4308);
and U4973 (N_4973,N_4497,N_4132);
nor U4974 (N_4974,N_4202,N_4063);
and U4975 (N_4975,N_4118,N_4104);
and U4976 (N_4976,N_4489,N_4495);
or U4977 (N_4977,N_4171,N_4093);
or U4978 (N_4978,N_4373,N_4137);
nor U4979 (N_4979,N_4252,N_4235);
nand U4980 (N_4980,N_4391,N_4258);
nor U4981 (N_4981,N_4164,N_4399);
xnor U4982 (N_4982,N_4312,N_4135);
xor U4983 (N_4983,N_4280,N_4114);
nor U4984 (N_4984,N_4378,N_4473);
or U4985 (N_4985,N_4458,N_4120);
and U4986 (N_4986,N_4286,N_4019);
xnor U4987 (N_4987,N_4455,N_4200);
nor U4988 (N_4988,N_4160,N_4165);
nor U4989 (N_4989,N_4220,N_4089);
or U4990 (N_4990,N_4083,N_4338);
xnor U4991 (N_4991,N_4388,N_4293);
or U4992 (N_4992,N_4419,N_4431);
or U4993 (N_4993,N_4062,N_4269);
and U4994 (N_4994,N_4490,N_4392);
and U4995 (N_4995,N_4238,N_4436);
or U4996 (N_4996,N_4255,N_4076);
or U4997 (N_4997,N_4226,N_4051);
nand U4998 (N_4998,N_4175,N_4124);
nand U4999 (N_4999,N_4095,N_4302);
nor U5000 (N_5000,N_4823,N_4842);
and U5001 (N_5001,N_4696,N_4604);
and U5002 (N_5002,N_4839,N_4652);
nand U5003 (N_5003,N_4924,N_4727);
or U5004 (N_5004,N_4755,N_4845);
nor U5005 (N_5005,N_4753,N_4664);
nand U5006 (N_5006,N_4894,N_4650);
or U5007 (N_5007,N_4951,N_4939);
or U5008 (N_5008,N_4521,N_4678);
nand U5009 (N_5009,N_4607,N_4904);
nand U5010 (N_5010,N_4587,N_4718);
nand U5011 (N_5011,N_4902,N_4527);
nand U5012 (N_5012,N_4712,N_4819);
xor U5013 (N_5013,N_4682,N_4513);
and U5014 (N_5014,N_4549,N_4877);
nand U5015 (N_5015,N_4929,N_4608);
nor U5016 (N_5016,N_4730,N_4990);
nor U5017 (N_5017,N_4618,N_4945);
or U5018 (N_5018,N_4593,N_4961);
and U5019 (N_5019,N_4956,N_4884);
nand U5020 (N_5020,N_4970,N_4706);
nand U5021 (N_5021,N_4594,N_4849);
nand U5022 (N_5022,N_4725,N_4556);
and U5023 (N_5023,N_4530,N_4954);
nand U5024 (N_5024,N_4704,N_4735);
nor U5025 (N_5025,N_4994,N_4509);
nand U5026 (N_5026,N_4835,N_4570);
nand U5027 (N_5027,N_4818,N_4564);
or U5028 (N_5028,N_4599,N_4827);
nand U5029 (N_5029,N_4757,N_4810);
nor U5030 (N_5030,N_4986,N_4680);
xor U5031 (N_5031,N_4825,N_4501);
nand U5032 (N_5032,N_4901,N_4559);
and U5033 (N_5033,N_4841,N_4947);
nor U5034 (N_5034,N_4623,N_4751);
nor U5035 (N_5035,N_4523,N_4703);
nand U5036 (N_5036,N_4790,N_4885);
or U5037 (N_5037,N_4806,N_4563);
nand U5038 (N_5038,N_4567,N_4701);
nand U5039 (N_5039,N_4848,N_4890);
and U5040 (N_5040,N_4948,N_4740);
nand U5041 (N_5041,N_4505,N_4989);
nand U5042 (N_5042,N_4940,N_4565);
nand U5043 (N_5043,N_4893,N_4869);
nor U5044 (N_5044,N_4524,N_4719);
nor U5045 (N_5045,N_4975,N_4714);
nand U5046 (N_5046,N_4526,N_4661);
or U5047 (N_5047,N_4761,N_4746);
or U5048 (N_5048,N_4566,N_4511);
nand U5049 (N_5049,N_4831,N_4871);
or U5050 (N_5050,N_4583,N_4649);
nor U5051 (N_5051,N_4996,N_4908);
or U5052 (N_5052,N_4872,N_4729);
or U5053 (N_5053,N_4504,N_4590);
or U5054 (N_5054,N_4648,N_4610);
or U5055 (N_5055,N_4912,N_4972);
nand U5056 (N_5056,N_4782,N_4540);
or U5057 (N_5057,N_4919,N_4809);
or U5058 (N_5058,N_4734,N_4721);
nor U5059 (N_5059,N_4829,N_4770);
nor U5060 (N_5060,N_4634,N_4744);
nand U5061 (N_5061,N_4942,N_4612);
or U5062 (N_5062,N_4969,N_4531);
nor U5063 (N_5063,N_4820,N_4837);
and U5064 (N_5064,N_4817,N_4539);
and U5065 (N_5065,N_4802,N_4597);
nand U5066 (N_5066,N_4516,N_4533);
or U5067 (N_5067,N_4974,N_4697);
or U5068 (N_5068,N_4798,N_4752);
nand U5069 (N_5069,N_4870,N_4762);
or U5070 (N_5070,N_4874,N_4868);
nor U5071 (N_5071,N_4949,N_4592);
nor U5072 (N_5072,N_4659,N_4569);
nor U5073 (N_5073,N_4671,N_4713);
and U5074 (N_5074,N_4911,N_4637);
and U5075 (N_5075,N_4535,N_4934);
and U5076 (N_5076,N_4875,N_4500);
and U5077 (N_5077,N_4621,N_4657);
and U5078 (N_5078,N_4510,N_4863);
nor U5079 (N_5079,N_4532,N_4591);
nor U5080 (N_5080,N_4813,N_4895);
nand U5081 (N_5081,N_4873,N_4957);
and U5082 (N_5082,N_4792,N_4838);
nor U5083 (N_5083,N_4794,N_4705);
nor U5084 (N_5084,N_4528,N_4596);
xor U5085 (N_5085,N_4546,N_4759);
nand U5086 (N_5086,N_4675,N_4936);
nor U5087 (N_5087,N_4891,N_4653);
nor U5088 (N_5088,N_4991,N_4976);
nor U5089 (N_5089,N_4545,N_4834);
nor U5090 (N_5090,N_4879,N_4828);
and U5091 (N_5091,N_4800,N_4844);
and U5092 (N_5092,N_4686,N_4937);
or U5093 (N_5093,N_4965,N_4950);
nor U5094 (N_5094,N_4958,N_4938);
and U5095 (N_5095,N_4690,N_4645);
xor U5096 (N_5096,N_4867,N_4995);
and U5097 (N_5097,N_4931,N_4896);
xor U5098 (N_5098,N_4581,N_4639);
or U5099 (N_5099,N_4773,N_4674);
or U5100 (N_5100,N_4625,N_4700);
and U5101 (N_5101,N_4677,N_4756);
or U5102 (N_5102,N_4771,N_4562);
nor U5103 (N_5103,N_4736,N_4585);
or U5104 (N_5104,N_4672,N_4638);
nand U5105 (N_5105,N_4611,N_4913);
and U5106 (N_5106,N_4508,N_4766);
and U5107 (N_5107,N_4855,N_4656);
and U5108 (N_5108,N_4830,N_4903);
nand U5109 (N_5109,N_4624,N_4886);
and U5110 (N_5110,N_4517,N_4915);
nor U5111 (N_5111,N_4507,N_4655);
nor U5112 (N_5112,N_4749,N_4676);
nand U5113 (N_5113,N_4693,N_4629);
nor U5114 (N_5114,N_4575,N_4742);
and U5115 (N_5115,N_4537,N_4925);
nor U5116 (N_5116,N_4804,N_4654);
xnor U5117 (N_5117,N_4963,N_4826);
and U5118 (N_5118,N_4843,N_4660);
or U5119 (N_5119,N_4574,N_4797);
nand U5120 (N_5120,N_4909,N_4640);
nor U5121 (N_5121,N_4600,N_4927);
nor U5122 (N_5122,N_4914,N_4750);
nand U5123 (N_5123,N_4850,N_4709);
or U5124 (N_5124,N_4987,N_4979);
nor U5125 (N_5125,N_4662,N_4998);
and U5126 (N_5126,N_4805,N_4907);
nor U5127 (N_5127,N_4864,N_4856);
or U5128 (N_5128,N_4905,N_4557);
xor U5129 (N_5129,N_4616,N_4635);
and U5130 (N_5130,N_4647,N_4821);
nor U5131 (N_5131,N_4941,N_4763);
and U5132 (N_5132,N_4738,N_4605);
nand U5133 (N_5133,N_4920,N_4555);
nor U5134 (N_5134,N_4775,N_4536);
nor U5135 (N_5135,N_4542,N_4568);
nand U5136 (N_5136,N_4964,N_4741);
or U5137 (N_5137,N_4959,N_4808);
and U5138 (N_5138,N_4966,N_4960);
xor U5139 (N_5139,N_4814,N_4632);
nor U5140 (N_5140,N_4999,N_4561);
nor U5141 (N_5141,N_4926,N_4514);
nor U5142 (N_5142,N_4681,N_4862);
or U5143 (N_5143,N_4900,N_4578);
nor U5144 (N_5144,N_4997,N_4589);
or U5145 (N_5145,N_4670,N_4883);
and U5146 (N_5146,N_4646,N_4962);
nand U5147 (N_5147,N_4717,N_4642);
nor U5148 (N_5148,N_4691,N_4620);
nor U5149 (N_5149,N_4627,N_4609);
nand U5150 (N_5150,N_4781,N_4933);
or U5151 (N_5151,N_4558,N_4506);
nor U5152 (N_5152,N_4853,N_4985);
and U5153 (N_5153,N_4622,N_4876);
nor U5154 (N_5154,N_4685,N_4636);
or U5155 (N_5155,N_4707,N_4765);
and U5156 (N_5156,N_4881,N_4538);
and U5157 (N_5157,N_4764,N_4550);
nor U5158 (N_5158,N_4784,N_4777);
xor U5159 (N_5159,N_4667,N_4586);
nand U5160 (N_5160,N_4518,N_4541);
and U5161 (N_5161,N_4923,N_4666);
xnor U5162 (N_5162,N_4577,N_4595);
and U5163 (N_5163,N_4882,N_4815);
nor U5164 (N_5164,N_4669,N_4836);
or U5165 (N_5165,N_4728,N_4534);
nand U5166 (N_5166,N_4613,N_4971);
and U5167 (N_5167,N_4519,N_4658);
or U5168 (N_5168,N_4711,N_4588);
nand U5169 (N_5169,N_4779,N_4822);
nor U5170 (N_5170,N_4952,N_4968);
nor U5171 (N_5171,N_4715,N_4633);
nand U5172 (N_5172,N_4854,N_4878);
or U5173 (N_5173,N_4967,N_4906);
nand U5174 (N_5174,N_4768,N_4643);
or U5175 (N_5175,N_4572,N_4816);
nand U5176 (N_5176,N_4791,N_4880);
nand U5177 (N_5177,N_4503,N_4598);
nand U5178 (N_5178,N_4930,N_4673);
nor U5179 (N_5179,N_4758,N_4573);
nor U5180 (N_5180,N_4796,N_4702);
nor U5181 (N_5181,N_4858,N_4847);
nor U5182 (N_5182,N_4603,N_4668);
or U5183 (N_5183,N_4793,N_4722);
nor U5184 (N_5184,N_4789,N_4552);
or U5185 (N_5185,N_4747,N_4774);
or U5186 (N_5186,N_4692,N_4888);
nand U5187 (N_5187,N_4543,N_4785);
or U5188 (N_5188,N_4724,N_4776);
or U5189 (N_5189,N_4512,N_4601);
and U5190 (N_5190,N_4644,N_4859);
nand U5191 (N_5191,N_4866,N_4992);
nor U5192 (N_5192,N_4628,N_4783);
nand U5193 (N_5193,N_4743,N_4795);
nor U5194 (N_5194,N_4665,N_4944);
or U5195 (N_5195,N_4619,N_4502);
nand U5196 (N_5196,N_4767,N_4739);
or U5197 (N_5197,N_4860,N_4731);
nand U5198 (N_5198,N_4547,N_4553);
nor U5199 (N_5199,N_4892,N_4695);
nor U5200 (N_5200,N_4571,N_4852);
or U5201 (N_5201,N_4641,N_4769);
and U5202 (N_5202,N_4544,N_4993);
and U5203 (N_5203,N_4584,N_4683);
and U5204 (N_5204,N_4694,N_4840);
and U5205 (N_5205,N_4529,N_4630);
and U5206 (N_5206,N_4811,N_4807);
nand U5207 (N_5207,N_4684,N_4617);
nand U5208 (N_5208,N_4861,N_4732);
or U5209 (N_5209,N_4663,N_4688);
or U5210 (N_5210,N_4955,N_4887);
nor U5211 (N_5211,N_4799,N_4928);
and U5212 (N_5212,N_4679,N_4716);
and U5213 (N_5213,N_4726,N_4626);
and U5214 (N_5214,N_4614,N_4921);
nor U5215 (N_5215,N_4548,N_4982);
nor U5216 (N_5216,N_4737,N_4778);
and U5217 (N_5217,N_4917,N_4788);
nor U5218 (N_5218,N_4978,N_4606);
and U5219 (N_5219,N_4922,N_4824);
nand U5220 (N_5220,N_4801,N_4710);
and U5221 (N_5221,N_4576,N_4720);
nor U5222 (N_5222,N_4897,N_4733);
nand U5223 (N_5223,N_4698,N_4832);
xor U5224 (N_5224,N_4651,N_4943);
and U5225 (N_5225,N_4786,N_4803);
and U5226 (N_5226,N_4515,N_4525);
and U5227 (N_5227,N_4946,N_4787);
or U5228 (N_5228,N_4580,N_4579);
nor U5229 (N_5229,N_4916,N_4602);
and U5230 (N_5230,N_4899,N_4699);
xor U5231 (N_5231,N_4889,N_4812);
nor U5232 (N_5232,N_4973,N_4551);
or U5233 (N_5233,N_4520,N_4865);
nand U5234 (N_5234,N_4745,N_4898);
or U5235 (N_5235,N_4932,N_4689);
nand U5236 (N_5236,N_4687,N_4615);
or U5237 (N_5237,N_4582,N_4983);
nor U5238 (N_5238,N_4723,N_4833);
nand U5239 (N_5239,N_4554,N_4953);
and U5240 (N_5240,N_4760,N_4748);
or U5241 (N_5241,N_4631,N_4772);
and U5242 (N_5242,N_4910,N_4918);
or U5243 (N_5243,N_4560,N_4857);
nor U5244 (N_5244,N_4851,N_4988);
or U5245 (N_5245,N_4935,N_4780);
nor U5246 (N_5246,N_4977,N_4984);
and U5247 (N_5247,N_4708,N_4981);
and U5248 (N_5248,N_4754,N_4522);
and U5249 (N_5249,N_4846,N_4980);
and U5250 (N_5250,N_4947,N_4533);
nor U5251 (N_5251,N_4888,N_4804);
nand U5252 (N_5252,N_4572,N_4825);
nor U5253 (N_5253,N_4956,N_4710);
nand U5254 (N_5254,N_4550,N_4657);
nand U5255 (N_5255,N_4683,N_4861);
or U5256 (N_5256,N_4787,N_4800);
or U5257 (N_5257,N_4963,N_4511);
nor U5258 (N_5258,N_4806,N_4786);
nand U5259 (N_5259,N_4807,N_4789);
or U5260 (N_5260,N_4684,N_4910);
nand U5261 (N_5261,N_4863,N_4719);
and U5262 (N_5262,N_4881,N_4817);
nor U5263 (N_5263,N_4643,N_4847);
nand U5264 (N_5264,N_4910,N_4570);
or U5265 (N_5265,N_4855,N_4622);
and U5266 (N_5266,N_4729,N_4657);
or U5267 (N_5267,N_4687,N_4662);
and U5268 (N_5268,N_4517,N_4960);
or U5269 (N_5269,N_4571,N_4983);
or U5270 (N_5270,N_4899,N_4732);
or U5271 (N_5271,N_4910,N_4957);
and U5272 (N_5272,N_4909,N_4617);
and U5273 (N_5273,N_4558,N_4902);
nand U5274 (N_5274,N_4973,N_4594);
nand U5275 (N_5275,N_4973,N_4527);
and U5276 (N_5276,N_4756,N_4520);
or U5277 (N_5277,N_4922,N_4664);
nor U5278 (N_5278,N_4740,N_4525);
and U5279 (N_5279,N_4808,N_4816);
nand U5280 (N_5280,N_4869,N_4717);
or U5281 (N_5281,N_4940,N_4856);
or U5282 (N_5282,N_4790,N_4898);
nor U5283 (N_5283,N_4655,N_4513);
nor U5284 (N_5284,N_4617,N_4813);
and U5285 (N_5285,N_4719,N_4993);
and U5286 (N_5286,N_4857,N_4904);
nand U5287 (N_5287,N_4671,N_4835);
and U5288 (N_5288,N_4748,N_4957);
or U5289 (N_5289,N_4537,N_4598);
or U5290 (N_5290,N_4880,N_4819);
nor U5291 (N_5291,N_4520,N_4745);
nor U5292 (N_5292,N_4886,N_4815);
and U5293 (N_5293,N_4964,N_4596);
or U5294 (N_5294,N_4690,N_4916);
nor U5295 (N_5295,N_4751,N_4687);
nor U5296 (N_5296,N_4712,N_4537);
and U5297 (N_5297,N_4957,N_4665);
nand U5298 (N_5298,N_4934,N_4929);
nor U5299 (N_5299,N_4674,N_4553);
or U5300 (N_5300,N_4971,N_4988);
nand U5301 (N_5301,N_4790,N_4783);
nand U5302 (N_5302,N_4570,N_4974);
and U5303 (N_5303,N_4867,N_4525);
nor U5304 (N_5304,N_4650,N_4967);
nor U5305 (N_5305,N_4790,N_4956);
nor U5306 (N_5306,N_4686,N_4766);
nand U5307 (N_5307,N_4641,N_4668);
or U5308 (N_5308,N_4850,N_4583);
nand U5309 (N_5309,N_4829,N_4712);
nand U5310 (N_5310,N_4694,N_4837);
nand U5311 (N_5311,N_4941,N_4520);
nor U5312 (N_5312,N_4872,N_4797);
nor U5313 (N_5313,N_4648,N_4923);
nor U5314 (N_5314,N_4973,N_4937);
nand U5315 (N_5315,N_4576,N_4525);
nor U5316 (N_5316,N_4801,N_4537);
or U5317 (N_5317,N_4679,N_4734);
nand U5318 (N_5318,N_4683,N_4854);
nand U5319 (N_5319,N_4994,N_4899);
nor U5320 (N_5320,N_4901,N_4509);
and U5321 (N_5321,N_4849,N_4872);
nor U5322 (N_5322,N_4746,N_4963);
nor U5323 (N_5323,N_4964,N_4947);
nand U5324 (N_5324,N_4906,N_4754);
xor U5325 (N_5325,N_4831,N_4887);
nand U5326 (N_5326,N_4564,N_4928);
or U5327 (N_5327,N_4660,N_4887);
and U5328 (N_5328,N_4980,N_4922);
nor U5329 (N_5329,N_4953,N_4569);
and U5330 (N_5330,N_4726,N_4603);
and U5331 (N_5331,N_4614,N_4763);
xnor U5332 (N_5332,N_4947,N_4881);
and U5333 (N_5333,N_4799,N_4597);
nand U5334 (N_5334,N_4770,N_4729);
and U5335 (N_5335,N_4985,N_4976);
nand U5336 (N_5336,N_4582,N_4681);
nand U5337 (N_5337,N_4855,N_4784);
and U5338 (N_5338,N_4767,N_4702);
and U5339 (N_5339,N_4752,N_4996);
and U5340 (N_5340,N_4600,N_4543);
and U5341 (N_5341,N_4726,N_4764);
and U5342 (N_5342,N_4861,N_4849);
and U5343 (N_5343,N_4733,N_4694);
nor U5344 (N_5344,N_4740,N_4512);
and U5345 (N_5345,N_4661,N_4514);
and U5346 (N_5346,N_4512,N_4834);
or U5347 (N_5347,N_4943,N_4657);
nor U5348 (N_5348,N_4659,N_4845);
and U5349 (N_5349,N_4856,N_4529);
or U5350 (N_5350,N_4933,N_4628);
nand U5351 (N_5351,N_4647,N_4507);
and U5352 (N_5352,N_4580,N_4978);
or U5353 (N_5353,N_4583,N_4723);
or U5354 (N_5354,N_4747,N_4783);
nor U5355 (N_5355,N_4574,N_4865);
and U5356 (N_5356,N_4694,N_4572);
nor U5357 (N_5357,N_4609,N_4731);
nor U5358 (N_5358,N_4563,N_4938);
nor U5359 (N_5359,N_4911,N_4549);
or U5360 (N_5360,N_4983,N_4990);
nand U5361 (N_5361,N_4964,N_4781);
or U5362 (N_5362,N_4972,N_4818);
nand U5363 (N_5363,N_4896,N_4870);
and U5364 (N_5364,N_4734,N_4939);
and U5365 (N_5365,N_4620,N_4584);
and U5366 (N_5366,N_4843,N_4545);
nor U5367 (N_5367,N_4706,N_4821);
xnor U5368 (N_5368,N_4604,N_4778);
nand U5369 (N_5369,N_4615,N_4913);
nor U5370 (N_5370,N_4675,N_4607);
nor U5371 (N_5371,N_4953,N_4531);
or U5372 (N_5372,N_4726,N_4790);
nand U5373 (N_5373,N_4788,N_4995);
nand U5374 (N_5374,N_4844,N_4591);
nor U5375 (N_5375,N_4918,N_4560);
or U5376 (N_5376,N_4734,N_4949);
nand U5377 (N_5377,N_4996,N_4784);
and U5378 (N_5378,N_4963,N_4670);
or U5379 (N_5379,N_4986,N_4597);
or U5380 (N_5380,N_4630,N_4514);
nor U5381 (N_5381,N_4711,N_4907);
nor U5382 (N_5382,N_4527,N_4630);
nand U5383 (N_5383,N_4764,N_4635);
xnor U5384 (N_5384,N_4741,N_4531);
nand U5385 (N_5385,N_4500,N_4984);
or U5386 (N_5386,N_4907,N_4703);
nand U5387 (N_5387,N_4623,N_4505);
nand U5388 (N_5388,N_4963,N_4855);
and U5389 (N_5389,N_4642,N_4960);
nand U5390 (N_5390,N_4976,N_4796);
nor U5391 (N_5391,N_4930,N_4847);
or U5392 (N_5392,N_4943,N_4542);
and U5393 (N_5393,N_4981,N_4600);
or U5394 (N_5394,N_4888,N_4731);
nand U5395 (N_5395,N_4850,N_4616);
nand U5396 (N_5396,N_4531,N_4942);
or U5397 (N_5397,N_4638,N_4772);
and U5398 (N_5398,N_4683,N_4746);
and U5399 (N_5399,N_4656,N_4981);
nor U5400 (N_5400,N_4907,N_4875);
or U5401 (N_5401,N_4509,N_4531);
or U5402 (N_5402,N_4587,N_4971);
or U5403 (N_5403,N_4521,N_4896);
nand U5404 (N_5404,N_4698,N_4932);
nand U5405 (N_5405,N_4675,N_4760);
and U5406 (N_5406,N_4944,N_4604);
nor U5407 (N_5407,N_4827,N_4746);
nor U5408 (N_5408,N_4735,N_4883);
nand U5409 (N_5409,N_4698,N_4911);
and U5410 (N_5410,N_4545,N_4711);
or U5411 (N_5411,N_4967,N_4689);
nand U5412 (N_5412,N_4742,N_4871);
and U5413 (N_5413,N_4840,N_4825);
nand U5414 (N_5414,N_4895,N_4788);
nor U5415 (N_5415,N_4719,N_4532);
nor U5416 (N_5416,N_4939,N_4526);
xnor U5417 (N_5417,N_4585,N_4911);
or U5418 (N_5418,N_4649,N_4926);
and U5419 (N_5419,N_4639,N_4842);
nor U5420 (N_5420,N_4553,N_4985);
and U5421 (N_5421,N_4771,N_4896);
nand U5422 (N_5422,N_4861,N_4531);
nand U5423 (N_5423,N_4546,N_4886);
or U5424 (N_5424,N_4868,N_4972);
nand U5425 (N_5425,N_4582,N_4712);
and U5426 (N_5426,N_4921,N_4667);
and U5427 (N_5427,N_4971,N_4860);
or U5428 (N_5428,N_4941,N_4762);
and U5429 (N_5429,N_4588,N_4604);
nor U5430 (N_5430,N_4704,N_4606);
and U5431 (N_5431,N_4524,N_4534);
nor U5432 (N_5432,N_4680,N_4575);
nor U5433 (N_5433,N_4594,N_4826);
nand U5434 (N_5434,N_4737,N_4692);
or U5435 (N_5435,N_4819,N_4536);
and U5436 (N_5436,N_4776,N_4940);
xor U5437 (N_5437,N_4873,N_4615);
nand U5438 (N_5438,N_4841,N_4731);
or U5439 (N_5439,N_4724,N_4568);
or U5440 (N_5440,N_4635,N_4842);
nor U5441 (N_5441,N_4854,N_4980);
nor U5442 (N_5442,N_4867,N_4511);
nor U5443 (N_5443,N_4707,N_4995);
or U5444 (N_5444,N_4788,N_4771);
or U5445 (N_5445,N_4972,N_4862);
xor U5446 (N_5446,N_4559,N_4613);
nand U5447 (N_5447,N_4865,N_4640);
or U5448 (N_5448,N_4777,N_4529);
and U5449 (N_5449,N_4618,N_4934);
nand U5450 (N_5450,N_4915,N_4997);
nand U5451 (N_5451,N_4761,N_4995);
and U5452 (N_5452,N_4841,N_4758);
or U5453 (N_5453,N_4932,N_4575);
nand U5454 (N_5454,N_4760,N_4672);
or U5455 (N_5455,N_4640,N_4889);
nand U5456 (N_5456,N_4628,N_4766);
nor U5457 (N_5457,N_4868,N_4635);
nand U5458 (N_5458,N_4768,N_4837);
and U5459 (N_5459,N_4504,N_4900);
and U5460 (N_5460,N_4726,N_4743);
nor U5461 (N_5461,N_4905,N_4606);
or U5462 (N_5462,N_4976,N_4721);
or U5463 (N_5463,N_4722,N_4900);
or U5464 (N_5464,N_4747,N_4979);
nand U5465 (N_5465,N_4664,N_4816);
or U5466 (N_5466,N_4918,N_4962);
nor U5467 (N_5467,N_4559,N_4793);
xnor U5468 (N_5468,N_4722,N_4964);
xnor U5469 (N_5469,N_4891,N_4682);
and U5470 (N_5470,N_4907,N_4819);
nand U5471 (N_5471,N_4565,N_4609);
and U5472 (N_5472,N_4946,N_4629);
or U5473 (N_5473,N_4951,N_4505);
and U5474 (N_5474,N_4611,N_4533);
nor U5475 (N_5475,N_4850,N_4660);
nand U5476 (N_5476,N_4513,N_4780);
xnor U5477 (N_5477,N_4753,N_4986);
and U5478 (N_5478,N_4507,N_4768);
and U5479 (N_5479,N_4830,N_4622);
or U5480 (N_5480,N_4822,N_4915);
nor U5481 (N_5481,N_4704,N_4738);
and U5482 (N_5482,N_4503,N_4610);
nor U5483 (N_5483,N_4733,N_4569);
nand U5484 (N_5484,N_4674,N_4573);
or U5485 (N_5485,N_4859,N_4526);
or U5486 (N_5486,N_4920,N_4507);
and U5487 (N_5487,N_4996,N_4766);
and U5488 (N_5488,N_4715,N_4604);
nor U5489 (N_5489,N_4793,N_4769);
nand U5490 (N_5490,N_4816,N_4575);
nand U5491 (N_5491,N_4785,N_4556);
nor U5492 (N_5492,N_4586,N_4895);
nor U5493 (N_5493,N_4641,N_4636);
xor U5494 (N_5494,N_4866,N_4605);
or U5495 (N_5495,N_4779,N_4856);
xor U5496 (N_5496,N_4801,N_4930);
nor U5497 (N_5497,N_4631,N_4526);
nor U5498 (N_5498,N_4915,N_4643);
nor U5499 (N_5499,N_4837,N_4588);
and U5500 (N_5500,N_5312,N_5152);
nand U5501 (N_5501,N_5403,N_5012);
or U5502 (N_5502,N_5347,N_5172);
nor U5503 (N_5503,N_5186,N_5179);
nor U5504 (N_5504,N_5359,N_5193);
nand U5505 (N_5505,N_5252,N_5076);
nor U5506 (N_5506,N_5308,N_5204);
nor U5507 (N_5507,N_5345,N_5091);
xnor U5508 (N_5508,N_5483,N_5142);
nor U5509 (N_5509,N_5155,N_5380);
and U5510 (N_5510,N_5078,N_5070);
nor U5511 (N_5511,N_5349,N_5048);
or U5512 (N_5512,N_5210,N_5052);
nand U5513 (N_5513,N_5125,N_5280);
xor U5514 (N_5514,N_5230,N_5087);
xnor U5515 (N_5515,N_5283,N_5160);
or U5516 (N_5516,N_5148,N_5336);
nor U5517 (N_5517,N_5479,N_5004);
nand U5518 (N_5518,N_5493,N_5121);
nand U5519 (N_5519,N_5399,N_5426);
and U5520 (N_5520,N_5147,N_5188);
nand U5521 (N_5521,N_5183,N_5221);
xnor U5522 (N_5522,N_5450,N_5243);
or U5523 (N_5523,N_5309,N_5303);
nand U5524 (N_5524,N_5397,N_5433);
xor U5525 (N_5525,N_5151,N_5115);
nor U5526 (N_5526,N_5126,N_5153);
or U5527 (N_5527,N_5042,N_5306);
nor U5528 (N_5528,N_5063,N_5109);
or U5529 (N_5529,N_5476,N_5353);
and U5530 (N_5530,N_5366,N_5299);
or U5531 (N_5531,N_5202,N_5059);
or U5532 (N_5532,N_5326,N_5377);
and U5533 (N_5533,N_5339,N_5219);
nand U5534 (N_5534,N_5488,N_5460);
or U5535 (N_5535,N_5143,N_5010);
nor U5536 (N_5536,N_5196,N_5064);
or U5537 (N_5537,N_5024,N_5105);
and U5538 (N_5538,N_5164,N_5051);
nand U5539 (N_5539,N_5067,N_5328);
or U5540 (N_5540,N_5400,N_5365);
and U5541 (N_5541,N_5368,N_5350);
nor U5542 (N_5542,N_5469,N_5200);
nor U5543 (N_5543,N_5158,N_5225);
or U5544 (N_5544,N_5390,N_5173);
or U5545 (N_5545,N_5319,N_5298);
nor U5546 (N_5546,N_5244,N_5223);
and U5547 (N_5547,N_5373,N_5285);
nor U5548 (N_5548,N_5075,N_5360);
nor U5549 (N_5549,N_5335,N_5379);
and U5550 (N_5550,N_5232,N_5402);
nor U5551 (N_5551,N_5393,N_5028);
nor U5552 (N_5552,N_5013,N_5464);
nor U5553 (N_5553,N_5430,N_5136);
or U5554 (N_5554,N_5275,N_5383);
or U5555 (N_5555,N_5362,N_5199);
nor U5556 (N_5556,N_5346,N_5082);
or U5557 (N_5557,N_5321,N_5094);
nor U5558 (N_5558,N_5046,N_5036);
xnor U5559 (N_5559,N_5029,N_5089);
and U5560 (N_5560,N_5385,N_5388);
and U5561 (N_5561,N_5408,N_5043);
and U5562 (N_5562,N_5103,N_5412);
and U5563 (N_5563,N_5175,N_5241);
and U5564 (N_5564,N_5471,N_5058);
nand U5565 (N_5565,N_5263,N_5442);
nand U5566 (N_5566,N_5047,N_5418);
nand U5567 (N_5567,N_5435,N_5170);
and U5568 (N_5568,N_5340,N_5239);
and U5569 (N_5569,N_5293,N_5135);
nand U5570 (N_5570,N_5203,N_5287);
or U5571 (N_5571,N_5166,N_5157);
nor U5572 (N_5572,N_5086,N_5330);
nor U5573 (N_5573,N_5182,N_5258);
and U5574 (N_5574,N_5332,N_5007);
nand U5575 (N_5575,N_5327,N_5267);
or U5576 (N_5576,N_5236,N_5238);
and U5577 (N_5577,N_5456,N_5113);
and U5578 (N_5578,N_5361,N_5475);
nand U5579 (N_5579,N_5249,N_5116);
xor U5580 (N_5580,N_5057,N_5008);
or U5581 (N_5581,N_5448,N_5144);
and U5582 (N_5582,N_5382,N_5304);
nand U5583 (N_5583,N_5259,N_5101);
and U5584 (N_5584,N_5296,N_5229);
nor U5585 (N_5585,N_5331,N_5441);
xor U5586 (N_5586,N_5053,N_5127);
or U5587 (N_5587,N_5455,N_5465);
nor U5588 (N_5588,N_5001,N_5311);
nand U5589 (N_5589,N_5484,N_5378);
nand U5590 (N_5590,N_5478,N_5301);
or U5591 (N_5591,N_5463,N_5054);
or U5592 (N_5592,N_5141,N_5253);
xnor U5593 (N_5593,N_5364,N_5178);
nor U5594 (N_5594,N_5080,N_5461);
nor U5595 (N_5595,N_5201,N_5401);
nor U5596 (N_5596,N_5088,N_5074);
and U5597 (N_5597,N_5235,N_5256);
nor U5598 (N_5598,N_5176,N_5406);
and U5599 (N_5599,N_5357,N_5137);
and U5600 (N_5600,N_5477,N_5133);
or U5601 (N_5601,N_5495,N_5034);
or U5602 (N_5602,N_5485,N_5363);
or U5603 (N_5603,N_5003,N_5209);
or U5604 (N_5604,N_5065,N_5445);
and U5605 (N_5605,N_5324,N_5061);
and U5606 (N_5606,N_5040,N_5458);
nand U5607 (N_5607,N_5104,N_5092);
or U5608 (N_5608,N_5315,N_5352);
nand U5609 (N_5609,N_5146,N_5023);
or U5610 (N_5610,N_5006,N_5314);
or U5611 (N_5611,N_5279,N_5468);
or U5612 (N_5612,N_5019,N_5031);
nand U5613 (N_5613,N_5389,N_5169);
nand U5614 (N_5614,N_5261,N_5248);
nor U5615 (N_5615,N_5318,N_5413);
or U5616 (N_5616,N_5457,N_5404);
and U5617 (N_5617,N_5228,N_5174);
nand U5618 (N_5618,N_5274,N_5271);
or U5619 (N_5619,N_5420,N_5452);
nand U5620 (N_5620,N_5185,N_5369);
or U5621 (N_5621,N_5022,N_5180);
or U5622 (N_5622,N_5156,N_5437);
and U5623 (N_5623,N_5292,N_5260);
and U5624 (N_5624,N_5112,N_5251);
and U5625 (N_5625,N_5351,N_5424);
or U5626 (N_5626,N_5071,N_5095);
or U5627 (N_5627,N_5073,N_5313);
nor U5628 (N_5628,N_5356,N_5438);
nand U5629 (N_5629,N_5436,N_5497);
nand U5630 (N_5630,N_5338,N_5494);
nand U5631 (N_5631,N_5425,N_5474);
nor U5632 (N_5632,N_5079,N_5462);
and U5633 (N_5633,N_5191,N_5100);
or U5634 (N_5634,N_5149,N_5282);
and U5635 (N_5635,N_5415,N_5419);
nor U5636 (N_5636,N_5120,N_5454);
and U5637 (N_5637,N_5168,N_5014);
nand U5638 (N_5638,N_5165,N_5266);
nand U5639 (N_5639,N_5325,N_5190);
and U5640 (N_5640,N_5355,N_5097);
nor U5641 (N_5641,N_5123,N_5410);
nand U5642 (N_5642,N_5288,N_5090);
and U5643 (N_5643,N_5498,N_5333);
nor U5644 (N_5644,N_5145,N_5265);
nand U5645 (N_5645,N_5015,N_5220);
nor U5646 (N_5646,N_5446,N_5026);
nand U5647 (N_5647,N_5119,N_5247);
and U5648 (N_5648,N_5214,N_5081);
and U5649 (N_5649,N_5222,N_5354);
xor U5650 (N_5650,N_5320,N_5375);
or U5651 (N_5651,N_5310,N_5035);
nand U5652 (N_5652,N_5434,N_5421);
nor U5653 (N_5653,N_5056,N_5177);
nand U5654 (N_5654,N_5187,N_5384);
or U5655 (N_5655,N_5163,N_5374);
nand U5656 (N_5656,N_5020,N_5207);
or U5657 (N_5657,N_5297,N_5205);
or U5658 (N_5658,N_5124,N_5428);
nand U5659 (N_5659,N_5482,N_5416);
nand U5660 (N_5660,N_5440,N_5499);
nor U5661 (N_5661,N_5041,N_5481);
or U5662 (N_5662,N_5489,N_5050);
xnor U5663 (N_5663,N_5030,N_5262);
nand U5664 (N_5664,N_5106,N_5432);
or U5665 (N_5665,N_5411,N_5009);
and U5666 (N_5666,N_5044,N_5281);
nand U5667 (N_5667,N_5197,N_5150);
nand U5668 (N_5668,N_5102,N_5302);
and U5669 (N_5669,N_5341,N_5409);
and U5670 (N_5670,N_5117,N_5130);
nand U5671 (N_5671,N_5154,N_5367);
nor U5672 (N_5672,N_5138,N_5140);
nand U5673 (N_5673,N_5002,N_5194);
xnor U5674 (N_5674,N_5118,N_5017);
xor U5675 (N_5675,N_5417,N_5322);
nor U5676 (N_5676,N_5184,N_5069);
and U5677 (N_5677,N_5427,N_5496);
nor U5678 (N_5678,N_5439,N_5342);
and U5679 (N_5679,N_5268,N_5348);
nand U5680 (N_5680,N_5470,N_5277);
or U5681 (N_5681,N_5407,N_5038);
and U5682 (N_5682,N_5198,N_5237);
or U5683 (N_5683,N_5216,N_5396);
or U5684 (N_5684,N_5316,N_5161);
or U5685 (N_5685,N_5334,N_5429);
and U5686 (N_5686,N_5084,N_5344);
and U5687 (N_5687,N_5016,N_5284);
and U5688 (N_5688,N_5264,N_5307);
nand U5689 (N_5689,N_5449,N_5467);
or U5690 (N_5690,N_5025,N_5005);
or U5691 (N_5691,N_5234,N_5018);
and U5692 (N_5692,N_5289,N_5276);
or U5693 (N_5693,N_5391,N_5211);
or U5694 (N_5694,N_5139,N_5111);
nand U5695 (N_5695,N_5134,N_5394);
and U5696 (N_5696,N_5066,N_5000);
nor U5697 (N_5697,N_5011,N_5195);
nand U5698 (N_5698,N_5098,N_5110);
or U5699 (N_5699,N_5294,N_5215);
or U5700 (N_5700,N_5077,N_5192);
nand U5701 (N_5701,N_5181,N_5386);
or U5702 (N_5702,N_5398,N_5358);
or U5703 (N_5703,N_5093,N_5208);
nand U5704 (N_5704,N_5206,N_5453);
or U5705 (N_5705,N_5226,N_5227);
nor U5706 (N_5706,N_5131,N_5387);
xnor U5707 (N_5707,N_5395,N_5122);
nor U5708 (N_5708,N_5422,N_5107);
or U5709 (N_5709,N_5159,N_5272);
nand U5710 (N_5710,N_5278,N_5250);
and U5711 (N_5711,N_5245,N_5300);
and U5712 (N_5712,N_5049,N_5062);
nand U5713 (N_5713,N_5473,N_5459);
and U5714 (N_5714,N_5083,N_5337);
and U5715 (N_5715,N_5217,N_5242);
or U5716 (N_5716,N_5128,N_5370);
nand U5717 (N_5717,N_5212,N_5027);
and U5718 (N_5718,N_5305,N_5343);
nand U5719 (N_5719,N_5213,N_5405);
or U5720 (N_5720,N_5273,N_5376);
and U5721 (N_5721,N_5045,N_5329);
or U5722 (N_5722,N_5466,N_5269);
nand U5723 (N_5723,N_5491,N_5257);
nand U5724 (N_5724,N_5381,N_5037);
and U5725 (N_5725,N_5096,N_5431);
nand U5726 (N_5726,N_5392,N_5189);
nor U5727 (N_5727,N_5423,N_5295);
nor U5728 (N_5728,N_5317,N_5480);
and U5729 (N_5729,N_5444,N_5039);
nor U5730 (N_5730,N_5255,N_5487);
or U5731 (N_5731,N_5447,N_5224);
nand U5732 (N_5732,N_5231,N_5218);
nor U5733 (N_5733,N_5171,N_5486);
nor U5734 (N_5734,N_5414,N_5472);
or U5735 (N_5735,N_5372,N_5068);
and U5736 (N_5736,N_5032,N_5033);
or U5737 (N_5737,N_5114,N_5290);
nand U5738 (N_5738,N_5286,N_5099);
and U5739 (N_5739,N_5129,N_5291);
nand U5740 (N_5740,N_5108,N_5167);
or U5741 (N_5741,N_5162,N_5085);
nand U5742 (N_5742,N_5254,N_5240);
nor U5743 (N_5743,N_5055,N_5323);
nand U5744 (N_5744,N_5021,N_5270);
nor U5745 (N_5745,N_5132,N_5443);
or U5746 (N_5746,N_5371,N_5060);
and U5747 (N_5747,N_5246,N_5451);
and U5748 (N_5748,N_5492,N_5233);
or U5749 (N_5749,N_5072,N_5490);
nor U5750 (N_5750,N_5043,N_5087);
nor U5751 (N_5751,N_5188,N_5177);
and U5752 (N_5752,N_5135,N_5297);
nor U5753 (N_5753,N_5258,N_5139);
nand U5754 (N_5754,N_5449,N_5261);
or U5755 (N_5755,N_5384,N_5260);
nand U5756 (N_5756,N_5101,N_5126);
nor U5757 (N_5757,N_5193,N_5333);
or U5758 (N_5758,N_5365,N_5341);
nor U5759 (N_5759,N_5067,N_5317);
and U5760 (N_5760,N_5267,N_5439);
or U5761 (N_5761,N_5112,N_5066);
or U5762 (N_5762,N_5351,N_5158);
nor U5763 (N_5763,N_5211,N_5478);
or U5764 (N_5764,N_5403,N_5120);
or U5765 (N_5765,N_5169,N_5179);
and U5766 (N_5766,N_5327,N_5094);
and U5767 (N_5767,N_5255,N_5018);
or U5768 (N_5768,N_5298,N_5383);
xor U5769 (N_5769,N_5057,N_5069);
or U5770 (N_5770,N_5030,N_5210);
or U5771 (N_5771,N_5177,N_5099);
nand U5772 (N_5772,N_5166,N_5168);
and U5773 (N_5773,N_5006,N_5466);
or U5774 (N_5774,N_5208,N_5013);
or U5775 (N_5775,N_5349,N_5181);
nand U5776 (N_5776,N_5273,N_5421);
or U5777 (N_5777,N_5109,N_5307);
nor U5778 (N_5778,N_5444,N_5118);
nor U5779 (N_5779,N_5292,N_5295);
xor U5780 (N_5780,N_5320,N_5381);
or U5781 (N_5781,N_5150,N_5001);
xnor U5782 (N_5782,N_5042,N_5156);
nor U5783 (N_5783,N_5105,N_5279);
and U5784 (N_5784,N_5433,N_5011);
and U5785 (N_5785,N_5355,N_5462);
or U5786 (N_5786,N_5449,N_5337);
and U5787 (N_5787,N_5434,N_5432);
or U5788 (N_5788,N_5176,N_5389);
and U5789 (N_5789,N_5055,N_5337);
nor U5790 (N_5790,N_5236,N_5151);
nor U5791 (N_5791,N_5205,N_5097);
and U5792 (N_5792,N_5193,N_5136);
nor U5793 (N_5793,N_5267,N_5241);
nand U5794 (N_5794,N_5436,N_5098);
nor U5795 (N_5795,N_5439,N_5290);
nor U5796 (N_5796,N_5416,N_5248);
nand U5797 (N_5797,N_5263,N_5465);
or U5798 (N_5798,N_5086,N_5476);
and U5799 (N_5799,N_5347,N_5158);
and U5800 (N_5800,N_5341,N_5479);
and U5801 (N_5801,N_5200,N_5029);
nand U5802 (N_5802,N_5204,N_5318);
nand U5803 (N_5803,N_5489,N_5444);
or U5804 (N_5804,N_5488,N_5192);
nor U5805 (N_5805,N_5396,N_5226);
and U5806 (N_5806,N_5354,N_5453);
and U5807 (N_5807,N_5383,N_5032);
xor U5808 (N_5808,N_5173,N_5441);
and U5809 (N_5809,N_5310,N_5181);
nor U5810 (N_5810,N_5098,N_5439);
or U5811 (N_5811,N_5166,N_5454);
nor U5812 (N_5812,N_5164,N_5129);
and U5813 (N_5813,N_5149,N_5473);
and U5814 (N_5814,N_5139,N_5227);
nor U5815 (N_5815,N_5059,N_5216);
or U5816 (N_5816,N_5106,N_5488);
and U5817 (N_5817,N_5468,N_5063);
and U5818 (N_5818,N_5141,N_5359);
or U5819 (N_5819,N_5159,N_5001);
nand U5820 (N_5820,N_5272,N_5444);
and U5821 (N_5821,N_5478,N_5142);
and U5822 (N_5822,N_5281,N_5013);
or U5823 (N_5823,N_5307,N_5363);
and U5824 (N_5824,N_5398,N_5001);
or U5825 (N_5825,N_5102,N_5451);
nand U5826 (N_5826,N_5328,N_5357);
nor U5827 (N_5827,N_5420,N_5011);
nand U5828 (N_5828,N_5129,N_5151);
nor U5829 (N_5829,N_5458,N_5271);
nand U5830 (N_5830,N_5146,N_5442);
nand U5831 (N_5831,N_5278,N_5431);
nand U5832 (N_5832,N_5041,N_5280);
and U5833 (N_5833,N_5081,N_5227);
and U5834 (N_5834,N_5136,N_5257);
and U5835 (N_5835,N_5481,N_5387);
and U5836 (N_5836,N_5224,N_5208);
xnor U5837 (N_5837,N_5219,N_5174);
nor U5838 (N_5838,N_5214,N_5245);
nand U5839 (N_5839,N_5244,N_5136);
or U5840 (N_5840,N_5364,N_5275);
nor U5841 (N_5841,N_5024,N_5092);
and U5842 (N_5842,N_5084,N_5266);
and U5843 (N_5843,N_5236,N_5369);
nor U5844 (N_5844,N_5217,N_5151);
xnor U5845 (N_5845,N_5496,N_5438);
and U5846 (N_5846,N_5414,N_5416);
or U5847 (N_5847,N_5219,N_5464);
or U5848 (N_5848,N_5066,N_5281);
and U5849 (N_5849,N_5144,N_5299);
and U5850 (N_5850,N_5242,N_5065);
nand U5851 (N_5851,N_5339,N_5264);
or U5852 (N_5852,N_5441,N_5218);
xnor U5853 (N_5853,N_5177,N_5290);
or U5854 (N_5854,N_5279,N_5073);
nand U5855 (N_5855,N_5469,N_5055);
or U5856 (N_5856,N_5096,N_5390);
nand U5857 (N_5857,N_5320,N_5102);
or U5858 (N_5858,N_5481,N_5407);
nor U5859 (N_5859,N_5290,N_5056);
nor U5860 (N_5860,N_5036,N_5317);
nand U5861 (N_5861,N_5463,N_5379);
nand U5862 (N_5862,N_5397,N_5104);
and U5863 (N_5863,N_5341,N_5020);
nor U5864 (N_5864,N_5322,N_5447);
and U5865 (N_5865,N_5097,N_5260);
nand U5866 (N_5866,N_5315,N_5089);
or U5867 (N_5867,N_5128,N_5217);
or U5868 (N_5868,N_5295,N_5486);
nand U5869 (N_5869,N_5286,N_5235);
nand U5870 (N_5870,N_5152,N_5446);
nor U5871 (N_5871,N_5102,N_5420);
or U5872 (N_5872,N_5442,N_5089);
xnor U5873 (N_5873,N_5110,N_5362);
and U5874 (N_5874,N_5258,N_5494);
nand U5875 (N_5875,N_5326,N_5246);
nor U5876 (N_5876,N_5449,N_5387);
and U5877 (N_5877,N_5410,N_5304);
nor U5878 (N_5878,N_5195,N_5430);
nand U5879 (N_5879,N_5294,N_5097);
and U5880 (N_5880,N_5151,N_5293);
and U5881 (N_5881,N_5464,N_5107);
or U5882 (N_5882,N_5188,N_5070);
or U5883 (N_5883,N_5313,N_5049);
nor U5884 (N_5884,N_5323,N_5239);
nor U5885 (N_5885,N_5305,N_5189);
nor U5886 (N_5886,N_5135,N_5189);
nand U5887 (N_5887,N_5429,N_5395);
nand U5888 (N_5888,N_5131,N_5403);
and U5889 (N_5889,N_5090,N_5015);
nand U5890 (N_5890,N_5071,N_5454);
nand U5891 (N_5891,N_5086,N_5265);
nor U5892 (N_5892,N_5312,N_5176);
nor U5893 (N_5893,N_5020,N_5150);
and U5894 (N_5894,N_5149,N_5243);
or U5895 (N_5895,N_5496,N_5383);
or U5896 (N_5896,N_5251,N_5344);
nor U5897 (N_5897,N_5033,N_5044);
or U5898 (N_5898,N_5301,N_5057);
xnor U5899 (N_5899,N_5092,N_5476);
nand U5900 (N_5900,N_5442,N_5105);
or U5901 (N_5901,N_5047,N_5125);
nand U5902 (N_5902,N_5105,N_5047);
nor U5903 (N_5903,N_5285,N_5046);
nor U5904 (N_5904,N_5010,N_5322);
or U5905 (N_5905,N_5407,N_5360);
or U5906 (N_5906,N_5127,N_5132);
nand U5907 (N_5907,N_5006,N_5385);
nor U5908 (N_5908,N_5108,N_5068);
nand U5909 (N_5909,N_5094,N_5420);
and U5910 (N_5910,N_5175,N_5422);
and U5911 (N_5911,N_5008,N_5115);
and U5912 (N_5912,N_5034,N_5131);
or U5913 (N_5913,N_5496,N_5166);
and U5914 (N_5914,N_5397,N_5193);
or U5915 (N_5915,N_5159,N_5362);
nand U5916 (N_5916,N_5434,N_5244);
nor U5917 (N_5917,N_5137,N_5170);
nor U5918 (N_5918,N_5039,N_5455);
nor U5919 (N_5919,N_5492,N_5208);
nand U5920 (N_5920,N_5262,N_5297);
nand U5921 (N_5921,N_5403,N_5031);
nand U5922 (N_5922,N_5069,N_5225);
or U5923 (N_5923,N_5242,N_5223);
nor U5924 (N_5924,N_5255,N_5269);
or U5925 (N_5925,N_5212,N_5047);
and U5926 (N_5926,N_5420,N_5249);
nor U5927 (N_5927,N_5398,N_5037);
nand U5928 (N_5928,N_5343,N_5468);
or U5929 (N_5929,N_5196,N_5170);
and U5930 (N_5930,N_5327,N_5151);
nor U5931 (N_5931,N_5332,N_5221);
and U5932 (N_5932,N_5052,N_5346);
and U5933 (N_5933,N_5218,N_5168);
nor U5934 (N_5934,N_5139,N_5256);
nand U5935 (N_5935,N_5070,N_5450);
nor U5936 (N_5936,N_5123,N_5274);
nor U5937 (N_5937,N_5487,N_5278);
nor U5938 (N_5938,N_5417,N_5267);
nand U5939 (N_5939,N_5075,N_5451);
nand U5940 (N_5940,N_5483,N_5117);
nand U5941 (N_5941,N_5261,N_5137);
and U5942 (N_5942,N_5381,N_5011);
and U5943 (N_5943,N_5218,N_5313);
or U5944 (N_5944,N_5490,N_5433);
nand U5945 (N_5945,N_5180,N_5120);
nor U5946 (N_5946,N_5225,N_5360);
nand U5947 (N_5947,N_5292,N_5090);
nor U5948 (N_5948,N_5485,N_5208);
nand U5949 (N_5949,N_5096,N_5373);
nor U5950 (N_5950,N_5477,N_5333);
nor U5951 (N_5951,N_5456,N_5224);
nor U5952 (N_5952,N_5295,N_5358);
or U5953 (N_5953,N_5430,N_5125);
and U5954 (N_5954,N_5491,N_5206);
and U5955 (N_5955,N_5351,N_5394);
and U5956 (N_5956,N_5205,N_5405);
and U5957 (N_5957,N_5107,N_5280);
nand U5958 (N_5958,N_5114,N_5247);
nor U5959 (N_5959,N_5033,N_5481);
and U5960 (N_5960,N_5156,N_5409);
nand U5961 (N_5961,N_5042,N_5000);
nand U5962 (N_5962,N_5461,N_5287);
nand U5963 (N_5963,N_5109,N_5035);
and U5964 (N_5964,N_5083,N_5243);
or U5965 (N_5965,N_5348,N_5297);
nor U5966 (N_5966,N_5109,N_5163);
nor U5967 (N_5967,N_5004,N_5289);
nor U5968 (N_5968,N_5246,N_5317);
nor U5969 (N_5969,N_5402,N_5014);
or U5970 (N_5970,N_5109,N_5123);
or U5971 (N_5971,N_5483,N_5305);
and U5972 (N_5972,N_5480,N_5177);
nor U5973 (N_5973,N_5176,N_5330);
nor U5974 (N_5974,N_5417,N_5490);
nor U5975 (N_5975,N_5318,N_5309);
and U5976 (N_5976,N_5092,N_5046);
and U5977 (N_5977,N_5037,N_5129);
and U5978 (N_5978,N_5074,N_5211);
nand U5979 (N_5979,N_5427,N_5441);
or U5980 (N_5980,N_5360,N_5371);
and U5981 (N_5981,N_5163,N_5148);
and U5982 (N_5982,N_5171,N_5261);
nor U5983 (N_5983,N_5249,N_5082);
nor U5984 (N_5984,N_5339,N_5420);
or U5985 (N_5985,N_5346,N_5471);
nor U5986 (N_5986,N_5278,N_5287);
nand U5987 (N_5987,N_5030,N_5122);
xor U5988 (N_5988,N_5212,N_5101);
nor U5989 (N_5989,N_5428,N_5152);
and U5990 (N_5990,N_5267,N_5057);
nand U5991 (N_5991,N_5233,N_5290);
nand U5992 (N_5992,N_5478,N_5423);
or U5993 (N_5993,N_5392,N_5096);
or U5994 (N_5994,N_5389,N_5186);
nor U5995 (N_5995,N_5081,N_5156);
nor U5996 (N_5996,N_5211,N_5397);
and U5997 (N_5997,N_5261,N_5281);
and U5998 (N_5998,N_5298,N_5309);
nand U5999 (N_5999,N_5343,N_5431);
or U6000 (N_6000,N_5806,N_5817);
or U6001 (N_6001,N_5826,N_5651);
or U6002 (N_6002,N_5699,N_5932);
or U6003 (N_6003,N_5884,N_5576);
nor U6004 (N_6004,N_5953,N_5694);
nand U6005 (N_6005,N_5773,N_5854);
nand U6006 (N_6006,N_5834,N_5527);
nor U6007 (N_6007,N_5794,N_5803);
and U6008 (N_6008,N_5838,N_5546);
or U6009 (N_6009,N_5606,N_5644);
nor U6010 (N_6010,N_5542,N_5859);
nand U6011 (N_6011,N_5610,N_5877);
nor U6012 (N_6012,N_5565,N_5825);
and U6013 (N_6013,N_5833,N_5870);
or U6014 (N_6014,N_5541,N_5663);
and U6015 (N_6015,N_5970,N_5689);
nor U6016 (N_6016,N_5521,N_5821);
nor U6017 (N_6017,N_5755,N_5731);
nor U6018 (N_6018,N_5963,N_5865);
or U6019 (N_6019,N_5635,N_5898);
or U6020 (N_6020,N_5510,N_5950);
nand U6021 (N_6021,N_5761,N_5904);
or U6022 (N_6022,N_5662,N_5553);
nand U6023 (N_6023,N_5743,N_5781);
nor U6024 (N_6024,N_5924,N_5560);
and U6025 (N_6025,N_5706,N_5780);
and U6026 (N_6026,N_5992,N_5595);
or U6027 (N_6027,N_5926,N_5547);
or U6028 (N_6028,N_5867,N_5664);
nor U6029 (N_6029,N_5738,N_5903);
and U6030 (N_6030,N_5646,N_5568);
nor U6031 (N_6031,N_5700,N_5899);
and U6032 (N_6032,N_5681,N_5976);
and U6033 (N_6033,N_5969,N_5787);
and U6034 (N_6034,N_5964,N_5954);
xor U6035 (N_6035,N_5863,N_5797);
nand U6036 (N_6036,N_5670,N_5557);
nand U6037 (N_6037,N_5637,N_5944);
nand U6038 (N_6038,N_5508,N_5989);
and U6039 (N_6039,N_5609,N_5686);
and U6040 (N_6040,N_5584,N_5840);
or U6041 (N_6041,N_5692,N_5878);
and U6042 (N_6042,N_5798,N_5575);
and U6043 (N_6043,N_5933,N_5939);
or U6044 (N_6044,N_5740,N_5795);
and U6045 (N_6045,N_5589,N_5974);
nor U6046 (N_6046,N_5608,N_5647);
or U6047 (N_6047,N_5828,N_5951);
or U6048 (N_6048,N_5843,N_5523);
xnor U6049 (N_6049,N_5571,N_5975);
and U6050 (N_6050,N_5791,N_5856);
or U6051 (N_6051,N_5894,N_5634);
or U6052 (N_6052,N_5650,N_5617);
or U6053 (N_6053,N_5759,N_5545);
and U6054 (N_6054,N_5813,N_5660);
or U6055 (N_6055,N_5580,N_5675);
nand U6056 (N_6056,N_5848,N_5752);
nand U6057 (N_6057,N_5912,N_5501);
nand U6058 (N_6058,N_5581,N_5889);
nor U6059 (N_6059,N_5996,N_5762);
and U6060 (N_6060,N_5629,N_5550);
and U6061 (N_6061,N_5613,N_5562);
xnor U6062 (N_6062,N_5707,N_5882);
and U6063 (N_6063,N_5742,N_5804);
and U6064 (N_6064,N_5881,N_5765);
and U6065 (N_6065,N_5980,N_5596);
nand U6066 (N_6066,N_5711,N_5533);
nor U6067 (N_6067,N_5793,N_5505);
or U6068 (N_6068,N_5966,N_5666);
nor U6069 (N_6069,N_5783,N_5910);
nor U6070 (N_6070,N_5535,N_5841);
or U6071 (N_6071,N_5516,N_5654);
and U6072 (N_6072,N_5993,N_5799);
or U6073 (N_6073,N_5927,N_5633);
and U6074 (N_6074,N_5582,N_5648);
and U6075 (N_6075,N_5973,N_5625);
or U6076 (N_6076,N_5957,N_5661);
nand U6077 (N_6077,N_5543,N_5921);
nand U6078 (N_6078,N_5754,N_5891);
or U6079 (N_6079,N_5688,N_5829);
nand U6080 (N_6080,N_5846,N_5880);
and U6081 (N_6081,N_5509,N_5757);
and U6082 (N_6082,N_5623,N_5929);
and U6083 (N_6083,N_5615,N_5522);
or U6084 (N_6084,N_5758,N_5790);
and U6085 (N_6085,N_5955,N_5869);
xnor U6086 (N_6086,N_5801,N_5500);
and U6087 (N_6087,N_5528,N_5655);
nand U6088 (N_6088,N_5671,N_5600);
and U6089 (N_6089,N_5937,N_5524);
and U6090 (N_6090,N_5721,N_5864);
nand U6091 (N_6091,N_5956,N_5642);
nor U6092 (N_6092,N_5786,N_5569);
xor U6093 (N_6093,N_5525,N_5777);
nor U6094 (N_6094,N_5529,N_5851);
nor U6095 (N_6095,N_5997,N_5552);
nand U6096 (N_6096,N_5872,N_5732);
nand U6097 (N_6097,N_5816,N_5747);
nand U6098 (N_6098,N_5815,N_5753);
and U6099 (N_6099,N_5638,N_5621);
or U6100 (N_6100,N_5632,N_5641);
and U6101 (N_6101,N_5734,N_5900);
nand U6102 (N_6102,N_5984,N_5897);
or U6103 (N_6103,N_5722,N_5824);
xor U6104 (N_6104,N_5696,N_5590);
nand U6105 (N_6105,N_5987,N_5549);
nor U6106 (N_6106,N_5946,N_5519);
and U6107 (N_6107,N_5728,N_5643);
nor U6108 (N_6108,N_5587,N_5938);
nor U6109 (N_6109,N_5611,N_5583);
and U6110 (N_6110,N_5756,N_5687);
nand U6111 (N_6111,N_5942,N_5701);
nor U6112 (N_6112,N_5916,N_5713);
nor U6113 (N_6113,N_5620,N_5673);
and U6114 (N_6114,N_5931,N_5985);
or U6115 (N_6115,N_5839,N_5923);
or U6116 (N_6116,N_5574,N_5888);
xnor U6117 (N_6117,N_5503,N_5855);
or U6118 (N_6118,N_5586,N_5695);
or U6119 (N_6119,N_5890,N_5750);
or U6120 (N_6120,N_5507,N_5626);
nand U6121 (N_6121,N_5934,N_5814);
and U6122 (N_6122,N_5925,N_5708);
nand U6123 (N_6123,N_5792,N_5809);
nor U6124 (N_6124,N_5896,N_5594);
or U6125 (N_6125,N_5979,N_5573);
or U6126 (N_6126,N_5918,N_5724);
nand U6127 (N_6127,N_5767,N_5674);
or U6128 (N_6128,N_5958,N_5669);
nand U6129 (N_6129,N_5748,N_5796);
nor U6130 (N_6130,N_5684,N_5567);
or U6131 (N_6131,N_5837,N_5668);
nand U6132 (N_6132,N_5819,N_5835);
nor U6133 (N_6133,N_5785,N_5538);
nand U6134 (N_6134,N_5778,N_5627);
nor U6135 (N_6135,N_5564,N_5920);
nor U6136 (N_6136,N_5591,N_5911);
nand U6137 (N_6137,N_5977,N_5892);
nor U6138 (N_6138,N_5725,N_5982);
and U6139 (N_6139,N_5531,N_5978);
nand U6140 (N_6140,N_5502,N_5810);
or U6141 (N_6141,N_5605,N_5685);
or U6142 (N_6142,N_5811,N_5842);
nor U6143 (N_6143,N_5619,N_5908);
and U6144 (N_6144,N_5727,N_5599);
or U6145 (N_6145,N_5802,N_5905);
and U6146 (N_6146,N_5733,N_5871);
or U6147 (N_6147,N_5769,N_5735);
nor U6148 (N_6148,N_5917,N_5990);
and U6149 (N_6149,N_5548,N_5639);
and U6150 (N_6150,N_5504,N_5818);
nor U6151 (N_6151,N_5913,N_5901);
and U6152 (N_6152,N_5554,N_5922);
and U6153 (N_6153,N_5822,N_5601);
nor U6154 (N_6154,N_5624,N_5879);
and U6155 (N_6155,N_5849,N_5857);
or U6156 (N_6156,N_5514,N_5534);
nand U6157 (N_6157,N_5719,N_5960);
nor U6158 (N_6158,N_5866,N_5526);
and U6159 (N_6159,N_5656,N_5506);
nand U6160 (N_6160,N_5775,N_5874);
and U6161 (N_6161,N_5572,N_5511);
and U6162 (N_6162,N_5709,N_5945);
nor U6163 (N_6163,N_5559,N_5789);
nand U6164 (N_6164,N_5537,N_5737);
and U6165 (N_6165,N_5820,N_5741);
or U6166 (N_6166,N_5860,N_5994);
or U6167 (N_6167,N_5805,N_5995);
nor U6168 (N_6168,N_5607,N_5578);
and U6169 (N_6169,N_5763,N_5784);
nor U6170 (N_6170,N_5652,N_5518);
or U6171 (N_6171,N_5850,N_5716);
nor U6172 (N_6172,N_5726,N_5530);
nor U6173 (N_6173,N_5788,N_5902);
nand U6174 (N_6174,N_5513,N_5614);
nand U6175 (N_6175,N_5693,N_5630);
nor U6176 (N_6176,N_5883,N_5736);
nor U6177 (N_6177,N_5680,N_5540);
nor U6178 (N_6178,N_5712,N_5679);
nor U6179 (N_6179,N_5965,N_5967);
and U6180 (N_6180,N_5986,N_5622);
nor U6181 (N_6181,N_5588,N_5603);
and U6182 (N_6182,N_5676,N_5555);
nand U6183 (N_6183,N_5909,N_5940);
nor U6184 (N_6184,N_5705,N_5585);
or U6185 (N_6185,N_5764,N_5710);
or U6186 (N_6186,N_5830,N_5919);
nand U6187 (N_6187,N_5928,N_5868);
or U6188 (N_6188,N_5690,N_5563);
nor U6189 (N_6189,N_5845,N_5715);
and U6190 (N_6190,N_5570,N_5847);
nand U6191 (N_6191,N_5703,N_5943);
nand U6192 (N_6192,N_5930,N_5906);
or U6193 (N_6193,N_5645,N_5640);
or U6194 (N_6194,N_5512,N_5593);
nand U6195 (N_6195,N_5592,N_5649);
or U6196 (N_6196,N_5730,N_5566);
nor U6197 (N_6197,N_5766,N_5771);
nand U6198 (N_6198,N_5672,N_5776);
nand U6199 (N_6199,N_5983,N_5532);
or U6200 (N_6200,N_5952,N_5539);
and U6201 (N_6201,N_5551,N_5968);
or U6202 (N_6202,N_5515,N_5628);
nand U6203 (N_6203,N_5875,N_5561);
and U6204 (N_6204,N_5683,N_5616);
nand U6205 (N_6205,N_5862,N_5947);
or U6206 (N_6206,N_5739,N_5885);
or U6207 (N_6207,N_5770,N_5915);
nor U6208 (N_6208,N_5935,N_5536);
nand U6209 (N_6209,N_5836,N_5999);
and U6210 (N_6210,N_5760,N_5636);
nor U6211 (N_6211,N_5682,N_5823);
and U6212 (N_6212,N_5729,N_5941);
nand U6213 (N_6213,N_5962,N_5812);
nand U6214 (N_6214,N_5658,N_5907);
and U6215 (N_6215,N_5749,N_5579);
nand U6216 (N_6216,N_5631,N_5807);
nand U6217 (N_6217,N_5657,N_5914);
nor U6218 (N_6218,N_5972,N_5988);
nor U6219 (N_6219,N_5827,N_5873);
and U6220 (N_6220,N_5844,N_5782);
or U6221 (N_6221,N_5618,N_5691);
nand U6222 (N_6222,N_5832,N_5779);
nand U6223 (N_6223,N_5949,N_5602);
nand U6224 (N_6224,N_5887,N_5677);
nand U6225 (N_6225,N_5971,N_5768);
or U6226 (N_6226,N_5667,N_5604);
nor U6227 (N_6227,N_5961,N_5774);
nand U6228 (N_6228,N_5744,N_5723);
nand U6229 (N_6229,N_5520,N_5697);
nand U6230 (N_6230,N_5653,N_5698);
nor U6231 (N_6231,N_5577,N_5831);
nand U6232 (N_6232,N_5808,N_5886);
nand U6233 (N_6233,N_5895,N_5981);
and U6234 (N_6234,N_5704,N_5991);
xnor U6235 (N_6235,N_5702,N_5746);
and U6236 (N_6236,N_5598,N_5597);
nand U6237 (N_6237,N_5959,N_5659);
or U6238 (N_6238,N_5876,N_5612);
or U6239 (N_6239,N_5556,N_5772);
nand U6240 (N_6240,N_5800,N_5720);
and U6241 (N_6241,N_5558,N_5717);
nor U6242 (N_6242,N_5714,N_5544);
nor U6243 (N_6243,N_5745,N_5665);
or U6244 (N_6244,N_5936,N_5893);
nor U6245 (N_6245,N_5858,N_5948);
or U6246 (N_6246,N_5853,N_5718);
or U6247 (N_6247,N_5998,N_5751);
xor U6248 (N_6248,N_5861,N_5678);
nand U6249 (N_6249,N_5852,N_5517);
or U6250 (N_6250,N_5946,N_5936);
nor U6251 (N_6251,N_5925,N_5835);
or U6252 (N_6252,N_5603,N_5567);
and U6253 (N_6253,N_5574,N_5761);
nor U6254 (N_6254,N_5653,N_5876);
nand U6255 (N_6255,N_5824,N_5919);
nand U6256 (N_6256,N_5500,N_5573);
and U6257 (N_6257,N_5869,N_5798);
nor U6258 (N_6258,N_5516,N_5838);
and U6259 (N_6259,N_5570,N_5547);
and U6260 (N_6260,N_5635,N_5534);
or U6261 (N_6261,N_5909,N_5541);
nand U6262 (N_6262,N_5566,N_5500);
nor U6263 (N_6263,N_5595,N_5611);
nand U6264 (N_6264,N_5736,N_5744);
nor U6265 (N_6265,N_5824,N_5742);
nand U6266 (N_6266,N_5773,N_5838);
nand U6267 (N_6267,N_5990,N_5902);
or U6268 (N_6268,N_5991,N_5602);
nand U6269 (N_6269,N_5851,N_5683);
nor U6270 (N_6270,N_5563,N_5924);
nand U6271 (N_6271,N_5542,N_5891);
or U6272 (N_6272,N_5767,N_5801);
xor U6273 (N_6273,N_5726,N_5998);
nor U6274 (N_6274,N_5629,N_5541);
nand U6275 (N_6275,N_5884,N_5688);
and U6276 (N_6276,N_5788,N_5860);
nand U6277 (N_6277,N_5616,N_5568);
nand U6278 (N_6278,N_5548,N_5776);
nand U6279 (N_6279,N_5965,N_5820);
and U6280 (N_6280,N_5886,N_5969);
or U6281 (N_6281,N_5542,N_5928);
or U6282 (N_6282,N_5500,N_5957);
nor U6283 (N_6283,N_5658,N_5753);
nor U6284 (N_6284,N_5963,N_5529);
or U6285 (N_6285,N_5554,N_5833);
nor U6286 (N_6286,N_5933,N_5528);
and U6287 (N_6287,N_5791,N_5684);
or U6288 (N_6288,N_5723,N_5874);
nand U6289 (N_6289,N_5739,N_5984);
or U6290 (N_6290,N_5872,N_5786);
nor U6291 (N_6291,N_5587,N_5935);
and U6292 (N_6292,N_5726,N_5747);
or U6293 (N_6293,N_5910,N_5926);
xor U6294 (N_6294,N_5747,N_5649);
and U6295 (N_6295,N_5671,N_5987);
or U6296 (N_6296,N_5896,N_5749);
and U6297 (N_6297,N_5539,N_5760);
nor U6298 (N_6298,N_5607,N_5534);
nor U6299 (N_6299,N_5642,N_5800);
or U6300 (N_6300,N_5600,N_5958);
or U6301 (N_6301,N_5662,N_5866);
xnor U6302 (N_6302,N_5835,N_5983);
nand U6303 (N_6303,N_5578,N_5749);
nand U6304 (N_6304,N_5532,N_5871);
or U6305 (N_6305,N_5519,N_5508);
nand U6306 (N_6306,N_5547,N_5726);
xor U6307 (N_6307,N_5999,N_5969);
or U6308 (N_6308,N_5775,N_5820);
xnor U6309 (N_6309,N_5587,N_5991);
nand U6310 (N_6310,N_5737,N_5743);
and U6311 (N_6311,N_5974,N_5874);
or U6312 (N_6312,N_5616,N_5970);
nand U6313 (N_6313,N_5882,N_5998);
nand U6314 (N_6314,N_5506,N_5526);
xor U6315 (N_6315,N_5742,N_5950);
nand U6316 (N_6316,N_5965,N_5983);
and U6317 (N_6317,N_5642,N_5983);
nor U6318 (N_6318,N_5883,N_5827);
or U6319 (N_6319,N_5542,N_5938);
nand U6320 (N_6320,N_5525,N_5980);
or U6321 (N_6321,N_5747,N_5766);
nor U6322 (N_6322,N_5982,N_5930);
or U6323 (N_6323,N_5829,N_5975);
nand U6324 (N_6324,N_5581,N_5612);
nor U6325 (N_6325,N_5677,N_5933);
nor U6326 (N_6326,N_5546,N_5737);
and U6327 (N_6327,N_5538,N_5585);
or U6328 (N_6328,N_5932,N_5895);
nand U6329 (N_6329,N_5655,N_5952);
and U6330 (N_6330,N_5837,N_5886);
or U6331 (N_6331,N_5873,N_5757);
xnor U6332 (N_6332,N_5836,N_5778);
nand U6333 (N_6333,N_5919,N_5687);
or U6334 (N_6334,N_5572,N_5872);
or U6335 (N_6335,N_5789,N_5981);
and U6336 (N_6336,N_5531,N_5762);
and U6337 (N_6337,N_5546,N_5943);
and U6338 (N_6338,N_5964,N_5862);
and U6339 (N_6339,N_5653,N_5835);
and U6340 (N_6340,N_5741,N_5941);
or U6341 (N_6341,N_5836,N_5946);
nand U6342 (N_6342,N_5962,N_5847);
and U6343 (N_6343,N_5860,N_5942);
or U6344 (N_6344,N_5701,N_5729);
and U6345 (N_6345,N_5599,N_5753);
nor U6346 (N_6346,N_5546,N_5562);
or U6347 (N_6347,N_5919,N_5951);
or U6348 (N_6348,N_5811,N_5918);
and U6349 (N_6349,N_5849,N_5759);
nor U6350 (N_6350,N_5539,N_5920);
nand U6351 (N_6351,N_5799,N_5545);
and U6352 (N_6352,N_5814,N_5907);
or U6353 (N_6353,N_5930,N_5853);
nand U6354 (N_6354,N_5541,N_5511);
nand U6355 (N_6355,N_5953,N_5525);
nand U6356 (N_6356,N_5717,N_5531);
nand U6357 (N_6357,N_5585,N_5533);
nor U6358 (N_6358,N_5537,N_5647);
and U6359 (N_6359,N_5896,N_5757);
or U6360 (N_6360,N_5521,N_5574);
nor U6361 (N_6361,N_5676,N_5847);
or U6362 (N_6362,N_5798,N_5844);
or U6363 (N_6363,N_5623,N_5724);
and U6364 (N_6364,N_5953,N_5620);
nor U6365 (N_6365,N_5720,N_5743);
and U6366 (N_6366,N_5693,N_5986);
or U6367 (N_6367,N_5546,N_5607);
nor U6368 (N_6368,N_5856,N_5747);
and U6369 (N_6369,N_5974,N_5574);
nor U6370 (N_6370,N_5661,N_5570);
nand U6371 (N_6371,N_5567,N_5637);
nand U6372 (N_6372,N_5595,N_5663);
or U6373 (N_6373,N_5678,N_5630);
xnor U6374 (N_6374,N_5914,N_5709);
and U6375 (N_6375,N_5891,N_5597);
nand U6376 (N_6376,N_5709,N_5550);
nor U6377 (N_6377,N_5711,N_5980);
nor U6378 (N_6378,N_5980,N_5806);
nand U6379 (N_6379,N_5577,N_5524);
nand U6380 (N_6380,N_5592,N_5653);
nand U6381 (N_6381,N_5729,N_5890);
and U6382 (N_6382,N_5541,N_5517);
nand U6383 (N_6383,N_5666,N_5901);
nand U6384 (N_6384,N_5909,N_5521);
nand U6385 (N_6385,N_5766,N_5929);
and U6386 (N_6386,N_5672,N_5724);
or U6387 (N_6387,N_5752,N_5651);
or U6388 (N_6388,N_5646,N_5643);
or U6389 (N_6389,N_5698,N_5943);
nor U6390 (N_6390,N_5992,N_5996);
or U6391 (N_6391,N_5507,N_5938);
or U6392 (N_6392,N_5857,N_5646);
nand U6393 (N_6393,N_5695,N_5696);
or U6394 (N_6394,N_5933,N_5514);
nor U6395 (N_6395,N_5789,N_5692);
or U6396 (N_6396,N_5723,N_5549);
nor U6397 (N_6397,N_5524,N_5973);
nand U6398 (N_6398,N_5694,N_5583);
or U6399 (N_6399,N_5640,N_5984);
nor U6400 (N_6400,N_5942,N_5693);
nor U6401 (N_6401,N_5894,N_5630);
nor U6402 (N_6402,N_5669,N_5997);
nand U6403 (N_6403,N_5683,N_5665);
and U6404 (N_6404,N_5623,N_5813);
or U6405 (N_6405,N_5569,N_5534);
nand U6406 (N_6406,N_5592,N_5933);
nor U6407 (N_6407,N_5632,N_5697);
nand U6408 (N_6408,N_5713,N_5907);
or U6409 (N_6409,N_5809,N_5721);
and U6410 (N_6410,N_5973,N_5640);
nand U6411 (N_6411,N_5677,N_5681);
xnor U6412 (N_6412,N_5799,N_5920);
nor U6413 (N_6413,N_5529,N_5514);
and U6414 (N_6414,N_5718,N_5521);
xor U6415 (N_6415,N_5970,N_5840);
or U6416 (N_6416,N_5626,N_5829);
nor U6417 (N_6417,N_5632,N_5569);
nand U6418 (N_6418,N_5591,N_5771);
or U6419 (N_6419,N_5607,N_5961);
nor U6420 (N_6420,N_5812,N_5850);
and U6421 (N_6421,N_5591,N_5969);
or U6422 (N_6422,N_5636,N_5581);
or U6423 (N_6423,N_5851,N_5649);
nor U6424 (N_6424,N_5567,N_5985);
or U6425 (N_6425,N_5564,N_5550);
nor U6426 (N_6426,N_5573,N_5698);
nand U6427 (N_6427,N_5680,N_5854);
or U6428 (N_6428,N_5544,N_5676);
or U6429 (N_6429,N_5616,N_5715);
or U6430 (N_6430,N_5968,N_5906);
or U6431 (N_6431,N_5703,N_5704);
or U6432 (N_6432,N_5522,N_5730);
nand U6433 (N_6433,N_5898,N_5633);
nor U6434 (N_6434,N_5662,N_5573);
nor U6435 (N_6435,N_5562,N_5947);
or U6436 (N_6436,N_5692,N_5726);
and U6437 (N_6437,N_5667,N_5705);
or U6438 (N_6438,N_5875,N_5965);
nor U6439 (N_6439,N_5547,N_5982);
nor U6440 (N_6440,N_5582,N_5819);
nor U6441 (N_6441,N_5993,N_5644);
nand U6442 (N_6442,N_5633,N_5648);
or U6443 (N_6443,N_5527,N_5890);
or U6444 (N_6444,N_5988,N_5650);
nand U6445 (N_6445,N_5757,N_5598);
nand U6446 (N_6446,N_5584,N_5908);
nor U6447 (N_6447,N_5703,N_5853);
nor U6448 (N_6448,N_5903,N_5600);
nand U6449 (N_6449,N_5508,N_5703);
nand U6450 (N_6450,N_5923,N_5954);
nand U6451 (N_6451,N_5873,N_5703);
xor U6452 (N_6452,N_5678,N_5594);
and U6453 (N_6453,N_5935,N_5544);
xnor U6454 (N_6454,N_5911,N_5774);
and U6455 (N_6455,N_5753,N_5737);
nor U6456 (N_6456,N_5552,N_5776);
or U6457 (N_6457,N_5861,N_5719);
xor U6458 (N_6458,N_5646,N_5508);
or U6459 (N_6459,N_5837,N_5866);
and U6460 (N_6460,N_5816,N_5568);
or U6461 (N_6461,N_5913,N_5931);
nor U6462 (N_6462,N_5959,N_5956);
and U6463 (N_6463,N_5740,N_5863);
nor U6464 (N_6464,N_5603,N_5739);
or U6465 (N_6465,N_5806,N_5847);
and U6466 (N_6466,N_5829,N_5991);
nor U6467 (N_6467,N_5778,N_5597);
or U6468 (N_6468,N_5800,N_5710);
nor U6469 (N_6469,N_5609,N_5906);
and U6470 (N_6470,N_5666,N_5766);
or U6471 (N_6471,N_5823,N_5803);
and U6472 (N_6472,N_5857,N_5720);
or U6473 (N_6473,N_5585,N_5586);
nand U6474 (N_6474,N_5999,N_5996);
nand U6475 (N_6475,N_5763,N_5721);
xor U6476 (N_6476,N_5587,N_5971);
and U6477 (N_6477,N_5779,N_5891);
or U6478 (N_6478,N_5772,N_5947);
and U6479 (N_6479,N_5551,N_5790);
nand U6480 (N_6480,N_5737,N_5584);
or U6481 (N_6481,N_5829,N_5539);
and U6482 (N_6482,N_5824,N_5848);
or U6483 (N_6483,N_5660,N_5607);
or U6484 (N_6484,N_5924,N_5512);
nor U6485 (N_6485,N_5806,N_5738);
and U6486 (N_6486,N_5834,N_5825);
nor U6487 (N_6487,N_5813,N_5647);
and U6488 (N_6488,N_5867,N_5535);
nor U6489 (N_6489,N_5899,N_5677);
or U6490 (N_6490,N_5956,N_5888);
or U6491 (N_6491,N_5883,N_5877);
and U6492 (N_6492,N_5638,N_5821);
nor U6493 (N_6493,N_5823,N_5667);
nor U6494 (N_6494,N_5864,N_5830);
xnor U6495 (N_6495,N_5581,N_5964);
or U6496 (N_6496,N_5799,N_5890);
and U6497 (N_6497,N_5518,N_5988);
or U6498 (N_6498,N_5870,N_5979);
nor U6499 (N_6499,N_5685,N_5828);
nor U6500 (N_6500,N_6271,N_6175);
nor U6501 (N_6501,N_6161,N_6221);
nand U6502 (N_6502,N_6337,N_6327);
and U6503 (N_6503,N_6371,N_6341);
nand U6504 (N_6504,N_6269,N_6007);
or U6505 (N_6505,N_6344,N_6101);
xnor U6506 (N_6506,N_6200,N_6331);
xnor U6507 (N_6507,N_6323,N_6381);
nor U6508 (N_6508,N_6495,N_6455);
nor U6509 (N_6509,N_6148,N_6472);
nand U6510 (N_6510,N_6287,N_6485);
and U6511 (N_6511,N_6017,N_6074);
xor U6512 (N_6512,N_6284,N_6235);
or U6513 (N_6513,N_6231,N_6185);
and U6514 (N_6514,N_6237,N_6443);
nor U6515 (N_6515,N_6088,N_6199);
or U6516 (N_6516,N_6095,N_6498);
or U6517 (N_6517,N_6251,N_6339);
nor U6518 (N_6518,N_6418,N_6034);
nand U6519 (N_6519,N_6187,N_6044);
nand U6520 (N_6520,N_6014,N_6479);
or U6521 (N_6521,N_6475,N_6273);
or U6522 (N_6522,N_6109,N_6283);
nor U6523 (N_6523,N_6459,N_6484);
or U6524 (N_6524,N_6093,N_6153);
nor U6525 (N_6525,N_6154,N_6480);
and U6526 (N_6526,N_6233,N_6321);
and U6527 (N_6527,N_6334,N_6328);
nand U6528 (N_6528,N_6388,N_6184);
and U6529 (N_6529,N_6340,N_6456);
and U6530 (N_6530,N_6057,N_6298);
and U6531 (N_6531,N_6083,N_6037);
nor U6532 (N_6532,N_6202,N_6322);
nor U6533 (N_6533,N_6238,N_6268);
and U6534 (N_6534,N_6402,N_6391);
or U6535 (N_6535,N_6280,N_6058);
nor U6536 (N_6536,N_6416,N_6397);
and U6537 (N_6537,N_6469,N_6038);
and U6538 (N_6538,N_6377,N_6068);
and U6539 (N_6539,N_6229,N_6216);
and U6540 (N_6540,N_6009,N_6055);
and U6541 (N_6541,N_6206,N_6129);
nor U6542 (N_6542,N_6299,N_6180);
and U6543 (N_6543,N_6019,N_6156);
and U6544 (N_6544,N_6252,N_6125);
nor U6545 (N_6545,N_6470,N_6174);
and U6546 (N_6546,N_6225,N_6390);
nand U6547 (N_6547,N_6304,N_6043);
or U6548 (N_6548,N_6031,N_6127);
nor U6549 (N_6549,N_6393,N_6433);
nand U6550 (N_6550,N_6330,N_6279);
and U6551 (N_6551,N_6369,N_6318);
nand U6552 (N_6552,N_6414,N_6305);
and U6553 (N_6553,N_6285,N_6030);
or U6554 (N_6554,N_6203,N_6438);
nor U6555 (N_6555,N_6210,N_6142);
nand U6556 (N_6556,N_6368,N_6296);
and U6557 (N_6557,N_6449,N_6073);
nand U6558 (N_6558,N_6158,N_6020);
or U6559 (N_6559,N_6473,N_6119);
nand U6560 (N_6560,N_6159,N_6496);
nor U6561 (N_6561,N_6167,N_6364);
and U6562 (N_6562,N_6071,N_6054);
nor U6563 (N_6563,N_6403,N_6214);
or U6564 (N_6564,N_6164,N_6080);
and U6565 (N_6565,N_6267,N_6482);
or U6566 (N_6566,N_6315,N_6316);
and U6567 (N_6567,N_6471,N_6489);
nand U6568 (N_6568,N_6442,N_6274);
and U6569 (N_6569,N_6089,N_6432);
or U6570 (N_6570,N_6060,N_6086);
or U6571 (N_6571,N_6295,N_6363);
nand U6572 (N_6572,N_6181,N_6049);
nor U6573 (N_6573,N_6146,N_6445);
and U6574 (N_6574,N_6145,N_6050);
nand U6575 (N_6575,N_6032,N_6103);
and U6576 (N_6576,N_6491,N_6487);
nor U6577 (N_6577,N_6224,N_6313);
nor U6578 (N_6578,N_6270,N_6400);
xor U6579 (N_6579,N_6041,N_6163);
nand U6580 (N_6580,N_6133,N_6178);
nand U6581 (N_6581,N_6292,N_6215);
nor U6582 (N_6582,N_6053,N_6128);
or U6583 (N_6583,N_6157,N_6326);
or U6584 (N_6584,N_6275,N_6162);
nor U6585 (N_6585,N_6423,N_6182);
or U6586 (N_6586,N_6309,N_6261);
nor U6587 (N_6587,N_6349,N_6065);
nand U6588 (N_6588,N_6205,N_6351);
and U6589 (N_6589,N_6490,N_6492);
and U6590 (N_6590,N_6176,N_6412);
nand U6591 (N_6591,N_6173,N_6421);
nand U6592 (N_6592,N_6462,N_6066);
nor U6593 (N_6593,N_6047,N_6311);
nand U6594 (N_6594,N_6481,N_6389);
nand U6595 (N_6595,N_6352,N_6499);
nand U6596 (N_6596,N_6383,N_6264);
and U6597 (N_6597,N_6144,N_6234);
and U6598 (N_6598,N_6107,N_6335);
nand U6599 (N_6599,N_6218,N_6370);
and U6600 (N_6600,N_6067,N_6282);
nor U6601 (N_6601,N_6121,N_6192);
nand U6602 (N_6602,N_6018,N_6426);
or U6603 (N_6603,N_6061,N_6168);
or U6604 (N_6604,N_6272,N_6072);
nand U6605 (N_6605,N_6276,N_6120);
nand U6606 (N_6606,N_6246,N_6110);
and U6607 (N_6607,N_6006,N_6406);
nand U6608 (N_6608,N_6422,N_6353);
nand U6609 (N_6609,N_6436,N_6413);
or U6610 (N_6610,N_6005,N_6076);
nand U6611 (N_6611,N_6004,N_6379);
or U6612 (N_6612,N_6293,N_6198);
nor U6613 (N_6613,N_6451,N_6035);
and U6614 (N_6614,N_6011,N_6317);
and U6615 (N_6615,N_6213,N_6189);
nor U6616 (N_6616,N_6427,N_6051);
nand U6617 (N_6617,N_6149,N_6130);
or U6618 (N_6618,N_6140,N_6244);
or U6619 (N_6619,N_6429,N_6171);
nor U6620 (N_6620,N_6376,N_6108);
nand U6621 (N_6621,N_6241,N_6294);
xnor U6622 (N_6622,N_6398,N_6036);
nand U6623 (N_6623,N_6113,N_6085);
or U6624 (N_6624,N_6118,N_6262);
and U6625 (N_6625,N_6424,N_6230);
or U6626 (N_6626,N_6139,N_6029);
and U6627 (N_6627,N_6342,N_6355);
nor U6628 (N_6628,N_6408,N_6420);
and U6629 (N_6629,N_6132,N_6466);
nor U6630 (N_6630,N_6314,N_6281);
and U6631 (N_6631,N_6301,N_6223);
or U6632 (N_6632,N_6105,N_6266);
or U6633 (N_6633,N_6114,N_6190);
nand U6634 (N_6634,N_6468,N_6117);
and U6635 (N_6635,N_6098,N_6253);
or U6636 (N_6636,N_6063,N_6493);
or U6637 (N_6637,N_6025,N_6361);
nand U6638 (N_6638,N_6405,N_6415);
and U6639 (N_6639,N_6291,N_6112);
nor U6640 (N_6640,N_6476,N_6226);
or U6641 (N_6641,N_6228,N_6012);
nor U6642 (N_6642,N_6106,N_6010);
and U6643 (N_6643,N_6082,N_6263);
and U6644 (N_6644,N_6141,N_6325);
and U6645 (N_6645,N_6197,N_6135);
nor U6646 (N_6646,N_6079,N_6245);
nor U6647 (N_6647,N_6399,N_6046);
nand U6648 (N_6648,N_6147,N_6052);
and U6649 (N_6649,N_6417,N_6434);
nor U6650 (N_6650,N_6394,N_6249);
nor U6651 (N_6651,N_6260,N_6166);
nor U6652 (N_6652,N_6392,N_6401);
or U6653 (N_6653,N_6457,N_6022);
nor U6654 (N_6654,N_6220,N_6155);
nand U6655 (N_6655,N_6099,N_6212);
and U6656 (N_6656,N_6123,N_6042);
and U6657 (N_6657,N_6409,N_6463);
nor U6658 (N_6658,N_6465,N_6336);
nor U6659 (N_6659,N_6345,N_6302);
and U6660 (N_6660,N_6346,N_6090);
xnor U6661 (N_6661,N_6453,N_6290);
or U6662 (N_6662,N_6458,N_6332);
and U6663 (N_6663,N_6454,N_6059);
nor U6664 (N_6664,N_6333,N_6039);
nand U6665 (N_6665,N_6188,N_6122);
or U6666 (N_6666,N_6186,N_6069);
or U6667 (N_6667,N_6040,N_6378);
nand U6668 (N_6668,N_6435,N_6385);
or U6669 (N_6669,N_6165,N_6239);
or U6670 (N_6670,N_6056,N_6021);
nor U6671 (N_6671,N_6460,N_6070);
and U6672 (N_6672,N_6115,N_6373);
or U6673 (N_6673,N_6307,N_6087);
nor U6674 (N_6674,N_6045,N_6000);
nor U6675 (N_6675,N_6134,N_6195);
or U6676 (N_6676,N_6138,N_6104);
and U6677 (N_6677,N_6124,N_6026);
or U6678 (N_6678,N_6137,N_6257);
and U6679 (N_6679,N_6191,N_6407);
and U6680 (N_6680,N_6348,N_6126);
nor U6681 (N_6681,N_6028,N_6209);
and U6682 (N_6682,N_6478,N_6467);
or U6683 (N_6683,N_6062,N_6419);
or U6684 (N_6684,N_6446,N_6078);
or U6685 (N_6685,N_6094,N_6372);
or U6686 (N_6686,N_6319,N_6461);
nor U6687 (N_6687,N_6360,N_6247);
nand U6688 (N_6688,N_6256,N_6300);
nand U6689 (N_6689,N_6359,N_6303);
and U6690 (N_6690,N_6324,N_6136);
nand U6691 (N_6691,N_6306,N_6013);
or U6692 (N_6692,N_6102,N_6227);
or U6693 (N_6693,N_6404,N_6365);
or U6694 (N_6694,N_6437,N_6312);
nor U6695 (N_6695,N_6248,N_6354);
or U6696 (N_6696,N_6236,N_6343);
and U6697 (N_6697,N_6177,N_6092);
nand U6698 (N_6698,N_6208,N_6152);
and U6699 (N_6699,N_6265,N_6183);
nand U6700 (N_6700,N_6425,N_6483);
and U6701 (N_6701,N_6016,N_6350);
nand U6702 (N_6702,N_6380,N_6320);
or U6703 (N_6703,N_6131,N_6447);
or U6704 (N_6704,N_6286,N_6477);
and U6705 (N_6705,N_6204,N_6064);
xor U6706 (N_6706,N_6410,N_6024);
nand U6707 (N_6707,N_6091,N_6362);
or U6708 (N_6708,N_6207,N_6075);
or U6709 (N_6709,N_6430,N_6096);
or U6710 (N_6710,N_6289,N_6366);
nor U6711 (N_6711,N_6201,N_6358);
nand U6712 (N_6712,N_6277,N_6193);
or U6713 (N_6713,N_6150,N_6452);
or U6714 (N_6714,N_6396,N_6243);
and U6715 (N_6715,N_6015,N_6081);
nand U6716 (N_6716,N_6440,N_6448);
or U6717 (N_6717,N_6329,N_6217);
nor U6718 (N_6718,N_6374,N_6367);
and U6719 (N_6719,N_6001,N_6084);
or U6720 (N_6720,N_6258,N_6464);
or U6721 (N_6721,N_6278,N_6003);
nor U6722 (N_6722,N_6211,N_6338);
nand U6723 (N_6723,N_6441,N_6387);
nand U6724 (N_6724,N_6310,N_6111);
nor U6725 (N_6725,N_6386,N_6116);
and U6726 (N_6726,N_6033,N_6497);
xnor U6727 (N_6727,N_6219,N_6488);
nand U6728 (N_6728,N_6382,N_6172);
or U6729 (N_6729,N_6194,N_6170);
and U6730 (N_6730,N_6431,N_6428);
nand U6731 (N_6731,N_6439,N_6048);
nor U6732 (N_6732,N_6395,N_6151);
xor U6733 (N_6733,N_6077,N_6232);
nor U6734 (N_6734,N_6384,N_6356);
or U6735 (N_6735,N_6242,N_6143);
or U6736 (N_6736,N_6160,N_6008);
or U6737 (N_6737,N_6023,N_6222);
nand U6738 (N_6738,N_6255,N_6100);
nand U6739 (N_6739,N_6254,N_6474);
or U6740 (N_6740,N_6288,N_6450);
and U6741 (N_6741,N_6297,N_6375);
nand U6742 (N_6742,N_6357,N_6444);
nor U6743 (N_6743,N_6411,N_6486);
and U6744 (N_6744,N_6097,N_6250);
nor U6745 (N_6745,N_6179,N_6002);
nand U6746 (N_6746,N_6494,N_6240);
nand U6747 (N_6747,N_6308,N_6347);
nor U6748 (N_6748,N_6196,N_6027);
nand U6749 (N_6749,N_6259,N_6169);
or U6750 (N_6750,N_6131,N_6025);
or U6751 (N_6751,N_6194,N_6035);
nand U6752 (N_6752,N_6155,N_6496);
or U6753 (N_6753,N_6444,N_6073);
xnor U6754 (N_6754,N_6070,N_6450);
or U6755 (N_6755,N_6438,N_6355);
or U6756 (N_6756,N_6113,N_6041);
and U6757 (N_6757,N_6124,N_6348);
and U6758 (N_6758,N_6459,N_6307);
and U6759 (N_6759,N_6371,N_6383);
nor U6760 (N_6760,N_6044,N_6188);
nor U6761 (N_6761,N_6457,N_6185);
nand U6762 (N_6762,N_6401,N_6263);
or U6763 (N_6763,N_6389,N_6295);
nand U6764 (N_6764,N_6255,N_6288);
and U6765 (N_6765,N_6112,N_6297);
nand U6766 (N_6766,N_6108,N_6195);
nand U6767 (N_6767,N_6427,N_6458);
or U6768 (N_6768,N_6353,N_6201);
nand U6769 (N_6769,N_6032,N_6228);
nor U6770 (N_6770,N_6201,N_6229);
nand U6771 (N_6771,N_6104,N_6005);
or U6772 (N_6772,N_6481,N_6224);
nor U6773 (N_6773,N_6479,N_6498);
nand U6774 (N_6774,N_6052,N_6272);
and U6775 (N_6775,N_6482,N_6404);
or U6776 (N_6776,N_6376,N_6032);
nand U6777 (N_6777,N_6273,N_6235);
nand U6778 (N_6778,N_6139,N_6160);
nor U6779 (N_6779,N_6473,N_6154);
nor U6780 (N_6780,N_6198,N_6412);
nand U6781 (N_6781,N_6000,N_6338);
or U6782 (N_6782,N_6293,N_6188);
and U6783 (N_6783,N_6201,N_6287);
nor U6784 (N_6784,N_6009,N_6407);
nor U6785 (N_6785,N_6436,N_6321);
nor U6786 (N_6786,N_6353,N_6106);
or U6787 (N_6787,N_6205,N_6376);
or U6788 (N_6788,N_6334,N_6349);
and U6789 (N_6789,N_6200,N_6375);
or U6790 (N_6790,N_6256,N_6454);
nor U6791 (N_6791,N_6151,N_6349);
nor U6792 (N_6792,N_6393,N_6376);
xor U6793 (N_6793,N_6284,N_6186);
nor U6794 (N_6794,N_6252,N_6376);
nor U6795 (N_6795,N_6116,N_6238);
and U6796 (N_6796,N_6246,N_6002);
nand U6797 (N_6797,N_6319,N_6050);
or U6798 (N_6798,N_6299,N_6115);
or U6799 (N_6799,N_6493,N_6166);
nor U6800 (N_6800,N_6208,N_6249);
nor U6801 (N_6801,N_6421,N_6076);
or U6802 (N_6802,N_6360,N_6114);
nand U6803 (N_6803,N_6026,N_6175);
nor U6804 (N_6804,N_6318,N_6036);
and U6805 (N_6805,N_6167,N_6135);
nor U6806 (N_6806,N_6317,N_6167);
or U6807 (N_6807,N_6031,N_6386);
or U6808 (N_6808,N_6120,N_6261);
xnor U6809 (N_6809,N_6216,N_6471);
nor U6810 (N_6810,N_6288,N_6377);
nand U6811 (N_6811,N_6023,N_6301);
and U6812 (N_6812,N_6453,N_6348);
nand U6813 (N_6813,N_6220,N_6298);
nand U6814 (N_6814,N_6229,N_6279);
nand U6815 (N_6815,N_6465,N_6056);
nor U6816 (N_6816,N_6090,N_6301);
or U6817 (N_6817,N_6053,N_6207);
and U6818 (N_6818,N_6337,N_6290);
and U6819 (N_6819,N_6026,N_6429);
nand U6820 (N_6820,N_6285,N_6307);
nor U6821 (N_6821,N_6038,N_6149);
and U6822 (N_6822,N_6306,N_6321);
and U6823 (N_6823,N_6112,N_6411);
or U6824 (N_6824,N_6012,N_6352);
nor U6825 (N_6825,N_6296,N_6364);
nand U6826 (N_6826,N_6384,N_6248);
nand U6827 (N_6827,N_6310,N_6397);
or U6828 (N_6828,N_6035,N_6251);
and U6829 (N_6829,N_6217,N_6350);
nor U6830 (N_6830,N_6490,N_6265);
or U6831 (N_6831,N_6244,N_6337);
and U6832 (N_6832,N_6279,N_6467);
and U6833 (N_6833,N_6144,N_6477);
and U6834 (N_6834,N_6104,N_6173);
nor U6835 (N_6835,N_6449,N_6154);
nor U6836 (N_6836,N_6054,N_6289);
or U6837 (N_6837,N_6064,N_6049);
and U6838 (N_6838,N_6019,N_6083);
nand U6839 (N_6839,N_6227,N_6357);
nand U6840 (N_6840,N_6240,N_6311);
nor U6841 (N_6841,N_6027,N_6475);
nand U6842 (N_6842,N_6229,N_6303);
or U6843 (N_6843,N_6191,N_6231);
and U6844 (N_6844,N_6412,N_6194);
and U6845 (N_6845,N_6112,N_6212);
nor U6846 (N_6846,N_6492,N_6215);
and U6847 (N_6847,N_6344,N_6229);
and U6848 (N_6848,N_6366,N_6284);
nand U6849 (N_6849,N_6208,N_6229);
and U6850 (N_6850,N_6193,N_6356);
or U6851 (N_6851,N_6497,N_6499);
and U6852 (N_6852,N_6182,N_6228);
or U6853 (N_6853,N_6216,N_6411);
nand U6854 (N_6854,N_6400,N_6311);
and U6855 (N_6855,N_6275,N_6369);
nand U6856 (N_6856,N_6352,N_6331);
xor U6857 (N_6857,N_6246,N_6166);
or U6858 (N_6858,N_6139,N_6395);
nor U6859 (N_6859,N_6385,N_6364);
and U6860 (N_6860,N_6290,N_6033);
and U6861 (N_6861,N_6499,N_6380);
nand U6862 (N_6862,N_6058,N_6459);
and U6863 (N_6863,N_6018,N_6177);
nor U6864 (N_6864,N_6383,N_6107);
and U6865 (N_6865,N_6491,N_6287);
and U6866 (N_6866,N_6485,N_6232);
and U6867 (N_6867,N_6220,N_6163);
nand U6868 (N_6868,N_6020,N_6136);
xnor U6869 (N_6869,N_6209,N_6185);
or U6870 (N_6870,N_6029,N_6247);
nor U6871 (N_6871,N_6000,N_6188);
and U6872 (N_6872,N_6296,N_6241);
nor U6873 (N_6873,N_6064,N_6274);
xor U6874 (N_6874,N_6377,N_6250);
and U6875 (N_6875,N_6148,N_6099);
and U6876 (N_6876,N_6445,N_6257);
nand U6877 (N_6877,N_6437,N_6120);
nor U6878 (N_6878,N_6030,N_6241);
or U6879 (N_6879,N_6013,N_6439);
or U6880 (N_6880,N_6009,N_6294);
nand U6881 (N_6881,N_6364,N_6161);
nor U6882 (N_6882,N_6152,N_6341);
or U6883 (N_6883,N_6065,N_6084);
or U6884 (N_6884,N_6160,N_6351);
nand U6885 (N_6885,N_6175,N_6163);
and U6886 (N_6886,N_6438,N_6252);
and U6887 (N_6887,N_6401,N_6028);
or U6888 (N_6888,N_6074,N_6158);
nor U6889 (N_6889,N_6322,N_6055);
and U6890 (N_6890,N_6077,N_6336);
xnor U6891 (N_6891,N_6255,N_6003);
or U6892 (N_6892,N_6309,N_6291);
nor U6893 (N_6893,N_6012,N_6113);
nand U6894 (N_6894,N_6283,N_6304);
or U6895 (N_6895,N_6279,N_6234);
nand U6896 (N_6896,N_6214,N_6062);
nand U6897 (N_6897,N_6289,N_6225);
nor U6898 (N_6898,N_6152,N_6069);
nor U6899 (N_6899,N_6422,N_6310);
nand U6900 (N_6900,N_6196,N_6413);
nor U6901 (N_6901,N_6191,N_6250);
xnor U6902 (N_6902,N_6239,N_6336);
or U6903 (N_6903,N_6233,N_6257);
and U6904 (N_6904,N_6285,N_6283);
xor U6905 (N_6905,N_6366,N_6272);
or U6906 (N_6906,N_6433,N_6176);
nor U6907 (N_6907,N_6271,N_6255);
nor U6908 (N_6908,N_6489,N_6011);
or U6909 (N_6909,N_6383,N_6327);
or U6910 (N_6910,N_6100,N_6267);
and U6911 (N_6911,N_6375,N_6243);
xnor U6912 (N_6912,N_6374,N_6379);
or U6913 (N_6913,N_6454,N_6214);
xor U6914 (N_6914,N_6095,N_6007);
nand U6915 (N_6915,N_6489,N_6178);
or U6916 (N_6916,N_6107,N_6281);
nor U6917 (N_6917,N_6455,N_6396);
nor U6918 (N_6918,N_6323,N_6435);
or U6919 (N_6919,N_6492,N_6495);
nand U6920 (N_6920,N_6462,N_6072);
nor U6921 (N_6921,N_6279,N_6255);
and U6922 (N_6922,N_6251,N_6445);
and U6923 (N_6923,N_6202,N_6125);
nor U6924 (N_6924,N_6193,N_6216);
nand U6925 (N_6925,N_6043,N_6358);
nor U6926 (N_6926,N_6155,N_6435);
xnor U6927 (N_6927,N_6199,N_6083);
xnor U6928 (N_6928,N_6278,N_6328);
nor U6929 (N_6929,N_6048,N_6247);
nor U6930 (N_6930,N_6168,N_6137);
nand U6931 (N_6931,N_6356,N_6443);
nor U6932 (N_6932,N_6174,N_6252);
and U6933 (N_6933,N_6370,N_6091);
nor U6934 (N_6934,N_6482,N_6230);
nand U6935 (N_6935,N_6201,N_6218);
or U6936 (N_6936,N_6132,N_6272);
or U6937 (N_6937,N_6313,N_6382);
nand U6938 (N_6938,N_6453,N_6059);
nand U6939 (N_6939,N_6044,N_6331);
nand U6940 (N_6940,N_6280,N_6374);
or U6941 (N_6941,N_6361,N_6382);
or U6942 (N_6942,N_6340,N_6398);
nor U6943 (N_6943,N_6119,N_6299);
nand U6944 (N_6944,N_6401,N_6036);
and U6945 (N_6945,N_6294,N_6333);
nand U6946 (N_6946,N_6264,N_6082);
xor U6947 (N_6947,N_6360,N_6190);
and U6948 (N_6948,N_6001,N_6166);
or U6949 (N_6949,N_6200,N_6121);
or U6950 (N_6950,N_6226,N_6292);
nor U6951 (N_6951,N_6326,N_6212);
and U6952 (N_6952,N_6402,N_6245);
and U6953 (N_6953,N_6050,N_6259);
and U6954 (N_6954,N_6027,N_6363);
nor U6955 (N_6955,N_6243,N_6258);
nor U6956 (N_6956,N_6377,N_6100);
xor U6957 (N_6957,N_6019,N_6299);
and U6958 (N_6958,N_6187,N_6107);
and U6959 (N_6959,N_6194,N_6388);
or U6960 (N_6960,N_6051,N_6018);
or U6961 (N_6961,N_6123,N_6022);
nor U6962 (N_6962,N_6038,N_6359);
xor U6963 (N_6963,N_6052,N_6067);
and U6964 (N_6964,N_6428,N_6389);
or U6965 (N_6965,N_6132,N_6279);
nand U6966 (N_6966,N_6262,N_6261);
xnor U6967 (N_6967,N_6429,N_6163);
xnor U6968 (N_6968,N_6003,N_6416);
nand U6969 (N_6969,N_6263,N_6482);
nand U6970 (N_6970,N_6060,N_6291);
and U6971 (N_6971,N_6069,N_6181);
or U6972 (N_6972,N_6347,N_6436);
nand U6973 (N_6973,N_6421,N_6265);
nand U6974 (N_6974,N_6363,N_6246);
nor U6975 (N_6975,N_6053,N_6089);
or U6976 (N_6976,N_6085,N_6054);
and U6977 (N_6977,N_6344,N_6287);
and U6978 (N_6978,N_6305,N_6332);
and U6979 (N_6979,N_6309,N_6052);
nor U6980 (N_6980,N_6109,N_6058);
and U6981 (N_6981,N_6022,N_6200);
or U6982 (N_6982,N_6143,N_6158);
nand U6983 (N_6983,N_6039,N_6408);
and U6984 (N_6984,N_6488,N_6400);
nor U6985 (N_6985,N_6011,N_6093);
or U6986 (N_6986,N_6346,N_6159);
nor U6987 (N_6987,N_6463,N_6042);
and U6988 (N_6988,N_6314,N_6287);
nor U6989 (N_6989,N_6352,N_6305);
or U6990 (N_6990,N_6092,N_6036);
nand U6991 (N_6991,N_6303,N_6155);
or U6992 (N_6992,N_6323,N_6338);
nand U6993 (N_6993,N_6169,N_6002);
and U6994 (N_6994,N_6484,N_6189);
or U6995 (N_6995,N_6152,N_6382);
nor U6996 (N_6996,N_6132,N_6489);
xor U6997 (N_6997,N_6347,N_6385);
nor U6998 (N_6998,N_6093,N_6416);
or U6999 (N_6999,N_6006,N_6010);
nand U7000 (N_7000,N_6836,N_6581);
and U7001 (N_7001,N_6860,N_6867);
or U7002 (N_7002,N_6864,N_6777);
or U7003 (N_7003,N_6800,N_6539);
or U7004 (N_7004,N_6805,N_6952);
nand U7005 (N_7005,N_6648,N_6826);
or U7006 (N_7006,N_6622,N_6594);
nor U7007 (N_7007,N_6775,N_6785);
nand U7008 (N_7008,N_6780,N_6715);
and U7009 (N_7009,N_6920,N_6948);
and U7010 (N_7010,N_6556,N_6956);
nand U7011 (N_7011,N_6778,N_6897);
and U7012 (N_7012,N_6570,N_6935);
or U7013 (N_7013,N_6963,N_6824);
xnor U7014 (N_7014,N_6861,N_6684);
nand U7015 (N_7015,N_6944,N_6585);
nor U7016 (N_7016,N_6662,N_6704);
nand U7017 (N_7017,N_6717,N_6808);
nand U7018 (N_7018,N_6750,N_6557);
nand U7019 (N_7019,N_6936,N_6908);
and U7020 (N_7020,N_6899,N_6840);
or U7021 (N_7021,N_6694,N_6880);
and U7022 (N_7022,N_6934,N_6979);
and U7023 (N_7023,N_6567,N_6960);
or U7024 (N_7024,N_6743,N_6900);
and U7025 (N_7025,N_6644,N_6655);
nor U7026 (N_7026,N_6583,N_6877);
and U7027 (N_7027,N_6997,N_6526);
or U7028 (N_7028,N_6533,N_6924);
nand U7029 (N_7029,N_6984,N_6951);
nand U7030 (N_7030,N_6815,N_6597);
or U7031 (N_7031,N_6548,N_6671);
and U7032 (N_7032,N_6766,N_6966);
nand U7033 (N_7033,N_6998,N_6507);
or U7034 (N_7034,N_6855,N_6504);
nor U7035 (N_7035,N_6927,N_6814);
or U7036 (N_7036,N_6933,N_6727);
nand U7037 (N_7037,N_6736,N_6573);
or U7038 (N_7038,N_6636,N_6532);
and U7039 (N_7039,N_6882,N_6500);
xor U7040 (N_7040,N_6969,N_6980);
nand U7041 (N_7041,N_6803,N_6953);
nor U7042 (N_7042,N_6914,N_6928);
nor U7043 (N_7043,N_6941,N_6901);
or U7044 (N_7044,N_6702,N_6865);
nand U7045 (N_7045,N_6930,N_6524);
or U7046 (N_7046,N_6765,N_6538);
nand U7047 (N_7047,N_6946,N_6572);
or U7048 (N_7048,N_6501,N_6962);
nand U7049 (N_7049,N_6722,N_6552);
nand U7050 (N_7050,N_6903,N_6733);
nand U7051 (N_7051,N_6858,N_6703);
nand U7052 (N_7052,N_6832,N_6641);
or U7053 (N_7053,N_6584,N_6834);
and U7054 (N_7054,N_6818,N_6620);
nor U7055 (N_7055,N_6839,N_6847);
and U7056 (N_7056,N_6918,N_6784);
xnor U7057 (N_7057,N_6673,N_6604);
nand U7058 (N_7058,N_6823,N_6838);
or U7059 (N_7059,N_6837,N_6821);
or U7060 (N_7060,N_6950,N_6626);
or U7061 (N_7061,N_6714,N_6536);
or U7062 (N_7062,N_6721,N_6608);
and U7063 (N_7063,N_6845,N_6931);
xnor U7064 (N_7064,N_6516,N_6994);
nor U7065 (N_7065,N_6764,N_6968);
and U7066 (N_7066,N_6651,N_6517);
nand U7067 (N_7067,N_6925,N_6659);
or U7068 (N_7068,N_6510,N_6866);
and U7069 (N_7069,N_6681,N_6569);
nand U7070 (N_7070,N_6791,N_6893);
or U7071 (N_7071,N_6697,N_6982);
or U7072 (N_7072,N_6844,N_6749);
and U7073 (N_7073,N_6735,N_6794);
and U7074 (N_7074,N_6521,N_6577);
and U7075 (N_7075,N_6658,N_6638);
nand U7076 (N_7076,N_6718,N_6670);
and U7077 (N_7077,N_6701,N_6896);
nand U7078 (N_7078,N_6725,N_6683);
xor U7079 (N_7079,N_6595,N_6745);
nor U7080 (N_7080,N_6522,N_6822);
or U7081 (N_7081,N_6862,N_6603);
nand U7082 (N_7082,N_6560,N_6959);
or U7083 (N_7083,N_6955,N_6787);
and U7084 (N_7084,N_6811,N_6796);
and U7085 (N_7085,N_6724,N_6964);
or U7086 (N_7086,N_6913,N_6881);
and U7087 (N_7087,N_6506,N_6712);
nor U7088 (N_7088,N_6543,N_6645);
or U7089 (N_7089,N_6910,N_6562);
or U7090 (N_7090,N_6992,N_6699);
and U7091 (N_7091,N_6661,N_6515);
nor U7092 (N_7092,N_6843,N_6664);
nor U7093 (N_7093,N_6518,N_6915);
xor U7094 (N_7094,N_6737,N_6906);
nor U7095 (N_7095,N_6761,N_6827);
nor U7096 (N_7096,N_6663,N_6898);
nand U7097 (N_7097,N_6841,N_6647);
and U7098 (N_7098,N_6523,N_6793);
or U7099 (N_7099,N_6879,N_6949);
and U7100 (N_7100,N_6688,N_6639);
and U7101 (N_7101,N_6576,N_6609);
nor U7102 (N_7102,N_6762,N_6601);
xnor U7103 (N_7103,N_6978,N_6873);
and U7104 (N_7104,N_6563,N_6973);
or U7105 (N_7105,N_6753,N_6876);
or U7106 (N_7106,N_6729,N_6829);
and U7107 (N_7107,N_6503,N_6580);
or U7108 (N_7108,N_6614,N_6961);
or U7109 (N_7109,N_6640,N_6752);
or U7110 (N_7110,N_6676,N_6875);
nand U7111 (N_7111,N_6972,N_6652);
and U7112 (N_7112,N_6687,N_6530);
nand U7113 (N_7113,N_6895,N_6977);
nand U7114 (N_7114,N_6565,N_6774);
nand U7115 (N_7115,N_6561,N_6911);
nor U7116 (N_7116,N_6600,N_6535);
nor U7117 (N_7117,N_6932,N_6617);
nand U7118 (N_7118,N_6891,N_6967);
nand U7119 (N_7119,N_6635,N_6546);
xnor U7120 (N_7120,N_6686,N_6923);
nor U7121 (N_7121,N_6942,N_6534);
or U7122 (N_7122,N_6654,N_6857);
nor U7123 (N_7123,N_6739,N_6642);
nor U7124 (N_7124,N_6947,N_6544);
and U7125 (N_7125,N_6842,N_6799);
nand U7126 (N_7126,N_6709,N_6741);
or U7127 (N_7127,N_6868,N_6682);
and U7128 (N_7128,N_6835,N_6767);
nor U7129 (N_7129,N_6631,N_6888);
nor U7130 (N_7130,N_6742,N_6731);
nor U7131 (N_7131,N_6940,N_6760);
nor U7132 (N_7132,N_6738,N_6678);
nand U7133 (N_7133,N_6666,N_6613);
and U7134 (N_7134,N_6730,N_6669);
or U7135 (N_7135,N_6574,N_6575);
nor U7136 (N_7136,N_6751,N_6586);
nor U7137 (N_7137,N_6553,N_6975);
and U7138 (N_7138,N_6549,N_6719);
nor U7139 (N_7139,N_6711,N_6945);
xor U7140 (N_7140,N_6525,N_6769);
and U7141 (N_7141,N_6619,N_6502);
or U7142 (N_7142,N_6590,N_6989);
nand U7143 (N_7143,N_6810,N_6887);
nor U7144 (N_7144,N_6537,N_6813);
and U7145 (N_7145,N_6917,N_6754);
nand U7146 (N_7146,N_6759,N_6716);
nand U7147 (N_7147,N_6792,N_6568);
nand U7148 (N_7148,N_6596,N_6675);
nor U7149 (N_7149,N_6606,N_6559);
nand U7150 (N_7150,N_6598,N_6564);
nand U7151 (N_7151,N_6825,N_6788);
nand U7152 (N_7152,N_6599,N_6587);
and U7153 (N_7153,N_6783,N_6612);
xor U7154 (N_7154,N_6710,N_6996);
nand U7155 (N_7155,N_6852,N_6804);
or U7156 (N_7156,N_6905,N_6909);
or U7157 (N_7157,N_6693,N_6912);
nor U7158 (N_7158,N_6939,N_6871);
or U7159 (N_7159,N_6519,N_6633);
nor U7160 (N_7160,N_6902,N_6732);
or U7161 (N_7161,N_6720,N_6520);
and U7162 (N_7162,N_6916,N_6801);
or U7163 (N_7163,N_6611,N_6929);
nand U7164 (N_7164,N_6831,N_6650);
nand U7165 (N_7165,N_6884,N_6665);
nand U7166 (N_7166,N_6547,N_6505);
nand U7167 (N_7167,N_6907,N_6630);
and U7168 (N_7168,N_6589,N_6615);
or U7169 (N_7169,N_6726,N_6554);
and U7170 (N_7170,N_6623,N_6634);
or U7171 (N_7171,N_6685,N_6734);
or U7172 (N_7172,N_6781,N_6758);
xnor U7173 (N_7173,N_6943,N_6723);
nor U7174 (N_7174,N_6593,N_6571);
nand U7175 (N_7175,N_6995,N_6856);
or U7176 (N_7176,N_6649,N_6629);
or U7177 (N_7177,N_6653,N_6886);
nand U7178 (N_7178,N_6894,N_6643);
nor U7179 (N_7179,N_6812,N_6610);
nor U7180 (N_7180,N_6987,N_6851);
nand U7181 (N_7181,N_6602,N_6981);
or U7182 (N_7182,N_6983,N_6846);
and U7183 (N_7183,N_6677,N_6954);
nand U7184 (N_7184,N_6999,N_6691);
and U7185 (N_7185,N_6582,N_6937);
and U7186 (N_7186,N_6779,N_6528);
nor U7187 (N_7187,N_6698,N_6773);
nor U7188 (N_7188,N_6957,N_6926);
or U7189 (N_7189,N_6668,N_6706);
nor U7190 (N_7190,N_6607,N_6705);
nand U7191 (N_7191,N_6807,N_6511);
or U7192 (N_7192,N_6890,N_6786);
nand U7193 (N_7193,N_6588,N_6904);
or U7194 (N_7194,N_6755,N_6798);
or U7195 (N_7195,N_6889,N_6993);
and U7196 (N_7196,N_6797,N_6551);
nand U7197 (N_7197,N_6820,N_6878);
or U7198 (N_7198,N_6744,N_6970);
nor U7199 (N_7199,N_6853,N_6508);
or U7200 (N_7200,N_6892,N_6768);
nor U7201 (N_7201,N_6618,N_6531);
nor U7202 (N_7202,N_6869,N_6833);
nor U7203 (N_7203,N_6605,N_6806);
and U7204 (N_7204,N_6632,N_6789);
nand U7205 (N_7205,N_6657,N_6828);
or U7206 (N_7206,N_6885,N_6819);
or U7207 (N_7207,N_6624,N_6692);
xor U7208 (N_7208,N_6919,N_6921);
and U7209 (N_7209,N_6541,N_6863);
nor U7210 (N_7210,N_6874,N_6859);
nand U7211 (N_7211,N_6848,N_6555);
and U7212 (N_7212,N_6816,N_6795);
nand U7213 (N_7213,N_6802,N_6625);
or U7214 (N_7214,N_6991,N_6696);
nand U7215 (N_7215,N_6747,N_6756);
nand U7216 (N_7216,N_6700,N_6646);
and U7217 (N_7217,N_6854,N_6512);
and U7218 (N_7218,N_6771,N_6509);
nand U7219 (N_7219,N_6637,N_6695);
and U7220 (N_7220,N_6990,N_6817);
or U7221 (N_7221,N_6757,N_6514);
and U7222 (N_7222,N_6772,N_6849);
xor U7223 (N_7223,N_6672,N_6986);
nand U7224 (N_7224,N_6690,N_6558);
and U7225 (N_7225,N_6621,N_6872);
and U7226 (N_7226,N_6850,N_6579);
and U7227 (N_7227,N_6922,N_6971);
nor U7228 (N_7228,N_6809,N_6965);
nor U7229 (N_7229,N_6988,N_6674);
or U7230 (N_7230,N_6776,N_6707);
nand U7231 (N_7231,N_6974,N_6770);
and U7232 (N_7232,N_6529,N_6870);
nand U7233 (N_7233,N_6628,N_6592);
nor U7234 (N_7234,N_6938,N_6708);
or U7235 (N_7235,N_6680,N_6790);
or U7236 (N_7236,N_6883,N_6830);
and U7237 (N_7237,N_6746,N_6679);
nand U7238 (N_7238,N_6740,N_6513);
nand U7239 (N_7239,N_6667,N_6542);
or U7240 (N_7240,N_6763,N_6748);
nand U7241 (N_7241,N_6540,N_6689);
nand U7242 (N_7242,N_6976,N_6591);
nor U7243 (N_7243,N_6578,N_6545);
nand U7244 (N_7244,N_6713,N_6566);
and U7245 (N_7245,N_6728,N_6550);
and U7246 (N_7246,N_6656,N_6958);
nand U7247 (N_7247,N_6527,N_6782);
or U7248 (N_7248,N_6660,N_6627);
and U7249 (N_7249,N_6616,N_6985);
nor U7250 (N_7250,N_6810,N_6531);
nand U7251 (N_7251,N_6835,N_6788);
or U7252 (N_7252,N_6589,N_6745);
nor U7253 (N_7253,N_6938,N_6773);
and U7254 (N_7254,N_6928,N_6523);
nor U7255 (N_7255,N_6766,N_6709);
and U7256 (N_7256,N_6810,N_6799);
nand U7257 (N_7257,N_6549,N_6831);
nand U7258 (N_7258,N_6652,N_6554);
or U7259 (N_7259,N_6572,N_6789);
and U7260 (N_7260,N_6964,N_6904);
or U7261 (N_7261,N_6733,N_6668);
nand U7262 (N_7262,N_6958,N_6951);
or U7263 (N_7263,N_6978,N_6664);
and U7264 (N_7264,N_6541,N_6909);
or U7265 (N_7265,N_6670,N_6819);
or U7266 (N_7266,N_6742,N_6818);
and U7267 (N_7267,N_6959,N_6752);
or U7268 (N_7268,N_6825,N_6710);
or U7269 (N_7269,N_6842,N_6834);
nor U7270 (N_7270,N_6511,N_6627);
nor U7271 (N_7271,N_6997,N_6616);
nor U7272 (N_7272,N_6784,N_6922);
or U7273 (N_7273,N_6807,N_6726);
and U7274 (N_7274,N_6681,N_6771);
and U7275 (N_7275,N_6932,N_6594);
nor U7276 (N_7276,N_6781,N_6833);
xnor U7277 (N_7277,N_6785,N_6514);
or U7278 (N_7278,N_6847,N_6794);
xnor U7279 (N_7279,N_6514,N_6863);
or U7280 (N_7280,N_6819,N_6800);
and U7281 (N_7281,N_6966,N_6667);
or U7282 (N_7282,N_6888,N_6955);
nor U7283 (N_7283,N_6990,N_6563);
nand U7284 (N_7284,N_6859,N_6909);
nor U7285 (N_7285,N_6788,N_6938);
or U7286 (N_7286,N_6880,N_6529);
nor U7287 (N_7287,N_6693,N_6781);
or U7288 (N_7288,N_6779,N_6929);
and U7289 (N_7289,N_6700,N_6625);
nor U7290 (N_7290,N_6776,N_6572);
and U7291 (N_7291,N_6744,N_6880);
xor U7292 (N_7292,N_6641,N_6752);
nand U7293 (N_7293,N_6568,N_6978);
nor U7294 (N_7294,N_6823,N_6623);
nand U7295 (N_7295,N_6802,N_6589);
or U7296 (N_7296,N_6953,N_6690);
and U7297 (N_7297,N_6607,N_6790);
and U7298 (N_7298,N_6801,N_6866);
or U7299 (N_7299,N_6528,N_6874);
nor U7300 (N_7300,N_6670,N_6926);
nand U7301 (N_7301,N_6917,N_6889);
nor U7302 (N_7302,N_6975,N_6537);
nand U7303 (N_7303,N_6657,N_6522);
nand U7304 (N_7304,N_6713,N_6919);
nor U7305 (N_7305,N_6825,N_6964);
nand U7306 (N_7306,N_6869,N_6664);
and U7307 (N_7307,N_6758,N_6809);
nor U7308 (N_7308,N_6946,N_6584);
nor U7309 (N_7309,N_6761,N_6809);
nand U7310 (N_7310,N_6624,N_6849);
nand U7311 (N_7311,N_6994,N_6549);
and U7312 (N_7312,N_6670,N_6773);
nand U7313 (N_7313,N_6703,N_6761);
or U7314 (N_7314,N_6742,N_6664);
and U7315 (N_7315,N_6918,N_6849);
nor U7316 (N_7316,N_6949,N_6553);
nor U7317 (N_7317,N_6661,N_6612);
nand U7318 (N_7318,N_6575,N_6619);
and U7319 (N_7319,N_6749,N_6978);
nand U7320 (N_7320,N_6613,N_6842);
and U7321 (N_7321,N_6690,N_6550);
or U7322 (N_7322,N_6511,N_6895);
and U7323 (N_7323,N_6505,N_6795);
and U7324 (N_7324,N_6849,N_6935);
or U7325 (N_7325,N_6867,N_6518);
and U7326 (N_7326,N_6839,N_6558);
or U7327 (N_7327,N_6786,N_6771);
nor U7328 (N_7328,N_6595,N_6961);
and U7329 (N_7329,N_6943,N_6724);
and U7330 (N_7330,N_6571,N_6757);
or U7331 (N_7331,N_6599,N_6573);
or U7332 (N_7332,N_6709,N_6654);
or U7333 (N_7333,N_6779,N_6751);
xnor U7334 (N_7334,N_6720,N_6967);
nand U7335 (N_7335,N_6933,N_6651);
and U7336 (N_7336,N_6625,N_6626);
nand U7337 (N_7337,N_6676,N_6963);
nor U7338 (N_7338,N_6630,N_6911);
nor U7339 (N_7339,N_6558,N_6597);
nand U7340 (N_7340,N_6554,N_6681);
or U7341 (N_7341,N_6846,N_6704);
nor U7342 (N_7342,N_6586,N_6599);
or U7343 (N_7343,N_6914,N_6850);
or U7344 (N_7344,N_6918,N_6868);
or U7345 (N_7345,N_6894,N_6535);
or U7346 (N_7346,N_6964,N_6996);
nor U7347 (N_7347,N_6608,N_6889);
or U7348 (N_7348,N_6956,N_6740);
and U7349 (N_7349,N_6990,N_6907);
nor U7350 (N_7350,N_6624,N_6580);
nand U7351 (N_7351,N_6525,N_6716);
nor U7352 (N_7352,N_6522,N_6967);
and U7353 (N_7353,N_6774,N_6670);
nor U7354 (N_7354,N_6818,N_6514);
nor U7355 (N_7355,N_6533,N_6819);
nand U7356 (N_7356,N_6546,N_6839);
nand U7357 (N_7357,N_6503,N_6955);
and U7358 (N_7358,N_6647,N_6762);
or U7359 (N_7359,N_6746,N_6701);
nand U7360 (N_7360,N_6857,N_6694);
nor U7361 (N_7361,N_6997,N_6808);
and U7362 (N_7362,N_6876,N_6821);
nand U7363 (N_7363,N_6984,N_6921);
nor U7364 (N_7364,N_6935,N_6520);
or U7365 (N_7365,N_6695,N_6697);
nor U7366 (N_7366,N_6595,N_6979);
and U7367 (N_7367,N_6849,N_6928);
or U7368 (N_7368,N_6574,N_6853);
xnor U7369 (N_7369,N_6636,N_6808);
nand U7370 (N_7370,N_6537,N_6720);
nand U7371 (N_7371,N_6600,N_6646);
or U7372 (N_7372,N_6580,N_6510);
nor U7373 (N_7373,N_6662,N_6750);
nand U7374 (N_7374,N_6874,N_6592);
and U7375 (N_7375,N_6640,N_6941);
or U7376 (N_7376,N_6829,N_6897);
or U7377 (N_7377,N_6723,N_6685);
nor U7378 (N_7378,N_6892,N_6987);
nand U7379 (N_7379,N_6991,N_6544);
or U7380 (N_7380,N_6701,N_6551);
or U7381 (N_7381,N_6714,N_6531);
or U7382 (N_7382,N_6700,N_6500);
and U7383 (N_7383,N_6743,N_6526);
nand U7384 (N_7384,N_6512,N_6804);
nand U7385 (N_7385,N_6768,N_6550);
or U7386 (N_7386,N_6837,N_6657);
nor U7387 (N_7387,N_6923,N_6989);
and U7388 (N_7388,N_6985,N_6651);
nor U7389 (N_7389,N_6575,N_6867);
and U7390 (N_7390,N_6556,N_6738);
or U7391 (N_7391,N_6708,N_6896);
nand U7392 (N_7392,N_6870,N_6533);
or U7393 (N_7393,N_6699,N_6501);
nor U7394 (N_7394,N_6685,N_6589);
and U7395 (N_7395,N_6531,N_6939);
nor U7396 (N_7396,N_6987,N_6543);
or U7397 (N_7397,N_6702,N_6905);
and U7398 (N_7398,N_6960,N_6693);
or U7399 (N_7399,N_6720,N_6947);
and U7400 (N_7400,N_6965,N_6963);
nand U7401 (N_7401,N_6624,N_6515);
nand U7402 (N_7402,N_6915,N_6859);
or U7403 (N_7403,N_6946,N_6803);
nand U7404 (N_7404,N_6655,N_6786);
nor U7405 (N_7405,N_6638,N_6721);
nand U7406 (N_7406,N_6551,N_6859);
and U7407 (N_7407,N_6617,N_6912);
nand U7408 (N_7408,N_6608,N_6836);
nand U7409 (N_7409,N_6848,N_6801);
and U7410 (N_7410,N_6657,N_6785);
nand U7411 (N_7411,N_6875,N_6691);
or U7412 (N_7412,N_6906,N_6776);
and U7413 (N_7413,N_6850,N_6866);
or U7414 (N_7414,N_6569,N_6965);
and U7415 (N_7415,N_6514,N_6974);
or U7416 (N_7416,N_6635,N_6616);
and U7417 (N_7417,N_6782,N_6512);
or U7418 (N_7418,N_6747,N_6657);
nor U7419 (N_7419,N_6946,N_6707);
and U7420 (N_7420,N_6569,N_6600);
nand U7421 (N_7421,N_6618,N_6784);
nor U7422 (N_7422,N_6523,N_6870);
nor U7423 (N_7423,N_6848,N_6807);
and U7424 (N_7424,N_6836,N_6770);
nor U7425 (N_7425,N_6874,N_6515);
or U7426 (N_7426,N_6685,N_6855);
nand U7427 (N_7427,N_6867,N_6865);
and U7428 (N_7428,N_6544,N_6569);
and U7429 (N_7429,N_6589,N_6585);
and U7430 (N_7430,N_6893,N_6760);
nor U7431 (N_7431,N_6793,N_6644);
and U7432 (N_7432,N_6831,N_6748);
nand U7433 (N_7433,N_6672,N_6603);
or U7434 (N_7434,N_6930,N_6853);
and U7435 (N_7435,N_6600,N_6774);
or U7436 (N_7436,N_6976,N_6735);
or U7437 (N_7437,N_6599,N_6906);
or U7438 (N_7438,N_6745,N_6671);
nor U7439 (N_7439,N_6713,N_6616);
nor U7440 (N_7440,N_6711,N_6987);
or U7441 (N_7441,N_6652,N_6627);
or U7442 (N_7442,N_6750,N_6916);
nor U7443 (N_7443,N_6735,N_6552);
xnor U7444 (N_7444,N_6812,N_6736);
and U7445 (N_7445,N_6609,N_6656);
nand U7446 (N_7446,N_6521,N_6952);
nand U7447 (N_7447,N_6943,N_6589);
nor U7448 (N_7448,N_6536,N_6786);
or U7449 (N_7449,N_6833,N_6650);
and U7450 (N_7450,N_6816,N_6824);
and U7451 (N_7451,N_6992,N_6528);
nor U7452 (N_7452,N_6966,N_6526);
and U7453 (N_7453,N_6910,N_6612);
nand U7454 (N_7454,N_6604,N_6829);
and U7455 (N_7455,N_6795,N_6606);
or U7456 (N_7456,N_6538,N_6709);
nand U7457 (N_7457,N_6911,N_6837);
nor U7458 (N_7458,N_6984,N_6512);
xnor U7459 (N_7459,N_6973,N_6730);
nor U7460 (N_7460,N_6980,N_6584);
nand U7461 (N_7461,N_6686,N_6535);
and U7462 (N_7462,N_6910,N_6682);
and U7463 (N_7463,N_6831,N_6672);
or U7464 (N_7464,N_6527,N_6978);
nand U7465 (N_7465,N_6594,N_6522);
nor U7466 (N_7466,N_6774,N_6901);
and U7467 (N_7467,N_6935,N_6693);
nand U7468 (N_7468,N_6844,N_6544);
nand U7469 (N_7469,N_6700,N_6784);
nor U7470 (N_7470,N_6621,N_6511);
and U7471 (N_7471,N_6795,N_6576);
nand U7472 (N_7472,N_6825,N_6730);
nand U7473 (N_7473,N_6706,N_6890);
nand U7474 (N_7474,N_6704,N_6592);
nor U7475 (N_7475,N_6882,N_6739);
nand U7476 (N_7476,N_6531,N_6649);
and U7477 (N_7477,N_6696,N_6789);
or U7478 (N_7478,N_6914,N_6540);
nor U7479 (N_7479,N_6916,N_6847);
or U7480 (N_7480,N_6954,N_6932);
nand U7481 (N_7481,N_6992,N_6606);
nor U7482 (N_7482,N_6999,N_6505);
and U7483 (N_7483,N_6579,N_6793);
or U7484 (N_7484,N_6746,N_6884);
or U7485 (N_7485,N_6912,N_6692);
or U7486 (N_7486,N_6951,N_6852);
and U7487 (N_7487,N_6974,N_6705);
or U7488 (N_7488,N_6629,N_6982);
nand U7489 (N_7489,N_6705,N_6598);
nor U7490 (N_7490,N_6878,N_6745);
and U7491 (N_7491,N_6517,N_6532);
and U7492 (N_7492,N_6994,N_6867);
nand U7493 (N_7493,N_6764,N_6791);
nand U7494 (N_7494,N_6573,N_6786);
or U7495 (N_7495,N_6971,N_6959);
nand U7496 (N_7496,N_6918,N_6778);
nand U7497 (N_7497,N_6913,N_6901);
or U7498 (N_7498,N_6805,N_6673);
or U7499 (N_7499,N_6731,N_6970);
nand U7500 (N_7500,N_7483,N_7257);
or U7501 (N_7501,N_7112,N_7078);
nor U7502 (N_7502,N_7044,N_7148);
nand U7503 (N_7503,N_7183,N_7052);
or U7504 (N_7504,N_7457,N_7166);
nand U7505 (N_7505,N_7201,N_7425);
nor U7506 (N_7506,N_7437,N_7102);
nand U7507 (N_7507,N_7247,N_7194);
nand U7508 (N_7508,N_7096,N_7448);
nor U7509 (N_7509,N_7222,N_7233);
and U7510 (N_7510,N_7465,N_7382);
and U7511 (N_7511,N_7270,N_7126);
nand U7512 (N_7512,N_7241,N_7008);
nand U7513 (N_7513,N_7197,N_7340);
xor U7514 (N_7514,N_7121,N_7424);
and U7515 (N_7515,N_7427,N_7151);
or U7516 (N_7516,N_7310,N_7309);
xor U7517 (N_7517,N_7317,N_7398);
or U7518 (N_7518,N_7307,N_7130);
nand U7519 (N_7519,N_7407,N_7447);
and U7520 (N_7520,N_7179,N_7205);
and U7521 (N_7521,N_7258,N_7288);
xnor U7522 (N_7522,N_7097,N_7279);
nor U7523 (N_7523,N_7423,N_7452);
nor U7524 (N_7524,N_7069,N_7381);
and U7525 (N_7525,N_7215,N_7024);
nor U7526 (N_7526,N_7314,N_7181);
nor U7527 (N_7527,N_7090,N_7421);
nand U7528 (N_7528,N_7083,N_7195);
nor U7529 (N_7529,N_7039,N_7054);
nor U7530 (N_7530,N_7167,N_7059);
or U7531 (N_7531,N_7162,N_7362);
nand U7532 (N_7532,N_7139,N_7359);
nand U7533 (N_7533,N_7220,N_7101);
and U7534 (N_7534,N_7445,N_7371);
or U7535 (N_7535,N_7210,N_7060);
nor U7536 (N_7536,N_7116,N_7107);
nor U7537 (N_7537,N_7497,N_7253);
nand U7538 (N_7538,N_7079,N_7113);
and U7539 (N_7539,N_7466,N_7429);
xor U7540 (N_7540,N_7211,N_7461);
or U7541 (N_7541,N_7003,N_7063);
nor U7542 (N_7542,N_7203,N_7485);
nand U7543 (N_7543,N_7152,N_7141);
nand U7544 (N_7544,N_7456,N_7185);
and U7545 (N_7545,N_7200,N_7088);
nand U7546 (N_7546,N_7093,N_7408);
nor U7547 (N_7547,N_7091,N_7396);
xnor U7548 (N_7548,N_7420,N_7482);
nor U7549 (N_7549,N_7490,N_7412);
or U7550 (N_7550,N_7099,N_7234);
and U7551 (N_7551,N_7388,N_7009);
xnor U7552 (N_7552,N_7277,N_7394);
and U7553 (N_7553,N_7391,N_7272);
nand U7554 (N_7554,N_7082,N_7037);
nand U7555 (N_7555,N_7468,N_7248);
or U7556 (N_7556,N_7496,N_7165);
nand U7557 (N_7557,N_7259,N_7287);
and U7558 (N_7558,N_7263,N_7454);
and U7559 (N_7559,N_7046,N_7393);
and U7560 (N_7560,N_7415,N_7467);
nand U7561 (N_7561,N_7012,N_7158);
or U7562 (N_7562,N_7308,N_7439);
or U7563 (N_7563,N_7401,N_7074);
and U7564 (N_7564,N_7295,N_7219);
and U7565 (N_7565,N_7299,N_7182);
nand U7566 (N_7566,N_7291,N_7389);
nand U7567 (N_7567,N_7418,N_7395);
or U7568 (N_7568,N_7062,N_7092);
nor U7569 (N_7569,N_7402,N_7020);
and U7570 (N_7570,N_7072,N_7123);
and U7571 (N_7571,N_7014,N_7264);
nand U7572 (N_7572,N_7055,N_7216);
nand U7573 (N_7573,N_7479,N_7489);
or U7574 (N_7574,N_7184,N_7202);
nand U7575 (N_7575,N_7084,N_7118);
and U7576 (N_7576,N_7328,N_7443);
or U7577 (N_7577,N_7019,N_7207);
and U7578 (N_7578,N_7385,N_7144);
nor U7579 (N_7579,N_7463,N_7089);
nand U7580 (N_7580,N_7323,N_7494);
or U7581 (N_7581,N_7224,N_7064);
nor U7582 (N_7582,N_7453,N_7322);
and U7583 (N_7583,N_7026,N_7305);
or U7584 (N_7584,N_7032,N_7127);
nand U7585 (N_7585,N_7278,N_7337);
and U7586 (N_7586,N_7364,N_7469);
nor U7587 (N_7587,N_7142,N_7232);
xor U7588 (N_7588,N_7285,N_7071);
and U7589 (N_7589,N_7329,N_7325);
nand U7590 (N_7590,N_7034,N_7297);
and U7591 (N_7591,N_7360,N_7397);
and U7592 (N_7592,N_7035,N_7392);
nor U7593 (N_7593,N_7106,N_7411);
or U7594 (N_7594,N_7251,N_7492);
and U7595 (N_7595,N_7372,N_7068);
or U7596 (N_7596,N_7140,N_7135);
nor U7597 (N_7597,N_7189,N_7378);
nand U7598 (N_7598,N_7261,N_7262);
nor U7599 (N_7599,N_7406,N_7004);
or U7600 (N_7600,N_7221,N_7174);
xor U7601 (N_7601,N_7256,N_7498);
nor U7602 (N_7602,N_7341,N_7146);
and U7603 (N_7603,N_7137,N_7336);
or U7604 (N_7604,N_7306,N_7414);
nor U7605 (N_7605,N_7073,N_7161);
nand U7606 (N_7606,N_7086,N_7348);
nor U7607 (N_7607,N_7041,N_7303);
and U7608 (N_7608,N_7001,N_7358);
or U7609 (N_7609,N_7376,N_7236);
and U7610 (N_7610,N_7000,N_7486);
nand U7611 (N_7611,N_7134,N_7300);
xor U7612 (N_7612,N_7168,N_7242);
nor U7613 (N_7613,N_7110,N_7190);
nand U7614 (N_7614,N_7380,N_7212);
nor U7615 (N_7615,N_7440,N_7171);
or U7616 (N_7616,N_7370,N_7361);
or U7617 (N_7617,N_7345,N_7192);
nand U7618 (N_7618,N_7246,N_7449);
and U7619 (N_7619,N_7390,N_7484);
nand U7620 (N_7620,N_7013,N_7301);
nand U7621 (N_7621,N_7087,N_7374);
nand U7622 (N_7622,N_7163,N_7157);
or U7623 (N_7623,N_7103,N_7217);
or U7624 (N_7624,N_7357,N_7373);
nor U7625 (N_7625,N_7386,N_7051);
nand U7626 (N_7626,N_7493,N_7455);
and U7627 (N_7627,N_7464,N_7172);
and U7628 (N_7628,N_7267,N_7255);
or U7629 (N_7629,N_7209,N_7442);
or U7630 (N_7630,N_7298,N_7472);
nand U7631 (N_7631,N_7413,N_7284);
nor U7632 (N_7632,N_7332,N_7023);
nor U7633 (N_7633,N_7047,N_7302);
nor U7634 (N_7634,N_7399,N_7354);
or U7635 (N_7635,N_7353,N_7477);
and U7636 (N_7636,N_7265,N_7153);
or U7637 (N_7637,N_7196,N_7094);
nand U7638 (N_7638,N_7237,N_7080);
nor U7639 (N_7639,N_7122,N_7027);
nor U7640 (N_7640,N_7108,N_7095);
or U7641 (N_7641,N_7231,N_7098);
or U7642 (N_7642,N_7347,N_7109);
nand U7643 (N_7643,N_7254,N_7434);
nor U7644 (N_7644,N_7030,N_7349);
and U7645 (N_7645,N_7160,N_7033);
nor U7646 (N_7646,N_7346,N_7495);
or U7647 (N_7647,N_7076,N_7104);
nor U7648 (N_7648,N_7176,N_7419);
and U7649 (N_7649,N_7159,N_7015);
nand U7650 (N_7650,N_7010,N_7316);
xor U7651 (N_7651,N_7198,N_7245);
or U7652 (N_7652,N_7487,N_7199);
xnor U7653 (N_7653,N_7066,N_7342);
nand U7654 (N_7654,N_7252,N_7249);
nor U7655 (N_7655,N_7131,N_7223);
and U7656 (N_7656,N_7040,N_7460);
or U7657 (N_7657,N_7475,N_7061);
and U7658 (N_7658,N_7471,N_7244);
and U7659 (N_7659,N_7450,N_7250);
nor U7660 (N_7660,N_7327,N_7204);
nor U7661 (N_7661,N_7011,N_7339);
and U7662 (N_7662,N_7147,N_7441);
or U7663 (N_7663,N_7124,N_7289);
and U7664 (N_7664,N_7100,N_7228);
or U7665 (N_7665,N_7227,N_7038);
and U7666 (N_7666,N_7433,N_7311);
and U7667 (N_7667,N_7006,N_7042);
nor U7668 (N_7668,N_7156,N_7180);
or U7669 (N_7669,N_7269,N_7114);
or U7670 (N_7670,N_7111,N_7164);
and U7671 (N_7671,N_7356,N_7286);
and U7672 (N_7672,N_7312,N_7025);
or U7673 (N_7673,N_7077,N_7384);
nand U7674 (N_7674,N_7375,N_7294);
nor U7675 (N_7675,N_7326,N_7075);
or U7676 (N_7676,N_7343,N_7007);
nor U7677 (N_7677,N_7186,N_7459);
nand U7678 (N_7678,N_7324,N_7155);
and U7679 (N_7679,N_7018,N_7260);
nor U7680 (N_7680,N_7335,N_7022);
nor U7681 (N_7681,N_7333,N_7473);
nor U7682 (N_7682,N_7214,N_7292);
nor U7683 (N_7683,N_7352,N_7321);
or U7684 (N_7684,N_7451,N_7017);
nor U7685 (N_7685,N_7048,N_7143);
nor U7686 (N_7686,N_7369,N_7053);
xnor U7687 (N_7687,N_7435,N_7320);
and U7688 (N_7688,N_7149,N_7235);
and U7689 (N_7689,N_7319,N_7383);
nor U7690 (N_7690,N_7191,N_7119);
and U7691 (N_7691,N_7028,N_7170);
and U7692 (N_7692,N_7428,N_7338);
and U7693 (N_7693,N_7276,N_7085);
xor U7694 (N_7694,N_7274,N_7056);
and U7695 (N_7695,N_7188,N_7315);
nand U7696 (N_7696,N_7462,N_7225);
or U7697 (N_7697,N_7128,N_7070);
nor U7698 (N_7698,N_7368,N_7036);
and U7699 (N_7699,N_7367,N_7243);
and U7700 (N_7700,N_7120,N_7363);
or U7701 (N_7701,N_7344,N_7387);
nor U7702 (N_7702,N_7350,N_7029);
and U7703 (N_7703,N_7230,N_7173);
or U7704 (N_7704,N_7005,N_7138);
and U7705 (N_7705,N_7043,N_7226);
nand U7706 (N_7706,N_7405,N_7175);
and U7707 (N_7707,N_7065,N_7403);
xor U7708 (N_7708,N_7436,N_7377);
nor U7709 (N_7709,N_7458,N_7355);
or U7710 (N_7710,N_7208,N_7187);
or U7711 (N_7711,N_7115,N_7240);
nor U7712 (N_7712,N_7273,N_7290);
nor U7713 (N_7713,N_7193,N_7281);
and U7714 (N_7714,N_7478,N_7050);
nor U7715 (N_7715,N_7266,N_7422);
nor U7716 (N_7716,N_7331,N_7431);
nor U7717 (N_7717,N_7499,N_7296);
and U7718 (N_7718,N_7271,N_7049);
and U7719 (N_7719,N_7379,N_7206);
nor U7720 (N_7720,N_7067,N_7409);
or U7721 (N_7721,N_7318,N_7238);
nor U7722 (N_7722,N_7432,N_7132);
nand U7723 (N_7723,N_7282,N_7145);
nand U7724 (N_7724,N_7304,N_7133);
or U7725 (N_7725,N_7438,N_7365);
nor U7726 (N_7726,N_7081,N_7117);
nor U7727 (N_7727,N_7351,N_7021);
or U7728 (N_7728,N_7045,N_7366);
nand U7729 (N_7729,N_7400,N_7031);
and U7730 (N_7730,N_7491,N_7275);
nand U7731 (N_7731,N_7426,N_7470);
nor U7732 (N_7732,N_7154,N_7169);
nand U7733 (N_7733,N_7330,N_7218);
and U7734 (N_7734,N_7016,N_7177);
and U7735 (N_7735,N_7178,N_7058);
nand U7736 (N_7736,N_7476,N_7481);
nand U7737 (N_7737,N_7129,N_7334);
nand U7738 (N_7738,N_7105,N_7239);
xnor U7739 (N_7739,N_7283,N_7444);
nand U7740 (N_7740,N_7002,N_7446);
or U7741 (N_7741,N_7404,N_7125);
nor U7742 (N_7742,N_7313,N_7268);
nand U7743 (N_7743,N_7474,N_7480);
and U7744 (N_7744,N_7430,N_7213);
and U7745 (N_7745,N_7136,N_7057);
nor U7746 (N_7746,N_7293,N_7417);
or U7747 (N_7747,N_7280,N_7416);
and U7748 (N_7748,N_7150,N_7410);
or U7749 (N_7749,N_7229,N_7488);
nand U7750 (N_7750,N_7142,N_7433);
or U7751 (N_7751,N_7008,N_7489);
and U7752 (N_7752,N_7216,N_7123);
nand U7753 (N_7753,N_7439,N_7353);
and U7754 (N_7754,N_7274,N_7435);
nand U7755 (N_7755,N_7265,N_7112);
and U7756 (N_7756,N_7434,N_7169);
nor U7757 (N_7757,N_7258,N_7090);
nor U7758 (N_7758,N_7169,N_7220);
or U7759 (N_7759,N_7176,N_7292);
and U7760 (N_7760,N_7146,N_7199);
or U7761 (N_7761,N_7111,N_7054);
nor U7762 (N_7762,N_7130,N_7425);
and U7763 (N_7763,N_7289,N_7318);
nor U7764 (N_7764,N_7022,N_7127);
or U7765 (N_7765,N_7069,N_7446);
and U7766 (N_7766,N_7474,N_7384);
and U7767 (N_7767,N_7365,N_7456);
nor U7768 (N_7768,N_7213,N_7422);
nand U7769 (N_7769,N_7316,N_7052);
and U7770 (N_7770,N_7050,N_7084);
nand U7771 (N_7771,N_7430,N_7204);
or U7772 (N_7772,N_7456,N_7401);
nor U7773 (N_7773,N_7435,N_7082);
nor U7774 (N_7774,N_7397,N_7240);
nand U7775 (N_7775,N_7192,N_7458);
nor U7776 (N_7776,N_7005,N_7159);
nor U7777 (N_7777,N_7466,N_7491);
nand U7778 (N_7778,N_7471,N_7296);
nand U7779 (N_7779,N_7419,N_7052);
nand U7780 (N_7780,N_7423,N_7373);
and U7781 (N_7781,N_7296,N_7299);
nor U7782 (N_7782,N_7332,N_7461);
and U7783 (N_7783,N_7191,N_7247);
or U7784 (N_7784,N_7342,N_7279);
nand U7785 (N_7785,N_7074,N_7468);
nand U7786 (N_7786,N_7469,N_7051);
nand U7787 (N_7787,N_7100,N_7334);
and U7788 (N_7788,N_7474,N_7121);
or U7789 (N_7789,N_7044,N_7430);
and U7790 (N_7790,N_7157,N_7025);
and U7791 (N_7791,N_7280,N_7149);
nor U7792 (N_7792,N_7173,N_7202);
and U7793 (N_7793,N_7133,N_7120);
nor U7794 (N_7794,N_7159,N_7442);
xnor U7795 (N_7795,N_7133,N_7329);
nor U7796 (N_7796,N_7432,N_7190);
or U7797 (N_7797,N_7320,N_7218);
nand U7798 (N_7798,N_7365,N_7417);
nand U7799 (N_7799,N_7484,N_7455);
nand U7800 (N_7800,N_7444,N_7452);
and U7801 (N_7801,N_7168,N_7084);
and U7802 (N_7802,N_7368,N_7032);
nand U7803 (N_7803,N_7454,N_7457);
nor U7804 (N_7804,N_7056,N_7457);
or U7805 (N_7805,N_7357,N_7183);
and U7806 (N_7806,N_7356,N_7160);
nor U7807 (N_7807,N_7083,N_7385);
nand U7808 (N_7808,N_7032,N_7238);
or U7809 (N_7809,N_7015,N_7337);
nor U7810 (N_7810,N_7241,N_7423);
and U7811 (N_7811,N_7075,N_7409);
nor U7812 (N_7812,N_7441,N_7328);
xnor U7813 (N_7813,N_7239,N_7462);
and U7814 (N_7814,N_7384,N_7447);
and U7815 (N_7815,N_7029,N_7060);
and U7816 (N_7816,N_7404,N_7330);
xnor U7817 (N_7817,N_7014,N_7158);
or U7818 (N_7818,N_7336,N_7483);
or U7819 (N_7819,N_7144,N_7437);
and U7820 (N_7820,N_7298,N_7060);
or U7821 (N_7821,N_7288,N_7210);
or U7822 (N_7822,N_7476,N_7314);
xor U7823 (N_7823,N_7359,N_7356);
or U7824 (N_7824,N_7001,N_7157);
nand U7825 (N_7825,N_7366,N_7348);
nand U7826 (N_7826,N_7466,N_7293);
and U7827 (N_7827,N_7388,N_7086);
or U7828 (N_7828,N_7189,N_7192);
nor U7829 (N_7829,N_7361,N_7303);
nand U7830 (N_7830,N_7094,N_7193);
or U7831 (N_7831,N_7402,N_7260);
nand U7832 (N_7832,N_7123,N_7045);
nand U7833 (N_7833,N_7127,N_7338);
nor U7834 (N_7834,N_7426,N_7415);
and U7835 (N_7835,N_7487,N_7423);
nor U7836 (N_7836,N_7047,N_7086);
or U7837 (N_7837,N_7484,N_7259);
nor U7838 (N_7838,N_7066,N_7370);
nand U7839 (N_7839,N_7488,N_7191);
nor U7840 (N_7840,N_7038,N_7031);
or U7841 (N_7841,N_7259,N_7167);
nor U7842 (N_7842,N_7184,N_7182);
nand U7843 (N_7843,N_7301,N_7392);
nand U7844 (N_7844,N_7409,N_7090);
and U7845 (N_7845,N_7062,N_7301);
and U7846 (N_7846,N_7271,N_7385);
xnor U7847 (N_7847,N_7072,N_7011);
nor U7848 (N_7848,N_7460,N_7116);
or U7849 (N_7849,N_7129,N_7463);
and U7850 (N_7850,N_7195,N_7077);
and U7851 (N_7851,N_7279,N_7281);
and U7852 (N_7852,N_7067,N_7412);
nor U7853 (N_7853,N_7081,N_7070);
nor U7854 (N_7854,N_7172,N_7118);
nor U7855 (N_7855,N_7263,N_7447);
nor U7856 (N_7856,N_7096,N_7277);
and U7857 (N_7857,N_7250,N_7178);
xnor U7858 (N_7858,N_7020,N_7431);
nand U7859 (N_7859,N_7030,N_7478);
nand U7860 (N_7860,N_7475,N_7332);
nor U7861 (N_7861,N_7208,N_7026);
and U7862 (N_7862,N_7219,N_7255);
or U7863 (N_7863,N_7288,N_7292);
and U7864 (N_7864,N_7209,N_7491);
and U7865 (N_7865,N_7188,N_7194);
xnor U7866 (N_7866,N_7356,N_7003);
and U7867 (N_7867,N_7156,N_7021);
nor U7868 (N_7868,N_7344,N_7460);
nor U7869 (N_7869,N_7475,N_7028);
nand U7870 (N_7870,N_7494,N_7088);
nor U7871 (N_7871,N_7055,N_7045);
xor U7872 (N_7872,N_7488,N_7328);
nor U7873 (N_7873,N_7010,N_7272);
or U7874 (N_7874,N_7359,N_7387);
nand U7875 (N_7875,N_7013,N_7213);
and U7876 (N_7876,N_7432,N_7034);
nand U7877 (N_7877,N_7149,N_7428);
xor U7878 (N_7878,N_7281,N_7200);
nand U7879 (N_7879,N_7170,N_7062);
nor U7880 (N_7880,N_7194,N_7039);
and U7881 (N_7881,N_7144,N_7362);
nor U7882 (N_7882,N_7058,N_7034);
and U7883 (N_7883,N_7002,N_7390);
nor U7884 (N_7884,N_7084,N_7335);
or U7885 (N_7885,N_7467,N_7345);
and U7886 (N_7886,N_7208,N_7383);
or U7887 (N_7887,N_7071,N_7142);
and U7888 (N_7888,N_7339,N_7134);
or U7889 (N_7889,N_7269,N_7352);
nor U7890 (N_7890,N_7319,N_7105);
or U7891 (N_7891,N_7251,N_7435);
nand U7892 (N_7892,N_7261,N_7113);
nand U7893 (N_7893,N_7279,N_7442);
nor U7894 (N_7894,N_7098,N_7029);
nand U7895 (N_7895,N_7432,N_7164);
or U7896 (N_7896,N_7068,N_7030);
nand U7897 (N_7897,N_7464,N_7229);
nand U7898 (N_7898,N_7442,N_7475);
nor U7899 (N_7899,N_7407,N_7107);
nor U7900 (N_7900,N_7388,N_7268);
or U7901 (N_7901,N_7274,N_7431);
or U7902 (N_7902,N_7380,N_7285);
or U7903 (N_7903,N_7454,N_7300);
and U7904 (N_7904,N_7053,N_7130);
and U7905 (N_7905,N_7157,N_7428);
nor U7906 (N_7906,N_7029,N_7322);
nand U7907 (N_7907,N_7397,N_7344);
nand U7908 (N_7908,N_7166,N_7437);
or U7909 (N_7909,N_7360,N_7289);
and U7910 (N_7910,N_7391,N_7421);
xnor U7911 (N_7911,N_7329,N_7239);
nor U7912 (N_7912,N_7344,N_7406);
and U7913 (N_7913,N_7227,N_7073);
nand U7914 (N_7914,N_7478,N_7335);
or U7915 (N_7915,N_7491,N_7437);
or U7916 (N_7916,N_7451,N_7489);
nand U7917 (N_7917,N_7252,N_7350);
nand U7918 (N_7918,N_7137,N_7375);
xnor U7919 (N_7919,N_7368,N_7447);
nand U7920 (N_7920,N_7123,N_7475);
or U7921 (N_7921,N_7042,N_7163);
nor U7922 (N_7922,N_7406,N_7187);
and U7923 (N_7923,N_7099,N_7042);
nor U7924 (N_7924,N_7156,N_7210);
nor U7925 (N_7925,N_7220,N_7281);
nor U7926 (N_7926,N_7484,N_7049);
or U7927 (N_7927,N_7474,N_7345);
or U7928 (N_7928,N_7139,N_7467);
and U7929 (N_7929,N_7398,N_7055);
and U7930 (N_7930,N_7072,N_7405);
nor U7931 (N_7931,N_7093,N_7198);
nor U7932 (N_7932,N_7282,N_7301);
nand U7933 (N_7933,N_7021,N_7191);
and U7934 (N_7934,N_7421,N_7053);
and U7935 (N_7935,N_7327,N_7145);
nand U7936 (N_7936,N_7474,N_7414);
nand U7937 (N_7937,N_7346,N_7493);
nand U7938 (N_7938,N_7232,N_7016);
and U7939 (N_7939,N_7454,N_7219);
or U7940 (N_7940,N_7246,N_7447);
and U7941 (N_7941,N_7067,N_7357);
and U7942 (N_7942,N_7321,N_7263);
xnor U7943 (N_7943,N_7032,N_7028);
or U7944 (N_7944,N_7041,N_7266);
nor U7945 (N_7945,N_7369,N_7224);
nand U7946 (N_7946,N_7144,N_7181);
or U7947 (N_7947,N_7312,N_7446);
nand U7948 (N_7948,N_7491,N_7121);
or U7949 (N_7949,N_7034,N_7358);
and U7950 (N_7950,N_7099,N_7052);
nor U7951 (N_7951,N_7117,N_7377);
nor U7952 (N_7952,N_7262,N_7291);
nand U7953 (N_7953,N_7309,N_7017);
nor U7954 (N_7954,N_7243,N_7327);
or U7955 (N_7955,N_7424,N_7034);
and U7956 (N_7956,N_7282,N_7347);
nand U7957 (N_7957,N_7355,N_7177);
or U7958 (N_7958,N_7122,N_7264);
nor U7959 (N_7959,N_7251,N_7339);
nor U7960 (N_7960,N_7061,N_7111);
nand U7961 (N_7961,N_7140,N_7318);
nand U7962 (N_7962,N_7339,N_7408);
and U7963 (N_7963,N_7458,N_7448);
nor U7964 (N_7964,N_7101,N_7338);
and U7965 (N_7965,N_7326,N_7202);
nor U7966 (N_7966,N_7313,N_7143);
nor U7967 (N_7967,N_7494,N_7322);
nand U7968 (N_7968,N_7399,N_7364);
nor U7969 (N_7969,N_7408,N_7442);
nor U7970 (N_7970,N_7346,N_7349);
nor U7971 (N_7971,N_7251,N_7344);
nor U7972 (N_7972,N_7467,N_7361);
and U7973 (N_7973,N_7335,N_7191);
nand U7974 (N_7974,N_7420,N_7324);
or U7975 (N_7975,N_7492,N_7432);
nor U7976 (N_7976,N_7028,N_7402);
or U7977 (N_7977,N_7058,N_7179);
and U7978 (N_7978,N_7319,N_7363);
and U7979 (N_7979,N_7035,N_7151);
nand U7980 (N_7980,N_7285,N_7405);
or U7981 (N_7981,N_7066,N_7318);
and U7982 (N_7982,N_7352,N_7222);
nand U7983 (N_7983,N_7135,N_7197);
or U7984 (N_7984,N_7370,N_7182);
nor U7985 (N_7985,N_7113,N_7266);
and U7986 (N_7986,N_7035,N_7492);
and U7987 (N_7987,N_7003,N_7384);
or U7988 (N_7988,N_7439,N_7295);
nor U7989 (N_7989,N_7428,N_7325);
nand U7990 (N_7990,N_7215,N_7104);
nor U7991 (N_7991,N_7259,N_7151);
nand U7992 (N_7992,N_7482,N_7402);
nand U7993 (N_7993,N_7085,N_7013);
or U7994 (N_7994,N_7188,N_7480);
and U7995 (N_7995,N_7026,N_7221);
or U7996 (N_7996,N_7025,N_7194);
nor U7997 (N_7997,N_7283,N_7293);
nand U7998 (N_7998,N_7308,N_7045);
nor U7999 (N_7999,N_7441,N_7173);
nor U8000 (N_8000,N_7606,N_7645);
and U8001 (N_8001,N_7509,N_7886);
nand U8002 (N_8002,N_7637,N_7848);
and U8003 (N_8003,N_7635,N_7858);
or U8004 (N_8004,N_7955,N_7535);
or U8005 (N_8005,N_7881,N_7783);
nand U8006 (N_8006,N_7945,N_7786);
or U8007 (N_8007,N_7524,N_7734);
nor U8008 (N_8008,N_7701,N_7632);
nor U8009 (N_8009,N_7984,N_7918);
nor U8010 (N_8010,N_7878,N_7800);
or U8011 (N_8011,N_7915,N_7827);
nand U8012 (N_8012,N_7767,N_7964);
or U8013 (N_8013,N_7591,N_7538);
xor U8014 (N_8014,N_7845,N_7888);
nor U8015 (N_8015,N_7722,N_7624);
nand U8016 (N_8016,N_7693,N_7705);
or U8017 (N_8017,N_7846,N_7715);
or U8018 (N_8018,N_7641,N_7612);
or U8019 (N_8019,N_7916,N_7738);
and U8020 (N_8020,N_7500,N_7691);
nor U8021 (N_8021,N_7835,N_7853);
nand U8022 (N_8022,N_7579,N_7811);
nor U8023 (N_8023,N_7920,N_7829);
nor U8024 (N_8024,N_7912,N_7669);
and U8025 (N_8025,N_7826,N_7904);
nor U8026 (N_8026,N_7993,N_7690);
nand U8027 (N_8027,N_7566,N_7539);
nor U8028 (N_8028,N_7860,N_7562);
nand U8029 (N_8029,N_7609,N_7717);
nor U8030 (N_8030,N_7563,N_7925);
nor U8031 (N_8031,N_7949,N_7678);
or U8032 (N_8032,N_7565,N_7516);
nand U8033 (N_8033,N_7699,N_7662);
nor U8034 (N_8034,N_7531,N_7590);
nor U8035 (N_8035,N_7607,N_7792);
nor U8036 (N_8036,N_7697,N_7782);
or U8037 (N_8037,N_7757,N_7601);
nand U8038 (N_8038,N_7766,N_7922);
nor U8039 (N_8039,N_7906,N_7968);
xor U8040 (N_8040,N_7659,N_7657);
nand U8041 (N_8041,N_7504,N_7997);
and U8042 (N_8042,N_7751,N_7876);
and U8043 (N_8043,N_7967,N_7506);
and U8044 (N_8044,N_7961,N_7864);
nand U8045 (N_8045,N_7508,N_7684);
nor U8046 (N_8046,N_7700,N_7573);
and U8047 (N_8047,N_7948,N_7541);
nand U8048 (N_8048,N_7520,N_7986);
or U8049 (N_8049,N_7615,N_7581);
or U8050 (N_8050,N_7973,N_7899);
nor U8051 (N_8051,N_7661,N_7988);
and U8052 (N_8052,N_7947,N_7614);
nand U8053 (N_8053,N_7586,N_7726);
nand U8054 (N_8054,N_7765,N_7784);
nor U8055 (N_8055,N_7851,N_7577);
nor U8056 (N_8056,N_7672,N_7771);
and U8057 (N_8057,N_7935,N_7849);
nand U8058 (N_8058,N_7901,N_7958);
and U8059 (N_8059,N_7698,N_7894);
nor U8060 (N_8060,N_7911,N_7668);
and U8061 (N_8061,N_7514,N_7806);
nand U8062 (N_8062,N_7503,N_7527);
or U8063 (N_8063,N_7626,N_7560);
or U8064 (N_8064,N_7869,N_7789);
or U8065 (N_8065,N_7640,N_7707);
nand U8066 (N_8066,N_7813,N_7622);
nand U8067 (N_8067,N_7728,N_7873);
or U8068 (N_8068,N_7528,N_7764);
nor U8069 (N_8069,N_7561,N_7512);
nand U8070 (N_8070,N_7544,N_7822);
nor U8071 (N_8071,N_7913,N_7970);
or U8072 (N_8072,N_7580,N_7628);
and U8073 (N_8073,N_7854,N_7694);
and U8074 (N_8074,N_7564,N_7688);
nor U8075 (N_8075,N_7518,N_7570);
or U8076 (N_8076,N_7996,N_7642);
xor U8077 (N_8077,N_7630,N_7517);
nor U8078 (N_8078,N_7594,N_7865);
and U8079 (N_8079,N_7725,N_7852);
xnor U8080 (N_8080,N_7529,N_7938);
xnor U8081 (N_8081,N_7875,N_7588);
or U8082 (N_8082,N_7867,N_7638);
nand U8083 (N_8083,N_7831,N_7521);
and U8084 (N_8084,N_7569,N_7934);
nor U8085 (N_8085,N_7999,N_7763);
nor U8086 (N_8086,N_7554,N_7990);
or U8087 (N_8087,N_7674,N_7952);
and U8088 (N_8088,N_7617,N_7780);
nand U8089 (N_8089,N_7709,N_7941);
nor U8090 (N_8090,N_7675,N_7507);
and U8091 (N_8091,N_7761,N_7682);
and U8092 (N_8092,N_7686,N_7957);
or U8093 (N_8093,N_7549,N_7572);
or U8094 (N_8094,N_7917,N_7823);
and U8095 (N_8095,N_7908,N_7924);
and U8096 (N_8096,N_7543,N_7724);
and U8097 (N_8097,N_7729,N_7832);
xnor U8098 (N_8098,N_7596,N_7787);
nand U8099 (N_8099,N_7712,N_7744);
nor U8100 (N_8100,N_7863,N_7850);
and U8101 (N_8101,N_7898,N_7903);
nor U8102 (N_8102,N_7511,N_7711);
nand U8103 (N_8103,N_7695,N_7627);
and U8104 (N_8104,N_7611,N_7872);
nand U8105 (N_8105,N_7733,N_7663);
and U8106 (N_8106,N_7805,N_7946);
nor U8107 (N_8107,N_7812,N_7855);
nand U8108 (N_8108,N_7798,N_7629);
and U8109 (N_8109,N_7773,N_7959);
or U8110 (N_8110,N_7862,N_7929);
nand U8111 (N_8111,N_7943,N_7884);
nand U8112 (N_8112,N_7992,N_7731);
nand U8113 (N_8113,N_7870,N_7779);
or U8114 (N_8114,N_7874,N_7809);
and U8115 (N_8115,N_7856,N_7623);
and U8116 (N_8116,N_7537,N_7654);
or U8117 (N_8117,N_7589,N_7652);
or U8118 (N_8118,N_7753,N_7793);
and U8119 (N_8119,N_7769,N_7533);
nand U8120 (N_8120,N_7840,N_7818);
and U8121 (N_8121,N_7892,N_7583);
nor U8122 (N_8122,N_7866,N_7844);
or U8123 (N_8123,N_7571,N_7593);
and U8124 (N_8124,N_7585,N_7972);
or U8125 (N_8125,N_7976,N_7987);
or U8126 (N_8126,N_7746,N_7759);
nor U8127 (N_8127,N_7551,N_7721);
xnor U8128 (N_8128,N_7807,N_7679);
and U8129 (N_8129,N_7825,N_7745);
and U8130 (N_8130,N_7727,N_7940);
or U8131 (N_8131,N_7556,N_7696);
nand U8132 (N_8132,N_7592,N_7755);
and U8133 (N_8133,N_7743,N_7859);
and U8134 (N_8134,N_7879,N_7975);
and U8135 (N_8135,N_7555,N_7921);
nand U8136 (N_8136,N_7814,N_7680);
or U8137 (N_8137,N_7983,N_7553);
and U8138 (N_8138,N_7877,N_7932);
nand U8139 (N_8139,N_7871,N_7616);
xnor U8140 (N_8140,N_7954,N_7605);
or U8141 (N_8141,N_7720,N_7736);
or U8142 (N_8142,N_7909,N_7923);
nor U8143 (N_8143,N_7708,N_7651);
nor U8144 (N_8144,N_7836,N_7971);
nand U8145 (N_8145,N_7716,N_7742);
or U8146 (N_8146,N_7597,N_7737);
and U8147 (N_8147,N_7534,N_7880);
and U8148 (N_8148,N_7927,N_7634);
nor U8149 (N_8149,N_7857,N_7703);
nand U8150 (N_8150,N_7683,N_7677);
nand U8151 (N_8151,N_7890,N_7781);
and U8152 (N_8152,N_7978,N_7648);
or U8153 (N_8153,N_7833,N_7584);
and U8154 (N_8154,N_7969,N_7750);
nor U8155 (N_8155,N_7895,N_7953);
nand U8156 (N_8156,N_7791,N_7778);
and U8157 (N_8157,N_7545,N_7749);
and U8158 (N_8158,N_7574,N_7723);
and U8159 (N_8159,N_7599,N_7974);
nor U8160 (N_8160,N_7681,N_7576);
nand U8161 (N_8161,N_7900,N_7944);
and U8162 (N_8162,N_7965,N_7525);
nor U8163 (N_8163,N_7519,N_7557);
and U8164 (N_8164,N_7982,N_7804);
or U8165 (N_8165,N_7928,N_7713);
and U8166 (N_8166,N_7802,N_7803);
nor U8167 (N_8167,N_7603,N_7931);
nand U8168 (N_8168,N_7550,N_7604);
nand U8169 (N_8169,N_7515,N_7808);
and U8170 (N_8170,N_7788,N_7891);
and U8171 (N_8171,N_7981,N_7885);
or U8172 (N_8172,N_7673,N_7977);
xor U8173 (N_8173,N_7625,N_7548);
or U8174 (N_8174,N_7559,N_7687);
or U8175 (N_8175,N_7747,N_7660);
or U8176 (N_8176,N_7608,N_7790);
and U8177 (N_8177,N_7810,N_7770);
nand U8178 (N_8178,N_7618,N_7735);
nor U8179 (N_8179,N_7905,N_7530);
or U8180 (N_8180,N_7842,N_7893);
nand U8181 (N_8181,N_7619,N_7794);
xnor U8182 (N_8182,N_7513,N_7760);
nor U8183 (N_8183,N_7649,N_7636);
or U8184 (N_8184,N_7546,N_7897);
nor U8185 (N_8185,N_7685,N_7998);
nand U8186 (N_8186,N_7985,N_7774);
nor U8187 (N_8187,N_7646,N_7882);
and U8188 (N_8188,N_7631,N_7739);
or U8189 (N_8189,N_7671,N_7939);
nor U8190 (N_8190,N_7838,N_7772);
and U8191 (N_8191,N_7843,N_7796);
nor U8192 (N_8192,N_7621,N_7960);
nor U8193 (N_8193,N_7536,N_7595);
nand U8194 (N_8194,N_7505,N_7989);
nand U8195 (N_8195,N_7658,N_7667);
and U8196 (N_8196,N_7502,N_7956);
or U8197 (N_8197,N_7839,N_7552);
or U8198 (N_8198,N_7748,N_7828);
nor U8199 (N_8199,N_7542,N_7785);
nand U8200 (N_8200,N_7666,N_7587);
or U8201 (N_8201,N_7837,N_7647);
nor U8202 (N_8202,N_7962,N_7610);
nor U8203 (N_8203,N_7820,N_7644);
or U8204 (N_8204,N_7752,N_7602);
xnor U8205 (N_8205,N_7933,N_7706);
nand U8206 (N_8206,N_7994,N_7719);
and U8207 (N_8207,N_7653,N_7942);
nor U8208 (N_8208,N_7834,N_7966);
or U8209 (N_8209,N_7861,N_7526);
and U8210 (N_8210,N_7643,N_7775);
or U8211 (N_8211,N_7914,N_7979);
or U8212 (N_8212,N_7664,N_7741);
or U8213 (N_8213,N_7902,N_7797);
nor U8214 (N_8214,N_7633,N_7830);
nand U8215 (N_8215,N_7676,N_7926);
nand U8216 (N_8216,N_7910,N_7639);
or U8217 (N_8217,N_7930,N_7689);
and U8218 (N_8218,N_7995,N_7919);
nand U8219 (N_8219,N_7501,N_7883);
nor U8220 (N_8220,N_7991,N_7575);
and U8221 (N_8221,N_7522,N_7523);
nand U8222 (N_8222,N_7754,N_7817);
and U8223 (N_8223,N_7704,N_7718);
nand U8224 (N_8224,N_7510,N_7889);
nor U8225 (N_8225,N_7714,N_7578);
nand U8226 (N_8226,N_7540,N_7887);
nand U8227 (N_8227,N_7656,N_7702);
and U8228 (N_8228,N_7730,N_7532);
nand U8229 (N_8229,N_7650,N_7547);
xor U8230 (N_8230,N_7758,N_7868);
or U8231 (N_8231,N_7582,N_7777);
nor U8232 (N_8232,N_7598,N_7620);
nor U8233 (N_8233,N_7568,N_7801);
or U8234 (N_8234,N_7950,N_7655);
xnor U8235 (N_8235,N_7710,N_7768);
or U8236 (N_8236,N_7762,N_7567);
or U8237 (N_8237,N_7740,N_7670);
and U8238 (N_8238,N_7600,N_7756);
and U8239 (N_8239,N_7980,N_7819);
and U8240 (N_8240,N_7732,N_7776);
and U8241 (N_8241,N_7558,N_7847);
and U8242 (N_8242,N_7799,N_7936);
nand U8243 (N_8243,N_7815,N_7665);
nand U8244 (N_8244,N_7951,N_7613);
and U8245 (N_8245,N_7937,N_7896);
or U8246 (N_8246,N_7692,N_7824);
or U8247 (N_8247,N_7821,N_7907);
or U8248 (N_8248,N_7841,N_7795);
nor U8249 (N_8249,N_7816,N_7963);
nor U8250 (N_8250,N_7952,N_7998);
nor U8251 (N_8251,N_7950,N_7547);
or U8252 (N_8252,N_7735,N_7696);
nand U8253 (N_8253,N_7902,N_7601);
or U8254 (N_8254,N_7532,N_7926);
or U8255 (N_8255,N_7975,N_7793);
or U8256 (N_8256,N_7570,N_7828);
and U8257 (N_8257,N_7796,N_7668);
and U8258 (N_8258,N_7555,N_7525);
nor U8259 (N_8259,N_7995,N_7822);
nand U8260 (N_8260,N_7917,N_7886);
or U8261 (N_8261,N_7820,N_7767);
or U8262 (N_8262,N_7607,N_7525);
or U8263 (N_8263,N_7525,N_7818);
or U8264 (N_8264,N_7867,N_7946);
and U8265 (N_8265,N_7790,N_7547);
or U8266 (N_8266,N_7634,N_7834);
nor U8267 (N_8267,N_7746,N_7665);
and U8268 (N_8268,N_7916,N_7620);
nand U8269 (N_8269,N_7781,N_7559);
and U8270 (N_8270,N_7947,N_7845);
or U8271 (N_8271,N_7904,N_7810);
nand U8272 (N_8272,N_7979,N_7931);
and U8273 (N_8273,N_7520,N_7900);
and U8274 (N_8274,N_7781,N_7690);
and U8275 (N_8275,N_7601,N_7503);
or U8276 (N_8276,N_7704,N_7586);
nand U8277 (N_8277,N_7545,N_7637);
nor U8278 (N_8278,N_7708,N_7818);
nor U8279 (N_8279,N_7835,N_7936);
xnor U8280 (N_8280,N_7848,N_7685);
or U8281 (N_8281,N_7554,N_7689);
xor U8282 (N_8282,N_7645,N_7947);
nand U8283 (N_8283,N_7971,N_7662);
and U8284 (N_8284,N_7635,N_7676);
or U8285 (N_8285,N_7797,N_7784);
and U8286 (N_8286,N_7959,N_7819);
nand U8287 (N_8287,N_7724,N_7757);
and U8288 (N_8288,N_7826,N_7936);
and U8289 (N_8289,N_7797,N_7729);
nand U8290 (N_8290,N_7535,N_7930);
nor U8291 (N_8291,N_7699,N_7900);
or U8292 (N_8292,N_7874,N_7638);
nand U8293 (N_8293,N_7811,N_7938);
nand U8294 (N_8294,N_7787,N_7851);
nor U8295 (N_8295,N_7980,N_7673);
and U8296 (N_8296,N_7546,N_7502);
nand U8297 (N_8297,N_7883,N_7711);
or U8298 (N_8298,N_7640,N_7578);
nand U8299 (N_8299,N_7823,N_7974);
and U8300 (N_8300,N_7887,N_7712);
or U8301 (N_8301,N_7655,N_7938);
or U8302 (N_8302,N_7948,N_7999);
nand U8303 (N_8303,N_7849,N_7515);
or U8304 (N_8304,N_7637,N_7964);
xnor U8305 (N_8305,N_7544,N_7517);
and U8306 (N_8306,N_7519,N_7587);
or U8307 (N_8307,N_7735,N_7795);
nand U8308 (N_8308,N_7898,N_7911);
nand U8309 (N_8309,N_7774,N_7734);
and U8310 (N_8310,N_7844,N_7667);
nor U8311 (N_8311,N_7876,N_7960);
or U8312 (N_8312,N_7788,N_7962);
or U8313 (N_8313,N_7867,N_7988);
or U8314 (N_8314,N_7868,N_7872);
xor U8315 (N_8315,N_7563,N_7986);
and U8316 (N_8316,N_7825,N_7893);
or U8317 (N_8317,N_7823,N_7695);
and U8318 (N_8318,N_7808,N_7763);
nand U8319 (N_8319,N_7964,N_7822);
nor U8320 (N_8320,N_7882,N_7857);
nand U8321 (N_8321,N_7541,N_7868);
or U8322 (N_8322,N_7978,N_7723);
and U8323 (N_8323,N_7537,N_7878);
or U8324 (N_8324,N_7784,N_7910);
or U8325 (N_8325,N_7624,N_7581);
or U8326 (N_8326,N_7878,N_7583);
nand U8327 (N_8327,N_7549,N_7770);
and U8328 (N_8328,N_7758,N_7763);
and U8329 (N_8329,N_7889,N_7896);
and U8330 (N_8330,N_7847,N_7882);
nor U8331 (N_8331,N_7838,N_7706);
nor U8332 (N_8332,N_7666,N_7767);
nand U8333 (N_8333,N_7560,N_7619);
or U8334 (N_8334,N_7959,N_7693);
nor U8335 (N_8335,N_7855,N_7813);
and U8336 (N_8336,N_7913,N_7790);
and U8337 (N_8337,N_7943,N_7625);
nor U8338 (N_8338,N_7525,N_7846);
nand U8339 (N_8339,N_7593,N_7924);
nor U8340 (N_8340,N_7598,N_7885);
nor U8341 (N_8341,N_7776,N_7970);
or U8342 (N_8342,N_7668,N_7798);
or U8343 (N_8343,N_7542,N_7694);
nor U8344 (N_8344,N_7636,N_7507);
nor U8345 (N_8345,N_7998,N_7948);
and U8346 (N_8346,N_7821,N_7665);
nor U8347 (N_8347,N_7850,N_7639);
nand U8348 (N_8348,N_7806,N_7601);
nand U8349 (N_8349,N_7700,N_7972);
and U8350 (N_8350,N_7526,N_7596);
or U8351 (N_8351,N_7931,N_7719);
or U8352 (N_8352,N_7526,N_7724);
or U8353 (N_8353,N_7737,N_7541);
nand U8354 (N_8354,N_7733,N_7890);
or U8355 (N_8355,N_7595,N_7770);
or U8356 (N_8356,N_7774,N_7581);
nor U8357 (N_8357,N_7889,N_7712);
and U8358 (N_8358,N_7548,N_7951);
nand U8359 (N_8359,N_7954,N_7882);
nand U8360 (N_8360,N_7573,N_7752);
or U8361 (N_8361,N_7611,N_7677);
or U8362 (N_8362,N_7678,N_7710);
nor U8363 (N_8363,N_7835,N_7678);
or U8364 (N_8364,N_7523,N_7767);
and U8365 (N_8365,N_7534,N_7798);
nand U8366 (N_8366,N_7996,N_7769);
xor U8367 (N_8367,N_7507,N_7776);
and U8368 (N_8368,N_7964,N_7589);
and U8369 (N_8369,N_7808,N_7526);
nor U8370 (N_8370,N_7992,N_7793);
and U8371 (N_8371,N_7681,N_7731);
or U8372 (N_8372,N_7968,N_7501);
and U8373 (N_8373,N_7635,N_7963);
xor U8374 (N_8374,N_7598,N_7652);
or U8375 (N_8375,N_7873,N_7634);
nor U8376 (N_8376,N_7999,N_7587);
nand U8377 (N_8377,N_7904,N_7720);
or U8378 (N_8378,N_7782,N_7596);
and U8379 (N_8379,N_7850,N_7984);
and U8380 (N_8380,N_7908,N_7518);
and U8381 (N_8381,N_7740,N_7870);
or U8382 (N_8382,N_7668,N_7526);
nand U8383 (N_8383,N_7651,N_7803);
and U8384 (N_8384,N_7947,N_7967);
nor U8385 (N_8385,N_7660,N_7997);
nor U8386 (N_8386,N_7832,N_7751);
and U8387 (N_8387,N_7886,N_7981);
or U8388 (N_8388,N_7912,N_7858);
nor U8389 (N_8389,N_7712,N_7789);
and U8390 (N_8390,N_7708,N_7521);
nor U8391 (N_8391,N_7525,N_7580);
or U8392 (N_8392,N_7723,N_7666);
nand U8393 (N_8393,N_7883,N_7815);
xnor U8394 (N_8394,N_7679,N_7764);
nand U8395 (N_8395,N_7890,N_7647);
or U8396 (N_8396,N_7649,N_7863);
nor U8397 (N_8397,N_7567,N_7898);
nor U8398 (N_8398,N_7757,N_7557);
nand U8399 (N_8399,N_7782,N_7568);
nand U8400 (N_8400,N_7998,N_7518);
or U8401 (N_8401,N_7899,N_7866);
or U8402 (N_8402,N_7547,N_7761);
nand U8403 (N_8403,N_7705,N_7586);
nor U8404 (N_8404,N_7925,N_7720);
nor U8405 (N_8405,N_7728,N_7609);
nor U8406 (N_8406,N_7943,N_7725);
nand U8407 (N_8407,N_7679,N_7951);
nor U8408 (N_8408,N_7870,N_7644);
nor U8409 (N_8409,N_7869,N_7610);
nand U8410 (N_8410,N_7784,N_7643);
or U8411 (N_8411,N_7908,N_7742);
nand U8412 (N_8412,N_7814,N_7941);
nor U8413 (N_8413,N_7625,N_7788);
or U8414 (N_8414,N_7558,N_7636);
nand U8415 (N_8415,N_7644,N_7668);
and U8416 (N_8416,N_7681,N_7775);
nand U8417 (N_8417,N_7989,N_7831);
and U8418 (N_8418,N_7853,N_7686);
or U8419 (N_8419,N_7956,N_7663);
nor U8420 (N_8420,N_7519,N_7949);
nor U8421 (N_8421,N_7844,N_7917);
or U8422 (N_8422,N_7681,N_7570);
nand U8423 (N_8423,N_7522,N_7609);
nand U8424 (N_8424,N_7867,N_7885);
and U8425 (N_8425,N_7847,N_7701);
nand U8426 (N_8426,N_7994,N_7850);
nor U8427 (N_8427,N_7871,N_7700);
nor U8428 (N_8428,N_7695,N_7870);
nor U8429 (N_8429,N_7821,N_7521);
or U8430 (N_8430,N_7991,N_7566);
or U8431 (N_8431,N_7800,N_7647);
or U8432 (N_8432,N_7945,N_7727);
nand U8433 (N_8433,N_7750,N_7799);
nand U8434 (N_8434,N_7649,N_7686);
and U8435 (N_8435,N_7684,N_7878);
nand U8436 (N_8436,N_7617,N_7867);
nand U8437 (N_8437,N_7817,N_7779);
nand U8438 (N_8438,N_7595,N_7604);
nand U8439 (N_8439,N_7752,N_7850);
nor U8440 (N_8440,N_7943,N_7540);
or U8441 (N_8441,N_7918,N_7601);
nor U8442 (N_8442,N_7554,N_7595);
nor U8443 (N_8443,N_7953,N_7888);
nor U8444 (N_8444,N_7775,N_7610);
nor U8445 (N_8445,N_7782,N_7681);
or U8446 (N_8446,N_7650,N_7518);
and U8447 (N_8447,N_7676,N_7565);
nand U8448 (N_8448,N_7632,N_7744);
nand U8449 (N_8449,N_7907,N_7632);
and U8450 (N_8450,N_7602,N_7873);
or U8451 (N_8451,N_7606,N_7728);
and U8452 (N_8452,N_7705,N_7841);
and U8453 (N_8453,N_7758,N_7605);
nand U8454 (N_8454,N_7885,N_7613);
xnor U8455 (N_8455,N_7946,N_7793);
nand U8456 (N_8456,N_7536,N_7577);
nand U8457 (N_8457,N_7651,N_7952);
and U8458 (N_8458,N_7751,N_7542);
nand U8459 (N_8459,N_7721,N_7808);
nand U8460 (N_8460,N_7691,N_7885);
or U8461 (N_8461,N_7797,N_7999);
nor U8462 (N_8462,N_7753,N_7922);
nor U8463 (N_8463,N_7799,N_7972);
nand U8464 (N_8464,N_7901,N_7623);
nand U8465 (N_8465,N_7607,N_7773);
and U8466 (N_8466,N_7685,N_7978);
nand U8467 (N_8467,N_7554,N_7763);
nand U8468 (N_8468,N_7781,N_7681);
or U8469 (N_8469,N_7602,N_7882);
and U8470 (N_8470,N_7790,N_7761);
nor U8471 (N_8471,N_7794,N_7730);
and U8472 (N_8472,N_7975,N_7541);
or U8473 (N_8473,N_7720,N_7687);
or U8474 (N_8474,N_7988,N_7694);
nor U8475 (N_8475,N_7930,N_7909);
nor U8476 (N_8476,N_7704,N_7833);
and U8477 (N_8477,N_7667,N_7792);
and U8478 (N_8478,N_7658,N_7604);
and U8479 (N_8479,N_7966,N_7645);
xor U8480 (N_8480,N_7967,N_7998);
nor U8481 (N_8481,N_7853,N_7760);
or U8482 (N_8482,N_7921,N_7825);
nor U8483 (N_8483,N_7831,N_7615);
or U8484 (N_8484,N_7941,N_7500);
or U8485 (N_8485,N_7730,N_7799);
nand U8486 (N_8486,N_7980,N_7816);
and U8487 (N_8487,N_7983,N_7863);
nand U8488 (N_8488,N_7965,N_7709);
and U8489 (N_8489,N_7657,N_7943);
nand U8490 (N_8490,N_7697,N_7824);
and U8491 (N_8491,N_7826,N_7909);
nor U8492 (N_8492,N_7563,N_7714);
and U8493 (N_8493,N_7930,N_7502);
and U8494 (N_8494,N_7963,N_7505);
nand U8495 (N_8495,N_7536,N_7872);
nor U8496 (N_8496,N_7705,N_7536);
nand U8497 (N_8497,N_7605,N_7858);
nor U8498 (N_8498,N_7900,N_7516);
and U8499 (N_8499,N_7733,N_7655);
nand U8500 (N_8500,N_8118,N_8328);
and U8501 (N_8501,N_8497,N_8481);
nor U8502 (N_8502,N_8198,N_8058);
nor U8503 (N_8503,N_8249,N_8094);
or U8504 (N_8504,N_8248,N_8212);
nor U8505 (N_8505,N_8342,N_8359);
nand U8506 (N_8506,N_8136,N_8037);
nor U8507 (N_8507,N_8370,N_8150);
or U8508 (N_8508,N_8146,N_8012);
and U8509 (N_8509,N_8394,N_8221);
nand U8510 (N_8510,N_8385,N_8326);
nor U8511 (N_8511,N_8382,N_8015);
and U8512 (N_8512,N_8308,N_8285);
or U8513 (N_8513,N_8369,N_8262);
and U8514 (N_8514,N_8304,N_8000);
and U8515 (N_8515,N_8440,N_8296);
or U8516 (N_8516,N_8353,N_8086);
nand U8517 (N_8517,N_8106,N_8111);
nor U8518 (N_8518,N_8235,N_8048);
nand U8519 (N_8519,N_8386,N_8241);
or U8520 (N_8520,N_8314,N_8339);
nor U8521 (N_8521,N_8350,N_8341);
and U8522 (N_8522,N_8306,N_8310);
nand U8523 (N_8523,N_8083,N_8471);
nor U8524 (N_8524,N_8056,N_8054);
and U8525 (N_8525,N_8287,N_8226);
and U8526 (N_8526,N_8464,N_8280);
and U8527 (N_8527,N_8158,N_8329);
or U8528 (N_8528,N_8364,N_8484);
nand U8529 (N_8529,N_8202,N_8438);
and U8530 (N_8530,N_8265,N_8052);
nor U8531 (N_8531,N_8008,N_8121);
nor U8532 (N_8532,N_8028,N_8185);
or U8533 (N_8533,N_8113,N_8416);
and U8534 (N_8534,N_8013,N_8325);
nor U8535 (N_8535,N_8026,N_8264);
and U8536 (N_8536,N_8465,N_8195);
or U8537 (N_8537,N_8096,N_8070);
nand U8538 (N_8538,N_8009,N_8422);
nor U8539 (N_8539,N_8401,N_8286);
xnor U8540 (N_8540,N_8311,N_8356);
and U8541 (N_8541,N_8489,N_8301);
nor U8542 (N_8542,N_8239,N_8205);
nand U8543 (N_8543,N_8003,N_8403);
nand U8544 (N_8544,N_8063,N_8294);
or U8545 (N_8545,N_8457,N_8035);
nand U8546 (N_8546,N_8055,N_8479);
or U8547 (N_8547,N_8454,N_8429);
and U8548 (N_8548,N_8125,N_8320);
xor U8549 (N_8549,N_8192,N_8477);
nand U8550 (N_8550,N_8418,N_8174);
and U8551 (N_8551,N_8298,N_8042);
nand U8552 (N_8552,N_8345,N_8159);
or U8553 (N_8553,N_8321,N_8162);
nor U8554 (N_8554,N_8421,N_8223);
or U8555 (N_8555,N_8439,N_8188);
or U8556 (N_8556,N_8152,N_8095);
nor U8557 (N_8557,N_8098,N_8045);
and U8558 (N_8558,N_8040,N_8128);
nor U8559 (N_8559,N_8216,N_8177);
and U8560 (N_8560,N_8127,N_8087);
and U8561 (N_8561,N_8130,N_8145);
or U8562 (N_8562,N_8378,N_8398);
nor U8563 (N_8563,N_8039,N_8024);
nand U8564 (N_8564,N_8148,N_8209);
and U8565 (N_8565,N_8181,N_8332);
and U8566 (N_8566,N_8272,N_8362);
nand U8567 (N_8567,N_8044,N_8103);
or U8568 (N_8568,N_8176,N_8186);
or U8569 (N_8569,N_8323,N_8441);
or U8570 (N_8570,N_8156,N_8315);
and U8571 (N_8571,N_8299,N_8388);
nor U8572 (N_8572,N_8112,N_8194);
nor U8573 (N_8573,N_8366,N_8279);
and U8574 (N_8574,N_8025,N_8290);
or U8575 (N_8575,N_8002,N_8090);
nand U8576 (N_8576,N_8049,N_8257);
or U8577 (N_8577,N_8317,N_8419);
nor U8578 (N_8578,N_8102,N_8448);
or U8579 (N_8579,N_8470,N_8069);
nor U8580 (N_8580,N_8007,N_8200);
xnor U8581 (N_8581,N_8004,N_8116);
nor U8582 (N_8582,N_8189,N_8447);
or U8583 (N_8583,N_8276,N_8021);
nor U8584 (N_8584,N_8230,N_8065);
or U8585 (N_8585,N_8201,N_8423);
nand U8586 (N_8586,N_8390,N_8085);
and U8587 (N_8587,N_8259,N_8377);
nand U8588 (N_8588,N_8089,N_8354);
or U8589 (N_8589,N_8051,N_8242);
and U8590 (N_8590,N_8488,N_8417);
nor U8591 (N_8591,N_8442,N_8316);
or U8592 (N_8592,N_8173,N_8478);
nand U8593 (N_8593,N_8164,N_8267);
nor U8594 (N_8594,N_8283,N_8074);
and U8595 (N_8595,N_8406,N_8413);
nor U8596 (N_8596,N_8224,N_8036);
nor U8597 (N_8597,N_8455,N_8046);
nor U8598 (N_8598,N_8238,N_8134);
or U8599 (N_8599,N_8319,N_8208);
and U8600 (N_8600,N_8031,N_8270);
and U8601 (N_8601,N_8172,N_8075);
nand U8602 (N_8602,N_8077,N_8081);
and U8603 (N_8603,N_8414,N_8180);
and U8604 (N_8604,N_8293,N_8435);
nand U8605 (N_8605,N_8142,N_8204);
nor U8606 (N_8606,N_8400,N_8494);
and U8607 (N_8607,N_8060,N_8459);
nand U8608 (N_8608,N_8193,N_8492);
and U8609 (N_8609,N_8227,N_8399);
nor U8610 (N_8610,N_8499,N_8255);
nor U8611 (N_8611,N_8466,N_8178);
nand U8612 (N_8612,N_8371,N_8260);
nor U8613 (N_8613,N_8425,N_8244);
and U8614 (N_8614,N_8302,N_8432);
and U8615 (N_8615,N_8225,N_8080);
or U8616 (N_8616,N_8473,N_8122);
nand U8617 (N_8617,N_8119,N_8073);
nor U8618 (N_8618,N_8105,N_8187);
or U8619 (N_8619,N_8171,N_8038);
or U8620 (N_8620,N_8082,N_8437);
nor U8621 (N_8621,N_8247,N_8402);
or U8622 (N_8622,N_8474,N_8360);
or U8623 (N_8623,N_8337,N_8047);
nand U8624 (N_8624,N_8289,N_8444);
and U8625 (N_8625,N_8236,N_8475);
nor U8626 (N_8626,N_8348,N_8335);
or U8627 (N_8627,N_8273,N_8263);
nor U8628 (N_8628,N_8232,N_8072);
nand U8629 (N_8629,N_8461,N_8424);
nand U8630 (N_8630,N_8100,N_8231);
and U8631 (N_8631,N_8214,N_8295);
nor U8632 (N_8632,N_8254,N_8436);
nand U8633 (N_8633,N_8109,N_8001);
or U8634 (N_8634,N_8071,N_8258);
nand U8635 (N_8635,N_8343,N_8114);
nor U8636 (N_8636,N_8373,N_8196);
and U8637 (N_8637,N_8281,N_8338);
nand U8638 (N_8638,N_8269,N_8154);
and U8639 (N_8639,N_8057,N_8020);
and U8640 (N_8640,N_8307,N_8284);
nor U8641 (N_8641,N_8117,N_8184);
or U8642 (N_8642,N_8483,N_8165);
and U8643 (N_8643,N_8210,N_8292);
nand U8644 (N_8644,N_8006,N_8218);
nand U8645 (N_8645,N_8110,N_8151);
or U8646 (N_8646,N_8068,N_8278);
or U8647 (N_8647,N_8389,N_8137);
nand U8648 (N_8648,N_8491,N_8374);
nand U8649 (N_8649,N_8076,N_8005);
nand U8650 (N_8650,N_8213,N_8139);
or U8651 (N_8651,N_8115,N_8415);
nand U8652 (N_8652,N_8309,N_8467);
or U8653 (N_8653,N_8357,N_8445);
nand U8654 (N_8654,N_8211,N_8271);
nor U8655 (N_8655,N_8407,N_8312);
and U8656 (N_8656,N_8496,N_8023);
or U8657 (N_8657,N_8014,N_8291);
or U8658 (N_8658,N_8027,N_8334);
nand U8659 (N_8659,N_8256,N_8222);
and U8660 (N_8660,N_8097,N_8160);
nand U8661 (N_8661,N_8372,N_8333);
nand U8662 (N_8662,N_8206,N_8404);
nand U8663 (N_8663,N_8300,N_8482);
and U8664 (N_8664,N_8099,N_8351);
nand U8665 (N_8665,N_8430,N_8228);
and U8666 (N_8666,N_8123,N_8199);
or U8667 (N_8667,N_8485,N_8380);
nand U8668 (N_8668,N_8059,N_8379);
nor U8669 (N_8669,N_8091,N_8412);
nand U8670 (N_8670,N_8234,N_8381);
nor U8671 (N_8671,N_8288,N_8183);
or U8672 (N_8672,N_8107,N_8088);
or U8673 (N_8673,N_8149,N_8463);
or U8674 (N_8674,N_8108,N_8450);
nand U8675 (N_8675,N_8084,N_8161);
or U8676 (N_8676,N_8062,N_8266);
or U8677 (N_8677,N_8392,N_8253);
nor U8678 (N_8678,N_8346,N_8361);
nand U8679 (N_8679,N_8324,N_8126);
and U8680 (N_8680,N_8397,N_8197);
nor U8681 (N_8681,N_8449,N_8066);
xor U8682 (N_8682,N_8147,N_8363);
xor U8683 (N_8683,N_8144,N_8458);
or U8684 (N_8684,N_8330,N_8219);
and U8685 (N_8685,N_8393,N_8443);
and U8686 (N_8686,N_8034,N_8453);
nand U8687 (N_8687,N_8019,N_8243);
nand U8688 (N_8688,N_8408,N_8168);
and U8689 (N_8689,N_8022,N_8451);
nand U8690 (N_8690,N_8480,N_8405);
nand U8691 (N_8691,N_8251,N_8383);
nand U8692 (N_8692,N_8349,N_8486);
nor U8693 (N_8693,N_8322,N_8433);
or U8694 (N_8694,N_8132,N_8033);
nor U8695 (N_8695,N_8093,N_8487);
or U8696 (N_8696,N_8141,N_8368);
nand U8697 (N_8697,N_8246,N_8409);
or U8698 (N_8698,N_8190,N_8133);
or U8699 (N_8699,N_8462,N_8017);
nand U8700 (N_8700,N_8395,N_8420);
nor U8701 (N_8701,N_8375,N_8428);
nor U8702 (N_8702,N_8367,N_8391);
and U8703 (N_8703,N_8153,N_8282);
and U8704 (N_8704,N_8365,N_8498);
and U8705 (N_8705,N_8240,N_8303);
nand U8706 (N_8706,N_8167,N_8041);
or U8707 (N_8707,N_8411,N_8138);
nor U8708 (N_8708,N_8166,N_8018);
nor U8709 (N_8709,N_8355,N_8426);
or U8710 (N_8710,N_8032,N_8469);
and U8711 (N_8711,N_8495,N_8434);
nor U8712 (N_8712,N_8163,N_8220);
nand U8713 (N_8713,N_8135,N_8313);
nand U8714 (N_8714,N_8237,N_8352);
nor U8715 (N_8715,N_8472,N_8446);
and U8716 (N_8716,N_8318,N_8336);
nor U8717 (N_8717,N_8120,N_8092);
nor U8718 (N_8718,N_8067,N_8233);
and U8719 (N_8719,N_8410,N_8157);
or U8720 (N_8720,N_8297,N_8305);
nand U8721 (N_8721,N_8140,N_8104);
and U8722 (N_8722,N_8468,N_8493);
nor U8723 (N_8723,N_8456,N_8053);
and U8724 (N_8724,N_8387,N_8061);
nand U8725 (N_8725,N_8175,N_8179);
nor U8726 (N_8726,N_8169,N_8016);
nand U8727 (N_8727,N_8131,N_8274);
nor U8728 (N_8728,N_8078,N_8396);
xnor U8729 (N_8729,N_8452,N_8064);
or U8730 (N_8730,N_8203,N_8384);
nor U8731 (N_8731,N_8431,N_8340);
nor U8732 (N_8732,N_8217,N_8011);
and U8733 (N_8733,N_8250,N_8182);
nand U8734 (N_8734,N_8155,N_8043);
and U8735 (N_8735,N_8460,N_8079);
xor U8736 (N_8736,N_8207,N_8215);
or U8737 (N_8737,N_8050,N_8358);
nand U8738 (N_8738,N_8490,N_8124);
nand U8739 (N_8739,N_8261,N_8275);
nand U8740 (N_8740,N_8029,N_8010);
nor U8741 (N_8741,N_8101,N_8170);
nand U8742 (N_8742,N_8347,N_8268);
xnor U8743 (N_8743,N_8191,N_8129);
xnor U8744 (N_8744,N_8252,N_8277);
nand U8745 (N_8745,N_8344,N_8327);
or U8746 (N_8746,N_8476,N_8427);
or U8747 (N_8747,N_8229,N_8030);
nor U8748 (N_8748,N_8245,N_8143);
and U8749 (N_8749,N_8376,N_8331);
nor U8750 (N_8750,N_8317,N_8319);
nor U8751 (N_8751,N_8028,N_8137);
or U8752 (N_8752,N_8424,N_8319);
nor U8753 (N_8753,N_8188,N_8058);
or U8754 (N_8754,N_8144,N_8478);
nand U8755 (N_8755,N_8273,N_8342);
or U8756 (N_8756,N_8020,N_8267);
and U8757 (N_8757,N_8168,N_8118);
and U8758 (N_8758,N_8463,N_8473);
nand U8759 (N_8759,N_8057,N_8244);
nor U8760 (N_8760,N_8475,N_8438);
nor U8761 (N_8761,N_8017,N_8333);
or U8762 (N_8762,N_8287,N_8196);
nand U8763 (N_8763,N_8456,N_8164);
and U8764 (N_8764,N_8403,N_8431);
nand U8765 (N_8765,N_8229,N_8460);
and U8766 (N_8766,N_8056,N_8442);
xnor U8767 (N_8767,N_8423,N_8318);
or U8768 (N_8768,N_8384,N_8411);
nor U8769 (N_8769,N_8379,N_8269);
and U8770 (N_8770,N_8217,N_8183);
nor U8771 (N_8771,N_8170,N_8225);
or U8772 (N_8772,N_8221,N_8025);
and U8773 (N_8773,N_8490,N_8443);
nand U8774 (N_8774,N_8487,N_8446);
nor U8775 (N_8775,N_8315,N_8016);
or U8776 (N_8776,N_8411,N_8494);
or U8777 (N_8777,N_8354,N_8370);
and U8778 (N_8778,N_8037,N_8427);
and U8779 (N_8779,N_8123,N_8226);
nand U8780 (N_8780,N_8022,N_8371);
and U8781 (N_8781,N_8092,N_8088);
and U8782 (N_8782,N_8007,N_8220);
and U8783 (N_8783,N_8251,N_8236);
nor U8784 (N_8784,N_8117,N_8487);
and U8785 (N_8785,N_8475,N_8375);
or U8786 (N_8786,N_8170,N_8486);
and U8787 (N_8787,N_8085,N_8445);
and U8788 (N_8788,N_8239,N_8353);
nor U8789 (N_8789,N_8330,N_8067);
nand U8790 (N_8790,N_8372,N_8158);
and U8791 (N_8791,N_8213,N_8294);
nor U8792 (N_8792,N_8374,N_8341);
or U8793 (N_8793,N_8281,N_8288);
or U8794 (N_8794,N_8342,N_8101);
nor U8795 (N_8795,N_8405,N_8102);
and U8796 (N_8796,N_8059,N_8305);
nor U8797 (N_8797,N_8312,N_8179);
and U8798 (N_8798,N_8101,N_8340);
nor U8799 (N_8799,N_8029,N_8378);
and U8800 (N_8800,N_8464,N_8328);
or U8801 (N_8801,N_8446,N_8426);
nor U8802 (N_8802,N_8051,N_8377);
nor U8803 (N_8803,N_8243,N_8247);
nand U8804 (N_8804,N_8119,N_8320);
nor U8805 (N_8805,N_8409,N_8299);
and U8806 (N_8806,N_8072,N_8265);
nor U8807 (N_8807,N_8329,N_8278);
nand U8808 (N_8808,N_8471,N_8171);
nor U8809 (N_8809,N_8059,N_8318);
nand U8810 (N_8810,N_8036,N_8120);
nand U8811 (N_8811,N_8331,N_8226);
or U8812 (N_8812,N_8079,N_8453);
nand U8813 (N_8813,N_8237,N_8075);
nor U8814 (N_8814,N_8306,N_8326);
nor U8815 (N_8815,N_8292,N_8455);
and U8816 (N_8816,N_8318,N_8023);
or U8817 (N_8817,N_8258,N_8436);
or U8818 (N_8818,N_8394,N_8458);
and U8819 (N_8819,N_8352,N_8185);
and U8820 (N_8820,N_8455,N_8364);
nand U8821 (N_8821,N_8337,N_8470);
nor U8822 (N_8822,N_8358,N_8034);
nand U8823 (N_8823,N_8435,N_8393);
and U8824 (N_8824,N_8004,N_8468);
nor U8825 (N_8825,N_8488,N_8137);
and U8826 (N_8826,N_8392,N_8226);
and U8827 (N_8827,N_8064,N_8422);
or U8828 (N_8828,N_8164,N_8259);
and U8829 (N_8829,N_8206,N_8382);
nand U8830 (N_8830,N_8339,N_8198);
or U8831 (N_8831,N_8287,N_8446);
and U8832 (N_8832,N_8267,N_8246);
or U8833 (N_8833,N_8484,N_8231);
nor U8834 (N_8834,N_8378,N_8226);
nand U8835 (N_8835,N_8398,N_8001);
or U8836 (N_8836,N_8172,N_8113);
nand U8837 (N_8837,N_8174,N_8364);
and U8838 (N_8838,N_8468,N_8255);
nand U8839 (N_8839,N_8027,N_8313);
or U8840 (N_8840,N_8075,N_8024);
and U8841 (N_8841,N_8064,N_8247);
nor U8842 (N_8842,N_8032,N_8383);
or U8843 (N_8843,N_8409,N_8272);
and U8844 (N_8844,N_8364,N_8413);
or U8845 (N_8845,N_8457,N_8025);
and U8846 (N_8846,N_8349,N_8286);
or U8847 (N_8847,N_8484,N_8088);
nand U8848 (N_8848,N_8030,N_8462);
xor U8849 (N_8849,N_8299,N_8116);
nand U8850 (N_8850,N_8103,N_8264);
xnor U8851 (N_8851,N_8247,N_8452);
nand U8852 (N_8852,N_8454,N_8186);
and U8853 (N_8853,N_8083,N_8123);
nand U8854 (N_8854,N_8034,N_8177);
nand U8855 (N_8855,N_8091,N_8025);
nand U8856 (N_8856,N_8278,N_8259);
or U8857 (N_8857,N_8319,N_8166);
nand U8858 (N_8858,N_8064,N_8248);
nor U8859 (N_8859,N_8214,N_8071);
and U8860 (N_8860,N_8270,N_8001);
nand U8861 (N_8861,N_8343,N_8411);
and U8862 (N_8862,N_8456,N_8172);
and U8863 (N_8863,N_8142,N_8140);
nand U8864 (N_8864,N_8473,N_8186);
or U8865 (N_8865,N_8126,N_8227);
nand U8866 (N_8866,N_8041,N_8455);
and U8867 (N_8867,N_8307,N_8410);
nor U8868 (N_8868,N_8092,N_8076);
or U8869 (N_8869,N_8298,N_8396);
nor U8870 (N_8870,N_8192,N_8464);
nand U8871 (N_8871,N_8330,N_8358);
nor U8872 (N_8872,N_8481,N_8437);
or U8873 (N_8873,N_8023,N_8198);
or U8874 (N_8874,N_8343,N_8171);
or U8875 (N_8875,N_8088,N_8315);
or U8876 (N_8876,N_8428,N_8117);
or U8877 (N_8877,N_8320,N_8190);
and U8878 (N_8878,N_8029,N_8148);
nor U8879 (N_8879,N_8273,N_8004);
and U8880 (N_8880,N_8117,N_8424);
and U8881 (N_8881,N_8416,N_8409);
and U8882 (N_8882,N_8289,N_8428);
and U8883 (N_8883,N_8079,N_8018);
or U8884 (N_8884,N_8409,N_8327);
nor U8885 (N_8885,N_8170,N_8443);
nand U8886 (N_8886,N_8262,N_8360);
nand U8887 (N_8887,N_8033,N_8497);
and U8888 (N_8888,N_8210,N_8496);
and U8889 (N_8889,N_8238,N_8205);
or U8890 (N_8890,N_8219,N_8210);
nand U8891 (N_8891,N_8445,N_8224);
nor U8892 (N_8892,N_8414,N_8068);
nand U8893 (N_8893,N_8490,N_8478);
and U8894 (N_8894,N_8233,N_8221);
xor U8895 (N_8895,N_8002,N_8292);
and U8896 (N_8896,N_8263,N_8146);
nor U8897 (N_8897,N_8389,N_8124);
and U8898 (N_8898,N_8220,N_8010);
and U8899 (N_8899,N_8199,N_8021);
and U8900 (N_8900,N_8253,N_8123);
or U8901 (N_8901,N_8234,N_8330);
nor U8902 (N_8902,N_8333,N_8273);
and U8903 (N_8903,N_8225,N_8003);
or U8904 (N_8904,N_8421,N_8102);
and U8905 (N_8905,N_8287,N_8433);
nand U8906 (N_8906,N_8084,N_8421);
nand U8907 (N_8907,N_8024,N_8382);
nand U8908 (N_8908,N_8094,N_8439);
nor U8909 (N_8909,N_8421,N_8345);
or U8910 (N_8910,N_8038,N_8304);
or U8911 (N_8911,N_8127,N_8264);
nor U8912 (N_8912,N_8284,N_8131);
nor U8913 (N_8913,N_8146,N_8016);
nor U8914 (N_8914,N_8457,N_8416);
or U8915 (N_8915,N_8183,N_8256);
nor U8916 (N_8916,N_8143,N_8047);
nor U8917 (N_8917,N_8320,N_8249);
or U8918 (N_8918,N_8237,N_8461);
nand U8919 (N_8919,N_8407,N_8177);
or U8920 (N_8920,N_8063,N_8359);
nand U8921 (N_8921,N_8321,N_8461);
or U8922 (N_8922,N_8342,N_8156);
nand U8923 (N_8923,N_8366,N_8250);
nor U8924 (N_8924,N_8368,N_8147);
or U8925 (N_8925,N_8409,N_8092);
and U8926 (N_8926,N_8310,N_8183);
nand U8927 (N_8927,N_8319,N_8269);
nor U8928 (N_8928,N_8087,N_8216);
nand U8929 (N_8929,N_8489,N_8133);
and U8930 (N_8930,N_8065,N_8309);
nor U8931 (N_8931,N_8290,N_8101);
and U8932 (N_8932,N_8167,N_8213);
and U8933 (N_8933,N_8037,N_8189);
and U8934 (N_8934,N_8441,N_8260);
and U8935 (N_8935,N_8049,N_8225);
or U8936 (N_8936,N_8470,N_8419);
nand U8937 (N_8937,N_8188,N_8406);
nand U8938 (N_8938,N_8344,N_8478);
nor U8939 (N_8939,N_8183,N_8274);
nand U8940 (N_8940,N_8313,N_8275);
xnor U8941 (N_8941,N_8235,N_8272);
or U8942 (N_8942,N_8378,N_8250);
nor U8943 (N_8943,N_8097,N_8296);
nor U8944 (N_8944,N_8255,N_8402);
nor U8945 (N_8945,N_8330,N_8073);
nor U8946 (N_8946,N_8399,N_8471);
nor U8947 (N_8947,N_8096,N_8436);
nor U8948 (N_8948,N_8173,N_8032);
nand U8949 (N_8949,N_8310,N_8172);
and U8950 (N_8950,N_8240,N_8082);
nand U8951 (N_8951,N_8203,N_8317);
nor U8952 (N_8952,N_8234,N_8262);
or U8953 (N_8953,N_8425,N_8273);
and U8954 (N_8954,N_8159,N_8133);
nor U8955 (N_8955,N_8401,N_8166);
and U8956 (N_8956,N_8149,N_8222);
or U8957 (N_8957,N_8299,N_8126);
or U8958 (N_8958,N_8177,N_8414);
nand U8959 (N_8959,N_8344,N_8075);
or U8960 (N_8960,N_8010,N_8103);
nand U8961 (N_8961,N_8359,N_8142);
nand U8962 (N_8962,N_8166,N_8075);
or U8963 (N_8963,N_8004,N_8335);
or U8964 (N_8964,N_8128,N_8197);
nor U8965 (N_8965,N_8414,N_8304);
or U8966 (N_8966,N_8445,N_8125);
nor U8967 (N_8967,N_8318,N_8222);
and U8968 (N_8968,N_8299,N_8393);
and U8969 (N_8969,N_8249,N_8312);
nand U8970 (N_8970,N_8102,N_8481);
or U8971 (N_8971,N_8400,N_8408);
or U8972 (N_8972,N_8425,N_8488);
and U8973 (N_8973,N_8145,N_8161);
nand U8974 (N_8974,N_8400,N_8041);
and U8975 (N_8975,N_8451,N_8052);
and U8976 (N_8976,N_8099,N_8249);
and U8977 (N_8977,N_8436,N_8093);
and U8978 (N_8978,N_8223,N_8477);
or U8979 (N_8979,N_8132,N_8302);
and U8980 (N_8980,N_8368,N_8166);
and U8981 (N_8981,N_8160,N_8253);
and U8982 (N_8982,N_8429,N_8178);
nand U8983 (N_8983,N_8139,N_8014);
nor U8984 (N_8984,N_8197,N_8002);
nand U8985 (N_8985,N_8200,N_8106);
xnor U8986 (N_8986,N_8001,N_8420);
nor U8987 (N_8987,N_8384,N_8072);
nand U8988 (N_8988,N_8351,N_8365);
nor U8989 (N_8989,N_8130,N_8021);
and U8990 (N_8990,N_8062,N_8022);
nor U8991 (N_8991,N_8334,N_8277);
and U8992 (N_8992,N_8185,N_8150);
nor U8993 (N_8993,N_8268,N_8029);
and U8994 (N_8994,N_8299,N_8382);
nand U8995 (N_8995,N_8452,N_8438);
nor U8996 (N_8996,N_8359,N_8013);
xor U8997 (N_8997,N_8363,N_8194);
and U8998 (N_8998,N_8323,N_8404);
nand U8999 (N_8999,N_8171,N_8219);
and U9000 (N_9000,N_8574,N_8597);
nor U9001 (N_9001,N_8664,N_8984);
nand U9002 (N_9002,N_8857,N_8925);
nand U9003 (N_9003,N_8906,N_8989);
nor U9004 (N_9004,N_8886,N_8983);
nand U9005 (N_9005,N_8666,N_8769);
or U9006 (N_9006,N_8627,N_8840);
or U9007 (N_9007,N_8905,N_8871);
nor U9008 (N_9008,N_8647,N_8918);
or U9009 (N_9009,N_8896,N_8941);
or U9010 (N_9010,N_8870,N_8963);
nand U9011 (N_9011,N_8598,N_8862);
or U9012 (N_9012,N_8690,N_8700);
nand U9013 (N_9013,N_8673,N_8907);
and U9014 (N_9014,N_8833,N_8736);
and U9015 (N_9015,N_8851,N_8694);
nand U9016 (N_9016,N_8646,N_8744);
nand U9017 (N_9017,N_8997,N_8590);
and U9018 (N_9018,N_8727,N_8572);
or U9019 (N_9019,N_8623,N_8708);
nand U9020 (N_9020,N_8578,N_8576);
nor U9021 (N_9021,N_8709,N_8934);
and U9022 (N_9022,N_8575,N_8781);
or U9023 (N_9023,N_8856,N_8930);
or U9024 (N_9024,N_8763,N_8844);
nand U9025 (N_9025,N_8835,N_8900);
nor U9026 (N_9026,N_8799,N_8739);
nand U9027 (N_9027,N_8832,N_8669);
nand U9028 (N_9028,N_8620,N_8848);
nand U9029 (N_9029,N_8991,N_8765);
or U9030 (N_9030,N_8797,N_8698);
nand U9031 (N_9031,N_8805,N_8704);
nor U9032 (N_9032,N_8823,N_8924);
and U9033 (N_9033,N_8845,N_8957);
nor U9034 (N_9034,N_8868,N_8699);
and U9035 (N_9035,N_8536,N_8839);
or U9036 (N_9036,N_8894,N_8585);
or U9037 (N_9037,N_8693,N_8611);
nor U9038 (N_9038,N_8766,N_8811);
and U9039 (N_9039,N_8786,N_8922);
nor U9040 (N_9040,N_8733,N_8770);
or U9041 (N_9041,N_8682,N_8943);
nand U9042 (N_9042,N_8773,N_8715);
or U9043 (N_9043,N_8538,N_8652);
nand U9044 (N_9044,N_8893,N_8517);
and U9045 (N_9045,N_8692,N_8942);
nor U9046 (N_9046,N_8768,N_8561);
or U9047 (N_9047,N_8954,N_8961);
and U9048 (N_9048,N_8509,N_8742);
nand U9049 (N_9049,N_8541,N_8842);
or U9050 (N_9050,N_8753,N_8684);
or U9051 (N_9051,N_8676,N_8818);
or U9052 (N_9052,N_8814,N_8858);
or U9053 (N_9053,N_8508,N_8558);
nor U9054 (N_9054,N_8677,N_8982);
or U9055 (N_9055,N_8792,N_8826);
and U9056 (N_9056,N_8582,N_8813);
and U9057 (N_9057,N_8969,N_8542);
nor U9058 (N_9058,N_8663,N_8780);
nor U9059 (N_9059,N_8820,N_8668);
nand U9060 (N_9060,N_8904,N_8951);
nand U9061 (N_9061,N_8606,N_8685);
nor U9062 (N_9062,N_8750,N_8625);
nor U9063 (N_9063,N_8808,N_8793);
nand U9064 (N_9064,N_8747,N_8824);
nand U9065 (N_9065,N_8819,N_8919);
and U9066 (N_9066,N_8847,N_8568);
nor U9067 (N_9067,N_8931,N_8630);
or U9068 (N_9068,N_8827,N_8605);
and U9069 (N_9069,N_8529,N_8595);
nand U9070 (N_9070,N_8571,N_8939);
and U9071 (N_9071,N_8998,N_8926);
nor U9072 (N_9072,N_8622,N_8658);
xnor U9073 (N_9073,N_8688,N_8557);
nor U9074 (N_9074,N_8881,N_8591);
or U9075 (N_9075,N_8874,N_8988);
or U9076 (N_9076,N_8701,N_8927);
nor U9077 (N_9077,N_8873,N_8539);
and U9078 (N_9078,N_8807,N_8959);
nor U9079 (N_9079,N_8566,N_8854);
nor U9080 (N_9080,N_8817,N_8644);
and U9081 (N_9081,N_8718,N_8626);
nor U9082 (N_9082,N_8635,N_8777);
or U9083 (N_9083,N_8801,N_8995);
or U9084 (N_9084,N_8902,N_8501);
nand U9085 (N_9085,N_8901,N_8810);
and U9086 (N_9086,N_8895,N_8994);
nand U9087 (N_9087,N_8899,N_8752);
or U9088 (N_9088,N_8686,N_8681);
and U9089 (N_9089,N_8678,N_8527);
nand U9090 (N_9090,N_8710,N_8608);
or U9091 (N_9091,N_8697,N_8592);
nand U9092 (N_9092,N_8916,N_8565);
nand U9093 (N_9093,N_8756,N_8973);
nand U9094 (N_9094,N_8522,N_8649);
or U9095 (N_9095,N_8860,N_8948);
and U9096 (N_9096,N_8639,N_8754);
and U9097 (N_9097,N_8962,N_8967);
or U9098 (N_9098,N_8788,N_8655);
nand U9099 (N_9099,N_8938,N_8530);
and U9100 (N_9100,N_8737,N_8841);
nor U9101 (N_9101,N_8974,N_8723);
nand U9102 (N_9102,N_8555,N_8535);
and U9103 (N_9103,N_8950,N_8534);
or U9104 (N_9104,N_8540,N_8993);
nand U9105 (N_9105,N_8774,N_8637);
nand U9106 (N_9106,N_8556,N_8712);
nor U9107 (N_9107,N_8936,N_8695);
or U9108 (N_9108,N_8751,N_8716);
nand U9109 (N_9109,N_8528,N_8828);
nand U9110 (N_9110,N_8720,N_8843);
or U9111 (N_9111,N_8779,N_8581);
or U9112 (N_9112,N_8859,N_8587);
or U9113 (N_9113,N_8577,N_8722);
or U9114 (N_9114,N_8641,N_8691);
or U9115 (N_9115,N_8849,N_8866);
and U9116 (N_9116,N_8913,N_8505);
nor U9117 (N_9117,N_8875,N_8564);
and U9118 (N_9118,N_8607,N_8724);
or U9119 (N_9119,N_8514,N_8759);
or U9120 (N_9120,N_8992,N_8762);
xor U9121 (N_9121,N_8729,N_8648);
and U9122 (N_9122,N_8795,N_8711);
or U9123 (N_9123,N_8889,N_8702);
nand U9124 (N_9124,N_8616,N_8563);
nand U9125 (N_9125,N_8589,N_8846);
nor U9126 (N_9126,N_8782,N_8730);
and U9127 (N_9127,N_8731,N_8549);
nand U9128 (N_9128,N_8660,N_8883);
or U9129 (N_9129,N_8800,N_8594);
and U9130 (N_9130,N_8834,N_8877);
nor U9131 (N_9131,N_8944,N_8500);
and U9132 (N_9132,N_8569,N_8515);
nand U9133 (N_9133,N_8532,N_8659);
or U9134 (N_9134,N_8772,N_8728);
nor U9135 (N_9135,N_8815,N_8816);
or U9136 (N_9136,N_8506,N_8657);
and U9137 (N_9137,N_8741,N_8533);
nor U9138 (N_9138,N_8651,N_8670);
xnor U9139 (N_9139,N_8619,N_8830);
and U9140 (N_9140,N_8865,N_8725);
or U9141 (N_9141,N_8952,N_8642);
and U9142 (N_9142,N_8547,N_8882);
nor U9143 (N_9143,N_8897,N_8852);
nor U9144 (N_9144,N_8749,N_8999);
nand U9145 (N_9145,N_8584,N_8764);
xor U9146 (N_9146,N_8884,N_8617);
and U9147 (N_9147,N_8634,N_8512);
nand U9148 (N_9148,N_8831,N_8559);
nor U9149 (N_9149,N_8794,N_8554);
or U9150 (N_9150,N_8504,N_8912);
and U9151 (N_9151,N_8789,N_8638);
nand U9152 (N_9152,N_8775,N_8806);
nand U9153 (N_9153,N_8654,N_8879);
or U9154 (N_9154,N_8560,N_8628);
or U9155 (N_9155,N_8864,N_8636);
nand U9156 (N_9156,N_8971,N_8932);
nor U9157 (N_9157,N_8996,N_8910);
or U9158 (N_9158,N_8940,N_8738);
or U9159 (N_9159,N_8872,N_8719);
nor U9160 (N_9160,N_8714,N_8914);
or U9161 (N_9161,N_8802,N_8543);
nand U9162 (N_9162,N_8545,N_8550);
and U9163 (N_9163,N_8632,N_8867);
nor U9164 (N_9164,N_8903,N_8825);
and U9165 (N_9165,N_8758,N_8562);
or U9166 (N_9166,N_8675,N_8975);
and U9167 (N_9167,N_8643,N_8829);
nor U9168 (N_9168,N_8890,N_8933);
nand U9169 (N_9169,N_8920,N_8911);
nand U9170 (N_9170,N_8885,N_8985);
or U9171 (N_9171,N_8946,N_8850);
and U9172 (N_9172,N_8672,N_8990);
nand U9173 (N_9173,N_8687,N_8612);
nand U9174 (N_9174,N_8705,N_8599);
or U9175 (N_9175,N_8537,N_8583);
nand U9176 (N_9176,N_8898,N_8548);
or U9177 (N_9177,N_8812,N_8965);
nor U9178 (N_9178,N_8978,N_8588);
and U9179 (N_9179,N_8908,N_8615);
nand U9180 (N_9180,N_8656,N_8503);
or U9181 (N_9181,N_8821,N_8665);
or U9182 (N_9182,N_8964,N_8757);
and U9183 (N_9183,N_8679,N_8523);
and U9184 (N_9184,N_8980,N_8502);
nor U9185 (N_9185,N_8979,N_8836);
xor U9186 (N_9186,N_8928,N_8546);
or U9187 (N_9187,N_8573,N_8531);
or U9188 (N_9188,N_8863,N_8683);
nand U9189 (N_9189,N_8618,N_8707);
and U9190 (N_9190,N_8853,N_8972);
or U9191 (N_9191,N_8519,N_8776);
or U9192 (N_9192,N_8633,N_8521);
or U9193 (N_9193,N_8680,N_8721);
nand U9194 (N_9194,N_8949,N_8955);
nand U9195 (N_9195,N_8524,N_8953);
or U9196 (N_9196,N_8511,N_8778);
nor U9197 (N_9197,N_8760,N_8703);
and U9198 (N_9198,N_8876,N_8966);
nor U9199 (N_9199,N_8551,N_8662);
and U9200 (N_9200,N_8614,N_8986);
nor U9201 (N_9201,N_8935,N_8790);
and U9202 (N_9202,N_8929,N_8609);
nand U9203 (N_9203,N_8604,N_8861);
and U9204 (N_9204,N_8706,N_8610);
or U9205 (N_9205,N_8987,N_8915);
or U9206 (N_9206,N_8645,N_8570);
nor U9207 (N_9207,N_8887,N_8796);
nor U9208 (N_9208,N_8970,N_8717);
and U9209 (N_9209,N_8785,N_8732);
or U9210 (N_9210,N_8809,N_8923);
or U9211 (N_9211,N_8981,N_8888);
nand U9212 (N_9212,N_8674,N_8621);
nor U9213 (N_9213,N_8783,N_8507);
nor U9214 (N_9214,N_8787,N_8804);
nor U9215 (N_9215,N_8603,N_8968);
nor U9216 (N_9216,N_8746,N_8956);
nand U9217 (N_9217,N_8629,N_8784);
nor U9218 (N_9218,N_8891,N_8650);
nand U9219 (N_9219,N_8520,N_8653);
nand U9220 (N_9220,N_8667,N_8977);
or U9221 (N_9221,N_8516,N_8713);
and U9222 (N_9222,N_8921,N_8593);
nand U9223 (N_9223,N_8518,N_8892);
nor U9224 (N_9224,N_8748,N_8771);
nor U9225 (N_9225,N_8880,N_8947);
nor U9226 (N_9226,N_8878,N_8798);
and U9227 (N_9227,N_8586,N_8937);
nor U9228 (N_9228,N_8726,N_8945);
nand U9229 (N_9229,N_8803,N_8745);
or U9230 (N_9230,N_8917,N_8838);
nand U9231 (N_9231,N_8761,N_8567);
nand U9232 (N_9232,N_8526,N_8855);
or U9233 (N_9233,N_8791,N_8544);
or U9234 (N_9234,N_8661,N_8631);
nor U9235 (N_9235,N_8960,N_8579);
or U9236 (N_9236,N_8767,N_8740);
nor U9237 (N_9237,N_8869,N_8958);
and U9238 (N_9238,N_8510,N_8743);
nand U9239 (N_9239,N_8596,N_8837);
nor U9240 (N_9240,N_8601,N_8689);
nand U9241 (N_9241,N_8735,N_8553);
or U9242 (N_9242,N_8513,N_8671);
and U9243 (N_9243,N_8755,N_8909);
nand U9244 (N_9244,N_8602,N_8613);
nand U9245 (N_9245,N_8696,N_8525);
nand U9246 (N_9246,N_8624,N_8976);
and U9247 (N_9247,N_8580,N_8734);
and U9248 (N_9248,N_8822,N_8552);
nor U9249 (N_9249,N_8640,N_8600);
and U9250 (N_9250,N_8820,N_8571);
and U9251 (N_9251,N_8917,N_8808);
or U9252 (N_9252,N_8625,N_8660);
nand U9253 (N_9253,N_8853,N_8814);
xnor U9254 (N_9254,N_8765,N_8944);
nor U9255 (N_9255,N_8660,N_8630);
or U9256 (N_9256,N_8907,N_8953);
nand U9257 (N_9257,N_8640,N_8692);
and U9258 (N_9258,N_8930,N_8989);
or U9259 (N_9259,N_8827,N_8686);
nor U9260 (N_9260,N_8722,N_8946);
nor U9261 (N_9261,N_8778,N_8919);
nand U9262 (N_9262,N_8889,N_8870);
nor U9263 (N_9263,N_8531,N_8631);
nand U9264 (N_9264,N_8804,N_8536);
nor U9265 (N_9265,N_8542,N_8775);
or U9266 (N_9266,N_8690,N_8726);
and U9267 (N_9267,N_8694,N_8531);
or U9268 (N_9268,N_8636,N_8971);
and U9269 (N_9269,N_8806,N_8677);
or U9270 (N_9270,N_8613,N_8871);
or U9271 (N_9271,N_8855,N_8854);
or U9272 (N_9272,N_8624,N_8738);
nand U9273 (N_9273,N_8724,N_8501);
nor U9274 (N_9274,N_8743,N_8948);
nand U9275 (N_9275,N_8759,N_8916);
nor U9276 (N_9276,N_8764,N_8861);
and U9277 (N_9277,N_8510,N_8651);
or U9278 (N_9278,N_8538,N_8846);
or U9279 (N_9279,N_8944,N_8519);
and U9280 (N_9280,N_8747,N_8846);
nand U9281 (N_9281,N_8907,N_8697);
and U9282 (N_9282,N_8688,N_8728);
nor U9283 (N_9283,N_8631,N_8535);
and U9284 (N_9284,N_8502,N_8750);
nor U9285 (N_9285,N_8844,N_8568);
and U9286 (N_9286,N_8583,N_8681);
nor U9287 (N_9287,N_8611,N_8811);
nand U9288 (N_9288,N_8529,N_8778);
nand U9289 (N_9289,N_8850,N_8969);
nor U9290 (N_9290,N_8714,N_8967);
or U9291 (N_9291,N_8860,N_8710);
nand U9292 (N_9292,N_8596,N_8600);
and U9293 (N_9293,N_8742,N_8837);
nor U9294 (N_9294,N_8844,N_8745);
and U9295 (N_9295,N_8864,N_8750);
or U9296 (N_9296,N_8640,N_8611);
or U9297 (N_9297,N_8658,N_8889);
nand U9298 (N_9298,N_8805,N_8955);
nor U9299 (N_9299,N_8659,N_8628);
and U9300 (N_9300,N_8588,N_8673);
and U9301 (N_9301,N_8624,N_8996);
or U9302 (N_9302,N_8545,N_8836);
nor U9303 (N_9303,N_8750,N_8598);
or U9304 (N_9304,N_8785,N_8546);
nor U9305 (N_9305,N_8986,N_8585);
nor U9306 (N_9306,N_8635,N_8651);
nor U9307 (N_9307,N_8917,N_8895);
nand U9308 (N_9308,N_8899,N_8556);
and U9309 (N_9309,N_8906,N_8516);
nor U9310 (N_9310,N_8861,N_8510);
and U9311 (N_9311,N_8841,N_8795);
nand U9312 (N_9312,N_8847,N_8684);
or U9313 (N_9313,N_8603,N_8637);
nor U9314 (N_9314,N_8558,N_8789);
and U9315 (N_9315,N_8890,N_8796);
nor U9316 (N_9316,N_8996,N_8930);
nor U9317 (N_9317,N_8738,N_8615);
xor U9318 (N_9318,N_8722,N_8705);
or U9319 (N_9319,N_8946,N_8952);
xor U9320 (N_9320,N_8738,N_8853);
and U9321 (N_9321,N_8751,N_8584);
nor U9322 (N_9322,N_8590,N_8616);
and U9323 (N_9323,N_8931,N_8918);
and U9324 (N_9324,N_8626,N_8862);
nor U9325 (N_9325,N_8884,N_8540);
xnor U9326 (N_9326,N_8821,N_8913);
nand U9327 (N_9327,N_8871,N_8879);
nand U9328 (N_9328,N_8725,N_8920);
nor U9329 (N_9329,N_8658,N_8775);
and U9330 (N_9330,N_8692,N_8603);
nor U9331 (N_9331,N_8828,N_8767);
and U9332 (N_9332,N_8978,N_8575);
or U9333 (N_9333,N_8960,N_8946);
or U9334 (N_9334,N_8602,N_8820);
and U9335 (N_9335,N_8578,N_8855);
nor U9336 (N_9336,N_8735,N_8783);
or U9337 (N_9337,N_8777,N_8541);
nor U9338 (N_9338,N_8802,N_8956);
nor U9339 (N_9339,N_8707,N_8508);
and U9340 (N_9340,N_8792,N_8841);
and U9341 (N_9341,N_8519,N_8752);
nand U9342 (N_9342,N_8611,N_8961);
or U9343 (N_9343,N_8593,N_8565);
and U9344 (N_9344,N_8565,N_8513);
nor U9345 (N_9345,N_8890,N_8685);
and U9346 (N_9346,N_8944,N_8810);
or U9347 (N_9347,N_8659,N_8866);
or U9348 (N_9348,N_8600,N_8850);
or U9349 (N_9349,N_8911,N_8696);
or U9350 (N_9350,N_8756,N_8948);
nand U9351 (N_9351,N_8767,N_8571);
or U9352 (N_9352,N_8772,N_8717);
and U9353 (N_9353,N_8751,N_8511);
and U9354 (N_9354,N_8698,N_8807);
or U9355 (N_9355,N_8953,N_8606);
nor U9356 (N_9356,N_8596,N_8788);
nand U9357 (N_9357,N_8600,N_8934);
nor U9358 (N_9358,N_8705,N_8615);
or U9359 (N_9359,N_8557,N_8949);
and U9360 (N_9360,N_8750,N_8874);
nand U9361 (N_9361,N_8802,N_8814);
nand U9362 (N_9362,N_8604,N_8907);
or U9363 (N_9363,N_8878,N_8583);
nor U9364 (N_9364,N_8864,N_8886);
or U9365 (N_9365,N_8879,N_8906);
and U9366 (N_9366,N_8882,N_8532);
or U9367 (N_9367,N_8567,N_8894);
nor U9368 (N_9368,N_8853,N_8848);
and U9369 (N_9369,N_8770,N_8977);
and U9370 (N_9370,N_8501,N_8819);
nand U9371 (N_9371,N_8805,N_8769);
or U9372 (N_9372,N_8616,N_8660);
or U9373 (N_9373,N_8782,N_8993);
nor U9374 (N_9374,N_8985,N_8832);
nor U9375 (N_9375,N_8509,N_8925);
and U9376 (N_9376,N_8832,N_8785);
nand U9377 (N_9377,N_8925,N_8592);
nor U9378 (N_9378,N_8732,N_8904);
and U9379 (N_9379,N_8695,N_8703);
nand U9380 (N_9380,N_8655,N_8720);
xor U9381 (N_9381,N_8650,N_8876);
or U9382 (N_9382,N_8686,N_8852);
and U9383 (N_9383,N_8732,N_8596);
nand U9384 (N_9384,N_8899,N_8603);
or U9385 (N_9385,N_8553,N_8803);
and U9386 (N_9386,N_8977,N_8695);
and U9387 (N_9387,N_8944,N_8853);
and U9388 (N_9388,N_8768,N_8741);
nand U9389 (N_9389,N_8620,N_8840);
and U9390 (N_9390,N_8736,N_8993);
and U9391 (N_9391,N_8855,N_8580);
or U9392 (N_9392,N_8649,N_8521);
and U9393 (N_9393,N_8670,N_8839);
nor U9394 (N_9394,N_8654,N_8858);
xnor U9395 (N_9395,N_8607,N_8625);
or U9396 (N_9396,N_8525,N_8917);
nor U9397 (N_9397,N_8981,N_8537);
nor U9398 (N_9398,N_8727,N_8620);
or U9399 (N_9399,N_8508,N_8939);
and U9400 (N_9400,N_8957,N_8925);
or U9401 (N_9401,N_8824,N_8983);
and U9402 (N_9402,N_8879,N_8658);
or U9403 (N_9403,N_8922,N_8566);
nand U9404 (N_9404,N_8824,N_8965);
or U9405 (N_9405,N_8522,N_8571);
nand U9406 (N_9406,N_8788,N_8837);
or U9407 (N_9407,N_8717,N_8529);
and U9408 (N_9408,N_8724,N_8892);
or U9409 (N_9409,N_8715,N_8910);
or U9410 (N_9410,N_8528,N_8692);
and U9411 (N_9411,N_8726,N_8581);
or U9412 (N_9412,N_8712,N_8812);
and U9413 (N_9413,N_8857,N_8798);
or U9414 (N_9414,N_8745,N_8522);
nor U9415 (N_9415,N_8989,N_8508);
and U9416 (N_9416,N_8662,N_8573);
nor U9417 (N_9417,N_8694,N_8948);
or U9418 (N_9418,N_8558,N_8545);
xnor U9419 (N_9419,N_8589,N_8867);
nor U9420 (N_9420,N_8829,N_8909);
and U9421 (N_9421,N_8544,N_8671);
nor U9422 (N_9422,N_8596,N_8628);
or U9423 (N_9423,N_8703,N_8652);
or U9424 (N_9424,N_8964,N_8674);
nand U9425 (N_9425,N_8771,N_8579);
or U9426 (N_9426,N_8604,N_8630);
and U9427 (N_9427,N_8551,N_8583);
and U9428 (N_9428,N_8936,N_8690);
or U9429 (N_9429,N_8507,N_8723);
or U9430 (N_9430,N_8546,N_8957);
nor U9431 (N_9431,N_8769,N_8633);
or U9432 (N_9432,N_8514,N_8933);
and U9433 (N_9433,N_8671,N_8972);
or U9434 (N_9434,N_8899,N_8632);
nor U9435 (N_9435,N_8696,N_8531);
nand U9436 (N_9436,N_8807,N_8568);
nand U9437 (N_9437,N_8593,N_8687);
or U9438 (N_9438,N_8521,N_8646);
nor U9439 (N_9439,N_8666,N_8655);
nand U9440 (N_9440,N_8505,N_8600);
and U9441 (N_9441,N_8608,N_8659);
or U9442 (N_9442,N_8771,N_8655);
nand U9443 (N_9443,N_8751,N_8904);
nor U9444 (N_9444,N_8760,N_8666);
nor U9445 (N_9445,N_8609,N_8796);
and U9446 (N_9446,N_8853,N_8692);
nand U9447 (N_9447,N_8752,N_8741);
nand U9448 (N_9448,N_8767,N_8613);
and U9449 (N_9449,N_8550,N_8659);
nor U9450 (N_9450,N_8613,N_8589);
nor U9451 (N_9451,N_8561,N_8866);
or U9452 (N_9452,N_8533,N_8695);
nor U9453 (N_9453,N_8851,N_8864);
or U9454 (N_9454,N_8948,N_8649);
nand U9455 (N_9455,N_8978,N_8618);
and U9456 (N_9456,N_8813,N_8666);
nor U9457 (N_9457,N_8725,N_8762);
or U9458 (N_9458,N_8687,N_8716);
and U9459 (N_9459,N_8776,N_8836);
nor U9460 (N_9460,N_8766,N_8872);
or U9461 (N_9461,N_8934,N_8758);
and U9462 (N_9462,N_8828,N_8707);
or U9463 (N_9463,N_8902,N_8893);
or U9464 (N_9464,N_8848,N_8874);
nand U9465 (N_9465,N_8843,N_8779);
and U9466 (N_9466,N_8875,N_8678);
nor U9467 (N_9467,N_8680,N_8528);
xor U9468 (N_9468,N_8552,N_8698);
nor U9469 (N_9469,N_8906,N_8994);
or U9470 (N_9470,N_8903,N_8953);
nor U9471 (N_9471,N_8930,N_8525);
nor U9472 (N_9472,N_8862,N_8967);
nor U9473 (N_9473,N_8888,N_8582);
nor U9474 (N_9474,N_8992,N_8793);
nor U9475 (N_9475,N_8647,N_8841);
or U9476 (N_9476,N_8792,N_8767);
and U9477 (N_9477,N_8728,N_8504);
nand U9478 (N_9478,N_8690,N_8637);
nor U9479 (N_9479,N_8805,N_8524);
and U9480 (N_9480,N_8703,N_8532);
nand U9481 (N_9481,N_8575,N_8774);
and U9482 (N_9482,N_8826,N_8699);
nor U9483 (N_9483,N_8618,N_8654);
and U9484 (N_9484,N_8590,N_8842);
or U9485 (N_9485,N_8900,N_8883);
xor U9486 (N_9486,N_8685,N_8689);
or U9487 (N_9487,N_8890,N_8543);
xnor U9488 (N_9488,N_8802,N_8857);
and U9489 (N_9489,N_8799,N_8700);
nor U9490 (N_9490,N_8785,N_8953);
nand U9491 (N_9491,N_8664,N_8862);
xor U9492 (N_9492,N_8584,N_8837);
or U9493 (N_9493,N_8746,N_8886);
nand U9494 (N_9494,N_8802,N_8702);
nand U9495 (N_9495,N_8763,N_8696);
xor U9496 (N_9496,N_8599,N_8692);
and U9497 (N_9497,N_8635,N_8646);
or U9498 (N_9498,N_8728,N_8963);
nand U9499 (N_9499,N_8783,N_8516);
or U9500 (N_9500,N_9403,N_9245);
nand U9501 (N_9501,N_9410,N_9421);
nor U9502 (N_9502,N_9334,N_9052);
nor U9503 (N_9503,N_9036,N_9125);
or U9504 (N_9504,N_9474,N_9121);
nor U9505 (N_9505,N_9089,N_9078);
or U9506 (N_9506,N_9023,N_9493);
nand U9507 (N_9507,N_9472,N_9006);
nor U9508 (N_9508,N_9058,N_9098);
or U9509 (N_9509,N_9473,N_9366);
and U9510 (N_9510,N_9271,N_9244);
or U9511 (N_9511,N_9181,N_9275);
or U9512 (N_9512,N_9306,N_9350);
or U9513 (N_9513,N_9320,N_9030);
and U9514 (N_9514,N_9080,N_9408);
xor U9515 (N_9515,N_9468,N_9242);
nor U9516 (N_9516,N_9295,N_9438);
nor U9517 (N_9517,N_9362,N_9377);
and U9518 (N_9518,N_9441,N_9364);
nor U9519 (N_9519,N_9489,N_9158);
nor U9520 (N_9520,N_9418,N_9307);
or U9521 (N_9521,N_9073,N_9356);
and U9522 (N_9522,N_9162,N_9127);
or U9523 (N_9523,N_9312,N_9458);
and U9524 (N_9524,N_9116,N_9259);
nand U9525 (N_9525,N_9147,N_9071);
nor U9526 (N_9526,N_9380,N_9016);
or U9527 (N_9527,N_9387,N_9015);
nor U9528 (N_9528,N_9084,N_9165);
and U9529 (N_9529,N_9417,N_9440);
or U9530 (N_9530,N_9237,N_9247);
nand U9531 (N_9531,N_9288,N_9390);
or U9532 (N_9532,N_9461,N_9140);
nand U9533 (N_9533,N_9037,N_9484);
or U9534 (N_9534,N_9207,N_9045);
or U9535 (N_9535,N_9251,N_9059);
nand U9536 (N_9536,N_9286,N_9117);
nand U9537 (N_9537,N_9270,N_9424);
or U9538 (N_9538,N_9012,N_9289);
nand U9539 (N_9539,N_9194,N_9075);
nand U9540 (N_9540,N_9197,N_9381);
and U9541 (N_9541,N_9300,N_9457);
or U9542 (N_9542,N_9278,N_9296);
or U9543 (N_9543,N_9298,N_9466);
nor U9544 (N_9544,N_9425,N_9105);
xnor U9545 (N_9545,N_9496,N_9238);
and U9546 (N_9546,N_9254,N_9463);
nor U9547 (N_9547,N_9445,N_9324);
or U9548 (N_9548,N_9217,N_9308);
nor U9549 (N_9549,N_9026,N_9335);
nand U9550 (N_9550,N_9476,N_9309);
nand U9551 (N_9551,N_9189,N_9253);
nand U9552 (N_9552,N_9109,N_9118);
nor U9553 (N_9553,N_9021,N_9280);
nand U9554 (N_9554,N_9164,N_9115);
nand U9555 (N_9555,N_9317,N_9363);
and U9556 (N_9556,N_9166,N_9339);
nor U9557 (N_9557,N_9120,N_9459);
and U9558 (N_9558,N_9234,N_9383);
or U9559 (N_9559,N_9348,N_9246);
nor U9560 (N_9560,N_9170,N_9240);
and U9561 (N_9561,N_9415,N_9337);
or U9562 (N_9562,N_9107,N_9430);
nor U9563 (N_9563,N_9231,N_9175);
and U9564 (N_9564,N_9358,N_9029);
and U9565 (N_9565,N_9393,N_9169);
nand U9566 (N_9566,N_9025,N_9227);
and U9567 (N_9567,N_9326,N_9018);
nor U9568 (N_9568,N_9149,N_9192);
or U9569 (N_9569,N_9310,N_9123);
nand U9570 (N_9570,N_9336,N_9276);
or U9571 (N_9571,N_9420,N_9272);
or U9572 (N_9572,N_9055,N_9104);
or U9573 (N_9573,N_9034,N_9316);
nor U9574 (N_9574,N_9004,N_9369);
or U9575 (N_9575,N_9382,N_9093);
nor U9576 (N_9576,N_9135,N_9223);
and U9577 (N_9577,N_9313,N_9401);
and U9578 (N_9578,N_9002,N_9428);
and U9579 (N_9579,N_9396,N_9322);
nor U9580 (N_9580,N_9152,N_9460);
or U9581 (N_9581,N_9102,N_9051);
or U9582 (N_9582,N_9357,N_9371);
nand U9583 (N_9583,N_9154,N_9434);
nor U9584 (N_9584,N_9222,N_9119);
and U9585 (N_9585,N_9454,N_9359);
nor U9586 (N_9586,N_9096,N_9367);
nor U9587 (N_9587,N_9114,N_9083);
or U9588 (N_9588,N_9103,N_9331);
or U9589 (N_9589,N_9482,N_9395);
nand U9590 (N_9590,N_9450,N_9293);
nor U9591 (N_9591,N_9236,N_9009);
nand U9592 (N_9592,N_9360,N_9038);
nand U9593 (N_9593,N_9294,N_9354);
nand U9594 (N_9594,N_9427,N_9255);
nand U9595 (N_9595,N_9304,N_9409);
and U9596 (N_9596,N_9206,N_9419);
nand U9597 (N_9597,N_9024,N_9475);
and U9598 (N_9598,N_9407,N_9325);
and U9599 (N_9599,N_9195,N_9469);
nor U9600 (N_9600,N_9008,N_9447);
nor U9601 (N_9601,N_9077,N_9049);
and U9602 (N_9602,N_9060,N_9101);
and U9603 (N_9603,N_9465,N_9173);
xnor U9604 (N_9604,N_9057,N_9453);
and U9605 (N_9605,N_9411,N_9133);
and U9606 (N_9606,N_9068,N_9228);
or U9607 (N_9607,N_9072,N_9185);
nand U9608 (N_9608,N_9379,N_9178);
or U9609 (N_9609,N_9292,N_9394);
nand U9610 (N_9610,N_9263,N_9001);
nand U9611 (N_9611,N_9190,N_9168);
or U9612 (N_9612,N_9398,N_9079);
nand U9613 (N_9613,N_9070,N_9128);
or U9614 (N_9614,N_9129,N_9368);
and U9615 (N_9615,N_9056,N_9488);
and U9616 (N_9616,N_9462,N_9157);
nand U9617 (N_9617,N_9215,N_9451);
nor U9618 (N_9618,N_9290,N_9402);
nor U9619 (N_9619,N_9014,N_9141);
or U9620 (N_9620,N_9282,N_9346);
and U9621 (N_9621,N_9048,N_9176);
or U9622 (N_9622,N_9497,N_9091);
nand U9623 (N_9623,N_9188,N_9266);
and U9624 (N_9624,N_9315,N_9318);
nand U9625 (N_9625,N_9097,N_9005);
nor U9626 (N_9626,N_9201,N_9405);
or U9627 (N_9627,N_9180,N_9392);
and U9628 (N_9628,N_9010,N_9376);
nor U9629 (N_9629,N_9239,N_9481);
xor U9630 (N_9630,N_9404,N_9327);
nand U9631 (N_9631,N_9142,N_9137);
nand U9632 (N_9632,N_9042,N_9375);
xnor U9633 (N_9633,N_9291,N_9136);
or U9634 (N_9634,N_9384,N_9446);
xnor U9635 (N_9635,N_9495,N_9491);
nor U9636 (N_9636,N_9439,N_9100);
and U9637 (N_9637,N_9130,N_9437);
nor U9638 (N_9638,N_9480,N_9455);
nand U9639 (N_9639,N_9186,N_9041);
or U9640 (N_9640,N_9456,N_9338);
or U9641 (N_9641,N_9494,N_9256);
and U9642 (N_9642,N_9349,N_9321);
nor U9643 (N_9643,N_9370,N_9126);
or U9644 (N_9644,N_9200,N_9039);
or U9645 (N_9645,N_9490,N_9423);
or U9646 (N_9646,N_9183,N_9066);
nand U9647 (N_9647,N_9297,N_9351);
nor U9648 (N_9648,N_9063,N_9262);
and U9649 (N_9649,N_9341,N_9171);
nand U9650 (N_9650,N_9074,N_9241);
nor U9651 (N_9651,N_9378,N_9330);
nand U9652 (N_9652,N_9145,N_9267);
and U9653 (N_9653,N_9210,N_9081);
nor U9654 (N_9654,N_9365,N_9213);
nor U9655 (N_9655,N_9232,N_9198);
or U9656 (N_9656,N_9429,N_9265);
or U9657 (N_9657,N_9167,N_9218);
or U9658 (N_9658,N_9281,N_9448);
and U9659 (N_9659,N_9478,N_9035);
or U9660 (N_9660,N_9172,N_9487);
and U9661 (N_9661,N_9179,N_9248);
and U9662 (N_9662,N_9143,N_9435);
nor U9663 (N_9663,N_9249,N_9040);
and U9664 (N_9664,N_9054,N_9260);
or U9665 (N_9665,N_9470,N_9323);
nor U9666 (N_9666,N_9412,N_9082);
or U9667 (N_9667,N_9193,N_9314);
and U9668 (N_9668,N_9062,N_9486);
and U9669 (N_9669,N_9416,N_9191);
nand U9670 (N_9670,N_9122,N_9144);
nand U9671 (N_9671,N_9088,N_9065);
nor U9672 (N_9672,N_9444,N_9400);
or U9673 (N_9673,N_9046,N_9344);
nand U9674 (N_9674,N_9146,N_9386);
nand U9675 (N_9675,N_9053,N_9220);
or U9676 (N_9676,N_9452,N_9011);
and U9677 (N_9677,N_9095,N_9233);
nand U9678 (N_9678,N_9433,N_9064);
nand U9679 (N_9679,N_9148,N_9050);
nor U9680 (N_9680,N_9027,N_9299);
nor U9681 (N_9681,N_9258,N_9092);
and U9682 (N_9682,N_9043,N_9264);
nand U9683 (N_9683,N_9216,N_9187);
or U9684 (N_9684,N_9174,N_9464);
or U9685 (N_9685,N_9340,N_9305);
nand U9686 (N_9686,N_9028,N_9328);
nand U9687 (N_9687,N_9044,N_9467);
nand U9688 (N_9688,N_9243,N_9199);
and U9689 (N_9689,N_9252,N_9414);
nor U9690 (N_9690,N_9150,N_9355);
nor U9691 (N_9691,N_9000,N_9373);
nand U9692 (N_9692,N_9449,N_9224);
nor U9693 (N_9693,N_9229,N_9431);
nor U9694 (N_9694,N_9153,N_9139);
or U9695 (N_9695,N_9221,N_9177);
and U9696 (N_9696,N_9069,N_9160);
or U9697 (N_9697,N_9283,N_9226);
nand U9698 (N_9698,N_9319,N_9332);
nand U9699 (N_9699,N_9397,N_9134);
and U9700 (N_9700,N_9204,N_9131);
nand U9701 (N_9701,N_9047,N_9273);
nor U9702 (N_9702,N_9436,N_9302);
or U9703 (N_9703,N_9061,N_9342);
or U9704 (N_9704,N_9261,N_9374);
nor U9705 (N_9705,N_9347,N_9003);
nor U9706 (N_9706,N_9017,N_9372);
nand U9707 (N_9707,N_9345,N_9301);
and U9708 (N_9708,N_9020,N_9269);
or U9709 (N_9709,N_9361,N_9113);
or U9710 (N_9710,N_9284,N_9333);
nand U9711 (N_9711,N_9067,N_9108);
and U9712 (N_9712,N_9426,N_9086);
and U9713 (N_9713,N_9219,N_9182);
or U9714 (N_9714,N_9399,N_9184);
nand U9715 (N_9715,N_9388,N_9479);
nor U9716 (N_9716,N_9099,N_9159);
nand U9717 (N_9717,N_9343,N_9498);
and U9718 (N_9718,N_9279,N_9155);
and U9719 (N_9719,N_9285,N_9211);
nand U9720 (N_9720,N_9033,N_9202);
nand U9721 (N_9721,N_9352,N_9353);
nand U9722 (N_9722,N_9031,N_9268);
nand U9723 (N_9723,N_9163,N_9230);
or U9724 (N_9724,N_9406,N_9257);
nand U9725 (N_9725,N_9007,N_9110);
nor U9726 (N_9726,N_9225,N_9311);
nor U9727 (N_9727,N_9492,N_9205);
nand U9728 (N_9728,N_9111,N_9303);
nand U9729 (N_9729,N_9391,N_9389);
nor U9730 (N_9730,N_9235,N_9499);
nand U9731 (N_9731,N_9432,N_9196);
nand U9732 (N_9732,N_9422,N_9090);
or U9733 (N_9733,N_9250,N_9094);
and U9734 (N_9734,N_9087,N_9329);
and U9735 (N_9735,N_9124,N_9274);
nand U9736 (N_9736,N_9022,N_9156);
nand U9737 (N_9737,N_9385,N_9076);
or U9738 (N_9738,N_9214,N_9203);
nor U9739 (N_9739,N_9106,N_9212);
nor U9740 (N_9740,N_9138,N_9019);
and U9741 (N_9741,N_9085,N_9442);
xnor U9742 (N_9742,N_9208,N_9485);
or U9743 (N_9743,N_9209,N_9483);
nand U9744 (N_9744,N_9443,N_9471);
nand U9745 (N_9745,N_9032,N_9013);
nor U9746 (N_9746,N_9161,N_9112);
and U9747 (N_9747,N_9287,N_9277);
and U9748 (N_9748,N_9413,N_9151);
and U9749 (N_9749,N_9477,N_9132);
nor U9750 (N_9750,N_9491,N_9030);
and U9751 (N_9751,N_9265,N_9103);
and U9752 (N_9752,N_9163,N_9110);
and U9753 (N_9753,N_9398,N_9055);
or U9754 (N_9754,N_9396,N_9061);
nor U9755 (N_9755,N_9151,N_9042);
nand U9756 (N_9756,N_9317,N_9181);
and U9757 (N_9757,N_9201,N_9030);
nand U9758 (N_9758,N_9225,N_9134);
and U9759 (N_9759,N_9233,N_9277);
nand U9760 (N_9760,N_9458,N_9180);
and U9761 (N_9761,N_9350,N_9189);
or U9762 (N_9762,N_9442,N_9462);
or U9763 (N_9763,N_9412,N_9211);
nor U9764 (N_9764,N_9093,N_9124);
nand U9765 (N_9765,N_9297,N_9195);
or U9766 (N_9766,N_9426,N_9028);
nor U9767 (N_9767,N_9440,N_9476);
nand U9768 (N_9768,N_9208,N_9314);
or U9769 (N_9769,N_9089,N_9159);
nand U9770 (N_9770,N_9498,N_9047);
or U9771 (N_9771,N_9035,N_9368);
nand U9772 (N_9772,N_9395,N_9051);
nand U9773 (N_9773,N_9438,N_9182);
nor U9774 (N_9774,N_9195,N_9420);
nor U9775 (N_9775,N_9469,N_9418);
nand U9776 (N_9776,N_9034,N_9457);
and U9777 (N_9777,N_9391,N_9303);
xor U9778 (N_9778,N_9447,N_9112);
xor U9779 (N_9779,N_9492,N_9167);
or U9780 (N_9780,N_9358,N_9454);
nor U9781 (N_9781,N_9026,N_9259);
nor U9782 (N_9782,N_9319,N_9125);
or U9783 (N_9783,N_9059,N_9248);
and U9784 (N_9784,N_9355,N_9447);
nand U9785 (N_9785,N_9301,N_9138);
or U9786 (N_9786,N_9309,N_9048);
or U9787 (N_9787,N_9306,N_9395);
or U9788 (N_9788,N_9412,N_9150);
or U9789 (N_9789,N_9379,N_9275);
or U9790 (N_9790,N_9462,N_9456);
or U9791 (N_9791,N_9419,N_9200);
nand U9792 (N_9792,N_9020,N_9127);
nor U9793 (N_9793,N_9029,N_9231);
nor U9794 (N_9794,N_9384,N_9341);
or U9795 (N_9795,N_9069,N_9429);
nor U9796 (N_9796,N_9100,N_9498);
nor U9797 (N_9797,N_9313,N_9432);
or U9798 (N_9798,N_9072,N_9468);
and U9799 (N_9799,N_9159,N_9065);
or U9800 (N_9800,N_9473,N_9270);
nor U9801 (N_9801,N_9441,N_9404);
nor U9802 (N_9802,N_9042,N_9174);
and U9803 (N_9803,N_9122,N_9077);
and U9804 (N_9804,N_9228,N_9263);
nand U9805 (N_9805,N_9209,N_9192);
nand U9806 (N_9806,N_9347,N_9209);
nor U9807 (N_9807,N_9275,N_9456);
nor U9808 (N_9808,N_9280,N_9120);
xor U9809 (N_9809,N_9086,N_9039);
nand U9810 (N_9810,N_9305,N_9498);
nor U9811 (N_9811,N_9152,N_9399);
or U9812 (N_9812,N_9066,N_9161);
nor U9813 (N_9813,N_9493,N_9191);
nand U9814 (N_9814,N_9436,N_9075);
or U9815 (N_9815,N_9059,N_9142);
nor U9816 (N_9816,N_9387,N_9307);
nor U9817 (N_9817,N_9066,N_9353);
and U9818 (N_9818,N_9426,N_9372);
or U9819 (N_9819,N_9053,N_9459);
and U9820 (N_9820,N_9317,N_9161);
and U9821 (N_9821,N_9335,N_9333);
or U9822 (N_9822,N_9134,N_9171);
or U9823 (N_9823,N_9353,N_9063);
nor U9824 (N_9824,N_9359,N_9090);
nand U9825 (N_9825,N_9105,N_9407);
or U9826 (N_9826,N_9481,N_9229);
and U9827 (N_9827,N_9226,N_9358);
and U9828 (N_9828,N_9258,N_9418);
nand U9829 (N_9829,N_9029,N_9030);
nor U9830 (N_9830,N_9238,N_9133);
and U9831 (N_9831,N_9173,N_9400);
nand U9832 (N_9832,N_9069,N_9345);
and U9833 (N_9833,N_9248,N_9057);
and U9834 (N_9834,N_9452,N_9245);
or U9835 (N_9835,N_9036,N_9372);
nand U9836 (N_9836,N_9078,N_9349);
and U9837 (N_9837,N_9281,N_9026);
nor U9838 (N_9838,N_9184,N_9253);
nor U9839 (N_9839,N_9205,N_9382);
nor U9840 (N_9840,N_9328,N_9399);
nand U9841 (N_9841,N_9405,N_9174);
nand U9842 (N_9842,N_9143,N_9489);
nor U9843 (N_9843,N_9385,N_9022);
nor U9844 (N_9844,N_9343,N_9071);
xor U9845 (N_9845,N_9234,N_9439);
xnor U9846 (N_9846,N_9466,N_9398);
and U9847 (N_9847,N_9018,N_9140);
nand U9848 (N_9848,N_9397,N_9113);
or U9849 (N_9849,N_9357,N_9228);
nor U9850 (N_9850,N_9498,N_9294);
nand U9851 (N_9851,N_9453,N_9143);
or U9852 (N_9852,N_9286,N_9224);
and U9853 (N_9853,N_9307,N_9277);
nor U9854 (N_9854,N_9222,N_9102);
or U9855 (N_9855,N_9133,N_9319);
or U9856 (N_9856,N_9216,N_9409);
or U9857 (N_9857,N_9474,N_9179);
or U9858 (N_9858,N_9241,N_9183);
nand U9859 (N_9859,N_9251,N_9443);
nand U9860 (N_9860,N_9235,N_9127);
and U9861 (N_9861,N_9056,N_9050);
nor U9862 (N_9862,N_9388,N_9119);
xor U9863 (N_9863,N_9267,N_9408);
nand U9864 (N_9864,N_9373,N_9222);
xor U9865 (N_9865,N_9097,N_9221);
nand U9866 (N_9866,N_9312,N_9316);
or U9867 (N_9867,N_9010,N_9403);
or U9868 (N_9868,N_9296,N_9351);
or U9869 (N_9869,N_9262,N_9252);
nand U9870 (N_9870,N_9351,N_9009);
nand U9871 (N_9871,N_9113,N_9240);
nor U9872 (N_9872,N_9407,N_9324);
and U9873 (N_9873,N_9466,N_9493);
nor U9874 (N_9874,N_9189,N_9098);
nand U9875 (N_9875,N_9482,N_9342);
nand U9876 (N_9876,N_9018,N_9022);
nand U9877 (N_9877,N_9219,N_9353);
or U9878 (N_9878,N_9277,N_9192);
or U9879 (N_9879,N_9424,N_9132);
nor U9880 (N_9880,N_9190,N_9455);
and U9881 (N_9881,N_9487,N_9014);
and U9882 (N_9882,N_9268,N_9141);
nor U9883 (N_9883,N_9241,N_9073);
nand U9884 (N_9884,N_9172,N_9430);
nand U9885 (N_9885,N_9183,N_9084);
and U9886 (N_9886,N_9415,N_9484);
nor U9887 (N_9887,N_9280,N_9306);
and U9888 (N_9888,N_9119,N_9108);
nand U9889 (N_9889,N_9084,N_9050);
or U9890 (N_9890,N_9434,N_9310);
and U9891 (N_9891,N_9295,N_9477);
and U9892 (N_9892,N_9121,N_9230);
nor U9893 (N_9893,N_9228,N_9199);
or U9894 (N_9894,N_9024,N_9089);
nand U9895 (N_9895,N_9447,N_9149);
nand U9896 (N_9896,N_9323,N_9272);
and U9897 (N_9897,N_9166,N_9080);
nor U9898 (N_9898,N_9120,N_9308);
and U9899 (N_9899,N_9301,N_9416);
nor U9900 (N_9900,N_9057,N_9062);
nand U9901 (N_9901,N_9177,N_9139);
nor U9902 (N_9902,N_9443,N_9123);
nor U9903 (N_9903,N_9472,N_9190);
and U9904 (N_9904,N_9253,N_9051);
or U9905 (N_9905,N_9013,N_9105);
nor U9906 (N_9906,N_9384,N_9301);
or U9907 (N_9907,N_9466,N_9087);
and U9908 (N_9908,N_9245,N_9054);
nor U9909 (N_9909,N_9466,N_9221);
and U9910 (N_9910,N_9456,N_9242);
nor U9911 (N_9911,N_9431,N_9395);
nor U9912 (N_9912,N_9116,N_9222);
nand U9913 (N_9913,N_9165,N_9128);
nor U9914 (N_9914,N_9128,N_9267);
or U9915 (N_9915,N_9102,N_9030);
or U9916 (N_9916,N_9213,N_9442);
or U9917 (N_9917,N_9415,N_9067);
or U9918 (N_9918,N_9136,N_9385);
nand U9919 (N_9919,N_9355,N_9004);
or U9920 (N_9920,N_9194,N_9295);
nor U9921 (N_9921,N_9413,N_9399);
nor U9922 (N_9922,N_9331,N_9359);
nand U9923 (N_9923,N_9487,N_9455);
or U9924 (N_9924,N_9244,N_9119);
nand U9925 (N_9925,N_9002,N_9055);
nand U9926 (N_9926,N_9262,N_9021);
and U9927 (N_9927,N_9395,N_9485);
or U9928 (N_9928,N_9292,N_9285);
nand U9929 (N_9929,N_9071,N_9408);
nand U9930 (N_9930,N_9305,N_9284);
nor U9931 (N_9931,N_9307,N_9059);
nand U9932 (N_9932,N_9344,N_9203);
nand U9933 (N_9933,N_9434,N_9323);
xnor U9934 (N_9934,N_9263,N_9139);
and U9935 (N_9935,N_9062,N_9142);
nor U9936 (N_9936,N_9217,N_9442);
and U9937 (N_9937,N_9018,N_9321);
nor U9938 (N_9938,N_9195,N_9461);
nor U9939 (N_9939,N_9080,N_9495);
nand U9940 (N_9940,N_9208,N_9442);
and U9941 (N_9941,N_9043,N_9414);
and U9942 (N_9942,N_9313,N_9312);
nor U9943 (N_9943,N_9014,N_9239);
and U9944 (N_9944,N_9231,N_9400);
and U9945 (N_9945,N_9149,N_9089);
nor U9946 (N_9946,N_9467,N_9153);
nor U9947 (N_9947,N_9054,N_9357);
or U9948 (N_9948,N_9145,N_9465);
nor U9949 (N_9949,N_9277,N_9257);
or U9950 (N_9950,N_9495,N_9346);
nor U9951 (N_9951,N_9047,N_9381);
nand U9952 (N_9952,N_9059,N_9284);
or U9953 (N_9953,N_9115,N_9365);
or U9954 (N_9954,N_9151,N_9247);
nand U9955 (N_9955,N_9244,N_9316);
or U9956 (N_9956,N_9221,N_9138);
nor U9957 (N_9957,N_9116,N_9325);
nor U9958 (N_9958,N_9011,N_9478);
and U9959 (N_9959,N_9043,N_9402);
and U9960 (N_9960,N_9349,N_9176);
nor U9961 (N_9961,N_9082,N_9252);
and U9962 (N_9962,N_9318,N_9100);
or U9963 (N_9963,N_9200,N_9461);
nand U9964 (N_9964,N_9029,N_9142);
and U9965 (N_9965,N_9366,N_9010);
and U9966 (N_9966,N_9246,N_9160);
or U9967 (N_9967,N_9133,N_9403);
nor U9968 (N_9968,N_9064,N_9463);
xnor U9969 (N_9969,N_9019,N_9277);
xor U9970 (N_9970,N_9476,N_9310);
nor U9971 (N_9971,N_9433,N_9363);
or U9972 (N_9972,N_9165,N_9353);
and U9973 (N_9973,N_9457,N_9212);
or U9974 (N_9974,N_9141,N_9286);
nand U9975 (N_9975,N_9326,N_9091);
nand U9976 (N_9976,N_9479,N_9141);
nand U9977 (N_9977,N_9424,N_9083);
or U9978 (N_9978,N_9247,N_9257);
nor U9979 (N_9979,N_9477,N_9036);
or U9980 (N_9980,N_9479,N_9347);
and U9981 (N_9981,N_9147,N_9243);
nand U9982 (N_9982,N_9417,N_9156);
and U9983 (N_9983,N_9324,N_9254);
and U9984 (N_9984,N_9284,N_9366);
nor U9985 (N_9985,N_9458,N_9452);
nand U9986 (N_9986,N_9053,N_9407);
nor U9987 (N_9987,N_9060,N_9418);
and U9988 (N_9988,N_9122,N_9169);
and U9989 (N_9989,N_9328,N_9426);
nand U9990 (N_9990,N_9178,N_9477);
or U9991 (N_9991,N_9085,N_9310);
nor U9992 (N_9992,N_9241,N_9049);
and U9993 (N_9993,N_9061,N_9216);
nor U9994 (N_9994,N_9165,N_9461);
xor U9995 (N_9995,N_9234,N_9023);
nand U9996 (N_9996,N_9134,N_9298);
nand U9997 (N_9997,N_9057,N_9264);
nor U9998 (N_9998,N_9059,N_9108);
nor U9999 (N_9999,N_9400,N_9498);
and UO_0 (O_0,N_9537,N_9970);
nand UO_1 (O_1,N_9919,N_9952);
and UO_2 (O_2,N_9555,N_9644);
nor UO_3 (O_3,N_9765,N_9725);
or UO_4 (O_4,N_9639,N_9532);
or UO_5 (O_5,N_9732,N_9674);
nor UO_6 (O_6,N_9773,N_9764);
or UO_7 (O_7,N_9958,N_9727);
nor UO_8 (O_8,N_9813,N_9662);
or UO_9 (O_9,N_9770,N_9801);
or UO_10 (O_10,N_9956,N_9830);
nor UO_11 (O_11,N_9720,N_9609);
nand UO_12 (O_12,N_9802,N_9516);
and UO_13 (O_13,N_9832,N_9972);
and UO_14 (O_14,N_9619,N_9892);
nand UO_15 (O_15,N_9845,N_9723);
and UO_16 (O_16,N_9736,N_9811);
nand UO_17 (O_17,N_9545,N_9640);
and UO_18 (O_18,N_9763,N_9594);
nand UO_19 (O_19,N_9940,N_9617);
nand UO_20 (O_20,N_9935,N_9843);
and UO_21 (O_21,N_9611,N_9547);
or UO_22 (O_22,N_9580,N_9641);
and UO_23 (O_23,N_9601,N_9597);
or UO_24 (O_24,N_9914,N_9598);
nor UO_25 (O_25,N_9932,N_9896);
nor UO_26 (O_26,N_9954,N_9867);
and UO_27 (O_27,N_9792,N_9837);
and UO_28 (O_28,N_9777,N_9904);
or UO_29 (O_29,N_9925,N_9587);
or UO_30 (O_30,N_9719,N_9791);
nand UO_31 (O_31,N_9689,N_9924);
nand UO_32 (O_32,N_9694,N_9602);
nand UO_33 (O_33,N_9766,N_9751);
and UO_34 (O_34,N_9968,N_9873);
xnor UO_35 (O_35,N_9746,N_9680);
nand UO_36 (O_36,N_9683,N_9558);
nand UO_37 (O_37,N_9629,N_9561);
and UO_38 (O_38,N_9739,N_9949);
and UO_39 (O_39,N_9622,N_9649);
nor UO_40 (O_40,N_9897,N_9983);
nand UO_41 (O_41,N_9964,N_9755);
and UO_42 (O_42,N_9578,N_9960);
or UO_43 (O_43,N_9633,N_9752);
nor UO_44 (O_44,N_9535,N_9572);
nor UO_45 (O_45,N_9818,N_9543);
nand UO_46 (O_46,N_9973,N_9544);
and UO_47 (O_47,N_9772,N_9605);
and UO_48 (O_48,N_9750,N_9655);
nand UO_49 (O_49,N_9666,N_9610);
and UO_50 (O_50,N_9980,N_9953);
or UO_51 (O_51,N_9883,N_9875);
nand UO_52 (O_52,N_9583,N_9786);
or UO_53 (O_53,N_9709,N_9806);
and UO_54 (O_54,N_9685,N_9691);
nor UO_55 (O_55,N_9592,N_9887);
nor UO_56 (O_56,N_9513,N_9955);
nor UO_57 (O_57,N_9877,N_9730);
or UO_58 (O_58,N_9638,N_9745);
or UO_59 (O_59,N_9963,N_9695);
or UO_60 (O_60,N_9567,N_9876);
and UO_61 (O_61,N_9621,N_9618);
nor UO_62 (O_62,N_9826,N_9705);
nor UO_63 (O_63,N_9804,N_9581);
or UO_64 (O_64,N_9500,N_9635);
and UO_65 (O_65,N_9501,N_9945);
or UO_66 (O_66,N_9737,N_9616);
or UO_67 (O_67,N_9686,N_9993);
and UO_68 (O_68,N_9760,N_9626);
nor UO_69 (O_69,N_9827,N_9878);
nand UO_70 (O_70,N_9679,N_9862);
nand UO_71 (O_71,N_9969,N_9508);
nand UO_72 (O_72,N_9669,N_9866);
nand UO_73 (O_73,N_9743,N_9756);
or UO_74 (O_74,N_9560,N_9754);
and UO_75 (O_75,N_9762,N_9967);
nand UO_76 (O_76,N_9753,N_9790);
and UO_77 (O_77,N_9823,N_9821);
and UO_78 (O_78,N_9902,N_9589);
and UO_79 (O_79,N_9844,N_9657);
nand UO_80 (O_80,N_9533,N_9828);
nor UO_81 (O_81,N_9808,N_9509);
nand UO_82 (O_82,N_9539,N_9631);
nand UO_83 (O_83,N_9659,N_9779);
or UO_84 (O_84,N_9985,N_9645);
nor UO_85 (O_85,N_9591,N_9707);
nor UO_86 (O_86,N_9849,N_9898);
and UO_87 (O_87,N_9907,N_9521);
nand UO_88 (O_88,N_9950,N_9671);
and UO_89 (O_89,N_9652,N_9554);
nand UO_90 (O_90,N_9556,N_9624);
and UO_91 (O_91,N_9549,N_9787);
and UO_92 (O_92,N_9824,N_9894);
and UO_93 (O_93,N_9913,N_9568);
nor UO_94 (O_94,N_9809,N_9653);
or UO_95 (O_95,N_9724,N_9929);
and UO_96 (O_96,N_9510,N_9576);
or UO_97 (O_97,N_9614,N_9978);
and UO_98 (O_98,N_9825,N_9901);
and UO_99 (O_99,N_9872,N_9584);
or UO_100 (O_100,N_9884,N_9620);
nor UO_101 (O_101,N_9735,N_9951);
and UO_102 (O_102,N_9998,N_9820);
nand UO_103 (O_103,N_9987,N_9548);
and UO_104 (O_104,N_9740,N_9852);
or UO_105 (O_105,N_9651,N_9630);
and UO_106 (O_106,N_9915,N_9793);
nor UO_107 (O_107,N_9923,N_9771);
nor UO_108 (O_108,N_9857,N_9710);
or UO_109 (O_109,N_9934,N_9517);
nand UO_110 (O_110,N_9822,N_9522);
or UO_111 (O_111,N_9526,N_9780);
or UO_112 (O_112,N_9899,N_9704);
or UO_113 (O_113,N_9895,N_9658);
or UO_114 (O_114,N_9678,N_9854);
nand UO_115 (O_115,N_9979,N_9853);
or UO_116 (O_116,N_9984,N_9569);
nand UO_117 (O_117,N_9713,N_9975);
and UO_118 (O_118,N_9603,N_9856);
nand UO_119 (O_119,N_9858,N_9906);
xnor UO_120 (O_120,N_9749,N_9938);
nor UO_121 (O_121,N_9926,N_9841);
or UO_122 (O_122,N_9829,N_9722);
and UO_123 (O_123,N_9868,N_9927);
and UO_124 (O_124,N_9846,N_9675);
or UO_125 (O_125,N_9976,N_9700);
or UO_126 (O_126,N_9885,N_9636);
or UO_127 (O_127,N_9921,N_9928);
or UO_128 (O_128,N_9997,N_9784);
nand UO_129 (O_129,N_9504,N_9552);
nor UO_130 (O_130,N_9733,N_9982);
or UO_131 (O_131,N_9660,N_9738);
and UO_132 (O_132,N_9870,N_9566);
nand UO_133 (O_133,N_9536,N_9531);
nand UO_134 (O_134,N_9797,N_9816);
nand UO_135 (O_135,N_9986,N_9865);
or UO_136 (O_136,N_9550,N_9965);
nand UO_137 (O_137,N_9959,N_9718);
and UO_138 (O_138,N_9668,N_9893);
and UO_139 (O_139,N_9528,N_9527);
nand UO_140 (O_140,N_9726,N_9687);
or UO_141 (O_141,N_9551,N_9595);
nor UO_142 (O_142,N_9988,N_9646);
nand UO_143 (O_143,N_9703,N_9812);
or UO_144 (O_144,N_9590,N_9661);
and UO_145 (O_145,N_9530,N_9788);
nand UO_146 (O_146,N_9514,N_9848);
or UO_147 (O_147,N_9995,N_9803);
nand UO_148 (O_148,N_9847,N_9775);
and UO_149 (O_149,N_9615,N_9918);
nor UO_150 (O_150,N_9701,N_9564);
and UO_151 (O_151,N_9708,N_9992);
and UO_152 (O_152,N_9839,N_9664);
nand UO_153 (O_153,N_9861,N_9627);
and UO_154 (O_154,N_9946,N_9831);
nor UO_155 (O_155,N_9936,N_9942);
or UO_156 (O_156,N_9905,N_9761);
nand UO_157 (O_157,N_9922,N_9903);
nand UO_158 (O_158,N_9684,N_9795);
nand UO_159 (O_159,N_9596,N_9721);
nand UO_160 (O_160,N_9717,N_9604);
nor UO_161 (O_161,N_9943,N_9647);
nor UO_162 (O_162,N_9758,N_9769);
nor UO_163 (O_163,N_9891,N_9742);
and UO_164 (O_164,N_9912,N_9570);
and UO_165 (O_165,N_9667,N_9542);
xnor UO_166 (O_166,N_9608,N_9835);
nor UO_167 (O_167,N_9511,N_9890);
nor UO_168 (O_168,N_9814,N_9833);
or UO_169 (O_169,N_9505,N_9512);
and UO_170 (O_170,N_9523,N_9520);
nand UO_171 (O_171,N_9663,N_9706);
and UO_172 (O_172,N_9794,N_9881);
nand UO_173 (O_173,N_9637,N_9991);
nor UO_174 (O_174,N_9502,N_9879);
or UO_175 (O_175,N_9634,N_9933);
nand UO_176 (O_176,N_9506,N_9757);
and UO_177 (O_177,N_9728,N_9961);
nor UO_178 (O_178,N_9916,N_9586);
nand UO_179 (O_179,N_9747,N_9799);
and UO_180 (O_180,N_9716,N_9889);
nor UO_181 (O_181,N_9677,N_9920);
nand UO_182 (O_182,N_9529,N_9702);
or UO_183 (O_183,N_9698,N_9930);
and UO_184 (O_184,N_9948,N_9990);
and UO_185 (O_185,N_9999,N_9748);
nor UO_186 (O_186,N_9682,N_9600);
nand UO_187 (O_187,N_9957,N_9800);
nor UO_188 (O_188,N_9782,N_9874);
nor UO_189 (O_189,N_9941,N_9642);
nand UO_190 (O_190,N_9575,N_9688);
nor UO_191 (O_191,N_9908,N_9966);
and UO_192 (O_192,N_9783,N_9917);
nor UO_193 (O_193,N_9863,N_9625);
nor UO_194 (O_194,N_9673,N_9785);
xnor UO_195 (O_195,N_9851,N_9562);
nand UO_196 (O_196,N_9729,N_9503);
nor UO_197 (O_197,N_9909,N_9778);
or UO_198 (O_198,N_9944,N_9815);
or UO_199 (O_199,N_9768,N_9534);
or UO_200 (O_200,N_9911,N_9518);
nor UO_201 (O_201,N_9643,N_9971);
nand UO_202 (O_202,N_9697,N_9859);
xnor UO_203 (O_203,N_9886,N_9774);
nand UO_204 (O_204,N_9676,N_9996);
or UO_205 (O_205,N_9546,N_9654);
nand UO_206 (O_206,N_9541,N_9507);
or UO_207 (O_207,N_9789,N_9540);
nand UO_208 (O_208,N_9681,N_9559);
or UO_209 (O_209,N_9515,N_9632);
nand UO_210 (O_210,N_9994,N_9693);
and UO_211 (O_211,N_9744,N_9690);
nor UO_212 (O_212,N_9810,N_9981);
nand UO_213 (O_213,N_9714,N_9612);
nand UO_214 (O_214,N_9807,N_9665);
nor UO_215 (O_215,N_9962,N_9977);
and UO_216 (O_216,N_9672,N_9579);
nand UO_217 (O_217,N_9798,N_9553);
or UO_218 (O_218,N_9871,N_9692);
and UO_219 (O_219,N_9588,N_9931);
and UO_220 (O_220,N_9571,N_9880);
and UO_221 (O_221,N_9699,N_9573);
and UO_222 (O_222,N_9613,N_9767);
nand UO_223 (O_223,N_9577,N_9711);
or UO_224 (O_224,N_9648,N_9607);
or UO_225 (O_225,N_9656,N_9606);
and UO_226 (O_226,N_9599,N_9805);
and UO_227 (O_227,N_9989,N_9628);
or UO_228 (O_228,N_9937,N_9819);
and UO_229 (O_229,N_9731,N_9593);
nand UO_230 (O_230,N_9574,N_9563);
and UO_231 (O_231,N_9670,N_9538);
nor UO_232 (O_232,N_9585,N_9869);
or UO_233 (O_233,N_9817,N_9524);
or UO_234 (O_234,N_9864,N_9900);
nor UO_235 (O_235,N_9947,N_9850);
or UO_236 (O_236,N_9734,N_9840);
nor UO_237 (O_237,N_9741,N_9939);
nand UO_238 (O_238,N_9525,N_9882);
and UO_239 (O_239,N_9838,N_9557);
nand UO_240 (O_240,N_9855,N_9759);
and UO_241 (O_241,N_9715,N_9696);
and UO_242 (O_242,N_9781,N_9565);
and UO_243 (O_243,N_9519,N_9836);
or UO_244 (O_244,N_9834,N_9582);
and UO_245 (O_245,N_9776,N_9712);
or UO_246 (O_246,N_9910,N_9650);
or UO_247 (O_247,N_9623,N_9842);
nor UO_248 (O_248,N_9888,N_9860);
and UO_249 (O_249,N_9796,N_9974);
nand UO_250 (O_250,N_9818,N_9808);
and UO_251 (O_251,N_9900,N_9612);
xnor UO_252 (O_252,N_9541,N_9780);
nor UO_253 (O_253,N_9777,N_9599);
or UO_254 (O_254,N_9705,N_9942);
or UO_255 (O_255,N_9571,N_9753);
or UO_256 (O_256,N_9911,N_9564);
nor UO_257 (O_257,N_9922,N_9971);
nand UO_258 (O_258,N_9634,N_9908);
xnor UO_259 (O_259,N_9754,N_9537);
or UO_260 (O_260,N_9824,N_9530);
nand UO_261 (O_261,N_9628,N_9623);
or UO_262 (O_262,N_9989,N_9940);
and UO_263 (O_263,N_9631,N_9950);
nor UO_264 (O_264,N_9898,N_9705);
or UO_265 (O_265,N_9753,N_9748);
and UO_266 (O_266,N_9717,N_9935);
or UO_267 (O_267,N_9511,N_9948);
and UO_268 (O_268,N_9697,N_9850);
and UO_269 (O_269,N_9842,N_9690);
nor UO_270 (O_270,N_9686,N_9540);
xor UO_271 (O_271,N_9711,N_9852);
and UO_272 (O_272,N_9557,N_9639);
or UO_273 (O_273,N_9580,N_9646);
or UO_274 (O_274,N_9646,N_9507);
or UO_275 (O_275,N_9545,N_9793);
nand UO_276 (O_276,N_9940,N_9967);
or UO_277 (O_277,N_9628,N_9543);
or UO_278 (O_278,N_9931,N_9893);
nand UO_279 (O_279,N_9667,N_9928);
nand UO_280 (O_280,N_9768,N_9623);
nor UO_281 (O_281,N_9941,N_9699);
nand UO_282 (O_282,N_9990,N_9825);
nand UO_283 (O_283,N_9710,N_9792);
nor UO_284 (O_284,N_9510,N_9807);
nor UO_285 (O_285,N_9532,N_9777);
nor UO_286 (O_286,N_9848,N_9516);
and UO_287 (O_287,N_9728,N_9765);
and UO_288 (O_288,N_9582,N_9575);
nor UO_289 (O_289,N_9730,N_9949);
nor UO_290 (O_290,N_9906,N_9872);
xnor UO_291 (O_291,N_9690,N_9895);
nor UO_292 (O_292,N_9834,N_9852);
and UO_293 (O_293,N_9728,N_9551);
nand UO_294 (O_294,N_9527,N_9592);
or UO_295 (O_295,N_9599,N_9603);
and UO_296 (O_296,N_9829,N_9551);
nand UO_297 (O_297,N_9921,N_9777);
nor UO_298 (O_298,N_9781,N_9725);
nand UO_299 (O_299,N_9698,N_9979);
nand UO_300 (O_300,N_9502,N_9683);
and UO_301 (O_301,N_9691,N_9763);
or UO_302 (O_302,N_9918,N_9712);
nand UO_303 (O_303,N_9664,N_9538);
nand UO_304 (O_304,N_9649,N_9998);
nor UO_305 (O_305,N_9827,N_9633);
nor UO_306 (O_306,N_9530,N_9844);
or UO_307 (O_307,N_9929,N_9948);
xnor UO_308 (O_308,N_9809,N_9669);
nand UO_309 (O_309,N_9879,N_9708);
or UO_310 (O_310,N_9953,N_9947);
nor UO_311 (O_311,N_9652,N_9827);
nor UO_312 (O_312,N_9724,N_9536);
nor UO_313 (O_313,N_9501,N_9813);
and UO_314 (O_314,N_9716,N_9827);
nand UO_315 (O_315,N_9974,N_9835);
nor UO_316 (O_316,N_9777,N_9568);
nand UO_317 (O_317,N_9671,N_9500);
nor UO_318 (O_318,N_9851,N_9739);
or UO_319 (O_319,N_9883,N_9544);
or UO_320 (O_320,N_9642,N_9539);
and UO_321 (O_321,N_9764,N_9670);
nand UO_322 (O_322,N_9713,N_9840);
xnor UO_323 (O_323,N_9504,N_9808);
or UO_324 (O_324,N_9799,N_9575);
nor UO_325 (O_325,N_9835,N_9876);
nand UO_326 (O_326,N_9579,N_9843);
nor UO_327 (O_327,N_9572,N_9967);
nand UO_328 (O_328,N_9778,N_9895);
and UO_329 (O_329,N_9591,N_9752);
nand UO_330 (O_330,N_9607,N_9857);
and UO_331 (O_331,N_9557,N_9672);
nor UO_332 (O_332,N_9656,N_9576);
nand UO_333 (O_333,N_9896,N_9877);
or UO_334 (O_334,N_9503,N_9997);
or UO_335 (O_335,N_9728,N_9880);
nor UO_336 (O_336,N_9516,N_9569);
or UO_337 (O_337,N_9843,N_9502);
nand UO_338 (O_338,N_9960,N_9950);
and UO_339 (O_339,N_9866,N_9555);
or UO_340 (O_340,N_9708,N_9558);
nand UO_341 (O_341,N_9754,N_9962);
or UO_342 (O_342,N_9933,N_9908);
or UO_343 (O_343,N_9889,N_9922);
nand UO_344 (O_344,N_9702,N_9700);
and UO_345 (O_345,N_9526,N_9933);
nor UO_346 (O_346,N_9609,N_9559);
and UO_347 (O_347,N_9791,N_9585);
nand UO_348 (O_348,N_9614,N_9773);
nor UO_349 (O_349,N_9688,N_9696);
nor UO_350 (O_350,N_9580,N_9925);
nand UO_351 (O_351,N_9985,N_9860);
nor UO_352 (O_352,N_9586,N_9517);
or UO_353 (O_353,N_9602,N_9833);
and UO_354 (O_354,N_9882,N_9906);
or UO_355 (O_355,N_9732,N_9815);
or UO_356 (O_356,N_9748,N_9528);
nand UO_357 (O_357,N_9994,N_9723);
nand UO_358 (O_358,N_9676,N_9874);
nor UO_359 (O_359,N_9516,N_9969);
xnor UO_360 (O_360,N_9847,N_9967);
and UO_361 (O_361,N_9599,N_9535);
nand UO_362 (O_362,N_9764,N_9822);
nand UO_363 (O_363,N_9588,N_9729);
and UO_364 (O_364,N_9859,N_9617);
or UO_365 (O_365,N_9891,N_9676);
nand UO_366 (O_366,N_9988,N_9947);
and UO_367 (O_367,N_9956,N_9528);
and UO_368 (O_368,N_9939,N_9756);
nand UO_369 (O_369,N_9669,N_9559);
or UO_370 (O_370,N_9996,N_9816);
or UO_371 (O_371,N_9759,N_9893);
xnor UO_372 (O_372,N_9908,N_9734);
and UO_373 (O_373,N_9964,N_9852);
and UO_374 (O_374,N_9884,N_9855);
or UO_375 (O_375,N_9926,N_9574);
nor UO_376 (O_376,N_9639,N_9640);
nor UO_377 (O_377,N_9771,N_9791);
or UO_378 (O_378,N_9511,N_9616);
or UO_379 (O_379,N_9892,N_9957);
nor UO_380 (O_380,N_9809,N_9977);
and UO_381 (O_381,N_9960,N_9712);
and UO_382 (O_382,N_9877,N_9638);
nand UO_383 (O_383,N_9965,N_9702);
or UO_384 (O_384,N_9854,N_9527);
and UO_385 (O_385,N_9871,N_9636);
and UO_386 (O_386,N_9774,N_9748);
and UO_387 (O_387,N_9607,N_9783);
nor UO_388 (O_388,N_9860,N_9967);
or UO_389 (O_389,N_9550,N_9504);
nor UO_390 (O_390,N_9814,N_9798);
and UO_391 (O_391,N_9776,N_9800);
nor UO_392 (O_392,N_9557,N_9506);
nand UO_393 (O_393,N_9846,N_9640);
or UO_394 (O_394,N_9663,N_9606);
and UO_395 (O_395,N_9515,N_9514);
nor UO_396 (O_396,N_9510,N_9828);
and UO_397 (O_397,N_9709,N_9814);
nor UO_398 (O_398,N_9540,N_9831);
nor UO_399 (O_399,N_9771,N_9646);
and UO_400 (O_400,N_9899,N_9931);
nand UO_401 (O_401,N_9540,N_9912);
and UO_402 (O_402,N_9541,N_9625);
and UO_403 (O_403,N_9879,N_9594);
or UO_404 (O_404,N_9915,N_9918);
and UO_405 (O_405,N_9651,N_9570);
nand UO_406 (O_406,N_9806,N_9674);
nor UO_407 (O_407,N_9696,N_9866);
nor UO_408 (O_408,N_9998,N_9682);
nor UO_409 (O_409,N_9859,N_9992);
nor UO_410 (O_410,N_9810,N_9714);
and UO_411 (O_411,N_9812,N_9935);
nor UO_412 (O_412,N_9971,N_9703);
and UO_413 (O_413,N_9776,N_9964);
and UO_414 (O_414,N_9689,N_9748);
nand UO_415 (O_415,N_9983,N_9971);
nand UO_416 (O_416,N_9941,N_9925);
and UO_417 (O_417,N_9542,N_9648);
nor UO_418 (O_418,N_9828,N_9743);
xnor UO_419 (O_419,N_9515,N_9705);
or UO_420 (O_420,N_9638,N_9943);
xor UO_421 (O_421,N_9833,N_9966);
nor UO_422 (O_422,N_9577,N_9651);
and UO_423 (O_423,N_9759,N_9649);
nand UO_424 (O_424,N_9827,N_9506);
nor UO_425 (O_425,N_9653,N_9760);
and UO_426 (O_426,N_9780,N_9894);
or UO_427 (O_427,N_9954,N_9832);
and UO_428 (O_428,N_9866,N_9888);
or UO_429 (O_429,N_9955,N_9759);
nor UO_430 (O_430,N_9853,N_9998);
nand UO_431 (O_431,N_9824,N_9508);
and UO_432 (O_432,N_9962,N_9586);
nand UO_433 (O_433,N_9922,N_9654);
nand UO_434 (O_434,N_9898,N_9967);
and UO_435 (O_435,N_9986,N_9715);
nand UO_436 (O_436,N_9917,N_9869);
nor UO_437 (O_437,N_9523,N_9734);
or UO_438 (O_438,N_9656,N_9981);
nor UO_439 (O_439,N_9825,N_9846);
or UO_440 (O_440,N_9502,N_9587);
nor UO_441 (O_441,N_9891,N_9846);
nor UO_442 (O_442,N_9576,N_9692);
or UO_443 (O_443,N_9633,N_9716);
or UO_444 (O_444,N_9566,N_9586);
nor UO_445 (O_445,N_9945,N_9825);
nor UO_446 (O_446,N_9994,N_9641);
and UO_447 (O_447,N_9975,N_9778);
and UO_448 (O_448,N_9686,N_9745);
nand UO_449 (O_449,N_9910,N_9673);
nand UO_450 (O_450,N_9951,N_9645);
nor UO_451 (O_451,N_9999,N_9997);
or UO_452 (O_452,N_9913,N_9918);
nor UO_453 (O_453,N_9589,N_9574);
xnor UO_454 (O_454,N_9806,N_9748);
or UO_455 (O_455,N_9985,N_9547);
nor UO_456 (O_456,N_9904,N_9608);
and UO_457 (O_457,N_9641,N_9538);
nor UO_458 (O_458,N_9894,N_9577);
and UO_459 (O_459,N_9873,N_9687);
and UO_460 (O_460,N_9872,N_9588);
and UO_461 (O_461,N_9586,N_9524);
nor UO_462 (O_462,N_9689,N_9523);
and UO_463 (O_463,N_9621,N_9993);
and UO_464 (O_464,N_9605,N_9810);
and UO_465 (O_465,N_9870,N_9638);
nand UO_466 (O_466,N_9956,N_9518);
nor UO_467 (O_467,N_9744,N_9856);
nand UO_468 (O_468,N_9862,N_9928);
or UO_469 (O_469,N_9882,N_9594);
and UO_470 (O_470,N_9736,N_9851);
nand UO_471 (O_471,N_9993,N_9580);
or UO_472 (O_472,N_9848,N_9685);
nand UO_473 (O_473,N_9584,N_9797);
nor UO_474 (O_474,N_9778,N_9766);
or UO_475 (O_475,N_9501,N_9726);
or UO_476 (O_476,N_9818,N_9599);
and UO_477 (O_477,N_9638,N_9505);
or UO_478 (O_478,N_9661,N_9869);
nand UO_479 (O_479,N_9989,N_9767);
nor UO_480 (O_480,N_9544,N_9747);
and UO_481 (O_481,N_9718,N_9655);
nand UO_482 (O_482,N_9699,N_9787);
nand UO_483 (O_483,N_9650,N_9681);
nand UO_484 (O_484,N_9661,N_9553);
and UO_485 (O_485,N_9807,N_9508);
and UO_486 (O_486,N_9814,N_9532);
nand UO_487 (O_487,N_9888,N_9751);
nor UO_488 (O_488,N_9787,N_9909);
xnor UO_489 (O_489,N_9839,N_9610);
or UO_490 (O_490,N_9852,N_9547);
nor UO_491 (O_491,N_9511,N_9633);
nor UO_492 (O_492,N_9999,N_9812);
nand UO_493 (O_493,N_9872,N_9939);
nor UO_494 (O_494,N_9619,N_9797);
and UO_495 (O_495,N_9518,N_9606);
nor UO_496 (O_496,N_9629,N_9729);
nand UO_497 (O_497,N_9979,N_9508);
nor UO_498 (O_498,N_9577,N_9899);
nor UO_499 (O_499,N_9594,N_9521);
nor UO_500 (O_500,N_9567,N_9801);
and UO_501 (O_501,N_9732,N_9617);
or UO_502 (O_502,N_9781,N_9917);
or UO_503 (O_503,N_9547,N_9726);
or UO_504 (O_504,N_9810,N_9666);
nand UO_505 (O_505,N_9821,N_9876);
nor UO_506 (O_506,N_9639,N_9536);
nand UO_507 (O_507,N_9557,N_9552);
nand UO_508 (O_508,N_9716,N_9603);
nand UO_509 (O_509,N_9507,N_9604);
and UO_510 (O_510,N_9736,N_9989);
nand UO_511 (O_511,N_9933,N_9856);
and UO_512 (O_512,N_9945,N_9587);
nand UO_513 (O_513,N_9553,N_9527);
and UO_514 (O_514,N_9665,N_9990);
and UO_515 (O_515,N_9800,N_9904);
or UO_516 (O_516,N_9572,N_9605);
nor UO_517 (O_517,N_9868,N_9566);
and UO_518 (O_518,N_9845,N_9739);
or UO_519 (O_519,N_9807,N_9820);
and UO_520 (O_520,N_9879,N_9617);
nand UO_521 (O_521,N_9852,N_9853);
and UO_522 (O_522,N_9876,N_9676);
and UO_523 (O_523,N_9873,N_9961);
and UO_524 (O_524,N_9655,N_9701);
nor UO_525 (O_525,N_9540,N_9885);
or UO_526 (O_526,N_9793,N_9623);
nor UO_527 (O_527,N_9960,N_9681);
or UO_528 (O_528,N_9986,N_9513);
nor UO_529 (O_529,N_9888,N_9941);
nor UO_530 (O_530,N_9871,N_9962);
or UO_531 (O_531,N_9916,N_9688);
nand UO_532 (O_532,N_9681,N_9519);
nand UO_533 (O_533,N_9997,N_9634);
and UO_534 (O_534,N_9864,N_9910);
nor UO_535 (O_535,N_9856,N_9589);
nor UO_536 (O_536,N_9726,N_9816);
nor UO_537 (O_537,N_9579,N_9521);
and UO_538 (O_538,N_9753,N_9639);
or UO_539 (O_539,N_9805,N_9612);
and UO_540 (O_540,N_9753,N_9833);
or UO_541 (O_541,N_9717,N_9640);
nor UO_542 (O_542,N_9690,N_9638);
and UO_543 (O_543,N_9545,N_9515);
or UO_544 (O_544,N_9714,N_9517);
nor UO_545 (O_545,N_9859,N_9570);
nor UO_546 (O_546,N_9876,N_9581);
nor UO_547 (O_547,N_9537,N_9504);
xnor UO_548 (O_548,N_9777,N_9889);
nor UO_549 (O_549,N_9807,N_9727);
nor UO_550 (O_550,N_9965,N_9737);
or UO_551 (O_551,N_9766,N_9581);
nor UO_552 (O_552,N_9865,N_9532);
or UO_553 (O_553,N_9968,N_9646);
or UO_554 (O_554,N_9962,N_9601);
xor UO_555 (O_555,N_9961,N_9593);
and UO_556 (O_556,N_9895,N_9882);
nand UO_557 (O_557,N_9759,N_9920);
nor UO_558 (O_558,N_9630,N_9977);
or UO_559 (O_559,N_9952,N_9856);
and UO_560 (O_560,N_9571,N_9797);
nor UO_561 (O_561,N_9563,N_9727);
nand UO_562 (O_562,N_9857,N_9929);
and UO_563 (O_563,N_9769,N_9863);
and UO_564 (O_564,N_9913,N_9639);
nor UO_565 (O_565,N_9853,N_9655);
or UO_566 (O_566,N_9996,N_9560);
nor UO_567 (O_567,N_9629,N_9951);
nand UO_568 (O_568,N_9672,N_9832);
or UO_569 (O_569,N_9946,N_9947);
and UO_570 (O_570,N_9928,N_9941);
and UO_571 (O_571,N_9811,N_9545);
and UO_572 (O_572,N_9982,N_9561);
and UO_573 (O_573,N_9854,N_9669);
or UO_574 (O_574,N_9565,N_9541);
and UO_575 (O_575,N_9600,N_9870);
and UO_576 (O_576,N_9657,N_9783);
nand UO_577 (O_577,N_9753,N_9890);
or UO_578 (O_578,N_9692,N_9990);
and UO_579 (O_579,N_9634,N_9503);
or UO_580 (O_580,N_9922,N_9955);
or UO_581 (O_581,N_9901,N_9603);
nand UO_582 (O_582,N_9998,N_9985);
and UO_583 (O_583,N_9745,N_9564);
and UO_584 (O_584,N_9985,N_9987);
nand UO_585 (O_585,N_9767,N_9651);
nand UO_586 (O_586,N_9849,N_9823);
or UO_587 (O_587,N_9910,N_9881);
nor UO_588 (O_588,N_9749,N_9926);
nand UO_589 (O_589,N_9636,N_9774);
or UO_590 (O_590,N_9729,N_9648);
nor UO_591 (O_591,N_9565,N_9555);
nand UO_592 (O_592,N_9958,N_9762);
nand UO_593 (O_593,N_9571,N_9959);
nor UO_594 (O_594,N_9513,N_9833);
nor UO_595 (O_595,N_9541,N_9576);
nand UO_596 (O_596,N_9832,N_9934);
nor UO_597 (O_597,N_9935,N_9531);
nand UO_598 (O_598,N_9952,N_9864);
and UO_599 (O_599,N_9556,N_9500);
xor UO_600 (O_600,N_9619,N_9810);
nand UO_601 (O_601,N_9767,N_9704);
nor UO_602 (O_602,N_9836,N_9914);
nand UO_603 (O_603,N_9901,N_9515);
and UO_604 (O_604,N_9799,N_9791);
nor UO_605 (O_605,N_9600,N_9587);
nor UO_606 (O_606,N_9847,N_9976);
nor UO_607 (O_607,N_9866,N_9947);
or UO_608 (O_608,N_9693,N_9855);
nand UO_609 (O_609,N_9835,N_9664);
or UO_610 (O_610,N_9564,N_9530);
nor UO_611 (O_611,N_9687,N_9644);
and UO_612 (O_612,N_9928,N_9721);
or UO_613 (O_613,N_9897,N_9702);
nor UO_614 (O_614,N_9737,N_9584);
nand UO_615 (O_615,N_9620,N_9661);
and UO_616 (O_616,N_9763,N_9664);
or UO_617 (O_617,N_9619,N_9745);
or UO_618 (O_618,N_9682,N_9714);
and UO_619 (O_619,N_9523,N_9746);
or UO_620 (O_620,N_9543,N_9967);
or UO_621 (O_621,N_9516,N_9677);
and UO_622 (O_622,N_9632,N_9585);
and UO_623 (O_623,N_9804,N_9604);
nand UO_624 (O_624,N_9790,N_9979);
and UO_625 (O_625,N_9720,N_9850);
nor UO_626 (O_626,N_9729,N_9515);
nor UO_627 (O_627,N_9895,N_9899);
nand UO_628 (O_628,N_9686,N_9607);
and UO_629 (O_629,N_9920,N_9510);
and UO_630 (O_630,N_9573,N_9908);
and UO_631 (O_631,N_9925,N_9634);
and UO_632 (O_632,N_9689,N_9992);
and UO_633 (O_633,N_9524,N_9916);
nand UO_634 (O_634,N_9901,N_9943);
nor UO_635 (O_635,N_9831,N_9763);
nand UO_636 (O_636,N_9785,N_9592);
or UO_637 (O_637,N_9644,N_9549);
nand UO_638 (O_638,N_9809,N_9631);
xor UO_639 (O_639,N_9801,N_9831);
or UO_640 (O_640,N_9593,N_9883);
nor UO_641 (O_641,N_9941,N_9660);
nand UO_642 (O_642,N_9945,N_9829);
or UO_643 (O_643,N_9521,N_9754);
or UO_644 (O_644,N_9772,N_9999);
or UO_645 (O_645,N_9926,N_9995);
nand UO_646 (O_646,N_9523,N_9860);
nor UO_647 (O_647,N_9507,N_9947);
nor UO_648 (O_648,N_9729,N_9889);
or UO_649 (O_649,N_9880,N_9801);
or UO_650 (O_650,N_9758,N_9594);
nand UO_651 (O_651,N_9573,N_9509);
nor UO_652 (O_652,N_9894,N_9688);
nor UO_653 (O_653,N_9751,N_9864);
nand UO_654 (O_654,N_9640,N_9949);
nor UO_655 (O_655,N_9660,N_9616);
or UO_656 (O_656,N_9539,N_9590);
nand UO_657 (O_657,N_9566,N_9957);
nand UO_658 (O_658,N_9531,N_9581);
xor UO_659 (O_659,N_9736,N_9612);
and UO_660 (O_660,N_9933,N_9757);
nand UO_661 (O_661,N_9712,N_9917);
or UO_662 (O_662,N_9727,N_9864);
and UO_663 (O_663,N_9681,N_9572);
or UO_664 (O_664,N_9556,N_9926);
or UO_665 (O_665,N_9634,N_9841);
or UO_666 (O_666,N_9929,N_9753);
or UO_667 (O_667,N_9979,N_9767);
or UO_668 (O_668,N_9938,N_9630);
nor UO_669 (O_669,N_9566,N_9635);
and UO_670 (O_670,N_9893,N_9849);
or UO_671 (O_671,N_9530,N_9711);
nor UO_672 (O_672,N_9595,N_9531);
and UO_673 (O_673,N_9561,N_9644);
or UO_674 (O_674,N_9631,N_9890);
xnor UO_675 (O_675,N_9863,N_9502);
nor UO_676 (O_676,N_9968,N_9792);
xor UO_677 (O_677,N_9627,N_9531);
nor UO_678 (O_678,N_9584,N_9843);
or UO_679 (O_679,N_9834,N_9924);
nor UO_680 (O_680,N_9533,N_9921);
nor UO_681 (O_681,N_9810,N_9914);
or UO_682 (O_682,N_9761,N_9882);
or UO_683 (O_683,N_9564,N_9866);
or UO_684 (O_684,N_9534,N_9802);
or UO_685 (O_685,N_9528,N_9828);
nand UO_686 (O_686,N_9799,N_9715);
nor UO_687 (O_687,N_9586,N_9990);
nand UO_688 (O_688,N_9873,N_9758);
nor UO_689 (O_689,N_9699,N_9559);
and UO_690 (O_690,N_9588,N_9565);
and UO_691 (O_691,N_9971,N_9808);
and UO_692 (O_692,N_9938,N_9736);
nor UO_693 (O_693,N_9931,N_9817);
and UO_694 (O_694,N_9556,N_9662);
and UO_695 (O_695,N_9616,N_9512);
and UO_696 (O_696,N_9880,N_9529);
nand UO_697 (O_697,N_9934,N_9817);
and UO_698 (O_698,N_9594,N_9960);
nand UO_699 (O_699,N_9847,N_9873);
nor UO_700 (O_700,N_9557,N_9703);
or UO_701 (O_701,N_9555,N_9759);
and UO_702 (O_702,N_9973,N_9514);
nor UO_703 (O_703,N_9526,N_9603);
nor UO_704 (O_704,N_9846,N_9763);
nand UO_705 (O_705,N_9647,N_9761);
or UO_706 (O_706,N_9912,N_9911);
or UO_707 (O_707,N_9965,N_9946);
or UO_708 (O_708,N_9831,N_9657);
xnor UO_709 (O_709,N_9844,N_9746);
or UO_710 (O_710,N_9929,N_9952);
and UO_711 (O_711,N_9558,N_9688);
and UO_712 (O_712,N_9601,N_9802);
or UO_713 (O_713,N_9852,N_9769);
and UO_714 (O_714,N_9677,N_9906);
nor UO_715 (O_715,N_9789,N_9908);
nand UO_716 (O_716,N_9681,N_9763);
or UO_717 (O_717,N_9653,N_9578);
or UO_718 (O_718,N_9852,N_9551);
and UO_719 (O_719,N_9553,N_9794);
and UO_720 (O_720,N_9593,N_9727);
nor UO_721 (O_721,N_9950,N_9528);
nor UO_722 (O_722,N_9700,N_9606);
nand UO_723 (O_723,N_9540,N_9846);
nor UO_724 (O_724,N_9732,N_9843);
or UO_725 (O_725,N_9699,N_9771);
nand UO_726 (O_726,N_9985,N_9556);
and UO_727 (O_727,N_9859,N_9536);
nor UO_728 (O_728,N_9673,N_9527);
and UO_729 (O_729,N_9719,N_9968);
or UO_730 (O_730,N_9985,N_9750);
or UO_731 (O_731,N_9880,N_9802);
and UO_732 (O_732,N_9574,N_9807);
and UO_733 (O_733,N_9523,N_9916);
and UO_734 (O_734,N_9806,N_9596);
and UO_735 (O_735,N_9651,N_9614);
and UO_736 (O_736,N_9627,N_9728);
and UO_737 (O_737,N_9720,N_9911);
nor UO_738 (O_738,N_9612,N_9981);
nor UO_739 (O_739,N_9741,N_9881);
or UO_740 (O_740,N_9950,N_9731);
or UO_741 (O_741,N_9663,N_9855);
nand UO_742 (O_742,N_9574,N_9756);
nor UO_743 (O_743,N_9544,N_9954);
and UO_744 (O_744,N_9771,N_9628);
or UO_745 (O_745,N_9716,N_9888);
or UO_746 (O_746,N_9518,N_9967);
nor UO_747 (O_747,N_9733,N_9792);
and UO_748 (O_748,N_9790,N_9807);
nor UO_749 (O_749,N_9743,N_9724);
or UO_750 (O_750,N_9657,N_9842);
or UO_751 (O_751,N_9870,N_9826);
and UO_752 (O_752,N_9941,N_9629);
nor UO_753 (O_753,N_9738,N_9731);
or UO_754 (O_754,N_9937,N_9788);
nand UO_755 (O_755,N_9863,N_9619);
nand UO_756 (O_756,N_9691,N_9656);
nand UO_757 (O_757,N_9927,N_9980);
or UO_758 (O_758,N_9573,N_9796);
nand UO_759 (O_759,N_9913,N_9730);
nor UO_760 (O_760,N_9679,N_9557);
nand UO_761 (O_761,N_9948,N_9845);
nor UO_762 (O_762,N_9928,N_9778);
nor UO_763 (O_763,N_9685,N_9982);
nor UO_764 (O_764,N_9833,N_9651);
nor UO_765 (O_765,N_9730,N_9623);
or UO_766 (O_766,N_9935,N_9607);
xor UO_767 (O_767,N_9547,N_9685);
or UO_768 (O_768,N_9623,N_9674);
nor UO_769 (O_769,N_9815,N_9658);
and UO_770 (O_770,N_9957,N_9711);
nand UO_771 (O_771,N_9789,N_9701);
nand UO_772 (O_772,N_9609,N_9866);
or UO_773 (O_773,N_9766,N_9594);
and UO_774 (O_774,N_9885,N_9554);
nand UO_775 (O_775,N_9716,N_9692);
and UO_776 (O_776,N_9710,N_9960);
or UO_777 (O_777,N_9691,N_9852);
nand UO_778 (O_778,N_9742,N_9615);
or UO_779 (O_779,N_9758,N_9978);
nand UO_780 (O_780,N_9720,N_9546);
and UO_781 (O_781,N_9921,N_9529);
or UO_782 (O_782,N_9834,N_9598);
nor UO_783 (O_783,N_9977,N_9713);
and UO_784 (O_784,N_9593,N_9831);
and UO_785 (O_785,N_9998,N_9956);
nor UO_786 (O_786,N_9703,N_9709);
and UO_787 (O_787,N_9852,N_9709);
or UO_788 (O_788,N_9878,N_9828);
or UO_789 (O_789,N_9722,N_9688);
nor UO_790 (O_790,N_9544,N_9578);
or UO_791 (O_791,N_9515,N_9830);
nand UO_792 (O_792,N_9874,N_9548);
and UO_793 (O_793,N_9758,N_9520);
nor UO_794 (O_794,N_9616,N_9910);
and UO_795 (O_795,N_9991,N_9921);
and UO_796 (O_796,N_9515,N_9595);
and UO_797 (O_797,N_9801,N_9851);
nand UO_798 (O_798,N_9776,N_9674);
and UO_799 (O_799,N_9865,N_9871);
or UO_800 (O_800,N_9992,N_9826);
and UO_801 (O_801,N_9608,N_9675);
or UO_802 (O_802,N_9887,N_9953);
or UO_803 (O_803,N_9813,N_9526);
or UO_804 (O_804,N_9506,N_9928);
nor UO_805 (O_805,N_9766,N_9597);
xnor UO_806 (O_806,N_9899,N_9855);
or UO_807 (O_807,N_9661,N_9962);
nor UO_808 (O_808,N_9568,N_9704);
nor UO_809 (O_809,N_9881,N_9792);
nand UO_810 (O_810,N_9896,N_9908);
nor UO_811 (O_811,N_9510,N_9852);
nor UO_812 (O_812,N_9607,N_9611);
nor UO_813 (O_813,N_9582,N_9533);
and UO_814 (O_814,N_9806,N_9773);
and UO_815 (O_815,N_9554,N_9840);
nand UO_816 (O_816,N_9834,N_9953);
nor UO_817 (O_817,N_9848,N_9861);
and UO_818 (O_818,N_9768,N_9900);
or UO_819 (O_819,N_9541,N_9870);
nand UO_820 (O_820,N_9867,N_9580);
nand UO_821 (O_821,N_9583,N_9987);
and UO_822 (O_822,N_9899,N_9814);
nor UO_823 (O_823,N_9734,N_9784);
or UO_824 (O_824,N_9650,N_9618);
or UO_825 (O_825,N_9645,N_9602);
or UO_826 (O_826,N_9865,N_9538);
nor UO_827 (O_827,N_9983,N_9735);
and UO_828 (O_828,N_9942,N_9788);
and UO_829 (O_829,N_9734,N_9852);
nand UO_830 (O_830,N_9835,N_9975);
nor UO_831 (O_831,N_9738,N_9872);
nor UO_832 (O_832,N_9586,N_9723);
nor UO_833 (O_833,N_9644,N_9854);
and UO_834 (O_834,N_9701,N_9620);
or UO_835 (O_835,N_9740,N_9696);
xnor UO_836 (O_836,N_9522,N_9748);
nor UO_837 (O_837,N_9681,N_9507);
or UO_838 (O_838,N_9913,N_9505);
and UO_839 (O_839,N_9856,N_9811);
or UO_840 (O_840,N_9762,N_9685);
or UO_841 (O_841,N_9599,N_9939);
and UO_842 (O_842,N_9516,N_9875);
and UO_843 (O_843,N_9786,N_9750);
nor UO_844 (O_844,N_9706,N_9847);
nor UO_845 (O_845,N_9679,N_9612);
nand UO_846 (O_846,N_9553,N_9524);
nor UO_847 (O_847,N_9608,N_9695);
nand UO_848 (O_848,N_9955,N_9605);
nand UO_849 (O_849,N_9848,N_9705);
nand UO_850 (O_850,N_9523,N_9843);
or UO_851 (O_851,N_9951,N_9952);
and UO_852 (O_852,N_9772,N_9500);
or UO_853 (O_853,N_9801,N_9788);
nand UO_854 (O_854,N_9814,N_9959);
or UO_855 (O_855,N_9529,N_9526);
nor UO_856 (O_856,N_9866,N_9943);
or UO_857 (O_857,N_9907,N_9842);
nand UO_858 (O_858,N_9789,N_9973);
nand UO_859 (O_859,N_9615,N_9760);
and UO_860 (O_860,N_9769,N_9780);
and UO_861 (O_861,N_9673,N_9511);
xnor UO_862 (O_862,N_9888,N_9865);
or UO_863 (O_863,N_9807,N_9838);
nand UO_864 (O_864,N_9992,N_9716);
and UO_865 (O_865,N_9900,N_9725);
nor UO_866 (O_866,N_9710,N_9990);
nand UO_867 (O_867,N_9985,N_9838);
nand UO_868 (O_868,N_9619,N_9937);
and UO_869 (O_869,N_9590,N_9971);
nor UO_870 (O_870,N_9506,N_9902);
or UO_871 (O_871,N_9915,N_9821);
nor UO_872 (O_872,N_9909,N_9989);
nand UO_873 (O_873,N_9669,N_9776);
and UO_874 (O_874,N_9806,N_9682);
or UO_875 (O_875,N_9609,N_9814);
and UO_876 (O_876,N_9712,N_9739);
nor UO_877 (O_877,N_9735,N_9984);
nor UO_878 (O_878,N_9781,N_9887);
and UO_879 (O_879,N_9934,N_9907);
nand UO_880 (O_880,N_9849,N_9643);
and UO_881 (O_881,N_9801,N_9511);
and UO_882 (O_882,N_9975,N_9588);
nand UO_883 (O_883,N_9674,N_9863);
nand UO_884 (O_884,N_9947,N_9694);
or UO_885 (O_885,N_9674,N_9745);
and UO_886 (O_886,N_9625,N_9789);
nor UO_887 (O_887,N_9736,N_9641);
nand UO_888 (O_888,N_9700,N_9666);
nand UO_889 (O_889,N_9764,N_9739);
and UO_890 (O_890,N_9990,N_9941);
nor UO_891 (O_891,N_9537,N_9638);
nor UO_892 (O_892,N_9807,N_9610);
xnor UO_893 (O_893,N_9677,N_9728);
and UO_894 (O_894,N_9780,N_9638);
nand UO_895 (O_895,N_9721,N_9515);
nor UO_896 (O_896,N_9920,N_9934);
or UO_897 (O_897,N_9949,N_9858);
and UO_898 (O_898,N_9988,N_9817);
nand UO_899 (O_899,N_9673,N_9784);
nand UO_900 (O_900,N_9643,N_9940);
nand UO_901 (O_901,N_9666,N_9582);
xnor UO_902 (O_902,N_9798,N_9844);
and UO_903 (O_903,N_9927,N_9898);
nand UO_904 (O_904,N_9737,N_9640);
or UO_905 (O_905,N_9969,N_9548);
nand UO_906 (O_906,N_9686,N_9557);
or UO_907 (O_907,N_9660,N_9873);
and UO_908 (O_908,N_9860,N_9553);
nand UO_909 (O_909,N_9572,N_9916);
nand UO_910 (O_910,N_9543,N_9566);
or UO_911 (O_911,N_9627,N_9678);
and UO_912 (O_912,N_9805,N_9840);
and UO_913 (O_913,N_9852,N_9948);
or UO_914 (O_914,N_9896,N_9888);
or UO_915 (O_915,N_9710,N_9755);
nor UO_916 (O_916,N_9947,N_9841);
or UO_917 (O_917,N_9629,N_9830);
xor UO_918 (O_918,N_9890,N_9794);
nand UO_919 (O_919,N_9589,N_9723);
nor UO_920 (O_920,N_9575,N_9861);
nor UO_921 (O_921,N_9815,N_9707);
nand UO_922 (O_922,N_9984,N_9905);
nor UO_923 (O_923,N_9614,N_9755);
nor UO_924 (O_924,N_9962,N_9561);
nand UO_925 (O_925,N_9654,N_9935);
nor UO_926 (O_926,N_9681,N_9630);
nand UO_927 (O_927,N_9921,N_9986);
nor UO_928 (O_928,N_9844,N_9936);
nor UO_929 (O_929,N_9844,N_9921);
and UO_930 (O_930,N_9965,N_9771);
nor UO_931 (O_931,N_9621,N_9934);
nor UO_932 (O_932,N_9976,N_9679);
nor UO_933 (O_933,N_9616,N_9990);
or UO_934 (O_934,N_9645,N_9978);
nor UO_935 (O_935,N_9853,N_9599);
nand UO_936 (O_936,N_9819,N_9849);
and UO_937 (O_937,N_9672,N_9604);
and UO_938 (O_938,N_9599,N_9945);
and UO_939 (O_939,N_9960,N_9608);
nor UO_940 (O_940,N_9649,N_9953);
and UO_941 (O_941,N_9734,N_9788);
or UO_942 (O_942,N_9731,N_9713);
nand UO_943 (O_943,N_9581,N_9521);
nor UO_944 (O_944,N_9530,N_9631);
or UO_945 (O_945,N_9605,N_9763);
nor UO_946 (O_946,N_9644,N_9873);
nand UO_947 (O_947,N_9794,N_9725);
and UO_948 (O_948,N_9945,N_9581);
nand UO_949 (O_949,N_9847,N_9880);
nand UO_950 (O_950,N_9882,N_9582);
and UO_951 (O_951,N_9508,N_9654);
nand UO_952 (O_952,N_9796,N_9770);
or UO_953 (O_953,N_9714,N_9772);
or UO_954 (O_954,N_9838,N_9885);
and UO_955 (O_955,N_9943,N_9531);
xor UO_956 (O_956,N_9534,N_9735);
or UO_957 (O_957,N_9682,N_9645);
and UO_958 (O_958,N_9521,N_9781);
or UO_959 (O_959,N_9927,N_9574);
nand UO_960 (O_960,N_9562,N_9619);
nand UO_961 (O_961,N_9736,N_9912);
and UO_962 (O_962,N_9866,N_9717);
nand UO_963 (O_963,N_9572,N_9826);
and UO_964 (O_964,N_9745,N_9544);
or UO_965 (O_965,N_9828,N_9555);
and UO_966 (O_966,N_9823,N_9623);
nor UO_967 (O_967,N_9940,N_9639);
or UO_968 (O_968,N_9532,N_9790);
nor UO_969 (O_969,N_9940,N_9909);
nand UO_970 (O_970,N_9518,N_9870);
and UO_971 (O_971,N_9600,N_9609);
or UO_972 (O_972,N_9791,N_9969);
nand UO_973 (O_973,N_9596,N_9762);
or UO_974 (O_974,N_9521,N_9576);
or UO_975 (O_975,N_9567,N_9724);
nor UO_976 (O_976,N_9705,N_9973);
or UO_977 (O_977,N_9756,N_9818);
nand UO_978 (O_978,N_9977,N_9708);
or UO_979 (O_979,N_9697,N_9965);
xnor UO_980 (O_980,N_9591,N_9540);
nor UO_981 (O_981,N_9578,N_9605);
nor UO_982 (O_982,N_9660,N_9886);
and UO_983 (O_983,N_9643,N_9783);
nand UO_984 (O_984,N_9783,N_9969);
or UO_985 (O_985,N_9990,N_9644);
nand UO_986 (O_986,N_9681,N_9922);
and UO_987 (O_987,N_9709,N_9547);
and UO_988 (O_988,N_9885,N_9973);
and UO_989 (O_989,N_9929,N_9774);
or UO_990 (O_990,N_9918,N_9598);
nor UO_991 (O_991,N_9595,N_9831);
nand UO_992 (O_992,N_9936,N_9957);
and UO_993 (O_993,N_9601,N_9862);
nor UO_994 (O_994,N_9545,N_9539);
nor UO_995 (O_995,N_9753,N_9504);
and UO_996 (O_996,N_9917,N_9784);
and UO_997 (O_997,N_9604,N_9967);
and UO_998 (O_998,N_9948,N_9569);
nor UO_999 (O_999,N_9989,N_9540);
and UO_1000 (O_1000,N_9514,N_9888);
or UO_1001 (O_1001,N_9837,N_9955);
nand UO_1002 (O_1002,N_9866,N_9730);
nand UO_1003 (O_1003,N_9587,N_9645);
and UO_1004 (O_1004,N_9654,N_9618);
nand UO_1005 (O_1005,N_9717,N_9777);
or UO_1006 (O_1006,N_9759,N_9742);
and UO_1007 (O_1007,N_9524,N_9948);
nor UO_1008 (O_1008,N_9596,N_9957);
nor UO_1009 (O_1009,N_9692,N_9768);
nor UO_1010 (O_1010,N_9781,N_9953);
nor UO_1011 (O_1011,N_9721,N_9551);
or UO_1012 (O_1012,N_9760,N_9810);
nor UO_1013 (O_1013,N_9523,N_9942);
nand UO_1014 (O_1014,N_9609,N_9884);
nand UO_1015 (O_1015,N_9903,N_9574);
nor UO_1016 (O_1016,N_9766,N_9745);
xor UO_1017 (O_1017,N_9658,N_9893);
nand UO_1018 (O_1018,N_9917,N_9849);
and UO_1019 (O_1019,N_9742,N_9798);
nand UO_1020 (O_1020,N_9517,N_9904);
nand UO_1021 (O_1021,N_9805,N_9776);
nand UO_1022 (O_1022,N_9784,N_9665);
or UO_1023 (O_1023,N_9868,N_9941);
or UO_1024 (O_1024,N_9744,N_9976);
nor UO_1025 (O_1025,N_9823,N_9654);
nand UO_1026 (O_1026,N_9960,N_9787);
xnor UO_1027 (O_1027,N_9781,N_9881);
nor UO_1028 (O_1028,N_9926,N_9708);
nand UO_1029 (O_1029,N_9927,N_9509);
xnor UO_1030 (O_1030,N_9849,N_9971);
nand UO_1031 (O_1031,N_9993,N_9934);
nand UO_1032 (O_1032,N_9951,N_9584);
nor UO_1033 (O_1033,N_9629,N_9617);
nand UO_1034 (O_1034,N_9888,N_9536);
nor UO_1035 (O_1035,N_9514,N_9872);
and UO_1036 (O_1036,N_9565,N_9920);
and UO_1037 (O_1037,N_9591,N_9731);
nand UO_1038 (O_1038,N_9786,N_9627);
nand UO_1039 (O_1039,N_9862,N_9840);
nor UO_1040 (O_1040,N_9831,N_9822);
or UO_1041 (O_1041,N_9900,N_9514);
nand UO_1042 (O_1042,N_9914,N_9972);
nand UO_1043 (O_1043,N_9608,N_9873);
or UO_1044 (O_1044,N_9828,N_9570);
and UO_1045 (O_1045,N_9759,N_9624);
and UO_1046 (O_1046,N_9860,N_9800);
nor UO_1047 (O_1047,N_9869,N_9723);
nor UO_1048 (O_1048,N_9801,N_9691);
or UO_1049 (O_1049,N_9655,N_9592);
and UO_1050 (O_1050,N_9553,N_9791);
and UO_1051 (O_1051,N_9567,N_9796);
or UO_1052 (O_1052,N_9837,N_9924);
and UO_1053 (O_1053,N_9559,N_9795);
or UO_1054 (O_1054,N_9835,N_9797);
nor UO_1055 (O_1055,N_9954,N_9994);
and UO_1056 (O_1056,N_9792,N_9750);
or UO_1057 (O_1057,N_9673,N_9632);
nor UO_1058 (O_1058,N_9667,N_9607);
xor UO_1059 (O_1059,N_9979,N_9965);
nor UO_1060 (O_1060,N_9646,N_9578);
nand UO_1061 (O_1061,N_9857,N_9837);
nor UO_1062 (O_1062,N_9748,N_9867);
nand UO_1063 (O_1063,N_9649,N_9947);
nand UO_1064 (O_1064,N_9786,N_9893);
nor UO_1065 (O_1065,N_9635,N_9761);
nor UO_1066 (O_1066,N_9636,N_9586);
nor UO_1067 (O_1067,N_9800,N_9949);
and UO_1068 (O_1068,N_9958,N_9770);
nand UO_1069 (O_1069,N_9649,N_9825);
or UO_1070 (O_1070,N_9781,N_9902);
xor UO_1071 (O_1071,N_9713,N_9829);
and UO_1072 (O_1072,N_9937,N_9835);
or UO_1073 (O_1073,N_9739,N_9896);
nand UO_1074 (O_1074,N_9585,N_9527);
nand UO_1075 (O_1075,N_9716,N_9928);
and UO_1076 (O_1076,N_9774,N_9807);
and UO_1077 (O_1077,N_9834,N_9676);
or UO_1078 (O_1078,N_9835,N_9795);
nand UO_1079 (O_1079,N_9804,N_9920);
and UO_1080 (O_1080,N_9553,N_9619);
or UO_1081 (O_1081,N_9811,N_9840);
or UO_1082 (O_1082,N_9760,N_9764);
and UO_1083 (O_1083,N_9927,N_9833);
nor UO_1084 (O_1084,N_9829,N_9626);
xnor UO_1085 (O_1085,N_9999,N_9960);
nor UO_1086 (O_1086,N_9753,N_9933);
and UO_1087 (O_1087,N_9550,N_9857);
or UO_1088 (O_1088,N_9801,N_9714);
nor UO_1089 (O_1089,N_9648,N_9889);
and UO_1090 (O_1090,N_9517,N_9970);
and UO_1091 (O_1091,N_9826,N_9528);
nor UO_1092 (O_1092,N_9648,N_9744);
or UO_1093 (O_1093,N_9633,N_9963);
nor UO_1094 (O_1094,N_9831,N_9875);
nand UO_1095 (O_1095,N_9522,N_9831);
nor UO_1096 (O_1096,N_9955,N_9813);
and UO_1097 (O_1097,N_9980,N_9516);
nor UO_1098 (O_1098,N_9825,N_9779);
nor UO_1099 (O_1099,N_9594,N_9776);
nand UO_1100 (O_1100,N_9996,N_9686);
or UO_1101 (O_1101,N_9788,N_9918);
nor UO_1102 (O_1102,N_9583,N_9871);
and UO_1103 (O_1103,N_9608,N_9563);
or UO_1104 (O_1104,N_9838,N_9538);
nor UO_1105 (O_1105,N_9632,N_9781);
or UO_1106 (O_1106,N_9902,N_9663);
or UO_1107 (O_1107,N_9576,N_9651);
nor UO_1108 (O_1108,N_9550,N_9571);
nand UO_1109 (O_1109,N_9551,N_9606);
nor UO_1110 (O_1110,N_9752,N_9678);
nor UO_1111 (O_1111,N_9668,N_9818);
nand UO_1112 (O_1112,N_9834,N_9916);
xnor UO_1113 (O_1113,N_9949,N_9986);
nor UO_1114 (O_1114,N_9504,N_9996);
and UO_1115 (O_1115,N_9589,N_9759);
xor UO_1116 (O_1116,N_9601,N_9690);
and UO_1117 (O_1117,N_9583,N_9948);
or UO_1118 (O_1118,N_9573,N_9881);
xnor UO_1119 (O_1119,N_9854,N_9957);
or UO_1120 (O_1120,N_9869,N_9792);
nand UO_1121 (O_1121,N_9757,N_9977);
nand UO_1122 (O_1122,N_9673,N_9517);
nor UO_1123 (O_1123,N_9610,N_9522);
nor UO_1124 (O_1124,N_9728,N_9506);
nor UO_1125 (O_1125,N_9938,N_9901);
and UO_1126 (O_1126,N_9606,N_9980);
nand UO_1127 (O_1127,N_9883,N_9907);
and UO_1128 (O_1128,N_9993,N_9665);
or UO_1129 (O_1129,N_9519,N_9537);
and UO_1130 (O_1130,N_9687,N_9548);
nand UO_1131 (O_1131,N_9644,N_9799);
nand UO_1132 (O_1132,N_9895,N_9913);
or UO_1133 (O_1133,N_9719,N_9735);
or UO_1134 (O_1134,N_9506,N_9628);
and UO_1135 (O_1135,N_9707,N_9768);
or UO_1136 (O_1136,N_9829,N_9724);
nor UO_1137 (O_1137,N_9878,N_9729);
and UO_1138 (O_1138,N_9812,N_9590);
and UO_1139 (O_1139,N_9671,N_9984);
or UO_1140 (O_1140,N_9923,N_9533);
nor UO_1141 (O_1141,N_9542,N_9668);
nand UO_1142 (O_1142,N_9653,N_9908);
or UO_1143 (O_1143,N_9528,N_9946);
or UO_1144 (O_1144,N_9787,N_9598);
nand UO_1145 (O_1145,N_9564,N_9931);
nand UO_1146 (O_1146,N_9744,N_9559);
nand UO_1147 (O_1147,N_9809,N_9747);
or UO_1148 (O_1148,N_9814,N_9842);
and UO_1149 (O_1149,N_9860,N_9903);
and UO_1150 (O_1150,N_9758,N_9633);
or UO_1151 (O_1151,N_9992,N_9857);
or UO_1152 (O_1152,N_9819,N_9787);
xor UO_1153 (O_1153,N_9915,N_9981);
nand UO_1154 (O_1154,N_9695,N_9713);
nand UO_1155 (O_1155,N_9563,N_9924);
nand UO_1156 (O_1156,N_9698,N_9623);
nor UO_1157 (O_1157,N_9698,N_9505);
and UO_1158 (O_1158,N_9725,N_9878);
nand UO_1159 (O_1159,N_9723,N_9742);
nand UO_1160 (O_1160,N_9840,N_9860);
or UO_1161 (O_1161,N_9571,N_9861);
nor UO_1162 (O_1162,N_9936,N_9551);
nand UO_1163 (O_1163,N_9785,N_9898);
nand UO_1164 (O_1164,N_9538,N_9810);
or UO_1165 (O_1165,N_9690,N_9560);
nor UO_1166 (O_1166,N_9511,N_9520);
nor UO_1167 (O_1167,N_9636,N_9621);
or UO_1168 (O_1168,N_9780,N_9789);
and UO_1169 (O_1169,N_9913,N_9737);
nand UO_1170 (O_1170,N_9990,N_9798);
or UO_1171 (O_1171,N_9730,N_9922);
xor UO_1172 (O_1172,N_9896,N_9925);
nor UO_1173 (O_1173,N_9801,N_9674);
nand UO_1174 (O_1174,N_9673,N_9840);
nand UO_1175 (O_1175,N_9548,N_9965);
or UO_1176 (O_1176,N_9680,N_9787);
or UO_1177 (O_1177,N_9616,N_9939);
or UO_1178 (O_1178,N_9789,N_9603);
and UO_1179 (O_1179,N_9750,N_9511);
and UO_1180 (O_1180,N_9740,N_9956);
nand UO_1181 (O_1181,N_9841,N_9515);
and UO_1182 (O_1182,N_9605,N_9677);
or UO_1183 (O_1183,N_9749,N_9580);
nand UO_1184 (O_1184,N_9929,N_9907);
or UO_1185 (O_1185,N_9894,N_9595);
nor UO_1186 (O_1186,N_9516,N_9660);
nand UO_1187 (O_1187,N_9803,N_9697);
nand UO_1188 (O_1188,N_9735,N_9810);
or UO_1189 (O_1189,N_9944,N_9610);
nand UO_1190 (O_1190,N_9957,N_9525);
or UO_1191 (O_1191,N_9559,N_9642);
or UO_1192 (O_1192,N_9663,N_9815);
and UO_1193 (O_1193,N_9785,N_9870);
nand UO_1194 (O_1194,N_9885,N_9813);
nor UO_1195 (O_1195,N_9852,N_9689);
xor UO_1196 (O_1196,N_9736,N_9769);
nor UO_1197 (O_1197,N_9667,N_9995);
or UO_1198 (O_1198,N_9525,N_9629);
nor UO_1199 (O_1199,N_9717,N_9903);
xnor UO_1200 (O_1200,N_9811,N_9744);
or UO_1201 (O_1201,N_9718,N_9684);
and UO_1202 (O_1202,N_9901,N_9627);
nand UO_1203 (O_1203,N_9575,N_9752);
nor UO_1204 (O_1204,N_9518,N_9525);
or UO_1205 (O_1205,N_9564,N_9561);
or UO_1206 (O_1206,N_9797,N_9961);
nor UO_1207 (O_1207,N_9979,N_9703);
nand UO_1208 (O_1208,N_9714,N_9814);
and UO_1209 (O_1209,N_9943,N_9646);
nand UO_1210 (O_1210,N_9831,N_9654);
and UO_1211 (O_1211,N_9949,N_9721);
nor UO_1212 (O_1212,N_9838,N_9650);
nor UO_1213 (O_1213,N_9598,N_9944);
or UO_1214 (O_1214,N_9909,N_9552);
nor UO_1215 (O_1215,N_9735,N_9568);
nand UO_1216 (O_1216,N_9760,N_9511);
or UO_1217 (O_1217,N_9608,N_9594);
nand UO_1218 (O_1218,N_9574,N_9768);
xnor UO_1219 (O_1219,N_9878,N_9869);
and UO_1220 (O_1220,N_9851,N_9513);
or UO_1221 (O_1221,N_9799,N_9798);
or UO_1222 (O_1222,N_9931,N_9844);
nor UO_1223 (O_1223,N_9948,N_9673);
or UO_1224 (O_1224,N_9985,N_9972);
nor UO_1225 (O_1225,N_9961,N_9580);
nor UO_1226 (O_1226,N_9651,N_9645);
nand UO_1227 (O_1227,N_9653,N_9520);
and UO_1228 (O_1228,N_9756,N_9645);
nand UO_1229 (O_1229,N_9501,N_9777);
or UO_1230 (O_1230,N_9685,N_9651);
nor UO_1231 (O_1231,N_9922,N_9666);
and UO_1232 (O_1232,N_9775,N_9715);
and UO_1233 (O_1233,N_9856,N_9774);
nand UO_1234 (O_1234,N_9607,N_9512);
nor UO_1235 (O_1235,N_9921,N_9860);
or UO_1236 (O_1236,N_9595,N_9949);
nor UO_1237 (O_1237,N_9601,N_9873);
or UO_1238 (O_1238,N_9821,N_9643);
nand UO_1239 (O_1239,N_9964,N_9661);
xnor UO_1240 (O_1240,N_9654,N_9703);
nand UO_1241 (O_1241,N_9998,N_9733);
nand UO_1242 (O_1242,N_9977,N_9573);
nand UO_1243 (O_1243,N_9620,N_9513);
or UO_1244 (O_1244,N_9555,N_9575);
nand UO_1245 (O_1245,N_9810,N_9949);
and UO_1246 (O_1246,N_9639,N_9568);
nor UO_1247 (O_1247,N_9897,N_9986);
nand UO_1248 (O_1248,N_9829,N_9894);
nand UO_1249 (O_1249,N_9762,N_9860);
xor UO_1250 (O_1250,N_9763,N_9771);
and UO_1251 (O_1251,N_9911,N_9843);
nand UO_1252 (O_1252,N_9832,N_9784);
nand UO_1253 (O_1253,N_9711,N_9717);
and UO_1254 (O_1254,N_9507,N_9981);
nand UO_1255 (O_1255,N_9865,N_9635);
nand UO_1256 (O_1256,N_9829,N_9522);
nand UO_1257 (O_1257,N_9531,N_9780);
or UO_1258 (O_1258,N_9647,N_9554);
and UO_1259 (O_1259,N_9527,N_9784);
nor UO_1260 (O_1260,N_9522,N_9895);
or UO_1261 (O_1261,N_9855,N_9784);
or UO_1262 (O_1262,N_9942,N_9927);
nand UO_1263 (O_1263,N_9591,N_9585);
and UO_1264 (O_1264,N_9928,N_9641);
or UO_1265 (O_1265,N_9739,N_9904);
nor UO_1266 (O_1266,N_9854,N_9864);
nor UO_1267 (O_1267,N_9515,N_9961);
nor UO_1268 (O_1268,N_9546,N_9574);
and UO_1269 (O_1269,N_9757,N_9719);
and UO_1270 (O_1270,N_9961,N_9872);
and UO_1271 (O_1271,N_9718,N_9594);
xnor UO_1272 (O_1272,N_9955,N_9601);
and UO_1273 (O_1273,N_9932,N_9517);
nand UO_1274 (O_1274,N_9643,N_9707);
nand UO_1275 (O_1275,N_9898,N_9728);
nor UO_1276 (O_1276,N_9784,N_9848);
nand UO_1277 (O_1277,N_9688,N_9852);
and UO_1278 (O_1278,N_9878,N_9925);
or UO_1279 (O_1279,N_9783,N_9504);
nor UO_1280 (O_1280,N_9738,N_9945);
and UO_1281 (O_1281,N_9760,N_9549);
nor UO_1282 (O_1282,N_9904,N_9843);
nand UO_1283 (O_1283,N_9811,N_9927);
and UO_1284 (O_1284,N_9783,N_9930);
and UO_1285 (O_1285,N_9636,N_9913);
nand UO_1286 (O_1286,N_9650,N_9830);
xor UO_1287 (O_1287,N_9543,N_9756);
and UO_1288 (O_1288,N_9937,N_9585);
nor UO_1289 (O_1289,N_9968,N_9570);
nor UO_1290 (O_1290,N_9889,N_9731);
nand UO_1291 (O_1291,N_9727,N_9550);
nor UO_1292 (O_1292,N_9771,N_9650);
or UO_1293 (O_1293,N_9526,N_9957);
nand UO_1294 (O_1294,N_9726,N_9793);
and UO_1295 (O_1295,N_9940,N_9769);
nor UO_1296 (O_1296,N_9816,N_9787);
xnor UO_1297 (O_1297,N_9610,N_9574);
nand UO_1298 (O_1298,N_9521,N_9897);
nor UO_1299 (O_1299,N_9586,N_9760);
nand UO_1300 (O_1300,N_9631,N_9873);
and UO_1301 (O_1301,N_9517,N_9500);
and UO_1302 (O_1302,N_9747,N_9737);
nand UO_1303 (O_1303,N_9551,N_9773);
nor UO_1304 (O_1304,N_9683,N_9713);
or UO_1305 (O_1305,N_9835,N_9692);
nor UO_1306 (O_1306,N_9820,N_9983);
or UO_1307 (O_1307,N_9782,N_9991);
nand UO_1308 (O_1308,N_9525,N_9536);
nand UO_1309 (O_1309,N_9762,N_9739);
and UO_1310 (O_1310,N_9674,N_9978);
nand UO_1311 (O_1311,N_9534,N_9840);
and UO_1312 (O_1312,N_9827,N_9974);
xor UO_1313 (O_1313,N_9715,N_9647);
nand UO_1314 (O_1314,N_9522,N_9742);
nor UO_1315 (O_1315,N_9865,N_9972);
and UO_1316 (O_1316,N_9873,N_9655);
and UO_1317 (O_1317,N_9630,N_9935);
and UO_1318 (O_1318,N_9527,N_9814);
nor UO_1319 (O_1319,N_9598,N_9661);
and UO_1320 (O_1320,N_9603,N_9791);
and UO_1321 (O_1321,N_9722,N_9849);
nand UO_1322 (O_1322,N_9802,N_9740);
nand UO_1323 (O_1323,N_9964,N_9844);
nand UO_1324 (O_1324,N_9799,N_9573);
and UO_1325 (O_1325,N_9511,N_9898);
nor UO_1326 (O_1326,N_9556,N_9805);
and UO_1327 (O_1327,N_9946,N_9583);
or UO_1328 (O_1328,N_9602,N_9513);
or UO_1329 (O_1329,N_9737,N_9614);
or UO_1330 (O_1330,N_9738,N_9873);
and UO_1331 (O_1331,N_9799,N_9765);
nand UO_1332 (O_1332,N_9610,N_9779);
nand UO_1333 (O_1333,N_9678,N_9972);
and UO_1334 (O_1334,N_9856,N_9696);
xnor UO_1335 (O_1335,N_9768,N_9932);
or UO_1336 (O_1336,N_9695,N_9806);
and UO_1337 (O_1337,N_9570,N_9779);
nor UO_1338 (O_1338,N_9723,N_9883);
or UO_1339 (O_1339,N_9606,N_9995);
or UO_1340 (O_1340,N_9677,N_9568);
nor UO_1341 (O_1341,N_9818,N_9974);
and UO_1342 (O_1342,N_9829,N_9669);
or UO_1343 (O_1343,N_9844,N_9665);
nand UO_1344 (O_1344,N_9623,N_9513);
and UO_1345 (O_1345,N_9736,N_9760);
or UO_1346 (O_1346,N_9901,N_9721);
nand UO_1347 (O_1347,N_9802,N_9733);
nand UO_1348 (O_1348,N_9939,N_9833);
nand UO_1349 (O_1349,N_9845,N_9997);
nor UO_1350 (O_1350,N_9821,N_9720);
nand UO_1351 (O_1351,N_9784,N_9687);
and UO_1352 (O_1352,N_9925,N_9909);
nand UO_1353 (O_1353,N_9944,N_9696);
and UO_1354 (O_1354,N_9570,N_9607);
or UO_1355 (O_1355,N_9879,N_9601);
and UO_1356 (O_1356,N_9558,N_9965);
or UO_1357 (O_1357,N_9851,N_9823);
and UO_1358 (O_1358,N_9646,N_9655);
and UO_1359 (O_1359,N_9778,N_9639);
nand UO_1360 (O_1360,N_9586,N_9974);
or UO_1361 (O_1361,N_9544,N_9957);
nor UO_1362 (O_1362,N_9633,N_9618);
and UO_1363 (O_1363,N_9550,N_9713);
or UO_1364 (O_1364,N_9504,N_9902);
and UO_1365 (O_1365,N_9939,N_9855);
or UO_1366 (O_1366,N_9862,N_9568);
nor UO_1367 (O_1367,N_9845,N_9577);
nand UO_1368 (O_1368,N_9963,N_9747);
or UO_1369 (O_1369,N_9887,N_9929);
nand UO_1370 (O_1370,N_9992,N_9730);
or UO_1371 (O_1371,N_9616,N_9857);
or UO_1372 (O_1372,N_9862,N_9953);
nand UO_1373 (O_1373,N_9708,N_9960);
or UO_1374 (O_1374,N_9734,N_9546);
and UO_1375 (O_1375,N_9622,N_9873);
and UO_1376 (O_1376,N_9980,N_9679);
nor UO_1377 (O_1377,N_9509,N_9930);
nor UO_1378 (O_1378,N_9768,N_9723);
or UO_1379 (O_1379,N_9686,N_9676);
nand UO_1380 (O_1380,N_9765,N_9707);
and UO_1381 (O_1381,N_9878,N_9753);
or UO_1382 (O_1382,N_9966,N_9591);
nand UO_1383 (O_1383,N_9960,N_9641);
or UO_1384 (O_1384,N_9709,N_9751);
nand UO_1385 (O_1385,N_9767,N_9659);
or UO_1386 (O_1386,N_9515,N_9532);
and UO_1387 (O_1387,N_9944,N_9889);
or UO_1388 (O_1388,N_9861,N_9657);
and UO_1389 (O_1389,N_9813,N_9907);
nand UO_1390 (O_1390,N_9656,N_9630);
nor UO_1391 (O_1391,N_9915,N_9599);
nand UO_1392 (O_1392,N_9532,N_9978);
and UO_1393 (O_1393,N_9705,N_9712);
or UO_1394 (O_1394,N_9718,N_9977);
nand UO_1395 (O_1395,N_9785,N_9561);
and UO_1396 (O_1396,N_9971,N_9520);
nor UO_1397 (O_1397,N_9642,N_9752);
and UO_1398 (O_1398,N_9635,N_9672);
nand UO_1399 (O_1399,N_9569,N_9588);
or UO_1400 (O_1400,N_9975,N_9819);
and UO_1401 (O_1401,N_9771,N_9820);
nor UO_1402 (O_1402,N_9977,N_9937);
or UO_1403 (O_1403,N_9584,N_9677);
or UO_1404 (O_1404,N_9782,N_9567);
nor UO_1405 (O_1405,N_9542,N_9614);
and UO_1406 (O_1406,N_9800,N_9573);
nand UO_1407 (O_1407,N_9528,N_9780);
and UO_1408 (O_1408,N_9872,N_9681);
or UO_1409 (O_1409,N_9868,N_9893);
or UO_1410 (O_1410,N_9656,N_9759);
and UO_1411 (O_1411,N_9635,N_9642);
nand UO_1412 (O_1412,N_9535,N_9601);
and UO_1413 (O_1413,N_9678,N_9717);
and UO_1414 (O_1414,N_9999,N_9998);
nor UO_1415 (O_1415,N_9889,N_9839);
or UO_1416 (O_1416,N_9662,N_9828);
or UO_1417 (O_1417,N_9711,N_9579);
and UO_1418 (O_1418,N_9511,N_9632);
or UO_1419 (O_1419,N_9703,N_9692);
or UO_1420 (O_1420,N_9767,N_9784);
nand UO_1421 (O_1421,N_9528,N_9589);
or UO_1422 (O_1422,N_9787,N_9580);
nand UO_1423 (O_1423,N_9976,N_9592);
nand UO_1424 (O_1424,N_9772,N_9979);
or UO_1425 (O_1425,N_9939,N_9740);
nor UO_1426 (O_1426,N_9594,N_9717);
and UO_1427 (O_1427,N_9832,N_9807);
or UO_1428 (O_1428,N_9891,N_9552);
and UO_1429 (O_1429,N_9878,N_9981);
or UO_1430 (O_1430,N_9945,N_9697);
nand UO_1431 (O_1431,N_9943,N_9974);
nand UO_1432 (O_1432,N_9768,N_9795);
and UO_1433 (O_1433,N_9926,N_9815);
or UO_1434 (O_1434,N_9811,N_9960);
or UO_1435 (O_1435,N_9573,N_9648);
nand UO_1436 (O_1436,N_9912,N_9835);
and UO_1437 (O_1437,N_9584,N_9596);
and UO_1438 (O_1438,N_9699,N_9703);
nand UO_1439 (O_1439,N_9828,N_9906);
nor UO_1440 (O_1440,N_9766,N_9828);
or UO_1441 (O_1441,N_9941,N_9502);
or UO_1442 (O_1442,N_9889,N_9560);
or UO_1443 (O_1443,N_9755,N_9885);
or UO_1444 (O_1444,N_9609,N_9594);
nand UO_1445 (O_1445,N_9781,N_9543);
nor UO_1446 (O_1446,N_9579,N_9917);
and UO_1447 (O_1447,N_9630,N_9723);
nor UO_1448 (O_1448,N_9605,N_9701);
and UO_1449 (O_1449,N_9533,N_9774);
nand UO_1450 (O_1450,N_9646,N_9737);
or UO_1451 (O_1451,N_9886,N_9723);
nor UO_1452 (O_1452,N_9837,N_9897);
nor UO_1453 (O_1453,N_9735,N_9814);
nor UO_1454 (O_1454,N_9509,N_9882);
nor UO_1455 (O_1455,N_9822,N_9788);
or UO_1456 (O_1456,N_9702,N_9845);
nand UO_1457 (O_1457,N_9506,N_9957);
and UO_1458 (O_1458,N_9834,N_9579);
or UO_1459 (O_1459,N_9913,N_9583);
or UO_1460 (O_1460,N_9951,N_9832);
or UO_1461 (O_1461,N_9859,N_9588);
nor UO_1462 (O_1462,N_9615,N_9643);
nand UO_1463 (O_1463,N_9546,N_9595);
nor UO_1464 (O_1464,N_9504,N_9694);
or UO_1465 (O_1465,N_9719,N_9753);
nor UO_1466 (O_1466,N_9786,N_9785);
or UO_1467 (O_1467,N_9607,N_9510);
nor UO_1468 (O_1468,N_9626,N_9967);
nand UO_1469 (O_1469,N_9938,N_9829);
nor UO_1470 (O_1470,N_9818,N_9769);
or UO_1471 (O_1471,N_9667,N_9789);
and UO_1472 (O_1472,N_9734,N_9654);
nand UO_1473 (O_1473,N_9991,N_9688);
or UO_1474 (O_1474,N_9796,N_9808);
nor UO_1475 (O_1475,N_9946,N_9738);
and UO_1476 (O_1476,N_9629,N_9666);
xor UO_1477 (O_1477,N_9521,N_9697);
or UO_1478 (O_1478,N_9577,N_9602);
and UO_1479 (O_1479,N_9679,N_9654);
nand UO_1480 (O_1480,N_9570,N_9916);
nor UO_1481 (O_1481,N_9517,N_9681);
nor UO_1482 (O_1482,N_9881,N_9812);
nor UO_1483 (O_1483,N_9674,N_9796);
nor UO_1484 (O_1484,N_9826,N_9997);
or UO_1485 (O_1485,N_9546,N_9777);
and UO_1486 (O_1486,N_9590,N_9791);
or UO_1487 (O_1487,N_9603,N_9762);
or UO_1488 (O_1488,N_9625,N_9694);
nand UO_1489 (O_1489,N_9840,N_9920);
nor UO_1490 (O_1490,N_9630,N_9724);
nor UO_1491 (O_1491,N_9776,N_9673);
xor UO_1492 (O_1492,N_9545,N_9557);
nand UO_1493 (O_1493,N_9782,N_9554);
nand UO_1494 (O_1494,N_9947,N_9611);
nand UO_1495 (O_1495,N_9685,N_9928);
nor UO_1496 (O_1496,N_9535,N_9701);
and UO_1497 (O_1497,N_9781,N_9758);
nor UO_1498 (O_1498,N_9957,N_9972);
or UO_1499 (O_1499,N_9780,N_9516);
endmodule