module basic_5000_50000_5000_200_levels_10xor_2(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,In_3000,In_3001,In_3002,In_3003,In_3004,In_3005,In_3006,In_3007,In_3008,In_3009,In_3010,In_3011,In_3012,In_3013,In_3014,In_3015,In_3016,In_3017,In_3018,In_3019,In_3020,In_3021,In_3022,In_3023,In_3024,In_3025,In_3026,In_3027,In_3028,In_3029,In_3030,In_3031,In_3032,In_3033,In_3034,In_3035,In_3036,In_3037,In_3038,In_3039,In_3040,In_3041,In_3042,In_3043,In_3044,In_3045,In_3046,In_3047,In_3048,In_3049,In_3050,In_3051,In_3052,In_3053,In_3054,In_3055,In_3056,In_3057,In_3058,In_3059,In_3060,In_3061,In_3062,In_3063,In_3064,In_3065,In_3066,In_3067,In_3068,In_3069,In_3070,In_3071,In_3072,In_3073,In_3074,In_3075,In_3076,In_3077,In_3078,In_3079,In_3080,In_3081,In_3082,In_3083,In_3084,In_3085,In_3086,In_3087,In_3088,In_3089,In_3090,In_3091,In_3092,In_3093,In_3094,In_3095,In_3096,In_3097,In_3098,In_3099,In_3100,In_3101,In_3102,In_3103,In_3104,In_3105,In_3106,In_3107,In_3108,In_3109,In_3110,In_3111,In_3112,In_3113,In_3114,In_3115,In_3116,In_3117,In_3118,In_3119,In_3120,In_3121,In_3122,In_3123,In_3124,In_3125,In_3126,In_3127,In_3128,In_3129,In_3130,In_3131,In_3132,In_3133,In_3134,In_3135,In_3136,In_3137,In_3138,In_3139,In_3140,In_3141,In_3142,In_3143,In_3144,In_3145,In_3146,In_3147,In_3148,In_3149,In_3150,In_3151,In_3152,In_3153,In_3154,In_3155,In_3156,In_3157,In_3158,In_3159,In_3160,In_3161,In_3162,In_3163,In_3164,In_3165,In_3166,In_3167,In_3168,In_3169,In_3170,In_3171,In_3172,In_3173,In_3174,In_3175,In_3176,In_3177,In_3178,In_3179,In_3180,In_3181,In_3182,In_3183,In_3184,In_3185,In_3186,In_3187,In_3188,In_3189,In_3190,In_3191,In_3192,In_3193,In_3194,In_3195,In_3196,In_3197,In_3198,In_3199,In_3200,In_3201,In_3202,In_3203,In_3204,In_3205,In_3206,In_3207,In_3208,In_3209,In_3210,In_3211,In_3212,In_3213,In_3214,In_3215,In_3216,In_3217,In_3218,In_3219,In_3220,In_3221,In_3222,In_3223,In_3224,In_3225,In_3226,In_3227,In_3228,In_3229,In_3230,In_3231,In_3232,In_3233,In_3234,In_3235,In_3236,In_3237,In_3238,In_3239,In_3240,In_3241,In_3242,In_3243,In_3244,In_3245,In_3246,In_3247,In_3248,In_3249,In_3250,In_3251,In_3252,In_3253,In_3254,In_3255,In_3256,In_3257,In_3258,In_3259,In_3260,In_3261,In_3262,In_3263,In_3264,In_3265,In_3266,In_3267,In_3268,In_3269,In_3270,In_3271,In_3272,In_3273,In_3274,In_3275,In_3276,In_3277,In_3278,In_3279,In_3280,In_3281,In_3282,In_3283,In_3284,In_3285,In_3286,In_3287,In_3288,In_3289,In_3290,In_3291,In_3292,In_3293,In_3294,In_3295,In_3296,In_3297,In_3298,In_3299,In_3300,In_3301,In_3302,In_3303,In_3304,In_3305,In_3306,In_3307,In_3308,In_3309,In_3310,In_3311,In_3312,In_3313,In_3314,In_3315,In_3316,In_3317,In_3318,In_3319,In_3320,In_3321,In_3322,In_3323,In_3324,In_3325,In_3326,In_3327,In_3328,In_3329,In_3330,In_3331,In_3332,In_3333,In_3334,In_3335,In_3336,In_3337,In_3338,In_3339,In_3340,In_3341,In_3342,In_3343,In_3344,In_3345,In_3346,In_3347,In_3348,In_3349,In_3350,In_3351,In_3352,In_3353,In_3354,In_3355,In_3356,In_3357,In_3358,In_3359,In_3360,In_3361,In_3362,In_3363,In_3364,In_3365,In_3366,In_3367,In_3368,In_3369,In_3370,In_3371,In_3372,In_3373,In_3374,In_3375,In_3376,In_3377,In_3378,In_3379,In_3380,In_3381,In_3382,In_3383,In_3384,In_3385,In_3386,In_3387,In_3388,In_3389,In_3390,In_3391,In_3392,In_3393,In_3394,In_3395,In_3396,In_3397,In_3398,In_3399,In_3400,In_3401,In_3402,In_3403,In_3404,In_3405,In_3406,In_3407,In_3408,In_3409,In_3410,In_3411,In_3412,In_3413,In_3414,In_3415,In_3416,In_3417,In_3418,In_3419,In_3420,In_3421,In_3422,In_3423,In_3424,In_3425,In_3426,In_3427,In_3428,In_3429,In_3430,In_3431,In_3432,In_3433,In_3434,In_3435,In_3436,In_3437,In_3438,In_3439,In_3440,In_3441,In_3442,In_3443,In_3444,In_3445,In_3446,In_3447,In_3448,In_3449,In_3450,In_3451,In_3452,In_3453,In_3454,In_3455,In_3456,In_3457,In_3458,In_3459,In_3460,In_3461,In_3462,In_3463,In_3464,In_3465,In_3466,In_3467,In_3468,In_3469,In_3470,In_3471,In_3472,In_3473,In_3474,In_3475,In_3476,In_3477,In_3478,In_3479,In_3480,In_3481,In_3482,In_3483,In_3484,In_3485,In_3486,In_3487,In_3488,In_3489,In_3490,In_3491,In_3492,In_3493,In_3494,In_3495,In_3496,In_3497,In_3498,In_3499,In_3500,In_3501,In_3502,In_3503,In_3504,In_3505,In_3506,In_3507,In_3508,In_3509,In_3510,In_3511,In_3512,In_3513,In_3514,In_3515,In_3516,In_3517,In_3518,In_3519,In_3520,In_3521,In_3522,In_3523,In_3524,In_3525,In_3526,In_3527,In_3528,In_3529,In_3530,In_3531,In_3532,In_3533,In_3534,In_3535,In_3536,In_3537,In_3538,In_3539,In_3540,In_3541,In_3542,In_3543,In_3544,In_3545,In_3546,In_3547,In_3548,In_3549,In_3550,In_3551,In_3552,In_3553,In_3554,In_3555,In_3556,In_3557,In_3558,In_3559,In_3560,In_3561,In_3562,In_3563,In_3564,In_3565,In_3566,In_3567,In_3568,In_3569,In_3570,In_3571,In_3572,In_3573,In_3574,In_3575,In_3576,In_3577,In_3578,In_3579,In_3580,In_3581,In_3582,In_3583,In_3584,In_3585,In_3586,In_3587,In_3588,In_3589,In_3590,In_3591,In_3592,In_3593,In_3594,In_3595,In_3596,In_3597,In_3598,In_3599,In_3600,In_3601,In_3602,In_3603,In_3604,In_3605,In_3606,In_3607,In_3608,In_3609,In_3610,In_3611,In_3612,In_3613,In_3614,In_3615,In_3616,In_3617,In_3618,In_3619,In_3620,In_3621,In_3622,In_3623,In_3624,In_3625,In_3626,In_3627,In_3628,In_3629,In_3630,In_3631,In_3632,In_3633,In_3634,In_3635,In_3636,In_3637,In_3638,In_3639,In_3640,In_3641,In_3642,In_3643,In_3644,In_3645,In_3646,In_3647,In_3648,In_3649,In_3650,In_3651,In_3652,In_3653,In_3654,In_3655,In_3656,In_3657,In_3658,In_3659,In_3660,In_3661,In_3662,In_3663,In_3664,In_3665,In_3666,In_3667,In_3668,In_3669,In_3670,In_3671,In_3672,In_3673,In_3674,In_3675,In_3676,In_3677,In_3678,In_3679,In_3680,In_3681,In_3682,In_3683,In_3684,In_3685,In_3686,In_3687,In_3688,In_3689,In_3690,In_3691,In_3692,In_3693,In_3694,In_3695,In_3696,In_3697,In_3698,In_3699,In_3700,In_3701,In_3702,In_3703,In_3704,In_3705,In_3706,In_3707,In_3708,In_3709,In_3710,In_3711,In_3712,In_3713,In_3714,In_3715,In_3716,In_3717,In_3718,In_3719,In_3720,In_3721,In_3722,In_3723,In_3724,In_3725,In_3726,In_3727,In_3728,In_3729,In_3730,In_3731,In_3732,In_3733,In_3734,In_3735,In_3736,In_3737,In_3738,In_3739,In_3740,In_3741,In_3742,In_3743,In_3744,In_3745,In_3746,In_3747,In_3748,In_3749,In_3750,In_3751,In_3752,In_3753,In_3754,In_3755,In_3756,In_3757,In_3758,In_3759,In_3760,In_3761,In_3762,In_3763,In_3764,In_3765,In_3766,In_3767,In_3768,In_3769,In_3770,In_3771,In_3772,In_3773,In_3774,In_3775,In_3776,In_3777,In_3778,In_3779,In_3780,In_3781,In_3782,In_3783,In_3784,In_3785,In_3786,In_3787,In_3788,In_3789,In_3790,In_3791,In_3792,In_3793,In_3794,In_3795,In_3796,In_3797,In_3798,In_3799,In_3800,In_3801,In_3802,In_3803,In_3804,In_3805,In_3806,In_3807,In_3808,In_3809,In_3810,In_3811,In_3812,In_3813,In_3814,In_3815,In_3816,In_3817,In_3818,In_3819,In_3820,In_3821,In_3822,In_3823,In_3824,In_3825,In_3826,In_3827,In_3828,In_3829,In_3830,In_3831,In_3832,In_3833,In_3834,In_3835,In_3836,In_3837,In_3838,In_3839,In_3840,In_3841,In_3842,In_3843,In_3844,In_3845,In_3846,In_3847,In_3848,In_3849,In_3850,In_3851,In_3852,In_3853,In_3854,In_3855,In_3856,In_3857,In_3858,In_3859,In_3860,In_3861,In_3862,In_3863,In_3864,In_3865,In_3866,In_3867,In_3868,In_3869,In_3870,In_3871,In_3872,In_3873,In_3874,In_3875,In_3876,In_3877,In_3878,In_3879,In_3880,In_3881,In_3882,In_3883,In_3884,In_3885,In_3886,In_3887,In_3888,In_3889,In_3890,In_3891,In_3892,In_3893,In_3894,In_3895,In_3896,In_3897,In_3898,In_3899,In_3900,In_3901,In_3902,In_3903,In_3904,In_3905,In_3906,In_3907,In_3908,In_3909,In_3910,In_3911,In_3912,In_3913,In_3914,In_3915,In_3916,In_3917,In_3918,In_3919,In_3920,In_3921,In_3922,In_3923,In_3924,In_3925,In_3926,In_3927,In_3928,In_3929,In_3930,In_3931,In_3932,In_3933,In_3934,In_3935,In_3936,In_3937,In_3938,In_3939,In_3940,In_3941,In_3942,In_3943,In_3944,In_3945,In_3946,In_3947,In_3948,In_3949,In_3950,In_3951,In_3952,In_3953,In_3954,In_3955,In_3956,In_3957,In_3958,In_3959,In_3960,In_3961,In_3962,In_3963,In_3964,In_3965,In_3966,In_3967,In_3968,In_3969,In_3970,In_3971,In_3972,In_3973,In_3974,In_3975,In_3976,In_3977,In_3978,In_3979,In_3980,In_3981,In_3982,In_3983,In_3984,In_3985,In_3986,In_3987,In_3988,In_3989,In_3990,In_3991,In_3992,In_3993,In_3994,In_3995,In_3996,In_3997,In_3998,In_3999,In_4000,In_4001,In_4002,In_4003,In_4004,In_4005,In_4006,In_4007,In_4008,In_4009,In_4010,In_4011,In_4012,In_4013,In_4014,In_4015,In_4016,In_4017,In_4018,In_4019,In_4020,In_4021,In_4022,In_4023,In_4024,In_4025,In_4026,In_4027,In_4028,In_4029,In_4030,In_4031,In_4032,In_4033,In_4034,In_4035,In_4036,In_4037,In_4038,In_4039,In_4040,In_4041,In_4042,In_4043,In_4044,In_4045,In_4046,In_4047,In_4048,In_4049,In_4050,In_4051,In_4052,In_4053,In_4054,In_4055,In_4056,In_4057,In_4058,In_4059,In_4060,In_4061,In_4062,In_4063,In_4064,In_4065,In_4066,In_4067,In_4068,In_4069,In_4070,In_4071,In_4072,In_4073,In_4074,In_4075,In_4076,In_4077,In_4078,In_4079,In_4080,In_4081,In_4082,In_4083,In_4084,In_4085,In_4086,In_4087,In_4088,In_4089,In_4090,In_4091,In_4092,In_4093,In_4094,In_4095,In_4096,In_4097,In_4098,In_4099,In_4100,In_4101,In_4102,In_4103,In_4104,In_4105,In_4106,In_4107,In_4108,In_4109,In_4110,In_4111,In_4112,In_4113,In_4114,In_4115,In_4116,In_4117,In_4118,In_4119,In_4120,In_4121,In_4122,In_4123,In_4124,In_4125,In_4126,In_4127,In_4128,In_4129,In_4130,In_4131,In_4132,In_4133,In_4134,In_4135,In_4136,In_4137,In_4138,In_4139,In_4140,In_4141,In_4142,In_4143,In_4144,In_4145,In_4146,In_4147,In_4148,In_4149,In_4150,In_4151,In_4152,In_4153,In_4154,In_4155,In_4156,In_4157,In_4158,In_4159,In_4160,In_4161,In_4162,In_4163,In_4164,In_4165,In_4166,In_4167,In_4168,In_4169,In_4170,In_4171,In_4172,In_4173,In_4174,In_4175,In_4176,In_4177,In_4178,In_4179,In_4180,In_4181,In_4182,In_4183,In_4184,In_4185,In_4186,In_4187,In_4188,In_4189,In_4190,In_4191,In_4192,In_4193,In_4194,In_4195,In_4196,In_4197,In_4198,In_4199,In_4200,In_4201,In_4202,In_4203,In_4204,In_4205,In_4206,In_4207,In_4208,In_4209,In_4210,In_4211,In_4212,In_4213,In_4214,In_4215,In_4216,In_4217,In_4218,In_4219,In_4220,In_4221,In_4222,In_4223,In_4224,In_4225,In_4226,In_4227,In_4228,In_4229,In_4230,In_4231,In_4232,In_4233,In_4234,In_4235,In_4236,In_4237,In_4238,In_4239,In_4240,In_4241,In_4242,In_4243,In_4244,In_4245,In_4246,In_4247,In_4248,In_4249,In_4250,In_4251,In_4252,In_4253,In_4254,In_4255,In_4256,In_4257,In_4258,In_4259,In_4260,In_4261,In_4262,In_4263,In_4264,In_4265,In_4266,In_4267,In_4268,In_4269,In_4270,In_4271,In_4272,In_4273,In_4274,In_4275,In_4276,In_4277,In_4278,In_4279,In_4280,In_4281,In_4282,In_4283,In_4284,In_4285,In_4286,In_4287,In_4288,In_4289,In_4290,In_4291,In_4292,In_4293,In_4294,In_4295,In_4296,In_4297,In_4298,In_4299,In_4300,In_4301,In_4302,In_4303,In_4304,In_4305,In_4306,In_4307,In_4308,In_4309,In_4310,In_4311,In_4312,In_4313,In_4314,In_4315,In_4316,In_4317,In_4318,In_4319,In_4320,In_4321,In_4322,In_4323,In_4324,In_4325,In_4326,In_4327,In_4328,In_4329,In_4330,In_4331,In_4332,In_4333,In_4334,In_4335,In_4336,In_4337,In_4338,In_4339,In_4340,In_4341,In_4342,In_4343,In_4344,In_4345,In_4346,In_4347,In_4348,In_4349,In_4350,In_4351,In_4352,In_4353,In_4354,In_4355,In_4356,In_4357,In_4358,In_4359,In_4360,In_4361,In_4362,In_4363,In_4364,In_4365,In_4366,In_4367,In_4368,In_4369,In_4370,In_4371,In_4372,In_4373,In_4374,In_4375,In_4376,In_4377,In_4378,In_4379,In_4380,In_4381,In_4382,In_4383,In_4384,In_4385,In_4386,In_4387,In_4388,In_4389,In_4390,In_4391,In_4392,In_4393,In_4394,In_4395,In_4396,In_4397,In_4398,In_4399,In_4400,In_4401,In_4402,In_4403,In_4404,In_4405,In_4406,In_4407,In_4408,In_4409,In_4410,In_4411,In_4412,In_4413,In_4414,In_4415,In_4416,In_4417,In_4418,In_4419,In_4420,In_4421,In_4422,In_4423,In_4424,In_4425,In_4426,In_4427,In_4428,In_4429,In_4430,In_4431,In_4432,In_4433,In_4434,In_4435,In_4436,In_4437,In_4438,In_4439,In_4440,In_4441,In_4442,In_4443,In_4444,In_4445,In_4446,In_4447,In_4448,In_4449,In_4450,In_4451,In_4452,In_4453,In_4454,In_4455,In_4456,In_4457,In_4458,In_4459,In_4460,In_4461,In_4462,In_4463,In_4464,In_4465,In_4466,In_4467,In_4468,In_4469,In_4470,In_4471,In_4472,In_4473,In_4474,In_4475,In_4476,In_4477,In_4478,In_4479,In_4480,In_4481,In_4482,In_4483,In_4484,In_4485,In_4486,In_4487,In_4488,In_4489,In_4490,In_4491,In_4492,In_4493,In_4494,In_4495,In_4496,In_4497,In_4498,In_4499,In_4500,In_4501,In_4502,In_4503,In_4504,In_4505,In_4506,In_4507,In_4508,In_4509,In_4510,In_4511,In_4512,In_4513,In_4514,In_4515,In_4516,In_4517,In_4518,In_4519,In_4520,In_4521,In_4522,In_4523,In_4524,In_4525,In_4526,In_4527,In_4528,In_4529,In_4530,In_4531,In_4532,In_4533,In_4534,In_4535,In_4536,In_4537,In_4538,In_4539,In_4540,In_4541,In_4542,In_4543,In_4544,In_4545,In_4546,In_4547,In_4548,In_4549,In_4550,In_4551,In_4552,In_4553,In_4554,In_4555,In_4556,In_4557,In_4558,In_4559,In_4560,In_4561,In_4562,In_4563,In_4564,In_4565,In_4566,In_4567,In_4568,In_4569,In_4570,In_4571,In_4572,In_4573,In_4574,In_4575,In_4576,In_4577,In_4578,In_4579,In_4580,In_4581,In_4582,In_4583,In_4584,In_4585,In_4586,In_4587,In_4588,In_4589,In_4590,In_4591,In_4592,In_4593,In_4594,In_4595,In_4596,In_4597,In_4598,In_4599,In_4600,In_4601,In_4602,In_4603,In_4604,In_4605,In_4606,In_4607,In_4608,In_4609,In_4610,In_4611,In_4612,In_4613,In_4614,In_4615,In_4616,In_4617,In_4618,In_4619,In_4620,In_4621,In_4622,In_4623,In_4624,In_4625,In_4626,In_4627,In_4628,In_4629,In_4630,In_4631,In_4632,In_4633,In_4634,In_4635,In_4636,In_4637,In_4638,In_4639,In_4640,In_4641,In_4642,In_4643,In_4644,In_4645,In_4646,In_4647,In_4648,In_4649,In_4650,In_4651,In_4652,In_4653,In_4654,In_4655,In_4656,In_4657,In_4658,In_4659,In_4660,In_4661,In_4662,In_4663,In_4664,In_4665,In_4666,In_4667,In_4668,In_4669,In_4670,In_4671,In_4672,In_4673,In_4674,In_4675,In_4676,In_4677,In_4678,In_4679,In_4680,In_4681,In_4682,In_4683,In_4684,In_4685,In_4686,In_4687,In_4688,In_4689,In_4690,In_4691,In_4692,In_4693,In_4694,In_4695,In_4696,In_4697,In_4698,In_4699,In_4700,In_4701,In_4702,In_4703,In_4704,In_4705,In_4706,In_4707,In_4708,In_4709,In_4710,In_4711,In_4712,In_4713,In_4714,In_4715,In_4716,In_4717,In_4718,In_4719,In_4720,In_4721,In_4722,In_4723,In_4724,In_4725,In_4726,In_4727,In_4728,In_4729,In_4730,In_4731,In_4732,In_4733,In_4734,In_4735,In_4736,In_4737,In_4738,In_4739,In_4740,In_4741,In_4742,In_4743,In_4744,In_4745,In_4746,In_4747,In_4748,In_4749,In_4750,In_4751,In_4752,In_4753,In_4754,In_4755,In_4756,In_4757,In_4758,In_4759,In_4760,In_4761,In_4762,In_4763,In_4764,In_4765,In_4766,In_4767,In_4768,In_4769,In_4770,In_4771,In_4772,In_4773,In_4774,In_4775,In_4776,In_4777,In_4778,In_4779,In_4780,In_4781,In_4782,In_4783,In_4784,In_4785,In_4786,In_4787,In_4788,In_4789,In_4790,In_4791,In_4792,In_4793,In_4794,In_4795,In_4796,In_4797,In_4798,In_4799,In_4800,In_4801,In_4802,In_4803,In_4804,In_4805,In_4806,In_4807,In_4808,In_4809,In_4810,In_4811,In_4812,In_4813,In_4814,In_4815,In_4816,In_4817,In_4818,In_4819,In_4820,In_4821,In_4822,In_4823,In_4824,In_4825,In_4826,In_4827,In_4828,In_4829,In_4830,In_4831,In_4832,In_4833,In_4834,In_4835,In_4836,In_4837,In_4838,In_4839,In_4840,In_4841,In_4842,In_4843,In_4844,In_4845,In_4846,In_4847,In_4848,In_4849,In_4850,In_4851,In_4852,In_4853,In_4854,In_4855,In_4856,In_4857,In_4858,In_4859,In_4860,In_4861,In_4862,In_4863,In_4864,In_4865,In_4866,In_4867,In_4868,In_4869,In_4870,In_4871,In_4872,In_4873,In_4874,In_4875,In_4876,In_4877,In_4878,In_4879,In_4880,In_4881,In_4882,In_4883,In_4884,In_4885,In_4886,In_4887,In_4888,In_4889,In_4890,In_4891,In_4892,In_4893,In_4894,In_4895,In_4896,In_4897,In_4898,In_4899,In_4900,In_4901,In_4902,In_4903,In_4904,In_4905,In_4906,In_4907,In_4908,In_4909,In_4910,In_4911,In_4912,In_4913,In_4914,In_4915,In_4916,In_4917,In_4918,In_4919,In_4920,In_4921,In_4922,In_4923,In_4924,In_4925,In_4926,In_4927,In_4928,In_4929,In_4930,In_4931,In_4932,In_4933,In_4934,In_4935,In_4936,In_4937,In_4938,In_4939,In_4940,In_4941,In_4942,In_4943,In_4944,In_4945,In_4946,In_4947,In_4948,In_4949,In_4950,In_4951,In_4952,In_4953,In_4954,In_4955,In_4956,In_4957,In_4958,In_4959,In_4960,In_4961,In_4962,In_4963,In_4964,In_4965,In_4966,In_4967,In_4968,In_4969,In_4970,In_4971,In_4972,In_4973,In_4974,In_4975,In_4976,In_4977,In_4978,In_4979,In_4980,In_4981,In_4982,In_4983,In_4984,In_4985,In_4986,In_4987,In_4988,In_4989,In_4990,In_4991,In_4992,In_4993,In_4994,In_4995,In_4996,In_4997,In_4998,In_4999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499,O_3500,O_3501,O_3502,O_3503,O_3504,O_3505,O_3506,O_3507,O_3508,O_3509,O_3510,O_3511,O_3512,O_3513,O_3514,O_3515,O_3516,O_3517,O_3518,O_3519,O_3520,O_3521,O_3522,O_3523,O_3524,O_3525,O_3526,O_3527,O_3528,O_3529,O_3530,O_3531,O_3532,O_3533,O_3534,O_3535,O_3536,O_3537,O_3538,O_3539,O_3540,O_3541,O_3542,O_3543,O_3544,O_3545,O_3546,O_3547,O_3548,O_3549,O_3550,O_3551,O_3552,O_3553,O_3554,O_3555,O_3556,O_3557,O_3558,O_3559,O_3560,O_3561,O_3562,O_3563,O_3564,O_3565,O_3566,O_3567,O_3568,O_3569,O_3570,O_3571,O_3572,O_3573,O_3574,O_3575,O_3576,O_3577,O_3578,O_3579,O_3580,O_3581,O_3582,O_3583,O_3584,O_3585,O_3586,O_3587,O_3588,O_3589,O_3590,O_3591,O_3592,O_3593,O_3594,O_3595,O_3596,O_3597,O_3598,O_3599,O_3600,O_3601,O_3602,O_3603,O_3604,O_3605,O_3606,O_3607,O_3608,O_3609,O_3610,O_3611,O_3612,O_3613,O_3614,O_3615,O_3616,O_3617,O_3618,O_3619,O_3620,O_3621,O_3622,O_3623,O_3624,O_3625,O_3626,O_3627,O_3628,O_3629,O_3630,O_3631,O_3632,O_3633,O_3634,O_3635,O_3636,O_3637,O_3638,O_3639,O_3640,O_3641,O_3642,O_3643,O_3644,O_3645,O_3646,O_3647,O_3648,O_3649,O_3650,O_3651,O_3652,O_3653,O_3654,O_3655,O_3656,O_3657,O_3658,O_3659,O_3660,O_3661,O_3662,O_3663,O_3664,O_3665,O_3666,O_3667,O_3668,O_3669,O_3670,O_3671,O_3672,O_3673,O_3674,O_3675,O_3676,O_3677,O_3678,O_3679,O_3680,O_3681,O_3682,O_3683,O_3684,O_3685,O_3686,O_3687,O_3688,O_3689,O_3690,O_3691,O_3692,O_3693,O_3694,O_3695,O_3696,O_3697,O_3698,O_3699,O_3700,O_3701,O_3702,O_3703,O_3704,O_3705,O_3706,O_3707,O_3708,O_3709,O_3710,O_3711,O_3712,O_3713,O_3714,O_3715,O_3716,O_3717,O_3718,O_3719,O_3720,O_3721,O_3722,O_3723,O_3724,O_3725,O_3726,O_3727,O_3728,O_3729,O_3730,O_3731,O_3732,O_3733,O_3734,O_3735,O_3736,O_3737,O_3738,O_3739,O_3740,O_3741,O_3742,O_3743,O_3744,O_3745,O_3746,O_3747,O_3748,O_3749,O_3750,O_3751,O_3752,O_3753,O_3754,O_3755,O_3756,O_3757,O_3758,O_3759,O_3760,O_3761,O_3762,O_3763,O_3764,O_3765,O_3766,O_3767,O_3768,O_3769,O_3770,O_3771,O_3772,O_3773,O_3774,O_3775,O_3776,O_3777,O_3778,O_3779,O_3780,O_3781,O_3782,O_3783,O_3784,O_3785,O_3786,O_3787,O_3788,O_3789,O_3790,O_3791,O_3792,O_3793,O_3794,O_3795,O_3796,O_3797,O_3798,O_3799,O_3800,O_3801,O_3802,O_3803,O_3804,O_3805,O_3806,O_3807,O_3808,O_3809,O_3810,O_3811,O_3812,O_3813,O_3814,O_3815,O_3816,O_3817,O_3818,O_3819,O_3820,O_3821,O_3822,O_3823,O_3824,O_3825,O_3826,O_3827,O_3828,O_3829,O_3830,O_3831,O_3832,O_3833,O_3834,O_3835,O_3836,O_3837,O_3838,O_3839,O_3840,O_3841,O_3842,O_3843,O_3844,O_3845,O_3846,O_3847,O_3848,O_3849,O_3850,O_3851,O_3852,O_3853,O_3854,O_3855,O_3856,O_3857,O_3858,O_3859,O_3860,O_3861,O_3862,O_3863,O_3864,O_3865,O_3866,O_3867,O_3868,O_3869,O_3870,O_3871,O_3872,O_3873,O_3874,O_3875,O_3876,O_3877,O_3878,O_3879,O_3880,O_3881,O_3882,O_3883,O_3884,O_3885,O_3886,O_3887,O_3888,O_3889,O_3890,O_3891,O_3892,O_3893,O_3894,O_3895,O_3896,O_3897,O_3898,O_3899,O_3900,O_3901,O_3902,O_3903,O_3904,O_3905,O_3906,O_3907,O_3908,O_3909,O_3910,O_3911,O_3912,O_3913,O_3914,O_3915,O_3916,O_3917,O_3918,O_3919,O_3920,O_3921,O_3922,O_3923,O_3924,O_3925,O_3926,O_3927,O_3928,O_3929,O_3930,O_3931,O_3932,O_3933,O_3934,O_3935,O_3936,O_3937,O_3938,O_3939,O_3940,O_3941,O_3942,O_3943,O_3944,O_3945,O_3946,O_3947,O_3948,O_3949,O_3950,O_3951,O_3952,O_3953,O_3954,O_3955,O_3956,O_3957,O_3958,O_3959,O_3960,O_3961,O_3962,O_3963,O_3964,O_3965,O_3966,O_3967,O_3968,O_3969,O_3970,O_3971,O_3972,O_3973,O_3974,O_3975,O_3976,O_3977,O_3978,O_3979,O_3980,O_3981,O_3982,O_3983,O_3984,O_3985,O_3986,O_3987,O_3988,O_3989,O_3990,O_3991,O_3992,O_3993,O_3994,O_3995,O_3996,O_3997,O_3998,O_3999,O_4000,O_4001,O_4002,O_4003,O_4004,O_4005,O_4006,O_4007,O_4008,O_4009,O_4010,O_4011,O_4012,O_4013,O_4014,O_4015,O_4016,O_4017,O_4018,O_4019,O_4020,O_4021,O_4022,O_4023,O_4024,O_4025,O_4026,O_4027,O_4028,O_4029,O_4030,O_4031,O_4032,O_4033,O_4034,O_4035,O_4036,O_4037,O_4038,O_4039,O_4040,O_4041,O_4042,O_4043,O_4044,O_4045,O_4046,O_4047,O_4048,O_4049,O_4050,O_4051,O_4052,O_4053,O_4054,O_4055,O_4056,O_4057,O_4058,O_4059,O_4060,O_4061,O_4062,O_4063,O_4064,O_4065,O_4066,O_4067,O_4068,O_4069,O_4070,O_4071,O_4072,O_4073,O_4074,O_4075,O_4076,O_4077,O_4078,O_4079,O_4080,O_4081,O_4082,O_4083,O_4084,O_4085,O_4086,O_4087,O_4088,O_4089,O_4090,O_4091,O_4092,O_4093,O_4094,O_4095,O_4096,O_4097,O_4098,O_4099,O_4100,O_4101,O_4102,O_4103,O_4104,O_4105,O_4106,O_4107,O_4108,O_4109,O_4110,O_4111,O_4112,O_4113,O_4114,O_4115,O_4116,O_4117,O_4118,O_4119,O_4120,O_4121,O_4122,O_4123,O_4124,O_4125,O_4126,O_4127,O_4128,O_4129,O_4130,O_4131,O_4132,O_4133,O_4134,O_4135,O_4136,O_4137,O_4138,O_4139,O_4140,O_4141,O_4142,O_4143,O_4144,O_4145,O_4146,O_4147,O_4148,O_4149,O_4150,O_4151,O_4152,O_4153,O_4154,O_4155,O_4156,O_4157,O_4158,O_4159,O_4160,O_4161,O_4162,O_4163,O_4164,O_4165,O_4166,O_4167,O_4168,O_4169,O_4170,O_4171,O_4172,O_4173,O_4174,O_4175,O_4176,O_4177,O_4178,O_4179,O_4180,O_4181,O_4182,O_4183,O_4184,O_4185,O_4186,O_4187,O_4188,O_4189,O_4190,O_4191,O_4192,O_4193,O_4194,O_4195,O_4196,O_4197,O_4198,O_4199,O_4200,O_4201,O_4202,O_4203,O_4204,O_4205,O_4206,O_4207,O_4208,O_4209,O_4210,O_4211,O_4212,O_4213,O_4214,O_4215,O_4216,O_4217,O_4218,O_4219,O_4220,O_4221,O_4222,O_4223,O_4224,O_4225,O_4226,O_4227,O_4228,O_4229,O_4230,O_4231,O_4232,O_4233,O_4234,O_4235,O_4236,O_4237,O_4238,O_4239,O_4240,O_4241,O_4242,O_4243,O_4244,O_4245,O_4246,O_4247,O_4248,O_4249,O_4250,O_4251,O_4252,O_4253,O_4254,O_4255,O_4256,O_4257,O_4258,O_4259,O_4260,O_4261,O_4262,O_4263,O_4264,O_4265,O_4266,O_4267,O_4268,O_4269,O_4270,O_4271,O_4272,O_4273,O_4274,O_4275,O_4276,O_4277,O_4278,O_4279,O_4280,O_4281,O_4282,O_4283,O_4284,O_4285,O_4286,O_4287,O_4288,O_4289,O_4290,O_4291,O_4292,O_4293,O_4294,O_4295,O_4296,O_4297,O_4298,O_4299,O_4300,O_4301,O_4302,O_4303,O_4304,O_4305,O_4306,O_4307,O_4308,O_4309,O_4310,O_4311,O_4312,O_4313,O_4314,O_4315,O_4316,O_4317,O_4318,O_4319,O_4320,O_4321,O_4322,O_4323,O_4324,O_4325,O_4326,O_4327,O_4328,O_4329,O_4330,O_4331,O_4332,O_4333,O_4334,O_4335,O_4336,O_4337,O_4338,O_4339,O_4340,O_4341,O_4342,O_4343,O_4344,O_4345,O_4346,O_4347,O_4348,O_4349,O_4350,O_4351,O_4352,O_4353,O_4354,O_4355,O_4356,O_4357,O_4358,O_4359,O_4360,O_4361,O_4362,O_4363,O_4364,O_4365,O_4366,O_4367,O_4368,O_4369,O_4370,O_4371,O_4372,O_4373,O_4374,O_4375,O_4376,O_4377,O_4378,O_4379,O_4380,O_4381,O_4382,O_4383,O_4384,O_4385,O_4386,O_4387,O_4388,O_4389,O_4390,O_4391,O_4392,O_4393,O_4394,O_4395,O_4396,O_4397,O_4398,O_4399,O_4400,O_4401,O_4402,O_4403,O_4404,O_4405,O_4406,O_4407,O_4408,O_4409,O_4410,O_4411,O_4412,O_4413,O_4414,O_4415,O_4416,O_4417,O_4418,O_4419,O_4420,O_4421,O_4422,O_4423,O_4424,O_4425,O_4426,O_4427,O_4428,O_4429,O_4430,O_4431,O_4432,O_4433,O_4434,O_4435,O_4436,O_4437,O_4438,O_4439,O_4440,O_4441,O_4442,O_4443,O_4444,O_4445,O_4446,O_4447,O_4448,O_4449,O_4450,O_4451,O_4452,O_4453,O_4454,O_4455,O_4456,O_4457,O_4458,O_4459,O_4460,O_4461,O_4462,O_4463,O_4464,O_4465,O_4466,O_4467,O_4468,O_4469,O_4470,O_4471,O_4472,O_4473,O_4474,O_4475,O_4476,O_4477,O_4478,O_4479,O_4480,O_4481,O_4482,O_4483,O_4484,O_4485,O_4486,O_4487,O_4488,O_4489,O_4490,O_4491,O_4492,O_4493,O_4494,O_4495,O_4496,O_4497,O_4498,O_4499,O_4500,O_4501,O_4502,O_4503,O_4504,O_4505,O_4506,O_4507,O_4508,O_4509,O_4510,O_4511,O_4512,O_4513,O_4514,O_4515,O_4516,O_4517,O_4518,O_4519,O_4520,O_4521,O_4522,O_4523,O_4524,O_4525,O_4526,O_4527,O_4528,O_4529,O_4530,O_4531,O_4532,O_4533,O_4534,O_4535,O_4536,O_4537,O_4538,O_4539,O_4540,O_4541,O_4542,O_4543,O_4544,O_4545,O_4546,O_4547,O_4548,O_4549,O_4550,O_4551,O_4552,O_4553,O_4554,O_4555,O_4556,O_4557,O_4558,O_4559,O_4560,O_4561,O_4562,O_4563,O_4564,O_4565,O_4566,O_4567,O_4568,O_4569,O_4570,O_4571,O_4572,O_4573,O_4574,O_4575,O_4576,O_4577,O_4578,O_4579,O_4580,O_4581,O_4582,O_4583,O_4584,O_4585,O_4586,O_4587,O_4588,O_4589,O_4590,O_4591,O_4592,O_4593,O_4594,O_4595,O_4596,O_4597,O_4598,O_4599,O_4600,O_4601,O_4602,O_4603,O_4604,O_4605,O_4606,O_4607,O_4608,O_4609,O_4610,O_4611,O_4612,O_4613,O_4614,O_4615,O_4616,O_4617,O_4618,O_4619,O_4620,O_4621,O_4622,O_4623,O_4624,O_4625,O_4626,O_4627,O_4628,O_4629,O_4630,O_4631,O_4632,O_4633,O_4634,O_4635,O_4636,O_4637,O_4638,O_4639,O_4640,O_4641,O_4642,O_4643,O_4644,O_4645,O_4646,O_4647,O_4648,O_4649,O_4650,O_4651,O_4652,O_4653,O_4654,O_4655,O_4656,O_4657,O_4658,O_4659,O_4660,O_4661,O_4662,O_4663,O_4664,O_4665,O_4666,O_4667,O_4668,O_4669,O_4670,O_4671,O_4672,O_4673,O_4674,O_4675,O_4676,O_4677,O_4678,O_4679,O_4680,O_4681,O_4682,O_4683,O_4684,O_4685,O_4686,O_4687,O_4688,O_4689,O_4690,O_4691,O_4692,O_4693,O_4694,O_4695,O_4696,O_4697,O_4698,O_4699,O_4700,O_4701,O_4702,O_4703,O_4704,O_4705,O_4706,O_4707,O_4708,O_4709,O_4710,O_4711,O_4712,O_4713,O_4714,O_4715,O_4716,O_4717,O_4718,O_4719,O_4720,O_4721,O_4722,O_4723,O_4724,O_4725,O_4726,O_4727,O_4728,O_4729,O_4730,O_4731,O_4732,O_4733,O_4734,O_4735,O_4736,O_4737,O_4738,O_4739,O_4740,O_4741,O_4742,O_4743,O_4744,O_4745,O_4746,O_4747,O_4748,O_4749,O_4750,O_4751,O_4752,O_4753,O_4754,O_4755,O_4756,O_4757,O_4758,O_4759,O_4760,O_4761,O_4762,O_4763,O_4764,O_4765,O_4766,O_4767,O_4768,O_4769,O_4770,O_4771,O_4772,O_4773,O_4774,O_4775,O_4776,O_4777,O_4778,O_4779,O_4780,O_4781,O_4782,O_4783,O_4784,O_4785,O_4786,O_4787,O_4788,O_4789,O_4790,O_4791,O_4792,O_4793,O_4794,O_4795,O_4796,O_4797,O_4798,O_4799,O_4800,O_4801,O_4802,O_4803,O_4804,O_4805,O_4806,O_4807,O_4808,O_4809,O_4810,O_4811,O_4812,O_4813,O_4814,O_4815,O_4816,O_4817,O_4818,O_4819,O_4820,O_4821,O_4822,O_4823,O_4824,O_4825,O_4826,O_4827,O_4828,O_4829,O_4830,O_4831,O_4832,O_4833,O_4834,O_4835,O_4836,O_4837,O_4838,O_4839,O_4840,O_4841,O_4842,O_4843,O_4844,O_4845,O_4846,O_4847,O_4848,O_4849,O_4850,O_4851,O_4852,O_4853,O_4854,O_4855,O_4856,O_4857,O_4858,O_4859,O_4860,O_4861,O_4862,O_4863,O_4864,O_4865,O_4866,O_4867,O_4868,O_4869,O_4870,O_4871,O_4872,O_4873,O_4874,O_4875,O_4876,O_4877,O_4878,O_4879,O_4880,O_4881,O_4882,O_4883,O_4884,O_4885,O_4886,O_4887,O_4888,O_4889,O_4890,O_4891,O_4892,O_4893,O_4894,O_4895,O_4896,O_4897,O_4898,O_4899,O_4900,O_4901,O_4902,O_4903,O_4904,O_4905,O_4906,O_4907,O_4908,O_4909,O_4910,O_4911,O_4912,O_4913,O_4914,O_4915,O_4916,O_4917,O_4918,O_4919,O_4920,O_4921,O_4922,O_4923,O_4924,O_4925,O_4926,O_4927,O_4928,O_4929,O_4930,O_4931,O_4932,O_4933,O_4934,O_4935,O_4936,O_4937,O_4938,O_4939,O_4940,O_4941,O_4942,O_4943,O_4944,O_4945,O_4946,O_4947,O_4948,O_4949,O_4950,O_4951,O_4952,O_4953,O_4954,O_4955,O_4956,O_4957,O_4958,O_4959,O_4960,O_4961,O_4962,O_4963,O_4964,O_4965,O_4966,O_4967,O_4968,O_4969,O_4970,O_4971,O_4972,O_4973,O_4974,O_4975,O_4976,O_4977,O_4978,O_4979,O_4980,O_4981,O_4982,O_4983,O_4984,O_4985,O_4986,O_4987,O_4988,O_4989,O_4990,O_4991,O_4992,O_4993,O_4994,O_4995,O_4996,O_4997,O_4998,O_4999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,In_3000,In_3001,In_3002,In_3003,In_3004,In_3005,In_3006,In_3007,In_3008,In_3009,In_3010,In_3011,In_3012,In_3013,In_3014,In_3015,In_3016,In_3017,In_3018,In_3019,In_3020,In_3021,In_3022,In_3023,In_3024,In_3025,In_3026,In_3027,In_3028,In_3029,In_3030,In_3031,In_3032,In_3033,In_3034,In_3035,In_3036,In_3037,In_3038,In_3039,In_3040,In_3041,In_3042,In_3043,In_3044,In_3045,In_3046,In_3047,In_3048,In_3049,In_3050,In_3051,In_3052,In_3053,In_3054,In_3055,In_3056,In_3057,In_3058,In_3059,In_3060,In_3061,In_3062,In_3063,In_3064,In_3065,In_3066,In_3067,In_3068,In_3069,In_3070,In_3071,In_3072,In_3073,In_3074,In_3075,In_3076,In_3077,In_3078,In_3079,In_3080,In_3081,In_3082,In_3083,In_3084,In_3085,In_3086,In_3087,In_3088,In_3089,In_3090,In_3091,In_3092,In_3093,In_3094,In_3095,In_3096,In_3097,In_3098,In_3099,In_3100,In_3101,In_3102,In_3103,In_3104,In_3105,In_3106,In_3107,In_3108,In_3109,In_3110,In_3111,In_3112,In_3113,In_3114,In_3115,In_3116,In_3117,In_3118,In_3119,In_3120,In_3121,In_3122,In_3123,In_3124,In_3125,In_3126,In_3127,In_3128,In_3129,In_3130,In_3131,In_3132,In_3133,In_3134,In_3135,In_3136,In_3137,In_3138,In_3139,In_3140,In_3141,In_3142,In_3143,In_3144,In_3145,In_3146,In_3147,In_3148,In_3149,In_3150,In_3151,In_3152,In_3153,In_3154,In_3155,In_3156,In_3157,In_3158,In_3159,In_3160,In_3161,In_3162,In_3163,In_3164,In_3165,In_3166,In_3167,In_3168,In_3169,In_3170,In_3171,In_3172,In_3173,In_3174,In_3175,In_3176,In_3177,In_3178,In_3179,In_3180,In_3181,In_3182,In_3183,In_3184,In_3185,In_3186,In_3187,In_3188,In_3189,In_3190,In_3191,In_3192,In_3193,In_3194,In_3195,In_3196,In_3197,In_3198,In_3199,In_3200,In_3201,In_3202,In_3203,In_3204,In_3205,In_3206,In_3207,In_3208,In_3209,In_3210,In_3211,In_3212,In_3213,In_3214,In_3215,In_3216,In_3217,In_3218,In_3219,In_3220,In_3221,In_3222,In_3223,In_3224,In_3225,In_3226,In_3227,In_3228,In_3229,In_3230,In_3231,In_3232,In_3233,In_3234,In_3235,In_3236,In_3237,In_3238,In_3239,In_3240,In_3241,In_3242,In_3243,In_3244,In_3245,In_3246,In_3247,In_3248,In_3249,In_3250,In_3251,In_3252,In_3253,In_3254,In_3255,In_3256,In_3257,In_3258,In_3259,In_3260,In_3261,In_3262,In_3263,In_3264,In_3265,In_3266,In_3267,In_3268,In_3269,In_3270,In_3271,In_3272,In_3273,In_3274,In_3275,In_3276,In_3277,In_3278,In_3279,In_3280,In_3281,In_3282,In_3283,In_3284,In_3285,In_3286,In_3287,In_3288,In_3289,In_3290,In_3291,In_3292,In_3293,In_3294,In_3295,In_3296,In_3297,In_3298,In_3299,In_3300,In_3301,In_3302,In_3303,In_3304,In_3305,In_3306,In_3307,In_3308,In_3309,In_3310,In_3311,In_3312,In_3313,In_3314,In_3315,In_3316,In_3317,In_3318,In_3319,In_3320,In_3321,In_3322,In_3323,In_3324,In_3325,In_3326,In_3327,In_3328,In_3329,In_3330,In_3331,In_3332,In_3333,In_3334,In_3335,In_3336,In_3337,In_3338,In_3339,In_3340,In_3341,In_3342,In_3343,In_3344,In_3345,In_3346,In_3347,In_3348,In_3349,In_3350,In_3351,In_3352,In_3353,In_3354,In_3355,In_3356,In_3357,In_3358,In_3359,In_3360,In_3361,In_3362,In_3363,In_3364,In_3365,In_3366,In_3367,In_3368,In_3369,In_3370,In_3371,In_3372,In_3373,In_3374,In_3375,In_3376,In_3377,In_3378,In_3379,In_3380,In_3381,In_3382,In_3383,In_3384,In_3385,In_3386,In_3387,In_3388,In_3389,In_3390,In_3391,In_3392,In_3393,In_3394,In_3395,In_3396,In_3397,In_3398,In_3399,In_3400,In_3401,In_3402,In_3403,In_3404,In_3405,In_3406,In_3407,In_3408,In_3409,In_3410,In_3411,In_3412,In_3413,In_3414,In_3415,In_3416,In_3417,In_3418,In_3419,In_3420,In_3421,In_3422,In_3423,In_3424,In_3425,In_3426,In_3427,In_3428,In_3429,In_3430,In_3431,In_3432,In_3433,In_3434,In_3435,In_3436,In_3437,In_3438,In_3439,In_3440,In_3441,In_3442,In_3443,In_3444,In_3445,In_3446,In_3447,In_3448,In_3449,In_3450,In_3451,In_3452,In_3453,In_3454,In_3455,In_3456,In_3457,In_3458,In_3459,In_3460,In_3461,In_3462,In_3463,In_3464,In_3465,In_3466,In_3467,In_3468,In_3469,In_3470,In_3471,In_3472,In_3473,In_3474,In_3475,In_3476,In_3477,In_3478,In_3479,In_3480,In_3481,In_3482,In_3483,In_3484,In_3485,In_3486,In_3487,In_3488,In_3489,In_3490,In_3491,In_3492,In_3493,In_3494,In_3495,In_3496,In_3497,In_3498,In_3499,In_3500,In_3501,In_3502,In_3503,In_3504,In_3505,In_3506,In_3507,In_3508,In_3509,In_3510,In_3511,In_3512,In_3513,In_3514,In_3515,In_3516,In_3517,In_3518,In_3519,In_3520,In_3521,In_3522,In_3523,In_3524,In_3525,In_3526,In_3527,In_3528,In_3529,In_3530,In_3531,In_3532,In_3533,In_3534,In_3535,In_3536,In_3537,In_3538,In_3539,In_3540,In_3541,In_3542,In_3543,In_3544,In_3545,In_3546,In_3547,In_3548,In_3549,In_3550,In_3551,In_3552,In_3553,In_3554,In_3555,In_3556,In_3557,In_3558,In_3559,In_3560,In_3561,In_3562,In_3563,In_3564,In_3565,In_3566,In_3567,In_3568,In_3569,In_3570,In_3571,In_3572,In_3573,In_3574,In_3575,In_3576,In_3577,In_3578,In_3579,In_3580,In_3581,In_3582,In_3583,In_3584,In_3585,In_3586,In_3587,In_3588,In_3589,In_3590,In_3591,In_3592,In_3593,In_3594,In_3595,In_3596,In_3597,In_3598,In_3599,In_3600,In_3601,In_3602,In_3603,In_3604,In_3605,In_3606,In_3607,In_3608,In_3609,In_3610,In_3611,In_3612,In_3613,In_3614,In_3615,In_3616,In_3617,In_3618,In_3619,In_3620,In_3621,In_3622,In_3623,In_3624,In_3625,In_3626,In_3627,In_3628,In_3629,In_3630,In_3631,In_3632,In_3633,In_3634,In_3635,In_3636,In_3637,In_3638,In_3639,In_3640,In_3641,In_3642,In_3643,In_3644,In_3645,In_3646,In_3647,In_3648,In_3649,In_3650,In_3651,In_3652,In_3653,In_3654,In_3655,In_3656,In_3657,In_3658,In_3659,In_3660,In_3661,In_3662,In_3663,In_3664,In_3665,In_3666,In_3667,In_3668,In_3669,In_3670,In_3671,In_3672,In_3673,In_3674,In_3675,In_3676,In_3677,In_3678,In_3679,In_3680,In_3681,In_3682,In_3683,In_3684,In_3685,In_3686,In_3687,In_3688,In_3689,In_3690,In_3691,In_3692,In_3693,In_3694,In_3695,In_3696,In_3697,In_3698,In_3699,In_3700,In_3701,In_3702,In_3703,In_3704,In_3705,In_3706,In_3707,In_3708,In_3709,In_3710,In_3711,In_3712,In_3713,In_3714,In_3715,In_3716,In_3717,In_3718,In_3719,In_3720,In_3721,In_3722,In_3723,In_3724,In_3725,In_3726,In_3727,In_3728,In_3729,In_3730,In_3731,In_3732,In_3733,In_3734,In_3735,In_3736,In_3737,In_3738,In_3739,In_3740,In_3741,In_3742,In_3743,In_3744,In_3745,In_3746,In_3747,In_3748,In_3749,In_3750,In_3751,In_3752,In_3753,In_3754,In_3755,In_3756,In_3757,In_3758,In_3759,In_3760,In_3761,In_3762,In_3763,In_3764,In_3765,In_3766,In_3767,In_3768,In_3769,In_3770,In_3771,In_3772,In_3773,In_3774,In_3775,In_3776,In_3777,In_3778,In_3779,In_3780,In_3781,In_3782,In_3783,In_3784,In_3785,In_3786,In_3787,In_3788,In_3789,In_3790,In_3791,In_3792,In_3793,In_3794,In_3795,In_3796,In_3797,In_3798,In_3799,In_3800,In_3801,In_3802,In_3803,In_3804,In_3805,In_3806,In_3807,In_3808,In_3809,In_3810,In_3811,In_3812,In_3813,In_3814,In_3815,In_3816,In_3817,In_3818,In_3819,In_3820,In_3821,In_3822,In_3823,In_3824,In_3825,In_3826,In_3827,In_3828,In_3829,In_3830,In_3831,In_3832,In_3833,In_3834,In_3835,In_3836,In_3837,In_3838,In_3839,In_3840,In_3841,In_3842,In_3843,In_3844,In_3845,In_3846,In_3847,In_3848,In_3849,In_3850,In_3851,In_3852,In_3853,In_3854,In_3855,In_3856,In_3857,In_3858,In_3859,In_3860,In_3861,In_3862,In_3863,In_3864,In_3865,In_3866,In_3867,In_3868,In_3869,In_3870,In_3871,In_3872,In_3873,In_3874,In_3875,In_3876,In_3877,In_3878,In_3879,In_3880,In_3881,In_3882,In_3883,In_3884,In_3885,In_3886,In_3887,In_3888,In_3889,In_3890,In_3891,In_3892,In_3893,In_3894,In_3895,In_3896,In_3897,In_3898,In_3899,In_3900,In_3901,In_3902,In_3903,In_3904,In_3905,In_3906,In_3907,In_3908,In_3909,In_3910,In_3911,In_3912,In_3913,In_3914,In_3915,In_3916,In_3917,In_3918,In_3919,In_3920,In_3921,In_3922,In_3923,In_3924,In_3925,In_3926,In_3927,In_3928,In_3929,In_3930,In_3931,In_3932,In_3933,In_3934,In_3935,In_3936,In_3937,In_3938,In_3939,In_3940,In_3941,In_3942,In_3943,In_3944,In_3945,In_3946,In_3947,In_3948,In_3949,In_3950,In_3951,In_3952,In_3953,In_3954,In_3955,In_3956,In_3957,In_3958,In_3959,In_3960,In_3961,In_3962,In_3963,In_3964,In_3965,In_3966,In_3967,In_3968,In_3969,In_3970,In_3971,In_3972,In_3973,In_3974,In_3975,In_3976,In_3977,In_3978,In_3979,In_3980,In_3981,In_3982,In_3983,In_3984,In_3985,In_3986,In_3987,In_3988,In_3989,In_3990,In_3991,In_3992,In_3993,In_3994,In_3995,In_3996,In_3997,In_3998,In_3999,In_4000,In_4001,In_4002,In_4003,In_4004,In_4005,In_4006,In_4007,In_4008,In_4009,In_4010,In_4011,In_4012,In_4013,In_4014,In_4015,In_4016,In_4017,In_4018,In_4019,In_4020,In_4021,In_4022,In_4023,In_4024,In_4025,In_4026,In_4027,In_4028,In_4029,In_4030,In_4031,In_4032,In_4033,In_4034,In_4035,In_4036,In_4037,In_4038,In_4039,In_4040,In_4041,In_4042,In_4043,In_4044,In_4045,In_4046,In_4047,In_4048,In_4049,In_4050,In_4051,In_4052,In_4053,In_4054,In_4055,In_4056,In_4057,In_4058,In_4059,In_4060,In_4061,In_4062,In_4063,In_4064,In_4065,In_4066,In_4067,In_4068,In_4069,In_4070,In_4071,In_4072,In_4073,In_4074,In_4075,In_4076,In_4077,In_4078,In_4079,In_4080,In_4081,In_4082,In_4083,In_4084,In_4085,In_4086,In_4087,In_4088,In_4089,In_4090,In_4091,In_4092,In_4093,In_4094,In_4095,In_4096,In_4097,In_4098,In_4099,In_4100,In_4101,In_4102,In_4103,In_4104,In_4105,In_4106,In_4107,In_4108,In_4109,In_4110,In_4111,In_4112,In_4113,In_4114,In_4115,In_4116,In_4117,In_4118,In_4119,In_4120,In_4121,In_4122,In_4123,In_4124,In_4125,In_4126,In_4127,In_4128,In_4129,In_4130,In_4131,In_4132,In_4133,In_4134,In_4135,In_4136,In_4137,In_4138,In_4139,In_4140,In_4141,In_4142,In_4143,In_4144,In_4145,In_4146,In_4147,In_4148,In_4149,In_4150,In_4151,In_4152,In_4153,In_4154,In_4155,In_4156,In_4157,In_4158,In_4159,In_4160,In_4161,In_4162,In_4163,In_4164,In_4165,In_4166,In_4167,In_4168,In_4169,In_4170,In_4171,In_4172,In_4173,In_4174,In_4175,In_4176,In_4177,In_4178,In_4179,In_4180,In_4181,In_4182,In_4183,In_4184,In_4185,In_4186,In_4187,In_4188,In_4189,In_4190,In_4191,In_4192,In_4193,In_4194,In_4195,In_4196,In_4197,In_4198,In_4199,In_4200,In_4201,In_4202,In_4203,In_4204,In_4205,In_4206,In_4207,In_4208,In_4209,In_4210,In_4211,In_4212,In_4213,In_4214,In_4215,In_4216,In_4217,In_4218,In_4219,In_4220,In_4221,In_4222,In_4223,In_4224,In_4225,In_4226,In_4227,In_4228,In_4229,In_4230,In_4231,In_4232,In_4233,In_4234,In_4235,In_4236,In_4237,In_4238,In_4239,In_4240,In_4241,In_4242,In_4243,In_4244,In_4245,In_4246,In_4247,In_4248,In_4249,In_4250,In_4251,In_4252,In_4253,In_4254,In_4255,In_4256,In_4257,In_4258,In_4259,In_4260,In_4261,In_4262,In_4263,In_4264,In_4265,In_4266,In_4267,In_4268,In_4269,In_4270,In_4271,In_4272,In_4273,In_4274,In_4275,In_4276,In_4277,In_4278,In_4279,In_4280,In_4281,In_4282,In_4283,In_4284,In_4285,In_4286,In_4287,In_4288,In_4289,In_4290,In_4291,In_4292,In_4293,In_4294,In_4295,In_4296,In_4297,In_4298,In_4299,In_4300,In_4301,In_4302,In_4303,In_4304,In_4305,In_4306,In_4307,In_4308,In_4309,In_4310,In_4311,In_4312,In_4313,In_4314,In_4315,In_4316,In_4317,In_4318,In_4319,In_4320,In_4321,In_4322,In_4323,In_4324,In_4325,In_4326,In_4327,In_4328,In_4329,In_4330,In_4331,In_4332,In_4333,In_4334,In_4335,In_4336,In_4337,In_4338,In_4339,In_4340,In_4341,In_4342,In_4343,In_4344,In_4345,In_4346,In_4347,In_4348,In_4349,In_4350,In_4351,In_4352,In_4353,In_4354,In_4355,In_4356,In_4357,In_4358,In_4359,In_4360,In_4361,In_4362,In_4363,In_4364,In_4365,In_4366,In_4367,In_4368,In_4369,In_4370,In_4371,In_4372,In_4373,In_4374,In_4375,In_4376,In_4377,In_4378,In_4379,In_4380,In_4381,In_4382,In_4383,In_4384,In_4385,In_4386,In_4387,In_4388,In_4389,In_4390,In_4391,In_4392,In_4393,In_4394,In_4395,In_4396,In_4397,In_4398,In_4399,In_4400,In_4401,In_4402,In_4403,In_4404,In_4405,In_4406,In_4407,In_4408,In_4409,In_4410,In_4411,In_4412,In_4413,In_4414,In_4415,In_4416,In_4417,In_4418,In_4419,In_4420,In_4421,In_4422,In_4423,In_4424,In_4425,In_4426,In_4427,In_4428,In_4429,In_4430,In_4431,In_4432,In_4433,In_4434,In_4435,In_4436,In_4437,In_4438,In_4439,In_4440,In_4441,In_4442,In_4443,In_4444,In_4445,In_4446,In_4447,In_4448,In_4449,In_4450,In_4451,In_4452,In_4453,In_4454,In_4455,In_4456,In_4457,In_4458,In_4459,In_4460,In_4461,In_4462,In_4463,In_4464,In_4465,In_4466,In_4467,In_4468,In_4469,In_4470,In_4471,In_4472,In_4473,In_4474,In_4475,In_4476,In_4477,In_4478,In_4479,In_4480,In_4481,In_4482,In_4483,In_4484,In_4485,In_4486,In_4487,In_4488,In_4489,In_4490,In_4491,In_4492,In_4493,In_4494,In_4495,In_4496,In_4497,In_4498,In_4499,In_4500,In_4501,In_4502,In_4503,In_4504,In_4505,In_4506,In_4507,In_4508,In_4509,In_4510,In_4511,In_4512,In_4513,In_4514,In_4515,In_4516,In_4517,In_4518,In_4519,In_4520,In_4521,In_4522,In_4523,In_4524,In_4525,In_4526,In_4527,In_4528,In_4529,In_4530,In_4531,In_4532,In_4533,In_4534,In_4535,In_4536,In_4537,In_4538,In_4539,In_4540,In_4541,In_4542,In_4543,In_4544,In_4545,In_4546,In_4547,In_4548,In_4549,In_4550,In_4551,In_4552,In_4553,In_4554,In_4555,In_4556,In_4557,In_4558,In_4559,In_4560,In_4561,In_4562,In_4563,In_4564,In_4565,In_4566,In_4567,In_4568,In_4569,In_4570,In_4571,In_4572,In_4573,In_4574,In_4575,In_4576,In_4577,In_4578,In_4579,In_4580,In_4581,In_4582,In_4583,In_4584,In_4585,In_4586,In_4587,In_4588,In_4589,In_4590,In_4591,In_4592,In_4593,In_4594,In_4595,In_4596,In_4597,In_4598,In_4599,In_4600,In_4601,In_4602,In_4603,In_4604,In_4605,In_4606,In_4607,In_4608,In_4609,In_4610,In_4611,In_4612,In_4613,In_4614,In_4615,In_4616,In_4617,In_4618,In_4619,In_4620,In_4621,In_4622,In_4623,In_4624,In_4625,In_4626,In_4627,In_4628,In_4629,In_4630,In_4631,In_4632,In_4633,In_4634,In_4635,In_4636,In_4637,In_4638,In_4639,In_4640,In_4641,In_4642,In_4643,In_4644,In_4645,In_4646,In_4647,In_4648,In_4649,In_4650,In_4651,In_4652,In_4653,In_4654,In_4655,In_4656,In_4657,In_4658,In_4659,In_4660,In_4661,In_4662,In_4663,In_4664,In_4665,In_4666,In_4667,In_4668,In_4669,In_4670,In_4671,In_4672,In_4673,In_4674,In_4675,In_4676,In_4677,In_4678,In_4679,In_4680,In_4681,In_4682,In_4683,In_4684,In_4685,In_4686,In_4687,In_4688,In_4689,In_4690,In_4691,In_4692,In_4693,In_4694,In_4695,In_4696,In_4697,In_4698,In_4699,In_4700,In_4701,In_4702,In_4703,In_4704,In_4705,In_4706,In_4707,In_4708,In_4709,In_4710,In_4711,In_4712,In_4713,In_4714,In_4715,In_4716,In_4717,In_4718,In_4719,In_4720,In_4721,In_4722,In_4723,In_4724,In_4725,In_4726,In_4727,In_4728,In_4729,In_4730,In_4731,In_4732,In_4733,In_4734,In_4735,In_4736,In_4737,In_4738,In_4739,In_4740,In_4741,In_4742,In_4743,In_4744,In_4745,In_4746,In_4747,In_4748,In_4749,In_4750,In_4751,In_4752,In_4753,In_4754,In_4755,In_4756,In_4757,In_4758,In_4759,In_4760,In_4761,In_4762,In_4763,In_4764,In_4765,In_4766,In_4767,In_4768,In_4769,In_4770,In_4771,In_4772,In_4773,In_4774,In_4775,In_4776,In_4777,In_4778,In_4779,In_4780,In_4781,In_4782,In_4783,In_4784,In_4785,In_4786,In_4787,In_4788,In_4789,In_4790,In_4791,In_4792,In_4793,In_4794,In_4795,In_4796,In_4797,In_4798,In_4799,In_4800,In_4801,In_4802,In_4803,In_4804,In_4805,In_4806,In_4807,In_4808,In_4809,In_4810,In_4811,In_4812,In_4813,In_4814,In_4815,In_4816,In_4817,In_4818,In_4819,In_4820,In_4821,In_4822,In_4823,In_4824,In_4825,In_4826,In_4827,In_4828,In_4829,In_4830,In_4831,In_4832,In_4833,In_4834,In_4835,In_4836,In_4837,In_4838,In_4839,In_4840,In_4841,In_4842,In_4843,In_4844,In_4845,In_4846,In_4847,In_4848,In_4849,In_4850,In_4851,In_4852,In_4853,In_4854,In_4855,In_4856,In_4857,In_4858,In_4859,In_4860,In_4861,In_4862,In_4863,In_4864,In_4865,In_4866,In_4867,In_4868,In_4869,In_4870,In_4871,In_4872,In_4873,In_4874,In_4875,In_4876,In_4877,In_4878,In_4879,In_4880,In_4881,In_4882,In_4883,In_4884,In_4885,In_4886,In_4887,In_4888,In_4889,In_4890,In_4891,In_4892,In_4893,In_4894,In_4895,In_4896,In_4897,In_4898,In_4899,In_4900,In_4901,In_4902,In_4903,In_4904,In_4905,In_4906,In_4907,In_4908,In_4909,In_4910,In_4911,In_4912,In_4913,In_4914,In_4915,In_4916,In_4917,In_4918,In_4919,In_4920,In_4921,In_4922,In_4923,In_4924,In_4925,In_4926,In_4927,In_4928,In_4929,In_4930,In_4931,In_4932,In_4933,In_4934,In_4935,In_4936,In_4937,In_4938,In_4939,In_4940,In_4941,In_4942,In_4943,In_4944,In_4945,In_4946,In_4947,In_4948,In_4949,In_4950,In_4951,In_4952,In_4953,In_4954,In_4955,In_4956,In_4957,In_4958,In_4959,In_4960,In_4961,In_4962,In_4963,In_4964,In_4965,In_4966,In_4967,In_4968,In_4969,In_4970,In_4971,In_4972,In_4973,In_4974,In_4975,In_4976,In_4977,In_4978,In_4979,In_4980,In_4981,In_4982,In_4983,In_4984,In_4985,In_4986,In_4987,In_4988,In_4989,In_4990,In_4991,In_4992,In_4993,In_4994,In_4995,In_4996,In_4997,In_4998,In_4999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499,O_3500,O_3501,O_3502,O_3503,O_3504,O_3505,O_3506,O_3507,O_3508,O_3509,O_3510,O_3511,O_3512,O_3513,O_3514,O_3515,O_3516,O_3517,O_3518,O_3519,O_3520,O_3521,O_3522,O_3523,O_3524,O_3525,O_3526,O_3527,O_3528,O_3529,O_3530,O_3531,O_3532,O_3533,O_3534,O_3535,O_3536,O_3537,O_3538,O_3539,O_3540,O_3541,O_3542,O_3543,O_3544,O_3545,O_3546,O_3547,O_3548,O_3549,O_3550,O_3551,O_3552,O_3553,O_3554,O_3555,O_3556,O_3557,O_3558,O_3559,O_3560,O_3561,O_3562,O_3563,O_3564,O_3565,O_3566,O_3567,O_3568,O_3569,O_3570,O_3571,O_3572,O_3573,O_3574,O_3575,O_3576,O_3577,O_3578,O_3579,O_3580,O_3581,O_3582,O_3583,O_3584,O_3585,O_3586,O_3587,O_3588,O_3589,O_3590,O_3591,O_3592,O_3593,O_3594,O_3595,O_3596,O_3597,O_3598,O_3599,O_3600,O_3601,O_3602,O_3603,O_3604,O_3605,O_3606,O_3607,O_3608,O_3609,O_3610,O_3611,O_3612,O_3613,O_3614,O_3615,O_3616,O_3617,O_3618,O_3619,O_3620,O_3621,O_3622,O_3623,O_3624,O_3625,O_3626,O_3627,O_3628,O_3629,O_3630,O_3631,O_3632,O_3633,O_3634,O_3635,O_3636,O_3637,O_3638,O_3639,O_3640,O_3641,O_3642,O_3643,O_3644,O_3645,O_3646,O_3647,O_3648,O_3649,O_3650,O_3651,O_3652,O_3653,O_3654,O_3655,O_3656,O_3657,O_3658,O_3659,O_3660,O_3661,O_3662,O_3663,O_3664,O_3665,O_3666,O_3667,O_3668,O_3669,O_3670,O_3671,O_3672,O_3673,O_3674,O_3675,O_3676,O_3677,O_3678,O_3679,O_3680,O_3681,O_3682,O_3683,O_3684,O_3685,O_3686,O_3687,O_3688,O_3689,O_3690,O_3691,O_3692,O_3693,O_3694,O_3695,O_3696,O_3697,O_3698,O_3699,O_3700,O_3701,O_3702,O_3703,O_3704,O_3705,O_3706,O_3707,O_3708,O_3709,O_3710,O_3711,O_3712,O_3713,O_3714,O_3715,O_3716,O_3717,O_3718,O_3719,O_3720,O_3721,O_3722,O_3723,O_3724,O_3725,O_3726,O_3727,O_3728,O_3729,O_3730,O_3731,O_3732,O_3733,O_3734,O_3735,O_3736,O_3737,O_3738,O_3739,O_3740,O_3741,O_3742,O_3743,O_3744,O_3745,O_3746,O_3747,O_3748,O_3749,O_3750,O_3751,O_3752,O_3753,O_3754,O_3755,O_3756,O_3757,O_3758,O_3759,O_3760,O_3761,O_3762,O_3763,O_3764,O_3765,O_3766,O_3767,O_3768,O_3769,O_3770,O_3771,O_3772,O_3773,O_3774,O_3775,O_3776,O_3777,O_3778,O_3779,O_3780,O_3781,O_3782,O_3783,O_3784,O_3785,O_3786,O_3787,O_3788,O_3789,O_3790,O_3791,O_3792,O_3793,O_3794,O_3795,O_3796,O_3797,O_3798,O_3799,O_3800,O_3801,O_3802,O_3803,O_3804,O_3805,O_3806,O_3807,O_3808,O_3809,O_3810,O_3811,O_3812,O_3813,O_3814,O_3815,O_3816,O_3817,O_3818,O_3819,O_3820,O_3821,O_3822,O_3823,O_3824,O_3825,O_3826,O_3827,O_3828,O_3829,O_3830,O_3831,O_3832,O_3833,O_3834,O_3835,O_3836,O_3837,O_3838,O_3839,O_3840,O_3841,O_3842,O_3843,O_3844,O_3845,O_3846,O_3847,O_3848,O_3849,O_3850,O_3851,O_3852,O_3853,O_3854,O_3855,O_3856,O_3857,O_3858,O_3859,O_3860,O_3861,O_3862,O_3863,O_3864,O_3865,O_3866,O_3867,O_3868,O_3869,O_3870,O_3871,O_3872,O_3873,O_3874,O_3875,O_3876,O_3877,O_3878,O_3879,O_3880,O_3881,O_3882,O_3883,O_3884,O_3885,O_3886,O_3887,O_3888,O_3889,O_3890,O_3891,O_3892,O_3893,O_3894,O_3895,O_3896,O_3897,O_3898,O_3899,O_3900,O_3901,O_3902,O_3903,O_3904,O_3905,O_3906,O_3907,O_3908,O_3909,O_3910,O_3911,O_3912,O_3913,O_3914,O_3915,O_3916,O_3917,O_3918,O_3919,O_3920,O_3921,O_3922,O_3923,O_3924,O_3925,O_3926,O_3927,O_3928,O_3929,O_3930,O_3931,O_3932,O_3933,O_3934,O_3935,O_3936,O_3937,O_3938,O_3939,O_3940,O_3941,O_3942,O_3943,O_3944,O_3945,O_3946,O_3947,O_3948,O_3949,O_3950,O_3951,O_3952,O_3953,O_3954,O_3955,O_3956,O_3957,O_3958,O_3959,O_3960,O_3961,O_3962,O_3963,O_3964,O_3965,O_3966,O_3967,O_3968,O_3969,O_3970,O_3971,O_3972,O_3973,O_3974,O_3975,O_3976,O_3977,O_3978,O_3979,O_3980,O_3981,O_3982,O_3983,O_3984,O_3985,O_3986,O_3987,O_3988,O_3989,O_3990,O_3991,O_3992,O_3993,O_3994,O_3995,O_3996,O_3997,O_3998,O_3999,O_4000,O_4001,O_4002,O_4003,O_4004,O_4005,O_4006,O_4007,O_4008,O_4009,O_4010,O_4011,O_4012,O_4013,O_4014,O_4015,O_4016,O_4017,O_4018,O_4019,O_4020,O_4021,O_4022,O_4023,O_4024,O_4025,O_4026,O_4027,O_4028,O_4029,O_4030,O_4031,O_4032,O_4033,O_4034,O_4035,O_4036,O_4037,O_4038,O_4039,O_4040,O_4041,O_4042,O_4043,O_4044,O_4045,O_4046,O_4047,O_4048,O_4049,O_4050,O_4051,O_4052,O_4053,O_4054,O_4055,O_4056,O_4057,O_4058,O_4059,O_4060,O_4061,O_4062,O_4063,O_4064,O_4065,O_4066,O_4067,O_4068,O_4069,O_4070,O_4071,O_4072,O_4073,O_4074,O_4075,O_4076,O_4077,O_4078,O_4079,O_4080,O_4081,O_4082,O_4083,O_4084,O_4085,O_4086,O_4087,O_4088,O_4089,O_4090,O_4091,O_4092,O_4093,O_4094,O_4095,O_4096,O_4097,O_4098,O_4099,O_4100,O_4101,O_4102,O_4103,O_4104,O_4105,O_4106,O_4107,O_4108,O_4109,O_4110,O_4111,O_4112,O_4113,O_4114,O_4115,O_4116,O_4117,O_4118,O_4119,O_4120,O_4121,O_4122,O_4123,O_4124,O_4125,O_4126,O_4127,O_4128,O_4129,O_4130,O_4131,O_4132,O_4133,O_4134,O_4135,O_4136,O_4137,O_4138,O_4139,O_4140,O_4141,O_4142,O_4143,O_4144,O_4145,O_4146,O_4147,O_4148,O_4149,O_4150,O_4151,O_4152,O_4153,O_4154,O_4155,O_4156,O_4157,O_4158,O_4159,O_4160,O_4161,O_4162,O_4163,O_4164,O_4165,O_4166,O_4167,O_4168,O_4169,O_4170,O_4171,O_4172,O_4173,O_4174,O_4175,O_4176,O_4177,O_4178,O_4179,O_4180,O_4181,O_4182,O_4183,O_4184,O_4185,O_4186,O_4187,O_4188,O_4189,O_4190,O_4191,O_4192,O_4193,O_4194,O_4195,O_4196,O_4197,O_4198,O_4199,O_4200,O_4201,O_4202,O_4203,O_4204,O_4205,O_4206,O_4207,O_4208,O_4209,O_4210,O_4211,O_4212,O_4213,O_4214,O_4215,O_4216,O_4217,O_4218,O_4219,O_4220,O_4221,O_4222,O_4223,O_4224,O_4225,O_4226,O_4227,O_4228,O_4229,O_4230,O_4231,O_4232,O_4233,O_4234,O_4235,O_4236,O_4237,O_4238,O_4239,O_4240,O_4241,O_4242,O_4243,O_4244,O_4245,O_4246,O_4247,O_4248,O_4249,O_4250,O_4251,O_4252,O_4253,O_4254,O_4255,O_4256,O_4257,O_4258,O_4259,O_4260,O_4261,O_4262,O_4263,O_4264,O_4265,O_4266,O_4267,O_4268,O_4269,O_4270,O_4271,O_4272,O_4273,O_4274,O_4275,O_4276,O_4277,O_4278,O_4279,O_4280,O_4281,O_4282,O_4283,O_4284,O_4285,O_4286,O_4287,O_4288,O_4289,O_4290,O_4291,O_4292,O_4293,O_4294,O_4295,O_4296,O_4297,O_4298,O_4299,O_4300,O_4301,O_4302,O_4303,O_4304,O_4305,O_4306,O_4307,O_4308,O_4309,O_4310,O_4311,O_4312,O_4313,O_4314,O_4315,O_4316,O_4317,O_4318,O_4319,O_4320,O_4321,O_4322,O_4323,O_4324,O_4325,O_4326,O_4327,O_4328,O_4329,O_4330,O_4331,O_4332,O_4333,O_4334,O_4335,O_4336,O_4337,O_4338,O_4339,O_4340,O_4341,O_4342,O_4343,O_4344,O_4345,O_4346,O_4347,O_4348,O_4349,O_4350,O_4351,O_4352,O_4353,O_4354,O_4355,O_4356,O_4357,O_4358,O_4359,O_4360,O_4361,O_4362,O_4363,O_4364,O_4365,O_4366,O_4367,O_4368,O_4369,O_4370,O_4371,O_4372,O_4373,O_4374,O_4375,O_4376,O_4377,O_4378,O_4379,O_4380,O_4381,O_4382,O_4383,O_4384,O_4385,O_4386,O_4387,O_4388,O_4389,O_4390,O_4391,O_4392,O_4393,O_4394,O_4395,O_4396,O_4397,O_4398,O_4399,O_4400,O_4401,O_4402,O_4403,O_4404,O_4405,O_4406,O_4407,O_4408,O_4409,O_4410,O_4411,O_4412,O_4413,O_4414,O_4415,O_4416,O_4417,O_4418,O_4419,O_4420,O_4421,O_4422,O_4423,O_4424,O_4425,O_4426,O_4427,O_4428,O_4429,O_4430,O_4431,O_4432,O_4433,O_4434,O_4435,O_4436,O_4437,O_4438,O_4439,O_4440,O_4441,O_4442,O_4443,O_4444,O_4445,O_4446,O_4447,O_4448,O_4449,O_4450,O_4451,O_4452,O_4453,O_4454,O_4455,O_4456,O_4457,O_4458,O_4459,O_4460,O_4461,O_4462,O_4463,O_4464,O_4465,O_4466,O_4467,O_4468,O_4469,O_4470,O_4471,O_4472,O_4473,O_4474,O_4475,O_4476,O_4477,O_4478,O_4479,O_4480,O_4481,O_4482,O_4483,O_4484,O_4485,O_4486,O_4487,O_4488,O_4489,O_4490,O_4491,O_4492,O_4493,O_4494,O_4495,O_4496,O_4497,O_4498,O_4499,O_4500,O_4501,O_4502,O_4503,O_4504,O_4505,O_4506,O_4507,O_4508,O_4509,O_4510,O_4511,O_4512,O_4513,O_4514,O_4515,O_4516,O_4517,O_4518,O_4519,O_4520,O_4521,O_4522,O_4523,O_4524,O_4525,O_4526,O_4527,O_4528,O_4529,O_4530,O_4531,O_4532,O_4533,O_4534,O_4535,O_4536,O_4537,O_4538,O_4539,O_4540,O_4541,O_4542,O_4543,O_4544,O_4545,O_4546,O_4547,O_4548,O_4549,O_4550,O_4551,O_4552,O_4553,O_4554,O_4555,O_4556,O_4557,O_4558,O_4559,O_4560,O_4561,O_4562,O_4563,O_4564,O_4565,O_4566,O_4567,O_4568,O_4569,O_4570,O_4571,O_4572,O_4573,O_4574,O_4575,O_4576,O_4577,O_4578,O_4579,O_4580,O_4581,O_4582,O_4583,O_4584,O_4585,O_4586,O_4587,O_4588,O_4589,O_4590,O_4591,O_4592,O_4593,O_4594,O_4595,O_4596,O_4597,O_4598,O_4599,O_4600,O_4601,O_4602,O_4603,O_4604,O_4605,O_4606,O_4607,O_4608,O_4609,O_4610,O_4611,O_4612,O_4613,O_4614,O_4615,O_4616,O_4617,O_4618,O_4619,O_4620,O_4621,O_4622,O_4623,O_4624,O_4625,O_4626,O_4627,O_4628,O_4629,O_4630,O_4631,O_4632,O_4633,O_4634,O_4635,O_4636,O_4637,O_4638,O_4639,O_4640,O_4641,O_4642,O_4643,O_4644,O_4645,O_4646,O_4647,O_4648,O_4649,O_4650,O_4651,O_4652,O_4653,O_4654,O_4655,O_4656,O_4657,O_4658,O_4659,O_4660,O_4661,O_4662,O_4663,O_4664,O_4665,O_4666,O_4667,O_4668,O_4669,O_4670,O_4671,O_4672,O_4673,O_4674,O_4675,O_4676,O_4677,O_4678,O_4679,O_4680,O_4681,O_4682,O_4683,O_4684,O_4685,O_4686,O_4687,O_4688,O_4689,O_4690,O_4691,O_4692,O_4693,O_4694,O_4695,O_4696,O_4697,O_4698,O_4699,O_4700,O_4701,O_4702,O_4703,O_4704,O_4705,O_4706,O_4707,O_4708,O_4709,O_4710,O_4711,O_4712,O_4713,O_4714,O_4715,O_4716,O_4717,O_4718,O_4719,O_4720,O_4721,O_4722,O_4723,O_4724,O_4725,O_4726,O_4727,O_4728,O_4729,O_4730,O_4731,O_4732,O_4733,O_4734,O_4735,O_4736,O_4737,O_4738,O_4739,O_4740,O_4741,O_4742,O_4743,O_4744,O_4745,O_4746,O_4747,O_4748,O_4749,O_4750,O_4751,O_4752,O_4753,O_4754,O_4755,O_4756,O_4757,O_4758,O_4759,O_4760,O_4761,O_4762,O_4763,O_4764,O_4765,O_4766,O_4767,O_4768,O_4769,O_4770,O_4771,O_4772,O_4773,O_4774,O_4775,O_4776,O_4777,O_4778,O_4779,O_4780,O_4781,O_4782,O_4783,O_4784,O_4785,O_4786,O_4787,O_4788,O_4789,O_4790,O_4791,O_4792,O_4793,O_4794,O_4795,O_4796,O_4797,O_4798,O_4799,O_4800,O_4801,O_4802,O_4803,O_4804,O_4805,O_4806,O_4807,O_4808,O_4809,O_4810,O_4811,O_4812,O_4813,O_4814,O_4815,O_4816,O_4817,O_4818,O_4819,O_4820,O_4821,O_4822,O_4823,O_4824,O_4825,O_4826,O_4827,O_4828,O_4829,O_4830,O_4831,O_4832,O_4833,O_4834,O_4835,O_4836,O_4837,O_4838,O_4839,O_4840,O_4841,O_4842,O_4843,O_4844,O_4845,O_4846,O_4847,O_4848,O_4849,O_4850,O_4851,O_4852,O_4853,O_4854,O_4855,O_4856,O_4857,O_4858,O_4859,O_4860,O_4861,O_4862,O_4863,O_4864,O_4865,O_4866,O_4867,O_4868,O_4869,O_4870,O_4871,O_4872,O_4873,O_4874,O_4875,O_4876,O_4877,O_4878,O_4879,O_4880,O_4881,O_4882,O_4883,O_4884,O_4885,O_4886,O_4887,O_4888,O_4889,O_4890,O_4891,O_4892,O_4893,O_4894,O_4895,O_4896,O_4897,O_4898,O_4899,O_4900,O_4901,O_4902,O_4903,O_4904,O_4905,O_4906,O_4907,O_4908,O_4909,O_4910,O_4911,O_4912,O_4913,O_4914,O_4915,O_4916,O_4917,O_4918,O_4919,O_4920,O_4921,O_4922,O_4923,O_4924,O_4925,O_4926,O_4927,O_4928,O_4929,O_4930,O_4931,O_4932,O_4933,O_4934,O_4935,O_4936,O_4937,O_4938,O_4939,O_4940,O_4941,O_4942,O_4943,O_4944,O_4945,O_4946,O_4947,O_4948,O_4949,O_4950,O_4951,O_4952,O_4953,O_4954,O_4955,O_4956,O_4957,O_4958,O_4959,O_4960,O_4961,O_4962,O_4963,O_4964,O_4965,O_4966,O_4967,O_4968,O_4969,O_4970,O_4971,O_4972,O_4973,O_4974,O_4975,O_4976,O_4977,O_4978,O_4979,O_4980,O_4981,O_4982,O_4983,O_4984,O_4985,O_4986,O_4987,O_4988,O_4989,O_4990,O_4991,O_4992,O_4993,O_4994,O_4995,O_4996,O_4997,O_4998,O_4999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999,N_25000,N_25001,N_25002,N_25003,N_25004,N_25005,N_25006,N_25007,N_25008,N_25009,N_25010,N_25011,N_25012,N_25013,N_25014,N_25015,N_25016,N_25017,N_25018,N_25019,N_25020,N_25021,N_25022,N_25023,N_25024,N_25025,N_25026,N_25027,N_25028,N_25029,N_25030,N_25031,N_25032,N_25033,N_25034,N_25035,N_25036,N_25037,N_25038,N_25039,N_25040,N_25041,N_25042,N_25043,N_25044,N_25045,N_25046,N_25047,N_25048,N_25049,N_25050,N_25051,N_25052,N_25053,N_25054,N_25055,N_25056,N_25057,N_25058,N_25059,N_25060,N_25061,N_25062,N_25063,N_25064,N_25065,N_25066,N_25067,N_25068,N_25069,N_25070,N_25071,N_25072,N_25073,N_25074,N_25075,N_25076,N_25077,N_25078,N_25079,N_25080,N_25081,N_25082,N_25083,N_25084,N_25085,N_25086,N_25087,N_25088,N_25089,N_25090,N_25091,N_25092,N_25093,N_25094,N_25095,N_25096,N_25097,N_25098,N_25099,N_25100,N_25101,N_25102,N_25103,N_25104,N_25105,N_25106,N_25107,N_25108,N_25109,N_25110,N_25111,N_25112,N_25113,N_25114,N_25115,N_25116,N_25117,N_25118,N_25119,N_25120,N_25121,N_25122,N_25123,N_25124,N_25125,N_25126,N_25127,N_25128,N_25129,N_25130,N_25131,N_25132,N_25133,N_25134,N_25135,N_25136,N_25137,N_25138,N_25139,N_25140,N_25141,N_25142,N_25143,N_25144,N_25145,N_25146,N_25147,N_25148,N_25149,N_25150,N_25151,N_25152,N_25153,N_25154,N_25155,N_25156,N_25157,N_25158,N_25159,N_25160,N_25161,N_25162,N_25163,N_25164,N_25165,N_25166,N_25167,N_25168,N_25169,N_25170,N_25171,N_25172,N_25173,N_25174,N_25175,N_25176,N_25177,N_25178,N_25179,N_25180,N_25181,N_25182,N_25183,N_25184,N_25185,N_25186,N_25187,N_25188,N_25189,N_25190,N_25191,N_25192,N_25193,N_25194,N_25195,N_25196,N_25197,N_25198,N_25199,N_25200,N_25201,N_25202,N_25203,N_25204,N_25205,N_25206,N_25207,N_25208,N_25209,N_25210,N_25211,N_25212,N_25213,N_25214,N_25215,N_25216,N_25217,N_25218,N_25219,N_25220,N_25221,N_25222,N_25223,N_25224,N_25225,N_25226,N_25227,N_25228,N_25229,N_25230,N_25231,N_25232,N_25233,N_25234,N_25235,N_25236,N_25237,N_25238,N_25239,N_25240,N_25241,N_25242,N_25243,N_25244,N_25245,N_25246,N_25247,N_25248,N_25249,N_25250,N_25251,N_25252,N_25253,N_25254,N_25255,N_25256,N_25257,N_25258,N_25259,N_25260,N_25261,N_25262,N_25263,N_25264,N_25265,N_25266,N_25267,N_25268,N_25269,N_25270,N_25271,N_25272,N_25273,N_25274,N_25275,N_25276,N_25277,N_25278,N_25279,N_25280,N_25281,N_25282,N_25283,N_25284,N_25285,N_25286,N_25287,N_25288,N_25289,N_25290,N_25291,N_25292,N_25293,N_25294,N_25295,N_25296,N_25297,N_25298,N_25299,N_25300,N_25301,N_25302,N_25303,N_25304,N_25305,N_25306,N_25307,N_25308,N_25309,N_25310,N_25311,N_25312,N_25313,N_25314,N_25315,N_25316,N_25317,N_25318,N_25319,N_25320,N_25321,N_25322,N_25323,N_25324,N_25325,N_25326,N_25327,N_25328,N_25329,N_25330,N_25331,N_25332,N_25333,N_25334,N_25335,N_25336,N_25337,N_25338,N_25339,N_25340,N_25341,N_25342,N_25343,N_25344,N_25345,N_25346,N_25347,N_25348,N_25349,N_25350,N_25351,N_25352,N_25353,N_25354,N_25355,N_25356,N_25357,N_25358,N_25359,N_25360,N_25361,N_25362,N_25363,N_25364,N_25365,N_25366,N_25367,N_25368,N_25369,N_25370,N_25371,N_25372,N_25373,N_25374,N_25375,N_25376,N_25377,N_25378,N_25379,N_25380,N_25381,N_25382,N_25383,N_25384,N_25385,N_25386,N_25387,N_25388,N_25389,N_25390,N_25391,N_25392,N_25393,N_25394,N_25395,N_25396,N_25397,N_25398,N_25399,N_25400,N_25401,N_25402,N_25403,N_25404,N_25405,N_25406,N_25407,N_25408,N_25409,N_25410,N_25411,N_25412,N_25413,N_25414,N_25415,N_25416,N_25417,N_25418,N_25419,N_25420,N_25421,N_25422,N_25423,N_25424,N_25425,N_25426,N_25427,N_25428,N_25429,N_25430,N_25431,N_25432,N_25433,N_25434,N_25435,N_25436,N_25437,N_25438,N_25439,N_25440,N_25441,N_25442,N_25443,N_25444,N_25445,N_25446,N_25447,N_25448,N_25449,N_25450,N_25451,N_25452,N_25453,N_25454,N_25455,N_25456,N_25457,N_25458,N_25459,N_25460,N_25461,N_25462,N_25463,N_25464,N_25465,N_25466,N_25467,N_25468,N_25469,N_25470,N_25471,N_25472,N_25473,N_25474,N_25475,N_25476,N_25477,N_25478,N_25479,N_25480,N_25481,N_25482,N_25483,N_25484,N_25485,N_25486,N_25487,N_25488,N_25489,N_25490,N_25491,N_25492,N_25493,N_25494,N_25495,N_25496,N_25497,N_25498,N_25499,N_25500,N_25501,N_25502,N_25503,N_25504,N_25505,N_25506,N_25507,N_25508,N_25509,N_25510,N_25511,N_25512,N_25513,N_25514,N_25515,N_25516,N_25517,N_25518,N_25519,N_25520,N_25521,N_25522,N_25523,N_25524,N_25525,N_25526,N_25527,N_25528,N_25529,N_25530,N_25531,N_25532,N_25533,N_25534,N_25535,N_25536,N_25537,N_25538,N_25539,N_25540,N_25541,N_25542,N_25543,N_25544,N_25545,N_25546,N_25547,N_25548,N_25549,N_25550,N_25551,N_25552,N_25553,N_25554,N_25555,N_25556,N_25557,N_25558,N_25559,N_25560,N_25561,N_25562,N_25563,N_25564,N_25565,N_25566,N_25567,N_25568,N_25569,N_25570,N_25571,N_25572,N_25573,N_25574,N_25575,N_25576,N_25577,N_25578,N_25579,N_25580,N_25581,N_25582,N_25583,N_25584,N_25585,N_25586,N_25587,N_25588,N_25589,N_25590,N_25591,N_25592,N_25593,N_25594,N_25595,N_25596,N_25597,N_25598,N_25599,N_25600,N_25601,N_25602,N_25603,N_25604,N_25605,N_25606,N_25607,N_25608,N_25609,N_25610,N_25611,N_25612,N_25613,N_25614,N_25615,N_25616,N_25617,N_25618,N_25619,N_25620,N_25621,N_25622,N_25623,N_25624,N_25625,N_25626,N_25627,N_25628,N_25629,N_25630,N_25631,N_25632,N_25633,N_25634,N_25635,N_25636,N_25637,N_25638,N_25639,N_25640,N_25641,N_25642,N_25643,N_25644,N_25645,N_25646,N_25647,N_25648,N_25649,N_25650,N_25651,N_25652,N_25653,N_25654,N_25655,N_25656,N_25657,N_25658,N_25659,N_25660,N_25661,N_25662,N_25663,N_25664,N_25665,N_25666,N_25667,N_25668,N_25669,N_25670,N_25671,N_25672,N_25673,N_25674,N_25675,N_25676,N_25677,N_25678,N_25679,N_25680,N_25681,N_25682,N_25683,N_25684,N_25685,N_25686,N_25687,N_25688,N_25689,N_25690,N_25691,N_25692,N_25693,N_25694,N_25695,N_25696,N_25697,N_25698,N_25699,N_25700,N_25701,N_25702,N_25703,N_25704,N_25705,N_25706,N_25707,N_25708,N_25709,N_25710,N_25711,N_25712,N_25713,N_25714,N_25715,N_25716,N_25717,N_25718,N_25719,N_25720,N_25721,N_25722,N_25723,N_25724,N_25725,N_25726,N_25727,N_25728,N_25729,N_25730,N_25731,N_25732,N_25733,N_25734,N_25735,N_25736,N_25737,N_25738,N_25739,N_25740,N_25741,N_25742,N_25743,N_25744,N_25745,N_25746,N_25747,N_25748,N_25749,N_25750,N_25751,N_25752,N_25753,N_25754,N_25755,N_25756,N_25757,N_25758,N_25759,N_25760,N_25761,N_25762,N_25763,N_25764,N_25765,N_25766,N_25767,N_25768,N_25769,N_25770,N_25771,N_25772,N_25773,N_25774,N_25775,N_25776,N_25777,N_25778,N_25779,N_25780,N_25781,N_25782,N_25783,N_25784,N_25785,N_25786,N_25787,N_25788,N_25789,N_25790,N_25791,N_25792,N_25793,N_25794,N_25795,N_25796,N_25797,N_25798,N_25799,N_25800,N_25801,N_25802,N_25803,N_25804,N_25805,N_25806,N_25807,N_25808,N_25809,N_25810,N_25811,N_25812,N_25813,N_25814,N_25815,N_25816,N_25817,N_25818,N_25819,N_25820,N_25821,N_25822,N_25823,N_25824,N_25825,N_25826,N_25827,N_25828,N_25829,N_25830,N_25831,N_25832,N_25833,N_25834,N_25835,N_25836,N_25837,N_25838,N_25839,N_25840,N_25841,N_25842,N_25843,N_25844,N_25845,N_25846,N_25847,N_25848,N_25849,N_25850,N_25851,N_25852,N_25853,N_25854,N_25855,N_25856,N_25857,N_25858,N_25859,N_25860,N_25861,N_25862,N_25863,N_25864,N_25865,N_25866,N_25867,N_25868,N_25869,N_25870,N_25871,N_25872,N_25873,N_25874,N_25875,N_25876,N_25877,N_25878,N_25879,N_25880,N_25881,N_25882,N_25883,N_25884,N_25885,N_25886,N_25887,N_25888,N_25889,N_25890,N_25891,N_25892,N_25893,N_25894,N_25895,N_25896,N_25897,N_25898,N_25899,N_25900,N_25901,N_25902,N_25903,N_25904,N_25905,N_25906,N_25907,N_25908,N_25909,N_25910,N_25911,N_25912,N_25913,N_25914,N_25915,N_25916,N_25917,N_25918,N_25919,N_25920,N_25921,N_25922,N_25923,N_25924,N_25925,N_25926,N_25927,N_25928,N_25929,N_25930,N_25931,N_25932,N_25933,N_25934,N_25935,N_25936,N_25937,N_25938,N_25939,N_25940,N_25941,N_25942,N_25943,N_25944,N_25945,N_25946,N_25947,N_25948,N_25949,N_25950,N_25951,N_25952,N_25953,N_25954,N_25955,N_25956,N_25957,N_25958,N_25959,N_25960,N_25961,N_25962,N_25963,N_25964,N_25965,N_25966,N_25967,N_25968,N_25969,N_25970,N_25971,N_25972,N_25973,N_25974,N_25975,N_25976,N_25977,N_25978,N_25979,N_25980,N_25981,N_25982,N_25983,N_25984,N_25985,N_25986,N_25987,N_25988,N_25989,N_25990,N_25991,N_25992,N_25993,N_25994,N_25995,N_25996,N_25997,N_25998,N_25999,N_26000,N_26001,N_26002,N_26003,N_26004,N_26005,N_26006,N_26007,N_26008,N_26009,N_26010,N_26011,N_26012,N_26013,N_26014,N_26015,N_26016,N_26017,N_26018,N_26019,N_26020,N_26021,N_26022,N_26023,N_26024,N_26025,N_26026,N_26027,N_26028,N_26029,N_26030,N_26031,N_26032,N_26033,N_26034,N_26035,N_26036,N_26037,N_26038,N_26039,N_26040,N_26041,N_26042,N_26043,N_26044,N_26045,N_26046,N_26047,N_26048,N_26049,N_26050,N_26051,N_26052,N_26053,N_26054,N_26055,N_26056,N_26057,N_26058,N_26059,N_26060,N_26061,N_26062,N_26063,N_26064,N_26065,N_26066,N_26067,N_26068,N_26069,N_26070,N_26071,N_26072,N_26073,N_26074,N_26075,N_26076,N_26077,N_26078,N_26079,N_26080,N_26081,N_26082,N_26083,N_26084,N_26085,N_26086,N_26087,N_26088,N_26089,N_26090,N_26091,N_26092,N_26093,N_26094,N_26095,N_26096,N_26097,N_26098,N_26099,N_26100,N_26101,N_26102,N_26103,N_26104,N_26105,N_26106,N_26107,N_26108,N_26109,N_26110,N_26111,N_26112,N_26113,N_26114,N_26115,N_26116,N_26117,N_26118,N_26119,N_26120,N_26121,N_26122,N_26123,N_26124,N_26125,N_26126,N_26127,N_26128,N_26129,N_26130,N_26131,N_26132,N_26133,N_26134,N_26135,N_26136,N_26137,N_26138,N_26139,N_26140,N_26141,N_26142,N_26143,N_26144,N_26145,N_26146,N_26147,N_26148,N_26149,N_26150,N_26151,N_26152,N_26153,N_26154,N_26155,N_26156,N_26157,N_26158,N_26159,N_26160,N_26161,N_26162,N_26163,N_26164,N_26165,N_26166,N_26167,N_26168,N_26169,N_26170,N_26171,N_26172,N_26173,N_26174,N_26175,N_26176,N_26177,N_26178,N_26179,N_26180,N_26181,N_26182,N_26183,N_26184,N_26185,N_26186,N_26187,N_26188,N_26189,N_26190,N_26191,N_26192,N_26193,N_26194,N_26195,N_26196,N_26197,N_26198,N_26199,N_26200,N_26201,N_26202,N_26203,N_26204,N_26205,N_26206,N_26207,N_26208,N_26209,N_26210,N_26211,N_26212,N_26213,N_26214,N_26215,N_26216,N_26217,N_26218,N_26219,N_26220,N_26221,N_26222,N_26223,N_26224,N_26225,N_26226,N_26227,N_26228,N_26229,N_26230,N_26231,N_26232,N_26233,N_26234,N_26235,N_26236,N_26237,N_26238,N_26239,N_26240,N_26241,N_26242,N_26243,N_26244,N_26245,N_26246,N_26247,N_26248,N_26249,N_26250,N_26251,N_26252,N_26253,N_26254,N_26255,N_26256,N_26257,N_26258,N_26259,N_26260,N_26261,N_26262,N_26263,N_26264,N_26265,N_26266,N_26267,N_26268,N_26269,N_26270,N_26271,N_26272,N_26273,N_26274,N_26275,N_26276,N_26277,N_26278,N_26279,N_26280,N_26281,N_26282,N_26283,N_26284,N_26285,N_26286,N_26287,N_26288,N_26289,N_26290,N_26291,N_26292,N_26293,N_26294,N_26295,N_26296,N_26297,N_26298,N_26299,N_26300,N_26301,N_26302,N_26303,N_26304,N_26305,N_26306,N_26307,N_26308,N_26309,N_26310,N_26311,N_26312,N_26313,N_26314,N_26315,N_26316,N_26317,N_26318,N_26319,N_26320,N_26321,N_26322,N_26323,N_26324,N_26325,N_26326,N_26327,N_26328,N_26329,N_26330,N_26331,N_26332,N_26333,N_26334,N_26335,N_26336,N_26337,N_26338,N_26339,N_26340,N_26341,N_26342,N_26343,N_26344,N_26345,N_26346,N_26347,N_26348,N_26349,N_26350,N_26351,N_26352,N_26353,N_26354,N_26355,N_26356,N_26357,N_26358,N_26359,N_26360,N_26361,N_26362,N_26363,N_26364,N_26365,N_26366,N_26367,N_26368,N_26369,N_26370,N_26371,N_26372,N_26373,N_26374,N_26375,N_26376,N_26377,N_26378,N_26379,N_26380,N_26381,N_26382,N_26383,N_26384,N_26385,N_26386,N_26387,N_26388,N_26389,N_26390,N_26391,N_26392,N_26393,N_26394,N_26395,N_26396,N_26397,N_26398,N_26399,N_26400,N_26401,N_26402,N_26403,N_26404,N_26405,N_26406,N_26407,N_26408,N_26409,N_26410,N_26411,N_26412,N_26413,N_26414,N_26415,N_26416,N_26417,N_26418,N_26419,N_26420,N_26421,N_26422,N_26423,N_26424,N_26425,N_26426,N_26427,N_26428,N_26429,N_26430,N_26431,N_26432,N_26433,N_26434,N_26435,N_26436,N_26437,N_26438,N_26439,N_26440,N_26441,N_26442,N_26443,N_26444,N_26445,N_26446,N_26447,N_26448,N_26449,N_26450,N_26451,N_26452,N_26453,N_26454,N_26455,N_26456,N_26457,N_26458,N_26459,N_26460,N_26461,N_26462,N_26463,N_26464,N_26465,N_26466,N_26467,N_26468,N_26469,N_26470,N_26471,N_26472,N_26473,N_26474,N_26475,N_26476,N_26477,N_26478,N_26479,N_26480,N_26481,N_26482,N_26483,N_26484,N_26485,N_26486,N_26487,N_26488,N_26489,N_26490,N_26491,N_26492,N_26493,N_26494,N_26495,N_26496,N_26497,N_26498,N_26499,N_26500,N_26501,N_26502,N_26503,N_26504,N_26505,N_26506,N_26507,N_26508,N_26509,N_26510,N_26511,N_26512,N_26513,N_26514,N_26515,N_26516,N_26517,N_26518,N_26519,N_26520,N_26521,N_26522,N_26523,N_26524,N_26525,N_26526,N_26527,N_26528,N_26529,N_26530,N_26531,N_26532,N_26533,N_26534,N_26535,N_26536,N_26537,N_26538,N_26539,N_26540,N_26541,N_26542,N_26543,N_26544,N_26545,N_26546,N_26547,N_26548,N_26549,N_26550,N_26551,N_26552,N_26553,N_26554,N_26555,N_26556,N_26557,N_26558,N_26559,N_26560,N_26561,N_26562,N_26563,N_26564,N_26565,N_26566,N_26567,N_26568,N_26569,N_26570,N_26571,N_26572,N_26573,N_26574,N_26575,N_26576,N_26577,N_26578,N_26579,N_26580,N_26581,N_26582,N_26583,N_26584,N_26585,N_26586,N_26587,N_26588,N_26589,N_26590,N_26591,N_26592,N_26593,N_26594,N_26595,N_26596,N_26597,N_26598,N_26599,N_26600,N_26601,N_26602,N_26603,N_26604,N_26605,N_26606,N_26607,N_26608,N_26609,N_26610,N_26611,N_26612,N_26613,N_26614,N_26615,N_26616,N_26617,N_26618,N_26619,N_26620,N_26621,N_26622,N_26623,N_26624,N_26625,N_26626,N_26627,N_26628,N_26629,N_26630,N_26631,N_26632,N_26633,N_26634,N_26635,N_26636,N_26637,N_26638,N_26639,N_26640,N_26641,N_26642,N_26643,N_26644,N_26645,N_26646,N_26647,N_26648,N_26649,N_26650,N_26651,N_26652,N_26653,N_26654,N_26655,N_26656,N_26657,N_26658,N_26659,N_26660,N_26661,N_26662,N_26663,N_26664,N_26665,N_26666,N_26667,N_26668,N_26669,N_26670,N_26671,N_26672,N_26673,N_26674,N_26675,N_26676,N_26677,N_26678,N_26679,N_26680,N_26681,N_26682,N_26683,N_26684,N_26685,N_26686,N_26687,N_26688,N_26689,N_26690,N_26691,N_26692,N_26693,N_26694,N_26695,N_26696,N_26697,N_26698,N_26699,N_26700,N_26701,N_26702,N_26703,N_26704,N_26705,N_26706,N_26707,N_26708,N_26709,N_26710,N_26711,N_26712,N_26713,N_26714,N_26715,N_26716,N_26717,N_26718,N_26719,N_26720,N_26721,N_26722,N_26723,N_26724,N_26725,N_26726,N_26727,N_26728,N_26729,N_26730,N_26731,N_26732,N_26733,N_26734,N_26735,N_26736,N_26737,N_26738,N_26739,N_26740,N_26741,N_26742,N_26743,N_26744,N_26745,N_26746,N_26747,N_26748,N_26749,N_26750,N_26751,N_26752,N_26753,N_26754,N_26755,N_26756,N_26757,N_26758,N_26759,N_26760,N_26761,N_26762,N_26763,N_26764,N_26765,N_26766,N_26767,N_26768,N_26769,N_26770,N_26771,N_26772,N_26773,N_26774,N_26775,N_26776,N_26777,N_26778,N_26779,N_26780,N_26781,N_26782,N_26783,N_26784,N_26785,N_26786,N_26787,N_26788,N_26789,N_26790,N_26791,N_26792,N_26793,N_26794,N_26795,N_26796,N_26797,N_26798,N_26799,N_26800,N_26801,N_26802,N_26803,N_26804,N_26805,N_26806,N_26807,N_26808,N_26809,N_26810,N_26811,N_26812,N_26813,N_26814,N_26815,N_26816,N_26817,N_26818,N_26819,N_26820,N_26821,N_26822,N_26823,N_26824,N_26825,N_26826,N_26827,N_26828,N_26829,N_26830,N_26831,N_26832,N_26833,N_26834,N_26835,N_26836,N_26837,N_26838,N_26839,N_26840,N_26841,N_26842,N_26843,N_26844,N_26845,N_26846,N_26847,N_26848,N_26849,N_26850,N_26851,N_26852,N_26853,N_26854,N_26855,N_26856,N_26857,N_26858,N_26859,N_26860,N_26861,N_26862,N_26863,N_26864,N_26865,N_26866,N_26867,N_26868,N_26869,N_26870,N_26871,N_26872,N_26873,N_26874,N_26875,N_26876,N_26877,N_26878,N_26879,N_26880,N_26881,N_26882,N_26883,N_26884,N_26885,N_26886,N_26887,N_26888,N_26889,N_26890,N_26891,N_26892,N_26893,N_26894,N_26895,N_26896,N_26897,N_26898,N_26899,N_26900,N_26901,N_26902,N_26903,N_26904,N_26905,N_26906,N_26907,N_26908,N_26909,N_26910,N_26911,N_26912,N_26913,N_26914,N_26915,N_26916,N_26917,N_26918,N_26919,N_26920,N_26921,N_26922,N_26923,N_26924,N_26925,N_26926,N_26927,N_26928,N_26929,N_26930,N_26931,N_26932,N_26933,N_26934,N_26935,N_26936,N_26937,N_26938,N_26939,N_26940,N_26941,N_26942,N_26943,N_26944,N_26945,N_26946,N_26947,N_26948,N_26949,N_26950,N_26951,N_26952,N_26953,N_26954,N_26955,N_26956,N_26957,N_26958,N_26959,N_26960,N_26961,N_26962,N_26963,N_26964,N_26965,N_26966,N_26967,N_26968,N_26969,N_26970,N_26971,N_26972,N_26973,N_26974,N_26975,N_26976,N_26977,N_26978,N_26979,N_26980,N_26981,N_26982,N_26983,N_26984,N_26985,N_26986,N_26987,N_26988,N_26989,N_26990,N_26991,N_26992,N_26993,N_26994,N_26995,N_26996,N_26997,N_26998,N_26999,N_27000,N_27001,N_27002,N_27003,N_27004,N_27005,N_27006,N_27007,N_27008,N_27009,N_27010,N_27011,N_27012,N_27013,N_27014,N_27015,N_27016,N_27017,N_27018,N_27019,N_27020,N_27021,N_27022,N_27023,N_27024,N_27025,N_27026,N_27027,N_27028,N_27029,N_27030,N_27031,N_27032,N_27033,N_27034,N_27035,N_27036,N_27037,N_27038,N_27039,N_27040,N_27041,N_27042,N_27043,N_27044,N_27045,N_27046,N_27047,N_27048,N_27049,N_27050,N_27051,N_27052,N_27053,N_27054,N_27055,N_27056,N_27057,N_27058,N_27059,N_27060,N_27061,N_27062,N_27063,N_27064,N_27065,N_27066,N_27067,N_27068,N_27069,N_27070,N_27071,N_27072,N_27073,N_27074,N_27075,N_27076,N_27077,N_27078,N_27079,N_27080,N_27081,N_27082,N_27083,N_27084,N_27085,N_27086,N_27087,N_27088,N_27089,N_27090,N_27091,N_27092,N_27093,N_27094,N_27095,N_27096,N_27097,N_27098,N_27099,N_27100,N_27101,N_27102,N_27103,N_27104,N_27105,N_27106,N_27107,N_27108,N_27109,N_27110,N_27111,N_27112,N_27113,N_27114,N_27115,N_27116,N_27117,N_27118,N_27119,N_27120,N_27121,N_27122,N_27123,N_27124,N_27125,N_27126,N_27127,N_27128,N_27129,N_27130,N_27131,N_27132,N_27133,N_27134,N_27135,N_27136,N_27137,N_27138,N_27139,N_27140,N_27141,N_27142,N_27143,N_27144,N_27145,N_27146,N_27147,N_27148,N_27149,N_27150,N_27151,N_27152,N_27153,N_27154,N_27155,N_27156,N_27157,N_27158,N_27159,N_27160,N_27161,N_27162,N_27163,N_27164,N_27165,N_27166,N_27167,N_27168,N_27169,N_27170,N_27171,N_27172,N_27173,N_27174,N_27175,N_27176,N_27177,N_27178,N_27179,N_27180,N_27181,N_27182,N_27183,N_27184,N_27185,N_27186,N_27187,N_27188,N_27189,N_27190,N_27191,N_27192,N_27193,N_27194,N_27195,N_27196,N_27197,N_27198,N_27199,N_27200,N_27201,N_27202,N_27203,N_27204,N_27205,N_27206,N_27207,N_27208,N_27209,N_27210,N_27211,N_27212,N_27213,N_27214,N_27215,N_27216,N_27217,N_27218,N_27219,N_27220,N_27221,N_27222,N_27223,N_27224,N_27225,N_27226,N_27227,N_27228,N_27229,N_27230,N_27231,N_27232,N_27233,N_27234,N_27235,N_27236,N_27237,N_27238,N_27239,N_27240,N_27241,N_27242,N_27243,N_27244,N_27245,N_27246,N_27247,N_27248,N_27249,N_27250,N_27251,N_27252,N_27253,N_27254,N_27255,N_27256,N_27257,N_27258,N_27259,N_27260,N_27261,N_27262,N_27263,N_27264,N_27265,N_27266,N_27267,N_27268,N_27269,N_27270,N_27271,N_27272,N_27273,N_27274,N_27275,N_27276,N_27277,N_27278,N_27279,N_27280,N_27281,N_27282,N_27283,N_27284,N_27285,N_27286,N_27287,N_27288,N_27289,N_27290,N_27291,N_27292,N_27293,N_27294,N_27295,N_27296,N_27297,N_27298,N_27299,N_27300,N_27301,N_27302,N_27303,N_27304,N_27305,N_27306,N_27307,N_27308,N_27309,N_27310,N_27311,N_27312,N_27313,N_27314,N_27315,N_27316,N_27317,N_27318,N_27319,N_27320,N_27321,N_27322,N_27323,N_27324,N_27325,N_27326,N_27327,N_27328,N_27329,N_27330,N_27331,N_27332,N_27333,N_27334,N_27335,N_27336,N_27337,N_27338,N_27339,N_27340,N_27341,N_27342,N_27343,N_27344,N_27345,N_27346,N_27347,N_27348,N_27349,N_27350,N_27351,N_27352,N_27353,N_27354,N_27355,N_27356,N_27357,N_27358,N_27359,N_27360,N_27361,N_27362,N_27363,N_27364,N_27365,N_27366,N_27367,N_27368,N_27369,N_27370,N_27371,N_27372,N_27373,N_27374,N_27375,N_27376,N_27377,N_27378,N_27379,N_27380,N_27381,N_27382,N_27383,N_27384,N_27385,N_27386,N_27387,N_27388,N_27389,N_27390,N_27391,N_27392,N_27393,N_27394,N_27395,N_27396,N_27397,N_27398,N_27399,N_27400,N_27401,N_27402,N_27403,N_27404,N_27405,N_27406,N_27407,N_27408,N_27409,N_27410,N_27411,N_27412,N_27413,N_27414,N_27415,N_27416,N_27417,N_27418,N_27419,N_27420,N_27421,N_27422,N_27423,N_27424,N_27425,N_27426,N_27427,N_27428,N_27429,N_27430,N_27431,N_27432,N_27433,N_27434,N_27435,N_27436,N_27437,N_27438,N_27439,N_27440,N_27441,N_27442,N_27443,N_27444,N_27445,N_27446,N_27447,N_27448,N_27449,N_27450,N_27451,N_27452,N_27453,N_27454,N_27455,N_27456,N_27457,N_27458,N_27459,N_27460,N_27461,N_27462,N_27463,N_27464,N_27465,N_27466,N_27467,N_27468,N_27469,N_27470,N_27471,N_27472,N_27473,N_27474,N_27475,N_27476,N_27477,N_27478,N_27479,N_27480,N_27481,N_27482,N_27483,N_27484,N_27485,N_27486,N_27487,N_27488,N_27489,N_27490,N_27491,N_27492,N_27493,N_27494,N_27495,N_27496,N_27497,N_27498,N_27499,N_27500,N_27501,N_27502,N_27503,N_27504,N_27505,N_27506,N_27507,N_27508,N_27509,N_27510,N_27511,N_27512,N_27513,N_27514,N_27515,N_27516,N_27517,N_27518,N_27519,N_27520,N_27521,N_27522,N_27523,N_27524,N_27525,N_27526,N_27527,N_27528,N_27529,N_27530,N_27531,N_27532,N_27533,N_27534,N_27535,N_27536,N_27537,N_27538,N_27539,N_27540,N_27541,N_27542,N_27543,N_27544,N_27545,N_27546,N_27547,N_27548,N_27549,N_27550,N_27551,N_27552,N_27553,N_27554,N_27555,N_27556,N_27557,N_27558,N_27559,N_27560,N_27561,N_27562,N_27563,N_27564,N_27565,N_27566,N_27567,N_27568,N_27569,N_27570,N_27571,N_27572,N_27573,N_27574,N_27575,N_27576,N_27577,N_27578,N_27579,N_27580,N_27581,N_27582,N_27583,N_27584,N_27585,N_27586,N_27587,N_27588,N_27589,N_27590,N_27591,N_27592,N_27593,N_27594,N_27595,N_27596,N_27597,N_27598,N_27599,N_27600,N_27601,N_27602,N_27603,N_27604,N_27605,N_27606,N_27607,N_27608,N_27609,N_27610,N_27611,N_27612,N_27613,N_27614,N_27615,N_27616,N_27617,N_27618,N_27619,N_27620,N_27621,N_27622,N_27623,N_27624,N_27625,N_27626,N_27627,N_27628,N_27629,N_27630,N_27631,N_27632,N_27633,N_27634,N_27635,N_27636,N_27637,N_27638,N_27639,N_27640,N_27641,N_27642,N_27643,N_27644,N_27645,N_27646,N_27647,N_27648,N_27649,N_27650,N_27651,N_27652,N_27653,N_27654,N_27655,N_27656,N_27657,N_27658,N_27659,N_27660,N_27661,N_27662,N_27663,N_27664,N_27665,N_27666,N_27667,N_27668,N_27669,N_27670,N_27671,N_27672,N_27673,N_27674,N_27675,N_27676,N_27677,N_27678,N_27679,N_27680,N_27681,N_27682,N_27683,N_27684,N_27685,N_27686,N_27687,N_27688,N_27689,N_27690,N_27691,N_27692,N_27693,N_27694,N_27695,N_27696,N_27697,N_27698,N_27699,N_27700,N_27701,N_27702,N_27703,N_27704,N_27705,N_27706,N_27707,N_27708,N_27709,N_27710,N_27711,N_27712,N_27713,N_27714,N_27715,N_27716,N_27717,N_27718,N_27719,N_27720,N_27721,N_27722,N_27723,N_27724,N_27725,N_27726,N_27727,N_27728,N_27729,N_27730,N_27731,N_27732,N_27733,N_27734,N_27735,N_27736,N_27737,N_27738,N_27739,N_27740,N_27741,N_27742,N_27743,N_27744,N_27745,N_27746,N_27747,N_27748,N_27749,N_27750,N_27751,N_27752,N_27753,N_27754,N_27755,N_27756,N_27757,N_27758,N_27759,N_27760,N_27761,N_27762,N_27763,N_27764,N_27765,N_27766,N_27767,N_27768,N_27769,N_27770,N_27771,N_27772,N_27773,N_27774,N_27775,N_27776,N_27777,N_27778,N_27779,N_27780,N_27781,N_27782,N_27783,N_27784,N_27785,N_27786,N_27787,N_27788,N_27789,N_27790,N_27791,N_27792,N_27793,N_27794,N_27795,N_27796,N_27797,N_27798,N_27799,N_27800,N_27801,N_27802,N_27803,N_27804,N_27805,N_27806,N_27807,N_27808,N_27809,N_27810,N_27811,N_27812,N_27813,N_27814,N_27815,N_27816,N_27817,N_27818,N_27819,N_27820,N_27821,N_27822,N_27823,N_27824,N_27825,N_27826,N_27827,N_27828,N_27829,N_27830,N_27831,N_27832,N_27833,N_27834,N_27835,N_27836,N_27837,N_27838,N_27839,N_27840,N_27841,N_27842,N_27843,N_27844,N_27845,N_27846,N_27847,N_27848,N_27849,N_27850,N_27851,N_27852,N_27853,N_27854,N_27855,N_27856,N_27857,N_27858,N_27859,N_27860,N_27861,N_27862,N_27863,N_27864,N_27865,N_27866,N_27867,N_27868,N_27869,N_27870,N_27871,N_27872,N_27873,N_27874,N_27875,N_27876,N_27877,N_27878,N_27879,N_27880,N_27881,N_27882,N_27883,N_27884,N_27885,N_27886,N_27887,N_27888,N_27889,N_27890,N_27891,N_27892,N_27893,N_27894,N_27895,N_27896,N_27897,N_27898,N_27899,N_27900,N_27901,N_27902,N_27903,N_27904,N_27905,N_27906,N_27907,N_27908,N_27909,N_27910,N_27911,N_27912,N_27913,N_27914,N_27915,N_27916,N_27917,N_27918,N_27919,N_27920,N_27921,N_27922,N_27923,N_27924,N_27925,N_27926,N_27927,N_27928,N_27929,N_27930,N_27931,N_27932,N_27933,N_27934,N_27935,N_27936,N_27937,N_27938,N_27939,N_27940,N_27941,N_27942,N_27943,N_27944,N_27945,N_27946,N_27947,N_27948,N_27949,N_27950,N_27951,N_27952,N_27953,N_27954,N_27955,N_27956,N_27957,N_27958,N_27959,N_27960,N_27961,N_27962,N_27963,N_27964,N_27965,N_27966,N_27967,N_27968,N_27969,N_27970,N_27971,N_27972,N_27973,N_27974,N_27975,N_27976,N_27977,N_27978,N_27979,N_27980,N_27981,N_27982,N_27983,N_27984,N_27985,N_27986,N_27987,N_27988,N_27989,N_27990,N_27991,N_27992,N_27993,N_27994,N_27995,N_27996,N_27997,N_27998,N_27999,N_28000,N_28001,N_28002,N_28003,N_28004,N_28005,N_28006,N_28007,N_28008,N_28009,N_28010,N_28011,N_28012,N_28013,N_28014,N_28015,N_28016,N_28017,N_28018,N_28019,N_28020,N_28021,N_28022,N_28023,N_28024,N_28025,N_28026,N_28027,N_28028,N_28029,N_28030,N_28031,N_28032,N_28033,N_28034,N_28035,N_28036,N_28037,N_28038,N_28039,N_28040,N_28041,N_28042,N_28043,N_28044,N_28045,N_28046,N_28047,N_28048,N_28049,N_28050,N_28051,N_28052,N_28053,N_28054,N_28055,N_28056,N_28057,N_28058,N_28059,N_28060,N_28061,N_28062,N_28063,N_28064,N_28065,N_28066,N_28067,N_28068,N_28069,N_28070,N_28071,N_28072,N_28073,N_28074,N_28075,N_28076,N_28077,N_28078,N_28079,N_28080,N_28081,N_28082,N_28083,N_28084,N_28085,N_28086,N_28087,N_28088,N_28089,N_28090,N_28091,N_28092,N_28093,N_28094,N_28095,N_28096,N_28097,N_28098,N_28099,N_28100,N_28101,N_28102,N_28103,N_28104,N_28105,N_28106,N_28107,N_28108,N_28109,N_28110,N_28111,N_28112,N_28113,N_28114,N_28115,N_28116,N_28117,N_28118,N_28119,N_28120,N_28121,N_28122,N_28123,N_28124,N_28125,N_28126,N_28127,N_28128,N_28129,N_28130,N_28131,N_28132,N_28133,N_28134,N_28135,N_28136,N_28137,N_28138,N_28139,N_28140,N_28141,N_28142,N_28143,N_28144,N_28145,N_28146,N_28147,N_28148,N_28149,N_28150,N_28151,N_28152,N_28153,N_28154,N_28155,N_28156,N_28157,N_28158,N_28159,N_28160,N_28161,N_28162,N_28163,N_28164,N_28165,N_28166,N_28167,N_28168,N_28169,N_28170,N_28171,N_28172,N_28173,N_28174,N_28175,N_28176,N_28177,N_28178,N_28179,N_28180,N_28181,N_28182,N_28183,N_28184,N_28185,N_28186,N_28187,N_28188,N_28189,N_28190,N_28191,N_28192,N_28193,N_28194,N_28195,N_28196,N_28197,N_28198,N_28199,N_28200,N_28201,N_28202,N_28203,N_28204,N_28205,N_28206,N_28207,N_28208,N_28209,N_28210,N_28211,N_28212,N_28213,N_28214,N_28215,N_28216,N_28217,N_28218,N_28219,N_28220,N_28221,N_28222,N_28223,N_28224,N_28225,N_28226,N_28227,N_28228,N_28229,N_28230,N_28231,N_28232,N_28233,N_28234,N_28235,N_28236,N_28237,N_28238,N_28239,N_28240,N_28241,N_28242,N_28243,N_28244,N_28245,N_28246,N_28247,N_28248,N_28249,N_28250,N_28251,N_28252,N_28253,N_28254,N_28255,N_28256,N_28257,N_28258,N_28259,N_28260,N_28261,N_28262,N_28263,N_28264,N_28265,N_28266,N_28267,N_28268,N_28269,N_28270,N_28271,N_28272,N_28273,N_28274,N_28275,N_28276,N_28277,N_28278,N_28279,N_28280,N_28281,N_28282,N_28283,N_28284,N_28285,N_28286,N_28287,N_28288,N_28289,N_28290,N_28291,N_28292,N_28293,N_28294,N_28295,N_28296,N_28297,N_28298,N_28299,N_28300,N_28301,N_28302,N_28303,N_28304,N_28305,N_28306,N_28307,N_28308,N_28309,N_28310,N_28311,N_28312,N_28313,N_28314,N_28315,N_28316,N_28317,N_28318,N_28319,N_28320,N_28321,N_28322,N_28323,N_28324,N_28325,N_28326,N_28327,N_28328,N_28329,N_28330,N_28331,N_28332,N_28333,N_28334,N_28335,N_28336,N_28337,N_28338,N_28339,N_28340,N_28341,N_28342,N_28343,N_28344,N_28345,N_28346,N_28347,N_28348,N_28349,N_28350,N_28351,N_28352,N_28353,N_28354,N_28355,N_28356,N_28357,N_28358,N_28359,N_28360,N_28361,N_28362,N_28363,N_28364,N_28365,N_28366,N_28367,N_28368,N_28369,N_28370,N_28371,N_28372,N_28373,N_28374,N_28375,N_28376,N_28377,N_28378,N_28379,N_28380,N_28381,N_28382,N_28383,N_28384,N_28385,N_28386,N_28387,N_28388,N_28389,N_28390,N_28391,N_28392,N_28393,N_28394,N_28395,N_28396,N_28397,N_28398,N_28399,N_28400,N_28401,N_28402,N_28403,N_28404,N_28405,N_28406,N_28407,N_28408,N_28409,N_28410,N_28411,N_28412,N_28413,N_28414,N_28415,N_28416,N_28417,N_28418,N_28419,N_28420,N_28421,N_28422,N_28423,N_28424,N_28425,N_28426,N_28427,N_28428,N_28429,N_28430,N_28431,N_28432,N_28433,N_28434,N_28435,N_28436,N_28437,N_28438,N_28439,N_28440,N_28441,N_28442,N_28443,N_28444,N_28445,N_28446,N_28447,N_28448,N_28449,N_28450,N_28451,N_28452,N_28453,N_28454,N_28455,N_28456,N_28457,N_28458,N_28459,N_28460,N_28461,N_28462,N_28463,N_28464,N_28465,N_28466,N_28467,N_28468,N_28469,N_28470,N_28471,N_28472,N_28473,N_28474,N_28475,N_28476,N_28477,N_28478,N_28479,N_28480,N_28481,N_28482,N_28483,N_28484,N_28485,N_28486,N_28487,N_28488,N_28489,N_28490,N_28491,N_28492,N_28493,N_28494,N_28495,N_28496,N_28497,N_28498,N_28499,N_28500,N_28501,N_28502,N_28503,N_28504,N_28505,N_28506,N_28507,N_28508,N_28509,N_28510,N_28511,N_28512,N_28513,N_28514,N_28515,N_28516,N_28517,N_28518,N_28519,N_28520,N_28521,N_28522,N_28523,N_28524,N_28525,N_28526,N_28527,N_28528,N_28529,N_28530,N_28531,N_28532,N_28533,N_28534,N_28535,N_28536,N_28537,N_28538,N_28539,N_28540,N_28541,N_28542,N_28543,N_28544,N_28545,N_28546,N_28547,N_28548,N_28549,N_28550,N_28551,N_28552,N_28553,N_28554,N_28555,N_28556,N_28557,N_28558,N_28559,N_28560,N_28561,N_28562,N_28563,N_28564,N_28565,N_28566,N_28567,N_28568,N_28569,N_28570,N_28571,N_28572,N_28573,N_28574,N_28575,N_28576,N_28577,N_28578,N_28579,N_28580,N_28581,N_28582,N_28583,N_28584,N_28585,N_28586,N_28587,N_28588,N_28589,N_28590,N_28591,N_28592,N_28593,N_28594,N_28595,N_28596,N_28597,N_28598,N_28599,N_28600,N_28601,N_28602,N_28603,N_28604,N_28605,N_28606,N_28607,N_28608,N_28609,N_28610,N_28611,N_28612,N_28613,N_28614,N_28615,N_28616,N_28617,N_28618,N_28619,N_28620,N_28621,N_28622,N_28623,N_28624,N_28625,N_28626,N_28627,N_28628,N_28629,N_28630,N_28631,N_28632,N_28633,N_28634,N_28635,N_28636,N_28637,N_28638,N_28639,N_28640,N_28641,N_28642,N_28643,N_28644,N_28645,N_28646,N_28647,N_28648,N_28649,N_28650,N_28651,N_28652,N_28653,N_28654,N_28655,N_28656,N_28657,N_28658,N_28659,N_28660,N_28661,N_28662,N_28663,N_28664,N_28665,N_28666,N_28667,N_28668,N_28669,N_28670,N_28671,N_28672,N_28673,N_28674,N_28675,N_28676,N_28677,N_28678,N_28679,N_28680,N_28681,N_28682,N_28683,N_28684,N_28685,N_28686,N_28687,N_28688,N_28689,N_28690,N_28691,N_28692,N_28693,N_28694,N_28695,N_28696,N_28697,N_28698,N_28699,N_28700,N_28701,N_28702,N_28703,N_28704,N_28705,N_28706,N_28707,N_28708,N_28709,N_28710,N_28711,N_28712,N_28713,N_28714,N_28715,N_28716,N_28717,N_28718,N_28719,N_28720,N_28721,N_28722,N_28723,N_28724,N_28725,N_28726,N_28727,N_28728,N_28729,N_28730,N_28731,N_28732,N_28733,N_28734,N_28735,N_28736,N_28737,N_28738,N_28739,N_28740,N_28741,N_28742,N_28743,N_28744,N_28745,N_28746,N_28747,N_28748,N_28749,N_28750,N_28751,N_28752,N_28753,N_28754,N_28755,N_28756,N_28757,N_28758,N_28759,N_28760,N_28761,N_28762,N_28763,N_28764,N_28765,N_28766,N_28767,N_28768,N_28769,N_28770,N_28771,N_28772,N_28773,N_28774,N_28775,N_28776,N_28777,N_28778,N_28779,N_28780,N_28781,N_28782,N_28783,N_28784,N_28785,N_28786,N_28787,N_28788,N_28789,N_28790,N_28791,N_28792,N_28793,N_28794,N_28795,N_28796,N_28797,N_28798,N_28799,N_28800,N_28801,N_28802,N_28803,N_28804,N_28805,N_28806,N_28807,N_28808,N_28809,N_28810,N_28811,N_28812,N_28813,N_28814,N_28815,N_28816,N_28817,N_28818,N_28819,N_28820,N_28821,N_28822,N_28823,N_28824,N_28825,N_28826,N_28827,N_28828,N_28829,N_28830,N_28831,N_28832,N_28833,N_28834,N_28835,N_28836,N_28837,N_28838,N_28839,N_28840,N_28841,N_28842,N_28843,N_28844,N_28845,N_28846,N_28847,N_28848,N_28849,N_28850,N_28851,N_28852,N_28853,N_28854,N_28855,N_28856,N_28857,N_28858,N_28859,N_28860,N_28861,N_28862,N_28863,N_28864,N_28865,N_28866,N_28867,N_28868,N_28869,N_28870,N_28871,N_28872,N_28873,N_28874,N_28875,N_28876,N_28877,N_28878,N_28879,N_28880,N_28881,N_28882,N_28883,N_28884,N_28885,N_28886,N_28887,N_28888,N_28889,N_28890,N_28891,N_28892,N_28893,N_28894,N_28895,N_28896,N_28897,N_28898,N_28899,N_28900,N_28901,N_28902,N_28903,N_28904,N_28905,N_28906,N_28907,N_28908,N_28909,N_28910,N_28911,N_28912,N_28913,N_28914,N_28915,N_28916,N_28917,N_28918,N_28919,N_28920,N_28921,N_28922,N_28923,N_28924,N_28925,N_28926,N_28927,N_28928,N_28929,N_28930,N_28931,N_28932,N_28933,N_28934,N_28935,N_28936,N_28937,N_28938,N_28939,N_28940,N_28941,N_28942,N_28943,N_28944,N_28945,N_28946,N_28947,N_28948,N_28949,N_28950,N_28951,N_28952,N_28953,N_28954,N_28955,N_28956,N_28957,N_28958,N_28959,N_28960,N_28961,N_28962,N_28963,N_28964,N_28965,N_28966,N_28967,N_28968,N_28969,N_28970,N_28971,N_28972,N_28973,N_28974,N_28975,N_28976,N_28977,N_28978,N_28979,N_28980,N_28981,N_28982,N_28983,N_28984,N_28985,N_28986,N_28987,N_28988,N_28989,N_28990,N_28991,N_28992,N_28993,N_28994,N_28995,N_28996,N_28997,N_28998,N_28999,N_29000,N_29001,N_29002,N_29003,N_29004,N_29005,N_29006,N_29007,N_29008,N_29009,N_29010,N_29011,N_29012,N_29013,N_29014,N_29015,N_29016,N_29017,N_29018,N_29019,N_29020,N_29021,N_29022,N_29023,N_29024,N_29025,N_29026,N_29027,N_29028,N_29029,N_29030,N_29031,N_29032,N_29033,N_29034,N_29035,N_29036,N_29037,N_29038,N_29039,N_29040,N_29041,N_29042,N_29043,N_29044,N_29045,N_29046,N_29047,N_29048,N_29049,N_29050,N_29051,N_29052,N_29053,N_29054,N_29055,N_29056,N_29057,N_29058,N_29059,N_29060,N_29061,N_29062,N_29063,N_29064,N_29065,N_29066,N_29067,N_29068,N_29069,N_29070,N_29071,N_29072,N_29073,N_29074,N_29075,N_29076,N_29077,N_29078,N_29079,N_29080,N_29081,N_29082,N_29083,N_29084,N_29085,N_29086,N_29087,N_29088,N_29089,N_29090,N_29091,N_29092,N_29093,N_29094,N_29095,N_29096,N_29097,N_29098,N_29099,N_29100,N_29101,N_29102,N_29103,N_29104,N_29105,N_29106,N_29107,N_29108,N_29109,N_29110,N_29111,N_29112,N_29113,N_29114,N_29115,N_29116,N_29117,N_29118,N_29119,N_29120,N_29121,N_29122,N_29123,N_29124,N_29125,N_29126,N_29127,N_29128,N_29129,N_29130,N_29131,N_29132,N_29133,N_29134,N_29135,N_29136,N_29137,N_29138,N_29139,N_29140,N_29141,N_29142,N_29143,N_29144,N_29145,N_29146,N_29147,N_29148,N_29149,N_29150,N_29151,N_29152,N_29153,N_29154,N_29155,N_29156,N_29157,N_29158,N_29159,N_29160,N_29161,N_29162,N_29163,N_29164,N_29165,N_29166,N_29167,N_29168,N_29169,N_29170,N_29171,N_29172,N_29173,N_29174,N_29175,N_29176,N_29177,N_29178,N_29179,N_29180,N_29181,N_29182,N_29183,N_29184,N_29185,N_29186,N_29187,N_29188,N_29189,N_29190,N_29191,N_29192,N_29193,N_29194,N_29195,N_29196,N_29197,N_29198,N_29199,N_29200,N_29201,N_29202,N_29203,N_29204,N_29205,N_29206,N_29207,N_29208,N_29209,N_29210,N_29211,N_29212,N_29213,N_29214,N_29215,N_29216,N_29217,N_29218,N_29219,N_29220,N_29221,N_29222,N_29223,N_29224,N_29225,N_29226,N_29227,N_29228,N_29229,N_29230,N_29231,N_29232,N_29233,N_29234,N_29235,N_29236,N_29237,N_29238,N_29239,N_29240,N_29241,N_29242,N_29243,N_29244,N_29245,N_29246,N_29247,N_29248,N_29249,N_29250,N_29251,N_29252,N_29253,N_29254,N_29255,N_29256,N_29257,N_29258,N_29259,N_29260,N_29261,N_29262,N_29263,N_29264,N_29265,N_29266,N_29267,N_29268,N_29269,N_29270,N_29271,N_29272,N_29273,N_29274,N_29275,N_29276,N_29277,N_29278,N_29279,N_29280,N_29281,N_29282,N_29283,N_29284,N_29285,N_29286,N_29287,N_29288,N_29289,N_29290,N_29291,N_29292,N_29293,N_29294,N_29295,N_29296,N_29297,N_29298,N_29299,N_29300,N_29301,N_29302,N_29303,N_29304,N_29305,N_29306,N_29307,N_29308,N_29309,N_29310,N_29311,N_29312,N_29313,N_29314,N_29315,N_29316,N_29317,N_29318,N_29319,N_29320,N_29321,N_29322,N_29323,N_29324,N_29325,N_29326,N_29327,N_29328,N_29329,N_29330,N_29331,N_29332,N_29333,N_29334,N_29335,N_29336,N_29337,N_29338,N_29339,N_29340,N_29341,N_29342,N_29343,N_29344,N_29345,N_29346,N_29347,N_29348,N_29349,N_29350,N_29351,N_29352,N_29353,N_29354,N_29355,N_29356,N_29357,N_29358,N_29359,N_29360,N_29361,N_29362,N_29363,N_29364,N_29365,N_29366,N_29367,N_29368,N_29369,N_29370,N_29371,N_29372,N_29373,N_29374,N_29375,N_29376,N_29377,N_29378,N_29379,N_29380,N_29381,N_29382,N_29383,N_29384,N_29385,N_29386,N_29387,N_29388,N_29389,N_29390,N_29391,N_29392,N_29393,N_29394,N_29395,N_29396,N_29397,N_29398,N_29399,N_29400,N_29401,N_29402,N_29403,N_29404,N_29405,N_29406,N_29407,N_29408,N_29409,N_29410,N_29411,N_29412,N_29413,N_29414,N_29415,N_29416,N_29417,N_29418,N_29419,N_29420,N_29421,N_29422,N_29423,N_29424,N_29425,N_29426,N_29427,N_29428,N_29429,N_29430,N_29431,N_29432,N_29433,N_29434,N_29435,N_29436,N_29437,N_29438,N_29439,N_29440,N_29441,N_29442,N_29443,N_29444,N_29445,N_29446,N_29447,N_29448,N_29449,N_29450,N_29451,N_29452,N_29453,N_29454,N_29455,N_29456,N_29457,N_29458,N_29459,N_29460,N_29461,N_29462,N_29463,N_29464,N_29465,N_29466,N_29467,N_29468,N_29469,N_29470,N_29471,N_29472,N_29473,N_29474,N_29475,N_29476,N_29477,N_29478,N_29479,N_29480,N_29481,N_29482,N_29483,N_29484,N_29485,N_29486,N_29487,N_29488,N_29489,N_29490,N_29491,N_29492,N_29493,N_29494,N_29495,N_29496,N_29497,N_29498,N_29499,N_29500,N_29501,N_29502,N_29503,N_29504,N_29505,N_29506,N_29507,N_29508,N_29509,N_29510,N_29511,N_29512,N_29513,N_29514,N_29515,N_29516,N_29517,N_29518,N_29519,N_29520,N_29521,N_29522,N_29523,N_29524,N_29525,N_29526,N_29527,N_29528,N_29529,N_29530,N_29531,N_29532,N_29533,N_29534,N_29535,N_29536,N_29537,N_29538,N_29539,N_29540,N_29541,N_29542,N_29543,N_29544,N_29545,N_29546,N_29547,N_29548,N_29549,N_29550,N_29551,N_29552,N_29553,N_29554,N_29555,N_29556,N_29557,N_29558,N_29559,N_29560,N_29561,N_29562,N_29563,N_29564,N_29565,N_29566,N_29567,N_29568,N_29569,N_29570,N_29571,N_29572,N_29573,N_29574,N_29575,N_29576,N_29577,N_29578,N_29579,N_29580,N_29581,N_29582,N_29583,N_29584,N_29585,N_29586,N_29587,N_29588,N_29589,N_29590,N_29591,N_29592,N_29593,N_29594,N_29595,N_29596,N_29597,N_29598,N_29599,N_29600,N_29601,N_29602,N_29603,N_29604,N_29605,N_29606,N_29607,N_29608,N_29609,N_29610,N_29611,N_29612,N_29613,N_29614,N_29615,N_29616,N_29617,N_29618,N_29619,N_29620,N_29621,N_29622,N_29623,N_29624,N_29625,N_29626,N_29627,N_29628,N_29629,N_29630,N_29631,N_29632,N_29633,N_29634,N_29635,N_29636,N_29637,N_29638,N_29639,N_29640,N_29641,N_29642,N_29643,N_29644,N_29645,N_29646,N_29647,N_29648,N_29649,N_29650,N_29651,N_29652,N_29653,N_29654,N_29655,N_29656,N_29657,N_29658,N_29659,N_29660,N_29661,N_29662,N_29663,N_29664,N_29665,N_29666,N_29667,N_29668,N_29669,N_29670,N_29671,N_29672,N_29673,N_29674,N_29675,N_29676,N_29677,N_29678,N_29679,N_29680,N_29681,N_29682,N_29683,N_29684,N_29685,N_29686,N_29687,N_29688,N_29689,N_29690,N_29691,N_29692,N_29693,N_29694,N_29695,N_29696,N_29697,N_29698,N_29699,N_29700,N_29701,N_29702,N_29703,N_29704,N_29705,N_29706,N_29707,N_29708,N_29709,N_29710,N_29711,N_29712,N_29713,N_29714,N_29715,N_29716,N_29717,N_29718,N_29719,N_29720,N_29721,N_29722,N_29723,N_29724,N_29725,N_29726,N_29727,N_29728,N_29729,N_29730,N_29731,N_29732,N_29733,N_29734,N_29735,N_29736,N_29737,N_29738,N_29739,N_29740,N_29741,N_29742,N_29743,N_29744,N_29745,N_29746,N_29747,N_29748,N_29749,N_29750,N_29751,N_29752,N_29753,N_29754,N_29755,N_29756,N_29757,N_29758,N_29759,N_29760,N_29761,N_29762,N_29763,N_29764,N_29765,N_29766,N_29767,N_29768,N_29769,N_29770,N_29771,N_29772,N_29773,N_29774,N_29775,N_29776,N_29777,N_29778,N_29779,N_29780,N_29781,N_29782,N_29783,N_29784,N_29785,N_29786,N_29787,N_29788,N_29789,N_29790,N_29791,N_29792,N_29793,N_29794,N_29795,N_29796,N_29797,N_29798,N_29799,N_29800,N_29801,N_29802,N_29803,N_29804,N_29805,N_29806,N_29807,N_29808,N_29809,N_29810,N_29811,N_29812,N_29813,N_29814,N_29815,N_29816,N_29817,N_29818,N_29819,N_29820,N_29821,N_29822,N_29823,N_29824,N_29825,N_29826,N_29827,N_29828,N_29829,N_29830,N_29831,N_29832,N_29833,N_29834,N_29835,N_29836,N_29837,N_29838,N_29839,N_29840,N_29841,N_29842,N_29843,N_29844,N_29845,N_29846,N_29847,N_29848,N_29849,N_29850,N_29851,N_29852,N_29853,N_29854,N_29855,N_29856,N_29857,N_29858,N_29859,N_29860,N_29861,N_29862,N_29863,N_29864,N_29865,N_29866,N_29867,N_29868,N_29869,N_29870,N_29871,N_29872,N_29873,N_29874,N_29875,N_29876,N_29877,N_29878,N_29879,N_29880,N_29881,N_29882,N_29883,N_29884,N_29885,N_29886,N_29887,N_29888,N_29889,N_29890,N_29891,N_29892,N_29893,N_29894,N_29895,N_29896,N_29897,N_29898,N_29899,N_29900,N_29901,N_29902,N_29903,N_29904,N_29905,N_29906,N_29907,N_29908,N_29909,N_29910,N_29911,N_29912,N_29913,N_29914,N_29915,N_29916,N_29917,N_29918,N_29919,N_29920,N_29921,N_29922,N_29923,N_29924,N_29925,N_29926,N_29927,N_29928,N_29929,N_29930,N_29931,N_29932,N_29933,N_29934,N_29935,N_29936,N_29937,N_29938,N_29939,N_29940,N_29941,N_29942,N_29943,N_29944,N_29945,N_29946,N_29947,N_29948,N_29949,N_29950,N_29951,N_29952,N_29953,N_29954,N_29955,N_29956,N_29957,N_29958,N_29959,N_29960,N_29961,N_29962,N_29963,N_29964,N_29965,N_29966,N_29967,N_29968,N_29969,N_29970,N_29971,N_29972,N_29973,N_29974,N_29975,N_29976,N_29977,N_29978,N_29979,N_29980,N_29981,N_29982,N_29983,N_29984,N_29985,N_29986,N_29987,N_29988,N_29989,N_29990,N_29991,N_29992,N_29993,N_29994,N_29995,N_29996,N_29997,N_29998,N_29999,N_30000,N_30001,N_30002,N_30003,N_30004,N_30005,N_30006,N_30007,N_30008,N_30009,N_30010,N_30011,N_30012,N_30013,N_30014,N_30015,N_30016,N_30017,N_30018,N_30019,N_30020,N_30021,N_30022,N_30023,N_30024,N_30025,N_30026,N_30027,N_30028,N_30029,N_30030,N_30031,N_30032,N_30033,N_30034,N_30035,N_30036,N_30037,N_30038,N_30039,N_30040,N_30041,N_30042,N_30043,N_30044,N_30045,N_30046,N_30047,N_30048,N_30049,N_30050,N_30051,N_30052,N_30053,N_30054,N_30055,N_30056,N_30057,N_30058,N_30059,N_30060,N_30061,N_30062,N_30063,N_30064,N_30065,N_30066,N_30067,N_30068,N_30069,N_30070,N_30071,N_30072,N_30073,N_30074,N_30075,N_30076,N_30077,N_30078,N_30079,N_30080,N_30081,N_30082,N_30083,N_30084,N_30085,N_30086,N_30087,N_30088,N_30089,N_30090,N_30091,N_30092,N_30093,N_30094,N_30095,N_30096,N_30097,N_30098,N_30099,N_30100,N_30101,N_30102,N_30103,N_30104,N_30105,N_30106,N_30107,N_30108,N_30109,N_30110,N_30111,N_30112,N_30113,N_30114,N_30115,N_30116,N_30117,N_30118,N_30119,N_30120,N_30121,N_30122,N_30123,N_30124,N_30125,N_30126,N_30127,N_30128,N_30129,N_30130,N_30131,N_30132,N_30133,N_30134,N_30135,N_30136,N_30137,N_30138,N_30139,N_30140,N_30141,N_30142,N_30143,N_30144,N_30145,N_30146,N_30147,N_30148,N_30149,N_30150,N_30151,N_30152,N_30153,N_30154,N_30155,N_30156,N_30157,N_30158,N_30159,N_30160,N_30161,N_30162,N_30163,N_30164,N_30165,N_30166,N_30167,N_30168,N_30169,N_30170,N_30171,N_30172,N_30173,N_30174,N_30175,N_30176,N_30177,N_30178,N_30179,N_30180,N_30181,N_30182,N_30183,N_30184,N_30185,N_30186,N_30187,N_30188,N_30189,N_30190,N_30191,N_30192,N_30193,N_30194,N_30195,N_30196,N_30197,N_30198,N_30199,N_30200,N_30201,N_30202,N_30203,N_30204,N_30205,N_30206,N_30207,N_30208,N_30209,N_30210,N_30211,N_30212,N_30213,N_30214,N_30215,N_30216,N_30217,N_30218,N_30219,N_30220,N_30221,N_30222,N_30223,N_30224,N_30225,N_30226,N_30227,N_30228,N_30229,N_30230,N_30231,N_30232,N_30233,N_30234,N_30235,N_30236,N_30237,N_30238,N_30239,N_30240,N_30241,N_30242,N_30243,N_30244,N_30245,N_30246,N_30247,N_30248,N_30249,N_30250,N_30251,N_30252,N_30253,N_30254,N_30255,N_30256,N_30257,N_30258,N_30259,N_30260,N_30261,N_30262,N_30263,N_30264,N_30265,N_30266,N_30267,N_30268,N_30269,N_30270,N_30271,N_30272,N_30273,N_30274,N_30275,N_30276,N_30277,N_30278,N_30279,N_30280,N_30281,N_30282,N_30283,N_30284,N_30285,N_30286,N_30287,N_30288,N_30289,N_30290,N_30291,N_30292,N_30293,N_30294,N_30295,N_30296,N_30297,N_30298,N_30299,N_30300,N_30301,N_30302,N_30303,N_30304,N_30305,N_30306,N_30307,N_30308,N_30309,N_30310,N_30311,N_30312,N_30313,N_30314,N_30315,N_30316,N_30317,N_30318,N_30319,N_30320,N_30321,N_30322,N_30323,N_30324,N_30325,N_30326,N_30327,N_30328,N_30329,N_30330,N_30331,N_30332,N_30333,N_30334,N_30335,N_30336,N_30337,N_30338,N_30339,N_30340,N_30341,N_30342,N_30343,N_30344,N_30345,N_30346,N_30347,N_30348,N_30349,N_30350,N_30351,N_30352,N_30353,N_30354,N_30355,N_30356,N_30357,N_30358,N_30359,N_30360,N_30361,N_30362,N_30363,N_30364,N_30365,N_30366,N_30367,N_30368,N_30369,N_30370,N_30371,N_30372,N_30373,N_30374,N_30375,N_30376,N_30377,N_30378,N_30379,N_30380,N_30381,N_30382,N_30383,N_30384,N_30385,N_30386,N_30387,N_30388,N_30389,N_30390,N_30391,N_30392,N_30393,N_30394,N_30395,N_30396,N_30397,N_30398,N_30399,N_30400,N_30401,N_30402,N_30403,N_30404,N_30405,N_30406,N_30407,N_30408,N_30409,N_30410,N_30411,N_30412,N_30413,N_30414,N_30415,N_30416,N_30417,N_30418,N_30419,N_30420,N_30421,N_30422,N_30423,N_30424,N_30425,N_30426,N_30427,N_30428,N_30429,N_30430,N_30431,N_30432,N_30433,N_30434,N_30435,N_30436,N_30437,N_30438,N_30439,N_30440,N_30441,N_30442,N_30443,N_30444,N_30445,N_30446,N_30447,N_30448,N_30449,N_30450,N_30451,N_30452,N_30453,N_30454,N_30455,N_30456,N_30457,N_30458,N_30459,N_30460,N_30461,N_30462,N_30463,N_30464,N_30465,N_30466,N_30467,N_30468,N_30469,N_30470,N_30471,N_30472,N_30473,N_30474,N_30475,N_30476,N_30477,N_30478,N_30479,N_30480,N_30481,N_30482,N_30483,N_30484,N_30485,N_30486,N_30487,N_30488,N_30489,N_30490,N_30491,N_30492,N_30493,N_30494,N_30495,N_30496,N_30497,N_30498,N_30499,N_30500,N_30501,N_30502,N_30503,N_30504,N_30505,N_30506,N_30507,N_30508,N_30509,N_30510,N_30511,N_30512,N_30513,N_30514,N_30515,N_30516,N_30517,N_30518,N_30519,N_30520,N_30521,N_30522,N_30523,N_30524,N_30525,N_30526,N_30527,N_30528,N_30529,N_30530,N_30531,N_30532,N_30533,N_30534,N_30535,N_30536,N_30537,N_30538,N_30539,N_30540,N_30541,N_30542,N_30543,N_30544,N_30545,N_30546,N_30547,N_30548,N_30549,N_30550,N_30551,N_30552,N_30553,N_30554,N_30555,N_30556,N_30557,N_30558,N_30559,N_30560,N_30561,N_30562,N_30563,N_30564,N_30565,N_30566,N_30567,N_30568,N_30569,N_30570,N_30571,N_30572,N_30573,N_30574,N_30575,N_30576,N_30577,N_30578,N_30579,N_30580,N_30581,N_30582,N_30583,N_30584,N_30585,N_30586,N_30587,N_30588,N_30589,N_30590,N_30591,N_30592,N_30593,N_30594,N_30595,N_30596,N_30597,N_30598,N_30599,N_30600,N_30601,N_30602,N_30603,N_30604,N_30605,N_30606,N_30607,N_30608,N_30609,N_30610,N_30611,N_30612,N_30613,N_30614,N_30615,N_30616,N_30617,N_30618,N_30619,N_30620,N_30621,N_30622,N_30623,N_30624,N_30625,N_30626,N_30627,N_30628,N_30629,N_30630,N_30631,N_30632,N_30633,N_30634,N_30635,N_30636,N_30637,N_30638,N_30639,N_30640,N_30641,N_30642,N_30643,N_30644,N_30645,N_30646,N_30647,N_30648,N_30649,N_30650,N_30651,N_30652,N_30653,N_30654,N_30655,N_30656,N_30657,N_30658,N_30659,N_30660,N_30661,N_30662,N_30663,N_30664,N_30665,N_30666,N_30667,N_30668,N_30669,N_30670,N_30671,N_30672,N_30673,N_30674,N_30675,N_30676,N_30677,N_30678,N_30679,N_30680,N_30681,N_30682,N_30683,N_30684,N_30685,N_30686,N_30687,N_30688,N_30689,N_30690,N_30691,N_30692,N_30693,N_30694,N_30695,N_30696,N_30697,N_30698,N_30699,N_30700,N_30701,N_30702,N_30703,N_30704,N_30705,N_30706,N_30707,N_30708,N_30709,N_30710,N_30711,N_30712,N_30713,N_30714,N_30715,N_30716,N_30717,N_30718,N_30719,N_30720,N_30721,N_30722,N_30723,N_30724,N_30725,N_30726,N_30727,N_30728,N_30729,N_30730,N_30731,N_30732,N_30733,N_30734,N_30735,N_30736,N_30737,N_30738,N_30739,N_30740,N_30741,N_30742,N_30743,N_30744,N_30745,N_30746,N_30747,N_30748,N_30749,N_30750,N_30751,N_30752,N_30753,N_30754,N_30755,N_30756,N_30757,N_30758,N_30759,N_30760,N_30761,N_30762,N_30763,N_30764,N_30765,N_30766,N_30767,N_30768,N_30769,N_30770,N_30771,N_30772,N_30773,N_30774,N_30775,N_30776,N_30777,N_30778,N_30779,N_30780,N_30781,N_30782,N_30783,N_30784,N_30785,N_30786,N_30787,N_30788,N_30789,N_30790,N_30791,N_30792,N_30793,N_30794,N_30795,N_30796,N_30797,N_30798,N_30799,N_30800,N_30801,N_30802,N_30803,N_30804,N_30805,N_30806,N_30807,N_30808,N_30809,N_30810,N_30811,N_30812,N_30813,N_30814,N_30815,N_30816,N_30817,N_30818,N_30819,N_30820,N_30821,N_30822,N_30823,N_30824,N_30825,N_30826,N_30827,N_30828,N_30829,N_30830,N_30831,N_30832,N_30833,N_30834,N_30835,N_30836,N_30837,N_30838,N_30839,N_30840,N_30841,N_30842,N_30843,N_30844,N_30845,N_30846,N_30847,N_30848,N_30849,N_30850,N_30851,N_30852,N_30853,N_30854,N_30855,N_30856,N_30857,N_30858,N_30859,N_30860,N_30861,N_30862,N_30863,N_30864,N_30865,N_30866,N_30867,N_30868,N_30869,N_30870,N_30871,N_30872,N_30873,N_30874,N_30875,N_30876,N_30877,N_30878,N_30879,N_30880,N_30881,N_30882,N_30883,N_30884,N_30885,N_30886,N_30887,N_30888,N_30889,N_30890,N_30891,N_30892,N_30893,N_30894,N_30895,N_30896,N_30897,N_30898,N_30899,N_30900,N_30901,N_30902,N_30903,N_30904,N_30905,N_30906,N_30907,N_30908,N_30909,N_30910,N_30911,N_30912,N_30913,N_30914,N_30915,N_30916,N_30917,N_30918,N_30919,N_30920,N_30921,N_30922,N_30923,N_30924,N_30925,N_30926,N_30927,N_30928,N_30929,N_30930,N_30931,N_30932,N_30933,N_30934,N_30935,N_30936,N_30937,N_30938,N_30939,N_30940,N_30941,N_30942,N_30943,N_30944,N_30945,N_30946,N_30947,N_30948,N_30949,N_30950,N_30951,N_30952,N_30953,N_30954,N_30955,N_30956,N_30957,N_30958,N_30959,N_30960,N_30961,N_30962,N_30963,N_30964,N_30965,N_30966,N_30967,N_30968,N_30969,N_30970,N_30971,N_30972,N_30973,N_30974,N_30975,N_30976,N_30977,N_30978,N_30979,N_30980,N_30981,N_30982,N_30983,N_30984,N_30985,N_30986,N_30987,N_30988,N_30989,N_30990,N_30991,N_30992,N_30993,N_30994,N_30995,N_30996,N_30997,N_30998,N_30999,N_31000,N_31001,N_31002,N_31003,N_31004,N_31005,N_31006,N_31007,N_31008,N_31009,N_31010,N_31011,N_31012,N_31013,N_31014,N_31015,N_31016,N_31017,N_31018,N_31019,N_31020,N_31021,N_31022,N_31023,N_31024,N_31025,N_31026,N_31027,N_31028,N_31029,N_31030,N_31031,N_31032,N_31033,N_31034,N_31035,N_31036,N_31037,N_31038,N_31039,N_31040,N_31041,N_31042,N_31043,N_31044,N_31045,N_31046,N_31047,N_31048,N_31049,N_31050,N_31051,N_31052,N_31053,N_31054,N_31055,N_31056,N_31057,N_31058,N_31059,N_31060,N_31061,N_31062,N_31063,N_31064,N_31065,N_31066,N_31067,N_31068,N_31069,N_31070,N_31071,N_31072,N_31073,N_31074,N_31075,N_31076,N_31077,N_31078,N_31079,N_31080,N_31081,N_31082,N_31083,N_31084,N_31085,N_31086,N_31087,N_31088,N_31089,N_31090,N_31091,N_31092,N_31093,N_31094,N_31095,N_31096,N_31097,N_31098,N_31099,N_31100,N_31101,N_31102,N_31103,N_31104,N_31105,N_31106,N_31107,N_31108,N_31109,N_31110,N_31111,N_31112,N_31113,N_31114,N_31115,N_31116,N_31117,N_31118,N_31119,N_31120,N_31121,N_31122,N_31123,N_31124,N_31125,N_31126,N_31127,N_31128,N_31129,N_31130,N_31131,N_31132,N_31133,N_31134,N_31135,N_31136,N_31137,N_31138,N_31139,N_31140,N_31141,N_31142,N_31143,N_31144,N_31145,N_31146,N_31147,N_31148,N_31149,N_31150,N_31151,N_31152,N_31153,N_31154,N_31155,N_31156,N_31157,N_31158,N_31159,N_31160,N_31161,N_31162,N_31163,N_31164,N_31165,N_31166,N_31167,N_31168,N_31169,N_31170,N_31171,N_31172,N_31173,N_31174,N_31175,N_31176,N_31177,N_31178,N_31179,N_31180,N_31181,N_31182,N_31183,N_31184,N_31185,N_31186,N_31187,N_31188,N_31189,N_31190,N_31191,N_31192,N_31193,N_31194,N_31195,N_31196,N_31197,N_31198,N_31199,N_31200,N_31201,N_31202,N_31203,N_31204,N_31205,N_31206,N_31207,N_31208,N_31209,N_31210,N_31211,N_31212,N_31213,N_31214,N_31215,N_31216,N_31217,N_31218,N_31219,N_31220,N_31221,N_31222,N_31223,N_31224,N_31225,N_31226,N_31227,N_31228,N_31229,N_31230,N_31231,N_31232,N_31233,N_31234,N_31235,N_31236,N_31237,N_31238,N_31239,N_31240,N_31241,N_31242,N_31243,N_31244,N_31245,N_31246,N_31247,N_31248,N_31249,N_31250,N_31251,N_31252,N_31253,N_31254,N_31255,N_31256,N_31257,N_31258,N_31259,N_31260,N_31261,N_31262,N_31263,N_31264,N_31265,N_31266,N_31267,N_31268,N_31269,N_31270,N_31271,N_31272,N_31273,N_31274,N_31275,N_31276,N_31277,N_31278,N_31279,N_31280,N_31281,N_31282,N_31283,N_31284,N_31285,N_31286,N_31287,N_31288,N_31289,N_31290,N_31291,N_31292,N_31293,N_31294,N_31295,N_31296,N_31297,N_31298,N_31299,N_31300,N_31301,N_31302,N_31303,N_31304,N_31305,N_31306,N_31307,N_31308,N_31309,N_31310,N_31311,N_31312,N_31313,N_31314,N_31315,N_31316,N_31317,N_31318,N_31319,N_31320,N_31321,N_31322,N_31323,N_31324,N_31325,N_31326,N_31327,N_31328,N_31329,N_31330,N_31331,N_31332,N_31333,N_31334,N_31335,N_31336,N_31337,N_31338,N_31339,N_31340,N_31341,N_31342,N_31343,N_31344,N_31345,N_31346,N_31347,N_31348,N_31349,N_31350,N_31351,N_31352,N_31353,N_31354,N_31355,N_31356,N_31357,N_31358,N_31359,N_31360,N_31361,N_31362,N_31363,N_31364,N_31365,N_31366,N_31367,N_31368,N_31369,N_31370,N_31371,N_31372,N_31373,N_31374,N_31375,N_31376,N_31377,N_31378,N_31379,N_31380,N_31381,N_31382,N_31383,N_31384,N_31385,N_31386,N_31387,N_31388,N_31389,N_31390,N_31391,N_31392,N_31393,N_31394,N_31395,N_31396,N_31397,N_31398,N_31399,N_31400,N_31401,N_31402,N_31403,N_31404,N_31405,N_31406,N_31407,N_31408,N_31409,N_31410,N_31411,N_31412,N_31413,N_31414,N_31415,N_31416,N_31417,N_31418,N_31419,N_31420,N_31421,N_31422,N_31423,N_31424,N_31425,N_31426,N_31427,N_31428,N_31429,N_31430,N_31431,N_31432,N_31433,N_31434,N_31435,N_31436,N_31437,N_31438,N_31439,N_31440,N_31441,N_31442,N_31443,N_31444,N_31445,N_31446,N_31447,N_31448,N_31449,N_31450,N_31451,N_31452,N_31453,N_31454,N_31455,N_31456,N_31457,N_31458,N_31459,N_31460,N_31461,N_31462,N_31463,N_31464,N_31465,N_31466,N_31467,N_31468,N_31469,N_31470,N_31471,N_31472,N_31473,N_31474,N_31475,N_31476,N_31477,N_31478,N_31479,N_31480,N_31481,N_31482,N_31483,N_31484,N_31485,N_31486,N_31487,N_31488,N_31489,N_31490,N_31491,N_31492,N_31493,N_31494,N_31495,N_31496,N_31497,N_31498,N_31499,N_31500,N_31501,N_31502,N_31503,N_31504,N_31505,N_31506,N_31507,N_31508,N_31509,N_31510,N_31511,N_31512,N_31513,N_31514,N_31515,N_31516,N_31517,N_31518,N_31519,N_31520,N_31521,N_31522,N_31523,N_31524,N_31525,N_31526,N_31527,N_31528,N_31529,N_31530,N_31531,N_31532,N_31533,N_31534,N_31535,N_31536,N_31537,N_31538,N_31539,N_31540,N_31541,N_31542,N_31543,N_31544,N_31545,N_31546,N_31547,N_31548,N_31549,N_31550,N_31551,N_31552,N_31553,N_31554,N_31555,N_31556,N_31557,N_31558,N_31559,N_31560,N_31561,N_31562,N_31563,N_31564,N_31565,N_31566,N_31567,N_31568,N_31569,N_31570,N_31571,N_31572,N_31573,N_31574,N_31575,N_31576,N_31577,N_31578,N_31579,N_31580,N_31581,N_31582,N_31583,N_31584,N_31585,N_31586,N_31587,N_31588,N_31589,N_31590,N_31591,N_31592,N_31593,N_31594,N_31595,N_31596,N_31597,N_31598,N_31599,N_31600,N_31601,N_31602,N_31603,N_31604,N_31605,N_31606,N_31607,N_31608,N_31609,N_31610,N_31611,N_31612,N_31613,N_31614,N_31615,N_31616,N_31617,N_31618,N_31619,N_31620,N_31621,N_31622,N_31623,N_31624,N_31625,N_31626,N_31627,N_31628,N_31629,N_31630,N_31631,N_31632,N_31633,N_31634,N_31635,N_31636,N_31637,N_31638,N_31639,N_31640,N_31641,N_31642,N_31643,N_31644,N_31645,N_31646,N_31647,N_31648,N_31649,N_31650,N_31651,N_31652,N_31653,N_31654,N_31655,N_31656,N_31657,N_31658,N_31659,N_31660,N_31661,N_31662,N_31663,N_31664,N_31665,N_31666,N_31667,N_31668,N_31669,N_31670,N_31671,N_31672,N_31673,N_31674,N_31675,N_31676,N_31677,N_31678,N_31679,N_31680,N_31681,N_31682,N_31683,N_31684,N_31685,N_31686,N_31687,N_31688,N_31689,N_31690,N_31691,N_31692,N_31693,N_31694,N_31695,N_31696,N_31697,N_31698,N_31699,N_31700,N_31701,N_31702,N_31703,N_31704,N_31705,N_31706,N_31707,N_31708,N_31709,N_31710,N_31711,N_31712,N_31713,N_31714,N_31715,N_31716,N_31717,N_31718,N_31719,N_31720,N_31721,N_31722,N_31723,N_31724,N_31725,N_31726,N_31727,N_31728,N_31729,N_31730,N_31731,N_31732,N_31733,N_31734,N_31735,N_31736,N_31737,N_31738,N_31739,N_31740,N_31741,N_31742,N_31743,N_31744,N_31745,N_31746,N_31747,N_31748,N_31749,N_31750,N_31751,N_31752,N_31753,N_31754,N_31755,N_31756,N_31757,N_31758,N_31759,N_31760,N_31761,N_31762,N_31763,N_31764,N_31765,N_31766,N_31767,N_31768,N_31769,N_31770,N_31771,N_31772,N_31773,N_31774,N_31775,N_31776,N_31777,N_31778,N_31779,N_31780,N_31781,N_31782,N_31783,N_31784,N_31785,N_31786,N_31787,N_31788,N_31789,N_31790,N_31791,N_31792,N_31793,N_31794,N_31795,N_31796,N_31797,N_31798,N_31799,N_31800,N_31801,N_31802,N_31803,N_31804,N_31805,N_31806,N_31807,N_31808,N_31809,N_31810,N_31811,N_31812,N_31813,N_31814,N_31815,N_31816,N_31817,N_31818,N_31819,N_31820,N_31821,N_31822,N_31823,N_31824,N_31825,N_31826,N_31827,N_31828,N_31829,N_31830,N_31831,N_31832,N_31833,N_31834,N_31835,N_31836,N_31837,N_31838,N_31839,N_31840,N_31841,N_31842,N_31843,N_31844,N_31845,N_31846,N_31847,N_31848,N_31849,N_31850,N_31851,N_31852,N_31853,N_31854,N_31855,N_31856,N_31857,N_31858,N_31859,N_31860,N_31861,N_31862,N_31863,N_31864,N_31865,N_31866,N_31867,N_31868,N_31869,N_31870,N_31871,N_31872,N_31873,N_31874,N_31875,N_31876,N_31877,N_31878,N_31879,N_31880,N_31881,N_31882,N_31883,N_31884,N_31885,N_31886,N_31887,N_31888,N_31889,N_31890,N_31891,N_31892,N_31893,N_31894,N_31895,N_31896,N_31897,N_31898,N_31899,N_31900,N_31901,N_31902,N_31903,N_31904,N_31905,N_31906,N_31907,N_31908,N_31909,N_31910,N_31911,N_31912,N_31913,N_31914,N_31915,N_31916,N_31917,N_31918,N_31919,N_31920,N_31921,N_31922,N_31923,N_31924,N_31925,N_31926,N_31927,N_31928,N_31929,N_31930,N_31931,N_31932,N_31933,N_31934,N_31935,N_31936,N_31937,N_31938,N_31939,N_31940,N_31941,N_31942,N_31943,N_31944,N_31945,N_31946,N_31947,N_31948,N_31949,N_31950,N_31951,N_31952,N_31953,N_31954,N_31955,N_31956,N_31957,N_31958,N_31959,N_31960,N_31961,N_31962,N_31963,N_31964,N_31965,N_31966,N_31967,N_31968,N_31969,N_31970,N_31971,N_31972,N_31973,N_31974,N_31975,N_31976,N_31977,N_31978,N_31979,N_31980,N_31981,N_31982,N_31983,N_31984,N_31985,N_31986,N_31987,N_31988,N_31989,N_31990,N_31991,N_31992,N_31993,N_31994,N_31995,N_31996,N_31997,N_31998,N_31999,N_32000,N_32001,N_32002,N_32003,N_32004,N_32005,N_32006,N_32007,N_32008,N_32009,N_32010,N_32011,N_32012,N_32013,N_32014,N_32015,N_32016,N_32017,N_32018,N_32019,N_32020,N_32021,N_32022,N_32023,N_32024,N_32025,N_32026,N_32027,N_32028,N_32029,N_32030,N_32031,N_32032,N_32033,N_32034,N_32035,N_32036,N_32037,N_32038,N_32039,N_32040,N_32041,N_32042,N_32043,N_32044,N_32045,N_32046,N_32047,N_32048,N_32049,N_32050,N_32051,N_32052,N_32053,N_32054,N_32055,N_32056,N_32057,N_32058,N_32059,N_32060,N_32061,N_32062,N_32063,N_32064,N_32065,N_32066,N_32067,N_32068,N_32069,N_32070,N_32071,N_32072,N_32073,N_32074,N_32075,N_32076,N_32077,N_32078,N_32079,N_32080,N_32081,N_32082,N_32083,N_32084,N_32085,N_32086,N_32087,N_32088,N_32089,N_32090,N_32091,N_32092,N_32093,N_32094,N_32095,N_32096,N_32097,N_32098,N_32099,N_32100,N_32101,N_32102,N_32103,N_32104,N_32105,N_32106,N_32107,N_32108,N_32109,N_32110,N_32111,N_32112,N_32113,N_32114,N_32115,N_32116,N_32117,N_32118,N_32119,N_32120,N_32121,N_32122,N_32123,N_32124,N_32125,N_32126,N_32127,N_32128,N_32129,N_32130,N_32131,N_32132,N_32133,N_32134,N_32135,N_32136,N_32137,N_32138,N_32139,N_32140,N_32141,N_32142,N_32143,N_32144,N_32145,N_32146,N_32147,N_32148,N_32149,N_32150,N_32151,N_32152,N_32153,N_32154,N_32155,N_32156,N_32157,N_32158,N_32159,N_32160,N_32161,N_32162,N_32163,N_32164,N_32165,N_32166,N_32167,N_32168,N_32169,N_32170,N_32171,N_32172,N_32173,N_32174,N_32175,N_32176,N_32177,N_32178,N_32179,N_32180,N_32181,N_32182,N_32183,N_32184,N_32185,N_32186,N_32187,N_32188,N_32189,N_32190,N_32191,N_32192,N_32193,N_32194,N_32195,N_32196,N_32197,N_32198,N_32199,N_32200,N_32201,N_32202,N_32203,N_32204,N_32205,N_32206,N_32207,N_32208,N_32209,N_32210,N_32211,N_32212,N_32213,N_32214,N_32215,N_32216,N_32217,N_32218,N_32219,N_32220,N_32221,N_32222,N_32223,N_32224,N_32225,N_32226,N_32227,N_32228,N_32229,N_32230,N_32231,N_32232,N_32233,N_32234,N_32235,N_32236,N_32237,N_32238,N_32239,N_32240,N_32241,N_32242,N_32243,N_32244,N_32245,N_32246,N_32247,N_32248,N_32249,N_32250,N_32251,N_32252,N_32253,N_32254,N_32255,N_32256,N_32257,N_32258,N_32259,N_32260,N_32261,N_32262,N_32263,N_32264,N_32265,N_32266,N_32267,N_32268,N_32269,N_32270,N_32271,N_32272,N_32273,N_32274,N_32275,N_32276,N_32277,N_32278,N_32279,N_32280,N_32281,N_32282,N_32283,N_32284,N_32285,N_32286,N_32287,N_32288,N_32289,N_32290,N_32291,N_32292,N_32293,N_32294,N_32295,N_32296,N_32297,N_32298,N_32299,N_32300,N_32301,N_32302,N_32303,N_32304,N_32305,N_32306,N_32307,N_32308,N_32309,N_32310,N_32311,N_32312,N_32313,N_32314,N_32315,N_32316,N_32317,N_32318,N_32319,N_32320,N_32321,N_32322,N_32323,N_32324,N_32325,N_32326,N_32327,N_32328,N_32329,N_32330,N_32331,N_32332,N_32333,N_32334,N_32335,N_32336,N_32337,N_32338,N_32339,N_32340,N_32341,N_32342,N_32343,N_32344,N_32345,N_32346,N_32347,N_32348,N_32349,N_32350,N_32351,N_32352,N_32353,N_32354,N_32355,N_32356,N_32357,N_32358,N_32359,N_32360,N_32361,N_32362,N_32363,N_32364,N_32365,N_32366,N_32367,N_32368,N_32369,N_32370,N_32371,N_32372,N_32373,N_32374,N_32375,N_32376,N_32377,N_32378,N_32379,N_32380,N_32381,N_32382,N_32383,N_32384,N_32385,N_32386,N_32387,N_32388,N_32389,N_32390,N_32391,N_32392,N_32393,N_32394,N_32395,N_32396,N_32397,N_32398,N_32399,N_32400,N_32401,N_32402,N_32403,N_32404,N_32405,N_32406,N_32407,N_32408,N_32409,N_32410,N_32411,N_32412,N_32413,N_32414,N_32415,N_32416,N_32417,N_32418,N_32419,N_32420,N_32421,N_32422,N_32423,N_32424,N_32425,N_32426,N_32427,N_32428,N_32429,N_32430,N_32431,N_32432,N_32433,N_32434,N_32435,N_32436,N_32437,N_32438,N_32439,N_32440,N_32441,N_32442,N_32443,N_32444,N_32445,N_32446,N_32447,N_32448,N_32449,N_32450,N_32451,N_32452,N_32453,N_32454,N_32455,N_32456,N_32457,N_32458,N_32459,N_32460,N_32461,N_32462,N_32463,N_32464,N_32465,N_32466,N_32467,N_32468,N_32469,N_32470,N_32471,N_32472,N_32473,N_32474,N_32475,N_32476,N_32477,N_32478,N_32479,N_32480,N_32481,N_32482,N_32483,N_32484,N_32485,N_32486,N_32487,N_32488,N_32489,N_32490,N_32491,N_32492,N_32493,N_32494,N_32495,N_32496,N_32497,N_32498,N_32499,N_32500,N_32501,N_32502,N_32503,N_32504,N_32505,N_32506,N_32507,N_32508,N_32509,N_32510,N_32511,N_32512,N_32513,N_32514,N_32515,N_32516,N_32517,N_32518,N_32519,N_32520,N_32521,N_32522,N_32523,N_32524,N_32525,N_32526,N_32527,N_32528,N_32529,N_32530,N_32531,N_32532,N_32533,N_32534,N_32535,N_32536,N_32537,N_32538,N_32539,N_32540,N_32541,N_32542,N_32543,N_32544,N_32545,N_32546,N_32547,N_32548,N_32549,N_32550,N_32551,N_32552,N_32553,N_32554,N_32555,N_32556,N_32557,N_32558,N_32559,N_32560,N_32561,N_32562,N_32563,N_32564,N_32565,N_32566,N_32567,N_32568,N_32569,N_32570,N_32571,N_32572,N_32573,N_32574,N_32575,N_32576,N_32577,N_32578,N_32579,N_32580,N_32581,N_32582,N_32583,N_32584,N_32585,N_32586,N_32587,N_32588,N_32589,N_32590,N_32591,N_32592,N_32593,N_32594,N_32595,N_32596,N_32597,N_32598,N_32599,N_32600,N_32601,N_32602,N_32603,N_32604,N_32605,N_32606,N_32607,N_32608,N_32609,N_32610,N_32611,N_32612,N_32613,N_32614,N_32615,N_32616,N_32617,N_32618,N_32619,N_32620,N_32621,N_32622,N_32623,N_32624,N_32625,N_32626,N_32627,N_32628,N_32629,N_32630,N_32631,N_32632,N_32633,N_32634,N_32635,N_32636,N_32637,N_32638,N_32639,N_32640,N_32641,N_32642,N_32643,N_32644,N_32645,N_32646,N_32647,N_32648,N_32649,N_32650,N_32651,N_32652,N_32653,N_32654,N_32655,N_32656,N_32657,N_32658,N_32659,N_32660,N_32661,N_32662,N_32663,N_32664,N_32665,N_32666,N_32667,N_32668,N_32669,N_32670,N_32671,N_32672,N_32673,N_32674,N_32675,N_32676,N_32677,N_32678,N_32679,N_32680,N_32681,N_32682,N_32683,N_32684,N_32685,N_32686,N_32687,N_32688,N_32689,N_32690,N_32691,N_32692,N_32693,N_32694,N_32695,N_32696,N_32697,N_32698,N_32699,N_32700,N_32701,N_32702,N_32703,N_32704,N_32705,N_32706,N_32707,N_32708,N_32709,N_32710,N_32711,N_32712,N_32713,N_32714,N_32715,N_32716,N_32717,N_32718,N_32719,N_32720,N_32721,N_32722,N_32723,N_32724,N_32725,N_32726,N_32727,N_32728,N_32729,N_32730,N_32731,N_32732,N_32733,N_32734,N_32735,N_32736,N_32737,N_32738,N_32739,N_32740,N_32741,N_32742,N_32743,N_32744,N_32745,N_32746,N_32747,N_32748,N_32749,N_32750,N_32751,N_32752,N_32753,N_32754,N_32755,N_32756,N_32757,N_32758,N_32759,N_32760,N_32761,N_32762,N_32763,N_32764,N_32765,N_32766,N_32767,N_32768,N_32769,N_32770,N_32771,N_32772,N_32773,N_32774,N_32775,N_32776,N_32777,N_32778,N_32779,N_32780,N_32781,N_32782,N_32783,N_32784,N_32785,N_32786,N_32787,N_32788,N_32789,N_32790,N_32791,N_32792,N_32793,N_32794,N_32795,N_32796,N_32797,N_32798,N_32799,N_32800,N_32801,N_32802,N_32803,N_32804,N_32805,N_32806,N_32807,N_32808,N_32809,N_32810,N_32811,N_32812,N_32813,N_32814,N_32815,N_32816,N_32817,N_32818,N_32819,N_32820,N_32821,N_32822,N_32823,N_32824,N_32825,N_32826,N_32827,N_32828,N_32829,N_32830,N_32831,N_32832,N_32833,N_32834,N_32835,N_32836,N_32837,N_32838,N_32839,N_32840,N_32841,N_32842,N_32843,N_32844,N_32845,N_32846,N_32847,N_32848,N_32849,N_32850,N_32851,N_32852,N_32853,N_32854,N_32855,N_32856,N_32857,N_32858,N_32859,N_32860,N_32861,N_32862,N_32863,N_32864,N_32865,N_32866,N_32867,N_32868,N_32869,N_32870,N_32871,N_32872,N_32873,N_32874,N_32875,N_32876,N_32877,N_32878,N_32879,N_32880,N_32881,N_32882,N_32883,N_32884,N_32885,N_32886,N_32887,N_32888,N_32889,N_32890,N_32891,N_32892,N_32893,N_32894,N_32895,N_32896,N_32897,N_32898,N_32899,N_32900,N_32901,N_32902,N_32903,N_32904,N_32905,N_32906,N_32907,N_32908,N_32909,N_32910,N_32911,N_32912,N_32913,N_32914,N_32915,N_32916,N_32917,N_32918,N_32919,N_32920,N_32921,N_32922,N_32923,N_32924,N_32925,N_32926,N_32927,N_32928,N_32929,N_32930,N_32931,N_32932,N_32933,N_32934,N_32935,N_32936,N_32937,N_32938,N_32939,N_32940,N_32941,N_32942,N_32943,N_32944,N_32945,N_32946,N_32947,N_32948,N_32949,N_32950,N_32951,N_32952,N_32953,N_32954,N_32955,N_32956,N_32957,N_32958,N_32959,N_32960,N_32961,N_32962,N_32963,N_32964,N_32965,N_32966,N_32967,N_32968,N_32969,N_32970,N_32971,N_32972,N_32973,N_32974,N_32975,N_32976,N_32977,N_32978,N_32979,N_32980,N_32981,N_32982,N_32983,N_32984,N_32985,N_32986,N_32987,N_32988,N_32989,N_32990,N_32991,N_32992,N_32993,N_32994,N_32995,N_32996,N_32997,N_32998,N_32999,N_33000,N_33001,N_33002,N_33003,N_33004,N_33005,N_33006,N_33007,N_33008,N_33009,N_33010,N_33011,N_33012,N_33013,N_33014,N_33015,N_33016,N_33017,N_33018,N_33019,N_33020,N_33021,N_33022,N_33023,N_33024,N_33025,N_33026,N_33027,N_33028,N_33029,N_33030,N_33031,N_33032,N_33033,N_33034,N_33035,N_33036,N_33037,N_33038,N_33039,N_33040,N_33041,N_33042,N_33043,N_33044,N_33045,N_33046,N_33047,N_33048,N_33049,N_33050,N_33051,N_33052,N_33053,N_33054,N_33055,N_33056,N_33057,N_33058,N_33059,N_33060,N_33061,N_33062,N_33063,N_33064,N_33065,N_33066,N_33067,N_33068,N_33069,N_33070,N_33071,N_33072,N_33073,N_33074,N_33075,N_33076,N_33077,N_33078,N_33079,N_33080,N_33081,N_33082,N_33083,N_33084,N_33085,N_33086,N_33087,N_33088,N_33089,N_33090,N_33091,N_33092,N_33093,N_33094,N_33095,N_33096,N_33097,N_33098,N_33099,N_33100,N_33101,N_33102,N_33103,N_33104,N_33105,N_33106,N_33107,N_33108,N_33109,N_33110,N_33111,N_33112,N_33113,N_33114,N_33115,N_33116,N_33117,N_33118,N_33119,N_33120,N_33121,N_33122,N_33123,N_33124,N_33125,N_33126,N_33127,N_33128,N_33129,N_33130,N_33131,N_33132,N_33133,N_33134,N_33135,N_33136,N_33137,N_33138,N_33139,N_33140,N_33141,N_33142,N_33143,N_33144,N_33145,N_33146,N_33147,N_33148,N_33149,N_33150,N_33151,N_33152,N_33153,N_33154,N_33155,N_33156,N_33157,N_33158,N_33159,N_33160,N_33161,N_33162,N_33163,N_33164,N_33165,N_33166,N_33167,N_33168,N_33169,N_33170,N_33171,N_33172,N_33173,N_33174,N_33175,N_33176,N_33177,N_33178,N_33179,N_33180,N_33181,N_33182,N_33183,N_33184,N_33185,N_33186,N_33187,N_33188,N_33189,N_33190,N_33191,N_33192,N_33193,N_33194,N_33195,N_33196,N_33197,N_33198,N_33199,N_33200,N_33201,N_33202,N_33203,N_33204,N_33205,N_33206,N_33207,N_33208,N_33209,N_33210,N_33211,N_33212,N_33213,N_33214,N_33215,N_33216,N_33217,N_33218,N_33219,N_33220,N_33221,N_33222,N_33223,N_33224,N_33225,N_33226,N_33227,N_33228,N_33229,N_33230,N_33231,N_33232,N_33233,N_33234,N_33235,N_33236,N_33237,N_33238,N_33239,N_33240,N_33241,N_33242,N_33243,N_33244,N_33245,N_33246,N_33247,N_33248,N_33249,N_33250,N_33251,N_33252,N_33253,N_33254,N_33255,N_33256,N_33257,N_33258,N_33259,N_33260,N_33261,N_33262,N_33263,N_33264,N_33265,N_33266,N_33267,N_33268,N_33269,N_33270,N_33271,N_33272,N_33273,N_33274,N_33275,N_33276,N_33277,N_33278,N_33279,N_33280,N_33281,N_33282,N_33283,N_33284,N_33285,N_33286,N_33287,N_33288,N_33289,N_33290,N_33291,N_33292,N_33293,N_33294,N_33295,N_33296,N_33297,N_33298,N_33299,N_33300,N_33301,N_33302,N_33303,N_33304,N_33305,N_33306,N_33307,N_33308,N_33309,N_33310,N_33311,N_33312,N_33313,N_33314,N_33315,N_33316,N_33317,N_33318,N_33319,N_33320,N_33321,N_33322,N_33323,N_33324,N_33325,N_33326,N_33327,N_33328,N_33329,N_33330,N_33331,N_33332,N_33333,N_33334,N_33335,N_33336,N_33337,N_33338,N_33339,N_33340,N_33341,N_33342,N_33343,N_33344,N_33345,N_33346,N_33347,N_33348,N_33349,N_33350,N_33351,N_33352,N_33353,N_33354,N_33355,N_33356,N_33357,N_33358,N_33359,N_33360,N_33361,N_33362,N_33363,N_33364,N_33365,N_33366,N_33367,N_33368,N_33369,N_33370,N_33371,N_33372,N_33373,N_33374,N_33375,N_33376,N_33377,N_33378,N_33379,N_33380,N_33381,N_33382,N_33383,N_33384,N_33385,N_33386,N_33387,N_33388,N_33389,N_33390,N_33391,N_33392,N_33393,N_33394,N_33395,N_33396,N_33397,N_33398,N_33399,N_33400,N_33401,N_33402,N_33403,N_33404,N_33405,N_33406,N_33407,N_33408,N_33409,N_33410,N_33411,N_33412,N_33413,N_33414,N_33415,N_33416,N_33417,N_33418,N_33419,N_33420,N_33421,N_33422,N_33423,N_33424,N_33425,N_33426,N_33427,N_33428,N_33429,N_33430,N_33431,N_33432,N_33433,N_33434,N_33435,N_33436,N_33437,N_33438,N_33439,N_33440,N_33441,N_33442,N_33443,N_33444,N_33445,N_33446,N_33447,N_33448,N_33449,N_33450,N_33451,N_33452,N_33453,N_33454,N_33455,N_33456,N_33457,N_33458,N_33459,N_33460,N_33461,N_33462,N_33463,N_33464,N_33465,N_33466,N_33467,N_33468,N_33469,N_33470,N_33471,N_33472,N_33473,N_33474,N_33475,N_33476,N_33477,N_33478,N_33479,N_33480,N_33481,N_33482,N_33483,N_33484,N_33485,N_33486,N_33487,N_33488,N_33489,N_33490,N_33491,N_33492,N_33493,N_33494,N_33495,N_33496,N_33497,N_33498,N_33499,N_33500,N_33501,N_33502,N_33503,N_33504,N_33505,N_33506,N_33507,N_33508,N_33509,N_33510,N_33511,N_33512,N_33513,N_33514,N_33515,N_33516,N_33517,N_33518,N_33519,N_33520,N_33521,N_33522,N_33523,N_33524,N_33525,N_33526,N_33527,N_33528,N_33529,N_33530,N_33531,N_33532,N_33533,N_33534,N_33535,N_33536,N_33537,N_33538,N_33539,N_33540,N_33541,N_33542,N_33543,N_33544,N_33545,N_33546,N_33547,N_33548,N_33549,N_33550,N_33551,N_33552,N_33553,N_33554,N_33555,N_33556,N_33557,N_33558,N_33559,N_33560,N_33561,N_33562,N_33563,N_33564,N_33565,N_33566,N_33567,N_33568,N_33569,N_33570,N_33571,N_33572,N_33573,N_33574,N_33575,N_33576,N_33577,N_33578,N_33579,N_33580,N_33581,N_33582,N_33583,N_33584,N_33585,N_33586,N_33587,N_33588,N_33589,N_33590,N_33591,N_33592,N_33593,N_33594,N_33595,N_33596,N_33597,N_33598,N_33599,N_33600,N_33601,N_33602,N_33603,N_33604,N_33605,N_33606,N_33607,N_33608,N_33609,N_33610,N_33611,N_33612,N_33613,N_33614,N_33615,N_33616,N_33617,N_33618,N_33619,N_33620,N_33621,N_33622,N_33623,N_33624,N_33625,N_33626,N_33627,N_33628,N_33629,N_33630,N_33631,N_33632,N_33633,N_33634,N_33635,N_33636,N_33637,N_33638,N_33639,N_33640,N_33641,N_33642,N_33643,N_33644,N_33645,N_33646,N_33647,N_33648,N_33649,N_33650,N_33651,N_33652,N_33653,N_33654,N_33655,N_33656,N_33657,N_33658,N_33659,N_33660,N_33661,N_33662,N_33663,N_33664,N_33665,N_33666,N_33667,N_33668,N_33669,N_33670,N_33671,N_33672,N_33673,N_33674,N_33675,N_33676,N_33677,N_33678,N_33679,N_33680,N_33681,N_33682,N_33683,N_33684,N_33685,N_33686,N_33687,N_33688,N_33689,N_33690,N_33691,N_33692,N_33693,N_33694,N_33695,N_33696,N_33697,N_33698,N_33699,N_33700,N_33701,N_33702,N_33703,N_33704,N_33705,N_33706,N_33707,N_33708,N_33709,N_33710,N_33711,N_33712,N_33713,N_33714,N_33715,N_33716,N_33717,N_33718,N_33719,N_33720,N_33721,N_33722,N_33723,N_33724,N_33725,N_33726,N_33727,N_33728,N_33729,N_33730,N_33731,N_33732,N_33733,N_33734,N_33735,N_33736,N_33737,N_33738,N_33739,N_33740,N_33741,N_33742,N_33743,N_33744,N_33745,N_33746,N_33747,N_33748,N_33749,N_33750,N_33751,N_33752,N_33753,N_33754,N_33755,N_33756,N_33757,N_33758,N_33759,N_33760,N_33761,N_33762,N_33763,N_33764,N_33765,N_33766,N_33767,N_33768,N_33769,N_33770,N_33771,N_33772,N_33773,N_33774,N_33775,N_33776,N_33777,N_33778,N_33779,N_33780,N_33781,N_33782,N_33783,N_33784,N_33785,N_33786,N_33787,N_33788,N_33789,N_33790,N_33791,N_33792,N_33793,N_33794,N_33795,N_33796,N_33797,N_33798,N_33799,N_33800,N_33801,N_33802,N_33803,N_33804,N_33805,N_33806,N_33807,N_33808,N_33809,N_33810,N_33811,N_33812,N_33813,N_33814,N_33815,N_33816,N_33817,N_33818,N_33819,N_33820,N_33821,N_33822,N_33823,N_33824,N_33825,N_33826,N_33827,N_33828,N_33829,N_33830,N_33831,N_33832,N_33833,N_33834,N_33835,N_33836,N_33837,N_33838,N_33839,N_33840,N_33841,N_33842,N_33843,N_33844,N_33845,N_33846,N_33847,N_33848,N_33849,N_33850,N_33851,N_33852,N_33853,N_33854,N_33855,N_33856,N_33857,N_33858,N_33859,N_33860,N_33861,N_33862,N_33863,N_33864,N_33865,N_33866,N_33867,N_33868,N_33869,N_33870,N_33871,N_33872,N_33873,N_33874,N_33875,N_33876,N_33877,N_33878,N_33879,N_33880,N_33881,N_33882,N_33883,N_33884,N_33885,N_33886,N_33887,N_33888,N_33889,N_33890,N_33891,N_33892,N_33893,N_33894,N_33895,N_33896,N_33897,N_33898,N_33899,N_33900,N_33901,N_33902,N_33903,N_33904,N_33905,N_33906,N_33907,N_33908,N_33909,N_33910,N_33911,N_33912,N_33913,N_33914,N_33915,N_33916,N_33917,N_33918,N_33919,N_33920,N_33921,N_33922,N_33923,N_33924,N_33925,N_33926,N_33927,N_33928,N_33929,N_33930,N_33931,N_33932,N_33933,N_33934,N_33935,N_33936,N_33937,N_33938,N_33939,N_33940,N_33941,N_33942,N_33943,N_33944,N_33945,N_33946,N_33947,N_33948,N_33949,N_33950,N_33951,N_33952,N_33953,N_33954,N_33955,N_33956,N_33957,N_33958,N_33959,N_33960,N_33961,N_33962,N_33963,N_33964,N_33965,N_33966,N_33967,N_33968,N_33969,N_33970,N_33971,N_33972,N_33973,N_33974,N_33975,N_33976,N_33977,N_33978,N_33979,N_33980,N_33981,N_33982,N_33983,N_33984,N_33985,N_33986,N_33987,N_33988,N_33989,N_33990,N_33991,N_33992,N_33993,N_33994,N_33995,N_33996,N_33997,N_33998,N_33999,N_34000,N_34001,N_34002,N_34003,N_34004,N_34005,N_34006,N_34007,N_34008,N_34009,N_34010,N_34011,N_34012,N_34013,N_34014,N_34015,N_34016,N_34017,N_34018,N_34019,N_34020,N_34021,N_34022,N_34023,N_34024,N_34025,N_34026,N_34027,N_34028,N_34029,N_34030,N_34031,N_34032,N_34033,N_34034,N_34035,N_34036,N_34037,N_34038,N_34039,N_34040,N_34041,N_34042,N_34043,N_34044,N_34045,N_34046,N_34047,N_34048,N_34049,N_34050,N_34051,N_34052,N_34053,N_34054,N_34055,N_34056,N_34057,N_34058,N_34059,N_34060,N_34061,N_34062,N_34063,N_34064,N_34065,N_34066,N_34067,N_34068,N_34069,N_34070,N_34071,N_34072,N_34073,N_34074,N_34075,N_34076,N_34077,N_34078,N_34079,N_34080,N_34081,N_34082,N_34083,N_34084,N_34085,N_34086,N_34087,N_34088,N_34089,N_34090,N_34091,N_34092,N_34093,N_34094,N_34095,N_34096,N_34097,N_34098,N_34099,N_34100,N_34101,N_34102,N_34103,N_34104,N_34105,N_34106,N_34107,N_34108,N_34109,N_34110,N_34111,N_34112,N_34113,N_34114,N_34115,N_34116,N_34117,N_34118,N_34119,N_34120,N_34121,N_34122,N_34123,N_34124,N_34125,N_34126,N_34127,N_34128,N_34129,N_34130,N_34131,N_34132,N_34133,N_34134,N_34135,N_34136,N_34137,N_34138,N_34139,N_34140,N_34141,N_34142,N_34143,N_34144,N_34145,N_34146,N_34147,N_34148,N_34149,N_34150,N_34151,N_34152,N_34153,N_34154,N_34155,N_34156,N_34157,N_34158,N_34159,N_34160,N_34161,N_34162,N_34163,N_34164,N_34165,N_34166,N_34167,N_34168,N_34169,N_34170,N_34171,N_34172,N_34173,N_34174,N_34175,N_34176,N_34177,N_34178,N_34179,N_34180,N_34181,N_34182,N_34183,N_34184,N_34185,N_34186,N_34187,N_34188,N_34189,N_34190,N_34191,N_34192,N_34193,N_34194,N_34195,N_34196,N_34197,N_34198,N_34199,N_34200,N_34201,N_34202,N_34203,N_34204,N_34205,N_34206,N_34207,N_34208,N_34209,N_34210,N_34211,N_34212,N_34213,N_34214,N_34215,N_34216,N_34217,N_34218,N_34219,N_34220,N_34221,N_34222,N_34223,N_34224,N_34225,N_34226,N_34227,N_34228,N_34229,N_34230,N_34231,N_34232,N_34233,N_34234,N_34235,N_34236,N_34237,N_34238,N_34239,N_34240,N_34241,N_34242,N_34243,N_34244,N_34245,N_34246,N_34247,N_34248,N_34249,N_34250,N_34251,N_34252,N_34253,N_34254,N_34255,N_34256,N_34257,N_34258,N_34259,N_34260,N_34261,N_34262,N_34263,N_34264,N_34265,N_34266,N_34267,N_34268,N_34269,N_34270,N_34271,N_34272,N_34273,N_34274,N_34275,N_34276,N_34277,N_34278,N_34279,N_34280,N_34281,N_34282,N_34283,N_34284,N_34285,N_34286,N_34287,N_34288,N_34289,N_34290,N_34291,N_34292,N_34293,N_34294,N_34295,N_34296,N_34297,N_34298,N_34299,N_34300,N_34301,N_34302,N_34303,N_34304,N_34305,N_34306,N_34307,N_34308,N_34309,N_34310,N_34311,N_34312,N_34313,N_34314,N_34315,N_34316,N_34317,N_34318,N_34319,N_34320,N_34321,N_34322,N_34323,N_34324,N_34325,N_34326,N_34327,N_34328,N_34329,N_34330,N_34331,N_34332,N_34333,N_34334,N_34335,N_34336,N_34337,N_34338,N_34339,N_34340,N_34341,N_34342,N_34343,N_34344,N_34345,N_34346,N_34347,N_34348,N_34349,N_34350,N_34351,N_34352,N_34353,N_34354,N_34355,N_34356,N_34357,N_34358,N_34359,N_34360,N_34361,N_34362,N_34363,N_34364,N_34365,N_34366,N_34367,N_34368,N_34369,N_34370,N_34371,N_34372,N_34373,N_34374,N_34375,N_34376,N_34377,N_34378,N_34379,N_34380,N_34381,N_34382,N_34383,N_34384,N_34385,N_34386,N_34387,N_34388,N_34389,N_34390,N_34391,N_34392,N_34393,N_34394,N_34395,N_34396,N_34397,N_34398,N_34399,N_34400,N_34401,N_34402,N_34403,N_34404,N_34405,N_34406,N_34407,N_34408,N_34409,N_34410,N_34411,N_34412,N_34413,N_34414,N_34415,N_34416,N_34417,N_34418,N_34419,N_34420,N_34421,N_34422,N_34423,N_34424,N_34425,N_34426,N_34427,N_34428,N_34429,N_34430,N_34431,N_34432,N_34433,N_34434,N_34435,N_34436,N_34437,N_34438,N_34439,N_34440,N_34441,N_34442,N_34443,N_34444,N_34445,N_34446,N_34447,N_34448,N_34449,N_34450,N_34451,N_34452,N_34453,N_34454,N_34455,N_34456,N_34457,N_34458,N_34459,N_34460,N_34461,N_34462,N_34463,N_34464,N_34465,N_34466,N_34467,N_34468,N_34469,N_34470,N_34471,N_34472,N_34473,N_34474,N_34475,N_34476,N_34477,N_34478,N_34479,N_34480,N_34481,N_34482,N_34483,N_34484,N_34485,N_34486,N_34487,N_34488,N_34489,N_34490,N_34491,N_34492,N_34493,N_34494,N_34495,N_34496,N_34497,N_34498,N_34499,N_34500,N_34501,N_34502,N_34503,N_34504,N_34505,N_34506,N_34507,N_34508,N_34509,N_34510,N_34511,N_34512,N_34513,N_34514,N_34515,N_34516,N_34517,N_34518,N_34519,N_34520,N_34521,N_34522,N_34523,N_34524,N_34525,N_34526,N_34527,N_34528,N_34529,N_34530,N_34531,N_34532,N_34533,N_34534,N_34535,N_34536,N_34537,N_34538,N_34539,N_34540,N_34541,N_34542,N_34543,N_34544,N_34545,N_34546,N_34547,N_34548,N_34549,N_34550,N_34551,N_34552,N_34553,N_34554,N_34555,N_34556,N_34557,N_34558,N_34559,N_34560,N_34561,N_34562,N_34563,N_34564,N_34565,N_34566,N_34567,N_34568,N_34569,N_34570,N_34571,N_34572,N_34573,N_34574,N_34575,N_34576,N_34577,N_34578,N_34579,N_34580,N_34581,N_34582,N_34583,N_34584,N_34585,N_34586,N_34587,N_34588,N_34589,N_34590,N_34591,N_34592,N_34593,N_34594,N_34595,N_34596,N_34597,N_34598,N_34599,N_34600,N_34601,N_34602,N_34603,N_34604,N_34605,N_34606,N_34607,N_34608,N_34609,N_34610,N_34611,N_34612,N_34613,N_34614,N_34615,N_34616,N_34617,N_34618,N_34619,N_34620,N_34621,N_34622,N_34623,N_34624,N_34625,N_34626,N_34627,N_34628,N_34629,N_34630,N_34631,N_34632,N_34633,N_34634,N_34635,N_34636,N_34637,N_34638,N_34639,N_34640,N_34641,N_34642,N_34643,N_34644,N_34645,N_34646,N_34647,N_34648,N_34649,N_34650,N_34651,N_34652,N_34653,N_34654,N_34655,N_34656,N_34657,N_34658,N_34659,N_34660,N_34661,N_34662,N_34663,N_34664,N_34665,N_34666,N_34667,N_34668,N_34669,N_34670,N_34671,N_34672,N_34673,N_34674,N_34675,N_34676,N_34677,N_34678,N_34679,N_34680,N_34681,N_34682,N_34683,N_34684,N_34685,N_34686,N_34687,N_34688,N_34689,N_34690,N_34691,N_34692,N_34693,N_34694,N_34695,N_34696,N_34697,N_34698,N_34699,N_34700,N_34701,N_34702,N_34703,N_34704,N_34705,N_34706,N_34707,N_34708,N_34709,N_34710,N_34711,N_34712,N_34713,N_34714,N_34715,N_34716,N_34717,N_34718,N_34719,N_34720,N_34721,N_34722,N_34723,N_34724,N_34725,N_34726,N_34727,N_34728,N_34729,N_34730,N_34731,N_34732,N_34733,N_34734,N_34735,N_34736,N_34737,N_34738,N_34739,N_34740,N_34741,N_34742,N_34743,N_34744,N_34745,N_34746,N_34747,N_34748,N_34749,N_34750,N_34751,N_34752,N_34753,N_34754,N_34755,N_34756,N_34757,N_34758,N_34759,N_34760,N_34761,N_34762,N_34763,N_34764,N_34765,N_34766,N_34767,N_34768,N_34769,N_34770,N_34771,N_34772,N_34773,N_34774,N_34775,N_34776,N_34777,N_34778,N_34779,N_34780,N_34781,N_34782,N_34783,N_34784,N_34785,N_34786,N_34787,N_34788,N_34789,N_34790,N_34791,N_34792,N_34793,N_34794,N_34795,N_34796,N_34797,N_34798,N_34799,N_34800,N_34801,N_34802,N_34803,N_34804,N_34805,N_34806,N_34807,N_34808,N_34809,N_34810,N_34811,N_34812,N_34813,N_34814,N_34815,N_34816,N_34817,N_34818,N_34819,N_34820,N_34821,N_34822,N_34823,N_34824,N_34825,N_34826,N_34827,N_34828,N_34829,N_34830,N_34831,N_34832,N_34833,N_34834,N_34835,N_34836,N_34837,N_34838,N_34839,N_34840,N_34841,N_34842,N_34843,N_34844,N_34845,N_34846,N_34847,N_34848,N_34849,N_34850,N_34851,N_34852,N_34853,N_34854,N_34855,N_34856,N_34857,N_34858,N_34859,N_34860,N_34861,N_34862,N_34863,N_34864,N_34865,N_34866,N_34867,N_34868,N_34869,N_34870,N_34871,N_34872,N_34873,N_34874,N_34875,N_34876,N_34877,N_34878,N_34879,N_34880,N_34881,N_34882,N_34883,N_34884,N_34885,N_34886,N_34887,N_34888,N_34889,N_34890,N_34891,N_34892,N_34893,N_34894,N_34895,N_34896,N_34897,N_34898,N_34899,N_34900,N_34901,N_34902,N_34903,N_34904,N_34905,N_34906,N_34907,N_34908,N_34909,N_34910,N_34911,N_34912,N_34913,N_34914,N_34915,N_34916,N_34917,N_34918,N_34919,N_34920,N_34921,N_34922,N_34923,N_34924,N_34925,N_34926,N_34927,N_34928,N_34929,N_34930,N_34931,N_34932,N_34933,N_34934,N_34935,N_34936,N_34937,N_34938,N_34939,N_34940,N_34941,N_34942,N_34943,N_34944,N_34945,N_34946,N_34947,N_34948,N_34949,N_34950,N_34951,N_34952,N_34953,N_34954,N_34955,N_34956,N_34957,N_34958,N_34959,N_34960,N_34961,N_34962,N_34963,N_34964,N_34965,N_34966,N_34967,N_34968,N_34969,N_34970,N_34971,N_34972,N_34973,N_34974,N_34975,N_34976,N_34977,N_34978,N_34979,N_34980,N_34981,N_34982,N_34983,N_34984,N_34985,N_34986,N_34987,N_34988,N_34989,N_34990,N_34991,N_34992,N_34993,N_34994,N_34995,N_34996,N_34997,N_34998,N_34999,N_35000,N_35001,N_35002,N_35003,N_35004,N_35005,N_35006,N_35007,N_35008,N_35009,N_35010,N_35011,N_35012,N_35013,N_35014,N_35015,N_35016,N_35017,N_35018,N_35019,N_35020,N_35021,N_35022,N_35023,N_35024,N_35025,N_35026,N_35027,N_35028,N_35029,N_35030,N_35031,N_35032,N_35033,N_35034,N_35035,N_35036,N_35037,N_35038,N_35039,N_35040,N_35041,N_35042,N_35043,N_35044,N_35045,N_35046,N_35047,N_35048,N_35049,N_35050,N_35051,N_35052,N_35053,N_35054,N_35055,N_35056,N_35057,N_35058,N_35059,N_35060,N_35061,N_35062,N_35063,N_35064,N_35065,N_35066,N_35067,N_35068,N_35069,N_35070,N_35071,N_35072,N_35073,N_35074,N_35075,N_35076,N_35077,N_35078,N_35079,N_35080,N_35081,N_35082,N_35083,N_35084,N_35085,N_35086,N_35087,N_35088,N_35089,N_35090,N_35091,N_35092,N_35093,N_35094,N_35095,N_35096,N_35097,N_35098,N_35099,N_35100,N_35101,N_35102,N_35103,N_35104,N_35105,N_35106,N_35107,N_35108,N_35109,N_35110,N_35111,N_35112,N_35113,N_35114,N_35115,N_35116,N_35117,N_35118,N_35119,N_35120,N_35121,N_35122,N_35123,N_35124,N_35125,N_35126,N_35127,N_35128,N_35129,N_35130,N_35131,N_35132,N_35133,N_35134,N_35135,N_35136,N_35137,N_35138,N_35139,N_35140,N_35141,N_35142,N_35143,N_35144,N_35145,N_35146,N_35147,N_35148,N_35149,N_35150,N_35151,N_35152,N_35153,N_35154,N_35155,N_35156,N_35157,N_35158,N_35159,N_35160,N_35161,N_35162,N_35163,N_35164,N_35165,N_35166,N_35167,N_35168,N_35169,N_35170,N_35171,N_35172,N_35173,N_35174,N_35175,N_35176,N_35177,N_35178,N_35179,N_35180,N_35181,N_35182,N_35183,N_35184,N_35185,N_35186,N_35187,N_35188,N_35189,N_35190,N_35191,N_35192,N_35193,N_35194,N_35195,N_35196,N_35197,N_35198,N_35199,N_35200,N_35201,N_35202,N_35203,N_35204,N_35205,N_35206,N_35207,N_35208,N_35209,N_35210,N_35211,N_35212,N_35213,N_35214,N_35215,N_35216,N_35217,N_35218,N_35219,N_35220,N_35221,N_35222,N_35223,N_35224,N_35225,N_35226,N_35227,N_35228,N_35229,N_35230,N_35231,N_35232,N_35233,N_35234,N_35235,N_35236,N_35237,N_35238,N_35239,N_35240,N_35241,N_35242,N_35243,N_35244,N_35245,N_35246,N_35247,N_35248,N_35249,N_35250,N_35251,N_35252,N_35253,N_35254,N_35255,N_35256,N_35257,N_35258,N_35259,N_35260,N_35261,N_35262,N_35263,N_35264,N_35265,N_35266,N_35267,N_35268,N_35269,N_35270,N_35271,N_35272,N_35273,N_35274,N_35275,N_35276,N_35277,N_35278,N_35279,N_35280,N_35281,N_35282,N_35283,N_35284,N_35285,N_35286,N_35287,N_35288,N_35289,N_35290,N_35291,N_35292,N_35293,N_35294,N_35295,N_35296,N_35297,N_35298,N_35299,N_35300,N_35301,N_35302,N_35303,N_35304,N_35305,N_35306,N_35307,N_35308,N_35309,N_35310,N_35311,N_35312,N_35313,N_35314,N_35315,N_35316,N_35317,N_35318,N_35319,N_35320,N_35321,N_35322,N_35323,N_35324,N_35325,N_35326,N_35327,N_35328,N_35329,N_35330,N_35331,N_35332,N_35333,N_35334,N_35335,N_35336,N_35337,N_35338,N_35339,N_35340,N_35341,N_35342,N_35343,N_35344,N_35345,N_35346,N_35347,N_35348,N_35349,N_35350,N_35351,N_35352,N_35353,N_35354,N_35355,N_35356,N_35357,N_35358,N_35359,N_35360,N_35361,N_35362,N_35363,N_35364,N_35365,N_35366,N_35367,N_35368,N_35369,N_35370,N_35371,N_35372,N_35373,N_35374,N_35375,N_35376,N_35377,N_35378,N_35379,N_35380,N_35381,N_35382,N_35383,N_35384,N_35385,N_35386,N_35387,N_35388,N_35389,N_35390,N_35391,N_35392,N_35393,N_35394,N_35395,N_35396,N_35397,N_35398,N_35399,N_35400,N_35401,N_35402,N_35403,N_35404,N_35405,N_35406,N_35407,N_35408,N_35409,N_35410,N_35411,N_35412,N_35413,N_35414,N_35415,N_35416,N_35417,N_35418,N_35419,N_35420,N_35421,N_35422,N_35423,N_35424,N_35425,N_35426,N_35427,N_35428,N_35429,N_35430,N_35431,N_35432,N_35433,N_35434,N_35435,N_35436,N_35437,N_35438,N_35439,N_35440,N_35441,N_35442,N_35443,N_35444,N_35445,N_35446,N_35447,N_35448,N_35449,N_35450,N_35451,N_35452,N_35453,N_35454,N_35455,N_35456,N_35457,N_35458,N_35459,N_35460,N_35461,N_35462,N_35463,N_35464,N_35465,N_35466,N_35467,N_35468,N_35469,N_35470,N_35471,N_35472,N_35473,N_35474,N_35475,N_35476,N_35477,N_35478,N_35479,N_35480,N_35481,N_35482,N_35483,N_35484,N_35485,N_35486,N_35487,N_35488,N_35489,N_35490,N_35491,N_35492,N_35493,N_35494,N_35495,N_35496,N_35497,N_35498,N_35499,N_35500,N_35501,N_35502,N_35503,N_35504,N_35505,N_35506,N_35507,N_35508,N_35509,N_35510,N_35511,N_35512,N_35513,N_35514,N_35515,N_35516,N_35517,N_35518,N_35519,N_35520,N_35521,N_35522,N_35523,N_35524,N_35525,N_35526,N_35527,N_35528,N_35529,N_35530,N_35531,N_35532,N_35533,N_35534,N_35535,N_35536,N_35537,N_35538,N_35539,N_35540,N_35541,N_35542,N_35543,N_35544,N_35545,N_35546,N_35547,N_35548,N_35549,N_35550,N_35551,N_35552,N_35553,N_35554,N_35555,N_35556,N_35557,N_35558,N_35559,N_35560,N_35561,N_35562,N_35563,N_35564,N_35565,N_35566,N_35567,N_35568,N_35569,N_35570,N_35571,N_35572,N_35573,N_35574,N_35575,N_35576,N_35577,N_35578,N_35579,N_35580,N_35581,N_35582,N_35583,N_35584,N_35585,N_35586,N_35587,N_35588,N_35589,N_35590,N_35591,N_35592,N_35593,N_35594,N_35595,N_35596,N_35597,N_35598,N_35599,N_35600,N_35601,N_35602,N_35603,N_35604,N_35605,N_35606,N_35607,N_35608,N_35609,N_35610,N_35611,N_35612,N_35613,N_35614,N_35615,N_35616,N_35617,N_35618,N_35619,N_35620,N_35621,N_35622,N_35623,N_35624,N_35625,N_35626,N_35627,N_35628,N_35629,N_35630,N_35631,N_35632,N_35633,N_35634,N_35635,N_35636,N_35637,N_35638,N_35639,N_35640,N_35641,N_35642,N_35643,N_35644,N_35645,N_35646,N_35647,N_35648,N_35649,N_35650,N_35651,N_35652,N_35653,N_35654,N_35655,N_35656,N_35657,N_35658,N_35659,N_35660,N_35661,N_35662,N_35663,N_35664,N_35665,N_35666,N_35667,N_35668,N_35669,N_35670,N_35671,N_35672,N_35673,N_35674,N_35675,N_35676,N_35677,N_35678,N_35679,N_35680,N_35681,N_35682,N_35683,N_35684,N_35685,N_35686,N_35687,N_35688,N_35689,N_35690,N_35691,N_35692,N_35693,N_35694,N_35695,N_35696,N_35697,N_35698,N_35699,N_35700,N_35701,N_35702,N_35703,N_35704,N_35705,N_35706,N_35707,N_35708,N_35709,N_35710,N_35711,N_35712,N_35713,N_35714,N_35715,N_35716,N_35717,N_35718,N_35719,N_35720,N_35721,N_35722,N_35723,N_35724,N_35725,N_35726,N_35727,N_35728,N_35729,N_35730,N_35731,N_35732,N_35733,N_35734,N_35735,N_35736,N_35737,N_35738,N_35739,N_35740,N_35741,N_35742,N_35743,N_35744,N_35745,N_35746,N_35747,N_35748,N_35749,N_35750,N_35751,N_35752,N_35753,N_35754,N_35755,N_35756,N_35757,N_35758,N_35759,N_35760,N_35761,N_35762,N_35763,N_35764,N_35765,N_35766,N_35767,N_35768,N_35769,N_35770,N_35771,N_35772,N_35773,N_35774,N_35775,N_35776,N_35777,N_35778,N_35779,N_35780,N_35781,N_35782,N_35783,N_35784,N_35785,N_35786,N_35787,N_35788,N_35789,N_35790,N_35791,N_35792,N_35793,N_35794,N_35795,N_35796,N_35797,N_35798,N_35799,N_35800,N_35801,N_35802,N_35803,N_35804,N_35805,N_35806,N_35807,N_35808,N_35809,N_35810,N_35811,N_35812,N_35813,N_35814,N_35815,N_35816,N_35817,N_35818,N_35819,N_35820,N_35821,N_35822,N_35823,N_35824,N_35825,N_35826,N_35827,N_35828,N_35829,N_35830,N_35831,N_35832,N_35833,N_35834,N_35835,N_35836,N_35837,N_35838,N_35839,N_35840,N_35841,N_35842,N_35843,N_35844,N_35845,N_35846,N_35847,N_35848,N_35849,N_35850,N_35851,N_35852,N_35853,N_35854,N_35855,N_35856,N_35857,N_35858,N_35859,N_35860,N_35861,N_35862,N_35863,N_35864,N_35865,N_35866,N_35867,N_35868,N_35869,N_35870,N_35871,N_35872,N_35873,N_35874,N_35875,N_35876,N_35877,N_35878,N_35879,N_35880,N_35881,N_35882,N_35883,N_35884,N_35885,N_35886,N_35887,N_35888,N_35889,N_35890,N_35891,N_35892,N_35893,N_35894,N_35895,N_35896,N_35897,N_35898,N_35899,N_35900,N_35901,N_35902,N_35903,N_35904,N_35905,N_35906,N_35907,N_35908,N_35909,N_35910,N_35911,N_35912,N_35913,N_35914,N_35915,N_35916,N_35917,N_35918,N_35919,N_35920,N_35921,N_35922,N_35923,N_35924,N_35925,N_35926,N_35927,N_35928,N_35929,N_35930,N_35931,N_35932,N_35933,N_35934,N_35935,N_35936,N_35937,N_35938,N_35939,N_35940,N_35941,N_35942,N_35943,N_35944,N_35945,N_35946,N_35947,N_35948,N_35949,N_35950,N_35951,N_35952,N_35953,N_35954,N_35955,N_35956,N_35957,N_35958,N_35959,N_35960,N_35961,N_35962,N_35963,N_35964,N_35965,N_35966,N_35967,N_35968,N_35969,N_35970,N_35971,N_35972,N_35973,N_35974,N_35975,N_35976,N_35977,N_35978,N_35979,N_35980,N_35981,N_35982,N_35983,N_35984,N_35985,N_35986,N_35987,N_35988,N_35989,N_35990,N_35991,N_35992,N_35993,N_35994,N_35995,N_35996,N_35997,N_35998,N_35999,N_36000,N_36001,N_36002,N_36003,N_36004,N_36005,N_36006,N_36007,N_36008,N_36009,N_36010,N_36011,N_36012,N_36013,N_36014,N_36015,N_36016,N_36017,N_36018,N_36019,N_36020,N_36021,N_36022,N_36023,N_36024,N_36025,N_36026,N_36027,N_36028,N_36029,N_36030,N_36031,N_36032,N_36033,N_36034,N_36035,N_36036,N_36037,N_36038,N_36039,N_36040,N_36041,N_36042,N_36043,N_36044,N_36045,N_36046,N_36047,N_36048,N_36049,N_36050,N_36051,N_36052,N_36053,N_36054,N_36055,N_36056,N_36057,N_36058,N_36059,N_36060,N_36061,N_36062,N_36063,N_36064,N_36065,N_36066,N_36067,N_36068,N_36069,N_36070,N_36071,N_36072,N_36073,N_36074,N_36075,N_36076,N_36077,N_36078,N_36079,N_36080,N_36081,N_36082,N_36083,N_36084,N_36085,N_36086,N_36087,N_36088,N_36089,N_36090,N_36091,N_36092,N_36093,N_36094,N_36095,N_36096,N_36097,N_36098,N_36099,N_36100,N_36101,N_36102,N_36103,N_36104,N_36105,N_36106,N_36107,N_36108,N_36109,N_36110,N_36111,N_36112,N_36113,N_36114,N_36115,N_36116,N_36117,N_36118,N_36119,N_36120,N_36121,N_36122,N_36123,N_36124,N_36125,N_36126,N_36127,N_36128,N_36129,N_36130,N_36131,N_36132,N_36133,N_36134,N_36135,N_36136,N_36137,N_36138,N_36139,N_36140,N_36141,N_36142,N_36143,N_36144,N_36145,N_36146,N_36147,N_36148,N_36149,N_36150,N_36151,N_36152,N_36153,N_36154,N_36155,N_36156,N_36157,N_36158,N_36159,N_36160,N_36161,N_36162,N_36163,N_36164,N_36165,N_36166,N_36167,N_36168,N_36169,N_36170,N_36171,N_36172,N_36173,N_36174,N_36175,N_36176,N_36177,N_36178,N_36179,N_36180,N_36181,N_36182,N_36183,N_36184,N_36185,N_36186,N_36187,N_36188,N_36189,N_36190,N_36191,N_36192,N_36193,N_36194,N_36195,N_36196,N_36197,N_36198,N_36199,N_36200,N_36201,N_36202,N_36203,N_36204,N_36205,N_36206,N_36207,N_36208,N_36209,N_36210,N_36211,N_36212,N_36213,N_36214,N_36215,N_36216,N_36217,N_36218,N_36219,N_36220,N_36221,N_36222,N_36223,N_36224,N_36225,N_36226,N_36227,N_36228,N_36229,N_36230,N_36231,N_36232,N_36233,N_36234,N_36235,N_36236,N_36237,N_36238,N_36239,N_36240,N_36241,N_36242,N_36243,N_36244,N_36245,N_36246,N_36247,N_36248,N_36249,N_36250,N_36251,N_36252,N_36253,N_36254,N_36255,N_36256,N_36257,N_36258,N_36259,N_36260,N_36261,N_36262,N_36263,N_36264,N_36265,N_36266,N_36267,N_36268,N_36269,N_36270,N_36271,N_36272,N_36273,N_36274,N_36275,N_36276,N_36277,N_36278,N_36279,N_36280,N_36281,N_36282,N_36283,N_36284,N_36285,N_36286,N_36287,N_36288,N_36289,N_36290,N_36291,N_36292,N_36293,N_36294,N_36295,N_36296,N_36297,N_36298,N_36299,N_36300,N_36301,N_36302,N_36303,N_36304,N_36305,N_36306,N_36307,N_36308,N_36309,N_36310,N_36311,N_36312,N_36313,N_36314,N_36315,N_36316,N_36317,N_36318,N_36319,N_36320,N_36321,N_36322,N_36323,N_36324,N_36325,N_36326,N_36327,N_36328,N_36329,N_36330,N_36331,N_36332,N_36333,N_36334,N_36335,N_36336,N_36337,N_36338,N_36339,N_36340,N_36341,N_36342,N_36343,N_36344,N_36345,N_36346,N_36347,N_36348,N_36349,N_36350,N_36351,N_36352,N_36353,N_36354,N_36355,N_36356,N_36357,N_36358,N_36359,N_36360,N_36361,N_36362,N_36363,N_36364,N_36365,N_36366,N_36367,N_36368,N_36369,N_36370,N_36371,N_36372,N_36373,N_36374,N_36375,N_36376,N_36377,N_36378,N_36379,N_36380,N_36381,N_36382,N_36383,N_36384,N_36385,N_36386,N_36387,N_36388,N_36389,N_36390,N_36391,N_36392,N_36393,N_36394,N_36395,N_36396,N_36397,N_36398,N_36399,N_36400,N_36401,N_36402,N_36403,N_36404,N_36405,N_36406,N_36407,N_36408,N_36409,N_36410,N_36411,N_36412,N_36413,N_36414,N_36415,N_36416,N_36417,N_36418,N_36419,N_36420,N_36421,N_36422,N_36423,N_36424,N_36425,N_36426,N_36427,N_36428,N_36429,N_36430,N_36431,N_36432,N_36433,N_36434,N_36435,N_36436,N_36437,N_36438,N_36439,N_36440,N_36441,N_36442,N_36443,N_36444,N_36445,N_36446,N_36447,N_36448,N_36449,N_36450,N_36451,N_36452,N_36453,N_36454,N_36455,N_36456,N_36457,N_36458,N_36459,N_36460,N_36461,N_36462,N_36463,N_36464,N_36465,N_36466,N_36467,N_36468,N_36469,N_36470,N_36471,N_36472,N_36473,N_36474,N_36475,N_36476,N_36477,N_36478,N_36479,N_36480,N_36481,N_36482,N_36483,N_36484,N_36485,N_36486,N_36487,N_36488,N_36489,N_36490,N_36491,N_36492,N_36493,N_36494,N_36495,N_36496,N_36497,N_36498,N_36499,N_36500,N_36501,N_36502,N_36503,N_36504,N_36505,N_36506,N_36507,N_36508,N_36509,N_36510,N_36511,N_36512,N_36513,N_36514,N_36515,N_36516,N_36517,N_36518,N_36519,N_36520,N_36521,N_36522,N_36523,N_36524,N_36525,N_36526,N_36527,N_36528,N_36529,N_36530,N_36531,N_36532,N_36533,N_36534,N_36535,N_36536,N_36537,N_36538,N_36539,N_36540,N_36541,N_36542,N_36543,N_36544,N_36545,N_36546,N_36547,N_36548,N_36549,N_36550,N_36551,N_36552,N_36553,N_36554,N_36555,N_36556,N_36557,N_36558,N_36559,N_36560,N_36561,N_36562,N_36563,N_36564,N_36565,N_36566,N_36567,N_36568,N_36569,N_36570,N_36571,N_36572,N_36573,N_36574,N_36575,N_36576,N_36577,N_36578,N_36579,N_36580,N_36581,N_36582,N_36583,N_36584,N_36585,N_36586,N_36587,N_36588,N_36589,N_36590,N_36591,N_36592,N_36593,N_36594,N_36595,N_36596,N_36597,N_36598,N_36599,N_36600,N_36601,N_36602,N_36603,N_36604,N_36605,N_36606,N_36607,N_36608,N_36609,N_36610,N_36611,N_36612,N_36613,N_36614,N_36615,N_36616,N_36617,N_36618,N_36619,N_36620,N_36621,N_36622,N_36623,N_36624,N_36625,N_36626,N_36627,N_36628,N_36629,N_36630,N_36631,N_36632,N_36633,N_36634,N_36635,N_36636,N_36637,N_36638,N_36639,N_36640,N_36641,N_36642,N_36643,N_36644,N_36645,N_36646,N_36647,N_36648,N_36649,N_36650,N_36651,N_36652,N_36653,N_36654,N_36655,N_36656,N_36657,N_36658,N_36659,N_36660,N_36661,N_36662,N_36663,N_36664,N_36665,N_36666,N_36667,N_36668,N_36669,N_36670,N_36671,N_36672,N_36673,N_36674,N_36675,N_36676,N_36677,N_36678,N_36679,N_36680,N_36681,N_36682,N_36683,N_36684,N_36685,N_36686,N_36687,N_36688,N_36689,N_36690,N_36691,N_36692,N_36693,N_36694,N_36695,N_36696,N_36697,N_36698,N_36699,N_36700,N_36701,N_36702,N_36703,N_36704,N_36705,N_36706,N_36707,N_36708,N_36709,N_36710,N_36711,N_36712,N_36713,N_36714,N_36715,N_36716,N_36717,N_36718,N_36719,N_36720,N_36721,N_36722,N_36723,N_36724,N_36725,N_36726,N_36727,N_36728,N_36729,N_36730,N_36731,N_36732,N_36733,N_36734,N_36735,N_36736,N_36737,N_36738,N_36739,N_36740,N_36741,N_36742,N_36743,N_36744,N_36745,N_36746,N_36747,N_36748,N_36749,N_36750,N_36751,N_36752,N_36753,N_36754,N_36755,N_36756,N_36757,N_36758,N_36759,N_36760,N_36761,N_36762,N_36763,N_36764,N_36765,N_36766,N_36767,N_36768,N_36769,N_36770,N_36771,N_36772,N_36773,N_36774,N_36775,N_36776,N_36777,N_36778,N_36779,N_36780,N_36781,N_36782,N_36783,N_36784,N_36785,N_36786,N_36787,N_36788,N_36789,N_36790,N_36791,N_36792,N_36793,N_36794,N_36795,N_36796,N_36797,N_36798,N_36799,N_36800,N_36801,N_36802,N_36803,N_36804,N_36805,N_36806,N_36807,N_36808,N_36809,N_36810,N_36811,N_36812,N_36813,N_36814,N_36815,N_36816,N_36817,N_36818,N_36819,N_36820,N_36821,N_36822,N_36823,N_36824,N_36825,N_36826,N_36827,N_36828,N_36829,N_36830,N_36831,N_36832,N_36833,N_36834,N_36835,N_36836,N_36837,N_36838,N_36839,N_36840,N_36841,N_36842,N_36843,N_36844,N_36845,N_36846,N_36847,N_36848,N_36849,N_36850,N_36851,N_36852,N_36853,N_36854,N_36855,N_36856,N_36857,N_36858,N_36859,N_36860,N_36861,N_36862,N_36863,N_36864,N_36865,N_36866,N_36867,N_36868,N_36869,N_36870,N_36871,N_36872,N_36873,N_36874,N_36875,N_36876,N_36877,N_36878,N_36879,N_36880,N_36881,N_36882,N_36883,N_36884,N_36885,N_36886,N_36887,N_36888,N_36889,N_36890,N_36891,N_36892,N_36893,N_36894,N_36895,N_36896,N_36897,N_36898,N_36899,N_36900,N_36901,N_36902,N_36903,N_36904,N_36905,N_36906,N_36907,N_36908,N_36909,N_36910,N_36911,N_36912,N_36913,N_36914,N_36915,N_36916,N_36917,N_36918,N_36919,N_36920,N_36921,N_36922,N_36923,N_36924,N_36925,N_36926,N_36927,N_36928,N_36929,N_36930,N_36931,N_36932,N_36933,N_36934,N_36935,N_36936,N_36937,N_36938,N_36939,N_36940,N_36941,N_36942,N_36943,N_36944,N_36945,N_36946,N_36947,N_36948,N_36949,N_36950,N_36951,N_36952,N_36953,N_36954,N_36955,N_36956,N_36957,N_36958,N_36959,N_36960,N_36961,N_36962,N_36963,N_36964,N_36965,N_36966,N_36967,N_36968,N_36969,N_36970,N_36971,N_36972,N_36973,N_36974,N_36975,N_36976,N_36977,N_36978,N_36979,N_36980,N_36981,N_36982,N_36983,N_36984,N_36985,N_36986,N_36987,N_36988,N_36989,N_36990,N_36991,N_36992,N_36993,N_36994,N_36995,N_36996,N_36997,N_36998,N_36999,N_37000,N_37001,N_37002,N_37003,N_37004,N_37005,N_37006,N_37007,N_37008,N_37009,N_37010,N_37011,N_37012,N_37013,N_37014,N_37015,N_37016,N_37017,N_37018,N_37019,N_37020,N_37021,N_37022,N_37023,N_37024,N_37025,N_37026,N_37027,N_37028,N_37029,N_37030,N_37031,N_37032,N_37033,N_37034,N_37035,N_37036,N_37037,N_37038,N_37039,N_37040,N_37041,N_37042,N_37043,N_37044,N_37045,N_37046,N_37047,N_37048,N_37049,N_37050,N_37051,N_37052,N_37053,N_37054,N_37055,N_37056,N_37057,N_37058,N_37059,N_37060,N_37061,N_37062,N_37063,N_37064,N_37065,N_37066,N_37067,N_37068,N_37069,N_37070,N_37071,N_37072,N_37073,N_37074,N_37075,N_37076,N_37077,N_37078,N_37079,N_37080,N_37081,N_37082,N_37083,N_37084,N_37085,N_37086,N_37087,N_37088,N_37089,N_37090,N_37091,N_37092,N_37093,N_37094,N_37095,N_37096,N_37097,N_37098,N_37099,N_37100,N_37101,N_37102,N_37103,N_37104,N_37105,N_37106,N_37107,N_37108,N_37109,N_37110,N_37111,N_37112,N_37113,N_37114,N_37115,N_37116,N_37117,N_37118,N_37119,N_37120,N_37121,N_37122,N_37123,N_37124,N_37125,N_37126,N_37127,N_37128,N_37129,N_37130,N_37131,N_37132,N_37133,N_37134,N_37135,N_37136,N_37137,N_37138,N_37139,N_37140,N_37141,N_37142,N_37143,N_37144,N_37145,N_37146,N_37147,N_37148,N_37149,N_37150,N_37151,N_37152,N_37153,N_37154,N_37155,N_37156,N_37157,N_37158,N_37159,N_37160,N_37161,N_37162,N_37163,N_37164,N_37165,N_37166,N_37167,N_37168,N_37169,N_37170,N_37171,N_37172,N_37173,N_37174,N_37175,N_37176,N_37177,N_37178,N_37179,N_37180,N_37181,N_37182,N_37183,N_37184,N_37185,N_37186,N_37187,N_37188,N_37189,N_37190,N_37191,N_37192,N_37193,N_37194,N_37195,N_37196,N_37197,N_37198,N_37199,N_37200,N_37201,N_37202,N_37203,N_37204,N_37205,N_37206,N_37207,N_37208,N_37209,N_37210,N_37211,N_37212,N_37213,N_37214,N_37215,N_37216,N_37217,N_37218,N_37219,N_37220,N_37221,N_37222,N_37223,N_37224,N_37225,N_37226,N_37227,N_37228,N_37229,N_37230,N_37231,N_37232,N_37233,N_37234,N_37235,N_37236,N_37237,N_37238,N_37239,N_37240,N_37241,N_37242,N_37243,N_37244,N_37245,N_37246,N_37247,N_37248,N_37249,N_37250,N_37251,N_37252,N_37253,N_37254,N_37255,N_37256,N_37257,N_37258,N_37259,N_37260,N_37261,N_37262,N_37263,N_37264,N_37265,N_37266,N_37267,N_37268,N_37269,N_37270,N_37271,N_37272,N_37273,N_37274,N_37275,N_37276,N_37277,N_37278,N_37279,N_37280,N_37281,N_37282,N_37283,N_37284,N_37285,N_37286,N_37287,N_37288,N_37289,N_37290,N_37291,N_37292,N_37293,N_37294,N_37295,N_37296,N_37297,N_37298,N_37299,N_37300,N_37301,N_37302,N_37303,N_37304,N_37305,N_37306,N_37307,N_37308,N_37309,N_37310,N_37311,N_37312,N_37313,N_37314,N_37315,N_37316,N_37317,N_37318,N_37319,N_37320,N_37321,N_37322,N_37323,N_37324,N_37325,N_37326,N_37327,N_37328,N_37329,N_37330,N_37331,N_37332,N_37333,N_37334,N_37335,N_37336,N_37337,N_37338,N_37339,N_37340,N_37341,N_37342,N_37343,N_37344,N_37345,N_37346,N_37347,N_37348,N_37349,N_37350,N_37351,N_37352,N_37353,N_37354,N_37355,N_37356,N_37357,N_37358,N_37359,N_37360,N_37361,N_37362,N_37363,N_37364,N_37365,N_37366,N_37367,N_37368,N_37369,N_37370,N_37371,N_37372,N_37373,N_37374,N_37375,N_37376,N_37377,N_37378,N_37379,N_37380,N_37381,N_37382,N_37383,N_37384,N_37385,N_37386,N_37387,N_37388,N_37389,N_37390,N_37391,N_37392,N_37393,N_37394,N_37395,N_37396,N_37397,N_37398,N_37399,N_37400,N_37401,N_37402,N_37403,N_37404,N_37405,N_37406,N_37407,N_37408,N_37409,N_37410,N_37411,N_37412,N_37413,N_37414,N_37415,N_37416,N_37417,N_37418,N_37419,N_37420,N_37421,N_37422,N_37423,N_37424,N_37425,N_37426,N_37427,N_37428,N_37429,N_37430,N_37431,N_37432,N_37433,N_37434,N_37435,N_37436,N_37437,N_37438,N_37439,N_37440,N_37441,N_37442,N_37443,N_37444,N_37445,N_37446,N_37447,N_37448,N_37449,N_37450,N_37451,N_37452,N_37453,N_37454,N_37455,N_37456,N_37457,N_37458,N_37459,N_37460,N_37461,N_37462,N_37463,N_37464,N_37465,N_37466,N_37467,N_37468,N_37469,N_37470,N_37471,N_37472,N_37473,N_37474,N_37475,N_37476,N_37477,N_37478,N_37479,N_37480,N_37481,N_37482,N_37483,N_37484,N_37485,N_37486,N_37487,N_37488,N_37489,N_37490,N_37491,N_37492,N_37493,N_37494,N_37495,N_37496,N_37497,N_37498,N_37499,N_37500,N_37501,N_37502,N_37503,N_37504,N_37505,N_37506,N_37507,N_37508,N_37509,N_37510,N_37511,N_37512,N_37513,N_37514,N_37515,N_37516,N_37517,N_37518,N_37519,N_37520,N_37521,N_37522,N_37523,N_37524,N_37525,N_37526,N_37527,N_37528,N_37529,N_37530,N_37531,N_37532,N_37533,N_37534,N_37535,N_37536,N_37537,N_37538,N_37539,N_37540,N_37541,N_37542,N_37543,N_37544,N_37545,N_37546,N_37547,N_37548,N_37549,N_37550,N_37551,N_37552,N_37553,N_37554,N_37555,N_37556,N_37557,N_37558,N_37559,N_37560,N_37561,N_37562,N_37563,N_37564,N_37565,N_37566,N_37567,N_37568,N_37569,N_37570,N_37571,N_37572,N_37573,N_37574,N_37575,N_37576,N_37577,N_37578,N_37579,N_37580,N_37581,N_37582,N_37583,N_37584,N_37585,N_37586,N_37587,N_37588,N_37589,N_37590,N_37591,N_37592,N_37593,N_37594,N_37595,N_37596,N_37597,N_37598,N_37599,N_37600,N_37601,N_37602,N_37603,N_37604,N_37605,N_37606,N_37607,N_37608,N_37609,N_37610,N_37611,N_37612,N_37613,N_37614,N_37615,N_37616,N_37617,N_37618,N_37619,N_37620,N_37621,N_37622,N_37623,N_37624,N_37625,N_37626,N_37627,N_37628,N_37629,N_37630,N_37631,N_37632,N_37633,N_37634,N_37635,N_37636,N_37637,N_37638,N_37639,N_37640,N_37641,N_37642,N_37643,N_37644,N_37645,N_37646,N_37647,N_37648,N_37649,N_37650,N_37651,N_37652,N_37653,N_37654,N_37655,N_37656,N_37657,N_37658,N_37659,N_37660,N_37661,N_37662,N_37663,N_37664,N_37665,N_37666,N_37667,N_37668,N_37669,N_37670,N_37671,N_37672,N_37673,N_37674,N_37675,N_37676,N_37677,N_37678,N_37679,N_37680,N_37681,N_37682,N_37683,N_37684,N_37685,N_37686,N_37687,N_37688,N_37689,N_37690,N_37691,N_37692,N_37693,N_37694,N_37695,N_37696,N_37697,N_37698,N_37699,N_37700,N_37701,N_37702,N_37703,N_37704,N_37705,N_37706,N_37707,N_37708,N_37709,N_37710,N_37711,N_37712,N_37713,N_37714,N_37715,N_37716,N_37717,N_37718,N_37719,N_37720,N_37721,N_37722,N_37723,N_37724,N_37725,N_37726,N_37727,N_37728,N_37729,N_37730,N_37731,N_37732,N_37733,N_37734,N_37735,N_37736,N_37737,N_37738,N_37739,N_37740,N_37741,N_37742,N_37743,N_37744,N_37745,N_37746,N_37747,N_37748,N_37749,N_37750,N_37751,N_37752,N_37753,N_37754,N_37755,N_37756,N_37757,N_37758,N_37759,N_37760,N_37761,N_37762,N_37763,N_37764,N_37765,N_37766,N_37767,N_37768,N_37769,N_37770,N_37771,N_37772,N_37773,N_37774,N_37775,N_37776,N_37777,N_37778,N_37779,N_37780,N_37781,N_37782,N_37783,N_37784,N_37785,N_37786,N_37787,N_37788,N_37789,N_37790,N_37791,N_37792,N_37793,N_37794,N_37795,N_37796,N_37797,N_37798,N_37799,N_37800,N_37801,N_37802,N_37803,N_37804,N_37805,N_37806,N_37807,N_37808,N_37809,N_37810,N_37811,N_37812,N_37813,N_37814,N_37815,N_37816,N_37817,N_37818,N_37819,N_37820,N_37821,N_37822,N_37823,N_37824,N_37825,N_37826,N_37827,N_37828,N_37829,N_37830,N_37831,N_37832,N_37833,N_37834,N_37835,N_37836,N_37837,N_37838,N_37839,N_37840,N_37841,N_37842,N_37843,N_37844,N_37845,N_37846,N_37847,N_37848,N_37849,N_37850,N_37851,N_37852,N_37853,N_37854,N_37855,N_37856,N_37857,N_37858,N_37859,N_37860,N_37861,N_37862,N_37863,N_37864,N_37865,N_37866,N_37867,N_37868,N_37869,N_37870,N_37871,N_37872,N_37873,N_37874,N_37875,N_37876,N_37877,N_37878,N_37879,N_37880,N_37881,N_37882,N_37883,N_37884,N_37885,N_37886,N_37887,N_37888,N_37889,N_37890,N_37891,N_37892,N_37893,N_37894,N_37895,N_37896,N_37897,N_37898,N_37899,N_37900,N_37901,N_37902,N_37903,N_37904,N_37905,N_37906,N_37907,N_37908,N_37909,N_37910,N_37911,N_37912,N_37913,N_37914,N_37915,N_37916,N_37917,N_37918,N_37919,N_37920,N_37921,N_37922,N_37923,N_37924,N_37925,N_37926,N_37927,N_37928,N_37929,N_37930,N_37931,N_37932,N_37933,N_37934,N_37935,N_37936,N_37937,N_37938,N_37939,N_37940,N_37941,N_37942,N_37943,N_37944,N_37945,N_37946,N_37947,N_37948,N_37949,N_37950,N_37951,N_37952,N_37953,N_37954,N_37955,N_37956,N_37957,N_37958,N_37959,N_37960,N_37961,N_37962,N_37963,N_37964,N_37965,N_37966,N_37967,N_37968,N_37969,N_37970,N_37971,N_37972,N_37973,N_37974,N_37975,N_37976,N_37977,N_37978,N_37979,N_37980,N_37981,N_37982,N_37983,N_37984,N_37985,N_37986,N_37987,N_37988,N_37989,N_37990,N_37991,N_37992,N_37993,N_37994,N_37995,N_37996,N_37997,N_37998,N_37999,N_38000,N_38001,N_38002,N_38003,N_38004,N_38005,N_38006,N_38007,N_38008,N_38009,N_38010,N_38011,N_38012,N_38013,N_38014,N_38015,N_38016,N_38017,N_38018,N_38019,N_38020,N_38021,N_38022,N_38023,N_38024,N_38025,N_38026,N_38027,N_38028,N_38029,N_38030,N_38031,N_38032,N_38033,N_38034,N_38035,N_38036,N_38037,N_38038,N_38039,N_38040,N_38041,N_38042,N_38043,N_38044,N_38045,N_38046,N_38047,N_38048,N_38049,N_38050,N_38051,N_38052,N_38053,N_38054,N_38055,N_38056,N_38057,N_38058,N_38059,N_38060,N_38061,N_38062,N_38063,N_38064,N_38065,N_38066,N_38067,N_38068,N_38069,N_38070,N_38071,N_38072,N_38073,N_38074,N_38075,N_38076,N_38077,N_38078,N_38079,N_38080,N_38081,N_38082,N_38083,N_38084,N_38085,N_38086,N_38087,N_38088,N_38089,N_38090,N_38091,N_38092,N_38093,N_38094,N_38095,N_38096,N_38097,N_38098,N_38099,N_38100,N_38101,N_38102,N_38103,N_38104,N_38105,N_38106,N_38107,N_38108,N_38109,N_38110,N_38111,N_38112,N_38113,N_38114,N_38115,N_38116,N_38117,N_38118,N_38119,N_38120,N_38121,N_38122,N_38123,N_38124,N_38125,N_38126,N_38127,N_38128,N_38129,N_38130,N_38131,N_38132,N_38133,N_38134,N_38135,N_38136,N_38137,N_38138,N_38139,N_38140,N_38141,N_38142,N_38143,N_38144,N_38145,N_38146,N_38147,N_38148,N_38149,N_38150,N_38151,N_38152,N_38153,N_38154,N_38155,N_38156,N_38157,N_38158,N_38159,N_38160,N_38161,N_38162,N_38163,N_38164,N_38165,N_38166,N_38167,N_38168,N_38169,N_38170,N_38171,N_38172,N_38173,N_38174,N_38175,N_38176,N_38177,N_38178,N_38179,N_38180,N_38181,N_38182,N_38183,N_38184,N_38185,N_38186,N_38187,N_38188,N_38189,N_38190,N_38191,N_38192,N_38193,N_38194,N_38195,N_38196,N_38197,N_38198,N_38199,N_38200,N_38201,N_38202,N_38203,N_38204,N_38205,N_38206,N_38207,N_38208,N_38209,N_38210,N_38211,N_38212,N_38213,N_38214,N_38215,N_38216,N_38217,N_38218,N_38219,N_38220,N_38221,N_38222,N_38223,N_38224,N_38225,N_38226,N_38227,N_38228,N_38229,N_38230,N_38231,N_38232,N_38233,N_38234,N_38235,N_38236,N_38237,N_38238,N_38239,N_38240,N_38241,N_38242,N_38243,N_38244,N_38245,N_38246,N_38247,N_38248,N_38249,N_38250,N_38251,N_38252,N_38253,N_38254,N_38255,N_38256,N_38257,N_38258,N_38259,N_38260,N_38261,N_38262,N_38263,N_38264,N_38265,N_38266,N_38267,N_38268,N_38269,N_38270,N_38271,N_38272,N_38273,N_38274,N_38275,N_38276,N_38277,N_38278,N_38279,N_38280,N_38281,N_38282,N_38283,N_38284,N_38285,N_38286,N_38287,N_38288,N_38289,N_38290,N_38291,N_38292,N_38293,N_38294,N_38295,N_38296,N_38297,N_38298,N_38299,N_38300,N_38301,N_38302,N_38303,N_38304,N_38305,N_38306,N_38307,N_38308,N_38309,N_38310,N_38311,N_38312,N_38313,N_38314,N_38315,N_38316,N_38317,N_38318,N_38319,N_38320,N_38321,N_38322,N_38323,N_38324,N_38325,N_38326,N_38327,N_38328,N_38329,N_38330,N_38331,N_38332,N_38333,N_38334,N_38335,N_38336,N_38337,N_38338,N_38339,N_38340,N_38341,N_38342,N_38343,N_38344,N_38345,N_38346,N_38347,N_38348,N_38349,N_38350,N_38351,N_38352,N_38353,N_38354,N_38355,N_38356,N_38357,N_38358,N_38359,N_38360,N_38361,N_38362,N_38363,N_38364,N_38365,N_38366,N_38367,N_38368,N_38369,N_38370,N_38371,N_38372,N_38373,N_38374,N_38375,N_38376,N_38377,N_38378,N_38379,N_38380,N_38381,N_38382,N_38383,N_38384,N_38385,N_38386,N_38387,N_38388,N_38389,N_38390,N_38391,N_38392,N_38393,N_38394,N_38395,N_38396,N_38397,N_38398,N_38399,N_38400,N_38401,N_38402,N_38403,N_38404,N_38405,N_38406,N_38407,N_38408,N_38409,N_38410,N_38411,N_38412,N_38413,N_38414,N_38415,N_38416,N_38417,N_38418,N_38419,N_38420,N_38421,N_38422,N_38423,N_38424,N_38425,N_38426,N_38427,N_38428,N_38429,N_38430,N_38431,N_38432,N_38433,N_38434,N_38435,N_38436,N_38437,N_38438,N_38439,N_38440,N_38441,N_38442,N_38443,N_38444,N_38445,N_38446,N_38447,N_38448,N_38449,N_38450,N_38451,N_38452,N_38453,N_38454,N_38455,N_38456,N_38457,N_38458,N_38459,N_38460,N_38461,N_38462,N_38463,N_38464,N_38465,N_38466,N_38467,N_38468,N_38469,N_38470,N_38471,N_38472,N_38473,N_38474,N_38475,N_38476,N_38477,N_38478,N_38479,N_38480,N_38481,N_38482,N_38483,N_38484,N_38485,N_38486,N_38487,N_38488,N_38489,N_38490,N_38491,N_38492,N_38493,N_38494,N_38495,N_38496,N_38497,N_38498,N_38499,N_38500,N_38501,N_38502,N_38503,N_38504,N_38505,N_38506,N_38507,N_38508,N_38509,N_38510,N_38511,N_38512,N_38513,N_38514,N_38515,N_38516,N_38517,N_38518,N_38519,N_38520,N_38521,N_38522,N_38523,N_38524,N_38525,N_38526,N_38527,N_38528,N_38529,N_38530,N_38531,N_38532,N_38533,N_38534,N_38535,N_38536,N_38537,N_38538,N_38539,N_38540,N_38541,N_38542,N_38543,N_38544,N_38545,N_38546,N_38547,N_38548,N_38549,N_38550,N_38551,N_38552,N_38553,N_38554,N_38555,N_38556,N_38557,N_38558,N_38559,N_38560,N_38561,N_38562,N_38563,N_38564,N_38565,N_38566,N_38567,N_38568,N_38569,N_38570,N_38571,N_38572,N_38573,N_38574,N_38575,N_38576,N_38577,N_38578,N_38579,N_38580,N_38581,N_38582,N_38583,N_38584,N_38585,N_38586,N_38587,N_38588,N_38589,N_38590,N_38591,N_38592,N_38593,N_38594,N_38595,N_38596,N_38597,N_38598,N_38599,N_38600,N_38601,N_38602,N_38603,N_38604,N_38605,N_38606,N_38607,N_38608,N_38609,N_38610,N_38611,N_38612,N_38613,N_38614,N_38615,N_38616,N_38617,N_38618,N_38619,N_38620,N_38621,N_38622,N_38623,N_38624,N_38625,N_38626,N_38627,N_38628,N_38629,N_38630,N_38631,N_38632,N_38633,N_38634,N_38635,N_38636,N_38637,N_38638,N_38639,N_38640,N_38641,N_38642,N_38643,N_38644,N_38645,N_38646,N_38647,N_38648,N_38649,N_38650,N_38651,N_38652,N_38653,N_38654,N_38655,N_38656,N_38657,N_38658,N_38659,N_38660,N_38661,N_38662,N_38663,N_38664,N_38665,N_38666,N_38667,N_38668,N_38669,N_38670,N_38671,N_38672,N_38673,N_38674,N_38675,N_38676,N_38677,N_38678,N_38679,N_38680,N_38681,N_38682,N_38683,N_38684,N_38685,N_38686,N_38687,N_38688,N_38689,N_38690,N_38691,N_38692,N_38693,N_38694,N_38695,N_38696,N_38697,N_38698,N_38699,N_38700,N_38701,N_38702,N_38703,N_38704,N_38705,N_38706,N_38707,N_38708,N_38709,N_38710,N_38711,N_38712,N_38713,N_38714,N_38715,N_38716,N_38717,N_38718,N_38719,N_38720,N_38721,N_38722,N_38723,N_38724,N_38725,N_38726,N_38727,N_38728,N_38729,N_38730,N_38731,N_38732,N_38733,N_38734,N_38735,N_38736,N_38737,N_38738,N_38739,N_38740,N_38741,N_38742,N_38743,N_38744,N_38745,N_38746,N_38747,N_38748,N_38749,N_38750,N_38751,N_38752,N_38753,N_38754,N_38755,N_38756,N_38757,N_38758,N_38759,N_38760,N_38761,N_38762,N_38763,N_38764,N_38765,N_38766,N_38767,N_38768,N_38769,N_38770,N_38771,N_38772,N_38773,N_38774,N_38775,N_38776,N_38777,N_38778,N_38779,N_38780,N_38781,N_38782,N_38783,N_38784,N_38785,N_38786,N_38787,N_38788,N_38789,N_38790,N_38791,N_38792,N_38793,N_38794,N_38795,N_38796,N_38797,N_38798,N_38799,N_38800,N_38801,N_38802,N_38803,N_38804,N_38805,N_38806,N_38807,N_38808,N_38809,N_38810,N_38811,N_38812,N_38813,N_38814,N_38815,N_38816,N_38817,N_38818,N_38819,N_38820,N_38821,N_38822,N_38823,N_38824,N_38825,N_38826,N_38827,N_38828,N_38829,N_38830,N_38831,N_38832,N_38833,N_38834,N_38835,N_38836,N_38837,N_38838,N_38839,N_38840,N_38841,N_38842,N_38843,N_38844,N_38845,N_38846,N_38847,N_38848,N_38849,N_38850,N_38851,N_38852,N_38853,N_38854,N_38855,N_38856,N_38857,N_38858,N_38859,N_38860,N_38861,N_38862,N_38863,N_38864,N_38865,N_38866,N_38867,N_38868,N_38869,N_38870,N_38871,N_38872,N_38873,N_38874,N_38875,N_38876,N_38877,N_38878,N_38879,N_38880,N_38881,N_38882,N_38883,N_38884,N_38885,N_38886,N_38887,N_38888,N_38889,N_38890,N_38891,N_38892,N_38893,N_38894,N_38895,N_38896,N_38897,N_38898,N_38899,N_38900,N_38901,N_38902,N_38903,N_38904,N_38905,N_38906,N_38907,N_38908,N_38909,N_38910,N_38911,N_38912,N_38913,N_38914,N_38915,N_38916,N_38917,N_38918,N_38919,N_38920,N_38921,N_38922,N_38923,N_38924,N_38925,N_38926,N_38927,N_38928,N_38929,N_38930,N_38931,N_38932,N_38933,N_38934,N_38935,N_38936,N_38937,N_38938,N_38939,N_38940,N_38941,N_38942,N_38943,N_38944,N_38945,N_38946,N_38947,N_38948,N_38949,N_38950,N_38951,N_38952,N_38953,N_38954,N_38955,N_38956,N_38957,N_38958,N_38959,N_38960,N_38961,N_38962,N_38963,N_38964,N_38965,N_38966,N_38967,N_38968,N_38969,N_38970,N_38971,N_38972,N_38973,N_38974,N_38975,N_38976,N_38977,N_38978,N_38979,N_38980,N_38981,N_38982,N_38983,N_38984,N_38985,N_38986,N_38987,N_38988,N_38989,N_38990,N_38991,N_38992,N_38993,N_38994,N_38995,N_38996,N_38997,N_38998,N_38999,N_39000,N_39001,N_39002,N_39003,N_39004,N_39005,N_39006,N_39007,N_39008,N_39009,N_39010,N_39011,N_39012,N_39013,N_39014,N_39015,N_39016,N_39017,N_39018,N_39019,N_39020,N_39021,N_39022,N_39023,N_39024,N_39025,N_39026,N_39027,N_39028,N_39029,N_39030,N_39031,N_39032,N_39033,N_39034,N_39035,N_39036,N_39037,N_39038,N_39039,N_39040,N_39041,N_39042,N_39043,N_39044,N_39045,N_39046,N_39047,N_39048,N_39049,N_39050,N_39051,N_39052,N_39053,N_39054,N_39055,N_39056,N_39057,N_39058,N_39059,N_39060,N_39061,N_39062,N_39063,N_39064,N_39065,N_39066,N_39067,N_39068,N_39069,N_39070,N_39071,N_39072,N_39073,N_39074,N_39075,N_39076,N_39077,N_39078,N_39079,N_39080,N_39081,N_39082,N_39083,N_39084,N_39085,N_39086,N_39087,N_39088,N_39089,N_39090,N_39091,N_39092,N_39093,N_39094,N_39095,N_39096,N_39097,N_39098,N_39099,N_39100,N_39101,N_39102,N_39103,N_39104,N_39105,N_39106,N_39107,N_39108,N_39109,N_39110,N_39111,N_39112,N_39113,N_39114,N_39115,N_39116,N_39117,N_39118,N_39119,N_39120,N_39121,N_39122,N_39123,N_39124,N_39125,N_39126,N_39127,N_39128,N_39129,N_39130,N_39131,N_39132,N_39133,N_39134,N_39135,N_39136,N_39137,N_39138,N_39139,N_39140,N_39141,N_39142,N_39143,N_39144,N_39145,N_39146,N_39147,N_39148,N_39149,N_39150,N_39151,N_39152,N_39153,N_39154,N_39155,N_39156,N_39157,N_39158,N_39159,N_39160,N_39161,N_39162,N_39163,N_39164,N_39165,N_39166,N_39167,N_39168,N_39169,N_39170,N_39171,N_39172,N_39173,N_39174,N_39175,N_39176,N_39177,N_39178,N_39179,N_39180,N_39181,N_39182,N_39183,N_39184,N_39185,N_39186,N_39187,N_39188,N_39189,N_39190,N_39191,N_39192,N_39193,N_39194,N_39195,N_39196,N_39197,N_39198,N_39199,N_39200,N_39201,N_39202,N_39203,N_39204,N_39205,N_39206,N_39207,N_39208,N_39209,N_39210,N_39211,N_39212,N_39213,N_39214,N_39215,N_39216,N_39217,N_39218,N_39219,N_39220,N_39221,N_39222,N_39223,N_39224,N_39225,N_39226,N_39227,N_39228,N_39229,N_39230,N_39231,N_39232,N_39233,N_39234,N_39235,N_39236,N_39237,N_39238,N_39239,N_39240,N_39241,N_39242,N_39243,N_39244,N_39245,N_39246,N_39247,N_39248,N_39249,N_39250,N_39251,N_39252,N_39253,N_39254,N_39255,N_39256,N_39257,N_39258,N_39259,N_39260,N_39261,N_39262,N_39263,N_39264,N_39265,N_39266,N_39267,N_39268,N_39269,N_39270,N_39271,N_39272,N_39273,N_39274,N_39275,N_39276,N_39277,N_39278,N_39279,N_39280,N_39281,N_39282,N_39283,N_39284,N_39285,N_39286,N_39287,N_39288,N_39289,N_39290,N_39291,N_39292,N_39293,N_39294,N_39295,N_39296,N_39297,N_39298,N_39299,N_39300,N_39301,N_39302,N_39303,N_39304,N_39305,N_39306,N_39307,N_39308,N_39309,N_39310,N_39311,N_39312,N_39313,N_39314,N_39315,N_39316,N_39317,N_39318,N_39319,N_39320,N_39321,N_39322,N_39323,N_39324,N_39325,N_39326,N_39327,N_39328,N_39329,N_39330,N_39331,N_39332,N_39333,N_39334,N_39335,N_39336,N_39337,N_39338,N_39339,N_39340,N_39341,N_39342,N_39343,N_39344,N_39345,N_39346,N_39347,N_39348,N_39349,N_39350,N_39351,N_39352,N_39353,N_39354,N_39355,N_39356,N_39357,N_39358,N_39359,N_39360,N_39361,N_39362,N_39363,N_39364,N_39365,N_39366,N_39367,N_39368,N_39369,N_39370,N_39371,N_39372,N_39373,N_39374,N_39375,N_39376,N_39377,N_39378,N_39379,N_39380,N_39381,N_39382,N_39383,N_39384,N_39385,N_39386,N_39387,N_39388,N_39389,N_39390,N_39391,N_39392,N_39393,N_39394,N_39395,N_39396,N_39397,N_39398,N_39399,N_39400,N_39401,N_39402,N_39403,N_39404,N_39405,N_39406,N_39407,N_39408,N_39409,N_39410,N_39411,N_39412,N_39413,N_39414,N_39415,N_39416,N_39417,N_39418,N_39419,N_39420,N_39421,N_39422,N_39423,N_39424,N_39425,N_39426,N_39427,N_39428,N_39429,N_39430,N_39431,N_39432,N_39433,N_39434,N_39435,N_39436,N_39437,N_39438,N_39439,N_39440,N_39441,N_39442,N_39443,N_39444,N_39445,N_39446,N_39447,N_39448,N_39449,N_39450,N_39451,N_39452,N_39453,N_39454,N_39455,N_39456,N_39457,N_39458,N_39459,N_39460,N_39461,N_39462,N_39463,N_39464,N_39465,N_39466,N_39467,N_39468,N_39469,N_39470,N_39471,N_39472,N_39473,N_39474,N_39475,N_39476,N_39477,N_39478,N_39479,N_39480,N_39481,N_39482,N_39483,N_39484,N_39485,N_39486,N_39487,N_39488,N_39489,N_39490,N_39491,N_39492,N_39493,N_39494,N_39495,N_39496,N_39497,N_39498,N_39499,N_39500,N_39501,N_39502,N_39503,N_39504,N_39505,N_39506,N_39507,N_39508,N_39509,N_39510,N_39511,N_39512,N_39513,N_39514,N_39515,N_39516,N_39517,N_39518,N_39519,N_39520,N_39521,N_39522,N_39523,N_39524,N_39525,N_39526,N_39527,N_39528,N_39529,N_39530,N_39531,N_39532,N_39533,N_39534,N_39535,N_39536,N_39537,N_39538,N_39539,N_39540,N_39541,N_39542,N_39543,N_39544,N_39545,N_39546,N_39547,N_39548,N_39549,N_39550,N_39551,N_39552,N_39553,N_39554,N_39555,N_39556,N_39557,N_39558,N_39559,N_39560,N_39561,N_39562,N_39563,N_39564,N_39565,N_39566,N_39567,N_39568,N_39569,N_39570,N_39571,N_39572,N_39573,N_39574,N_39575,N_39576,N_39577,N_39578,N_39579,N_39580,N_39581,N_39582,N_39583,N_39584,N_39585,N_39586,N_39587,N_39588,N_39589,N_39590,N_39591,N_39592,N_39593,N_39594,N_39595,N_39596,N_39597,N_39598,N_39599,N_39600,N_39601,N_39602,N_39603,N_39604,N_39605,N_39606,N_39607,N_39608,N_39609,N_39610,N_39611,N_39612,N_39613,N_39614,N_39615,N_39616,N_39617,N_39618,N_39619,N_39620,N_39621,N_39622,N_39623,N_39624,N_39625,N_39626,N_39627,N_39628,N_39629,N_39630,N_39631,N_39632,N_39633,N_39634,N_39635,N_39636,N_39637,N_39638,N_39639,N_39640,N_39641,N_39642,N_39643,N_39644,N_39645,N_39646,N_39647,N_39648,N_39649,N_39650,N_39651,N_39652,N_39653,N_39654,N_39655,N_39656,N_39657,N_39658,N_39659,N_39660,N_39661,N_39662,N_39663,N_39664,N_39665,N_39666,N_39667,N_39668,N_39669,N_39670,N_39671,N_39672,N_39673,N_39674,N_39675,N_39676,N_39677,N_39678,N_39679,N_39680,N_39681,N_39682,N_39683,N_39684,N_39685,N_39686,N_39687,N_39688,N_39689,N_39690,N_39691,N_39692,N_39693,N_39694,N_39695,N_39696,N_39697,N_39698,N_39699,N_39700,N_39701,N_39702,N_39703,N_39704,N_39705,N_39706,N_39707,N_39708,N_39709,N_39710,N_39711,N_39712,N_39713,N_39714,N_39715,N_39716,N_39717,N_39718,N_39719,N_39720,N_39721,N_39722,N_39723,N_39724,N_39725,N_39726,N_39727,N_39728,N_39729,N_39730,N_39731,N_39732,N_39733,N_39734,N_39735,N_39736,N_39737,N_39738,N_39739,N_39740,N_39741,N_39742,N_39743,N_39744,N_39745,N_39746,N_39747,N_39748,N_39749,N_39750,N_39751,N_39752,N_39753,N_39754,N_39755,N_39756,N_39757,N_39758,N_39759,N_39760,N_39761,N_39762,N_39763,N_39764,N_39765,N_39766,N_39767,N_39768,N_39769,N_39770,N_39771,N_39772,N_39773,N_39774,N_39775,N_39776,N_39777,N_39778,N_39779,N_39780,N_39781,N_39782,N_39783,N_39784,N_39785,N_39786,N_39787,N_39788,N_39789,N_39790,N_39791,N_39792,N_39793,N_39794,N_39795,N_39796,N_39797,N_39798,N_39799,N_39800,N_39801,N_39802,N_39803,N_39804,N_39805,N_39806,N_39807,N_39808,N_39809,N_39810,N_39811,N_39812,N_39813,N_39814,N_39815,N_39816,N_39817,N_39818,N_39819,N_39820,N_39821,N_39822,N_39823,N_39824,N_39825,N_39826,N_39827,N_39828,N_39829,N_39830,N_39831,N_39832,N_39833,N_39834,N_39835,N_39836,N_39837,N_39838,N_39839,N_39840,N_39841,N_39842,N_39843,N_39844,N_39845,N_39846,N_39847,N_39848,N_39849,N_39850,N_39851,N_39852,N_39853,N_39854,N_39855,N_39856,N_39857,N_39858,N_39859,N_39860,N_39861,N_39862,N_39863,N_39864,N_39865,N_39866,N_39867,N_39868,N_39869,N_39870,N_39871,N_39872,N_39873,N_39874,N_39875,N_39876,N_39877,N_39878,N_39879,N_39880,N_39881,N_39882,N_39883,N_39884,N_39885,N_39886,N_39887,N_39888,N_39889,N_39890,N_39891,N_39892,N_39893,N_39894,N_39895,N_39896,N_39897,N_39898,N_39899,N_39900,N_39901,N_39902,N_39903,N_39904,N_39905,N_39906,N_39907,N_39908,N_39909,N_39910,N_39911,N_39912,N_39913,N_39914,N_39915,N_39916,N_39917,N_39918,N_39919,N_39920,N_39921,N_39922,N_39923,N_39924,N_39925,N_39926,N_39927,N_39928,N_39929,N_39930,N_39931,N_39932,N_39933,N_39934,N_39935,N_39936,N_39937,N_39938,N_39939,N_39940,N_39941,N_39942,N_39943,N_39944,N_39945,N_39946,N_39947,N_39948,N_39949,N_39950,N_39951,N_39952,N_39953,N_39954,N_39955,N_39956,N_39957,N_39958,N_39959,N_39960,N_39961,N_39962,N_39963,N_39964,N_39965,N_39966,N_39967,N_39968,N_39969,N_39970,N_39971,N_39972,N_39973,N_39974,N_39975,N_39976,N_39977,N_39978,N_39979,N_39980,N_39981,N_39982,N_39983,N_39984,N_39985,N_39986,N_39987,N_39988,N_39989,N_39990,N_39991,N_39992,N_39993,N_39994,N_39995,N_39996,N_39997,N_39998,N_39999,N_40000,N_40001,N_40002,N_40003,N_40004,N_40005,N_40006,N_40007,N_40008,N_40009,N_40010,N_40011,N_40012,N_40013,N_40014,N_40015,N_40016,N_40017,N_40018,N_40019,N_40020,N_40021,N_40022,N_40023,N_40024,N_40025,N_40026,N_40027,N_40028,N_40029,N_40030,N_40031,N_40032,N_40033,N_40034,N_40035,N_40036,N_40037,N_40038,N_40039,N_40040,N_40041,N_40042,N_40043,N_40044,N_40045,N_40046,N_40047,N_40048,N_40049,N_40050,N_40051,N_40052,N_40053,N_40054,N_40055,N_40056,N_40057,N_40058,N_40059,N_40060,N_40061,N_40062,N_40063,N_40064,N_40065,N_40066,N_40067,N_40068,N_40069,N_40070,N_40071,N_40072,N_40073,N_40074,N_40075,N_40076,N_40077,N_40078,N_40079,N_40080,N_40081,N_40082,N_40083,N_40084,N_40085,N_40086,N_40087,N_40088,N_40089,N_40090,N_40091,N_40092,N_40093,N_40094,N_40095,N_40096,N_40097,N_40098,N_40099,N_40100,N_40101,N_40102,N_40103,N_40104,N_40105,N_40106,N_40107,N_40108,N_40109,N_40110,N_40111,N_40112,N_40113,N_40114,N_40115,N_40116,N_40117,N_40118,N_40119,N_40120,N_40121,N_40122,N_40123,N_40124,N_40125,N_40126,N_40127,N_40128,N_40129,N_40130,N_40131,N_40132,N_40133,N_40134,N_40135,N_40136,N_40137,N_40138,N_40139,N_40140,N_40141,N_40142,N_40143,N_40144,N_40145,N_40146,N_40147,N_40148,N_40149,N_40150,N_40151,N_40152,N_40153,N_40154,N_40155,N_40156,N_40157,N_40158,N_40159,N_40160,N_40161,N_40162,N_40163,N_40164,N_40165,N_40166,N_40167,N_40168,N_40169,N_40170,N_40171,N_40172,N_40173,N_40174,N_40175,N_40176,N_40177,N_40178,N_40179,N_40180,N_40181,N_40182,N_40183,N_40184,N_40185,N_40186,N_40187,N_40188,N_40189,N_40190,N_40191,N_40192,N_40193,N_40194,N_40195,N_40196,N_40197,N_40198,N_40199,N_40200,N_40201,N_40202,N_40203,N_40204,N_40205,N_40206,N_40207,N_40208,N_40209,N_40210,N_40211,N_40212,N_40213,N_40214,N_40215,N_40216,N_40217,N_40218,N_40219,N_40220,N_40221,N_40222,N_40223,N_40224,N_40225,N_40226,N_40227,N_40228,N_40229,N_40230,N_40231,N_40232,N_40233,N_40234,N_40235,N_40236,N_40237,N_40238,N_40239,N_40240,N_40241,N_40242,N_40243,N_40244,N_40245,N_40246,N_40247,N_40248,N_40249,N_40250,N_40251,N_40252,N_40253,N_40254,N_40255,N_40256,N_40257,N_40258,N_40259,N_40260,N_40261,N_40262,N_40263,N_40264,N_40265,N_40266,N_40267,N_40268,N_40269,N_40270,N_40271,N_40272,N_40273,N_40274,N_40275,N_40276,N_40277,N_40278,N_40279,N_40280,N_40281,N_40282,N_40283,N_40284,N_40285,N_40286,N_40287,N_40288,N_40289,N_40290,N_40291,N_40292,N_40293,N_40294,N_40295,N_40296,N_40297,N_40298,N_40299,N_40300,N_40301,N_40302,N_40303,N_40304,N_40305,N_40306,N_40307,N_40308,N_40309,N_40310,N_40311,N_40312,N_40313,N_40314,N_40315,N_40316,N_40317,N_40318,N_40319,N_40320,N_40321,N_40322,N_40323,N_40324,N_40325,N_40326,N_40327,N_40328,N_40329,N_40330,N_40331,N_40332,N_40333,N_40334,N_40335,N_40336,N_40337,N_40338,N_40339,N_40340,N_40341,N_40342,N_40343,N_40344,N_40345,N_40346,N_40347,N_40348,N_40349,N_40350,N_40351,N_40352,N_40353,N_40354,N_40355,N_40356,N_40357,N_40358,N_40359,N_40360,N_40361,N_40362,N_40363,N_40364,N_40365,N_40366,N_40367,N_40368,N_40369,N_40370,N_40371,N_40372,N_40373,N_40374,N_40375,N_40376,N_40377,N_40378,N_40379,N_40380,N_40381,N_40382,N_40383,N_40384,N_40385,N_40386,N_40387,N_40388,N_40389,N_40390,N_40391,N_40392,N_40393,N_40394,N_40395,N_40396,N_40397,N_40398,N_40399,N_40400,N_40401,N_40402,N_40403,N_40404,N_40405,N_40406,N_40407,N_40408,N_40409,N_40410,N_40411,N_40412,N_40413,N_40414,N_40415,N_40416,N_40417,N_40418,N_40419,N_40420,N_40421,N_40422,N_40423,N_40424,N_40425,N_40426,N_40427,N_40428,N_40429,N_40430,N_40431,N_40432,N_40433,N_40434,N_40435,N_40436,N_40437,N_40438,N_40439,N_40440,N_40441,N_40442,N_40443,N_40444,N_40445,N_40446,N_40447,N_40448,N_40449,N_40450,N_40451,N_40452,N_40453,N_40454,N_40455,N_40456,N_40457,N_40458,N_40459,N_40460,N_40461,N_40462,N_40463,N_40464,N_40465,N_40466,N_40467,N_40468,N_40469,N_40470,N_40471,N_40472,N_40473,N_40474,N_40475,N_40476,N_40477,N_40478,N_40479,N_40480,N_40481,N_40482,N_40483,N_40484,N_40485,N_40486,N_40487,N_40488,N_40489,N_40490,N_40491,N_40492,N_40493,N_40494,N_40495,N_40496,N_40497,N_40498,N_40499,N_40500,N_40501,N_40502,N_40503,N_40504,N_40505,N_40506,N_40507,N_40508,N_40509,N_40510,N_40511,N_40512,N_40513,N_40514,N_40515,N_40516,N_40517,N_40518,N_40519,N_40520,N_40521,N_40522,N_40523,N_40524,N_40525,N_40526,N_40527,N_40528,N_40529,N_40530,N_40531,N_40532,N_40533,N_40534,N_40535,N_40536,N_40537,N_40538,N_40539,N_40540,N_40541,N_40542,N_40543,N_40544,N_40545,N_40546,N_40547,N_40548,N_40549,N_40550,N_40551,N_40552,N_40553,N_40554,N_40555,N_40556,N_40557,N_40558,N_40559,N_40560,N_40561,N_40562,N_40563,N_40564,N_40565,N_40566,N_40567,N_40568,N_40569,N_40570,N_40571,N_40572,N_40573,N_40574,N_40575,N_40576,N_40577,N_40578,N_40579,N_40580,N_40581,N_40582,N_40583,N_40584,N_40585,N_40586,N_40587,N_40588,N_40589,N_40590,N_40591,N_40592,N_40593,N_40594,N_40595,N_40596,N_40597,N_40598,N_40599,N_40600,N_40601,N_40602,N_40603,N_40604,N_40605,N_40606,N_40607,N_40608,N_40609,N_40610,N_40611,N_40612,N_40613,N_40614,N_40615,N_40616,N_40617,N_40618,N_40619,N_40620,N_40621,N_40622,N_40623,N_40624,N_40625,N_40626,N_40627,N_40628,N_40629,N_40630,N_40631,N_40632,N_40633,N_40634,N_40635,N_40636,N_40637,N_40638,N_40639,N_40640,N_40641,N_40642,N_40643,N_40644,N_40645,N_40646,N_40647,N_40648,N_40649,N_40650,N_40651,N_40652,N_40653,N_40654,N_40655,N_40656,N_40657,N_40658,N_40659,N_40660,N_40661,N_40662,N_40663,N_40664,N_40665,N_40666,N_40667,N_40668,N_40669,N_40670,N_40671,N_40672,N_40673,N_40674,N_40675,N_40676,N_40677,N_40678,N_40679,N_40680,N_40681,N_40682,N_40683,N_40684,N_40685,N_40686,N_40687,N_40688,N_40689,N_40690,N_40691,N_40692,N_40693,N_40694,N_40695,N_40696,N_40697,N_40698,N_40699,N_40700,N_40701,N_40702,N_40703,N_40704,N_40705,N_40706,N_40707,N_40708,N_40709,N_40710,N_40711,N_40712,N_40713,N_40714,N_40715,N_40716,N_40717,N_40718,N_40719,N_40720,N_40721,N_40722,N_40723,N_40724,N_40725,N_40726,N_40727,N_40728,N_40729,N_40730,N_40731,N_40732,N_40733,N_40734,N_40735,N_40736,N_40737,N_40738,N_40739,N_40740,N_40741,N_40742,N_40743,N_40744,N_40745,N_40746,N_40747,N_40748,N_40749,N_40750,N_40751,N_40752,N_40753,N_40754,N_40755,N_40756,N_40757,N_40758,N_40759,N_40760,N_40761,N_40762,N_40763,N_40764,N_40765,N_40766,N_40767,N_40768,N_40769,N_40770,N_40771,N_40772,N_40773,N_40774,N_40775,N_40776,N_40777,N_40778,N_40779,N_40780,N_40781,N_40782,N_40783,N_40784,N_40785,N_40786,N_40787,N_40788,N_40789,N_40790,N_40791,N_40792,N_40793,N_40794,N_40795,N_40796,N_40797,N_40798,N_40799,N_40800,N_40801,N_40802,N_40803,N_40804,N_40805,N_40806,N_40807,N_40808,N_40809,N_40810,N_40811,N_40812,N_40813,N_40814,N_40815,N_40816,N_40817,N_40818,N_40819,N_40820,N_40821,N_40822,N_40823,N_40824,N_40825,N_40826,N_40827,N_40828,N_40829,N_40830,N_40831,N_40832,N_40833,N_40834,N_40835,N_40836,N_40837,N_40838,N_40839,N_40840,N_40841,N_40842,N_40843,N_40844,N_40845,N_40846,N_40847,N_40848,N_40849,N_40850,N_40851,N_40852,N_40853,N_40854,N_40855,N_40856,N_40857,N_40858,N_40859,N_40860,N_40861,N_40862,N_40863,N_40864,N_40865,N_40866,N_40867,N_40868,N_40869,N_40870,N_40871,N_40872,N_40873,N_40874,N_40875,N_40876,N_40877,N_40878,N_40879,N_40880,N_40881,N_40882,N_40883,N_40884,N_40885,N_40886,N_40887,N_40888,N_40889,N_40890,N_40891,N_40892,N_40893,N_40894,N_40895,N_40896,N_40897,N_40898,N_40899,N_40900,N_40901,N_40902,N_40903,N_40904,N_40905,N_40906,N_40907,N_40908,N_40909,N_40910,N_40911,N_40912,N_40913,N_40914,N_40915,N_40916,N_40917,N_40918,N_40919,N_40920,N_40921,N_40922,N_40923,N_40924,N_40925,N_40926,N_40927,N_40928,N_40929,N_40930,N_40931,N_40932,N_40933,N_40934,N_40935,N_40936,N_40937,N_40938,N_40939,N_40940,N_40941,N_40942,N_40943,N_40944,N_40945,N_40946,N_40947,N_40948,N_40949,N_40950,N_40951,N_40952,N_40953,N_40954,N_40955,N_40956,N_40957,N_40958,N_40959,N_40960,N_40961,N_40962,N_40963,N_40964,N_40965,N_40966,N_40967,N_40968,N_40969,N_40970,N_40971,N_40972,N_40973,N_40974,N_40975,N_40976,N_40977,N_40978,N_40979,N_40980,N_40981,N_40982,N_40983,N_40984,N_40985,N_40986,N_40987,N_40988,N_40989,N_40990,N_40991,N_40992,N_40993,N_40994,N_40995,N_40996,N_40997,N_40998,N_40999,N_41000,N_41001,N_41002,N_41003,N_41004,N_41005,N_41006,N_41007,N_41008,N_41009,N_41010,N_41011,N_41012,N_41013,N_41014,N_41015,N_41016,N_41017,N_41018,N_41019,N_41020,N_41021,N_41022,N_41023,N_41024,N_41025,N_41026,N_41027,N_41028,N_41029,N_41030,N_41031,N_41032,N_41033,N_41034,N_41035,N_41036,N_41037,N_41038,N_41039,N_41040,N_41041,N_41042,N_41043,N_41044,N_41045,N_41046,N_41047,N_41048,N_41049,N_41050,N_41051,N_41052,N_41053,N_41054,N_41055,N_41056,N_41057,N_41058,N_41059,N_41060,N_41061,N_41062,N_41063,N_41064,N_41065,N_41066,N_41067,N_41068,N_41069,N_41070,N_41071,N_41072,N_41073,N_41074,N_41075,N_41076,N_41077,N_41078,N_41079,N_41080,N_41081,N_41082,N_41083,N_41084,N_41085,N_41086,N_41087,N_41088,N_41089,N_41090,N_41091,N_41092,N_41093,N_41094,N_41095,N_41096,N_41097,N_41098,N_41099,N_41100,N_41101,N_41102,N_41103,N_41104,N_41105,N_41106,N_41107,N_41108,N_41109,N_41110,N_41111,N_41112,N_41113,N_41114,N_41115,N_41116,N_41117,N_41118,N_41119,N_41120,N_41121,N_41122,N_41123,N_41124,N_41125,N_41126,N_41127,N_41128,N_41129,N_41130,N_41131,N_41132,N_41133,N_41134,N_41135,N_41136,N_41137,N_41138,N_41139,N_41140,N_41141,N_41142,N_41143,N_41144,N_41145,N_41146,N_41147,N_41148,N_41149,N_41150,N_41151,N_41152,N_41153,N_41154,N_41155,N_41156,N_41157,N_41158,N_41159,N_41160,N_41161,N_41162,N_41163,N_41164,N_41165,N_41166,N_41167,N_41168,N_41169,N_41170,N_41171,N_41172,N_41173,N_41174,N_41175,N_41176,N_41177,N_41178,N_41179,N_41180,N_41181,N_41182,N_41183,N_41184,N_41185,N_41186,N_41187,N_41188,N_41189,N_41190,N_41191,N_41192,N_41193,N_41194,N_41195,N_41196,N_41197,N_41198,N_41199,N_41200,N_41201,N_41202,N_41203,N_41204,N_41205,N_41206,N_41207,N_41208,N_41209,N_41210,N_41211,N_41212,N_41213,N_41214,N_41215,N_41216,N_41217,N_41218,N_41219,N_41220,N_41221,N_41222,N_41223,N_41224,N_41225,N_41226,N_41227,N_41228,N_41229,N_41230,N_41231,N_41232,N_41233,N_41234,N_41235,N_41236,N_41237,N_41238,N_41239,N_41240,N_41241,N_41242,N_41243,N_41244,N_41245,N_41246,N_41247,N_41248,N_41249,N_41250,N_41251,N_41252,N_41253,N_41254,N_41255,N_41256,N_41257,N_41258,N_41259,N_41260,N_41261,N_41262,N_41263,N_41264,N_41265,N_41266,N_41267,N_41268,N_41269,N_41270,N_41271,N_41272,N_41273,N_41274,N_41275,N_41276,N_41277,N_41278,N_41279,N_41280,N_41281,N_41282,N_41283,N_41284,N_41285,N_41286,N_41287,N_41288,N_41289,N_41290,N_41291,N_41292,N_41293,N_41294,N_41295,N_41296,N_41297,N_41298,N_41299,N_41300,N_41301,N_41302,N_41303,N_41304,N_41305,N_41306,N_41307,N_41308,N_41309,N_41310,N_41311,N_41312,N_41313,N_41314,N_41315,N_41316,N_41317,N_41318,N_41319,N_41320,N_41321,N_41322,N_41323,N_41324,N_41325,N_41326,N_41327,N_41328,N_41329,N_41330,N_41331,N_41332,N_41333,N_41334,N_41335,N_41336,N_41337,N_41338,N_41339,N_41340,N_41341,N_41342,N_41343,N_41344,N_41345,N_41346,N_41347,N_41348,N_41349,N_41350,N_41351,N_41352,N_41353,N_41354,N_41355,N_41356,N_41357,N_41358,N_41359,N_41360,N_41361,N_41362,N_41363,N_41364,N_41365,N_41366,N_41367,N_41368,N_41369,N_41370,N_41371,N_41372,N_41373,N_41374,N_41375,N_41376,N_41377,N_41378,N_41379,N_41380,N_41381,N_41382,N_41383,N_41384,N_41385,N_41386,N_41387,N_41388,N_41389,N_41390,N_41391,N_41392,N_41393,N_41394,N_41395,N_41396,N_41397,N_41398,N_41399,N_41400,N_41401,N_41402,N_41403,N_41404,N_41405,N_41406,N_41407,N_41408,N_41409,N_41410,N_41411,N_41412,N_41413,N_41414,N_41415,N_41416,N_41417,N_41418,N_41419,N_41420,N_41421,N_41422,N_41423,N_41424,N_41425,N_41426,N_41427,N_41428,N_41429,N_41430,N_41431,N_41432,N_41433,N_41434,N_41435,N_41436,N_41437,N_41438,N_41439,N_41440,N_41441,N_41442,N_41443,N_41444,N_41445,N_41446,N_41447,N_41448,N_41449,N_41450,N_41451,N_41452,N_41453,N_41454,N_41455,N_41456,N_41457,N_41458,N_41459,N_41460,N_41461,N_41462,N_41463,N_41464,N_41465,N_41466,N_41467,N_41468,N_41469,N_41470,N_41471,N_41472,N_41473,N_41474,N_41475,N_41476,N_41477,N_41478,N_41479,N_41480,N_41481,N_41482,N_41483,N_41484,N_41485,N_41486,N_41487,N_41488,N_41489,N_41490,N_41491,N_41492,N_41493,N_41494,N_41495,N_41496,N_41497,N_41498,N_41499,N_41500,N_41501,N_41502,N_41503,N_41504,N_41505,N_41506,N_41507,N_41508,N_41509,N_41510,N_41511,N_41512,N_41513,N_41514,N_41515,N_41516,N_41517,N_41518,N_41519,N_41520,N_41521,N_41522,N_41523,N_41524,N_41525,N_41526,N_41527,N_41528,N_41529,N_41530,N_41531,N_41532,N_41533,N_41534,N_41535,N_41536,N_41537,N_41538,N_41539,N_41540,N_41541,N_41542,N_41543,N_41544,N_41545,N_41546,N_41547,N_41548,N_41549,N_41550,N_41551,N_41552,N_41553,N_41554,N_41555,N_41556,N_41557,N_41558,N_41559,N_41560,N_41561,N_41562,N_41563,N_41564,N_41565,N_41566,N_41567,N_41568,N_41569,N_41570,N_41571,N_41572,N_41573,N_41574,N_41575,N_41576,N_41577,N_41578,N_41579,N_41580,N_41581,N_41582,N_41583,N_41584,N_41585,N_41586,N_41587,N_41588,N_41589,N_41590,N_41591,N_41592,N_41593,N_41594,N_41595,N_41596,N_41597,N_41598,N_41599,N_41600,N_41601,N_41602,N_41603,N_41604,N_41605,N_41606,N_41607,N_41608,N_41609,N_41610,N_41611,N_41612,N_41613,N_41614,N_41615,N_41616,N_41617,N_41618,N_41619,N_41620,N_41621,N_41622,N_41623,N_41624,N_41625,N_41626,N_41627,N_41628,N_41629,N_41630,N_41631,N_41632,N_41633,N_41634,N_41635,N_41636,N_41637,N_41638,N_41639,N_41640,N_41641,N_41642,N_41643,N_41644,N_41645,N_41646,N_41647,N_41648,N_41649,N_41650,N_41651,N_41652,N_41653,N_41654,N_41655,N_41656,N_41657,N_41658,N_41659,N_41660,N_41661,N_41662,N_41663,N_41664,N_41665,N_41666,N_41667,N_41668,N_41669,N_41670,N_41671,N_41672,N_41673,N_41674,N_41675,N_41676,N_41677,N_41678,N_41679,N_41680,N_41681,N_41682,N_41683,N_41684,N_41685,N_41686,N_41687,N_41688,N_41689,N_41690,N_41691,N_41692,N_41693,N_41694,N_41695,N_41696,N_41697,N_41698,N_41699,N_41700,N_41701,N_41702,N_41703,N_41704,N_41705,N_41706,N_41707,N_41708,N_41709,N_41710,N_41711,N_41712,N_41713,N_41714,N_41715,N_41716,N_41717,N_41718,N_41719,N_41720,N_41721,N_41722,N_41723,N_41724,N_41725,N_41726,N_41727,N_41728,N_41729,N_41730,N_41731,N_41732,N_41733,N_41734,N_41735,N_41736,N_41737,N_41738,N_41739,N_41740,N_41741,N_41742,N_41743,N_41744,N_41745,N_41746,N_41747,N_41748,N_41749,N_41750,N_41751,N_41752,N_41753,N_41754,N_41755,N_41756,N_41757,N_41758,N_41759,N_41760,N_41761,N_41762,N_41763,N_41764,N_41765,N_41766,N_41767,N_41768,N_41769,N_41770,N_41771,N_41772,N_41773,N_41774,N_41775,N_41776,N_41777,N_41778,N_41779,N_41780,N_41781,N_41782,N_41783,N_41784,N_41785,N_41786,N_41787,N_41788,N_41789,N_41790,N_41791,N_41792,N_41793,N_41794,N_41795,N_41796,N_41797,N_41798,N_41799,N_41800,N_41801,N_41802,N_41803,N_41804,N_41805,N_41806,N_41807,N_41808,N_41809,N_41810,N_41811,N_41812,N_41813,N_41814,N_41815,N_41816,N_41817,N_41818,N_41819,N_41820,N_41821,N_41822,N_41823,N_41824,N_41825,N_41826,N_41827,N_41828,N_41829,N_41830,N_41831,N_41832,N_41833,N_41834,N_41835,N_41836,N_41837,N_41838,N_41839,N_41840,N_41841,N_41842,N_41843,N_41844,N_41845,N_41846,N_41847,N_41848,N_41849,N_41850,N_41851,N_41852,N_41853,N_41854,N_41855,N_41856,N_41857,N_41858,N_41859,N_41860,N_41861,N_41862,N_41863,N_41864,N_41865,N_41866,N_41867,N_41868,N_41869,N_41870,N_41871,N_41872,N_41873,N_41874,N_41875,N_41876,N_41877,N_41878,N_41879,N_41880,N_41881,N_41882,N_41883,N_41884,N_41885,N_41886,N_41887,N_41888,N_41889,N_41890,N_41891,N_41892,N_41893,N_41894,N_41895,N_41896,N_41897,N_41898,N_41899,N_41900,N_41901,N_41902,N_41903,N_41904,N_41905,N_41906,N_41907,N_41908,N_41909,N_41910,N_41911,N_41912,N_41913,N_41914,N_41915,N_41916,N_41917,N_41918,N_41919,N_41920,N_41921,N_41922,N_41923,N_41924,N_41925,N_41926,N_41927,N_41928,N_41929,N_41930,N_41931,N_41932,N_41933,N_41934,N_41935,N_41936,N_41937,N_41938,N_41939,N_41940,N_41941,N_41942,N_41943,N_41944,N_41945,N_41946,N_41947,N_41948,N_41949,N_41950,N_41951,N_41952,N_41953,N_41954,N_41955,N_41956,N_41957,N_41958,N_41959,N_41960,N_41961,N_41962,N_41963,N_41964,N_41965,N_41966,N_41967,N_41968,N_41969,N_41970,N_41971,N_41972,N_41973,N_41974,N_41975,N_41976,N_41977,N_41978,N_41979,N_41980,N_41981,N_41982,N_41983,N_41984,N_41985,N_41986,N_41987,N_41988,N_41989,N_41990,N_41991,N_41992,N_41993,N_41994,N_41995,N_41996,N_41997,N_41998,N_41999,N_42000,N_42001,N_42002,N_42003,N_42004,N_42005,N_42006,N_42007,N_42008,N_42009,N_42010,N_42011,N_42012,N_42013,N_42014,N_42015,N_42016,N_42017,N_42018,N_42019,N_42020,N_42021,N_42022,N_42023,N_42024,N_42025,N_42026,N_42027,N_42028,N_42029,N_42030,N_42031,N_42032,N_42033,N_42034,N_42035,N_42036,N_42037,N_42038,N_42039,N_42040,N_42041,N_42042,N_42043,N_42044,N_42045,N_42046,N_42047,N_42048,N_42049,N_42050,N_42051,N_42052,N_42053,N_42054,N_42055,N_42056,N_42057,N_42058,N_42059,N_42060,N_42061,N_42062,N_42063,N_42064,N_42065,N_42066,N_42067,N_42068,N_42069,N_42070,N_42071,N_42072,N_42073,N_42074,N_42075,N_42076,N_42077,N_42078,N_42079,N_42080,N_42081,N_42082,N_42083,N_42084,N_42085,N_42086,N_42087,N_42088,N_42089,N_42090,N_42091,N_42092,N_42093,N_42094,N_42095,N_42096,N_42097,N_42098,N_42099,N_42100,N_42101,N_42102,N_42103,N_42104,N_42105,N_42106,N_42107,N_42108,N_42109,N_42110,N_42111,N_42112,N_42113,N_42114,N_42115,N_42116,N_42117,N_42118,N_42119,N_42120,N_42121,N_42122,N_42123,N_42124,N_42125,N_42126,N_42127,N_42128,N_42129,N_42130,N_42131,N_42132,N_42133,N_42134,N_42135,N_42136,N_42137,N_42138,N_42139,N_42140,N_42141,N_42142,N_42143,N_42144,N_42145,N_42146,N_42147,N_42148,N_42149,N_42150,N_42151,N_42152,N_42153,N_42154,N_42155,N_42156,N_42157,N_42158,N_42159,N_42160,N_42161,N_42162,N_42163,N_42164,N_42165,N_42166,N_42167,N_42168,N_42169,N_42170,N_42171,N_42172,N_42173,N_42174,N_42175,N_42176,N_42177,N_42178,N_42179,N_42180,N_42181,N_42182,N_42183,N_42184,N_42185,N_42186,N_42187,N_42188,N_42189,N_42190,N_42191,N_42192,N_42193,N_42194,N_42195,N_42196,N_42197,N_42198,N_42199,N_42200,N_42201,N_42202,N_42203,N_42204,N_42205,N_42206,N_42207,N_42208,N_42209,N_42210,N_42211,N_42212,N_42213,N_42214,N_42215,N_42216,N_42217,N_42218,N_42219,N_42220,N_42221,N_42222,N_42223,N_42224,N_42225,N_42226,N_42227,N_42228,N_42229,N_42230,N_42231,N_42232,N_42233,N_42234,N_42235,N_42236,N_42237,N_42238,N_42239,N_42240,N_42241,N_42242,N_42243,N_42244,N_42245,N_42246,N_42247,N_42248,N_42249,N_42250,N_42251,N_42252,N_42253,N_42254,N_42255,N_42256,N_42257,N_42258,N_42259,N_42260,N_42261,N_42262,N_42263,N_42264,N_42265,N_42266,N_42267,N_42268,N_42269,N_42270,N_42271,N_42272,N_42273,N_42274,N_42275,N_42276,N_42277,N_42278,N_42279,N_42280,N_42281,N_42282,N_42283,N_42284,N_42285,N_42286,N_42287,N_42288,N_42289,N_42290,N_42291,N_42292,N_42293,N_42294,N_42295,N_42296,N_42297,N_42298,N_42299,N_42300,N_42301,N_42302,N_42303,N_42304,N_42305,N_42306,N_42307,N_42308,N_42309,N_42310,N_42311,N_42312,N_42313,N_42314,N_42315,N_42316,N_42317,N_42318,N_42319,N_42320,N_42321,N_42322,N_42323,N_42324,N_42325,N_42326,N_42327,N_42328,N_42329,N_42330,N_42331,N_42332,N_42333,N_42334,N_42335,N_42336,N_42337,N_42338,N_42339,N_42340,N_42341,N_42342,N_42343,N_42344,N_42345,N_42346,N_42347,N_42348,N_42349,N_42350,N_42351,N_42352,N_42353,N_42354,N_42355,N_42356,N_42357,N_42358,N_42359,N_42360,N_42361,N_42362,N_42363,N_42364,N_42365,N_42366,N_42367,N_42368,N_42369,N_42370,N_42371,N_42372,N_42373,N_42374,N_42375,N_42376,N_42377,N_42378,N_42379,N_42380,N_42381,N_42382,N_42383,N_42384,N_42385,N_42386,N_42387,N_42388,N_42389,N_42390,N_42391,N_42392,N_42393,N_42394,N_42395,N_42396,N_42397,N_42398,N_42399,N_42400,N_42401,N_42402,N_42403,N_42404,N_42405,N_42406,N_42407,N_42408,N_42409,N_42410,N_42411,N_42412,N_42413,N_42414,N_42415,N_42416,N_42417,N_42418,N_42419,N_42420,N_42421,N_42422,N_42423,N_42424,N_42425,N_42426,N_42427,N_42428,N_42429,N_42430,N_42431,N_42432,N_42433,N_42434,N_42435,N_42436,N_42437,N_42438,N_42439,N_42440,N_42441,N_42442,N_42443,N_42444,N_42445,N_42446,N_42447,N_42448,N_42449,N_42450,N_42451,N_42452,N_42453,N_42454,N_42455,N_42456,N_42457,N_42458,N_42459,N_42460,N_42461,N_42462,N_42463,N_42464,N_42465,N_42466,N_42467,N_42468,N_42469,N_42470,N_42471,N_42472,N_42473,N_42474,N_42475,N_42476,N_42477,N_42478,N_42479,N_42480,N_42481,N_42482,N_42483,N_42484,N_42485,N_42486,N_42487,N_42488,N_42489,N_42490,N_42491,N_42492,N_42493,N_42494,N_42495,N_42496,N_42497,N_42498,N_42499,N_42500,N_42501,N_42502,N_42503,N_42504,N_42505,N_42506,N_42507,N_42508,N_42509,N_42510,N_42511,N_42512,N_42513,N_42514,N_42515,N_42516,N_42517,N_42518,N_42519,N_42520,N_42521,N_42522,N_42523,N_42524,N_42525,N_42526,N_42527,N_42528,N_42529,N_42530,N_42531,N_42532,N_42533,N_42534,N_42535,N_42536,N_42537,N_42538,N_42539,N_42540,N_42541,N_42542,N_42543,N_42544,N_42545,N_42546,N_42547,N_42548,N_42549,N_42550,N_42551,N_42552,N_42553,N_42554,N_42555,N_42556,N_42557,N_42558,N_42559,N_42560,N_42561,N_42562,N_42563,N_42564,N_42565,N_42566,N_42567,N_42568,N_42569,N_42570,N_42571,N_42572,N_42573,N_42574,N_42575,N_42576,N_42577,N_42578,N_42579,N_42580,N_42581,N_42582,N_42583,N_42584,N_42585,N_42586,N_42587,N_42588,N_42589,N_42590,N_42591,N_42592,N_42593,N_42594,N_42595,N_42596,N_42597,N_42598,N_42599,N_42600,N_42601,N_42602,N_42603,N_42604,N_42605,N_42606,N_42607,N_42608,N_42609,N_42610,N_42611,N_42612,N_42613,N_42614,N_42615,N_42616,N_42617,N_42618,N_42619,N_42620,N_42621,N_42622,N_42623,N_42624,N_42625,N_42626,N_42627,N_42628,N_42629,N_42630,N_42631,N_42632,N_42633,N_42634,N_42635,N_42636,N_42637,N_42638,N_42639,N_42640,N_42641,N_42642,N_42643,N_42644,N_42645,N_42646,N_42647,N_42648,N_42649,N_42650,N_42651,N_42652,N_42653,N_42654,N_42655,N_42656,N_42657,N_42658,N_42659,N_42660,N_42661,N_42662,N_42663,N_42664,N_42665,N_42666,N_42667,N_42668,N_42669,N_42670,N_42671,N_42672,N_42673,N_42674,N_42675,N_42676,N_42677,N_42678,N_42679,N_42680,N_42681,N_42682,N_42683,N_42684,N_42685,N_42686,N_42687,N_42688,N_42689,N_42690,N_42691,N_42692,N_42693,N_42694,N_42695,N_42696,N_42697,N_42698,N_42699,N_42700,N_42701,N_42702,N_42703,N_42704,N_42705,N_42706,N_42707,N_42708,N_42709,N_42710,N_42711,N_42712,N_42713,N_42714,N_42715,N_42716,N_42717,N_42718,N_42719,N_42720,N_42721,N_42722,N_42723,N_42724,N_42725,N_42726,N_42727,N_42728,N_42729,N_42730,N_42731,N_42732,N_42733,N_42734,N_42735,N_42736,N_42737,N_42738,N_42739,N_42740,N_42741,N_42742,N_42743,N_42744,N_42745,N_42746,N_42747,N_42748,N_42749,N_42750,N_42751,N_42752,N_42753,N_42754,N_42755,N_42756,N_42757,N_42758,N_42759,N_42760,N_42761,N_42762,N_42763,N_42764,N_42765,N_42766,N_42767,N_42768,N_42769,N_42770,N_42771,N_42772,N_42773,N_42774,N_42775,N_42776,N_42777,N_42778,N_42779,N_42780,N_42781,N_42782,N_42783,N_42784,N_42785,N_42786,N_42787,N_42788,N_42789,N_42790,N_42791,N_42792,N_42793,N_42794,N_42795,N_42796,N_42797,N_42798,N_42799,N_42800,N_42801,N_42802,N_42803,N_42804,N_42805,N_42806,N_42807,N_42808,N_42809,N_42810,N_42811,N_42812,N_42813,N_42814,N_42815,N_42816,N_42817,N_42818,N_42819,N_42820,N_42821,N_42822,N_42823,N_42824,N_42825,N_42826,N_42827,N_42828,N_42829,N_42830,N_42831,N_42832,N_42833,N_42834,N_42835,N_42836,N_42837,N_42838,N_42839,N_42840,N_42841,N_42842,N_42843,N_42844,N_42845,N_42846,N_42847,N_42848,N_42849,N_42850,N_42851,N_42852,N_42853,N_42854,N_42855,N_42856,N_42857,N_42858,N_42859,N_42860,N_42861,N_42862,N_42863,N_42864,N_42865,N_42866,N_42867,N_42868,N_42869,N_42870,N_42871,N_42872,N_42873,N_42874,N_42875,N_42876,N_42877,N_42878,N_42879,N_42880,N_42881,N_42882,N_42883,N_42884,N_42885,N_42886,N_42887,N_42888,N_42889,N_42890,N_42891,N_42892,N_42893,N_42894,N_42895,N_42896,N_42897,N_42898,N_42899,N_42900,N_42901,N_42902,N_42903,N_42904,N_42905,N_42906,N_42907,N_42908,N_42909,N_42910,N_42911,N_42912,N_42913,N_42914,N_42915,N_42916,N_42917,N_42918,N_42919,N_42920,N_42921,N_42922,N_42923,N_42924,N_42925,N_42926,N_42927,N_42928,N_42929,N_42930,N_42931,N_42932,N_42933,N_42934,N_42935,N_42936,N_42937,N_42938,N_42939,N_42940,N_42941,N_42942,N_42943,N_42944,N_42945,N_42946,N_42947,N_42948,N_42949,N_42950,N_42951,N_42952,N_42953,N_42954,N_42955,N_42956,N_42957,N_42958,N_42959,N_42960,N_42961,N_42962,N_42963,N_42964,N_42965,N_42966,N_42967,N_42968,N_42969,N_42970,N_42971,N_42972,N_42973,N_42974,N_42975,N_42976,N_42977,N_42978,N_42979,N_42980,N_42981,N_42982,N_42983,N_42984,N_42985,N_42986,N_42987,N_42988,N_42989,N_42990,N_42991,N_42992,N_42993,N_42994,N_42995,N_42996,N_42997,N_42998,N_42999,N_43000,N_43001,N_43002,N_43003,N_43004,N_43005,N_43006,N_43007,N_43008,N_43009,N_43010,N_43011,N_43012,N_43013,N_43014,N_43015,N_43016,N_43017,N_43018,N_43019,N_43020,N_43021,N_43022,N_43023,N_43024,N_43025,N_43026,N_43027,N_43028,N_43029,N_43030,N_43031,N_43032,N_43033,N_43034,N_43035,N_43036,N_43037,N_43038,N_43039,N_43040,N_43041,N_43042,N_43043,N_43044,N_43045,N_43046,N_43047,N_43048,N_43049,N_43050,N_43051,N_43052,N_43053,N_43054,N_43055,N_43056,N_43057,N_43058,N_43059,N_43060,N_43061,N_43062,N_43063,N_43064,N_43065,N_43066,N_43067,N_43068,N_43069,N_43070,N_43071,N_43072,N_43073,N_43074,N_43075,N_43076,N_43077,N_43078,N_43079,N_43080,N_43081,N_43082,N_43083,N_43084,N_43085,N_43086,N_43087,N_43088,N_43089,N_43090,N_43091,N_43092,N_43093,N_43094,N_43095,N_43096,N_43097,N_43098,N_43099,N_43100,N_43101,N_43102,N_43103,N_43104,N_43105,N_43106,N_43107,N_43108,N_43109,N_43110,N_43111,N_43112,N_43113,N_43114,N_43115,N_43116,N_43117,N_43118,N_43119,N_43120,N_43121,N_43122,N_43123,N_43124,N_43125,N_43126,N_43127,N_43128,N_43129,N_43130,N_43131,N_43132,N_43133,N_43134,N_43135,N_43136,N_43137,N_43138,N_43139,N_43140,N_43141,N_43142,N_43143,N_43144,N_43145,N_43146,N_43147,N_43148,N_43149,N_43150,N_43151,N_43152,N_43153,N_43154,N_43155,N_43156,N_43157,N_43158,N_43159,N_43160,N_43161,N_43162,N_43163,N_43164,N_43165,N_43166,N_43167,N_43168,N_43169,N_43170,N_43171,N_43172,N_43173,N_43174,N_43175,N_43176,N_43177,N_43178,N_43179,N_43180,N_43181,N_43182,N_43183,N_43184,N_43185,N_43186,N_43187,N_43188,N_43189,N_43190,N_43191,N_43192,N_43193,N_43194,N_43195,N_43196,N_43197,N_43198,N_43199,N_43200,N_43201,N_43202,N_43203,N_43204,N_43205,N_43206,N_43207,N_43208,N_43209,N_43210,N_43211,N_43212,N_43213,N_43214,N_43215,N_43216,N_43217,N_43218,N_43219,N_43220,N_43221,N_43222,N_43223,N_43224,N_43225,N_43226,N_43227,N_43228,N_43229,N_43230,N_43231,N_43232,N_43233,N_43234,N_43235,N_43236,N_43237,N_43238,N_43239,N_43240,N_43241,N_43242,N_43243,N_43244,N_43245,N_43246,N_43247,N_43248,N_43249,N_43250,N_43251,N_43252,N_43253,N_43254,N_43255,N_43256,N_43257,N_43258,N_43259,N_43260,N_43261,N_43262,N_43263,N_43264,N_43265,N_43266,N_43267,N_43268,N_43269,N_43270,N_43271,N_43272,N_43273,N_43274,N_43275,N_43276,N_43277,N_43278,N_43279,N_43280,N_43281,N_43282,N_43283,N_43284,N_43285,N_43286,N_43287,N_43288,N_43289,N_43290,N_43291,N_43292,N_43293,N_43294,N_43295,N_43296,N_43297,N_43298,N_43299,N_43300,N_43301,N_43302,N_43303,N_43304,N_43305,N_43306,N_43307,N_43308,N_43309,N_43310,N_43311,N_43312,N_43313,N_43314,N_43315,N_43316,N_43317,N_43318,N_43319,N_43320,N_43321,N_43322,N_43323,N_43324,N_43325,N_43326,N_43327,N_43328,N_43329,N_43330,N_43331,N_43332,N_43333,N_43334,N_43335,N_43336,N_43337,N_43338,N_43339,N_43340,N_43341,N_43342,N_43343,N_43344,N_43345,N_43346,N_43347,N_43348,N_43349,N_43350,N_43351,N_43352,N_43353,N_43354,N_43355,N_43356,N_43357,N_43358,N_43359,N_43360,N_43361,N_43362,N_43363,N_43364,N_43365,N_43366,N_43367,N_43368,N_43369,N_43370,N_43371,N_43372,N_43373,N_43374,N_43375,N_43376,N_43377,N_43378,N_43379,N_43380,N_43381,N_43382,N_43383,N_43384,N_43385,N_43386,N_43387,N_43388,N_43389,N_43390,N_43391,N_43392,N_43393,N_43394,N_43395,N_43396,N_43397,N_43398,N_43399,N_43400,N_43401,N_43402,N_43403,N_43404,N_43405,N_43406,N_43407,N_43408,N_43409,N_43410,N_43411,N_43412,N_43413,N_43414,N_43415,N_43416,N_43417,N_43418,N_43419,N_43420,N_43421,N_43422,N_43423,N_43424,N_43425,N_43426,N_43427,N_43428,N_43429,N_43430,N_43431,N_43432,N_43433,N_43434,N_43435,N_43436,N_43437,N_43438,N_43439,N_43440,N_43441,N_43442,N_43443,N_43444,N_43445,N_43446,N_43447,N_43448,N_43449,N_43450,N_43451,N_43452,N_43453,N_43454,N_43455,N_43456,N_43457,N_43458,N_43459,N_43460,N_43461,N_43462,N_43463,N_43464,N_43465,N_43466,N_43467,N_43468,N_43469,N_43470,N_43471,N_43472,N_43473,N_43474,N_43475,N_43476,N_43477,N_43478,N_43479,N_43480,N_43481,N_43482,N_43483,N_43484,N_43485,N_43486,N_43487,N_43488,N_43489,N_43490,N_43491,N_43492,N_43493,N_43494,N_43495,N_43496,N_43497,N_43498,N_43499,N_43500,N_43501,N_43502,N_43503,N_43504,N_43505,N_43506,N_43507,N_43508,N_43509,N_43510,N_43511,N_43512,N_43513,N_43514,N_43515,N_43516,N_43517,N_43518,N_43519,N_43520,N_43521,N_43522,N_43523,N_43524,N_43525,N_43526,N_43527,N_43528,N_43529,N_43530,N_43531,N_43532,N_43533,N_43534,N_43535,N_43536,N_43537,N_43538,N_43539,N_43540,N_43541,N_43542,N_43543,N_43544,N_43545,N_43546,N_43547,N_43548,N_43549,N_43550,N_43551,N_43552,N_43553,N_43554,N_43555,N_43556,N_43557,N_43558,N_43559,N_43560,N_43561,N_43562,N_43563,N_43564,N_43565,N_43566,N_43567,N_43568,N_43569,N_43570,N_43571,N_43572,N_43573,N_43574,N_43575,N_43576,N_43577,N_43578,N_43579,N_43580,N_43581,N_43582,N_43583,N_43584,N_43585,N_43586,N_43587,N_43588,N_43589,N_43590,N_43591,N_43592,N_43593,N_43594,N_43595,N_43596,N_43597,N_43598,N_43599,N_43600,N_43601,N_43602,N_43603,N_43604,N_43605,N_43606,N_43607,N_43608,N_43609,N_43610,N_43611,N_43612,N_43613,N_43614,N_43615,N_43616,N_43617,N_43618,N_43619,N_43620,N_43621,N_43622,N_43623,N_43624,N_43625,N_43626,N_43627,N_43628,N_43629,N_43630,N_43631,N_43632,N_43633,N_43634,N_43635,N_43636,N_43637,N_43638,N_43639,N_43640,N_43641,N_43642,N_43643,N_43644,N_43645,N_43646,N_43647,N_43648,N_43649,N_43650,N_43651,N_43652,N_43653,N_43654,N_43655,N_43656,N_43657,N_43658,N_43659,N_43660,N_43661,N_43662,N_43663,N_43664,N_43665,N_43666,N_43667,N_43668,N_43669,N_43670,N_43671,N_43672,N_43673,N_43674,N_43675,N_43676,N_43677,N_43678,N_43679,N_43680,N_43681,N_43682,N_43683,N_43684,N_43685,N_43686,N_43687,N_43688,N_43689,N_43690,N_43691,N_43692,N_43693,N_43694,N_43695,N_43696,N_43697,N_43698,N_43699,N_43700,N_43701,N_43702,N_43703,N_43704,N_43705,N_43706,N_43707,N_43708,N_43709,N_43710,N_43711,N_43712,N_43713,N_43714,N_43715,N_43716,N_43717,N_43718,N_43719,N_43720,N_43721,N_43722,N_43723,N_43724,N_43725,N_43726,N_43727,N_43728,N_43729,N_43730,N_43731,N_43732,N_43733,N_43734,N_43735,N_43736,N_43737,N_43738,N_43739,N_43740,N_43741,N_43742,N_43743,N_43744,N_43745,N_43746,N_43747,N_43748,N_43749,N_43750,N_43751,N_43752,N_43753,N_43754,N_43755,N_43756,N_43757,N_43758,N_43759,N_43760,N_43761,N_43762,N_43763,N_43764,N_43765,N_43766,N_43767,N_43768,N_43769,N_43770,N_43771,N_43772,N_43773,N_43774,N_43775,N_43776,N_43777,N_43778,N_43779,N_43780,N_43781,N_43782,N_43783,N_43784,N_43785,N_43786,N_43787,N_43788,N_43789,N_43790,N_43791,N_43792,N_43793,N_43794,N_43795,N_43796,N_43797,N_43798,N_43799,N_43800,N_43801,N_43802,N_43803,N_43804,N_43805,N_43806,N_43807,N_43808,N_43809,N_43810,N_43811,N_43812,N_43813,N_43814,N_43815,N_43816,N_43817,N_43818,N_43819,N_43820,N_43821,N_43822,N_43823,N_43824,N_43825,N_43826,N_43827,N_43828,N_43829,N_43830,N_43831,N_43832,N_43833,N_43834,N_43835,N_43836,N_43837,N_43838,N_43839,N_43840,N_43841,N_43842,N_43843,N_43844,N_43845,N_43846,N_43847,N_43848,N_43849,N_43850,N_43851,N_43852,N_43853,N_43854,N_43855,N_43856,N_43857,N_43858,N_43859,N_43860,N_43861,N_43862,N_43863,N_43864,N_43865,N_43866,N_43867,N_43868,N_43869,N_43870,N_43871,N_43872,N_43873,N_43874,N_43875,N_43876,N_43877,N_43878,N_43879,N_43880,N_43881,N_43882,N_43883,N_43884,N_43885,N_43886,N_43887,N_43888,N_43889,N_43890,N_43891,N_43892,N_43893,N_43894,N_43895,N_43896,N_43897,N_43898,N_43899,N_43900,N_43901,N_43902,N_43903,N_43904,N_43905,N_43906,N_43907,N_43908,N_43909,N_43910,N_43911,N_43912,N_43913,N_43914,N_43915,N_43916,N_43917,N_43918,N_43919,N_43920,N_43921,N_43922,N_43923,N_43924,N_43925,N_43926,N_43927,N_43928,N_43929,N_43930,N_43931,N_43932,N_43933,N_43934,N_43935,N_43936,N_43937,N_43938,N_43939,N_43940,N_43941,N_43942,N_43943,N_43944,N_43945,N_43946,N_43947,N_43948,N_43949,N_43950,N_43951,N_43952,N_43953,N_43954,N_43955,N_43956,N_43957,N_43958,N_43959,N_43960,N_43961,N_43962,N_43963,N_43964,N_43965,N_43966,N_43967,N_43968,N_43969,N_43970,N_43971,N_43972,N_43973,N_43974,N_43975,N_43976,N_43977,N_43978,N_43979,N_43980,N_43981,N_43982,N_43983,N_43984,N_43985,N_43986,N_43987,N_43988,N_43989,N_43990,N_43991,N_43992,N_43993,N_43994,N_43995,N_43996,N_43997,N_43998,N_43999,N_44000,N_44001,N_44002,N_44003,N_44004,N_44005,N_44006,N_44007,N_44008,N_44009,N_44010,N_44011,N_44012,N_44013,N_44014,N_44015,N_44016,N_44017,N_44018,N_44019,N_44020,N_44021,N_44022,N_44023,N_44024,N_44025,N_44026,N_44027,N_44028,N_44029,N_44030,N_44031,N_44032,N_44033,N_44034,N_44035,N_44036,N_44037,N_44038,N_44039,N_44040,N_44041,N_44042,N_44043,N_44044,N_44045,N_44046,N_44047,N_44048,N_44049,N_44050,N_44051,N_44052,N_44053,N_44054,N_44055,N_44056,N_44057,N_44058,N_44059,N_44060,N_44061,N_44062,N_44063,N_44064,N_44065,N_44066,N_44067,N_44068,N_44069,N_44070,N_44071,N_44072,N_44073,N_44074,N_44075,N_44076,N_44077,N_44078,N_44079,N_44080,N_44081,N_44082,N_44083,N_44084,N_44085,N_44086,N_44087,N_44088,N_44089,N_44090,N_44091,N_44092,N_44093,N_44094,N_44095,N_44096,N_44097,N_44098,N_44099,N_44100,N_44101,N_44102,N_44103,N_44104,N_44105,N_44106,N_44107,N_44108,N_44109,N_44110,N_44111,N_44112,N_44113,N_44114,N_44115,N_44116,N_44117,N_44118,N_44119,N_44120,N_44121,N_44122,N_44123,N_44124,N_44125,N_44126,N_44127,N_44128,N_44129,N_44130,N_44131,N_44132,N_44133,N_44134,N_44135,N_44136,N_44137,N_44138,N_44139,N_44140,N_44141,N_44142,N_44143,N_44144,N_44145,N_44146,N_44147,N_44148,N_44149,N_44150,N_44151,N_44152,N_44153,N_44154,N_44155,N_44156,N_44157,N_44158,N_44159,N_44160,N_44161,N_44162,N_44163,N_44164,N_44165,N_44166,N_44167,N_44168,N_44169,N_44170,N_44171,N_44172,N_44173,N_44174,N_44175,N_44176,N_44177,N_44178,N_44179,N_44180,N_44181,N_44182,N_44183,N_44184,N_44185,N_44186,N_44187,N_44188,N_44189,N_44190,N_44191,N_44192,N_44193,N_44194,N_44195,N_44196,N_44197,N_44198,N_44199,N_44200,N_44201,N_44202,N_44203,N_44204,N_44205,N_44206,N_44207,N_44208,N_44209,N_44210,N_44211,N_44212,N_44213,N_44214,N_44215,N_44216,N_44217,N_44218,N_44219,N_44220,N_44221,N_44222,N_44223,N_44224,N_44225,N_44226,N_44227,N_44228,N_44229,N_44230,N_44231,N_44232,N_44233,N_44234,N_44235,N_44236,N_44237,N_44238,N_44239,N_44240,N_44241,N_44242,N_44243,N_44244,N_44245,N_44246,N_44247,N_44248,N_44249,N_44250,N_44251,N_44252,N_44253,N_44254,N_44255,N_44256,N_44257,N_44258,N_44259,N_44260,N_44261,N_44262,N_44263,N_44264,N_44265,N_44266,N_44267,N_44268,N_44269,N_44270,N_44271,N_44272,N_44273,N_44274,N_44275,N_44276,N_44277,N_44278,N_44279,N_44280,N_44281,N_44282,N_44283,N_44284,N_44285,N_44286,N_44287,N_44288,N_44289,N_44290,N_44291,N_44292,N_44293,N_44294,N_44295,N_44296,N_44297,N_44298,N_44299,N_44300,N_44301,N_44302,N_44303,N_44304,N_44305,N_44306,N_44307,N_44308,N_44309,N_44310,N_44311,N_44312,N_44313,N_44314,N_44315,N_44316,N_44317,N_44318,N_44319,N_44320,N_44321,N_44322,N_44323,N_44324,N_44325,N_44326,N_44327,N_44328,N_44329,N_44330,N_44331,N_44332,N_44333,N_44334,N_44335,N_44336,N_44337,N_44338,N_44339,N_44340,N_44341,N_44342,N_44343,N_44344,N_44345,N_44346,N_44347,N_44348,N_44349,N_44350,N_44351,N_44352,N_44353,N_44354,N_44355,N_44356,N_44357,N_44358,N_44359,N_44360,N_44361,N_44362,N_44363,N_44364,N_44365,N_44366,N_44367,N_44368,N_44369,N_44370,N_44371,N_44372,N_44373,N_44374,N_44375,N_44376,N_44377,N_44378,N_44379,N_44380,N_44381,N_44382,N_44383,N_44384,N_44385,N_44386,N_44387,N_44388,N_44389,N_44390,N_44391,N_44392,N_44393,N_44394,N_44395,N_44396,N_44397,N_44398,N_44399,N_44400,N_44401,N_44402,N_44403,N_44404,N_44405,N_44406,N_44407,N_44408,N_44409,N_44410,N_44411,N_44412,N_44413,N_44414,N_44415,N_44416,N_44417,N_44418,N_44419,N_44420,N_44421,N_44422,N_44423,N_44424,N_44425,N_44426,N_44427,N_44428,N_44429,N_44430,N_44431,N_44432,N_44433,N_44434,N_44435,N_44436,N_44437,N_44438,N_44439,N_44440,N_44441,N_44442,N_44443,N_44444,N_44445,N_44446,N_44447,N_44448,N_44449,N_44450,N_44451,N_44452,N_44453,N_44454,N_44455,N_44456,N_44457,N_44458,N_44459,N_44460,N_44461,N_44462,N_44463,N_44464,N_44465,N_44466,N_44467,N_44468,N_44469,N_44470,N_44471,N_44472,N_44473,N_44474,N_44475,N_44476,N_44477,N_44478,N_44479,N_44480,N_44481,N_44482,N_44483,N_44484,N_44485,N_44486,N_44487,N_44488,N_44489,N_44490,N_44491,N_44492,N_44493,N_44494,N_44495,N_44496,N_44497,N_44498,N_44499,N_44500,N_44501,N_44502,N_44503,N_44504,N_44505,N_44506,N_44507,N_44508,N_44509,N_44510,N_44511,N_44512,N_44513,N_44514,N_44515,N_44516,N_44517,N_44518,N_44519,N_44520,N_44521,N_44522,N_44523,N_44524,N_44525,N_44526,N_44527,N_44528,N_44529,N_44530,N_44531,N_44532,N_44533,N_44534,N_44535,N_44536,N_44537,N_44538,N_44539,N_44540,N_44541,N_44542,N_44543,N_44544,N_44545,N_44546,N_44547,N_44548,N_44549,N_44550,N_44551,N_44552,N_44553,N_44554,N_44555,N_44556,N_44557,N_44558,N_44559,N_44560,N_44561,N_44562,N_44563,N_44564,N_44565,N_44566,N_44567,N_44568,N_44569,N_44570,N_44571,N_44572,N_44573,N_44574,N_44575,N_44576,N_44577,N_44578,N_44579,N_44580,N_44581,N_44582,N_44583,N_44584,N_44585,N_44586,N_44587,N_44588,N_44589,N_44590,N_44591,N_44592,N_44593,N_44594,N_44595,N_44596,N_44597,N_44598,N_44599,N_44600,N_44601,N_44602,N_44603,N_44604,N_44605,N_44606,N_44607,N_44608,N_44609,N_44610,N_44611,N_44612,N_44613,N_44614,N_44615,N_44616,N_44617,N_44618,N_44619,N_44620,N_44621,N_44622,N_44623,N_44624,N_44625,N_44626,N_44627,N_44628,N_44629,N_44630,N_44631,N_44632,N_44633,N_44634,N_44635,N_44636,N_44637,N_44638,N_44639,N_44640,N_44641,N_44642,N_44643,N_44644,N_44645,N_44646,N_44647,N_44648,N_44649,N_44650,N_44651,N_44652,N_44653,N_44654,N_44655,N_44656,N_44657,N_44658,N_44659,N_44660,N_44661,N_44662,N_44663,N_44664,N_44665,N_44666,N_44667,N_44668,N_44669,N_44670,N_44671,N_44672,N_44673,N_44674,N_44675,N_44676,N_44677,N_44678,N_44679,N_44680,N_44681,N_44682,N_44683,N_44684,N_44685,N_44686,N_44687,N_44688,N_44689,N_44690,N_44691,N_44692,N_44693,N_44694,N_44695,N_44696,N_44697,N_44698,N_44699,N_44700,N_44701,N_44702,N_44703,N_44704,N_44705,N_44706,N_44707,N_44708,N_44709,N_44710,N_44711,N_44712,N_44713,N_44714,N_44715,N_44716,N_44717,N_44718,N_44719,N_44720,N_44721,N_44722,N_44723,N_44724,N_44725,N_44726,N_44727,N_44728,N_44729,N_44730,N_44731,N_44732,N_44733,N_44734,N_44735,N_44736,N_44737,N_44738,N_44739,N_44740,N_44741,N_44742,N_44743,N_44744,N_44745,N_44746,N_44747,N_44748,N_44749,N_44750,N_44751,N_44752,N_44753,N_44754,N_44755,N_44756,N_44757,N_44758,N_44759,N_44760,N_44761,N_44762,N_44763,N_44764,N_44765,N_44766,N_44767,N_44768,N_44769,N_44770,N_44771,N_44772,N_44773,N_44774,N_44775,N_44776,N_44777,N_44778,N_44779,N_44780,N_44781,N_44782,N_44783,N_44784,N_44785,N_44786,N_44787,N_44788,N_44789,N_44790,N_44791,N_44792,N_44793,N_44794,N_44795,N_44796,N_44797,N_44798,N_44799,N_44800,N_44801,N_44802,N_44803,N_44804,N_44805,N_44806,N_44807,N_44808,N_44809,N_44810,N_44811,N_44812,N_44813,N_44814,N_44815,N_44816,N_44817,N_44818,N_44819,N_44820,N_44821,N_44822,N_44823,N_44824,N_44825,N_44826,N_44827,N_44828,N_44829,N_44830,N_44831,N_44832,N_44833,N_44834,N_44835,N_44836,N_44837,N_44838,N_44839,N_44840,N_44841,N_44842,N_44843,N_44844,N_44845,N_44846,N_44847,N_44848,N_44849,N_44850,N_44851,N_44852,N_44853,N_44854,N_44855,N_44856,N_44857,N_44858,N_44859,N_44860,N_44861,N_44862,N_44863,N_44864,N_44865,N_44866,N_44867,N_44868,N_44869,N_44870,N_44871,N_44872,N_44873,N_44874,N_44875,N_44876,N_44877,N_44878,N_44879,N_44880,N_44881,N_44882,N_44883,N_44884,N_44885,N_44886,N_44887,N_44888,N_44889,N_44890,N_44891,N_44892,N_44893,N_44894,N_44895,N_44896,N_44897,N_44898,N_44899,N_44900,N_44901,N_44902,N_44903,N_44904,N_44905,N_44906,N_44907,N_44908,N_44909,N_44910,N_44911,N_44912,N_44913,N_44914,N_44915,N_44916,N_44917,N_44918,N_44919,N_44920,N_44921,N_44922,N_44923,N_44924,N_44925,N_44926,N_44927,N_44928,N_44929,N_44930,N_44931,N_44932,N_44933,N_44934,N_44935,N_44936,N_44937,N_44938,N_44939,N_44940,N_44941,N_44942,N_44943,N_44944,N_44945,N_44946,N_44947,N_44948,N_44949,N_44950,N_44951,N_44952,N_44953,N_44954,N_44955,N_44956,N_44957,N_44958,N_44959,N_44960,N_44961,N_44962,N_44963,N_44964,N_44965,N_44966,N_44967,N_44968,N_44969,N_44970,N_44971,N_44972,N_44973,N_44974,N_44975,N_44976,N_44977,N_44978,N_44979,N_44980,N_44981,N_44982,N_44983,N_44984,N_44985,N_44986,N_44987,N_44988,N_44989,N_44990,N_44991,N_44992,N_44993,N_44994,N_44995,N_44996,N_44997,N_44998,N_44999,N_45000,N_45001,N_45002,N_45003,N_45004,N_45005,N_45006,N_45007,N_45008,N_45009,N_45010,N_45011,N_45012,N_45013,N_45014,N_45015,N_45016,N_45017,N_45018,N_45019,N_45020,N_45021,N_45022,N_45023,N_45024,N_45025,N_45026,N_45027,N_45028,N_45029,N_45030,N_45031,N_45032,N_45033,N_45034,N_45035,N_45036,N_45037,N_45038,N_45039,N_45040,N_45041,N_45042,N_45043,N_45044,N_45045,N_45046,N_45047,N_45048,N_45049,N_45050,N_45051,N_45052,N_45053,N_45054,N_45055,N_45056,N_45057,N_45058,N_45059,N_45060,N_45061,N_45062,N_45063,N_45064,N_45065,N_45066,N_45067,N_45068,N_45069,N_45070,N_45071,N_45072,N_45073,N_45074,N_45075,N_45076,N_45077,N_45078,N_45079,N_45080,N_45081,N_45082,N_45083,N_45084,N_45085,N_45086,N_45087,N_45088,N_45089,N_45090,N_45091,N_45092,N_45093,N_45094,N_45095,N_45096,N_45097,N_45098,N_45099,N_45100,N_45101,N_45102,N_45103,N_45104,N_45105,N_45106,N_45107,N_45108,N_45109,N_45110,N_45111,N_45112,N_45113,N_45114,N_45115,N_45116,N_45117,N_45118,N_45119,N_45120,N_45121,N_45122,N_45123,N_45124,N_45125,N_45126,N_45127,N_45128,N_45129,N_45130,N_45131,N_45132,N_45133,N_45134,N_45135,N_45136,N_45137,N_45138,N_45139,N_45140,N_45141,N_45142,N_45143,N_45144,N_45145,N_45146,N_45147,N_45148,N_45149,N_45150,N_45151,N_45152,N_45153,N_45154,N_45155,N_45156,N_45157,N_45158,N_45159,N_45160,N_45161,N_45162,N_45163,N_45164,N_45165,N_45166,N_45167,N_45168,N_45169,N_45170,N_45171,N_45172,N_45173,N_45174,N_45175,N_45176,N_45177,N_45178,N_45179,N_45180,N_45181,N_45182,N_45183,N_45184,N_45185,N_45186,N_45187,N_45188,N_45189,N_45190,N_45191,N_45192,N_45193,N_45194,N_45195,N_45196,N_45197,N_45198,N_45199,N_45200,N_45201,N_45202,N_45203,N_45204,N_45205,N_45206,N_45207,N_45208,N_45209,N_45210,N_45211,N_45212,N_45213,N_45214,N_45215,N_45216,N_45217,N_45218,N_45219,N_45220,N_45221,N_45222,N_45223,N_45224,N_45225,N_45226,N_45227,N_45228,N_45229,N_45230,N_45231,N_45232,N_45233,N_45234,N_45235,N_45236,N_45237,N_45238,N_45239,N_45240,N_45241,N_45242,N_45243,N_45244,N_45245,N_45246,N_45247,N_45248,N_45249,N_45250,N_45251,N_45252,N_45253,N_45254,N_45255,N_45256,N_45257,N_45258,N_45259,N_45260,N_45261,N_45262,N_45263,N_45264,N_45265,N_45266,N_45267,N_45268,N_45269,N_45270,N_45271,N_45272,N_45273,N_45274,N_45275,N_45276,N_45277,N_45278,N_45279,N_45280,N_45281,N_45282,N_45283,N_45284,N_45285,N_45286,N_45287,N_45288,N_45289,N_45290,N_45291,N_45292,N_45293,N_45294,N_45295,N_45296,N_45297,N_45298,N_45299,N_45300,N_45301,N_45302,N_45303,N_45304,N_45305,N_45306,N_45307,N_45308,N_45309,N_45310,N_45311,N_45312,N_45313,N_45314,N_45315,N_45316,N_45317,N_45318,N_45319,N_45320,N_45321,N_45322,N_45323,N_45324,N_45325,N_45326,N_45327,N_45328,N_45329,N_45330,N_45331,N_45332,N_45333,N_45334,N_45335,N_45336,N_45337,N_45338,N_45339,N_45340,N_45341,N_45342,N_45343,N_45344,N_45345,N_45346,N_45347,N_45348,N_45349,N_45350,N_45351,N_45352,N_45353,N_45354,N_45355,N_45356,N_45357,N_45358,N_45359,N_45360,N_45361,N_45362,N_45363,N_45364,N_45365,N_45366,N_45367,N_45368,N_45369,N_45370,N_45371,N_45372,N_45373,N_45374,N_45375,N_45376,N_45377,N_45378,N_45379,N_45380,N_45381,N_45382,N_45383,N_45384,N_45385,N_45386,N_45387,N_45388,N_45389,N_45390,N_45391,N_45392,N_45393,N_45394,N_45395,N_45396,N_45397,N_45398,N_45399,N_45400,N_45401,N_45402,N_45403,N_45404,N_45405,N_45406,N_45407,N_45408,N_45409,N_45410,N_45411,N_45412,N_45413,N_45414,N_45415,N_45416,N_45417,N_45418,N_45419,N_45420,N_45421,N_45422,N_45423,N_45424,N_45425,N_45426,N_45427,N_45428,N_45429,N_45430,N_45431,N_45432,N_45433,N_45434,N_45435,N_45436,N_45437,N_45438,N_45439,N_45440,N_45441,N_45442,N_45443,N_45444,N_45445,N_45446,N_45447,N_45448,N_45449,N_45450,N_45451,N_45452,N_45453,N_45454,N_45455,N_45456,N_45457,N_45458,N_45459,N_45460,N_45461,N_45462,N_45463,N_45464,N_45465,N_45466,N_45467,N_45468,N_45469,N_45470,N_45471,N_45472,N_45473,N_45474,N_45475,N_45476,N_45477,N_45478,N_45479,N_45480,N_45481,N_45482,N_45483,N_45484,N_45485,N_45486,N_45487,N_45488,N_45489,N_45490,N_45491,N_45492,N_45493,N_45494,N_45495,N_45496,N_45497,N_45498,N_45499,N_45500,N_45501,N_45502,N_45503,N_45504,N_45505,N_45506,N_45507,N_45508,N_45509,N_45510,N_45511,N_45512,N_45513,N_45514,N_45515,N_45516,N_45517,N_45518,N_45519,N_45520,N_45521,N_45522,N_45523,N_45524,N_45525,N_45526,N_45527,N_45528,N_45529,N_45530,N_45531,N_45532,N_45533,N_45534,N_45535,N_45536,N_45537,N_45538,N_45539,N_45540,N_45541,N_45542,N_45543,N_45544,N_45545,N_45546,N_45547,N_45548,N_45549,N_45550,N_45551,N_45552,N_45553,N_45554,N_45555,N_45556,N_45557,N_45558,N_45559,N_45560,N_45561,N_45562,N_45563,N_45564,N_45565,N_45566,N_45567,N_45568,N_45569,N_45570,N_45571,N_45572,N_45573,N_45574,N_45575,N_45576,N_45577,N_45578,N_45579,N_45580,N_45581,N_45582,N_45583,N_45584,N_45585,N_45586,N_45587,N_45588,N_45589,N_45590,N_45591,N_45592,N_45593,N_45594,N_45595,N_45596,N_45597,N_45598,N_45599,N_45600,N_45601,N_45602,N_45603,N_45604,N_45605,N_45606,N_45607,N_45608,N_45609,N_45610,N_45611,N_45612,N_45613,N_45614,N_45615,N_45616,N_45617,N_45618,N_45619,N_45620,N_45621,N_45622,N_45623,N_45624,N_45625,N_45626,N_45627,N_45628,N_45629,N_45630,N_45631,N_45632,N_45633,N_45634,N_45635,N_45636,N_45637,N_45638,N_45639,N_45640,N_45641,N_45642,N_45643,N_45644,N_45645,N_45646,N_45647,N_45648,N_45649,N_45650,N_45651,N_45652,N_45653,N_45654,N_45655,N_45656,N_45657,N_45658,N_45659,N_45660,N_45661,N_45662,N_45663,N_45664,N_45665,N_45666,N_45667,N_45668,N_45669,N_45670,N_45671,N_45672,N_45673,N_45674,N_45675,N_45676,N_45677,N_45678,N_45679,N_45680,N_45681,N_45682,N_45683,N_45684,N_45685,N_45686,N_45687,N_45688,N_45689,N_45690,N_45691,N_45692,N_45693,N_45694,N_45695,N_45696,N_45697,N_45698,N_45699,N_45700,N_45701,N_45702,N_45703,N_45704,N_45705,N_45706,N_45707,N_45708,N_45709,N_45710,N_45711,N_45712,N_45713,N_45714,N_45715,N_45716,N_45717,N_45718,N_45719,N_45720,N_45721,N_45722,N_45723,N_45724,N_45725,N_45726,N_45727,N_45728,N_45729,N_45730,N_45731,N_45732,N_45733,N_45734,N_45735,N_45736,N_45737,N_45738,N_45739,N_45740,N_45741,N_45742,N_45743,N_45744,N_45745,N_45746,N_45747,N_45748,N_45749,N_45750,N_45751,N_45752,N_45753,N_45754,N_45755,N_45756,N_45757,N_45758,N_45759,N_45760,N_45761,N_45762,N_45763,N_45764,N_45765,N_45766,N_45767,N_45768,N_45769,N_45770,N_45771,N_45772,N_45773,N_45774,N_45775,N_45776,N_45777,N_45778,N_45779,N_45780,N_45781,N_45782,N_45783,N_45784,N_45785,N_45786,N_45787,N_45788,N_45789,N_45790,N_45791,N_45792,N_45793,N_45794,N_45795,N_45796,N_45797,N_45798,N_45799,N_45800,N_45801,N_45802,N_45803,N_45804,N_45805,N_45806,N_45807,N_45808,N_45809,N_45810,N_45811,N_45812,N_45813,N_45814,N_45815,N_45816,N_45817,N_45818,N_45819,N_45820,N_45821,N_45822,N_45823,N_45824,N_45825,N_45826,N_45827,N_45828,N_45829,N_45830,N_45831,N_45832,N_45833,N_45834,N_45835,N_45836,N_45837,N_45838,N_45839,N_45840,N_45841,N_45842,N_45843,N_45844,N_45845,N_45846,N_45847,N_45848,N_45849,N_45850,N_45851,N_45852,N_45853,N_45854,N_45855,N_45856,N_45857,N_45858,N_45859,N_45860,N_45861,N_45862,N_45863,N_45864,N_45865,N_45866,N_45867,N_45868,N_45869,N_45870,N_45871,N_45872,N_45873,N_45874,N_45875,N_45876,N_45877,N_45878,N_45879,N_45880,N_45881,N_45882,N_45883,N_45884,N_45885,N_45886,N_45887,N_45888,N_45889,N_45890,N_45891,N_45892,N_45893,N_45894,N_45895,N_45896,N_45897,N_45898,N_45899,N_45900,N_45901,N_45902,N_45903,N_45904,N_45905,N_45906,N_45907,N_45908,N_45909,N_45910,N_45911,N_45912,N_45913,N_45914,N_45915,N_45916,N_45917,N_45918,N_45919,N_45920,N_45921,N_45922,N_45923,N_45924,N_45925,N_45926,N_45927,N_45928,N_45929,N_45930,N_45931,N_45932,N_45933,N_45934,N_45935,N_45936,N_45937,N_45938,N_45939,N_45940,N_45941,N_45942,N_45943,N_45944,N_45945,N_45946,N_45947,N_45948,N_45949,N_45950,N_45951,N_45952,N_45953,N_45954,N_45955,N_45956,N_45957,N_45958,N_45959,N_45960,N_45961,N_45962,N_45963,N_45964,N_45965,N_45966,N_45967,N_45968,N_45969,N_45970,N_45971,N_45972,N_45973,N_45974,N_45975,N_45976,N_45977,N_45978,N_45979,N_45980,N_45981,N_45982,N_45983,N_45984,N_45985,N_45986,N_45987,N_45988,N_45989,N_45990,N_45991,N_45992,N_45993,N_45994,N_45995,N_45996,N_45997,N_45998,N_45999,N_46000,N_46001,N_46002,N_46003,N_46004,N_46005,N_46006,N_46007,N_46008,N_46009,N_46010,N_46011,N_46012,N_46013,N_46014,N_46015,N_46016,N_46017,N_46018,N_46019,N_46020,N_46021,N_46022,N_46023,N_46024,N_46025,N_46026,N_46027,N_46028,N_46029,N_46030,N_46031,N_46032,N_46033,N_46034,N_46035,N_46036,N_46037,N_46038,N_46039,N_46040,N_46041,N_46042,N_46043,N_46044,N_46045,N_46046,N_46047,N_46048,N_46049,N_46050,N_46051,N_46052,N_46053,N_46054,N_46055,N_46056,N_46057,N_46058,N_46059,N_46060,N_46061,N_46062,N_46063,N_46064,N_46065,N_46066,N_46067,N_46068,N_46069,N_46070,N_46071,N_46072,N_46073,N_46074,N_46075,N_46076,N_46077,N_46078,N_46079,N_46080,N_46081,N_46082,N_46083,N_46084,N_46085,N_46086,N_46087,N_46088,N_46089,N_46090,N_46091,N_46092,N_46093,N_46094,N_46095,N_46096,N_46097,N_46098,N_46099,N_46100,N_46101,N_46102,N_46103,N_46104,N_46105,N_46106,N_46107,N_46108,N_46109,N_46110,N_46111,N_46112,N_46113,N_46114,N_46115,N_46116,N_46117,N_46118,N_46119,N_46120,N_46121,N_46122,N_46123,N_46124,N_46125,N_46126,N_46127,N_46128,N_46129,N_46130,N_46131,N_46132,N_46133,N_46134,N_46135,N_46136,N_46137,N_46138,N_46139,N_46140,N_46141,N_46142,N_46143,N_46144,N_46145,N_46146,N_46147,N_46148,N_46149,N_46150,N_46151,N_46152,N_46153,N_46154,N_46155,N_46156,N_46157,N_46158,N_46159,N_46160,N_46161,N_46162,N_46163,N_46164,N_46165,N_46166,N_46167,N_46168,N_46169,N_46170,N_46171,N_46172,N_46173,N_46174,N_46175,N_46176,N_46177,N_46178,N_46179,N_46180,N_46181,N_46182,N_46183,N_46184,N_46185,N_46186,N_46187,N_46188,N_46189,N_46190,N_46191,N_46192,N_46193,N_46194,N_46195,N_46196,N_46197,N_46198,N_46199,N_46200,N_46201,N_46202,N_46203,N_46204,N_46205,N_46206,N_46207,N_46208,N_46209,N_46210,N_46211,N_46212,N_46213,N_46214,N_46215,N_46216,N_46217,N_46218,N_46219,N_46220,N_46221,N_46222,N_46223,N_46224,N_46225,N_46226,N_46227,N_46228,N_46229,N_46230,N_46231,N_46232,N_46233,N_46234,N_46235,N_46236,N_46237,N_46238,N_46239,N_46240,N_46241,N_46242,N_46243,N_46244,N_46245,N_46246,N_46247,N_46248,N_46249,N_46250,N_46251,N_46252,N_46253,N_46254,N_46255,N_46256,N_46257,N_46258,N_46259,N_46260,N_46261,N_46262,N_46263,N_46264,N_46265,N_46266,N_46267,N_46268,N_46269,N_46270,N_46271,N_46272,N_46273,N_46274,N_46275,N_46276,N_46277,N_46278,N_46279,N_46280,N_46281,N_46282,N_46283,N_46284,N_46285,N_46286,N_46287,N_46288,N_46289,N_46290,N_46291,N_46292,N_46293,N_46294,N_46295,N_46296,N_46297,N_46298,N_46299,N_46300,N_46301,N_46302,N_46303,N_46304,N_46305,N_46306,N_46307,N_46308,N_46309,N_46310,N_46311,N_46312,N_46313,N_46314,N_46315,N_46316,N_46317,N_46318,N_46319,N_46320,N_46321,N_46322,N_46323,N_46324,N_46325,N_46326,N_46327,N_46328,N_46329,N_46330,N_46331,N_46332,N_46333,N_46334,N_46335,N_46336,N_46337,N_46338,N_46339,N_46340,N_46341,N_46342,N_46343,N_46344,N_46345,N_46346,N_46347,N_46348,N_46349,N_46350,N_46351,N_46352,N_46353,N_46354,N_46355,N_46356,N_46357,N_46358,N_46359,N_46360,N_46361,N_46362,N_46363,N_46364,N_46365,N_46366,N_46367,N_46368,N_46369,N_46370,N_46371,N_46372,N_46373,N_46374,N_46375,N_46376,N_46377,N_46378,N_46379,N_46380,N_46381,N_46382,N_46383,N_46384,N_46385,N_46386,N_46387,N_46388,N_46389,N_46390,N_46391,N_46392,N_46393,N_46394,N_46395,N_46396,N_46397,N_46398,N_46399,N_46400,N_46401,N_46402,N_46403,N_46404,N_46405,N_46406,N_46407,N_46408,N_46409,N_46410,N_46411,N_46412,N_46413,N_46414,N_46415,N_46416,N_46417,N_46418,N_46419,N_46420,N_46421,N_46422,N_46423,N_46424,N_46425,N_46426,N_46427,N_46428,N_46429,N_46430,N_46431,N_46432,N_46433,N_46434,N_46435,N_46436,N_46437,N_46438,N_46439,N_46440,N_46441,N_46442,N_46443,N_46444,N_46445,N_46446,N_46447,N_46448,N_46449,N_46450,N_46451,N_46452,N_46453,N_46454,N_46455,N_46456,N_46457,N_46458,N_46459,N_46460,N_46461,N_46462,N_46463,N_46464,N_46465,N_46466,N_46467,N_46468,N_46469,N_46470,N_46471,N_46472,N_46473,N_46474,N_46475,N_46476,N_46477,N_46478,N_46479,N_46480,N_46481,N_46482,N_46483,N_46484,N_46485,N_46486,N_46487,N_46488,N_46489,N_46490,N_46491,N_46492,N_46493,N_46494,N_46495,N_46496,N_46497,N_46498,N_46499,N_46500,N_46501,N_46502,N_46503,N_46504,N_46505,N_46506,N_46507,N_46508,N_46509,N_46510,N_46511,N_46512,N_46513,N_46514,N_46515,N_46516,N_46517,N_46518,N_46519,N_46520,N_46521,N_46522,N_46523,N_46524,N_46525,N_46526,N_46527,N_46528,N_46529,N_46530,N_46531,N_46532,N_46533,N_46534,N_46535,N_46536,N_46537,N_46538,N_46539,N_46540,N_46541,N_46542,N_46543,N_46544,N_46545,N_46546,N_46547,N_46548,N_46549,N_46550,N_46551,N_46552,N_46553,N_46554,N_46555,N_46556,N_46557,N_46558,N_46559,N_46560,N_46561,N_46562,N_46563,N_46564,N_46565,N_46566,N_46567,N_46568,N_46569,N_46570,N_46571,N_46572,N_46573,N_46574,N_46575,N_46576,N_46577,N_46578,N_46579,N_46580,N_46581,N_46582,N_46583,N_46584,N_46585,N_46586,N_46587,N_46588,N_46589,N_46590,N_46591,N_46592,N_46593,N_46594,N_46595,N_46596,N_46597,N_46598,N_46599,N_46600,N_46601,N_46602,N_46603,N_46604,N_46605,N_46606,N_46607,N_46608,N_46609,N_46610,N_46611,N_46612,N_46613,N_46614,N_46615,N_46616,N_46617,N_46618,N_46619,N_46620,N_46621,N_46622,N_46623,N_46624,N_46625,N_46626,N_46627,N_46628,N_46629,N_46630,N_46631,N_46632,N_46633,N_46634,N_46635,N_46636,N_46637,N_46638,N_46639,N_46640,N_46641,N_46642,N_46643,N_46644,N_46645,N_46646,N_46647,N_46648,N_46649,N_46650,N_46651,N_46652,N_46653,N_46654,N_46655,N_46656,N_46657,N_46658,N_46659,N_46660,N_46661,N_46662,N_46663,N_46664,N_46665,N_46666,N_46667,N_46668,N_46669,N_46670,N_46671,N_46672,N_46673,N_46674,N_46675,N_46676,N_46677,N_46678,N_46679,N_46680,N_46681,N_46682,N_46683,N_46684,N_46685,N_46686,N_46687,N_46688,N_46689,N_46690,N_46691,N_46692,N_46693,N_46694,N_46695,N_46696,N_46697,N_46698,N_46699,N_46700,N_46701,N_46702,N_46703,N_46704,N_46705,N_46706,N_46707,N_46708,N_46709,N_46710,N_46711,N_46712,N_46713,N_46714,N_46715,N_46716,N_46717,N_46718,N_46719,N_46720,N_46721,N_46722,N_46723,N_46724,N_46725,N_46726,N_46727,N_46728,N_46729,N_46730,N_46731,N_46732,N_46733,N_46734,N_46735,N_46736,N_46737,N_46738,N_46739,N_46740,N_46741,N_46742,N_46743,N_46744,N_46745,N_46746,N_46747,N_46748,N_46749,N_46750,N_46751,N_46752,N_46753,N_46754,N_46755,N_46756,N_46757,N_46758,N_46759,N_46760,N_46761,N_46762,N_46763,N_46764,N_46765,N_46766,N_46767,N_46768,N_46769,N_46770,N_46771,N_46772,N_46773,N_46774,N_46775,N_46776,N_46777,N_46778,N_46779,N_46780,N_46781,N_46782,N_46783,N_46784,N_46785,N_46786,N_46787,N_46788,N_46789,N_46790,N_46791,N_46792,N_46793,N_46794,N_46795,N_46796,N_46797,N_46798,N_46799,N_46800,N_46801,N_46802,N_46803,N_46804,N_46805,N_46806,N_46807,N_46808,N_46809,N_46810,N_46811,N_46812,N_46813,N_46814,N_46815,N_46816,N_46817,N_46818,N_46819,N_46820,N_46821,N_46822,N_46823,N_46824,N_46825,N_46826,N_46827,N_46828,N_46829,N_46830,N_46831,N_46832,N_46833,N_46834,N_46835,N_46836,N_46837,N_46838,N_46839,N_46840,N_46841,N_46842,N_46843,N_46844,N_46845,N_46846,N_46847,N_46848,N_46849,N_46850,N_46851,N_46852,N_46853,N_46854,N_46855,N_46856,N_46857,N_46858,N_46859,N_46860,N_46861,N_46862,N_46863,N_46864,N_46865,N_46866,N_46867,N_46868,N_46869,N_46870,N_46871,N_46872,N_46873,N_46874,N_46875,N_46876,N_46877,N_46878,N_46879,N_46880,N_46881,N_46882,N_46883,N_46884,N_46885,N_46886,N_46887,N_46888,N_46889,N_46890,N_46891,N_46892,N_46893,N_46894,N_46895,N_46896,N_46897,N_46898,N_46899,N_46900,N_46901,N_46902,N_46903,N_46904,N_46905,N_46906,N_46907,N_46908,N_46909,N_46910,N_46911,N_46912,N_46913,N_46914,N_46915,N_46916,N_46917,N_46918,N_46919,N_46920,N_46921,N_46922,N_46923,N_46924,N_46925,N_46926,N_46927,N_46928,N_46929,N_46930,N_46931,N_46932,N_46933,N_46934,N_46935,N_46936,N_46937,N_46938,N_46939,N_46940,N_46941,N_46942,N_46943,N_46944,N_46945,N_46946,N_46947,N_46948,N_46949,N_46950,N_46951,N_46952,N_46953,N_46954,N_46955,N_46956,N_46957,N_46958,N_46959,N_46960,N_46961,N_46962,N_46963,N_46964,N_46965,N_46966,N_46967,N_46968,N_46969,N_46970,N_46971,N_46972,N_46973,N_46974,N_46975,N_46976,N_46977,N_46978,N_46979,N_46980,N_46981,N_46982,N_46983,N_46984,N_46985,N_46986,N_46987,N_46988,N_46989,N_46990,N_46991,N_46992,N_46993,N_46994,N_46995,N_46996,N_46997,N_46998,N_46999,N_47000,N_47001,N_47002,N_47003,N_47004,N_47005,N_47006,N_47007,N_47008,N_47009,N_47010,N_47011,N_47012,N_47013,N_47014,N_47015,N_47016,N_47017,N_47018,N_47019,N_47020,N_47021,N_47022,N_47023,N_47024,N_47025,N_47026,N_47027,N_47028,N_47029,N_47030,N_47031,N_47032,N_47033,N_47034,N_47035,N_47036,N_47037,N_47038,N_47039,N_47040,N_47041,N_47042,N_47043,N_47044,N_47045,N_47046,N_47047,N_47048,N_47049,N_47050,N_47051,N_47052,N_47053,N_47054,N_47055,N_47056,N_47057,N_47058,N_47059,N_47060,N_47061,N_47062,N_47063,N_47064,N_47065,N_47066,N_47067,N_47068,N_47069,N_47070,N_47071,N_47072,N_47073,N_47074,N_47075,N_47076,N_47077,N_47078,N_47079,N_47080,N_47081,N_47082,N_47083,N_47084,N_47085,N_47086,N_47087,N_47088,N_47089,N_47090,N_47091,N_47092,N_47093,N_47094,N_47095,N_47096,N_47097,N_47098,N_47099,N_47100,N_47101,N_47102,N_47103,N_47104,N_47105,N_47106,N_47107,N_47108,N_47109,N_47110,N_47111,N_47112,N_47113,N_47114,N_47115,N_47116,N_47117,N_47118,N_47119,N_47120,N_47121,N_47122,N_47123,N_47124,N_47125,N_47126,N_47127,N_47128,N_47129,N_47130,N_47131,N_47132,N_47133,N_47134,N_47135,N_47136,N_47137,N_47138,N_47139,N_47140,N_47141,N_47142,N_47143,N_47144,N_47145,N_47146,N_47147,N_47148,N_47149,N_47150,N_47151,N_47152,N_47153,N_47154,N_47155,N_47156,N_47157,N_47158,N_47159,N_47160,N_47161,N_47162,N_47163,N_47164,N_47165,N_47166,N_47167,N_47168,N_47169,N_47170,N_47171,N_47172,N_47173,N_47174,N_47175,N_47176,N_47177,N_47178,N_47179,N_47180,N_47181,N_47182,N_47183,N_47184,N_47185,N_47186,N_47187,N_47188,N_47189,N_47190,N_47191,N_47192,N_47193,N_47194,N_47195,N_47196,N_47197,N_47198,N_47199,N_47200,N_47201,N_47202,N_47203,N_47204,N_47205,N_47206,N_47207,N_47208,N_47209,N_47210,N_47211,N_47212,N_47213,N_47214,N_47215,N_47216,N_47217,N_47218,N_47219,N_47220,N_47221,N_47222,N_47223,N_47224,N_47225,N_47226,N_47227,N_47228,N_47229,N_47230,N_47231,N_47232,N_47233,N_47234,N_47235,N_47236,N_47237,N_47238,N_47239,N_47240,N_47241,N_47242,N_47243,N_47244,N_47245,N_47246,N_47247,N_47248,N_47249,N_47250,N_47251,N_47252,N_47253,N_47254,N_47255,N_47256,N_47257,N_47258,N_47259,N_47260,N_47261,N_47262,N_47263,N_47264,N_47265,N_47266,N_47267,N_47268,N_47269,N_47270,N_47271,N_47272,N_47273,N_47274,N_47275,N_47276,N_47277,N_47278,N_47279,N_47280,N_47281,N_47282,N_47283,N_47284,N_47285,N_47286,N_47287,N_47288,N_47289,N_47290,N_47291,N_47292,N_47293,N_47294,N_47295,N_47296,N_47297,N_47298,N_47299,N_47300,N_47301,N_47302,N_47303,N_47304,N_47305,N_47306,N_47307,N_47308,N_47309,N_47310,N_47311,N_47312,N_47313,N_47314,N_47315,N_47316,N_47317,N_47318,N_47319,N_47320,N_47321,N_47322,N_47323,N_47324,N_47325,N_47326,N_47327,N_47328,N_47329,N_47330,N_47331,N_47332,N_47333,N_47334,N_47335,N_47336,N_47337,N_47338,N_47339,N_47340,N_47341,N_47342,N_47343,N_47344,N_47345,N_47346,N_47347,N_47348,N_47349,N_47350,N_47351,N_47352,N_47353,N_47354,N_47355,N_47356,N_47357,N_47358,N_47359,N_47360,N_47361,N_47362,N_47363,N_47364,N_47365,N_47366,N_47367,N_47368,N_47369,N_47370,N_47371,N_47372,N_47373,N_47374,N_47375,N_47376,N_47377,N_47378,N_47379,N_47380,N_47381,N_47382,N_47383,N_47384,N_47385,N_47386,N_47387,N_47388,N_47389,N_47390,N_47391,N_47392,N_47393,N_47394,N_47395,N_47396,N_47397,N_47398,N_47399,N_47400,N_47401,N_47402,N_47403,N_47404,N_47405,N_47406,N_47407,N_47408,N_47409,N_47410,N_47411,N_47412,N_47413,N_47414,N_47415,N_47416,N_47417,N_47418,N_47419,N_47420,N_47421,N_47422,N_47423,N_47424,N_47425,N_47426,N_47427,N_47428,N_47429,N_47430,N_47431,N_47432,N_47433,N_47434,N_47435,N_47436,N_47437,N_47438,N_47439,N_47440,N_47441,N_47442,N_47443,N_47444,N_47445,N_47446,N_47447,N_47448,N_47449,N_47450,N_47451,N_47452,N_47453,N_47454,N_47455,N_47456,N_47457,N_47458,N_47459,N_47460,N_47461,N_47462,N_47463,N_47464,N_47465,N_47466,N_47467,N_47468,N_47469,N_47470,N_47471,N_47472,N_47473,N_47474,N_47475,N_47476,N_47477,N_47478,N_47479,N_47480,N_47481,N_47482,N_47483,N_47484,N_47485,N_47486,N_47487,N_47488,N_47489,N_47490,N_47491,N_47492,N_47493,N_47494,N_47495,N_47496,N_47497,N_47498,N_47499,N_47500,N_47501,N_47502,N_47503,N_47504,N_47505,N_47506,N_47507,N_47508,N_47509,N_47510,N_47511,N_47512,N_47513,N_47514,N_47515,N_47516,N_47517,N_47518,N_47519,N_47520,N_47521,N_47522,N_47523,N_47524,N_47525,N_47526,N_47527,N_47528,N_47529,N_47530,N_47531,N_47532,N_47533,N_47534,N_47535,N_47536,N_47537,N_47538,N_47539,N_47540,N_47541,N_47542,N_47543,N_47544,N_47545,N_47546,N_47547,N_47548,N_47549,N_47550,N_47551,N_47552,N_47553,N_47554,N_47555,N_47556,N_47557,N_47558,N_47559,N_47560,N_47561,N_47562,N_47563,N_47564,N_47565,N_47566,N_47567,N_47568,N_47569,N_47570,N_47571,N_47572,N_47573,N_47574,N_47575,N_47576,N_47577,N_47578,N_47579,N_47580,N_47581,N_47582,N_47583,N_47584,N_47585,N_47586,N_47587,N_47588,N_47589,N_47590,N_47591,N_47592,N_47593,N_47594,N_47595,N_47596,N_47597,N_47598,N_47599,N_47600,N_47601,N_47602,N_47603,N_47604,N_47605,N_47606,N_47607,N_47608,N_47609,N_47610,N_47611,N_47612,N_47613,N_47614,N_47615,N_47616,N_47617,N_47618,N_47619,N_47620,N_47621,N_47622,N_47623,N_47624,N_47625,N_47626,N_47627,N_47628,N_47629,N_47630,N_47631,N_47632,N_47633,N_47634,N_47635,N_47636,N_47637,N_47638,N_47639,N_47640,N_47641,N_47642,N_47643,N_47644,N_47645,N_47646,N_47647,N_47648,N_47649,N_47650,N_47651,N_47652,N_47653,N_47654,N_47655,N_47656,N_47657,N_47658,N_47659,N_47660,N_47661,N_47662,N_47663,N_47664,N_47665,N_47666,N_47667,N_47668,N_47669,N_47670,N_47671,N_47672,N_47673,N_47674,N_47675,N_47676,N_47677,N_47678,N_47679,N_47680,N_47681,N_47682,N_47683,N_47684,N_47685,N_47686,N_47687,N_47688,N_47689,N_47690,N_47691,N_47692,N_47693,N_47694,N_47695,N_47696,N_47697,N_47698,N_47699,N_47700,N_47701,N_47702,N_47703,N_47704,N_47705,N_47706,N_47707,N_47708,N_47709,N_47710,N_47711,N_47712,N_47713,N_47714,N_47715,N_47716,N_47717,N_47718,N_47719,N_47720,N_47721,N_47722,N_47723,N_47724,N_47725,N_47726,N_47727,N_47728,N_47729,N_47730,N_47731,N_47732,N_47733,N_47734,N_47735,N_47736,N_47737,N_47738,N_47739,N_47740,N_47741,N_47742,N_47743,N_47744,N_47745,N_47746,N_47747,N_47748,N_47749,N_47750,N_47751,N_47752,N_47753,N_47754,N_47755,N_47756,N_47757,N_47758,N_47759,N_47760,N_47761,N_47762,N_47763,N_47764,N_47765,N_47766,N_47767,N_47768,N_47769,N_47770,N_47771,N_47772,N_47773,N_47774,N_47775,N_47776,N_47777,N_47778,N_47779,N_47780,N_47781,N_47782,N_47783,N_47784,N_47785,N_47786,N_47787,N_47788,N_47789,N_47790,N_47791,N_47792,N_47793,N_47794,N_47795,N_47796,N_47797,N_47798,N_47799,N_47800,N_47801,N_47802,N_47803,N_47804,N_47805,N_47806,N_47807,N_47808,N_47809,N_47810,N_47811,N_47812,N_47813,N_47814,N_47815,N_47816,N_47817,N_47818,N_47819,N_47820,N_47821,N_47822,N_47823,N_47824,N_47825,N_47826,N_47827,N_47828,N_47829,N_47830,N_47831,N_47832,N_47833,N_47834,N_47835,N_47836,N_47837,N_47838,N_47839,N_47840,N_47841,N_47842,N_47843,N_47844,N_47845,N_47846,N_47847,N_47848,N_47849,N_47850,N_47851,N_47852,N_47853,N_47854,N_47855,N_47856,N_47857,N_47858,N_47859,N_47860,N_47861,N_47862,N_47863,N_47864,N_47865,N_47866,N_47867,N_47868,N_47869,N_47870,N_47871,N_47872,N_47873,N_47874,N_47875,N_47876,N_47877,N_47878,N_47879,N_47880,N_47881,N_47882,N_47883,N_47884,N_47885,N_47886,N_47887,N_47888,N_47889,N_47890,N_47891,N_47892,N_47893,N_47894,N_47895,N_47896,N_47897,N_47898,N_47899,N_47900,N_47901,N_47902,N_47903,N_47904,N_47905,N_47906,N_47907,N_47908,N_47909,N_47910,N_47911,N_47912,N_47913,N_47914,N_47915,N_47916,N_47917,N_47918,N_47919,N_47920,N_47921,N_47922,N_47923,N_47924,N_47925,N_47926,N_47927,N_47928,N_47929,N_47930,N_47931,N_47932,N_47933,N_47934,N_47935,N_47936,N_47937,N_47938,N_47939,N_47940,N_47941,N_47942,N_47943,N_47944,N_47945,N_47946,N_47947,N_47948,N_47949,N_47950,N_47951,N_47952,N_47953,N_47954,N_47955,N_47956,N_47957,N_47958,N_47959,N_47960,N_47961,N_47962,N_47963,N_47964,N_47965,N_47966,N_47967,N_47968,N_47969,N_47970,N_47971,N_47972,N_47973,N_47974,N_47975,N_47976,N_47977,N_47978,N_47979,N_47980,N_47981,N_47982,N_47983,N_47984,N_47985,N_47986,N_47987,N_47988,N_47989,N_47990,N_47991,N_47992,N_47993,N_47994,N_47995,N_47996,N_47997,N_47998,N_47999,N_48000,N_48001,N_48002,N_48003,N_48004,N_48005,N_48006,N_48007,N_48008,N_48009,N_48010,N_48011,N_48012,N_48013,N_48014,N_48015,N_48016,N_48017,N_48018,N_48019,N_48020,N_48021,N_48022,N_48023,N_48024,N_48025,N_48026,N_48027,N_48028,N_48029,N_48030,N_48031,N_48032,N_48033,N_48034,N_48035,N_48036,N_48037,N_48038,N_48039,N_48040,N_48041,N_48042,N_48043,N_48044,N_48045,N_48046,N_48047,N_48048,N_48049,N_48050,N_48051,N_48052,N_48053,N_48054,N_48055,N_48056,N_48057,N_48058,N_48059,N_48060,N_48061,N_48062,N_48063,N_48064,N_48065,N_48066,N_48067,N_48068,N_48069,N_48070,N_48071,N_48072,N_48073,N_48074,N_48075,N_48076,N_48077,N_48078,N_48079,N_48080,N_48081,N_48082,N_48083,N_48084,N_48085,N_48086,N_48087,N_48088,N_48089,N_48090,N_48091,N_48092,N_48093,N_48094,N_48095,N_48096,N_48097,N_48098,N_48099,N_48100,N_48101,N_48102,N_48103,N_48104,N_48105,N_48106,N_48107,N_48108,N_48109,N_48110,N_48111,N_48112,N_48113,N_48114,N_48115,N_48116,N_48117,N_48118,N_48119,N_48120,N_48121,N_48122,N_48123,N_48124,N_48125,N_48126,N_48127,N_48128,N_48129,N_48130,N_48131,N_48132,N_48133,N_48134,N_48135,N_48136,N_48137,N_48138,N_48139,N_48140,N_48141,N_48142,N_48143,N_48144,N_48145,N_48146,N_48147,N_48148,N_48149,N_48150,N_48151,N_48152,N_48153,N_48154,N_48155,N_48156,N_48157,N_48158,N_48159,N_48160,N_48161,N_48162,N_48163,N_48164,N_48165,N_48166,N_48167,N_48168,N_48169,N_48170,N_48171,N_48172,N_48173,N_48174,N_48175,N_48176,N_48177,N_48178,N_48179,N_48180,N_48181,N_48182,N_48183,N_48184,N_48185,N_48186,N_48187,N_48188,N_48189,N_48190,N_48191,N_48192,N_48193,N_48194,N_48195,N_48196,N_48197,N_48198,N_48199,N_48200,N_48201,N_48202,N_48203,N_48204,N_48205,N_48206,N_48207,N_48208,N_48209,N_48210,N_48211,N_48212,N_48213,N_48214,N_48215,N_48216,N_48217,N_48218,N_48219,N_48220,N_48221,N_48222,N_48223,N_48224,N_48225,N_48226,N_48227,N_48228,N_48229,N_48230,N_48231,N_48232,N_48233,N_48234,N_48235,N_48236,N_48237,N_48238,N_48239,N_48240,N_48241,N_48242,N_48243,N_48244,N_48245,N_48246,N_48247,N_48248,N_48249,N_48250,N_48251,N_48252,N_48253,N_48254,N_48255,N_48256,N_48257,N_48258,N_48259,N_48260,N_48261,N_48262,N_48263,N_48264,N_48265,N_48266,N_48267,N_48268,N_48269,N_48270,N_48271,N_48272,N_48273,N_48274,N_48275,N_48276,N_48277,N_48278,N_48279,N_48280,N_48281,N_48282,N_48283,N_48284,N_48285,N_48286,N_48287,N_48288,N_48289,N_48290,N_48291,N_48292,N_48293,N_48294,N_48295,N_48296,N_48297,N_48298,N_48299,N_48300,N_48301,N_48302,N_48303,N_48304,N_48305,N_48306,N_48307,N_48308,N_48309,N_48310,N_48311,N_48312,N_48313,N_48314,N_48315,N_48316,N_48317,N_48318,N_48319,N_48320,N_48321,N_48322,N_48323,N_48324,N_48325,N_48326,N_48327,N_48328,N_48329,N_48330,N_48331,N_48332,N_48333,N_48334,N_48335,N_48336,N_48337,N_48338,N_48339,N_48340,N_48341,N_48342,N_48343,N_48344,N_48345,N_48346,N_48347,N_48348,N_48349,N_48350,N_48351,N_48352,N_48353,N_48354,N_48355,N_48356,N_48357,N_48358,N_48359,N_48360,N_48361,N_48362,N_48363,N_48364,N_48365,N_48366,N_48367,N_48368,N_48369,N_48370,N_48371,N_48372,N_48373,N_48374,N_48375,N_48376,N_48377,N_48378,N_48379,N_48380,N_48381,N_48382,N_48383,N_48384,N_48385,N_48386,N_48387,N_48388,N_48389,N_48390,N_48391,N_48392,N_48393,N_48394,N_48395,N_48396,N_48397,N_48398,N_48399,N_48400,N_48401,N_48402,N_48403,N_48404,N_48405,N_48406,N_48407,N_48408,N_48409,N_48410,N_48411,N_48412,N_48413,N_48414,N_48415,N_48416,N_48417,N_48418,N_48419,N_48420,N_48421,N_48422,N_48423,N_48424,N_48425,N_48426,N_48427,N_48428,N_48429,N_48430,N_48431,N_48432,N_48433,N_48434,N_48435,N_48436,N_48437,N_48438,N_48439,N_48440,N_48441,N_48442,N_48443,N_48444,N_48445,N_48446,N_48447,N_48448,N_48449,N_48450,N_48451,N_48452,N_48453,N_48454,N_48455,N_48456,N_48457,N_48458,N_48459,N_48460,N_48461,N_48462,N_48463,N_48464,N_48465,N_48466,N_48467,N_48468,N_48469,N_48470,N_48471,N_48472,N_48473,N_48474,N_48475,N_48476,N_48477,N_48478,N_48479,N_48480,N_48481,N_48482,N_48483,N_48484,N_48485,N_48486,N_48487,N_48488,N_48489,N_48490,N_48491,N_48492,N_48493,N_48494,N_48495,N_48496,N_48497,N_48498,N_48499,N_48500,N_48501,N_48502,N_48503,N_48504,N_48505,N_48506,N_48507,N_48508,N_48509,N_48510,N_48511,N_48512,N_48513,N_48514,N_48515,N_48516,N_48517,N_48518,N_48519,N_48520,N_48521,N_48522,N_48523,N_48524,N_48525,N_48526,N_48527,N_48528,N_48529,N_48530,N_48531,N_48532,N_48533,N_48534,N_48535,N_48536,N_48537,N_48538,N_48539,N_48540,N_48541,N_48542,N_48543,N_48544,N_48545,N_48546,N_48547,N_48548,N_48549,N_48550,N_48551,N_48552,N_48553,N_48554,N_48555,N_48556,N_48557,N_48558,N_48559,N_48560,N_48561,N_48562,N_48563,N_48564,N_48565,N_48566,N_48567,N_48568,N_48569,N_48570,N_48571,N_48572,N_48573,N_48574,N_48575,N_48576,N_48577,N_48578,N_48579,N_48580,N_48581,N_48582,N_48583,N_48584,N_48585,N_48586,N_48587,N_48588,N_48589,N_48590,N_48591,N_48592,N_48593,N_48594,N_48595,N_48596,N_48597,N_48598,N_48599,N_48600,N_48601,N_48602,N_48603,N_48604,N_48605,N_48606,N_48607,N_48608,N_48609,N_48610,N_48611,N_48612,N_48613,N_48614,N_48615,N_48616,N_48617,N_48618,N_48619,N_48620,N_48621,N_48622,N_48623,N_48624,N_48625,N_48626,N_48627,N_48628,N_48629,N_48630,N_48631,N_48632,N_48633,N_48634,N_48635,N_48636,N_48637,N_48638,N_48639,N_48640,N_48641,N_48642,N_48643,N_48644,N_48645,N_48646,N_48647,N_48648,N_48649,N_48650,N_48651,N_48652,N_48653,N_48654,N_48655,N_48656,N_48657,N_48658,N_48659,N_48660,N_48661,N_48662,N_48663,N_48664,N_48665,N_48666,N_48667,N_48668,N_48669,N_48670,N_48671,N_48672,N_48673,N_48674,N_48675,N_48676,N_48677,N_48678,N_48679,N_48680,N_48681,N_48682,N_48683,N_48684,N_48685,N_48686,N_48687,N_48688,N_48689,N_48690,N_48691,N_48692,N_48693,N_48694,N_48695,N_48696,N_48697,N_48698,N_48699,N_48700,N_48701,N_48702,N_48703,N_48704,N_48705,N_48706,N_48707,N_48708,N_48709,N_48710,N_48711,N_48712,N_48713,N_48714,N_48715,N_48716,N_48717,N_48718,N_48719,N_48720,N_48721,N_48722,N_48723,N_48724,N_48725,N_48726,N_48727,N_48728,N_48729,N_48730,N_48731,N_48732,N_48733,N_48734,N_48735,N_48736,N_48737,N_48738,N_48739,N_48740,N_48741,N_48742,N_48743,N_48744,N_48745,N_48746,N_48747,N_48748,N_48749,N_48750,N_48751,N_48752,N_48753,N_48754,N_48755,N_48756,N_48757,N_48758,N_48759,N_48760,N_48761,N_48762,N_48763,N_48764,N_48765,N_48766,N_48767,N_48768,N_48769,N_48770,N_48771,N_48772,N_48773,N_48774,N_48775,N_48776,N_48777,N_48778,N_48779,N_48780,N_48781,N_48782,N_48783,N_48784,N_48785,N_48786,N_48787,N_48788,N_48789,N_48790,N_48791,N_48792,N_48793,N_48794,N_48795,N_48796,N_48797,N_48798,N_48799,N_48800,N_48801,N_48802,N_48803,N_48804,N_48805,N_48806,N_48807,N_48808,N_48809,N_48810,N_48811,N_48812,N_48813,N_48814,N_48815,N_48816,N_48817,N_48818,N_48819,N_48820,N_48821,N_48822,N_48823,N_48824,N_48825,N_48826,N_48827,N_48828,N_48829,N_48830,N_48831,N_48832,N_48833,N_48834,N_48835,N_48836,N_48837,N_48838,N_48839,N_48840,N_48841,N_48842,N_48843,N_48844,N_48845,N_48846,N_48847,N_48848,N_48849,N_48850,N_48851,N_48852,N_48853,N_48854,N_48855,N_48856,N_48857,N_48858,N_48859,N_48860,N_48861,N_48862,N_48863,N_48864,N_48865,N_48866,N_48867,N_48868,N_48869,N_48870,N_48871,N_48872,N_48873,N_48874,N_48875,N_48876,N_48877,N_48878,N_48879,N_48880,N_48881,N_48882,N_48883,N_48884,N_48885,N_48886,N_48887,N_48888,N_48889,N_48890,N_48891,N_48892,N_48893,N_48894,N_48895,N_48896,N_48897,N_48898,N_48899,N_48900,N_48901,N_48902,N_48903,N_48904,N_48905,N_48906,N_48907,N_48908,N_48909,N_48910,N_48911,N_48912,N_48913,N_48914,N_48915,N_48916,N_48917,N_48918,N_48919,N_48920,N_48921,N_48922,N_48923,N_48924,N_48925,N_48926,N_48927,N_48928,N_48929,N_48930,N_48931,N_48932,N_48933,N_48934,N_48935,N_48936,N_48937,N_48938,N_48939,N_48940,N_48941,N_48942,N_48943,N_48944,N_48945,N_48946,N_48947,N_48948,N_48949,N_48950,N_48951,N_48952,N_48953,N_48954,N_48955,N_48956,N_48957,N_48958,N_48959,N_48960,N_48961,N_48962,N_48963,N_48964,N_48965,N_48966,N_48967,N_48968,N_48969,N_48970,N_48971,N_48972,N_48973,N_48974,N_48975,N_48976,N_48977,N_48978,N_48979,N_48980,N_48981,N_48982,N_48983,N_48984,N_48985,N_48986,N_48987,N_48988,N_48989,N_48990,N_48991,N_48992,N_48993,N_48994,N_48995,N_48996,N_48997,N_48998,N_48999,N_49000,N_49001,N_49002,N_49003,N_49004,N_49005,N_49006,N_49007,N_49008,N_49009,N_49010,N_49011,N_49012,N_49013,N_49014,N_49015,N_49016,N_49017,N_49018,N_49019,N_49020,N_49021,N_49022,N_49023,N_49024,N_49025,N_49026,N_49027,N_49028,N_49029,N_49030,N_49031,N_49032,N_49033,N_49034,N_49035,N_49036,N_49037,N_49038,N_49039,N_49040,N_49041,N_49042,N_49043,N_49044,N_49045,N_49046,N_49047,N_49048,N_49049,N_49050,N_49051,N_49052,N_49053,N_49054,N_49055,N_49056,N_49057,N_49058,N_49059,N_49060,N_49061,N_49062,N_49063,N_49064,N_49065,N_49066,N_49067,N_49068,N_49069,N_49070,N_49071,N_49072,N_49073,N_49074,N_49075,N_49076,N_49077,N_49078,N_49079,N_49080,N_49081,N_49082,N_49083,N_49084,N_49085,N_49086,N_49087,N_49088,N_49089,N_49090,N_49091,N_49092,N_49093,N_49094,N_49095,N_49096,N_49097,N_49098,N_49099,N_49100,N_49101,N_49102,N_49103,N_49104,N_49105,N_49106,N_49107,N_49108,N_49109,N_49110,N_49111,N_49112,N_49113,N_49114,N_49115,N_49116,N_49117,N_49118,N_49119,N_49120,N_49121,N_49122,N_49123,N_49124,N_49125,N_49126,N_49127,N_49128,N_49129,N_49130,N_49131,N_49132,N_49133,N_49134,N_49135,N_49136,N_49137,N_49138,N_49139,N_49140,N_49141,N_49142,N_49143,N_49144,N_49145,N_49146,N_49147,N_49148,N_49149,N_49150,N_49151,N_49152,N_49153,N_49154,N_49155,N_49156,N_49157,N_49158,N_49159,N_49160,N_49161,N_49162,N_49163,N_49164,N_49165,N_49166,N_49167,N_49168,N_49169,N_49170,N_49171,N_49172,N_49173,N_49174,N_49175,N_49176,N_49177,N_49178,N_49179,N_49180,N_49181,N_49182,N_49183,N_49184,N_49185,N_49186,N_49187,N_49188,N_49189,N_49190,N_49191,N_49192,N_49193,N_49194,N_49195,N_49196,N_49197,N_49198,N_49199,N_49200,N_49201,N_49202,N_49203,N_49204,N_49205,N_49206,N_49207,N_49208,N_49209,N_49210,N_49211,N_49212,N_49213,N_49214,N_49215,N_49216,N_49217,N_49218,N_49219,N_49220,N_49221,N_49222,N_49223,N_49224,N_49225,N_49226,N_49227,N_49228,N_49229,N_49230,N_49231,N_49232,N_49233,N_49234,N_49235,N_49236,N_49237,N_49238,N_49239,N_49240,N_49241,N_49242,N_49243,N_49244,N_49245,N_49246,N_49247,N_49248,N_49249,N_49250,N_49251,N_49252,N_49253,N_49254,N_49255,N_49256,N_49257,N_49258,N_49259,N_49260,N_49261,N_49262,N_49263,N_49264,N_49265,N_49266,N_49267,N_49268,N_49269,N_49270,N_49271,N_49272,N_49273,N_49274,N_49275,N_49276,N_49277,N_49278,N_49279,N_49280,N_49281,N_49282,N_49283,N_49284,N_49285,N_49286,N_49287,N_49288,N_49289,N_49290,N_49291,N_49292,N_49293,N_49294,N_49295,N_49296,N_49297,N_49298,N_49299,N_49300,N_49301,N_49302,N_49303,N_49304,N_49305,N_49306,N_49307,N_49308,N_49309,N_49310,N_49311,N_49312,N_49313,N_49314,N_49315,N_49316,N_49317,N_49318,N_49319,N_49320,N_49321,N_49322,N_49323,N_49324,N_49325,N_49326,N_49327,N_49328,N_49329,N_49330,N_49331,N_49332,N_49333,N_49334,N_49335,N_49336,N_49337,N_49338,N_49339,N_49340,N_49341,N_49342,N_49343,N_49344,N_49345,N_49346,N_49347,N_49348,N_49349,N_49350,N_49351,N_49352,N_49353,N_49354,N_49355,N_49356,N_49357,N_49358,N_49359,N_49360,N_49361,N_49362,N_49363,N_49364,N_49365,N_49366,N_49367,N_49368,N_49369,N_49370,N_49371,N_49372,N_49373,N_49374,N_49375,N_49376,N_49377,N_49378,N_49379,N_49380,N_49381,N_49382,N_49383,N_49384,N_49385,N_49386,N_49387,N_49388,N_49389,N_49390,N_49391,N_49392,N_49393,N_49394,N_49395,N_49396,N_49397,N_49398,N_49399,N_49400,N_49401,N_49402,N_49403,N_49404,N_49405,N_49406,N_49407,N_49408,N_49409,N_49410,N_49411,N_49412,N_49413,N_49414,N_49415,N_49416,N_49417,N_49418,N_49419,N_49420,N_49421,N_49422,N_49423,N_49424,N_49425,N_49426,N_49427,N_49428,N_49429,N_49430,N_49431,N_49432,N_49433,N_49434,N_49435,N_49436,N_49437,N_49438,N_49439,N_49440,N_49441,N_49442,N_49443,N_49444,N_49445,N_49446,N_49447,N_49448,N_49449,N_49450,N_49451,N_49452,N_49453,N_49454,N_49455,N_49456,N_49457,N_49458,N_49459,N_49460,N_49461,N_49462,N_49463,N_49464,N_49465,N_49466,N_49467,N_49468,N_49469,N_49470,N_49471,N_49472,N_49473,N_49474,N_49475,N_49476,N_49477,N_49478,N_49479,N_49480,N_49481,N_49482,N_49483,N_49484,N_49485,N_49486,N_49487,N_49488,N_49489,N_49490,N_49491,N_49492,N_49493,N_49494,N_49495,N_49496,N_49497,N_49498,N_49499,N_49500,N_49501,N_49502,N_49503,N_49504,N_49505,N_49506,N_49507,N_49508,N_49509,N_49510,N_49511,N_49512,N_49513,N_49514,N_49515,N_49516,N_49517,N_49518,N_49519,N_49520,N_49521,N_49522,N_49523,N_49524,N_49525,N_49526,N_49527,N_49528,N_49529,N_49530,N_49531,N_49532,N_49533,N_49534,N_49535,N_49536,N_49537,N_49538,N_49539,N_49540,N_49541,N_49542,N_49543,N_49544,N_49545,N_49546,N_49547,N_49548,N_49549,N_49550,N_49551,N_49552,N_49553,N_49554,N_49555,N_49556,N_49557,N_49558,N_49559,N_49560,N_49561,N_49562,N_49563,N_49564,N_49565,N_49566,N_49567,N_49568,N_49569,N_49570,N_49571,N_49572,N_49573,N_49574,N_49575,N_49576,N_49577,N_49578,N_49579,N_49580,N_49581,N_49582,N_49583,N_49584,N_49585,N_49586,N_49587,N_49588,N_49589,N_49590,N_49591,N_49592,N_49593,N_49594,N_49595,N_49596,N_49597,N_49598,N_49599,N_49600,N_49601,N_49602,N_49603,N_49604,N_49605,N_49606,N_49607,N_49608,N_49609,N_49610,N_49611,N_49612,N_49613,N_49614,N_49615,N_49616,N_49617,N_49618,N_49619,N_49620,N_49621,N_49622,N_49623,N_49624,N_49625,N_49626,N_49627,N_49628,N_49629,N_49630,N_49631,N_49632,N_49633,N_49634,N_49635,N_49636,N_49637,N_49638,N_49639,N_49640,N_49641,N_49642,N_49643,N_49644,N_49645,N_49646,N_49647,N_49648,N_49649,N_49650,N_49651,N_49652,N_49653,N_49654,N_49655,N_49656,N_49657,N_49658,N_49659,N_49660,N_49661,N_49662,N_49663,N_49664,N_49665,N_49666,N_49667,N_49668,N_49669,N_49670,N_49671,N_49672,N_49673,N_49674,N_49675,N_49676,N_49677,N_49678,N_49679,N_49680,N_49681,N_49682,N_49683,N_49684,N_49685,N_49686,N_49687,N_49688,N_49689,N_49690,N_49691,N_49692,N_49693,N_49694,N_49695,N_49696,N_49697,N_49698,N_49699,N_49700,N_49701,N_49702,N_49703,N_49704,N_49705,N_49706,N_49707,N_49708,N_49709,N_49710,N_49711,N_49712,N_49713,N_49714,N_49715,N_49716,N_49717,N_49718,N_49719,N_49720,N_49721,N_49722,N_49723,N_49724,N_49725,N_49726,N_49727,N_49728,N_49729,N_49730,N_49731,N_49732,N_49733,N_49734,N_49735,N_49736,N_49737,N_49738,N_49739,N_49740,N_49741,N_49742,N_49743,N_49744,N_49745,N_49746,N_49747,N_49748,N_49749,N_49750,N_49751,N_49752,N_49753,N_49754,N_49755,N_49756,N_49757,N_49758,N_49759,N_49760,N_49761,N_49762,N_49763,N_49764,N_49765,N_49766,N_49767,N_49768,N_49769,N_49770,N_49771,N_49772,N_49773,N_49774,N_49775,N_49776,N_49777,N_49778,N_49779,N_49780,N_49781,N_49782,N_49783,N_49784,N_49785,N_49786,N_49787,N_49788,N_49789,N_49790,N_49791,N_49792,N_49793,N_49794,N_49795,N_49796,N_49797,N_49798,N_49799,N_49800,N_49801,N_49802,N_49803,N_49804,N_49805,N_49806,N_49807,N_49808,N_49809,N_49810,N_49811,N_49812,N_49813,N_49814,N_49815,N_49816,N_49817,N_49818,N_49819,N_49820,N_49821,N_49822,N_49823,N_49824,N_49825,N_49826,N_49827,N_49828,N_49829,N_49830,N_49831,N_49832,N_49833,N_49834,N_49835,N_49836,N_49837,N_49838,N_49839,N_49840,N_49841,N_49842,N_49843,N_49844,N_49845,N_49846,N_49847,N_49848,N_49849,N_49850,N_49851,N_49852,N_49853,N_49854,N_49855,N_49856,N_49857,N_49858,N_49859,N_49860,N_49861,N_49862,N_49863,N_49864,N_49865,N_49866,N_49867,N_49868,N_49869,N_49870,N_49871,N_49872,N_49873,N_49874,N_49875,N_49876,N_49877,N_49878,N_49879,N_49880,N_49881,N_49882,N_49883,N_49884,N_49885,N_49886,N_49887,N_49888,N_49889,N_49890,N_49891,N_49892,N_49893,N_49894,N_49895,N_49896,N_49897,N_49898,N_49899,N_49900,N_49901,N_49902,N_49903,N_49904,N_49905,N_49906,N_49907,N_49908,N_49909,N_49910,N_49911,N_49912,N_49913,N_49914,N_49915,N_49916,N_49917,N_49918,N_49919,N_49920,N_49921,N_49922,N_49923,N_49924,N_49925,N_49926,N_49927,N_49928,N_49929,N_49930,N_49931,N_49932,N_49933,N_49934,N_49935,N_49936,N_49937,N_49938,N_49939,N_49940,N_49941,N_49942,N_49943,N_49944,N_49945,N_49946,N_49947,N_49948,N_49949,N_49950,N_49951,N_49952,N_49953,N_49954,N_49955,N_49956,N_49957,N_49958,N_49959,N_49960,N_49961,N_49962,N_49963,N_49964,N_49965,N_49966,N_49967,N_49968,N_49969,N_49970,N_49971,N_49972,N_49973,N_49974,N_49975,N_49976,N_49977,N_49978,N_49979,N_49980,N_49981,N_49982,N_49983,N_49984,N_49985,N_49986,N_49987,N_49988,N_49989,N_49990,N_49991,N_49992,N_49993,N_49994,N_49995,N_49996,N_49997,N_49998,N_49999;
and U0 (N_0,In_2855,In_4037);
nand U1 (N_1,In_1330,In_1416);
nand U2 (N_2,In_3950,In_4796);
xnor U3 (N_3,In_4291,In_1362);
nand U4 (N_4,In_1260,In_2255);
and U5 (N_5,In_2417,In_3802);
nor U6 (N_6,In_412,In_3600);
xor U7 (N_7,In_2474,In_3880);
and U8 (N_8,In_2846,In_4385);
xnor U9 (N_9,In_4682,In_1156);
and U10 (N_10,In_975,In_2912);
nor U11 (N_11,In_2445,In_1149);
nand U12 (N_12,In_4940,In_3921);
nor U13 (N_13,In_993,In_3580);
xnor U14 (N_14,In_4775,In_1994);
and U15 (N_15,In_4142,In_65);
and U16 (N_16,In_1973,In_3556);
nand U17 (N_17,In_4692,In_3213);
nand U18 (N_18,In_735,In_3332);
nor U19 (N_19,In_4333,In_3986);
xnor U20 (N_20,In_4585,In_4124);
and U21 (N_21,In_671,In_1244);
and U22 (N_22,In_3043,In_3496);
and U23 (N_23,In_1352,In_2719);
nand U24 (N_24,In_4563,In_1089);
nand U25 (N_25,In_2231,In_893);
and U26 (N_26,In_1694,In_3671);
and U27 (N_27,In_4542,In_1036);
and U28 (N_28,In_3861,In_2318);
nor U29 (N_29,In_4571,In_2394);
xor U30 (N_30,In_4902,In_2539);
nand U31 (N_31,In_3319,In_1006);
and U32 (N_32,In_1502,In_1841);
xor U33 (N_33,In_3073,In_3778);
nand U34 (N_34,In_1842,In_1030);
xnor U35 (N_35,In_3212,In_3529);
nor U36 (N_36,In_4387,In_3981);
nor U37 (N_37,In_703,In_689);
and U38 (N_38,In_3665,In_2325);
or U39 (N_39,In_1458,In_566);
nor U40 (N_40,In_2631,In_2742);
nor U41 (N_41,In_3731,In_3780);
or U42 (N_42,In_743,In_1726);
xnor U43 (N_43,In_1853,In_1474);
xnor U44 (N_44,In_1160,In_4624);
xnor U45 (N_45,In_3104,In_3293);
nand U46 (N_46,In_235,In_285);
nand U47 (N_47,In_4709,In_4031);
and U48 (N_48,In_2448,In_1775);
nor U49 (N_49,In_2213,In_3226);
xnor U50 (N_50,In_1222,In_685);
nand U51 (N_51,In_4306,In_2296);
and U52 (N_52,In_3014,In_3983);
or U53 (N_53,In_1887,In_4664);
nand U54 (N_54,In_4521,In_3416);
xnor U55 (N_55,In_81,In_2570);
or U56 (N_56,In_1417,In_4995);
xnor U57 (N_57,In_4413,In_3174);
nor U58 (N_58,In_632,In_2586);
nor U59 (N_59,In_2739,In_2425);
xnor U60 (N_60,In_3454,In_3973);
or U61 (N_61,In_3412,In_1930);
or U62 (N_62,In_2970,In_612);
nand U63 (N_63,In_4767,In_4164);
and U64 (N_64,In_4791,In_4113);
nor U65 (N_65,In_4093,In_3866);
nor U66 (N_66,In_586,In_3375);
nand U67 (N_67,In_3022,In_3990);
nand U68 (N_68,In_3697,In_1283);
nand U69 (N_69,In_2841,In_2070);
nor U70 (N_70,In_3417,In_4858);
or U71 (N_71,In_2308,In_4803);
and U72 (N_72,In_1540,In_2200);
xor U73 (N_73,In_2391,In_1335);
and U74 (N_74,In_202,In_3009);
nor U75 (N_75,In_2331,In_3456);
nand U76 (N_76,In_3193,In_4684);
or U77 (N_77,In_4356,In_508);
and U78 (N_78,In_4708,In_1146);
or U79 (N_79,In_2625,In_201);
xor U80 (N_80,In_4653,In_1798);
and U81 (N_81,In_705,In_436);
nor U82 (N_82,In_797,In_1159);
or U83 (N_83,In_2190,In_4944);
nor U84 (N_84,In_430,In_2393);
and U85 (N_85,In_1262,In_1252);
xor U86 (N_86,In_867,In_1444);
or U87 (N_87,In_3602,In_114);
or U88 (N_88,In_4513,In_94);
nand U89 (N_89,In_2799,In_2724);
nand U90 (N_90,In_4439,In_2357);
and U91 (N_91,In_3614,In_2864);
and U92 (N_92,In_543,In_4371);
and U93 (N_93,In_2373,In_1738);
xor U94 (N_94,In_3736,In_1210);
nor U95 (N_95,In_719,In_3759);
nor U96 (N_96,In_296,In_2303);
and U97 (N_97,In_1295,In_814);
nand U98 (N_98,In_2648,In_2827);
nor U99 (N_99,In_2085,In_2201);
nor U100 (N_100,In_4667,In_4885);
or U101 (N_101,In_4301,In_681);
nand U102 (N_102,In_3794,In_1009);
nor U103 (N_103,In_1375,In_585);
xnor U104 (N_104,In_1523,In_1715);
nor U105 (N_105,In_70,In_1025);
and U106 (N_106,In_3249,In_223);
or U107 (N_107,In_515,In_832);
and U108 (N_108,In_4710,In_377);
nand U109 (N_109,In_1372,In_4838);
nor U110 (N_110,In_2214,In_781);
nor U111 (N_111,In_1062,In_83);
nand U112 (N_112,In_3534,In_2828);
xnor U113 (N_113,In_1257,In_3808);
nor U114 (N_114,In_3399,In_2588);
nor U115 (N_115,In_315,In_1091);
xor U116 (N_116,In_2626,In_4421);
or U117 (N_117,In_3349,In_2179);
nand U118 (N_118,In_4311,In_4337);
nand U119 (N_119,In_505,In_590);
xor U120 (N_120,In_286,In_3613);
and U121 (N_121,In_644,In_2371);
nand U122 (N_122,In_3976,In_1854);
xnor U123 (N_123,In_297,In_2336);
or U124 (N_124,In_589,In_3136);
nand U125 (N_125,In_3383,In_805);
nor U126 (N_126,In_607,In_2385);
xnor U127 (N_127,In_4038,In_763);
nand U128 (N_128,In_3132,In_3275);
and U129 (N_129,In_654,In_527);
or U130 (N_130,In_1535,In_4140);
nor U131 (N_131,In_4582,In_4888);
nand U132 (N_132,In_4661,In_4131);
and U133 (N_133,In_3724,In_4564);
or U134 (N_134,In_2199,In_2863);
xor U135 (N_135,In_3915,In_1913);
nor U136 (N_136,In_608,In_2156);
or U137 (N_137,In_2203,In_4862);
or U138 (N_138,In_1927,In_1473);
nor U139 (N_139,In_3934,In_3011);
xnor U140 (N_140,In_349,In_1693);
or U141 (N_141,In_427,In_2495);
and U142 (N_142,In_2390,In_599);
nand U143 (N_143,In_876,In_3047);
nor U144 (N_144,In_439,In_3883);
or U145 (N_145,In_3230,In_1341);
xor U146 (N_146,In_629,In_2444);
nand U147 (N_147,In_4778,In_4170);
xor U148 (N_148,In_2433,In_2197);
xor U149 (N_149,In_971,In_4535);
or U150 (N_150,In_2321,In_1097);
and U151 (N_151,In_4242,In_4615);
nand U152 (N_152,In_1580,In_200);
xor U153 (N_153,In_2008,In_1179);
and U154 (N_154,In_4633,In_985);
nor U155 (N_155,In_4467,In_1247);
or U156 (N_156,In_4631,In_3405);
and U157 (N_157,In_4003,In_121);
nand U158 (N_158,In_537,In_3352);
nand U159 (N_159,In_3636,In_1958);
and U160 (N_160,In_4383,In_166);
and U161 (N_161,In_3669,In_4780);
or U162 (N_162,In_2655,In_4919);
nor U163 (N_163,In_1253,In_2581);
nor U164 (N_164,In_2472,In_115);
nand U165 (N_165,In_1668,In_1196);
nand U166 (N_166,In_4695,In_1037);
xnor U167 (N_167,In_2059,In_4688);
nor U168 (N_168,In_718,In_1358);
or U169 (N_169,In_2701,In_1704);
nor U170 (N_170,In_3608,In_1618);
nor U171 (N_171,In_2237,In_3310);
nor U172 (N_172,In_3844,In_2192);
nand U173 (N_173,In_1041,In_4698);
and U174 (N_174,In_1483,In_2731);
nand U175 (N_175,In_791,In_3607);
or U176 (N_176,In_2364,In_4506);
nand U177 (N_177,In_146,In_4915);
nor U178 (N_178,In_1155,In_2830);
or U179 (N_179,In_3453,In_1492);
nand U180 (N_180,In_4308,In_3867);
nor U181 (N_181,In_3092,In_3729);
or U182 (N_182,In_4351,In_597);
xor U183 (N_183,In_2781,In_572);
or U184 (N_184,In_15,In_1943);
or U185 (N_185,In_3234,In_2591);
xor U186 (N_186,In_3793,In_3070);
nand U187 (N_187,In_2412,In_3576);
nor U188 (N_188,In_1129,In_4852);
nand U189 (N_189,In_3348,In_3322);
nor U190 (N_190,In_425,In_1585);
nor U191 (N_191,In_3659,In_4194);
nand U192 (N_192,In_3080,In_1381);
and U193 (N_193,In_402,In_2699);
or U194 (N_194,In_3959,In_1804);
or U195 (N_195,In_1365,In_533);
and U196 (N_196,In_244,In_287);
or U197 (N_197,In_4787,In_3077);
nor U198 (N_198,In_951,In_884);
nand U199 (N_199,In_4686,In_3205);
or U200 (N_200,In_2821,In_2766);
nand U201 (N_201,In_2265,In_3274);
or U202 (N_202,In_7,In_3532);
xor U203 (N_203,In_35,In_38);
and U204 (N_204,In_820,In_2777);
nor U205 (N_205,In_4568,In_1302);
xor U206 (N_206,In_3800,In_101);
xor U207 (N_207,In_2118,In_630);
and U208 (N_208,In_2061,In_3712);
xnor U209 (N_209,In_2587,In_2757);
and U210 (N_210,In_811,In_4908);
nor U211 (N_211,In_3220,In_3864);
nor U212 (N_212,In_4674,In_3770);
or U213 (N_213,In_386,In_856);
and U214 (N_214,In_2184,In_3917);
xnor U215 (N_215,In_2413,In_934);
and U216 (N_216,In_3215,In_2753);
nand U217 (N_217,In_2613,In_25);
or U218 (N_218,In_952,In_1451);
nor U219 (N_219,In_4323,In_2517);
or U220 (N_220,In_3143,In_4580);
or U221 (N_221,In_1370,In_4499);
xnor U222 (N_222,In_1086,In_3173);
or U223 (N_223,In_4445,In_281);
xnor U224 (N_224,In_3579,In_542);
xor U225 (N_225,In_1354,In_1665);
or U226 (N_226,In_3735,In_1412);
nor U227 (N_227,In_963,In_3521);
and U228 (N_228,In_3666,In_1460);
nand U229 (N_229,In_3191,In_451);
and U230 (N_230,In_4732,In_4101);
or U231 (N_231,In_504,In_2131);
or U232 (N_232,In_1655,In_90);
and U233 (N_233,In_3422,In_981);
or U234 (N_234,In_611,In_229);
and U235 (N_235,In_1819,In_4419);
xnor U236 (N_236,In_1767,In_2593);
nor U237 (N_237,In_3895,In_3457);
xor U238 (N_238,In_3195,In_1268);
xor U239 (N_239,In_2353,In_4806);
nor U240 (N_240,In_3640,In_4899);
nand U241 (N_241,In_2469,In_618);
nand U242 (N_242,In_3771,In_1163);
xnor U243 (N_243,In_2531,In_372);
nor U244 (N_244,In_84,In_13);
nor U245 (N_245,In_4330,In_4011);
xor U246 (N_246,In_4001,In_1980);
nand U247 (N_247,In_2801,In_561);
and U248 (N_248,In_306,In_2687);
or U249 (N_249,In_3506,In_4092);
and U250 (N_250,In_110,N_228);
nor U251 (N_251,In_2512,In_3403);
nand U252 (N_252,In_4478,In_4120);
or U253 (N_253,In_4353,In_1939);
nand U254 (N_254,In_2767,In_1813);
and U255 (N_255,In_3218,In_1448);
and U256 (N_256,In_3649,In_1735);
and U257 (N_257,In_2288,In_4203);
nor U258 (N_258,N_10,In_61);
and U259 (N_259,In_1870,In_155);
and U260 (N_260,In_4221,In_1703);
and U261 (N_261,In_12,In_4240);
nand U262 (N_262,In_3936,In_1307);
or U263 (N_263,In_3638,In_3189);
and U264 (N_264,In_1713,In_4596);
or U265 (N_265,In_4953,In_3593);
or U266 (N_266,In_1791,In_2804);
nor U267 (N_267,In_3920,In_1431);
nand U268 (N_268,In_4628,In_2212);
nor U269 (N_269,In_3164,In_4454);
xor U270 (N_270,In_2166,In_4973);
nor U271 (N_271,In_3647,In_2647);
and U272 (N_272,In_1134,In_3054);
and U273 (N_273,In_156,In_2232);
nor U274 (N_274,In_3970,In_3763);
nand U275 (N_275,In_4477,In_4189);
xor U276 (N_276,In_4084,In_391);
nor U277 (N_277,In_2968,In_2260);
xnor U278 (N_278,In_3358,In_3106);
nor U279 (N_279,In_466,In_3592);
nor U280 (N_280,In_1393,In_796);
or U281 (N_281,In_3026,In_3680);
nor U282 (N_282,N_246,In_1578);
or U283 (N_283,In_4462,In_4339);
nand U284 (N_284,In_2065,In_2662);
xnor U285 (N_285,In_3128,In_1424);
and U286 (N_286,In_845,N_144);
nand U287 (N_287,In_2143,In_2868);
or U288 (N_288,In_2481,In_1998);
and U289 (N_289,In_2033,In_1369);
or U290 (N_290,In_1084,In_2350);
xor U291 (N_291,In_4494,In_2494);
or U292 (N_292,In_903,In_3824);
nand U293 (N_293,In_4705,In_4096);
nand U294 (N_294,In_4678,In_905);
xnor U295 (N_295,In_2508,In_2119);
nand U296 (N_296,In_756,In_3367);
and U297 (N_297,In_2461,In_1220);
nand U298 (N_298,N_127,In_481);
and U299 (N_299,In_4157,In_4446);
nand U300 (N_300,N_211,In_4144);
or U301 (N_301,In_852,In_4064);
xor U302 (N_302,N_220,In_844);
and U303 (N_303,In_641,In_4522);
xnor U304 (N_304,In_3338,In_1017);
nor U305 (N_305,In_1374,N_82);
nor U306 (N_306,In_4551,In_2530);
xnor U307 (N_307,In_2025,In_3594);
or U308 (N_308,In_2929,In_4452);
and U309 (N_309,In_779,In_1186);
xor U310 (N_310,In_2022,In_906);
and U311 (N_311,In_2341,In_2520);
nor U312 (N_312,In_950,In_960);
xnor U313 (N_313,In_4177,In_1255);
or U314 (N_314,In_1661,In_4669);
and U315 (N_315,In_2204,In_3281);
xor U316 (N_316,In_4702,In_1422);
nor U317 (N_317,In_4916,In_4008);
nor U318 (N_318,In_2905,In_1629);
nand U319 (N_319,In_1290,In_421);
or U320 (N_320,In_1140,In_2423);
nand U321 (N_321,In_1078,In_2432);
and U322 (N_322,N_131,In_4181);
xor U323 (N_323,In_1581,In_32);
nand U324 (N_324,In_4270,In_765);
or U325 (N_325,In_2458,In_4072);
and U326 (N_326,In_3439,In_4925);
xor U327 (N_327,In_1926,In_1301);
nor U328 (N_328,In_674,In_2479);
nor U329 (N_329,In_67,In_3643);
xnor U330 (N_330,In_4364,In_3084);
xnor U331 (N_331,In_1481,In_4456);
xnor U332 (N_332,In_148,In_2068);
and U333 (N_333,In_2842,In_526);
nand U334 (N_334,In_988,In_2510);
or U335 (N_335,In_638,In_4389);
nor U336 (N_336,In_3152,In_816);
and U337 (N_337,In_4138,In_2723);
and U338 (N_338,In_920,In_4819);
nor U339 (N_339,In_3387,In_3312);
and U340 (N_340,In_4265,In_6);
nand U341 (N_341,In_4483,In_655);
nor U342 (N_342,In_1304,In_2457);
xor U343 (N_343,In_130,In_2388);
or U344 (N_344,In_4079,In_3400);
nor U345 (N_345,In_2568,In_3441);
nor U346 (N_346,In_3503,In_4948);
and U347 (N_347,In_3543,In_3708);
or U348 (N_348,In_569,In_2138);
xor U349 (N_349,In_3407,In_3365);
xnor U350 (N_350,In_2511,In_957);
and U351 (N_351,In_3408,In_2941);
nor U352 (N_352,In_2238,In_3992);
or U353 (N_353,In_2460,In_1122);
xor U354 (N_354,In_2761,In_3085);
xnor U355 (N_355,In_4267,N_68);
nand U356 (N_356,In_167,In_2806);
nor U357 (N_357,In_1048,In_3745);
or U358 (N_358,In_369,N_203);
nor U359 (N_359,In_2148,In_2704);
nor U360 (N_360,In_40,In_2683);
and U361 (N_361,In_1805,In_24);
xnor U362 (N_362,In_497,In_2721);
nor U363 (N_363,In_1872,In_1878);
and U364 (N_364,In_4962,In_2882);
and U365 (N_365,In_2748,In_2125);
nand U366 (N_366,In_2442,In_2285);
and U367 (N_367,In_2465,In_3458);
xnor U368 (N_368,In_2677,In_3185);
nor U369 (N_369,In_3517,In_4062);
or U370 (N_370,In_3393,In_670);
xnor U371 (N_371,In_2410,In_2848);
or U372 (N_372,In_546,In_2538);
nor U373 (N_373,In_302,In_2126);
or U374 (N_374,In_465,In_3072);
nand U375 (N_375,In_915,In_4614);
or U376 (N_376,In_1935,In_716);
and U377 (N_377,In_1909,In_4269);
nand U378 (N_378,In_1031,In_4937);
nand U379 (N_379,In_4500,In_72);
and U380 (N_380,In_753,In_1034);
or U381 (N_381,In_3324,In_3334);
xor U382 (N_382,In_4997,In_3991);
or U383 (N_383,In_1227,In_748);
nand U384 (N_384,In_2694,In_3670);
or U385 (N_385,In_2880,In_2980);
and U386 (N_386,In_2745,In_4466);
and U387 (N_387,In_2159,In_3818);
nor U388 (N_388,In_4910,In_3424);
and U389 (N_389,In_1938,In_3177);
or U390 (N_390,In_2399,In_3364);
or U391 (N_391,In_2437,In_1890);
nor U392 (N_392,In_3301,In_4552);
nand U393 (N_393,In_472,In_3832);
or U394 (N_394,In_3509,In_1243);
or U395 (N_395,In_555,In_2619);
nor U396 (N_396,In_4056,In_2903);
or U397 (N_397,In_1725,In_4459);
xor U398 (N_398,In_1029,In_493);
or U399 (N_399,In_3235,In_1346);
nor U400 (N_400,In_3568,In_2491);
or U401 (N_401,In_3342,In_2650);
nand U402 (N_402,In_978,In_3966);
nand U403 (N_403,In_442,In_2706);
nor U404 (N_404,In_4325,In_606);
xnor U405 (N_405,In_996,In_2076);
and U406 (N_406,In_318,In_274);
xnor U407 (N_407,In_2031,In_1322);
and U408 (N_408,In_4147,In_1357);
nand U409 (N_409,In_1627,In_75);
nor U410 (N_410,In_4475,In_4172);
nor U411 (N_411,In_2895,In_4597);
nand U412 (N_412,In_3756,In_650);
nand U413 (N_413,In_4825,In_517);
xnor U414 (N_414,N_130,In_532);
nand U415 (N_415,In_1053,In_2058);
xor U416 (N_416,In_3696,In_4518);
and U417 (N_417,In_4685,In_4956);
nand U418 (N_418,In_4360,In_1670);
or U419 (N_419,In_463,In_112);
xnor U420 (N_420,In_1808,In_3601);
and U421 (N_421,In_4618,In_3836);
and U422 (N_422,In_2974,In_2326);
xnor U423 (N_423,In_4469,In_4549);
nand U424 (N_424,In_4508,In_2686);
xor U425 (N_425,In_239,In_2775);
or U426 (N_426,In_4436,In_330);
nor U427 (N_427,In_2969,In_3374);
or U428 (N_428,In_4961,In_2533);
nand U429 (N_429,In_4550,In_2947);
or U430 (N_430,In_10,In_2667);
xnor U431 (N_431,In_2555,In_2356);
and U432 (N_432,In_4476,In_2063);
nor U433 (N_433,In_3784,In_4577);
xor U434 (N_434,In_969,In_1136);
or U435 (N_435,In_209,In_3550);
nand U436 (N_436,In_441,In_1166);
xor U437 (N_437,In_1532,In_1686);
or U438 (N_438,In_4137,In_3838);
nand U439 (N_439,In_4813,In_1708);
nand U440 (N_440,In_2840,In_4380);
and U441 (N_441,N_5,In_4800);
or U442 (N_442,In_3748,In_1399);
nor U443 (N_443,In_2612,In_3148);
xor U444 (N_444,In_4130,In_4707);
or U445 (N_445,In_1075,In_185);
nand U446 (N_446,In_3604,N_229);
nor U447 (N_447,In_138,In_1954);
and U448 (N_448,In_687,In_173);
nand U449 (N_449,In_1952,In_1741);
and U450 (N_450,In_4607,In_3535);
nor U451 (N_451,In_1194,In_1530);
xnor U452 (N_452,In_3198,In_1067);
or U453 (N_453,In_2311,In_3062);
nor U454 (N_454,In_690,In_3562);
xor U455 (N_455,In_310,In_1131);
and U456 (N_456,In_2091,In_3008);
and U457 (N_457,In_1669,N_19);
nand U458 (N_458,In_4271,In_639);
or U459 (N_459,In_3237,In_4673);
and U460 (N_460,In_326,In_3385);
nand U461 (N_461,In_3795,In_883);
nor U462 (N_462,In_3524,In_4376);
nand U463 (N_463,In_2547,In_3020);
and U464 (N_464,In_1640,N_181);
nand U465 (N_465,In_2154,In_2716);
nand U466 (N_466,In_2805,In_2219);
or U467 (N_467,In_99,In_1632);
nand U468 (N_468,In_187,In_4158);
nor U469 (N_469,In_2810,In_3757);
xor U470 (N_470,In_2189,In_4790);
nor U471 (N_471,In_849,In_3806);
nand U472 (N_472,In_853,In_2595);
and U473 (N_473,In_1246,N_83);
and U474 (N_474,In_4052,In_534);
and U475 (N_475,In_591,In_1656);
or U476 (N_476,In_3318,In_3609);
nor U477 (N_477,N_158,In_633);
or U478 (N_478,In_2249,In_3672);
and U479 (N_479,In_3380,In_694);
and U480 (N_480,In_1279,In_422);
nor U481 (N_481,N_174,In_2);
or U482 (N_482,In_435,In_2850);
or U483 (N_483,In_2935,In_2602);
xor U484 (N_484,In_243,In_3108);
or U485 (N_485,In_2218,In_1043);
nand U486 (N_486,In_1382,In_3470);
nand U487 (N_487,In_1182,In_4135);
xor U488 (N_488,In_995,In_1527);
xor U489 (N_489,In_2837,In_1486);
or U490 (N_490,In_139,N_31);
xor U491 (N_491,In_1452,In_1800);
xor U492 (N_492,In_1681,In_1742);
nor U493 (N_493,In_3118,In_9);
xor U494 (N_494,N_221,In_376);
or U495 (N_495,In_923,In_3150);
and U496 (N_496,In_4759,In_660);
and U497 (N_497,In_3586,In_1054);
xor U498 (N_498,In_1153,In_4805);
nand U499 (N_499,In_1104,In_1968);
nand U500 (N_500,In_413,N_118);
nand U501 (N_501,In_496,In_3993);
and U502 (N_502,N_22,In_3548);
or U503 (N_503,In_2797,N_58);
nor U504 (N_504,In_445,In_4901);
nand U505 (N_505,In_1019,In_1442);
nor U506 (N_506,In_525,In_3662);
nand U507 (N_507,In_3898,In_4417);
or U508 (N_508,N_477,In_3270);
xnor U509 (N_509,In_429,In_3982);
or U510 (N_510,In_1493,In_3829);
nand U511 (N_511,N_194,In_3569);
nor U512 (N_512,In_3814,N_435);
nand U513 (N_513,In_1617,In_821);
or U514 (N_514,In_4815,N_441);
and U515 (N_515,In_193,In_4126);
xnor U516 (N_516,In_344,In_3553);
nor U517 (N_517,In_1401,In_3239);
or U518 (N_518,In_4715,In_1101);
nand U519 (N_519,In_2525,In_4230);
nor U520 (N_520,In_1730,In_2114);
nand U521 (N_521,In_4763,In_4139);
nor U522 (N_522,N_303,N_451);
nand U523 (N_523,In_3858,N_88);
xnor U524 (N_524,In_4604,N_286);
xnor U525 (N_525,N_80,In_2104);
nor U526 (N_526,In_1045,In_388);
and U527 (N_527,In_490,In_2858);
xor U528 (N_528,In_1482,In_2026);
and U529 (N_529,In_4335,In_3648);
nand U530 (N_530,In_521,In_3112);
nor U531 (N_531,In_3055,In_1436);
nor U532 (N_532,In_3511,In_407);
xor U533 (N_533,In_2529,In_4220);
nor U534 (N_534,In_1112,In_4169);
nand U535 (N_535,In_3980,In_468);
or U536 (N_536,N_92,In_2047);
nor U537 (N_537,In_1165,N_288);
or U538 (N_538,N_425,In_1117);
or U539 (N_539,In_2195,In_1420);
nor U540 (N_540,In_4855,In_4256);
and U541 (N_541,In_4952,In_913);
nor U542 (N_542,In_946,In_4703);
nor U543 (N_543,In_2292,In_1537);
nand U544 (N_544,In_503,N_155);
or U545 (N_545,In_866,In_4262);
nand U546 (N_546,In_1300,In_499);
xnor U547 (N_547,In_181,In_3726);
or U548 (N_548,In_4470,In_935);
nand U549 (N_549,In_2426,In_1941);
nor U550 (N_550,In_3036,In_153);
nand U551 (N_551,N_148,In_2659);
and U552 (N_552,In_4321,In_2055);
xnor U553 (N_553,In_2165,In_2466);
nor U554 (N_554,In_2024,In_4013);
nor U555 (N_555,In_3706,In_1705);
and U556 (N_556,In_3946,In_665);
and U557 (N_557,In_1653,In_3660);
or U558 (N_558,In_2653,In_2916);
xor U559 (N_559,In_838,In_911);
xor U560 (N_560,In_4753,In_4216);
nor U561 (N_561,In_1737,In_3969);
and U562 (N_562,In_4903,In_2149);
or U563 (N_563,In_2594,In_3443);
nor U564 (N_564,In_785,In_4706);
or U565 (N_565,N_372,In_896);
or U566 (N_566,In_1551,In_2488);
and U567 (N_567,In_889,In_2924);
and U568 (N_568,In_478,In_1876);
and U569 (N_569,In_1512,In_3718);
nor U570 (N_570,In_4495,In_224);
xor U571 (N_571,In_1649,In_396);
nor U572 (N_572,In_1541,N_335);
or U573 (N_573,In_3216,In_1749);
or U574 (N_574,In_4350,In_3803);
and U575 (N_575,In_841,N_492);
or U576 (N_576,In_1986,In_1611);
nor U577 (N_577,In_4377,In_368);
or U578 (N_578,In_1193,In_4689);
xor U579 (N_579,In_2136,In_1121);
xnor U580 (N_580,In_3146,In_2036);
and U581 (N_581,In_2869,In_571);
xor U582 (N_582,In_4828,In_3120);
nor U583 (N_583,In_4213,In_1001);
nor U584 (N_584,N_223,In_1667);
nor U585 (N_585,In_1191,In_373);
or U586 (N_586,In_4776,In_1345);
nand U587 (N_587,In_2351,In_788);
xor U588 (N_588,N_409,In_3501);
nand U589 (N_589,In_2281,In_2439);
or U590 (N_590,In_2856,In_144);
and U591 (N_591,N_292,In_1609);
xor U592 (N_592,In_4545,N_287);
or U593 (N_593,In_4457,In_2637);
xnor U594 (N_594,In_2215,In_2576);
or U595 (N_595,In_4666,In_3462);
xor U596 (N_596,In_4965,In_4635);
and U597 (N_597,In_3674,In_2407);
nor U598 (N_598,In_1394,In_2870);
or U599 (N_599,In_3153,In_2345);
xnor U600 (N_600,In_2562,In_564);
and U601 (N_601,In_2178,In_4823);
nand U602 (N_602,In_1409,In_4151);
nand U603 (N_603,N_266,In_1641);
nand U604 (N_604,In_1962,In_1688);
nand U605 (N_605,In_2693,N_54);
and U606 (N_606,In_3279,In_2915);
and U607 (N_607,In_3316,N_281);
and U608 (N_608,In_80,In_2526);
xnor U609 (N_609,In_836,In_3626);
xor U610 (N_610,In_19,In_4829);
xnor U611 (N_611,In_584,In_3523);
and U612 (N_612,In_4020,In_1050);
xnor U613 (N_613,N_14,N_436);
nor U614 (N_614,In_4334,In_4045);
and U615 (N_615,In_4529,In_4771);
nand U616 (N_616,In_1849,In_3109);
nand U617 (N_617,In_404,In_4264);
nor U618 (N_618,In_79,In_0);
nand U619 (N_619,In_2640,In_2352);
or U620 (N_620,In_1893,In_3746);
nand U621 (N_621,In_4832,In_3490);
xnor U622 (N_622,N_362,In_4025);
nand U623 (N_623,In_2583,In_2266);
nand U624 (N_624,In_2630,N_140);
or U625 (N_625,In_3304,In_2770);
nor U626 (N_626,In_118,In_4379);
and U627 (N_627,In_3512,In_741);
or U628 (N_628,In_4282,In_4600);
nand U629 (N_629,In_1100,In_3527);
or U630 (N_630,In_1783,In_1999);
nor U631 (N_631,In_3927,In_3186);
xor U632 (N_632,In_3489,In_2083);
or U633 (N_633,In_1498,In_1896);
xnor U634 (N_634,In_2832,In_4165);
nor U635 (N_635,In_4032,In_3985);
nand U636 (N_636,In_2780,In_833);
nor U637 (N_637,In_4520,In_773);
nor U638 (N_638,In_998,In_4437);
and U639 (N_639,In_3325,In_220);
or U640 (N_640,In_734,In_1151);
nor U641 (N_641,In_953,In_1338);
nor U642 (N_642,In_780,In_3837);
nand U643 (N_643,In_3492,In_4792);
nor U644 (N_644,In_3083,In_3520);
or U645 (N_645,In_4565,In_695);
and U646 (N_646,In_2635,In_1780);
nand U647 (N_647,In_1671,In_1270);
xor U648 (N_648,In_1026,In_3932);
and U649 (N_649,In_3050,In_60);
or U650 (N_650,In_2489,In_4996);
nand U651 (N_651,In_325,N_400);
nand U652 (N_652,In_3192,In_3583);
xor U653 (N_653,In_3488,In_2944);
and U654 (N_654,In_3519,In_916);
and U655 (N_655,In_3840,In_538);
nor U656 (N_656,In_1215,In_4760);
and U657 (N_657,In_4854,In_3874);
or U658 (N_658,In_551,In_2592);
xor U659 (N_659,In_1934,N_166);
nand U660 (N_660,N_164,In_2884);
or U661 (N_661,N_479,In_2191);
and U662 (N_662,In_1079,In_2932);
nor U663 (N_663,In_4382,In_3271);
and U664 (N_664,In_1558,In_4433);
nor U665 (N_665,In_1171,In_410);
nor U666 (N_666,N_66,In_3918);
xnor U667 (N_667,In_3183,In_2956);
or U668 (N_668,In_2559,In_307);
and U669 (N_669,In_1779,In_4438);
nand U670 (N_670,In_2333,In_3370);
nor U671 (N_671,In_2329,In_4224);
and U672 (N_672,In_26,N_231);
nor U673 (N_673,In_3533,In_4894);
xor U674 (N_674,In_102,In_1901);
nand U675 (N_675,In_453,In_4817);
or U676 (N_676,In_3831,In_4091);
or U677 (N_677,N_471,In_3815);
nor U678 (N_678,In_4426,N_306);
nand U679 (N_679,In_862,In_737);
nor U680 (N_680,In_3041,In_1209);
nand U681 (N_681,In_2248,In_4590);
nand U682 (N_682,N_52,In_1709);
or U683 (N_683,In_331,In_3307);
nor U684 (N_684,In_4125,In_1229);
xor U685 (N_685,In_3487,In_4253);
or U686 (N_686,In_4014,In_1894);
nand U687 (N_687,In_899,In_4128);
or U688 (N_688,In_2169,In_236);
nand U689 (N_689,In_2992,In_4517);
or U690 (N_690,In_1747,In_823);
xor U691 (N_691,In_3179,In_1630);
or U692 (N_692,N_375,In_2174);
or U693 (N_693,In_174,In_2392);
xor U694 (N_694,In_4204,In_2017);
or U695 (N_695,In_4583,In_2081);
and U696 (N_696,In_2643,In_720);
nor U697 (N_697,In_987,In_1744);
nand U698 (N_698,In_2816,In_4117);
xor U699 (N_699,In_828,In_4863);
and U700 (N_700,In_4795,In_2454);
nand U701 (N_701,In_1599,In_617);
nand U702 (N_702,In_66,In_4060);
xnor U703 (N_703,In_3833,In_2406);
or U704 (N_704,In_3354,In_3088);
and U705 (N_705,In_338,In_1584);
nand U706 (N_706,In_4726,In_2039);
nand U707 (N_707,In_870,In_4818);
or U708 (N_708,In_2451,In_4028);
nand U709 (N_709,N_332,N_137);
nand U710 (N_710,In_839,In_4842);
xor U711 (N_711,In_147,In_2173);
or U712 (N_712,In_4002,In_1843);
nand U713 (N_713,In_4430,N_485);
or U714 (N_714,In_134,In_2161);
and U715 (N_715,In_4022,In_11);
xor U716 (N_716,In_4704,In_3345);
or U717 (N_717,N_353,N_341);
and U718 (N_718,In_2866,In_3151);
nand U719 (N_719,In_4451,In_4741);
or U720 (N_720,In_1992,In_2194);
and U721 (N_721,In_4789,In_4762);
nor U722 (N_722,In_42,In_4886);
or U723 (N_723,In_4205,In_226);
or U724 (N_724,In_2383,In_4481);
nand U725 (N_725,In_1698,In_2150);
nor U726 (N_726,In_415,In_2235);
nand U727 (N_727,In_1970,In_3886);
and U728 (N_728,In_786,In_2940);
and U729 (N_729,In_383,In_1439);
nor U730 (N_730,In_991,In_2239);
or U731 (N_731,In_1757,In_2106);
or U732 (N_732,In_3446,In_4619);
or U733 (N_733,In_4227,In_2140);
or U734 (N_734,In_4912,In_3116);
nor U735 (N_735,In_4626,In_2242);
and U736 (N_736,In_3907,In_4801);
and U737 (N_737,N_57,In_1566);
or U738 (N_738,In_46,In_312);
xnor U739 (N_739,In_776,In_2902);
nand U740 (N_740,In_4000,In_3021);
and U741 (N_741,In_1177,In_2447);
nand U742 (N_742,In_1543,In_2550);
or U743 (N_743,N_430,In_3048);
nand U744 (N_744,In_4248,In_1339);
and U745 (N_745,In_471,In_3086);
nand U746 (N_746,In_2913,In_3479);
or U747 (N_747,In_1218,N_124);
nand U748 (N_748,In_2558,In_4992);
nand U749 (N_749,In_1786,In_3779);
nor U750 (N_750,In_3438,In_3567);
or U751 (N_751,In_4042,N_588);
xnor U752 (N_752,In_3910,N_365);
xnor U753 (N_753,In_2921,In_190);
and U754 (N_754,In_1175,In_2907);
xnor U755 (N_755,In_1687,In_3952);
nand U756 (N_756,In_2098,In_2086);
or U757 (N_757,In_4332,In_251);
nor U758 (N_758,In_1421,In_1949);
and U759 (N_759,In_4251,In_4979);
xor U760 (N_760,In_1306,In_140);
and U761 (N_761,In_4954,N_621);
nand U762 (N_762,In_4121,In_738);
nand U763 (N_763,In_2290,In_4059);
nor U764 (N_764,In_2270,In_3246);
or U765 (N_765,In_3502,In_818);
and U766 (N_766,In_2812,In_567);
nand U767 (N_767,In_488,In_1398);
or U768 (N_768,In_2134,In_3865);
and U769 (N_769,In_3431,In_770);
nand U770 (N_770,In_2034,In_725);
nor U771 (N_771,In_677,In_736);
nand U772 (N_772,In_4947,In_2524);
nand U773 (N_773,In_1162,In_3373);
or U774 (N_774,In_2395,In_4739);
or U775 (N_775,In_1261,In_3125);
xor U776 (N_776,In_473,In_3835);
and U777 (N_777,In_3225,In_4358);
nor U778 (N_778,In_1405,In_869);
and U779 (N_779,In_3755,In_4747);
nand U780 (N_780,In_1180,In_1024);
nand U781 (N_781,In_1231,N_649);
nand U782 (N_782,In_959,In_228);
and U783 (N_783,In_293,In_4425);
nand U784 (N_784,In_2175,In_2549);
xor U785 (N_785,In_958,In_4700);
and U786 (N_786,In_4810,In_395);
and U787 (N_787,In_300,N_339);
xor U788 (N_788,In_4699,In_2355);
or U789 (N_789,In_1400,In_4694);
and U790 (N_790,In_2691,In_3889);
nor U791 (N_791,In_414,In_50);
and U792 (N_792,In_4352,In_4613);
nor U793 (N_793,In_457,In_1740);
nand U794 (N_794,N_154,In_1418);
nor U795 (N_795,In_4183,In_4843);
and U796 (N_796,In_455,N_299);
or U797 (N_797,In_405,In_850);
nand U798 (N_798,In_3938,In_3327);
or U799 (N_799,In_4869,In_2639);
xnor U800 (N_800,In_1594,In_2823);
or U801 (N_801,In_529,In_3930);
nor U802 (N_802,In_2240,In_3903);
nand U803 (N_803,In_1116,In_1937);
nor U804 (N_804,In_1552,In_1673);
and U805 (N_805,In_4432,In_1951);
nand U806 (N_806,In_4648,In_1081);
or U807 (N_807,In_1505,In_4219);
nand U808 (N_808,In_1862,In_880);
and U809 (N_809,In_3255,In_1010);
xnor U810 (N_810,In_511,In_4543);
nor U811 (N_811,N_578,In_4200);
or U812 (N_812,In_4826,In_1947);
or U813 (N_813,In_2419,In_1087);
nand U814 (N_814,In_2582,In_1823);
nand U815 (N_815,In_1425,In_848);
and U816 (N_816,In_2185,In_4641);
and U817 (N_817,In_1821,In_627);
nor U818 (N_818,In_277,N_738);
or U819 (N_819,In_2875,In_3046);
nand U820 (N_820,In_3162,In_3273);
nor U821 (N_821,In_278,In_2067);
xnor U822 (N_822,In_2785,In_1211);
nand U823 (N_823,In_8,N_147);
nand U824 (N_824,N_172,In_2611);
nor U825 (N_825,N_399,In_1874);
nor U826 (N_826,In_2105,In_1793);
xnor U827 (N_827,In_2943,In_4198);
xnor U828 (N_828,In_4570,In_1454);
xnor U829 (N_829,In_1296,N_422);
or U830 (N_830,N_412,N_689);
or U831 (N_831,In_874,In_3394);
nand U832 (N_832,In_4567,In_672);
nor U833 (N_833,In_1110,In_4289);
and U834 (N_834,In_2347,In_3853);
or U835 (N_835,In_1734,In_4560);
xnor U836 (N_836,In_1965,In_1645);
and U837 (N_837,In_1794,N_606);
nand U838 (N_838,In_1192,In_2089);
xnor U839 (N_839,In_3251,In_3111);
nand U840 (N_840,In_3337,N_648);
xor U841 (N_841,In_3355,In_1500);
and U842 (N_842,In_3896,In_2930);
nor U843 (N_843,In_762,In_3326);
xnor U844 (N_844,In_2003,In_2084);
and U845 (N_845,In_3710,In_1173);
and U846 (N_846,In_4785,In_3471);
xnor U847 (N_847,In_1899,In_728);
xor U848 (N_848,In_1051,In_2142);
xor U849 (N_849,In_808,In_2887);
xor U850 (N_850,In_1835,In_4285);
xor U851 (N_851,N_193,In_1776);
nand U852 (N_852,In_1152,In_3366);
nand U853 (N_853,In_394,In_4073);
and U854 (N_854,N_618,In_1990);
and U855 (N_855,In_370,In_4734);
nor U856 (N_856,In_3634,In_3749);
or U857 (N_857,In_4774,N_289);
or U858 (N_858,In_1508,In_4878);
nor U859 (N_859,In_4553,In_276);
or U860 (N_860,In_3039,In_419);
nor U861 (N_861,In_1202,In_3612);
nor U862 (N_862,In_2793,N_468);
xnor U863 (N_863,In_3254,In_4132);
or U864 (N_864,In_885,In_1837);
nand U865 (N_865,In_603,In_47);
nand U866 (N_866,In_804,In_2756);
xor U867 (N_867,N_535,In_1124);
xor U868 (N_868,N_595,In_613);
and U869 (N_869,In_3811,In_854);
nand U870 (N_870,In_2372,In_891);
nand U871 (N_871,In_3103,In_3415);
or U872 (N_872,In_782,In_136);
nand U873 (N_873,In_1232,In_1976);
and U874 (N_874,In_2962,In_4053);
and U875 (N_875,In_2344,In_2983);
xor U876 (N_876,In_1867,In_2141);
or U877 (N_877,In_4765,In_1602);
or U878 (N_878,In_4866,In_4443);
or U879 (N_879,In_4175,N_37);
nor U880 (N_880,In_3056,In_1240);
nand U881 (N_881,N_391,In_1133);
or U882 (N_882,N_98,In_3804);
or U883 (N_883,In_3061,In_3469);
nor U884 (N_884,In_2945,N_524);
xor U885 (N_885,In_4017,In_3890);
nand U886 (N_886,In_2340,In_4441);
nor U887 (N_887,In_652,N_693);
nand U888 (N_888,In_2965,N_607);
nand U889 (N_889,In_2964,In_4429);
nor U890 (N_890,In_4647,In_1851);
or U891 (N_891,N_671,In_3652);
and U892 (N_892,In_3219,N_668);
or U893 (N_893,In_1190,N_78);
xnor U894 (N_894,In_3909,In_489);
and U895 (N_895,In_2543,In_2702);
or U896 (N_896,In_2540,In_2674);
and U897 (N_897,In_1259,In_518);
nand U898 (N_898,In_604,N_337);
xnor U899 (N_899,In_2977,In_1682);
nand U900 (N_900,In_772,N_102);
xnor U901 (N_901,In_2117,In_4196);
or U902 (N_902,In_456,N_513);
nor U903 (N_903,In_1707,In_1371);
xnor U904 (N_904,In_3611,N_628);
or U905 (N_905,In_4414,In_2979);
or U906 (N_906,In_316,In_4907);
xnor U907 (N_907,In_4864,In_3692);
and U908 (N_908,In_917,In_2224);
nand U909 (N_909,N_568,In_4742);
or U910 (N_910,In_2917,In_382);
nor U911 (N_911,In_3280,N_491);
or U912 (N_912,In_361,In_1093);
xnor U913 (N_913,In_2480,In_2450);
nand U914 (N_914,In_1950,In_2295);
or U915 (N_915,In_1717,In_3821);
or U916 (N_916,In_4779,In_640);
nand U917 (N_917,In_3409,In_3114);
or U918 (N_918,In_1342,In_4629);
and U919 (N_919,In_31,In_1663);
nor U920 (N_920,In_1539,N_176);
nand U921 (N_921,In_1525,In_3870);
nor U922 (N_922,In_2709,N_146);
nand U923 (N_923,In_942,In_4035);
or U924 (N_924,In_2302,In_2103);
and U925 (N_925,In_4788,In_3984);
nand U926 (N_926,N_151,N_70);
or U927 (N_927,In_2306,In_4039);
or U928 (N_928,In_168,N_113);
nor U929 (N_929,In_4328,In_1900);
nand U930 (N_930,In_1105,In_4960);
nor U931 (N_931,N_539,In_2075);
nor U932 (N_932,In_203,In_141);
and U933 (N_933,In_2343,In_771);
xor U934 (N_934,In_2102,In_3528);
nor U935 (N_935,In_4616,In_580);
and U936 (N_936,In_824,In_2464);
xor U937 (N_937,In_789,In_4455);
and U938 (N_938,N_305,In_4407);
or U939 (N_939,In_4086,In_2942);
or U940 (N_940,In_2155,In_2991);
and U941 (N_941,In_3633,In_3598);
nand U942 (N_942,In_3774,In_125);
nor U943 (N_943,In_1479,In_2405);
and U944 (N_944,In_91,In_4578);
or U945 (N_945,In_2483,In_746);
nor U946 (N_946,In_143,N_133);
xor U947 (N_947,In_594,In_999);
nand U948 (N_948,In_1604,In_177);
or U949 (N_949,In_1188,In_3291);
and U950 (N_950,In_653,In_4955);
nand U951 (N_951,In_4918,In_375);
nand U952 (N_952,In_2628,In_3842);
or U953 (N_953,N_660,In_803);
xor U954 (N_954,In_3495,In_2553);
nor U955 (N_955,In_766,In_1565);
and U956 (N_956,In_2914,N_403);
nor U957 (N_957,In_3852,In_3933);
nor U958 (N_958,In_398,In_592);
xnor U959 (N_959,In_619,In_2513);
xor U960 (N_960,In_2901,N_189);
or U961 (N_961,In_280,In_262);
xnor U962 (N_962,In_1569,In_1195);
and U963 (N_963,In_596,N_548);
xnor U964 (N_964,In_4388,In_4720);
and U965 (N_965,In_1921,N_313);
nor U966 (N_966,In_1971,In_3905);
nor U967 (N_967,In_2004,In_4365);
or U968 (N_968,In_2441,In_2015);
or U969 (N_969,In_1865,In_601);
or U970 (N_970,In_2692,In_3734);
nand U971 (N_971,In_3099,In_3472);
xnor U972 (N_972,In_730,In_4909);
xnor U973 (N_973,In_313,In_3244);
or U974 (N_974,In_759,In_2182);
nand U975 (N_975,In_2988,In_4275);
nor U976 (N_976,In_3421,In_3711);
nand U977 (N_977,In_492,In_409);
nor U978 (N_978,N_531,N_324);
nor U979 (N_979,In_2334,In_3767);
nand U980 (N_980,In_1450,N_583);
nor U981 (N_981,In_4561,In_807);
or U982 (N_982,In_3994,In_4598);
nor U983 (N_983,In_3376,In_937);
nand U984 (N_984,In_4835,In_2627);
xnor U985 (N_985,In_1993,In_536);
xor U986 (N_986,In_4636,In_44);
and U987 (N_987,In_3141,In_3082);
xor U988 (N_988,In_1511,In_4584);
and U989 (N_989,In_3683,In_1606);
xnor U990 (N_990,In_4811,In_1612);
and U991 (N_991,In_755,In_4814);
nor U992 (N_992,In_3641,In_1510);
or U993 (N_993,In_1600,In_1648);
nand U994 (N_994,N_608,In_3728);
nand U995 (N_995,In_4300,In_4872);
nor U996 (N_996,In_157,In_1877);
and U997 (N_997,In_2431,In_3060);
xnor U998 (N_998,In_954,In_4502);
or U999 (N_999,In_1478,In_1833);
and U1000 (N_1000,In_4949,In_3248);
nor U1001 (N_1001,In_4186,N_741);
and U1002 (N_1002,In_1123,In_2108);
xor U1003 (N_1003,In_3003,In_1464);
and U1004 (N_1004,In_506,In_4612);
and U1005 (N_1005,In_3515,In_1343);
xor U1006 (N_1006,In_3761,In_3657);
nand U1007 (N_1007,In_2851,In_4276);
nand U1008 (N_1008,In_1183,N_676);
and U1009 (N_1009,In_2661,In_837);
and U1010 (N_1010,In_374,N_967);
nand U1011 (N_1011,In_1360,In_479);
nor U1012 (N_1012,In_1864,In_2397);
xor U1013 (N_1013,In_4773,In_2931);
xnor U1014 (N_1014,In_2471,N_724);
or U1015 (N_1015,In_3178,In_3154);
nor U1016 (N_1016,In_666,N_675);
xnor U1017 (N_1017,In_3695,In_693);
xor U1018 (N_1018,In_3559,In_2835);
or U1019 (N_1019,In_4041,N_690);
or U1020 (N_1020,In_4523,In_2287);
nor U1021 (N_1021,In_4115,In_2629);
nor U1022 (N_1022,N_114,In_1654);
xor U1023 (N_1023,In_2300,In_1658);
nor U1024 (N_1024,In_1546,In_3742);
nand U1025 (N_1025,In_1413,N_887);
nand U1026 (N_1026,In_2786,In_4770);
or U1027 (N_1027,In_4016,In_164);
nand U1028 (N_1028,N_502,In_3691);
nor U1029 (N_1029,In_1605,In_2206);
or U1030 (N_1030,In_1200,In_4679);
nor U1031 (N_1031,In_1758,In_3560);
nand U1032 (N_1032,In_3988,N_418);
nand U1033 (N_1033,In_990,In_1293);
nand U1034 (N_1034,In_1564,In_4677);
nand U1035 (N_1035,In_21,In_222);
xnor U1036 (N_1036,N_881,In_1083);
nor U1037 (N_1037,In_2367,In_4722);
nand U1038 (N_1038,In_336,In_1680);
nand U1039 (N_1039,In_4259,In_4098);
nor U1040 (N_1040,In_100,In_3155);
xnor U1041 (N_1041,In_1003,In_2571);
and U1042 (N_1042,In_2453,In_179);
or U1043 (N_1043,In_3513,N_134);
and U1044 (N_1044,In_2700,In_1320);
nor U1045 (N_1045,In_4724,In_1714);
xor U1046 (N_1046,In_3058,In_2177);
nor U1047 (N_1047,In_1995,In_4994);
nor U1048 (N_1048,In_3940,In_1015);
nor U1049 (N_1049,In_1521,In_2163);
xor U1050 (N_1050,In_4163,In_605);
nand U1051 (N_1051,In_4047,In_3701);
and U1052 (N_1052,N_802,N_517);
nand U1053 (N_1053,In_4680,In_2656);
nor U1054 (N_1054,In_4192,In_3372);
nor U1055 (N_1055,In_2668,N_500);
nor U1056 (N_1056,In_1692,In_4516);
nor U1057 (N_1057,N_538,N_630);
xor U1058 (N_1058,In_1732,N_843);
nor U1059 (N_1059,In_3738,In_3733);
xnor U1060 (N_1060,In_3787,N_759);
nor U1061 (N_1061,In_3159,N_464);
and U1062 (N_1062,In_2633,In_879);
nor U1063 (N_1063,N_792,In_4737);
nor U1064 (N_1064,N_987,In_4748);
xor U1065 (N_1065,In_359,In_362);
xor U1066 (N_1066,In_3330,N_81);
xor U1067 (N_1067,In_4743,In_2152);
nor U1068 (N_1068,In_562,In_3796);
nand U1069 (N_1069,In_1435,In_2527);
xor U1070 (N_1070,In_2985,N_216);
nor U1071 (N_1071,In_4754,In_4280);
or U1072 (N_1072,In_4634,In_3526);
nor U1073 (N_1073,In_2107,N_888);
xor U1074 (N_1074,In_1403,In_4318);
nand U1075 (N_1075,N_566,In_2564);
xor U1076 (N_1076,In_1419,In_3450);
and U1077 (N_1077,In_4893,N_239);
xor U1078 (N_1078,N_632,In_1586);
nor U1079 (N_1079,In_4993,In_2028);
nand U1080 (N_1080,N_95,In_20);
xnor U1081 (N_1081,N_977,In_4964);
or U1082 (N_1082,In_1223,In_3505);
nor U1083 (N_1083,N_960,In_64);
or U1084 (N_1084,In_1816,N_141);
nand U1085 (N_1085,In_440,In_170);
nand U1086 (N_1086,In_3823,N_786);
xnor U1087 (N_1087,N_62,In_2228);
nor U1088 (N_1088,In_1044,In_4191);
or U1089 (N_1089,In_4404,In_895);
nor U1090 (N_1090,In_2193,In_4736);
and U1091 (N_1091,In_4548,N_268);
nor U1092 (N_1092,In_4786,In_3707);
nor U1093 (N_1093,In_2598,In_3482);
xnor U1094 (N_1094,In_1312,In_1);
or U1095 (N_1095,In_2144,In_4304);
and U1096 (N_1096,In_1787,In_2563);
nand U1097 (N_1097,N_599,In_3314);
xnor U1098 (N_1098,In_1724,In_4687);
and U1099 (N_1099,In_3025,In_2429);
and U1100 (N_1100,In_2561,In_1021);
xnor U1101 (N_1101,In_1353,In_4296);
nand U1102 (N_1102,In_1891,In_423);
xnor U1103 (N_1103,In_1472,In_4544);
or U1104 (N_1104,In_1555,In_393);
nor U1105 (N_1105,In_1073,In_3360);
and U1106 (N_1106,In_4156,In_3196);
xor U1107 (N_1107,In_3006,N_765);
xnor U1108 (N_1108,In_4394,In_2016);
xor U1109 (N_1109,In_3351,In_1528);
nor U1110 (N_1110,In_1298,In_1059);
nor U1111 (N_1111,In_2361,In_744);
nor U1112 (N_1112,N_336,In_1098);
xor U1113 (N_1113,In_2283,In_938);
xor U1114 (N_1114,In_732,In_4110);
nand U1115 (N_1115,In_625,In_4851);
or U1116 (N_1116,In_3053,In_4099);
nor U1117 (N_1117,N_282,N_537);
nand U1118 (N_1118,In_556,In_965);
or U1119 (N_1119,N_645,N_476);
nand U1120 (N_1120,N_704,In_1731);
nand U1121 (N_1121,N_858,In_4769);
nand U1122 (N_1122,N_467,In_2789);
nand U1123 (N_1123,In_2726,N_575);
nor U1124 (N_1124,In_2541,In_2111);
nand U1125 (N_1125,In_1674,In_1204);
or U1126 (N_1126,In_2710,N_758);
and U1127 (N_1127,In_2254,In_3635);
nand U1128 (N_1128,In_4207,N_753);
nor U1129 (N_1129,In_4480,In_822);
nor U1130 (N_1130,In_2514,In_2146);
or U1131 (N_1131,In_1347,In_2052);
or U1132 (N_1132,In_502,In_1313);
or U1133 (N_1133,In_3893,N_414);
nor U1134 (N_1134,N_190,N_707);
nor U1135 (N_1135,In_3571,In_2836);
xor U1136 (N_1136,In_3436,In_563);
xor U1137 (N_1137,In_3591,In_2299);
xnor U1138 (N_1138,N_863,In_3584);
nand U1139 (N_1139,In_1462,In_851);
or U1140 (N_1140,In_39,In_800);
and U1141 (N_1141,N_717,N_395);
nor U1142 (N_1142,In_4821,In_1225);
or U1143 (N_1143,In_1942,In_389);
or U1144 (N_1144,N_235,In_4804);
or U1145 (N_1145,N_781,N_434);
xor U1146 (N_1146,In_2455,In_4312);
or U1147 (N_1147,N_665,In_2845);
and U1148 (N_1148,In_1005,N_504);
nand U1149 (N_1149,In_2380,N_705);
nand U1150 (N_1150,In_1719,In_4405);
and U1151 (N_1151,In_1289,In_4654);
or U1152 (N_1152,In_3541,In_2280);
nand U1153 (N_1153,In_4558,In_1868);
nor U1154 (N_1154,In_4222,In_4900);
nand U1155 (N_1155,In_2542,In_600);
nor U1156 (N_1156,In_2427,In_3595);
or U1157 (N_1157,N_136,N_801);
nand U1158 (N_1158,N_943,In_171);
and U1159 (N_1159,In_840,In_3032);
nor U1160 (N_1160,In_33,In_2462);
and U1161 (N_1161,N_25,In_700);
nor U1162 (N_1162,In_1562,In_1788);
or U1163 (N_1163,In_4807,N_277);
nor U1164 (N_1164,In_215,In_2718);
nor U1165 (N_1165,In_3494,In_2035);
and U1166 (N_1166,In_261,In_1174);
xnor U1167 (N_1167,N_909,In_579);
and U1168 (N_1168,In_2452,N_420);
xnor U1169 (N_1169,In_1348,In_1164);
nand U1170 (N_1170,In_2073,In_4197);
or U1171 (N_1171,In_1961,In_2071);
nand U1172 (N_1172,In_1476,In_3765);
xnor U1173 (N_1173,N_710,In_3484);
nor U1174 (N_1174,N_4,In_1294);
or U1175 (N_1175,N_200,In_3972);
xnor U1176 (N_1176,N_844,In_4070);
and U1177 (N_1177,In_1233,N_319);
nand U1178 (N_1178,N_32,In_3854);
nand U1179 (N_1179,In_3211,In_3435);
and U1180 (N_1180,In_624,In_3906);
nor U1181 (N_1181,In_2069,In_873);
nand U1182 (N_1182,In_4112,In_3432);
nand U1183 (N_1183,In_4479,In_63);
xor U1184 (N_1184,In_1912,In_3813);
xor U1185 (N_1185,In_1485,N_63);
or U1186 (N_1186,In_3224,In_4307);
nor U1187 (N_1187,N_859,In_3564);
or U1188 (N_1188,N_634,In_4740);
nor U1189 (N_1189,N_273,In_14);
and U1190 (N_1190,N_815,In_476);
or U1191 (N_1191,N_226,In_986);
or U1192 (N_1192,In_1187,In_3002);
nand U1193 (N_1193,In_813,N_940);
and U1194 (N_1194,In_930,In_4696);
nor U1195 (N_1195,In_1642,In_3369);
nor U1196 (N_1196,In_4418,In_2874);
and U1197 (N_1197,In_4950,N_768);
or U1198 (N_1198,In_3998,N_866);
or U1199 (N_1199,In_2703,In_2713);
or U1200 (N_1200,N_86,In_1497);
nand U1201 (N_1201,In_3019,In_2783);
or U1202 (N_1202,In_1766,In_4228);
xnor U1203 (N_1203,In_178,N_358);
and U1204 (N_1204,In_2037,N_816);
nor U1205 (N_1205,In_1109,N_679);
nand U1206 (N_1206,In_2428,In_1277);
and U1207 (N_1207,In_3267,In_131);
or U1208 (N_1208,In_2275,In_1150);
and U1209 (N_1209,In_2220,N_998);
or U1210 (N_1210,In_575,In_2808);
nand U1211 (N_1211,N_508,In_1315);
or U1212 (N_1212,N_67,In_3944);
nand U1213 (N_1213,In_2271,N_49);
nor U1214 (N_1214,In_4007,In_2261);
or U1215 (N_1215,In_3135,In_1120);
or U1216 (N_1216,N_896,N_656);
nor U1217 (N_1217,In_798,In_2377);
xor U1218 (N_1218,In_983,In_309);
and U1219 (N_1219,In_3068,In_2348);
or U1220 (N_1220,In_1636,In_4257);
or U1221 (N_1221,N_874,N_514);
nor U1222 (N_1222,In_909,In_1845);
xnor U1223 (N_1223,In_4921,In_1914);
xor U1224 (N_1224,In_3382,N_647);
nor U1225 (N_1225,In_4606,In_1792);
nor U1226 (N_1226,In_892,In_2839);
or U1227 (N_1227,In_2993,In_616);
xnor U1228 (N_1228,In_2362,In_4797);
nand U1229 (N_1229,In_52,N_822);
xnor U1230 (N_1230,N_951,In_2305);
xor U1231 (N_1231,In_4395,In_1828);
or U1232 (N_1232,In_1675,In_1588);
nor U1233 (N_1233,N_677,In_4048);
xor U1234 (N_1234,In_2554,N_830);
and U1235 (N_1235,In_4261,In_4733);
xnor U1236 (N_1236,In_859,In_3016);
nand U1237 (N_1237,In_1226,N_553);
and U1238 (N_1238,N_958,In_3445);
or U1239 (N_1239,N_18,In_1201);
and U1240 (N_1240,In_1310,In_452);
nand U1241 (N_1241,In_3536,N_29);
nand U1242 (N_1242,In_1007,In_3974);
xor U1243 (N_1243,In_2608,In_4460);
and U1244 (N_1244,N_300,N_549);
nand U1245 (N_1245,In_4294,In_4055);
or U1246 (N_1246,In_3939,In_1889);
xor U1247 (N_1247,In_2807,In_4024);
or U1248 (N_1248,In_1414,In_3406);
nand U1249 (N_1249,In_2252,In_3090);
nand U1250 (N_1250,In_2776,N_934);
nand U1251 (N_1251,In_23,In_2857);
or U1252 (N_1252,In_3028,In_4374);
nand U1253 (N_1253,In_4920,In_3161);
nand U1254 (N_1254,In_4106,N_853);
nor U1255 (N_1255,In_4174,In_871);
nand U1256 (N_1256,In_4830,N_854);
and U1257 (N_1257,In_4608,In_218);
nor U1258 (N_1258,N_96,In_570);
and U1259 (N_1259,In_3900,In_1545);
nor U1260 (N_1260,In_2346,N_308);
and U1261 (N_1261,N_243,In_2358);
xor U1262 (N_1262,In_1879,In_2695);
and U1263 (N_1263,N_340,In_448);
nand U1264 (N_1264,In_3180,In_3599);
nor U1265 (N_1265,In_3754,N_215);
nor U1266 (N_1266,N_501,In_2738);
or U1267 (N_1267,In_2157,In_4936);
nand U1268 (N_1268,In_4399,N_1128);
or U1269 (N_1269,In_2116,In_3289);
or U1270 (N_1270,In_1060,In_3891);
xnor U1271 (N_1271,In_2051,In_2618);
nand U1272 (N_1272,N_346,N_55);
and U1273 (N_1273,In_2045,In_1633);
or U1274 (N_1274,In_528,N_139);
nand U1275 (N_1275,N_232,In_1438);
nor U1276 (N_1276,In_82,In_1230);
xnor U1277 (N_1277,In_1272,N_864);
and U1278 (N_1278,In_3663,N_580);
nor U1279 (N_1279,In_636,In_2043);
or U1280 (N_1280,N_487,In_4283);
xnor U1281 (N_1281,In_3098,In_1721);
xor U1282 (N_1282,N_680,N_1247);
xnor U1283 (N_1283,In_4076,In_3362);
or U1284 (N_1284,In_192,In_548);
nor U1285 (N_1285,In_1314,In_4988);
or U1286 (N_1286,In_2957,In_2876);
nor U1287 (N_1287,In_645,In_2649);
nand U1288 (N_1288,In_582,In_4427);
nor U1289 (N_1289,In_752,In_3395);
or U1290 (N_1290,In_2291,In_1626);
and U1291 (N_1291,N_506,In_3411);
xor U1292 (N_1292,In_3181,N_370);
xor U1293 (N_1293,In_507,In_3485);
and U1294 (N_1294,In_3621,N_117);
and U1295 (N_1295,N_454,N_488);
and U1296 (N_1296,In_3347,In_4268);
and U1297 (N_1297,In_922,In_4655);
or U1298 (N_1298,In_460,In_3623);
nand U1299 (N_1299,In_760,N_163);
nand U1300 (N_1300,In_3925,In_4620);
xnor U1301 (N_1301,In_2606,N_316);
and U1302 (N_1302,In_3943,In_4572);
nand U1303 (N_1303,In_1959,In_2387);
nor U1304 (N_1304,N_429,In_284);
nor U1305 (N_1305,In_1513,In_109);
and U1306 (N_1306,N_667,In_3144);
nand U1307 (N_1307,N_344,N_882);
or U1308 (N_1308,In_1094,N_377);
or U1309 (N_1309,In_1883,In_2315);
nand U1310 (N_1310,In_3290,In_1066);
nand U1311 (N_1311,In_3015,In_2987);
and U1312 (N_1312,In_4971,In_3862);
nand U1313 (N_1313,In_4252,In_3551);
or U1314 (N_1314,N_1096,In_2791);
nand U1315 (N_1315,In_1396,N_36);
xor U1316 (N_1316,In_3545,In_3546);
xor U1317 (N_1317,N_1107,In_1773);
xnor U1318 (N_1318,N_725,In_129);
and U1319 (N_1319,In_4836,In_2802);
xnor U1320 (N_1320,In_3121,In_2181);
xnor U1321 (N_1321,In_2535,N_730);
nor U1322 (N_1322,In_1906,In_1333);
and U1323 (N_1323,In_4303,In_4892);
or U1324 (N_1324,N_752,N_312);
or U1325 (N_1325,In_2443,N_600);
and U1326 (N_1326,In_3188,N_132);
nand U1327 (N_1327,N_769,N_1068);
or U1328 (N_1328,N_108,N_90);
and U1329 (N_1329,In_2014,In_715);
and U1330 (N_1330,In_2322,In_3554);
nor U1331 (N_1331,N_1215,In_3194);
nand U1332 (N_1332,N_692,In_4645);
xnor U1333 (N_1333,N_348,In_3306);
nand U1334 (N_1334,In_1299,In_4005);
or U1335 (N_1335,N_809,In_2459);
and U1336 (N_1336,In_2680,In_2297);
xor U1337 (N_1337,N_1225,In_2509);
xor U1338 (N_1338,N_589,In_2368);
xnor U1339 (N_1339,N_1174,N_763);
xor U1340 (N_1340,In_3741,In_183);
xor U1341 (N_1341,In_2032,In_2366);
xor U1342 (N_1342,N_661,In_1556);
or U1343 (N_1343,In_926,N_819);
nor U1344 (N_1344,N_994,In_1979);
xnor U1345 (N_1345,In_434,In_3074);
nand U1346 (N_1346,In_956,In_93);
xnor U1347 (N_1347,In_159,In_2312);
or U1348 (N_1348,N_590,N_530);
or U1349 (N_1349,In_365,N_361);
or U1350 (N_1350,In_1297,In_3260);
nand U1351 (N_1351,In_2113,N_1218);
xnor U1352 (N_1352,N_619,In_3667);
and U1353 (N_1353,N_610,In_34);
xor U1354 (N_1354,In_4397,In_3777);
or U1355 (N_1355,In_2714,In_1754);
or U1356 (N_1356,In_3768,In_3963);
and U1357 (N_1357,In_2012,In_2638);
nor U1358 (N_1358,In_1154,N_933);
xor U1359 (N_1359,N_106,In_4336);
nand U1360 (N_1360,In_4095,In_1929);
nor U1361 (N_1361,N_53,In_1997);
nand U1362 (N_1362,In_2147,In_2205);
or U1363 (N_1363,In_3884,N_900);
xor U1364 (N_1364,N_245,In_2877);
or U1365 (N_1365,In_4329,In_2897);
nor U1366 (N_1366,In_1852,In_1660);
nand U1367 (N_1367,In_2078,In_2363);
and U1368 (N_1368,In_385,N_826);
or U1369 (N_1369,In_4279,In_4327);
nor U1370 (N_1370,In_3157,In_4018);
nor U1371 (N_1371,In_1466,In_2729);
and U1372 (N_1372,In_882,In_2006);
or U1373 (N_1373,In_1554,In_1022);
nor U1374 (N_1374,In_1241,N_94);
nand U1375 (N_1375,N_256,N_405);
nand U1376 (N_1376,In_1615,In_1366);
xnor U1377 (N_1377,In_1363,In_2599);
nor U1378 (N_1378,N_222,In_1217);
xor U1379 (N_1379,In_4129,N_1181);
xor U1380 (N_1380,In_1996,In_4396);
xnor U1381 (N_1381,N_386,In_927);
xnor U1382 (N_1382,In_1768,N_452);
xnor U1383 (N_1383,N_914,N_159);
nor U1384 (N_1384,N_1027,In_4134);
and U1385 (N_1385,N_637,In_3410);
and U1386 (N_1386,In_2122,In_3126);
and U1387 (N_1387,In_544,N_1190);
nand U1388 (N_1388,In_4012,In_2301);
xnor U1389 (N_1389,N_574,N_597);
xnor U1390 (N_1390,N_1062,N_961);
nand U1391 (N_1391,In_4004,In_1631);
nand U1392 (N_1392,In_3418,In_815);
xor U1393 (N_1393,In_4882,In_347);
nand U1394 (N_1394,In_2337,In_213);
and U1395 (N_1395,N_271,In_1457);
nor U1396 (N_1396,In_522,In_2663);
xnor U1397 (N_1397,In_890,N_351);
and U1398 (N_1398,In_2434,In_1070);
xor U1399 (N_1399,N_654,In_749);
nor U1400 (N_1400,In_790,In_1815);
nor U1401 (N_1401,In_1027,In_3175);
xor U1402 (N_1402,In_767,N_244);
nor U1403 (N_1403,In_3888,In_2002);
nor U1404 (N_1404,In_211,In_2516);
nand U1405 (N_1405,N_1131,In_22);
xnor U1406 (N_1406,In_3877,In_2536);
xor U1407 (N_1407,In_976,In_2170);
and U1408 (N_1408,In_180,N_41);
and U1409 (N_1409,In_3816,In_3850);
nand U1410 (N_1410,In_4484,In_279);
and U1411 (N_1411,N_895,In_810);
nand U1412 (N_1412,In_3951,In_4363);
nor U1413 (N_1413,In_459,In_1571);
nor U1414 (N_1414,In_1803,In_4185);
nand U1415 (N_1415,In_1251,In_2468);
xor U1416 (N_1416,In_1321,In_4537);
xor U1417 (N_1417,In_1088,In_4258);
and U1418 (N_1418,N_1103,In_2482);
xnor U1419 (N_1419,N_267,In_4370);
and U1420 (N_1420,N_354,N_440);
nor U1421 (N_1421,In_2728,In_3261);
xnor U1422 (N_1422,In_2532,In_3228);
and U1423 (N_1423,In_3752,In_1518);
or U1424 (N_1424,In_3642,In_1443);
and U1425 (N_1425,In_2523,In_4932);
xnor U1426 (N_1426,N_811,In_2537);
xnor U1427 (N_1427,In_2744,N_91);
or U1428 (N_1428,In_2153,In_3294);
or U1429 (N_1429,In_4554,In_4412);
nand U1430 (N_1430,N_742,In_547);
nand U1431 (N_1431,In_3138,In_3876);
nand U1432 (N_1432,N_1013,In_3451);
nor U1433 (N_1433,N_257,In_2463);
and U1434 (N_1434,N_426,N_544);
nor U1435 (N_1435,N_701,In_3197);
nand U1436 (N_1436,In_1208,N_1110);
nor U1437 (N_1437,In_2651,In_2620);
nand U1438 (N_1438,N_352,In_2044);
nand U1439 (N_1439,In_657,In_4292);
or U1440 (N_1440,In_1903,In_2256);
or U1441 (N_1441,In_2233,N_554);
xnor U1442 (N_1442,In_4299,N_1163);
or U1443 (N_1443,In_2545,In_1572);
and U1444 (N_1444,In_1318,In_1142);
nor U1445 (N_1445,N_162,In_1774);
and U1446 (N_1446,In_857,In_498);
nor U1447 (N_1447,In_2948,N_995);
xnor U1448 (N_1448,In_3130,In_4234);
nand U1449 (N_1449,In_352,In_2167);
nor U1450 (N_1450,In_2580,In_2422);
and U1451 (N_1451,In_230,N_651);
xnor U1452 (N_1452,In_688,In_3846);
xor U1453 (N_1453,In_339,N_458);
xnor U1454 (N_1454,In_947,In_3140);
xnor U1455 (N_1455,In_1639,N_702);
xor U1456 (N_1456,In_401,In_392);
or U1457 (N_1457,N_7,In_711);
or U1458 (N_1458,N_396,In_2528);
or U1459 (N_1459,In_2666,In_3344);
nand U1460 (N_1460,In_881,In_1795);
or U1461 (N_1461,In_2202,N_489);
xnor U1462 (N_1462,N_837,In_3202);
and U1463 (N_1463,In_1392,N_1184);
or U1464 (N_1464,In_3115,In_4);
nor U1465 (N_1465,N_571,In_3134);
or U1466 (N_1466,In_3071,In_3137);
or U1467 (N_1467,In_3913,In_2725);
nor U1468 (N_1468,N_879,In_1570);
and U1469 (N_1469,N_891,N_263);
xor U1470 (N_1470,N_1137,N_1043);
nand U1471 (N_1471,In_4941,In_4026);
nor U1472 (N_1472,In_3388,N_953);
or U1473 (N_1473,In_3333,N_635);
xnor U1474 (N_1474,In_2579,N_808);
and U1475 (N_1475,In_4357,In_273);
or U1476 (N_1476,In_2521,In_3052);
or U1477 (N_1477,In_3845,In_3096);
xnor U1478 (N_1478,In_4313,In_1496);
or U1479 (N_1479,In_2751,In_2614);
or U1480 (N_1480,N_1111,In_2873);
xnor U1481 (N_1481,N_1040,In_4525);
nand U1482 (N_1482,In_2168,In_3483);
nor U1483 (N_1483,In_1329,N_521);
nand U1484 (N_1484,N_551,In_2269);
nand U1485 (N_1485,In_1677,In_3679);
or U1486 (N_1486,N_371,In_3057);
nor U1487 (N_1487,In_2953,In_366);
xor U1488 (N_1488,In_4989,In_4744);
nor U1489 (N_1489,In_1531,In_1826);
xnor U1490 (N_1490,In_2707,N_1173);
or U1491 (N_1491,In_2369,In_4254);
nor U1492 (N_1492,In_3740,In_4725);
nor U1493 (N_1493,In_2600,In_248);
or U1494 (N_1494,In_4853,In_1922);
nand U1495 (N_1495,In_324,In_4519);
nand U1496 (N_1496,In_3158,N_727);
xnor U1497 (N_1497,In_4496,In_2849);
or U1498 (N_1498,In_1340,In_1748);
xnor U1499 (N_1499,N_573,In_3753);
nor U1500 (N_1500,In_1700,N_804);
xnor U1501 (N_1501,N_1223,In_4143);
xnor U1502 (N_1502,In_3122,In_524);
nor U1503 (N_1503,N_546,N_307);
nand U1504 (N_1504,In_3468,In_420);
and U1505 (N_1505,N_911,N_1341);
xor U1506 (N_1506,In_1953,In_539);
and U1507 (N_1507,N_296,N_684);
and U1508 (N_1508,In_2705,In_43);
and U1509 (N_1509,N_1354,In_3452);
or U1510 (N_1510,In_2127,In_2772);
or U1511 (N_1511,In_3585,N_1246);
xor U1512 (N_1512,N_907,In_1983);
and U1513 (N_1513,In_4293,In_3531);
nand U1514 (N_1514,In_1625,In_2221);
nor U1515 (N_1515,In_3646,N_1313);
nand U1516 (N_1516,In_142,N_1070);
or U1517 (N_1517,In_1397,N_1217);
nand U1518 (N_1518,In_288,In_1484);
xor U1519 (N_1519,In_3516,In_3473);
nor U1520 (N_1520,In_1092,In_2698);
xnor U1521 (N_1521,In_240,In_242);
or U1522 (N_1522,In_646,In_4066);
and U1523 (N_1523,N_1031,N_1286);
or U1524 (N_1524,In_4538,N_875);
nor U1525 (N_1525,N_964,In_197);
and U1526 (N_1526,N_1254,In_475);
nor U1527 (N_1527,N_982,N_1431);
and U1528 (N_1528,In_1168,In_531);
nand U1529 (N_1529,N_1032,In_2546);
or U1530 (N_1530,N_392,N_857);
xnor U1531 (N_1531,In_4097,In_3999);
nor U1532 (N_1532,In_1236,In_751);
nor U1533 (N_1533,In_2774,N_217);
nor U1534 (N_1534,N_278,In_1491);
nand U1535 (N_1535,N_746,In_588);
nand U1536 (N_1536,N_76,N_122);
nor U1537 (N_1537,N_260,N_1350);
nand U1538 (N_1538,In_1838,N_275);
or U1539 (N_1539,N_302,In_1624);
nand U1540 (N_1540,In_1507,In_1147);
nor U1541 (N_1541,In_4486,In_2826);
nand U1542 (N_1542,In_2796,N_1033);
or U1543 (N_1543,N_1058,In_1978);
and U1544 (N_1544,N_1376,In_2551);
xor U1545 (N_1545,In_565,N_197);
or U1546 (N_1546,In_1561,N_3);
or U1547 (N_1547,N_1370,N_171);
nand U1548 (N_1548,In_4586,In_875);
xor U1549 (N_1549,In_679,N_984);
nor U1550 (N_1550,In_4409,In_4111);
nor U1551 (N_1551,N_1165,N_1314);
nand U1552 (N_1552,In_4527,In_3522);
and U1553 (N_1553,N_1030,N_764);
nand U1554 (N_1554,In_2696,N_1000);
nor U1555 (N_1555,In_3384,N_1044);
or U1556 (N_1556,N_45,In_1975);
xor U1557 (N_1557,In_967,In_161);
nand U1558 (N_1558,In_4782,N_1240);
nand U1559 (N_1559,N_989,In_2389);
nand U1560 (N_1560,N_591,In_317);
nand U1561 (N_1561,N_999,In_4368);
nand U1562 (N_1562,In_4226,In_1859);
or U1563 (N_1563,In_3033,In_2747);
xor U1564 (N_1564,N_1282,In_1855);
xor U1565 (N_1565,In_2885,In_3675);
nand U1566 (N_1566,N_1392,N_213);
nand U1567 (N_1567,N_1328,N_625);
or U1568 (N_1568,N_290,In_27);
xor U1569 (N_1569,In_1772,In_3232);
xnor U1570 (N_1570,In_4006,In_1736);
nor U1571 (N_1571,N_331,In_1810);
or U1572 (N_1572,In_4341,In_1830);
or U1573 (N_1573,In_2485,In_2982);
and U1574 (N_1574,N_767,N_931);
nand U1575 (N_1575,N_206,In_4576);
nor U1576 (N_1576,In_1453,In_3537);
nor U1577 (N_1577,N_1320,In_904);
and U1578 (N_1578,N_1171,In_1285);
nor U1579 (N_1579,In_1197,In_587);
xnor U1580 (N_1580,In_4391,In_2370);
xnor U1581 (N_1581,N_1220,N_1372);
and U1582 (N_1582,N_309,In_249);
xnor U1583 (N_1583,In_4153,In_3171);
nand U1584 (N_1584,In_2567,In_4431);
xnor U1585 (N_1585,N_1197,In_4691);
or U1586 (N_1586,N_735,N_15);
and U1587 (N_1587,N_259,N_908);
and U1588 (N_1588,In_4884,N_65);
and U1589 (N_1589,In_1696,In_2359);
nor U1590 (N_1590,N_1479,In_120);
nand U1591 (N_1591,N_797,In_3430);
and U1592 (N_1592,N_328,N_713);
or U1593 (N_1593,In_2752,In_1429);
and U1594 (N_1594,N_1010,In_4752);
and U1595 (N_1595,N_380,N_43);
nor U1596 (N_1596,N_188,In_5);
or U1597 (N_1597,In_3024,N_720);
or U1598 (N_1598,N_1243,In_1303);
nor U1599 (N_1599,In_3873,In_2565);
xor U1600 (N_1600,In_1760,In_1946);
nor U1601 (N_1601,In_2954,In_3209);
or U1602 (N_1602,In_3142,In_4094);
xor U1603 (N_1603,In_1434,N_515);
nand U1604 (N_1604,N_899,In_1487);
nor U1605 (N_1605,N_1344,N_902);
nand U1606 (N_1606,N_1408,In_4355);
or U1607 (N_1607,N_598,N_1393);
and U1608 (N_1608,N_428,In_2814);
or U1609 (N_1609,In_4650,N_1463);
xor U1610 (N_1610,In_4938,In_1350);
and U1611 (N_1611,In_263,In_4108);
or U1612 (N_1612,N_169,In_172);
or U1613 (N_1613,In_48,In_1238);
nor U1614 (N_1614,In_74,In_1685);
nor U1615 (N_1615,In_3897,In_3257);
and U1616 (N_1616,In_3834,N_1374);
or U1617 (N_1617,In_403,In_1770);
nor U1618 (N_1618,In_4103,N_952);
and U1619 (N_1619,In_464,In_4751);
xor U1620 (N_1620,In_2230,In_3463);
or U1621 (N_1621,In_4651,N_695);
or U1622 (N_1622,N_417,In_3283);
and U1623 (N_1623,In_3989,In_4784);
or U1624 (N_1624,In_2416,In_1695);
and U1625 (N_1625,In_4298,In_204);
nand U1626 (N_1626,In_2330,In_4044);
and U1627 (N_1627,N_927,In_4671);
nor U1628 (N_1628,In_444,N_207);
and U1629 (N_1629,In_2196,In_2492);
nand U1630 (N_1630,In_2978,In_4489);
and U1631 (N_1631,In_4766,In_4755);
or U1632 (N_1632,N_111,In_2274);
nor U1633 (N_1633,N_208,N_1063);
xnor U1634 (N_1634,In_3051,In_2316);
nand U1635 (N_1635,N_1204,In_678);
nand U1636 (N_1636,N_1389,In_888);
nor U1637 (N_1637,N_1429,In_1650);
nand U1638 (N_1638,In_1311,In_2101);
or U1639 (N_1639,In_1679,In_3561);
and U1640 (N_1640,N_1385,N_562);
and U1641 (N_1641,In_238,In_970);
nand U1642 (N_1642,In_2712,In_799);
and U1643 (N_1643,N_1424,In_3826);
and U1644 (N_1644,N_1390,In_4487);
xor U1645 (N_1645,In_1806,In_3739);
xor U1646 (N_1646,N_484,In_3798);
nand U1647 (N_1647,N_482,N_378);
nor U1648 (N_1648,In_1047,N_674);
and U1649 (N_1649,In_3848,In_3276);
and U1650 (N_1650,In_3964,N_1416);
nor U1651 (N_1651,In_4411,In_2080);
nor U1652 (N_1652,In_1974,N_1296);
and U1653 (N_1653,N_823,In_2652);
or U1654 (N_1654,In_4061,In_1258);
or U1655 (N_1655,In_4247,N_125);
or U1656 (N_1656,N_1308,N_1443);
and U1657 (N_1657,In_1759,N_528);
or U1658 (N_1658,In_784,In_2926);
or U1659 (N_1659,In_724,In_76);
nor U1660 (N_1660,In_1820,N_1456);
nand U1661 (N_1661,N_79,In_622);
or U1662 (N_1662,In_701,In_3066);
or U1663 (N_1663,In_323,In_4617);
or U1664 (N_1664,In_574,In_552);
nand U1665 (N_1665,In_304,In_2381);
nor U1666 (N_1666,In_332,In_3717);
and U1667 (N_1667,In_3565,In_2740);
nor U1668 (N_1668,N_1109,In_1239);
and U1669 (N_1669,In_3799,In_4237);
and U1670 (N_1670,In_4463,N_1140);
and U1671 (N_1671,In_1378,In_1269);
or U1672 (N_1672,In_2262,In_3377);
nor U1673 (N_1673,In_353,In_2556);
nand U1674 (N_1674,In_921,In_1074);
xor U1675 (N_1675,N_210,In_2645);
nand U1676 (N_1676,In_637,In_321);
or U1677 (N_1677,In_2720,In_484);
and U1678 (N_1678,In_1052,N_330);
xnor U1679 (N_1679,In_656,N_1433);
xnor U1680 (N_1680,N_1325,In_3204);
or U1681 (N_1681,N_719,N_276);
and U1682 (N_1682,In_682,In_3957);
or U1683 (N_1683,In_4366,In_1522);
xnor U1684 (N_1684,In_390,In_1634);
and U1685 (N_1685,In_364,In_3100);
xor U1686 (N_1686,In_2323,N_1012);
nor U1687 (N_1687,N_227,In_4211);
nand U1688 (N_1688,In_777,In_3924);
or U1689 (N_1689,In_968,In_4090);
xor U1690 (N_1690,N_847,In_3341);
xnor U1691 (N_1691,N_636,In_4911);
nand U1692 (N_1692,N_1337,In_227);
xnor U1693 (N_1693,In_4146,N_1118);
or U1694 (N_1694,In_4581,In_1756);
and U1695 (N_1695,N_121,In_3650);
xor U1696 (N_1696,N_1400,In_367);
nand U1697 (N_1697,In_4683,In_2456);
nor U1698 (N_1698,In_4290,N_183);
nand U1699 (N_1699,In_3941,In_267);
or U1700 (N_1700,N_683,N_1052);
and U1701 (N_1701,In_4974,In_2727);
or U1702 (N_1702,In_3005,In_4663);
nor U1703 (N_1703,In_122,In_3499);
and U1704 (N_1704,In_1904,In_1789);
xnor U1705 (N_1705,In_901,In_1016);
or U1706 (N_1706,N_374,In_2342);
xor U1707 (N_1707,In_1056,In_399);
nor U1708 (N_1708,In_3922,N_825);
nand U1709 (N_1709,N_928,In_615);
and U1710 (N_1710,N_447,In_3987);
xor U1711 (N_1711,N_38,In_3478);
nand U1712 (N_1712,In_684,In_2644);
and U1713 (N_1713,In_1911,In_1706);
or U1714 (N_1714,In_56,N_1066);
nand U1715 (N_1715,N_469,In_1471);
or U1716 (N_1716,In_4201,N_766);
xor U1717 (N_1717,In_1722,In_2110);
nor U1718 (N_1718,In_3447,In_3256);
or U1719 (N_1719,In_4051,In_308);
or U1720 (N_1720,In_1172,N_21);
nand U1721 (N_1721,In_4027,In_3292);
nand U1722 (N_1722,N_917,In_1096);
nand U1723 (N_1723,N_565,In_494);
and U1724 (N_1724,In_4860,In_158);
nand U1725 (N_1725,N_1437,N_706);
xor U1726 (N_1726,In_847,N_533);
xor U1727 (N_1727,In_327,In_3010);
nor U1728 (N_1728,N_623,N_1316);
or U1729 (N_1729,N_1373,In_3442);
nand U1730 (N_1730,In_834,In_264);
or U1731 (N_1731,N_165,In_2998);
nor U1732 (N_1732,In_4898,N_814);
nor U1733 (N_1733,In_2501,In_1144);
xor U1734 (N_1734,In_598,In_2360);
xor U1735 (N_1735,In_2502,In_4874);
or U1736 (N_1736,N_916,In_2402);
or U1737 (N_1737,In_1697,In_1455);
nor U1738 (N_1738,N_805,N_406);
nor U1739 (N_1739,In_29,In_1423);
and U1740 (N_1740,N_212,N_1279);
or U1741 (N_1741,N_40,In_2507);
xnor U1742 (N_1742,N_1135,In_37);
xnor U1743 (N_1743,In_268,In_3628);
and U1744 (N_1744,N_442,In_2223);
xor U1745 (N_1745,In_4579,In_4316);
nor U1746 (N_1746,In_3606,N_1363);
nand U1747 (N_1747,In_1542,N_44);
nand U1748 (N_1748,In_1114,In_4392);
and U1749 (N_1749,N_1494,N_780);
or U1750 (N_1750,N_143,In_2660);
or U1751 (N_1751,In_994,In_2186);
nor U1752 (N_1752,N_878,In_3830);
nand U1753 (N_1753,In_1184,In_3686);
nand U1754 (N_1754,In_4354,N_1206);
and U1755 (N_1755,N_497,N_966);
and U1756 (N_1756,In_2951,In_4067);
xnor U1757 (N_1757,In_4809,N_1391);
nor U1758 (N_1758,In_621,In_1924);
or U1759 (N_1759,In_4917,In_4761);
nor U1760 (N_1760,In_1699,N_1594);
or U1761 (N_1761,N_1239,N_1547);
nand U1762 (N_1762,In_2834,In_1984);
nand U1763 (N_1763,N_1343,In_4036);
nor U1764 (N_1764,N_744,N_1426);
and U1765 (N_1765,In_4406,N_323);
or U1766 (N_1766,In_1553,In_2971);
xor U1767 (N_1767,In_2304,In_4588);
and U1768 (N_1768,N_315,N_1668);
and U1769 (N_1769,In_3477,N_241);
xor U1770 (N_1770,N_359,N_620);
nor U1771 (N_1771,N_1037,N_1445);
or U1772 (N_1772,N_321,In_2411);
nand U1773 (N_1773,In_4422,N_1235);
nand U1774 (N_1774,In_3391,In_2552);
and U1775 (N_1775,N_622,In_3737);
or U1776 (N_1776,In_1516,In_745);
xor U1777 (N_1777,In_237,In_2898);
xor U1778 (N_1778,In_1287,N_1491);
nand U1779 (N_1779,N_1459,N_772);
or U1780 (N_1780,In_2151,In_4556);
nand U1781 (N_1781,N_1511,N_1176);
xor U1782 (N_1782,N_1529,N_1434);
and U1783 (N_1783,In_291,N_1536);
or U1784 (N_1784,N_1048,In_2669);
nor U1785 (N_1785,In_2937,N_1546);
or U1786 (N_1786,N_1419,In_3996);
and U1787 (N_1787,In_4840,In_3782);
or U1788 (N_1788,In_154,In_1723);
and U1789 (N_1789,N_1233,In_4342);
xnor U1790 (N_1790,N_1597,N_1614);
nand U1791 (N_1791,In_3425,In_4870);
or U1792 (N_1792,N_1116,In_162);
and U1793 (N_1793,In_2062,N_1075);
nand U1794 (N_1794,In_4030,In_3720);
nor U1795 (N_1795,In_4658,In_3480);
nand U1796 (N_1796,N_1101,N_525);
nor U1797 (N_1797,N_1561,In_250);
nand U1798 (N_1798,In_4386,In_3639);
nor U1799 (N_1799,N_470,N_1086);
xnor U1800 (N_1800,N_349,In_512);
xor U1801 (N_1801,N_937,In_4546);
and U1802 (N_1802,N_153,In_3687);
and U1803 (N_1803,In_1379,In_1291);
nand U1804 (N_1804,In_4167,In_2732);
and U1805 (N_1805,In_557,N_1089);
xor U1806 (N_1806,In_53,N_283);
or U1807 (N_1807,In_4273,In_3045);
nand U1808 (N_1808,In_2918,N_1402);
xor U1809 (N_1809,In_1831,N_1381);
nand U1810 (N_1810,N_1652,In_4453);
nand U1811 (N_1811,N_1222,In_4594);
nor U1812 (N_1812,N_1015,In_89);
nor U1813 (N_1813,In_595,In_3962);
or U1814 (N_1814,In_1573,N_1563);
and U1815 (N_1815,In_3208,In_4532);
nor U1816 (N_1816,N_1074,In_4075);
xnor U1817 (N_1817,N_1427,In_4697);
nand U1818 (N_1818,N_1151,N_1380);
and U1819 (N_1819,In_188,N_672);
xor U1820 (N_1820,N_1020,In_4887);
or U1821 (N_1821,In_1212,N_957);
and U1822 (N_1822,In_2276,In_1960);
xor U1823 (N_1823,In_2029,N_1407);
xnor U1824 (N_1824,N_978,In_4054);
or U1825 (N_1825,N_871,In_984);
xnor U1826 (N_1826,In_1046,In_2904);
or U1827 (N_1827,N_138,In_3603);
nor U1828 (N_1828,In_2658,In_1802);
nor U1829 (N_1829,In_4986,N_1495);
and U1830 (N_1830,N_696,N_1411);
xnor U1831 (N_1831,In_2087,N_1142);
and U1832 (N_1832,In_3429,In_1065);
xnor U1833 (N_1833,In_4972,In_2715);
nand U1834 (N_1834,N_490,In_4009);
xor U1835 (N_1835,In_4021,N_1745);
nand U1836 (N_1836,N_1001,N_1535);
nand U1837 (N_1837,In_4231,N_1195);
nor U1838 (N_1838,N_327,N_157);
and U1839 (N_1839,In_2120,In_62);
nand U1840 (N_1840,N_1193,In_4148);
xor U1841 (N_1841,In_4627,In_558);
xor U1842 (N_1842,In_4890,N_700);
and U1843 (N_1843,In_1777,In_241);
nor U1844 (N_1844,In_919,N_285);
and U1845 (N_1845,In_4082,In_355);
nand U1846 (N_1846,N_107,N_754);
or U1847 (N_1847,In_2730,N_270);
nand U1848 (N_1848,N_1351,In_2436);
nand U1849 (N_1849,In_1115,In_3508);
xnor U1850 (N_1850,In_3582,In_406);
nand U1851 (N_1851,In_3139,In_861);
and U1852 (N_1852,N_1045,In_4229);
xor U1853 (N_1853,In_2831,In_73);
and U1854 (N_1854,N_284,In_3203);
or U1855 (N_1855,In_1533,In_4263);
and U1856 (N_1856,In_1822,N_1039);
or U1857 (N_1857,In_3776,In_2589);
and U1858 (N_1858,In_2294,In_4746);
and U1859 (N_1859,In_328,In_1662);
nor U1860 (N_1860,In_1824,N_1);
and U1861 (N_1861,N_317,N_1519);
xor U1862 (N_1862,In_4474,In_4023);
nand U1863 (N_1863,In_3698,In_2139);
xnor U1864 (N_1864,In_1376,N_1290);
nand U1865 (N_1865,N_1057,In_1118);
nand U1866 (N_1866,In_1796,In_3859);
or U1867 (N_1867,In_2604,In_1130);
nor U1868 (N_1868,N_939,In_4482);
or U1869 (N_1869,In_1085,N_369);
nor U1870 (N_1870,In_3879,In_4998);
nand U1871 (N_1871,N_996,N_360);
or U1872 (N_1872,In_4906,In_1103);
or U1873 (N_1873,N_732,N_659);
nand U1874 (N_1874,N_1317,In_3801);
nand U1875 (N_1875,In_1181,In_2560);
or U1876 (N_1876,In_1582,In_4897);
xnor U1877 (N_1877,In_4415,In_2717);
nand U1878 (N_1878,N_1178,N_218);
nor U1879 (N_1879,In_3684,N_736);
and U1880 (N_1880,In_2889,In_2923);
nand U1881 (N_1881,N_1356,In_3792);
nand U1882 (N_1882,N_1633,N_1613);
nor U1883 (N_1883,N_1683,N_773);
or U1884 (N_1884,In_2123,N_186);
nor U1885 (N_1885,In_28,In_2378);
nor U1886 (N_1886,In_2077,In_4868);
or U1887 (N_1887,N_1081,N_1345);
or U1888 (N_1888,In_3914,N_252);
xnor U1889 (N_1889,N_295,In_2050);
and U1890 (N_1890,In_4559,In_614);
xnor U1891 (N_1891,N_657,N_975);
nor U1892 (N_1892,N_77,In_4928);
nor U1893 (N_1893,N_751,N_382);
xnor U1894 (N_1894,In_4372,In_1167);
and U1895 (N_1895,In_36,N_1714);
and U1896 (N_1896,In_329,N_1441);
nand U1897 (N_1897,In_2487,In_4424);
nand U1898 (N_1898,In_3781,In_207);
xor U1899 (N_1899,In_1189,In_1579);
and U1900 (N_1900,In_447,In_1011);
xnor U1901 (N_1901,In_739,N_893);
nand U1902 (N_1902,In_438,N_532);
nor U1903 (N_1903,N_461,In_3201);
nand U1904 (N_1904,In_1267,N_1686);
and U1905 (N_1905,N_1601,In_206);
or U1906 (N_1906,N_1289,In_4777);
or U1907 (N_1907,In_2999,In_4923);
nand U1908 (N_1908,In_3199,In_2211);
nand U1909 (N_1909,In_3655,In_4501);
and U1910 (N_1910,In_962,In_2690);
nor U1911 (N_1911,In_3699,In_1701);
or U1912 (N_1912,In_2484,N_865);
nor U1913 (N_1913,N_1146,In_1568);
and U1914 (N_1914,In_1515,N_570);
and U1915 (N_1915,In_3094,N_495);
or U1916 (N_1916,N_1508,In_2415);
nor U1917 (N_1917,N_465,In_3027);
xnor U1918 (N_1918,In_2996,In_3557);
or U1919 (N_1919,In_1132,In_446);
xor U1920 (N_1920,In_1061,In_3123);
nor U1921 (N_1921,In_2046,N_810);
nor U1922 (N_1922,N_579,In_3379);
and U1923 (N_1923,In_1623,N_234);
nor U1924 (N_1924,N_1315,N_1700);
and U1925 (N_1925,In_3381,In_1863);
and U1926 (N_1926,In_673,In_964);
xor U1927 (N_1927,N_552,In_186);
and U1928 (N_1928,N_1100,N_432);
nand U1929 (N_1929,N_829,In_2867);
and U1930 (N_1930,In_3722,In_2268);
xor U1931 (N_1931,N_686,In_3305);
or U1932 (N_1932,N_1136,In_2298);
xnor U1933 (N_1933,In_4877,N_1552);
or U1934 (N_1934,N_868,N_1169);
nor U1935 (N_1935,N_1259,In_4088);
and U1936 (N_1936,N_100,N_962);
nand U1937 (N_1937,In_4168,In_458);
xnor U1938 (N_1938,In_2314,N_493);
and U1939 (N_1939,N_59,In_3119);
and U1940 (N_1940,In_4735,N_1092);
or U1941 (N_1941,N_718,N_542);
nand U1942 (N_1942,N_1046,In_2171);
or U1943 (N_1943,In_92,In_4566);
xor U1944 (N_1944,N_1016,N_832);
nor U1945 (N_1945,In_1449,In_4820);
nor U1946 (N_1946,N_1347,N_1080);
or U1947 (N_1947,N_1663,In_2603);
xnor U1948 (N_1948,In_2011,N_367);
nand U1949 (N_1949,N_664,N_1166);
nor U1950 (N_1950,N_225,N_1466);
and U1951 (N_1951,N_366,In_4609);
or U1952 (N_1952,N_529,In_54);
nand U1953 (N_1953,N_1256,In_1652);
and U1954 (N_1954,N_855,In_483);
xnor U1955 (N_1955,N_1106,In_2818);
or U1956 (N_1956,N_817,In_231);
or U1957 (N_1957,In_469,In_4176);
and U1958 (N_1958,In_3855,In_1254);
nand U1959 (N_1959,In_4533,N_1742);
xor U1960 (N_1960,In_4981,In_941);
nor U1961 (N_1961,N_475,In_929);
and U1962 (N_1962,In_2100,In_160);
nor U1963 (N_1963,In_2277,N_694);
nand U1964 (N_1964,N_1608,In_3357);
or U1965 (N_1965,In_3544,In_3396);
nand U1966 (N_1966,N_191,In_3264);
or U1967 (N_1967,N_1602,N_1504);
nor U1968 (N_1968,N_556,In_1778);
or U1969 (N_1969,N_27,N_342);
nor U1970 (N_1970,N_1236,In_2060);
and U1971 (N_1971,In_4190,In_4029);
xnor U1972 (N_1972,N_898,In_4173);
nand U1973 (N_1973,In_704,N_1694);
xor U1974 (N_1974,N_1005,In_4622);
and U1975 (N_1975,In_4555,N_1025);
and U1976 (N_1976,In_1049,In_4384);
xor U1977 (N_1977,N_1452,In_2183);
or U1978 (N_1978,In_246,In_4272);
nand U1979 (N_1979,In_768,In_1271);
nand U1980 (N_1980,N_1104,In_1309);
nand U1981 (N_1981,In_4223,In_3809);
nand U1982 (N_1982,N_1549,N_1368);
nor U1983 (N_1983,In_2624,In_2986);
xnor U1984 (N_1984,In_4540,In_3163);
nor U1985 (N_1985,In_2093,In_3004);
or U1986 (N_1986,N_1626,N_1425);
xnor U1987 (N_1987,In_363,N_1702);
and U1988 (N_1988,In_4401,N_253);
or U1989 (N_1989,In_661,N_1177);
and U1990 (N_1990,In_4043,In_4046);
nor U1991 (N_1991,In_710,N_1119);
nor U1992 (N_1992,In_2798,In_3788);
nor U1993 (N_1993,N_1387,In_1647);
or U1994 (N_1994,In_255,In_4639);
and U1995 (N_1995,N_1014,In_3245);
xnor U1996 (N_1996,In_3434,In_343);
xnor U1997 (N_1997,N_1467,N_156);
or U1998 (N_1998,In_4179,In_86);
nor U1999 (N_1999,In_1860,In_2617);
nor U2000 (N_2000,N_1923,N_1454);
or U2001 (N_2001,In_2000,In_1733);
nand U2002 (N_2002,In_4468,N_1201);
nand U2003 (N_2003,In_1559,In_691);
or U2004 (N_2004,In_358,In_1337);
nor U2005 (N_2005,In_4721,In_283);
xor U2006 (N_2006,N_1500,In_4107);
or U2007 (N_2007,In_3678,N_272);
nand U2008 (N_2008,In_714,N_703);
xnor U2009 (N_2009,N_1658,In_4250);
nor U2010 (N_2010,In_1753,N_1267);
nand U2011 (N_2011,In_1344,In_2092);
nand U2012 (N_2012,In_2005,In_1426);
xnor U2013 (N_2013,N_291,In_4150);
and U2014 (N_2014,In_1614,In_3682);
and U2015 (N_2015,N_1278,In_2879);
and U2016 (N_2016,N_1641,In_2557);
xor U2017 (N_2017,In_1323,In_4592);
nor U2018 (N_2018,In_4846,In_1762);
nor U2019 (N_2019,N_1567,N_849);
xnor U2020 (N_2020,In_3597,In_3277);
and U2021 (N_2021,In_1712,In_1509);
or U2022 (N_2022,N_1468,N_1133);
xnor U2023 (N_2023,N_1497,N_1348);
nand U2024 (N_2024,N_1327,N_1023);
nor U2025 (N_2025,N_1484,N_1576);
xor U2026 (N_2026,N_1183,N_1853);
xor U2027 (N_2027,N_142,N_1329);
or U2028 (N_2028,N_1338,In_443);
or U2029 (N_2029,In_928,In_992);
nor U2030 (N_2030,N_762,In_680);
nand U2031 (N_2031,In_4215,In_2319);
nand U2032 (N_2032,In_1948,In_2010);
and U2033 (N_2033,In_4595,In_4672);
xor U2034 (N_2034,N_841,In_371);
nor U2035 (N_2035,In_668,N_1907);
nor U2036 (N_2036,In_4238,N_950);
nand U2037 (N_2037,N_1762,In_2634);
nor U2038 (N_2038,In_314,In_2418);
or U2039 (N_2039,N_71,In_1266);
nand U2040 (N_2040,N_1172,N_770);
nand U2041 (N_2041,In_1106,In_2135);
or U2042 (N_2042,In_3590,In_381);
xor U2043 (N_2043,N_416,N_1170);
nand U2044 (N_2044,In_2615,N_885);
or U2045 (N_2045,In_2681,In_3311);
nand U2046 (N_2046,In_3822,N_1026);
nor U2047 (N_2047,In_2401,In_2743);
xor U2048 (N_2048,N_1417,In_1459);
xor U2049 (N_2049,In_1203,In_1213);
nor U2050 (N_2050,In_4632,N_60);
or U2051 (N_2051,In_4346,In_2886);
or U2052 (N_2052,N_1530,In_3790);
nor U2053 (N_2053,In_58,In_3419);
nand U2054 (N_2054,In_2722,In_2952);
and U2055 (N_2055,N_510,In_294);
or U2056 (N_2056,In_319,N_1245);
or U2057 (N_2057,N_569,N_1738);
nand U2058 (N_2058,N_453,N_1531);
and U2059 (N_2059,In_4847,In_1069);
and U2060 (N_2060,In_4122,N_1418);
or U2061 (N_2061,In_3187,In_1441);
and U2062 (N_2062,In_2504,In_4562);
nor U2063 (N_2063,In_1763,In_4844);
or U2064 (N_2064,In_2243,In_3575);
and U2065 (N_2065,N_1506,N_1436);
nor U2066 (N_2066,In_4281,In_4504);
xor U2067 (N_2067,In_2496,In_311);
nor U2068 (N_2068,In_1918,In_2911);
xor U2069 (N_2069,In_3581,N_280);
nand U2070 (N_2070,N_903,N_687);
nand U2071 (N_2071,N_1073,In_3849);
xnor U2072 (N_2072,In_4507,N_1986);
xnor U2073 (N_2073,N_1792,In_1038);
nor U2074 (N_2074,In_2596,N_279);
or U2075 (N_2075,In_3819,N_756);
nor U2076 (N_2076,In_2020,N_1977);
nor U2077 (N_2077,N_1695,N_1573);
and U2078 (N_2078,N_1285,N_1743);
and U2079 (N_2079,In_708,In_3929);
xnor U2080 (N_2080,N_985,In_1176);
or U2081 (N_2081,In_3361,N_1649);
or U2082 (N_2082,N_2,N_1098);
and U2083 (N_2083,N_972,N_51);
and U2084 (N_2084,N_1874,In_4420);
or U2085 (N_2085,N_1963,N_304);
or U2086 (N_2086,In_2386,N_1301);
and U2087 (N_2087,N_1998,In_4764);
xor U2088 (N_2088,N_1252,In_4074);
nand U2089 (N_2089,N_1298,N_1718);
or U2090 (N_2090,N_1273,N_946);
nor U2091 (N_2091,N_1514,In_1028);
xor U2092 (N_2092,In_3871,N_1330);
or U2093 (N_2093,N_161,In_3719);
and U2094 (N_2094,In_2844,In_4348);
and U2095 (N_2095,In_4514,In_2976);
and U2096 (N_2096,N_1238,In_898);
or U2097 (N_2097,N_729,In_3448);
and U2098 (N_2098,In_305,N_581);
or U2099 (N_2099,In_4873,In_610);
and U2100 (N_2100,In_417,N_611);
nand U2101 (N_2101,In_2689,In_4033);
or U2102 (N_2102,In_1524,In_733);
nor U2103 (N_2103,In_4711,In_216);
or U2104 (N_2104,N_1192,In_1751);
and U2105 (N_2105,N_1938,N_1910);
xnor U2106 (N_2106,N_559,N_209);
or U2107 (N_2107,N_519,N_851);
and U2108 (N_2108,In_384,N_1890);
xor U2109 (N_2109,N_789,N_1518);
and U2110 (N_2110,In_2320,N_1229);
nor U2111 (N_2111,N_1661,In_1782);
and U2112 (N_2112,N_42,In_2313);
or U2113 (N_2113,N_423,In_1138);
xor U2114 (N_2114,In_4320,N_1332);
or U2115 (N_2115,In_4344,N_373);
or U2116 (N_2116,In_864,N_1930);
nand U2117 (N_2117,N_383,In_1324);
xor U2118 (N_2118,N_601,In_912);
nor U2119 (N_2119,N_1640,In_333);
xor U2120 (N_2120,N_258,N_1637);
nand U2121 (N_2121,N_254,In_1848);
nor U2122 (N_2122,In_4510,N_1553);
and U2123 (N_2123,In_894,N_986);
and U2124 (N_2124,In_3894,In_1113);
nor U2125 (N_2125,In_568,N_1969);
xnor U2126 (N_2126,In_4509,N_1842);
or U2127 (N_2127,In_4867,N_1571);
xor U2128 (N_2128,N_1199,In_2041);
xor U2129 (N_2129,In_3095,In_2862);
nor U2130 (N_2130,In_806,N_1420);
xnor U2131 (N_2131,In_354,N_1481);
or U2132 (N_2132,In_301,In_2605);
and U2133 (N_2133,In_292,In_3856);
nor U2134 (N_2134,N_650,N_1295);
nand U2135 (N_2135,N_880,In_1940);
or U2136 (N_2136,In_2621,In_2746);
nor U2137 (N_2137,In_4236,In_2384);
and U2138 (N_2138,N_884,In_3839);
nor U2139 (N_2139,N_1648,In_4646);
xnor U2140 (N_2140,In_2379,In_3627);
or U2141 (N_2141,In_3210,In_3156);
nor U2142 (N_2142,N_1731,N_1579);
nor U2143 (N_2143,N_644,N_167);
or U2144 (N_2144,N_1947,N_1292);
or U2145 (N_2145,N_924,In_4934);
and U2146 (N_2146,N_481,In_3588);
xor U2147 (N_2147,In_908,N_1784);
nor U2148 (N_2148,In_1234,N_1855);
and U2149 (N_2149,N_1616,In_3184);
and U2150 (N_2150,N_1360,N_1617);
or U2151 (N_2151,In_2518,N_75);
and U2152 (N_2152,N_1059,In_1923);
nor U2153 (N_2153,In_1817,N_1786);
nor U2154 (N_2154,N_1898,In_3658);
nor U2155 (N_2155,In_583,N_1944);
and U2156 (N_2156,In_4104,In_3714);
xnor U2157 (N_2157,N_1397,N_1167);
nand U2158 (N_2158,In_4447,N_1526);
or U2159 (N_2159,In_2096,N_1158);
xor U2160 (N_2160,In_2865,N_1022);
xnor U2161 (N_2161,In_350,In_208);
nor U2162 (N_2162,In_3732,N_1876);
xnor U2163 (N_2163,In_1622,In_560);
xnor U2164 (N_2164,N_1713,In_3709);
and U2165 (N_2165,N_584,In_3904);
xor U2166 (N_2166,In_1161,N_800);
nor U2167 (N_2167,N_1095,N_1837);
and U2168 (N_2168,N_1386,N_224);
nor U2169 (N_2169,In_4057,In_1137);
xor U2170 (N_2170,In_2054,N_1639);
and U2171 (N_2171,In_2990,N_1496);
xnor U2172 (N_2172,In_902,N_93);
nand U2173 (N_2173,In_3335,In_1764);
or U2174 (N_2174,N_615,In_4539);
nand U2175 (N_2175,N_1523,N_269);
and U2176 (N_2176,In_4723,In_4824);
xnor U2177 (N_2177,N_1153,In_322);
or U2178 (N_2178,In_1499,N_1283);
nor U2179 (N_2179,In_2676,N_1843);
and U2180 (N_2180,In_4991,In_4816);
or U2181 (N_2181,N_1928,N_1924);
or U2182 (N_2182,In_1411,In_2900);
and U2183 (N_2183,In_4644,N_1715);
and U2184 (N_2184,N_1265,N_1804);
nor U2185 (N_2185,In_3278,In_980);
nor U2186 (N_2186,N_1864,N_1091);
nand U2187 (N_2187,N_1395,In_1720);
or U2188 (N_2188,In_3467,In_3427);
nand U2189 (N_2189,In_4659,In_2654);
xnor U2190 (N_2190,N_1179,N_1905);
and U2191 (N_2191,In_1465,In_3300);
and U2192 (N_2192,In_2758,In_4526);
nor U2193 (N_2193,In_2896,In_3947);
nand U2194 (N_2194,In_1076,In_49);
nor U2195 (N_2195,In_1829,In_1895);
and U2196 (N_2196,In_1884,In_2609);
nand U2197 (N_2197,In_4857,In_4295);
nor U2198 (N_2198,N_333,N_24);
nor U2199 (N_2199,N_175,In_4827);
xnor U2200 (N_2200,N_670,N_1809);
and U2201 (N_2201,N_1994,In_4114);
nand U2202 (N_2202,In_4879,N_543);
and U2203 (N_2203,In_2959,In_4187);
and U2204 (N_2204,In_924,N_201);
or U2205 (N_2205,In_1126,In_802);
nor U2206 (N_2206,In_4369,In_1477);
nand U2207 (N_2207,In_1727,N_1747);
nor U2208 (N_2208,N_1302,N_1974);
xor U2209 (N_2209,In_2094,In_977);
xor U2210 (N_2210,In_4449,N_1666);
and U2211 (N_2211,In_1869,In_128);
or U2212 (N_2212,N_1968,N_912);
or U2213 (N_2213,N_921,In_3236);
or U2214 (N_2214,In_165,In_3751);
and U2215 (N_2215,In_474,N_1664);
xnor U2216 (N_2216,N_1995,In_103);
nor U2217 (N_2217,In_1157,In_4243);
nor U2218 (N_2218,In_3149,N_182);
and U2219 (N_2219,In_1659,N_1852);
and U2220 (N_2220,In_2534,In_4241);
and U2221 (N_2221,In_1095,N_56);
xnor U2222 (N_2222,N_775,In_787);
xnor U2223 (N_2223,In_3105,In_1292);
and U2224 (N_2224,N_1849,In_3389);
xnor U2225 (N_2225,N_1940,N_247);
nor U2226 (N_2226,N_983,N_388);
nor U2227 (N_2227,In_1547,N_1055);
xor U2228 (N_2228,In_4278,In_4305);
nor U2229 (N_2229,In_3461,N_1667);
xnor U2230 (N_2230,N_1965,N_1446);
xnor U2231 (N_2231,N_749,N_776);
nand U2232 (N_2232,In_2258,In_4019);
nand U2233 (N_2233,In_1275,N_1194);
and U2234 (N_2234,In_1470,N_1857);
or U2235 (N_2235,N_1807,In_1389);
or U2236 (N_2236,In_272,In_2519);
xnor U2237 (N_2237,N_1440,In_3214);
nor U2238 (N_2238,N_1801,N_740);
xor U2239 (N_2239,In_4361,In_1446);
xnor U2240 (N_2240,In_2176,N_1188);
or U2241 (N_2241,N_145,In_1141);
nand U2242 (N_2242,In_4428,In_3491);
nand U2243 (N_2243,In_2066,N_1544);
or U2244 (N_2244,In_1538,N_1087);
or U2245 (N_2245,N_697,In_2665);
xor U2246 (N_2246,N_242,N_774);
nor U2247 (N_2247,In_4331,In_2642);
nor U2248 (N_2248,N_177,In_3605);
xor U2249 (N_2249,In_1214,N_1765);
xor U2250 (N_2250,In_3398,N_1357);
xor U2251 (N_2251,In_3685,N_1478);
nor U2252 (N_2252,In_4569,N_1226);
nor U2253 (N_2253,In_3958,N_2205);
xnor U2254 (N_2254,In_1619,In_835);
and U2255 (N_2255,In_2435,N_1469);
nand U2256 (N_2256,N_11,In_2566);
xnor U2257 (N_2257,In_2682,In_4927);
nand U2258 (N_2258,In_2217,In_3619);
and U2259 (N_2259,In_1526,In_3812);
nand U2260 (N_2260,In_96,N_2173);
nor U2261 (N_2261,In_4969,In_2048);
and U2262 (N_2262,In_2843,In_3331);
nor U2263 (N_2263,N_1097,In_189);
xor U2264 (N_2264,N_1779,N_782);
nor U2265 (N_2265,In_3287,N_944);
or U2266 (N_2266,In_2515,N_1219);
nand U2267 (N_2267,In_2675,In_2115);
nor U2268 (N_2268,In_1784,In_400);
nor U2269 (N_2269,In_2813,In_1920);
xnor U2270 (N_2270,In_4152,In_2544);
xor U2271 (N_2271,In_541,In_3926);
xnor U2272 (N_2272,In_2697,N_2094);
xor U2273 (N_2273,In_3518,In_2053);
nand U2274 (N_2274,N_2039,N_1967);
nor U2275 (N_2275,N_1934,N_640);
and U2276 (N_2276,N_1921,In_4400);
nor U2277 (N_2277,N_646,N_1946);
nand U2278 (N_2278,N_1486,In_4524);
nor U2279 (N_2279,N_2121,In_3783);
nand U2280 (N_2280,N_1775,In_932);
nand U2281 (N_2281,In_1185,In_3176);
xnor U2282 (N_2282,N_1560,N_2105);
xor U2283 (N_2283,In_3,N_1076);
and U2284 (N_2284,In_4182,N_437);
xnor U2285 (N_2285,In_348,N_1846);
nor U2286 (N_2286,N_617,In_3820);
nor U2287 (N_2287,In_3555,N_2136);
or U2288 (N_2288,N_2059,In_1936);
or U2289 (N_2289,In_482,N_1629);
or U2290 (N_2290,In_4662,In_1282);
or U2291 (N_2291,In_3656,N_1502);
nor U2292 (N_2292,In_4068,N_788);
or U2293 (N_2293,N_990,In_3878);
or U2294 (N_2294,N_1232,N_1093);
and U2295 (N_2295,In_4931,In_2499);
xnor U2296 (N_2296,N_1945,In_4491);
and U2297 (N_2297,In_1560,In_3616);
nand U2298 (N_2298,N_202,N_385);
xnor U2299 (N_2299,In_3651,In_1355);
nand U2300 (N_2300,N_1028,In_2522);
and U2301 (N_2301,N_932,N_1671);
and U2302 (N_2302,In_3542,N_1489);
nand U2303 (N_2303,N_1979,In_1583);
xnor U2304 (N_2304,In_3460,In_3723);
xnor U2305 (N_2305,N_1124,N_1704);
xnor U2306 (N_2306,In_523,N_1077);
xnor U2307 (N_2307,In_647,In_4266);
xor U2308 (N_2308,In_2398,In_2664);
or U2309 (N_2309,In_3238,In_4599);
and U2310 (N_2310,In_3107,In_4593);
xor U2311 (N_2311,In_2400,N_1729);
nor U2312 (N_2312,N_1352,In_2922);
xor U2313 (N_2313,In_3076,In_1596);
or U2314 (N_2314,In_3747,N_856);
nor U2315 (N_2315,N_1677,N_673);
nand U2316 (N_2316,N_1827,In_3549);
xor U2317 (N_2317,In_3899,In_1857);
nor U2318 (N_2318,In_4209,In_1158);
or U2319 (N_2319,In_2975,In_997);
nor U2320 (N_2320,In_1591,N_2082);
xnor U2321 (N_2321,In_3694,In_1111);
or U2322 (N_2322,N_20,In_3242);
xnor U2323 (N_2323,N_1312,In_111);
and U2324 (N_2324,N_2244,N_149);
and U2325 (N_2325,N_1604,N_747);
xnor U2326 (N_2326,In_4105,N_1464);
xor U2327 (N_2327,In_887,In_4939);
nor U2328 (N_2328,In_3350,In_3791);
nand U2329 (N_2329,N_2087,N_1674);
and U2330 (N_2330,In_3960,N_402);
nor U2331 (N_2331,N_314,N_653);
xnor U2332 (N_2332,N_1379,N_1654);
xor U2333 (N_2333,N_1237,In_2072);
nor U2334 (N_2334,N_459,In_4171);
xnor U2335 (N_2335,In_1809,In_855);
nand U2336 (N_2336,In_3129,In_3229);
or U2337 (N_2337,N_685,In_2963);
nor U2338 (N_2338,N_384,In_1957);
nor U2339 (N_2339,N_712,N_1660);
nor U2340 (N_2340,N_1324,N_1125);
nor U2341 (N_2341,N_824,In_628);
nor U2342 (N_2342,N_1862,In_2950);
nor U2343 (N_2343,In_3725,In_3807);
and U2344 (N_2344,N_1018,In_1746);
xnor U2345 (N_2345,N_2152,In_2476);
nand U2346 (N_2346,In_3547,In_4749);
or U2347 (N_2347,In_1385,In_3034);
or U2348 (N_2348,N_795,In_4637);
xor U2349 (N_2349,N_1721,N_1241);
and U2350 (N_2350,N_1642,N_1471);
or U2351 (N_2351,N_1605,N_1904);
nand U2352 (N_2352,In_1245,N_1108);
nor U2353 (N_2353,In_2787,N_1681);
xor U2354 (N_2354,In_2679,N_1004);
xnor U2355 (N_2355,N_862,N_662);
and U2356 (N_2356,In_2859,N_1528);
xnor U2357 (N_2357,N_709,In_4980);
nand U2358 (N_2358,In_1592,In_578);
nor U2359 (N_2359,N_1072,N_1367);
nand U2360 (N_2360,N_2103,N_904);
nor U2361 (N_2361,In_4573,N_1207);
nand U2362 (N_2362,N_251,In_1327);
or U2363 (N_2363,In_1415,In_3017);
xor U2364 (N_2364,In_2493,N_1250);
nand U2365 (N_2365,In_3475,In_886);
or U2366 (N_2366,N_381,In_635);
xnor U2367 (N_2367,N_1079,N_1688);
nand U2368 (N_2368,In_2112,N_1992);
or U2369 (N_2369,In_3570,N_1186);
nor U2370 (N_2370,In_1467,N_325);
nand U2371 (N_2371,In_256,In_3681);
nand U2372 (N_2372,In_2317,In_3956);
or U2373 (N_2373,N_2091,In_4861);
nor U2374 (N_2374,N_1834,N_1817);
nor U2375 (N_2375,In_658,In_1620);
nor U2376 (N_2376,N_1808,N_2016);
or U2377 (N_2377,In_4390,N_1656);
nor U2378 (N_2378,N_1556,N_1949);
or U2379 (N_2379,In_4141,N_1720);
and U2380 (N_2380,N_2145,In_1402);
nor U2381 (N_2381,N_2068,In_4408);
and U2382 (N_2382,N_2146,In_1489);
nor U2383 (N_2383,N_2116,In_1846);
nor U2384 (N_2384,In_2403,In_4889);
or U2385 (N_2385,N_1515,In_4492);
nand U2386 (N_2386,N_357,In_2284);
and U2387 (N_2387,N_1691,N_2164);
or U2388 (N_2388,In_335,N_1692);
nor U2389 (N_2389,In_387,In_1988);
and U2390 (N_2390,N_655,In_126);
xnor U2391 (N_2391,N_1148,N_1631);
nor U2392 (N_2392,N_2003,In_1536);
nor U2393 (N_2393,N_1662,In_3578);
and U2394 (N_2394,In_3693,N_820);
xor U2395 (N_2395,In_4162,N_2010);
xor U2396 (N_2396,In_826,N_1507);
xnor U2397 (N_2397,N_1261,N_2129);
xnor U2398 (N_2398,In_4180,In_426);
xor U2399 (N_2399,In_2960,In_2180);
nand U2400 (N_2400,In_944,In_2771);
and U2401 (N_2401,In_2227,N_1791);
or U2402 (N_2402,N_861,In_943);
nor U2403 (N_2403,In_3466,N_1568);
xnor U2404 (N_2404,In_723,In_2282);
nand U2405 (N_2405,N_1823,In_271);
or U2406 (N_2406,N_596,In_2949);
nor U2407 (N_2407,In_378,In_2782);
or U2408 (N_2408,N_965,In_4966);
and U2409 (N_2409,In_88,In_3919);
xor U2410 (N_2410,N_1421,In_4621);
nand U2411 (N_2411,N_2018,N_460);
xnor U2412 (N_2412,N_691,In_1206);
xor U2413 (N_2413,N_1595,In_3059);
nor U2414 (N_2414,N_1274,N_1919);
xor U2415 (N_2415,In_1237,N_329);
nor U2416 (N_2416,In_1064,In_712);
and U2417 (N_2417,In_4488,N_743);
nor U2418 (N_2418,N_1740,N_2017);
nand U2419 (N_2419,In_221,N_1970);
and U2420 (N_2420,In_259,In_2671);
and U2421 (N_2421,In_1249,In_2590);
nor U2422 (N_2422,In_3223,In_1866);
xnor U2423 (N_2423,In_1490,N_2229);
nor U2424 (N_2424,N_1679,N_1462);
nor U2425 (N_2425,In_4794,In_1907);
nor U2426 (N_2426,N_1475,In_4603);
and U2427 (N_2427,N_2156,N_2077);
or U2428 (N_2428,In_4245,In_530);
and U2429 (N_2429,In_3810,In_1902);
xnor U2430 (N_2430,In_1550,In_1684);
and U2431 (N_2431,In_4505,N_1996);
nor U2432 (N_2432,N_1916,N_1620);
and U2433 (N_2433,In_1613,In_4315);
xor U2434 (N_2434,N_1512,In_3631);
or U2435 (N_2435,N_2166,N_2246);
and U2436 (N_2436,In_184,N_498);
xor U2437 (N_2437,N_1772,N_1493);
nor U2438 (N_2438,In_1139,N_1593);
nor U2439 (N_2439,In_2374,In_3030);
or U2440 (N_2440,N_1266,In_961);
and U2441 (N_2441,In_107,N_2028);
and U2442 (N_2442,N_1366,N_2047);
xor U2443 (N_2443,N_1006,In_3705);
or U2444 (N_2444,N_1612,In_3428);
and U2445 (N_2445,N_629,In_3444);
nor U2446 (N_2446,N_2199,N_1918);
nand U2447 (N_2447,In_2872,N_28);
xor U2448 (N_2448,In_623,N_2153);
xnor U2449 (N_2449,In_4970,In_1729);
nand U2450 (N_2450,In_357,In_4676);
xnor U2451 (N_2451,In_124,In_1349);
or U2452 (N_2452,In_252,N_2073);
xnor U2453 (N_2453,In_3704,N_1589);
nand U2454 (N_2454,In_1145,N_1861);
or U2455 (N_2455,In_843,In_1765);
nor U2456 (N_2456,N_1942,In_3775);
xor U2457 (N_2457,N_1956,N_1187);
or U2458 (N_2458,In_2577,N_1403);
and U2459 (N_2459,In_334,In_1544);
or U2460 (N_2460,N_1659,N_462);
and U2461 (N_2461,In_2861,In_106);
nor U2462 (N_2462,In_1207,In_3997);
or U2463 (N_2463,N_1856,In_2440);
and U2464 (N_2464,In_3596,In_4314);
xnor U2465 (N_2465,In_133,In_2708);
and U2466 (N_2466,In_1406,N_1796);
nand U2467 (N_2467,In_2891,N_1802);
nand U2468 (N_2468,In_3200,N_1488);
or U2469 (N_2469,In_897,N_1983);
or U2470 (N_2470,N_47,N_1287);
or U2471 (N_2471,In_4822,N_1094);
nand U2472 (N_2472,N_1414,N_1908);
nand U2473 (N_2473,N_2151,In_3902);
nand U2474 (N_2474,In_1199,N_2167);
nor U2475 (N_2475,N_2192,In_3117);
xor U2476 (N_2476,In_4297,In_4255);
and U2477 (N_2477,In_214,N_1734);
or U2478 (N_2478,N_1726,N_320);
xor U2479 (N_2479,In_4471,N_2114);
or U2480 (N_2480,In_2328,N_297);
nand U2481 (N_2481,N_2025,In_2273);
nor U2482 (N_2482,N_979,N_2074);
and U2483 (N_2483,In_1797,N_2212);
nand U2484 (N_2484,N_2030,N_499);
nor U2485 (N_2485,N_557,N_605);
nor U2486 (N_2486,In_2657,N_941);
and U2487 (N_2487,N_785,In_3530);
nor U2488 (N_2488,In_4393,N_1154);
xnor U2489 (N_2489,N_1735,In_3507);
nor U2490 (N_2490,N_473,N_1625);
nor U2491 (N_2491,N_956,In_4904);
nand U2492 (N_2492,In_1108,N_639);
or U2493 (N_2493,In_3572,In_2162);
nor U2494 (N_2494,In_397,N_925);
or U2495 (N_2495,N_516,N_219);
or U2496 (N_2496,In_97,In_1495);
xnor U2497 (N_2497,In_1818,N_1732);
or U2498 (N_2498,In_3977,In_290);
nor U2499 (N_2499,N_1878,In_4080);
nand U2500 (N_2500,N_845,In_4381);
or U2501 (N_2501,In_341,In_3622);
or U2502 (N_2502,N_1585,In_145);
nor U2503 (N_2503,In_1390,In_3872);
and U2504 (N_2504,In_4883,In_4515);
or U2505 (N_2505,N_906,N_478);
and U2506 (N_2506,In_4193,N_1689);
and U2507 (N_2507,N_981,N_681);
nand U2508 (N_2508,In_4324,In_485);
nor U2509 (N_2509,In_3743,N_807);
xnor U2510 (N_2510,In_4859,N_1888);
nand U2511 (N_2511,N_236,N_545);
xnor U2512 (N_2512,N_2429,In_1504);
nand U2513 (N_2513,N_97,In_1603);
and U2514 (N_2514,In_2741,In_4322);
nor U2515 (N_2515,N_991,N_448);
nand U2516 (N_2516,N_2348,N_1954);
or U2517 (N_2517,N_1042,In_4896);
nand U2518 (N_2518,In_1728,In_2074);
nor U2519 (N_2519,N_1300,N_1388);
xor U2520 (N_2520,N_1150,In_2133);
nand U2521 (N_2521,In_1281,N_1244);
nand U2522 (N_2522,In_4302,In_4472);
xnor U2523 (N_2523,N_2014,In_4442);
or U2524 (N_2524,N_920,In_4772);
and U2525 (N_2525,N_2482,In_1850);
or U2526 (N_2526,N_2428,In_4310);
or U2527 (N_2527,In_1969,N_2194);
and U2528 (N_2528,In_3390,N_1650);
and U2529 (N_2529,In_1364,N_2215);
and U2530 (N_2530,N_1242,In_1917);
nor U2531 (N_2531,N_1448,N_1705);
xor U2532 (N_2532,In_2090,N_1961);
xor U2533 (N_2533,In_2919,N_1914);
or U2534 (N_2534,In_2475,N_2271);
nor U2535 (N_2535,In_1068,N_2230);
nand U2536 (N_2536,N_1727,N_968);
nand U2537 (N_2537,In_2241,N_2457);
and U2538 (N_2538,In_1501,N_1845);
nor U2539 (N_2539,N_1430,In_4208);
nand U2540 (N_2540,In_931,In_257);
or U2541 (N_2541,In_3875,N_1582);
or U2542 (N_2542,In_4184,In_4199);
xnor U2543 (N_2543,In_3079,In_3916);
nor U2544 (N_2544,N_494,In_4729);
nand U2545 (N_2545,In_1567,In_2607);
or U2546 (N_2546,N_1682,In_3945);
or U2547 (N_2547,In_2994,N_2499);
nor U2548 (N_2548,In_1331,N_1234);
nand U2549 (N_2549,In_3268,In_620);
nor U2550 (N_2550,N_901,In_3857);
nand U2551 (N_2551,In_4875,N_1264);
nor U2552 (N_2552,N_860,In_1834);
or U2553 (N_2553,N_838,N_1404);
nand U2554 (N_2554,N_179,N_652);
or U2555 (N_2555,N_1865,In_85);
and U2556 (N_2556,In_581,N_1971);
or U2557 (N_2557,N_2162,In_108);
and U2558 (N_2558,In_2811,In_4977);
nand U2559 (N_2559,N_1707,In_1781);
and U2560 (N_2560,In_1427,N_2132);
nor U2561 (N_2561,N_1147,In_1480);
nor U2562 (N_2562,N_1262,In_4714);
xnor U2563 (N_2563,N_1800,In_3744);
or U2564 (N_2564,In_972,N_2339);
xnor U2565 (N_2565,N_1299,N_2040);
nor U2566 (N_2566,N_1570,In_4656);
nand U2567 (N_2567,N_1564,In_2734);
xnor U2568 (N_2568,N_1205,N_1019);
or U2569 (N_2569,N_1221,N_2083);
nor U2570 (N_2570,N_1889,N_2004);
nand U2571 (N_2571,In_2824,N_2005);
xor U2572 (N_2572,In_1646,N_1029);
and U2573 (N_2573,N_2384,N_1575);
and U2574 (N_2574,N_2401,N_2044);
and U2575 (N_2575,N_1798,N_1310);
xor U2576 (N_2576,In_1916,N_1920);
nand U2577 (N_2577,N_2315,N_2317);
nor U2578 (N_2578,N_627,In_78);
xnor U2579 (N_2579,In_4876,In_4575);
nor U2580 (N_2580,In_4178,In_16);
and U2581 (N_2581,In_793,In_4719);
or U2582 (N_2582,In_783,In_356);
nand U2583 (N_2583,N_1690,In_519);
nor U2584 (N_2584,N_2308,N_748);
or U2585 (N_2585,N_103,In_4930);
nand U2586 (N_2586,N_1915,N_1056);
nor U2587 (N_2587,In_2264,In_199);
xnor U2588 (N_2588,N_1336,N_1657);
xor U2589 (N_2589,N_2396,In_1574);
xor U2590 (N_2590,In_1033,In_2365);
or U2591 (N_2591,In_2763,N_2042);
and U2592 (N_2592,N_1451,In_4591);
xor U2593 (N_2593,N_2050,N_1143);
nand U2594 (N_2594,In_1325,N_737);
xnor U2595 (N_2595,N_2374,N_2024);
nor U2596 (N_2596,N_2235,In_2573);
or U2597 (N_2597,In_298,N_2201);
and U2598 (N_2598,In_3668,N_2494);
nor U2599 (N_2599,N_778,In_3702);
and U2600 (N_2600,In_152,In_4630);
nand U2601 (N_2601,In_2018,N_1785);
nor U2602 (N_2602,In_2646,In_3426);
and U2603 (N_2603,In_4968,N_2365);
nand U2604 (N_2604,N_850,In_3577);
nor U2605 (N_2605,N_536,N_2430);
and U2606 (N_2606,In_1785,In_4547);
nor U2607 (N_2607,In_4848,N_1795);
xor U2608 (N_2608,In_2097,In_2019);
nor U2609 (N_2609,In_626,N_918);
xnor U2610 (N_2610,In_2795,In_1989);
nand U2611 (N_2611,N_2112,In_1317);
nand U2612 (N_2612,N_2184,In_1858);
xor U2613 (N_2613,In_57,In_1032);
or U2614 (N_2614,In_1002,In_2056);
and U2615 (N_2615,In_4730,N_61);
or U2616 (N_2616,In_2286,N_1566);
and U2617 (N_2617,N_1083,In_3721);
and U2618 (N_2618,N_1580,N_699);
or U2619 (N_2619,In_634,N_2345);
nor U2620 (N_2620,N_2225,N_1558);
nand U2621 (N_2621,In_1395,In_4416);
or U2622 (N_2622,In_722,In_2498);
xnor U2623 (N_2623,N_1926,N_2193);
nor U2624 (N_2624,In_4690,In_1018);
or U2625 (N_2625,In_1991,N_2075);
and U2626 (N_2626,In_2892,N_1958);
xnor U2627 (N_2627,N_1847,N_771);
nand U2628 (N_2628,N_2263,N_1331);
and U2629 (N_2629,N_1323,In_2906);
xnor U2630 (N_2630,In_2852,N_1723);
and U2631 (N_2631,In_1825,In_2711);
nor U2632 (N_2632,In_3789,N_2375);
nand U2633 (N_2633,N_1840,N_834);
xnor U2634 (N_2634,N_1733,In_1755);
nand U2635 (N_2635,In_1055,N_678);
or U2636 (N_2636,In_2246,N_443);
or U2637 (N_2637,In_4465,In_3539);
nand U2638 (N_2638,In_2253,In_3630);
xor U2639 (N_2639,In_1447,N_2218);
and U2640 (N_2640,In_3828,N_2158);
nor U2641 (N_2641,N_1024,In_1265);
nor U2642 (N_2642,In_4717,In_2335);
nand U2643 (N_2643,N_1708,In_1844);
or U2644 (N_2644,In_877,N_2475);
and U2645 (N_2645,N_1216,In_3131);
xor U2646 (N_2646,In_2198,N_311);
nor U2647 (N_2647,In_1597,In_1102);
xnor U2648 (N_2648,N_1643,In_550);
or U2649 (N_2649,N_2282,N_1902);
nor U2650 (N_2650,N_2321,In_649);
or U2651 (N_2651,In_282,In_132);
or U2652 (N_2652,N_99,In_2899);
nor U2653 (N_2653,N_2045,In_642);
or U2654 (N_2654,N_2422,N_2256);
and U2655 (N_2655,In_831,In_1090);
xor U2656 (N_2656,N_1517,N_1540);
nor U2657 (N_2657,In_3589,In_2548);
or U2658 (N_2658,N_1306,N_2251);
xor U2659 (N_2659,N_1985,In_4473);
or U2660 (N_2660,N_1872,In_4758);
and U2661 (N_2661,N_2496,In_2145);
and U2662 (N_2662,In_4895,N_2334);
nor U2663 (N_2663,N_2487,In_1919);
nand U2664 (N_2664,N_1335,N_2481);
or U2665 (N_2665,In_699,N_2022);
xnor U2666 (N_2666,In_4498,In_3423);
and U2667 (N_2667,In_3500,N_322);
nor U2668 (N_2668,In_4926,In_1388);
nor U2669 (N_2669,In_1082,In_3031);
xnor U2670 (N_2670,N_152,In_4574);
and U2671 (N_2671,N_1960,N_2471);
or U2672 (N_2672,N_2426,N_1258);
xnor U2673 (N_2673,N_1185,In_4087);
nor U2674 (N_2674,N_1394,N_631);
or U2675 (N_2675,N_2247,N_1532);
and U2676 (N_2676,In_2478,N_2392);
or U2677 (N_2677,N_1307,In_3296);
or U2678 (N_2678,N_1548,In_3949);
nor U2679 (N_2679,In_4340,In_4050);
nand U2680 (N_2680,In_4123,In_3063);
xnor U2681 (N_2681,In_1228,In_4287);
or U2682 (N_2682,N_796,In_4738);
nor U2683 (N_2683,In_4841,N_2438);
nand U2684 (N_2684,In_669,In_4745);
and U2685 (N_2685,N_2020,In_4214);
or U2686 (N_2686,N_1893,N_74);
nor U2687 (N_2687,In_3133,In_3207);
nor U2688 (N_2688,N_1161,In_1847);
xnor U2689 (N_2689,N_2061,N_1838);
nor U2690 (N_2690,In_4865,In_2981);
and U2691 (N_2691,N_30,N_638);
xor U2692 (N_2692,In_2187,In_1000);
nand U2693 (N_2693,In_169,N_2483);
xor U2694 (N_2694,In_4605,In_175);
nor U2695 (N_2695,In_1170,N_2117);
nor U2696 (N_2696,N_2188,N_2120);
or U2697 (N_2697,In_3885,In_868);
and U2698 (N_2698,N_393,In_4946);
and U2699 (N_2699,In_4288,In_2164);
or U2700 (N_2700,N_2388,In_3703);
nor U2701 (N_2701,N_980,N_2272);
nor U2702 (N_2702,N_2382,N_2486);
nand U2703 (N_2703,N_35,In_2673);
nor U2704 (N_2704,N_1868,N_2147);
xnor U2705 (N_2705,N_938,N_2160);
and U2706 (N_2706,N_750,N_389);
nor U2707 (N_2707,N_1773,In_3713);
and U2708 (N_2708,N_1210,N_310);
and U2709 (N_2709,N_1988,N_1953);
and U2710 (N_2710,N_1049,In_4871);
or U2711 (N_2711,In_3001,In_4343);
nor U2712 (N_2712,N_2233,In_1248);
nand U2713 (N_2713,In_1058,N_2393);
nor U2714 (N_2714,In_4657,In_2349);
or U2715 (N_2715,In_2610,In_1332);
and U2716 (N_2716,N_350,N_2180);
nor U2717 (N_2717,In_1601,In_4812);
and U2718 (N_2718,N_1277,In_4065);
xor U2719 (N_2719,N_1305,N_2257);
and U2720 (N_2720,In_742,In_1790);
nand U2721 (N_2721,In_4713,N_2019);
nand U2722 (N_2722,In_940,N_2108);
nand U2723 (N_2723,In_1107,N_1569);
or U2724 (N_2724,In_3081,In_360);
nand U2725 (N_2725,In_1305,In_2247);
and U2726 (N_2726,In_3298,In_4541);
xnor U2727 (N_2727,In_809,N_1516);
nand U2728 (N_2728,N_2411,In_1811);
nor U2729 (N_2729,N_1825,N_2473);
xnor U2730 (N_2730,N_2155,In_842);
and U2731 (N_2731,N_2335,In_1621);
xor U2732 (N_2732,N_2128,N_1766);
and U2733 (N_2733,N_50,In_1739);
or U2734 (N_2734,N_39,In_1216);
nand U2735 (N_2735,N_1895,In_3644);
and U2736 (N_2736,In_3272,N_1065);
nand U2737 (N_2737,N_1922,In_431);
and U2738 (N_2738,In_4945,N_1678);
and U2739 (N_2739,In_3243,N_2432);
nand U2740 (N_2740,In_3018,In_3975);
and U2741 (N_2741,In_2764,In_3689);
and U2742 (N_2742,In_3168,N_2367);
xnor U2743 (N_2743,N_604,In_4922);
and U2744 (N_2744,In_433,In_149);
and U2745 (N_2745,In_2961,N_1966);
and U2746 (N_2746,In_1836,In_462);
nand U2747 (N_2747,N_1297,In_3552);
and U2748 (N_2748,N_2451,N_1951);
nor U2749 (N_2749,In_3923,N_2444);
xnor U2750 (N_2750,In_1169,In_577);
and U2751 (N_2751,N_1249,N_1263);
or U2752 (N_2752,In_3169,N_561);
nand U2753 (N_2753,N_2351,N_1203);
or U2754 (N_2754,In_2853,N_1814);
and U2755 (N_2755,N_2029,In_4831);
or U2756 (N_2756,In_1224,N_2489);
or U2757 (N_2757,N_446,In_1931);
nor U2758 (N_2758,N_2608,In_1463);
xor U2759 (N_2759,N_1841,N_2400);
nor U2760 (N_2760,N_2353,In_1328);
xnor U2761 (N_2761,N_1931,N_1730);
xor U2762 (N_2762,N_721,N_1439);
or U2763 (N_2763,In_686,N_1435);
nor U2764 (N_2764,N_2423,In_1519);
nand U2765 (N_2765,In_491,N_2719);
nand U2766 (N_2766,N_612,In_3029);
xor U2767 (N_2767,N_2349,In_1135);
xnor U2768 (N_2768,N_2242,N_2466);
or U2769 (N_2769,In_3624,In_683);
and U2770 (N_2770,In_3097,N_2372);
and U2771 (N_2771,N_602,N_1943);
or U2772 (N_2772,N_1793,In_2838);
and U2773 (N_2773,N_2267,In_1638);
nor U2774 (N_2774,N_293,In_2584);
nand U2775 (N_2775,N_2046,N_2236);
and U2776 (N_2776,In_4218,N_2186);
or U2777 (N_2777,N_2222,N_2616);
xor U2778 (N_2778,N_1816,N_1937);
and U2779 (N_2779,N_2559,N_1470);
nor U2780 (N_2780,N_1334,In_2088);
nor U2781 (N_2781,In_1445,In_721);
xnor U2782 (N_2782,In_2890,N_2098);
nor U2783 (N_2783,N_2133,N_2302);
nand U2784 (N_2784,N_2605,N_2270);
and U2785 (N_2785,In_4206,N_1474);
nor U2786 (N_2786,In_4982,N_2591);
or U2787 (N_2787,In_2829,N_1449);
xnor U2788 (N_2788,N_1009,N_2652);
xor U2789 (N_2789,In_2822,N_2389);
xnor U2790 (N_2790,N_2595,In_3233);
nand U2791 (N_2791,N_1084,N_1275);
and U2792 (N_2792,In_4166,In_449);
or U2793 (N_2793,In_3397,N_1211);
and U2794 (N_2794,N_192,In_509);
xnor U2795 (N_2795,In_3632,N_2130);
xnor U2796 (N_2796,N_150,N_1586);
or U2797 (N_2797,In_3967,In_4531);
xor U2798 (N_2798,N_2662,N_2101);
and U2799 (N_2799,N_1651,N_449);
and U2800 (N_2800,N_2043,N_1777);
and U2801 (N_2801,In_4983,N_2294);
xor U2802 (N_2802,N_2581,N_2630);
nor U2803 (N_2803,N_1653,N_2560);
xor U2804 (N_2804,N_2051,In_1077);
xor U2805 (N_2805,N_2012,In_71);
and U2806 (N_2806,N_2649,In_4049);
xnor U2807 (N_2807,In_795,In_4643);
or U2808 (N_2808,In_1956,N_505);
or U2809 (N_2809,N_1554,N_2240);
or U2810 (N_2810,N_2099,N_2285);
nand U2811 (N_2811,In_3285,In_1635);
and U2812 (N_2812,N_711,N_1160);
nor U2813 (N_2813,N_1990,N_1472);
and U2814 (N_2814,In_4718,N_1476);
xor U2815 (N_2815,N_1848,N_633);
nor U2816 (N_2816,In_1391,N_2443);
or U2817 (N_2817,N_1716,In_1807);
xnor U2818 (N_2818,In_495,In_2803);
xor U2819 (N_2819,N_2544,N_2524);
and U2820 (N_2820,N_2419,In_3629);
xnor U2821 (N_2821,In_3297,In_2569);
and U2822 (N_2822,N_2154,N_2726);
or U2823 (N_2823,N_558,In_910);
xor U2824 (N_2824,N_2331,N_2406);
and U2825 (N_2825,N_2724,N_1453);
nand U2826 (N_2826,In_3465,N_922);
or U2827 (N_2827,N_576,N_1406);
xnor U2828 (N_2828,In_2997,In_1198);
and U2829 (N_2829,N_2528,N_2690);
nor U2830 (N_2830,N_261,In_2420);
nor U2831 (N_2831,In_1383,N_2546);
nand U2832 (N_2832,In_212,N_936);
or U2833 (N_2833,N_1490,In_1651);
xor U2834 (N_2834,N_2227,In_4345);
xor U2835 (N_2835,In_3065,N_1741);
or U2836 (N_2836,N_2296,In_1367);
xor U2837 (N_2837,In_2023,In_2574);
and U2838 (N_2838,N_2456,In_437);
xor U2839 (N_2839,N_2134,N_2361);
nor U2840 (N_2840,In_559,In_1308);
nor U2841 (N_2841,In_3618,N_1061);
and U2842 (N_2842,N_2624,N_2555);
nor U2843 (N_2843,N_2739,N_1359);
and U2844 (N_2844,N_1346,In_4990);
xnor U2845 (N_2845,N_626,In_520);
or U2846 (N_2846,N_2424,N_2569);
or U2847 (N_2847,In_1221,In_98);
and U2848 (N_2848,N_2542,N_2410);
nor U2849 (N_2849,In_4987,In_487);
or U2850 (N_2850,N_2027,N_1770);
nor U2851 (N_2851,N_2175,N_2611);
nor U2852 (N_2852,N_1903,N_1776);
or U2853 (N_2853,N_1127,In_380);
xor U2854 (N_2854,N_1672,N_2467);
nand U2855 (N_2855,N_2703,In_2128);
nor U2856 (N_2856,N_2448,N_1722);
nand U2857 (N_2857,N_2359,N_1778);
xnor U2858 (N_2858,In_41,In_2229);
nor U2859 (N_2859,N_1948,N_1303);
or U2860 (N_2860,N_1583,In_210);
nor U2861 (N_2861,In_949,In_702);
xor U2862 (N_2862,N_472,In_3240);
and U2863 (N_2863,In_104,N_2329);
or U2864 (N_2864,In_2733,In_761);
xnor U2865 (N_2865,N_2708,N_345);
nand U2866 (N_2866,In_4160,N_2021);
xor U2867 (N_2867,N_2248,N_2749);
or U2868 (N_2868,In_966,N_1805);
nor U2869 (N_2869,In_1148,N_2434);
nor U2870 (N_2870,In_69,In_1178);
or U2871 (N_2871,N_2268,N_585);
xor U2872 (N_2872,N_2553,N_2283);
nor U2873 (N_2873,In_4783,In_1336);
and U2874 (N_2874,In_2878,In_1432);
nor U2875 (N_2875,N_2119,In_3476);
xor U2876 (N_2876,N_2033,N_2060);
nor U2877 (N_2877,N_1746,In_2137);
nand U2878 (N_2878,N_1120,N_1941);
or U2879 (N_2879,In_3170,N_1321);
nand U2880 (N_2880,In_3558,In_4935);
and U2881 (N_2881,In_4235,In_2339);
and U2882 (N_2882,N_2122,N_419);
nor U2883 (N_2883,N_2510,In_3023);
xnor U2884 (N_2884,In_2670,In_270);
or U2885 (N_2885,N_2550,In_1718);
or U2886 (N_2886,N_338,N_173);
nor U2887 (N_2887,In_3040,N_2239);
nor U2888 (N_2888,N_2295,N_1750);
and U2889 (N_2889,N_1962,N_73);
or U2890 (N_2890,N_2562,N_2354);
nand U2891 (N_2891,In_1071,In_3172);
xnor U2892 (N_2892,N_2007,In_4756);
xnor U2893 (N_2893,In_812,N_839);
and U2894 (N_2894,N_889,In_2503);
nor U2895 (N_2895,N_2191,N_722);
xnor U2896 (N_2896,N_1925,N_2523);
xor U2897 (N_2897,N_1371,In_576);
nand U2898 (N_2898,In_1072,N_2399);
and U2899 (N_2899,N_1767,N_2588);
and U2900 (N_2900,N_1831,N_2450);
nand U2901 (N_2901,N_1078,N_2300);
nor U2902 (N_2902,In_2404,N_2452);
xnor U2903 (N_2903,In_3227,N_2479);
nor U2904 (N_2904,In_4246,N_2730);
or U2905 (N_2905,N_1873,N_2326);
or U2906 (N_2906,N_1839,In_4102);
xnor U2907 (N_2907,N_2086,In_3252);
or U2908 (N_2908,N_2181,N_1565);
nor U2909 (N_2909,N_716,N_708);
or U2910 (N_2910,N_2609,N_1997);
nor U2911 (N_2911,In_2251,In_254);
xnor U2912 (N_2912,In_4942,N_262);
xor U2913 (N_2913,In_1908,N_433);
xor U2914 (N_2914,N_1450,N_1180);
xnor U2915 (N_2915,N_1980,N_1409);
nand U2916 (N_2916,In_939,N_1863);
xor U2917 (N_2917,N_101,In_3766);
and U2918 (N_2918,N_34,In_2800);
and U2919 (N_2919,N_523,In_4845);
or U2920 (N_2920,N_1533,N_1311);
nand U2921 (N_2921,In_2209,In_1273);
or U2922 (N_2922,N_1284,N_2474);
or U2923 (N_2923,In_1520,N_1543);
and U2924 (N_2924,N_2165,N_2304);
or U2925 (N_2925,N_198,In_3653);
and U2926 (N_2926,N_2123,In_1351);
or U2927 (N_2927,In_454,N_930);
nor U2928 (N_2928,In_4109,N_2597);
and U2929 (N_2929,N_1442,N_1482);
nor U2930 (N_2930,N_407,In_3574);
and U2931 (N_2931,N_2187,N_1465);
nand U2932 (N_2932,N_2532,N_1787);
nor U2933 (N_2933,N_204,In_3329);
and U2934 (N_2934,In_573,N_415);
nor U2935 (N_2935,N_2065,In_2623);
or U2936 (N_2936,In_2825,In_2972);
or U2937 (N_2937,N_199,In_3892);
nor U2938 (N_2938,N_1375,N_739);
or U2939 (N_2939,N_828,In_1888);
nor U2940 (N_2940,In_2130,In_45);
nor U2941 (N_2941,In_1955,N_1423);
nor U2942 (N_2942,N_2379,N_48);
xor U2943 (N_2943,In_3504,In_2601);
and U2944 (N_2944,In_2244,N_593);
xnor U2945 (N_2945,In_2245,N_2278);
nor U2946 (N_2946,N_913,N_2403);
nor U2947 (N_2947,In_1644,N_2420);
nand U2948 (N_2948,In_470,N_2643);
or U2949 (N_2949,N_205,N_541);
or U2950 (N_2950,In_3069,In_4833);
and U2951 (N_2951,N_2677,In_1587);
nand U2952 (N_2952,N_2177,In_2289);
and U2953 (N_2953,N_2536,In_2636);
and U2954 (N_2954,N_2298,N_586);
nor U2955 (N_2955,In_4728,In_740);
and U2956 (N_2956,In_2505,N_2220);
and U2957 (N_2957,In_1319,N_195);
or U2958 (N_2958,N_2115,In_3617);
or U2959 (N_2959,In_2408,N_777);
xor U2960 (N_2960,N_1288,In_191);
and U2961 (N_2961,N_1141,N_6);
nor U2962 (N_2962,In_1437,N_1003);
nand U2963 (N_2963,In_4849,N_1309);
nor U2964 (N_2964,In_3954,In_3676);
xor U2965 (N_2965,N_1684,N_438);
nor U2966 (N_2966,N_2319,In_3093);
or U2967 (N_2967,N_105,In_1925);
nand U2968 (N_2968,In_4951,N_2113);
or U2969 (N_2969,N_2386,N_33);
and U2970 (N_2970,In_3433,N_910);
xnor U2971 (N_2971,N_2655,In_3315);
nor U2972 (N_2972,In_3087,N_2213);
xnor U2973 (N_2973,N_2525,In_667);
and U2974 (N_2974,N_2656,N_2737);
nor U2975 (N_2975,In_3664,In_3166);
or U2976 (N_2976,N_2437,N_2000);
nor U2977 (N_2977,N_2207,In_3760);
and U2978 (N_2978,N_954,In_4793);
nand U2979 (N_2979,N_1132,In_295);
xor U2980 (N_2980,N_2587,In_4034);
and U2981 (N_2981,In_119,N_2718);
or U2982 (N_2982,N_376,N_2425);
or U2983 (N_2983,In_4155,In_320);
and U2984 (N_2984,In_247,N_2287);
nand U2985 (N_2985,N_1754,In_4601);
nand U2986 (N_2986,N_2357,N_1901);
nor U2987 (N_2987,In_1610,N_463);
nor U2988 (N_2988,N_2501,N_368);
xnor U2989 (N_2989,N_1541,N_2157);
or U2990 (N_2990,N_2069,In_3101);
nor U2991 (N_2991,N_1623,N_2026);
nand U2992 (N_2992,N_1168,In_3785);
xnor U2993 (N_2993,N_2540,N_1326);
nand U2994 (N_2994,N_2249,In_659);
and U2995 (N_2995,N_2390,N_2538);
xor U2996 (N_2996,N_2380,N_1709);
xnor U2997 (N_2997,N_2053,In_4534);
nor U2998 (N_2998,N_2404,In_1468);
or U2999 (N_2999,N_1859,In_1242);
xor U3000 (N_3000,In_30,N_1126);
xnor U3001 (N_3001,N_812,N_2898);
nor U3002 (N_3002,N_2210,N_2100);
nor U3003 (N_3003,In_1676,N_2791);
nand U3004 (N_3004,In_4975,N_135);
nor U3005 (N_3005,In_163,In_1014);
nor U3006 (N_3006,In_4367,N_160);
nor U3007 (N_3007,N_2816,In_2267);
xor U3008 (N_3008,In_1517,N_2826);
or U3009 (N_3009,N_2691,N_2760);
nor U3010 (N_3010,N_2169,N_1191);
nor U3011 (N_3011,In_299,In_4444);
nor U3012 (N_3012,N_2862,N_1680);
and U3013 (N_3013,N_2506,N_1978);
and U3014 (N_3014,N_870,N_2934);
nor U3015 (N_3015,N_2290,In_4133);
nor U3016 (N_3016,In_17,N_439);
nor U3017 (N_3017,N_2877,N_2977);
nand U3018 (N_3018,N_803,N_2385);
nand U3019 (N_3019,N_783,N_2095);
nor U3020 (N_3020,In_3401,N_1067);
or U3021 (N_3021,In_2414,N_2551);
nor U3022 (N_3022,N_17,N_2773);
and U3023 (N_3023,In_3868,In_233);
and U3024 (N_3024,N_2918,N_2221);
or U3025 (N_3025,In_4078,N_2607);
nand U3026 (N_3026,In_1386,In_2129);
nor U3027 (N_3027,In_3750,N_2284);
xor U3028 (N_3028,N_1383,N_806);
nor U3029 (N_3029,In_4881,N_969);
and U3030 (N_3030,In_4202,N_2964);
nor U3031 (N_3031,N_1710,In_176);
nor U3032 (N_3032,In_4530,N_1017);
nor U3033 (N_3033,N_2262,N_2337);
xnor U3034 (N_3034,N_1053,N_2096);
nand U3035 (N_3035,N_2698,N_1578);
nor U3036 (N_3036,In_3147,N_1627);
or U3037 (N_3037,In_3978,In_3402);
and U3038 (N_3038,N_1835,N_2276);
and U3039 (N_3039,N_669,N_948);
nand U3040 (N_3040,N_2092,N_2837);
nand U3041 (N_3041,In_979,In_717);
xnor U3042 (N_3042,In_4642,N_2545);
nor U3043 (N_3043,In_4914,N_2808);
or U3044 (N_3044,N_520,In_4277);
nand U3045 (N_3045,In_1042,N_2747);
nand U3046 (N_3046,N_798,In_1666);
or U3047 (N_3047,N_1224,N_663);
and U3048 (N_3048,In_3356,N_821);
and U3049 (N_3049,N_2505,In_1128);
nor U3050 (N_3050,N_1189,In_3124);
xor U3051 (N_3051,In_3320,N_2681);
or U3052 (N_3052,N_1398,N_1769);
nand U3053 (N_3053,In_1880,N_2371);
nor U3054 (N_3054,N_603,In_467);
or U3055 (N_3055,N_2322,N_1759);
or U3056 (N_3056,N_2847,N_1487);
nor U3057 (N_3057,N_2347,In_778);
and U3058 (N_3058,N_249,N_1760);
or U3059 (N_3059,N_2995,N_688);
or U3060 (N_3060,In_2009,In_1219);
nor U3061 (N_3061,N_1900,In_2473);
nor U3062 (N_3062,N_2878,In_801);
xnor U3063 (N_3063,N_2672,N_1182);
or U3064 (N_3064,N_1162,In_2778);
xor U3065 (N_3065,In_2575,In_1945);
nand U3066 (N_3066,In_4493,N_1157);
nand U3067 (N_3067,In_1801,N_2980);
nor U3068 (N_3068,In_1595,In_3437);
and U3069 (N_3069,N_1697,N_2413);
and U3070 (N_3070,N_2224,In_1910);
nor U3071 (N_3071,N_46,N_2855);
nand U3072 (N_3072,In_4212,N_2102);
nor U3073 (N_3073,In_2332,N_2813);
and U3074 (N_3074,N_64,N_2814);
xor U3075 (N_3075,In_4359,N_2131);
nand U3076 (N_3076,N_2189,N_1114);
or U3077 (N_3077,N_923,N_2346);
nand U3078 (N_3078,N_2350,In_2132);
nor U3079 (N_3079,In_2486,N_1208);
nand U3080 (N_3080,In_4286,In_3250);
or U3081 (N_3081,N_2880,N_2418);
nand U3082 (N_3082,N_2873,In_3286);
or U3083 (N_3083,N_2956,N_2762);
or U3084 (N_3084,N_2851,N_2414);
xnor U3085 (N_3085,N_2840,N_240);
xnor U3086 (N_3086,N_411,N_2159);
nor U3087 (N_3087,N_1577,In_2854);
nand U3088 (N_3088,N_1269,N_2775);
and U3089 (N_3089,N_2497,In_4757);
nand U3090 (N_3090,N_2572,N_84);
or U3091 (N_3091,N_1230,In_4768);
and U3092 (N_3092,In_1710,In_2809);
nor U3093 (N_3093,N_1152,N_1428);
nand U3094 (N_3094,In_3449,N_2049);
nor U3095 (N_3095,N_2634,In_4660);
xor U3096 (N_3096,In_3620,N_2732);
or U3097 (N_3097,N_2311,In_709);
nand U3098 (N_3098,N_1748,In_4161);
and U3099 (N_3099,N_2919,In_3288);
and U3100 (N_3100,In_1967,N_2740);
nand U3101 (N_3101,N_2125,N_2107);
and U3102 (N_3102,N_1799,In_4701);
nor U3103 (N_3103,N_109,N_1129);
or U3104 (N_3104,N_2498,N_526);
or U3105 (N_3105,N_2197,N_1751);
nand U3106 (N_3106,In_675,N_2692);
and U3107 (N_3107,N_1047,N_2111);
xor U3108 (N_3108,N_2369,In_1839);
xor U3109 (N_3109,In_933,N_2200);
and U3110 (N_3110,N_1412,N_1342);
nor U3111 (N_3111,N_2325,N_2635);
xnor U3112 (N_3112,In_4681,N_2863);
and U3113 (N_3113,In_105,In_4891);
and U3114 (N_3114,In_794,N_2907);
xor U3115 (N_3115,N_2577,In_1593);
nand U3116 (N_3116,N_129,In_2597);
and U3117 (N_3117,In_1628,N_1333);
nor U3118 (N_3118,In_4232,In_4625);
and U3119 (N_3119,N_2618,In_1814);
nor U3120 (N_3120,In_4839,In_817);
nand U3121 (N_3121,N_1432,N_2453);
or U3122 (N_3122,In_4967,N_2756);
and U3123 (N_3123,In_3231,N_1213);
nor U3124 (N_3124,In_4458,N_2514);
nand U3125 (N_3125,In_4668,N_394);
or U3126 (N_3126,In_1377,In_514);
and U3127 (N_3127,N_734,N_2064);
nand U3128 (N_3128,In_1745,In_4640);
xor U3129 (N_3129,N_2590,In_1985);
nand U3130 (N_3130,N_794,N_2171);
and U3131 (N_3131,In_4375,In_2263);
or U3132 (N_3132,N_450,N_2796);
and U3133 (N_3133,N_2534,N_2066);
xnor U3134 (N_3134,N_2202,In_3764);
xor U3135 (N_3135,In_408,In_3637);
nand U3136 (N_3136,N_1782,N_2176);
or U3137 (N_3137,In_4373,In_1514);
nor U3138 (N_3138,N_1458,N_2395);
or U3139 (N_3139,In_2188,N_2243);
nand U3140 (N_3140,In_4984,In_4490);
and U3141 (N_3141,N_2674,N_2829);
xor U3142 (N_3142,In_4440,N_745);
or U3143 (N_3143,N_1599,In_3688);
and U3144 (N_3144,N_1090,In_4119);
nor U3145 (N_3145,In_4716,N_2054);
and U3146 (N_3146,N_852,N_2564);
xor U3147 (N_3147,N_1550,In_1690);
or U3148 (N_3148,N_2817,In_3404);
and U3149 (N_3149,In_3266,N_726);
xor U3150 (N_3150,N_1538,In_501);
nand U3151 (N_3151,N_1897,N_1138);
nand U3152 (N_3152,In_4798,N_2273);
or U3153 (N_3153,In_3881,N_1011);
nor U3154 (N_3154,N_2779,N_2582);
or U3155 (N_3155,N_2554,N_2352);
xnor U3156 (N_3156,In_1334,N_2944);
or U3157 (N_3157,N_2598,N_2872);
nor U3158 (N_3158,N_2127,N_2913);
nand U3159 (N_3159,N_1349,N_1460);
nor U3160 (N_3160,In_609,In_2737);
or U3161 (N_3161,In_1933,N_2978);
and U3162 (N_3162,N_905,In_974);
or U3163 (N_3163,N_455,In_2934);
xor U3164 (N_3164,In_2470,In_549);
xnor U3165 (N_3165,N_2067,N_387);
nand U3166 (N_3166,N_1885,In_3968);
or U3167 (N_3167,N_1503,N_2416);
and U3168 (N_3168,N_1744,N_2520);
or U3169 (N_3169,N_1212,In_4071);
or U3170 (N_3170,N_2277,N_2439);
and U3171 (N_3171,N_364,N_1510);
xor U3172 (N_3172,N_892,N_2109);
nand U3173 (N_3173,N_2417,N_2895);
and U3174 (N_3174,N_2810,N_2957);
nand U3175 (N_3175,In_3931,N_2149);
nand U3176 (N_3176,N_1444,N_2265);
nand U3177 (N_3177,N_2948,N_2667);
xor U3178 (N_3178,N_836,In_3869);
nor U3179 (N_3179,In_982,In_3042);
nand U3180 (N_3180,In_907,N_334);
or U3181 (N_3181,N_2792,N_2812);
or U3182 (N_3182,N_2849,In_3386);
xor U3183 (N_3183,In_676,In_1433);
or U3184 (N_3184,N_1644,N_1251);
nor U3185 (N_3185,In_829,In_1356);
nand U3186 (N_3186,In_3336,In_194);
and U3187 (N_3187,N_2997,N_1584);
nor U3188 (N_3188,N_2811,In_1590);
xnor U3189 (N_3189,N_408,N_1609);
xnor U3190 (N_3190,N_2204,In_4905);
and U3191 (N_3191,In_1099,N_2472);
nor U3192 (N_3192,N_2927,In_59);
nand U3193 (N_3193,N_2599,In_342);
nor U3194 (N_3194,In_4557,In_1494);
or U3195 (N_3195,In_2769,N_2945);
nor U3196 (N_3196,In_4010,In_4675);
nand U3197 (N_3197,In_825,N_1780);
or U3198 (N_3198,In_3827,In_2272);
nand U3199 (N_3199,N_1687,N_555);
and U3200 (N_3200,In_3953,In_2765);
or U3201 (N_3201,N_550,N_682);
xnor U3202 (N_3202,N_2561,In_3206);
nand U3203 (N_3203,N_2216,N_2642);
or U3204 (N_3204,N_2340,N_2833);
or U3205 (N_3205,N_2938,N_2818);
or U3206 (N_3206,N_2804,N_2198);
xor U3207 (N_3207,In_3673,N_2402);
or U3208 (N_3208,N_2318,N_2827);
or U3209 (N_3209,In_4649,N_2993);
nand U3210 (N_3210,In_3847,N_1693);
or U3211 (N_3211,N_2912,In_3247);
nor U3212 (N_3212,N_1820,In_4957);
nor U3213 (N_3213,N_2986,In_411);
or U3214 (N_3214,In_1576,N_1520);
or U3215 (N_3215,N_1145,N_2279);
and U3216 (N_3216,In_2109,In_3625);
and U3217 (N_3217,N_180,N_1112);
and U3218 (N_3218,N_2694,In_3645);
xnor U3219 (N_3219,N_2875,In_3000);
nand U3220 (N_3220,In_3498,N_2892);
nand U3221 (N_3221,In_3700,In_2216);
nand U3222 (N_3222,N_2341,N_1035);
nand U3223 (N_3223,N_2745,In_4083);
and U3224 (N_3224,In_4118,N_886);
or U3225 (N_3225,In_2989,N_540);
nand U3226 (N_3226,In_1799,N_1737);
and U3227 (N_3227,N_1836,N_2920);
and U3228 (N_3228,N_1964,N_2800);
xor U3229 (N_3229,In_2688,N_2950);
nor U3230 (N_3230,In_2966,In_3805);
nor U3231 (N_3231,N_2488,In_2910);
nor U3232 (N_3232,N_2834,N_2743);
or U3233 (N_3233,In_2158,N_2231);
or U3234 (N_3234,N_2110,N_2260);
nand U3235 (N_3235,In_2338,N_2785);
nand U3236 (N_3236,N_959,In_2936);
xnor U3237 (N_3237,N_2576,N_2883);
xor U3238 (N_3238,In_2578,N_2515);
nand U3239 (N_3239,N_1611,In_1039);
or U3240 (N_3240,N_318,N_2394);
nor U3241 (N_3241,N_942,N_2610);
xnor U3242 (N_3242,N_2613,In_2208);
nand U3243 (N_3243,N_2781,In_1020);
xor U3244 (N_3244,N_2750,N_1164);
xor U3245 (N_3245,In_3955,In_2500);
or U3246 (N_3246,N_2366,In_2973);
or U3247 (N_3247,N_2949,In_2210);
nand U3248 (N_3248,In_345,In_116);
and U3249 (N_3249,N_592,In_4069);
nor U3250 (N_3250,In_418,N_1880);
and U3251 (N_3251,N_2377,N_3063);
xor U3252 (N_3252,In_2755,N_3095);
and U3253 (N_3253,In_4837,In_87);
nand U3254 (N_3254,N_2871,N_2038);
or U3255 (N_3255,N_2759,N_2654);
or U3256 (N_3256,In_729,In_245);
or U3257 (N_3257,N_1812,N_3127);
nand U3258 (N_3258,N_2223,In_706);
nand U3259 (N_3259,In_137,N_3187);
xnor U3260 (N_3260,N_3211,N_2293);
nand U3261 (N_3261,N_784,N_1788);
nand U3262 (N_3262,N_3135,N_2633);
and U3263 (N_3263,N_2289,In_3262);
nand U3264 (N_3264,N_2992,N_2442);
nor U3265 (N_3265,N_2788,N_2436);
or U3266 (N_3266,In_3843,N_698);
xnor U3267 (N_3267,N_2683,N_3042);
nor U3268 (N_3268,N_3184,In_4933);
nand U3269 (N_3269,N_2615,N_1630);
and U3270 (N_3270,N_2567,N_2751);
xnor U3271 (N_3271,N_897,In_1875);
xnor U3272 (N_3272,N_2509,N_445);
nand U3273 (N_3273,In_3935,N_2644);
xnor U3274 (N_3274,N_833,In_696);
nor U3275 (N_3275,N_379,N_2923);
nand U3276 (N_3276,In_3113,N_1002);
nor U3277 (N_3277,In_4750,N_3097);
xor U3278 (N_3278,In_4448,In_500);
or U3279 (N_3279,N_2234,N_1591);
nor U3280 (N_3280,In_3308,N_1606);
or U3281 (N_3281,N_2991,In_3481);
nor U3282 (N_3282,N_2330,In_2833);
xnor U3283 (N_3283,N_1253,N_2678);
and U3284 (N_3284,In_1881,N_3078);
nand U3285 (N_3285,N_1339,N_3083);
xnor U3286 (N_3286,N_2627,N_2464);
or U3287 (N_3287,In_2792,N_2795);
nor U3288 (N_3288,In_3817,N_2172);
nor U3289 (N_3289,In_3222,N_3112);
nor U3290 (N_3290,N_1829,N_230);
xnor U3291 (N_3291,N_715,N_988);
or U3292 (N_3292,N_641,N_2052);
or U3293 (N_3293,In_217,In_754);
xnor U3294 (N_3294,N_3024,N_2902);
nor U3295 (N_3295,In_2013,N_2093);
xor U3296 (N_3296,N_168,N_779);
nand U3297 (N_3297,In_3035,N_1989);
xor U3298 (N_3298,In_4317,N_2807);
xnor U3299 (N_3299,N_2011,In_2396);
xor U3300 (N_3300,In_3263,N_2928);
nand U3301 (N_3301,N_2790,In_1359);
and U3302 (N_3302,N_2070,N_616);
nand U3303 (N_3303,In_1616,N_1622);
nand U3304 (N_3304,N_3222,N_1534);
or U3305 (N_3305,In_1832,In_1897);
nor U3306 (N_3306,N_3203,In_4670);
nand U3307 (N_3307,N_1322,N_2885);
or U3308 (N_3308,N_2876,N_1525);
and U3309 (N_3309,N_1991,In_827);
or U3310 (N_3310,In_1898,In_3110);
nor U3311 (N_3311,In_1469,N_2548);
or U3312 (N_3312,In_3587,N_2583);
nor U3313 (N_3313,In_3363,N_1879);
or U3314 (N_3314,N_2663,N_3220);
nand U3315 (N_3315,N_355,In_4274);
or U3316 (N_3316,N_2668,N_3200);
or U3317 (N_3317,N_2163,In_4154);
nor U3318 (N_3318,N_3143,N_2500);
or U3319 (N_3319,In_860,In_432);
or U3320 (N_3320,N_2721,In_1143);
or U3321 (N_3321,N_2421,N_2879);
xnor U3322 (N_3322,In_664,N_2391);
and U3323 (N_3323,N_1851,N_915);
nor U3324 (N_3324,N_992,N_3009);
nand U3325 (N_3325,N_214,N_2619);
nor U3326 (N_3326,In_3420,N_2770);
or U3327 (N_3327,N_3105,N_522);
xor U3328 (N_3328,N_1724,N_2517);
and U3329 (N_3329,In_4423,In_3961);
or U3330 (N_3330,N_1797,N_1008);
or U3331 (N_3331,In_3965,N_3114);
or U3332 (N_3332,In_4244,N_2714);
nand U3333 (N_3333,In_2382,In_651);
nor U3334 (N_3334,N_3088,N_2823);
xnor U3335 (N_3335,N_3074,N_2632);
and U3336 (N_3336,N_2081,N_2660);
nand U3337 (N_3337,N_1875,In_3145);
or U3338 (N_3338,In_1871,N_3172);
or U3339 (N_3339,N_3236,N_1670);
xnor U3340 (N_3340,N_2537,N_3006);
nor U3341 (N_3341,N_1634,N_3056);
nand U3342 (N_3342,N_2255,In_2925);
or U3343 (N_3343,N_1783,N_624);
or U3344 (N_3344,N_1457,N_1645);
xnor U3345 (N_3345,N_1819,In_3165);
xor U3346 (N_3346,N_3091,N_3010);
or U3347 (N_3347,N_2757,N_1725);
and U3348 (N_3348,N_3029,N_1319);
and U3349 (N_3349,N_728,N_3087);
nand U3350 (N_3350,N_3034,N_2629);
nor U3351 (N_3351,N_2622,In_4319);
nor U3352 (N_3352,N_1522,In_4638);
nand U3353 (N_3353,In_3455,In_3979);
xor U3354 (N_3354,N_2952,N_1590);
xor U3355 (N_3355,N_2217,In_4985);
xor U3356 (N_3356,In_219,N_3113);
nor U3357 (N_3357,In_2324,N_723);
xor U3358 (N_3358,N_2575,N_2568);
nor U3359 (N_3359,In_750,N_2002);
nand U3360 (N_3360,In_648,N_1950);
and U3361 (N_3361,N_1669,N_1521);
or U3362 (N_3362,In_2040,In_918);
or U3363 (N_3363,N_2292,In_4349);
or U3364 (N_3364,N_104,In_3299);
nand U3365 (N_3365,N_3073,N_2344);
nor U3366 (N_3366,In_2467,In_1404);
nor U3367 (N_3367,In_2234,In_4077);
xnor U3368 (N_3368,In_2424,In_4450);
xor U3369 (N_3369,In_1607,In_234);
nand U3370 (N_3370,N_3177,In_1013);
nand U3371 (N_3371,N_2035,In_4089);
nand U3372 (N_3372,N_2648,N_431);
or U3373 (N_3373,In_535,In_2354);
or U3374 (N_3374,N_2925,N_2338);
and U3375 (N_3375,In_545,In_2309);
or U3376 (N_3376,N_2786,N_2975);
or U3377 (N_3377,N_2324,N_2707);
nor U3378 (N_3378,N_2360,N_3053);
and U3379 (N_3379,In_182,N_3241);
nand U3380 (N_3380,In_713,N_2513);
xor U3381 (N_3381,N_1621,N_1159);
and U3382 (N_3382,N_2178,In_540);
nand U3383 (N_3383,N_1271,N_2041);
or U3384 (N_3384,N_2736,N_3089);
xor U3385 (N_3385,N_1102,N_3108);
xnor U3386 (N_3386,In_1683,N_1415);
and U3387 (N_3387,N_2998,N_2967);
nor U3388 (N_3388,In_3459,In_379);
nand U3389 (N_3389,In_1771,N_1758);
nor U3390 (N_3390,N_2996,N_2015);
nand U3391 (N_3391,N_3153,N_2954);
or U3392 (N_3392,In_3654,N_2603);
nor U3393 (N_3393,N_976,N_3046);
nor U3394 (N_3394,N_2250,In_4731);
nand U3395 (N_3395,N_2535,N_23);
xnor U3396 (N_3396,N_3179,N_2614);
nor U3397 (N_3397,N_1665,N_363);
nor U3398 (N_3398,N_926,N_3195);
xor U3399 (N_3399,N_2617,In_2376);
or U3400 (N_3400,N_2651,N_1587);
or U3401 (N_3401,N_2689,N_2929);
and U3402 (N_3402,N_3119,N_3084);
nor U3403 (N_3403,N_1696,N_2921);
xor U3404 (N_3404,In_196,N_2985);
xor U3405 (N_3405,N_2645,In_2446);
xnor U3406 (N_3406,N_2604,N_3246);
xor U3407 (N_3407,N_2687,N_2671);
nand U3408 (N_3408,In_3303,N_347);
or U3409 (N_3409,N_1999,In_340);
and U3410 (N_3410,N_2917,N_1405);
or U3411 (N_3411,In_3887,In_1276);
xnor U3412 (N_3412,N_1891,N_123);
xnor U3413 (N_3413,N_3094,N_3018);
xnor U3414 (N_3414,N_2638,N_1542);
or U3415 (N_3415,N_2963,N_1753);
xnor U3416 (N_3416,In_865,N_3201);
nand U3417 (N_3417,N_2857,In_4402);
nand U3418 (N_3418,N_2858,In_1250);
nor U3419 (N_3419,N_2946,In_1529);
nor U3420 (N_3420,In_1035,N_1685);
xor U3421 (N_3421,N_3017,N_2266);
xnor U3422 (N_3422,N_567,N_3023);
or U3423 (N_3423,In_205,N_2305);
or U3424 (N_3424,In_1752,N_3199);
nor U3425 (N_3425,N_2547,N_2772);
nor U3426 (N_3426,In_3190,In_3368);
nor U3427 (N_3427,N_1270,N_3014);
nand U3428 (N_3428,N_1701,N_413);
or U3429 (N_3429,N_185,N_507);
or U3430 (N_3430,N_3231,N_2072);
or U3431 (N_3431,In_2773,N_69);
xor U3432 (N_3432,N_2819,N_3205);
and U3433 (N_3433,N_2526,In_4958);
and U3434 (N_3434,In_303,In_2790);
nor U3435 (N_3435,N_1123,N_3123);
and U3436 (N_3436,N_1364,N_2310);
and U3437 (N_3437,N_3142,N_3049);
nand U3438 (N_3438,N_2254,N_2628);
or U3439 (N_3439,N_3248,In_1012);
xnor U3440 (N_3440,In_731,N_496);
or U3441 (N_3441,N_2710,N_1896);
nor U3442 (N_3442,N_2894,N_2140);
and U3443 (N_3443,In_2685,In_2860);
and U3444 (N_3444,In_764,N_3244);
and U3445 (N_3445,N_3133,N_1867);
xnor U3446 (N_3446,N_2784,N_1144);
and U3447 (N_3447,N_2405,In_198);
or U3448 (N_3448,N_2541,In_1373);
nor U3449 (N_3449,N_2343,N_1358);
nor U3450 (N_3450,In_989,In_1080);
and U3451 (N_3451,In_4623,N_872);
or U3452 (N_3452,N_2034,N_3186);
nor U3453 (N_3453,N_3025,N_2031);
or U3454 (N_3454,N_2381,N_3191);
nand U3455 (N_3455,N_2566,N_2673);
and U3456 (N_3456,N_2805,N_1815);
and U3457 (N_3457,N_2228,N_2071);
xnor U3458 (N_3458,In_4217,N_3233);
and U3459 (N_3459,N_2647,In_1263);
and U3460 (N_3460,N_1884,In_3860);
or U3461 (N_3461,In_1387,N_3229);
xnor U3462 (N_3462,N_2973,N_3111);
or U3463 (N_3463,N_2981,In_2327);
xnor U3464 (N_3464,N_2793,N_2848);
xor U3465 (N_3465,In_1987,N_3213);
or U3466 (N_3466,N_2657,In_3690);
and U3467 (N_3467,N_2214,N_2794);
nand U3468 (N_3468,In_3313,In_554);
nand U3469 (N_3469,In_18,N_3079);
and U3470 (N_3470,N_3061,N_2373);
xor U3471 (N_3471,N_2078,N_2531);
and U3472 (N_3472,N_1122,N_1477);
nor U3473 (N_3473,In_1977,N_2853);
nor U3474 (N_3474,N_2281,N_1850);
xnor U3475 (N_3475,N_2435,N_2076);
or U3476 (N_3476,N_1757,N_2013);
or U3477 (N_3477,N_2008,N_3237);
xnor U3478 (N_3478,N_2780,N_2626);
xor U3479 (N_3479,N_1280,In_973);
xor U3480 (N_3480,N_2908,N_2445);
nor U3481 (N_3481,N_3156,N_1712);
and U3482 (N_3482,N_3057,In_2768);
nor U3483 (N_3483,N_3206,N_8);
nor U3484 (N_3484,N_3144,N_2782);
and U3485 (N_3485,N_813,N_2558);
and U3486 (N_3486,In_1380,N_760);
nand U3487 (N_3487,N_3174,N_2765);
or U3488 (N_3488,N_3038,N_1557);
and U3489 (N_3489,In_4249,N_3030);
nand U3490 (N_3490,In_878,N_2933);
nand U3491 (N_3491,N_2485,N_2574);
nor U3492 (N_3492,N_2915,In_55);
or U3493 (N_3493,N_1768,N_3149);
nor U3494 (N_3494,N_1673,In_258);
nor U3495 (N_3495,In_2939,N_238);
nand U3496 (N_3496,N_2440,In_662);
xnor U3497 (N_3497,N_3027,N_3036);
or U3498 (N_3498,In_2226,N_2953);
or U3499 (N_3499,In_4136,N_2623);
or U3500 (N_3500,N_1647,N_1866);
nor U3501 (N_3501,N_1574,In_1637);
xor U3502 (N_3502,N_2738,N_3425);
nor U3503 (N_3503,N_2940,N_3168);
xnor U3504 (N_3504,N_2699,In_4712);
nor U3505 (N_3505,N_1789,N_1304);
nor U3506 (N_3506,In_1840,In_2121);
nand U3507 (N_3507,N_3051,In_4398);
nor U3508 (N_3508,N_3256,N_3475);
nand U3509 (N_3509,N_2048,N_1972);
nand U3510 (N_3510,N_3401,N_3151);
and U3511 (N_3511,N_2679,N_2280);
xor U3512 (N_3512,N_2852,In_1456);
nor U3513 (N_3513,In_1428,N_294);
nor U3514 (N_3514,N_3202,In_1702);
nand U3515 (N_3515,N_2512,N_848);
or U3516 (N_3516,N_955,N_2836);
nand U3517 (N_3517,N_2664,In_3841);
nand U3518 (N_3518,N_534,In_416);
nor U3519 (N_3519,N_842,In_3091);
and U3520 (N_3520,N_1377,N_3161);
and U3521 (N_3521,N_1255,In_123);
nand U3522 (N_3522,N_3284,N_1396);
or U3523 (N_3523,N_3426,N_2170);
xor U3524 (N_3524,N_1936,In_4528);
or U3525 (N_3525,N_2983,N_112);
nand U3526 (N_3526,In_4610,N_2080);
nand U3527 (N_3527,N_3317,N_2735);
nor U3528 (N_3528,N_3304,N_128);
nor U3529 (N_3529,In_77,N_2700);
and U3530 (N_3530,N_3122,N_398);
or U3531 (N_3531,N_3118,N_2764);
or U3532 (N_3532,N_2370,N_1362);
nor U3533 (N_3533,N_2815,N_474);
nand U3534 (N_3534,N_184,In_2585);
nand U3535 (N_3535,N_2713,In_135);
xor U3536 (N_3536,In_4781,In_4497);
nand U3537 (N_3537,N_3369,N_2333);
or U3538 (N_3538,N_3257,N_791);
xnor U3539 (N_3539,In_2760,N_2962);
xor U3540 (N_3540,N_2090,In_3677);
nand U3541 (N_3541,N_3085,In_2278);
nand U3542 (N_3542,N_3002,N_1539);
and U3543 (N_3543,In_4924,In_516);
or U3544 (N_3544,N_3381,N_2478);
nor U3545 (N_3545,N_3442,N_3380);
nor U3546 (N_3546,N_3155,N_0);
nand U3547 (N_3547,N_3066,N_1870);
and U3548 (N_3548,N_2798,N_1361);
nand U3549 (N_3549,N_2144,In_1672);
nor U3550 (N_3550,N_894,N_89);
xor U3551 (N_3551,N_2383,N_1717);
nor U3552 (N_3552,N_3499,N_1675);
nor U3553 (N_3553,In_3346,N_1527);
and U3554 (N_3554,N_2313,In_2678);
and U3555 (N_3555,N_1929,N_3216);
or U3556 (N_3556,N_3055,N_3267);
xor U3557 (N_3557,In_4284,In_1678);
and U3558 (N_3558,In_4149,N_511);
nand U3559 (N_3559,N_3272,N_3337);
nand U3560 (N_3560,N_3402,N_1899);
and U3561 (N_3561,N_3166,N_2530);
nor U3562 (N_3562,N_397,N_3159);
nand U3563 (N_3563,In_4378,N_2676);
xnor U3564 (N_3564,N_1771,N_3209);
nand U3565 (N_3565,In_1982,N_410);
nand U3566 (N_3566,N_1384,N_1355);
xor U3567 (N_3567,In_4802,In_2310);
xnor U3568 (N_3568,N_3165,N_3363);
nand U3569 (N_3569,N_846,In_3901);
or U3570 (N_3570,N_945,In_4435);
or U3571 (N_3571,N_486,N_2036);
and U3572 (N_3572,N_3224,In_480);
or U3573 (N_3573,In_1608,N_3117);
xnor U3574 (N_3574,N_642,N_3344);
nor U3575 (N_3575,In_2955,N_2702);
xnor U3576 (N_3576,N_503,N_2306);
nand U3577 (N_3577,N_2675,N_3329);
nor U3578 (N_3578,N_1293,In_1503);
or U3579 (N_3579,N_3418,N_3086);
and U3580 (N_3580,N_3496,N_3132);
nor U3581 (N_3581,N_1214,N_3370);
xor U3582 (N_3582,N_3242,N_2904);
nor U3583 (N_3583,In_3343,N_3441);
xnor U3584 (N_3584,N_2874,In_1711);
and U3585 (N_3585,In_4943,N_2195);
and U3586 (N_3586,N_2612,N_3464);
and U3587 (N_3587,In_2007,N_1794);
xnor U3588 (N_3588,N_1912,N_2565);
nand U3589 (N_3589,N_3310,N_1038);
and U3590 (N_3590,In_1256,In_792);
or U3591 (N_3591,N_2899,N_2637);
and U3592 (N_3592,N_1975,N_947);
or U3593 (N_3593,In_3486,N_2744);
xor U3594 (N_3594,In_1368,N_3240);
or U3595 (N_3595,N_3492,N_3423);
nand U3596 (N_3596,In_2684,N_1410);
and U3597 (N_3597,In_900,N_1007);
and U3598 (N_3598,N_3352,N_1551);
and U3599 (N_3599,N_2516,N_2378);
or U3600 (N_3600,In_51,In_4127);
or U3601 (N_3601,N_2909,In_2881);
xor U3602 (N_3602,N_582,In_1657);
xor U3603 (N_3603,N_3255,N_3121);
or U3604 (N_3604,N_1655,N_1756);
and U3605 (N_3605,N_3130,N_666);
and U3606 (N_3606,In_3493,N_2468);
and U3607 (N_3607,N_3489,In_1205);
or U3608 (N_3608,In_4403,N_1134);
or U3609 (N_3609,N_3410,In_698);
nor U3610 (N_3610,N_1935,In_225);
nor U3611 (N_3611,N_2589,In_2641);
and U3612 (N_3612,N_1860,N_755);
or U3613 (N_3613,In_3758,N_572);
or U3614 (N_3614,N_3343,N_2415);
or U3615 (N_3615,In_3540,N_1844);
nor U3616 (N_3616,N_3280,N_3481);
and U3617 (N_3617,N_2459,N_3354);
nor U3618 (N_3618,In_3241,In_275);
xnor U3619 (N_3619,N_2585,N_3384);
nand U3620 (N_3620,N_26,In_4589);
and U3621 (N_3621,N_3035,In_3317);
nand U3622 (N_3622,In_2572,N_2850);
nor U3623 (N_3623,N_2922,N_2118);
nor U3624 (N_3624,N_3164,N_2984);
and U3625 (N_3625,In_1063,N_3052);
and U3626 (N_3626,In_3328,N_1706);
nand U3627 (N_3627,In_4602,In_2172);
and U3628 (N_3628,N_2097,In_1915);
nand U3629 (N_3629,N_2891,In_351);
or U3630 (N_3630,In_2759,N_3428);
nand U3631 (N_3631,N_1228,N_2023);
nor U3632 (N_3632,N_2659,N_274);
xnor U3633 (N_3633,N_187,In_2057);
or U3634 (N_3634,N_250,In_4260);
nor U3635 (N_3635,N_1524,In_3295);
and U3636 (N_3636,N_1117,N_2533);
nor U3637 (N_3637,N_3269,N_2631);
nor U3638 (N_3638,N_2150,N_3479);
xnor U3639 (N_3639,N_356,N_2552);
and U3640 (N_3640,N_3245,In_4434);
nor U3641 (N_3641,N_3045,In_1384);
and U3642 (N_3642,N_3315,N_2839);
or U3643 (N_3643,N_3062,N_3361);
and U3644 (N_3644,N_935,N_3460);
xor U3645 (N_3645,N_2802,N_1624);
and U3646 (N_3646,N_3314,N_3092);
nand U3647 (N_3647,N_2838,In_3038);
and U3648 (N_3648,In_775,N_3435);
nor U3649 (N_3649,N_2881,N_3332);
nor U3650 (N_3650,N_3385,N_2252);
and U3651 (N_3651,N_2748,N_3044);
nor U3652 (N_3652,N_3077,In_510);
nand U3653 (N_3653,N_2507,N_456);
xor U3654 (N_3654,N_3291,In_2908);
and U3655 (N_3655,N_3171,In_4116);
nor U3656 (N_3656,N_1447,In_3259);
nand U3657 (N_3657,N_3005,N_3037);
and U3658 (N_3658,In_1856,In_2909);
and U3659 (N_3659,N_2563,N_2596);
xor U3660 (N_3660,N_2407,N_2914);
nor U3661 (N_3661,N_1774,N_3181);
or U3662 (N_3662,N_3128,N_3375);
nor U3663 (N_3663,N_1318,N_3480);
nand U3664 (N_3664,N_3274,N_2799);
nand U3665 (N_3665,N_787,N_2238);
xor U3666 (N_3666,N_1196,In_692);
or U3667 (N_3667,N_3331,N_2006);
xnor U3668 (N_3668,N_3413,N_3447);
and U3669 (N_3669,N_2085,N_2969);
xor U3670 (N_3670,N_2665,N_1562);
nor U3671 (N_3671,N_1378,In_2421);
and U3672 (N_3672,In_2250,N_3342);
or U3673 (N_3673,In_2160,In_1326);
and U3674 (N_3674,N_2182,N_2936);
nand U3675 (N_3675,In_1577,N_2527);
and U3676 (N_3676,In_2438,N_1149);
nand U3677 (N_3677,N_3210,N_1034);
nand U3678 (N_3678,N_3217,In_726);
and U3679 (N_3679,N_3146,N_3008);
nand U3680 (N_3680,In_3610,In_4159);
and U3681 (N_3681,N_2910,N_963);
nor U3682 (N_3682,In_697,N_1906);
nand U3683 (N_3683,N_1781,N_3194);
nand U3684 (N_3684,N_2859,N_2758);
and U3685 (N_3685,N_2037,N_1060);
xnor U3686 (N_3686,In_3863,N_3474);
nor U3687 (N_3687,In_553,In_4485);
and U3688 (N_3688,N_3311,N_3115);
and U3689 (N_3689,N_2592,N_564);
and U3690 (N_3690,N_2723,N_2888);
and U3691 (N_3691,In_2497,In_3786);
nor U3692 (N_3692,N_609,In_1008);
or U3693 (N_3693,In_2995,N_3182);
nor U3694 (N_3694,N_2835,N_1894);
and U3695 (N_3695,N_2492,N_3293);
xnor U3696 (N_3696,N_2704,N_2190);
nand U3697 (N_3697,N_3134,N_577);
and U3698 (N_3698,In_3217,N_3253);
nand U3699 (N_3699,N_2783,N_3355);
nor U3700 (N_3700,N_1869,N_1646);
or U3701 (N_3701,N_3391,N_3406);
and U3702 (N_3702,N_919,N_3075);
and U3703 (N_3703,N_1413,N_3491);
nor U3704 (N_3704,In_150,N_3101);
nor U3705 (N_3705,N_3249,N_3417);
nor U3706 (N_3706,N_2900,N_3129);
nor U3707 (N_3707,N_1818,In_3995);
and U3708 (N_3708,N_2926,N_1505);
or U3709 (N_3709,In_3928,N_3399);
or U3710 (N_3710,In_1410,In_4880);
xnor U3711 (N_3711,N_237,In_1761);
and U3712 (N_3712,N_1982,In_858);
nor U3713 (N_3713,N_3349,N_3448);
nand U3714 (N_3714,N_12,N_3324);
nor U3715 (N_3715,N_1483,In_4040);
nor U3716 (N_3716,In_1407,In_3340);
and U3717 (N_3717,In_4100,N_3243);
or U3718 (N_3718,N_3022,N_3106);
nor U3719 (N_3719,In_2920,N_1703);
or U3720 (N_3720,N_1438,N_3093);
or U3721 (N_3721,In_2001,N_2761);
nor U3722 (N_3722,N_1509,In_2784);
xor U3723 (N_3723,N_1763,N_3283);
nor U3724 (N_3724,N_2062,N_178);
and U3725 (N_3725,In_4309,In_4978);
and U3726 (N_3726,N_3483,N_3292);
and U3727 (N_3727,N_2801,N_2860);
nor U3728 (N_3728,N_3412,N_3316);
or U3729 (N_3729,N_2937,N_2942);
xor U3730 (N_3730,N_3360,N_587);
nand U3731 (N_3731,N_2960,In_2279);
xor U3732 (N_3732,N_3462,In_2099);
nand U3733 (N_3733,N_2601,In_4347);
and U3734 (N_3734,N_2625,N_1911);
or U3735 (N_3735,N_2828,In_113);
nand U3736 (N_3736,N_3068,N_3411);
or U3737 (N_3737,N_3414,N_2854);
nor U3738 (N_3738,N_2303,In_3339);
or U3739 (N_3739,In_4976,N_2449);
nand U3740 (N_3740,N_3225,In_707);
and U3741 (N_3741,N_2696,N_16);
and U3742 (N_3742,N_3482,N_2778);
nand U3743 (N_3743,In_1861,In_3525);
nand U3744 (N_3744,N_1628,N_974);
or U3745 (N_3745,In_3371,N_2958);
nand U3746 (N_3746,N_3169,In_2820);
nand U3747 (N_3747,N_1209,N_2208);
xor U3748 (N_3748,N_2911,N_3394);
nor U3749 (N_3749,N_3463,N_1257);
xor U3750 (N_3750,N_3282,N_1021);
xnor U3751 (N_3751,N_3434,N_3319);
and U3752 (N_3752,N_3320,N_3614);
xnor U3753 (N_3753,N_2725,N_2580);
nand U3754 (N_3754,N_3275,N_3596);
nand U3755 (N_3755,N_2143,N_2460);
nor U3756 (N_3756,In_1127,N_3671);
and U3757 (N_3757,N_3580,N_2774);
nand U3758 (N_3758,N_3259,N_3189);
nand U3759 (N_3759,N_3145,N_2570);
nor U3760 (N_3760,In_3012,N_2503);
or U3761 (N_3761,N_3570,N_3549);
nand U3762 (N_3762,N_3743,In_1827);
nor U3763 (N_3763,N_3595,N_3472);
xnor U3764 (N_3764,N_2398,N_2706);
nor U3765 (N_3765,In_4929,N_876);
nand U3766 (N_3766,N_3581,N_3263);
nor U3767 (N_3767,N_3054,N_2104);
xnor U3768 (N_3768,In_4058,N_2686);
or U3769 (N_3769,N_3396,N_3350);
and U3770 (N_3770,In_4693,N_3693);
and U3771 (N_3771,In_289,N_3395);
and U3772 (N_3772,N_480,N_2861);
or U3773 (N_3773,N_2931,N_3565);
nand U3774 (N_3774,N_3554,N_2593);
nor U3775 (N_3775,N_3080,N_2988);
xor U3776 (N_3776,In_1506,N_1592);
nor U3777 (N_3777,N_1268,N_3440);
and U3778 (N_3778,N_3325,N_466);
or U3779 (N_3779,N_3744,N_1455);
nand U3780 (N_3780,N_1600,N_3470);
nor U3781 (N_3781,N_3323,In_68);
xor U3782 (N_3782,N_2089,N_2138);
and U3783 (N_3783,N_3535,N_3589);
nand U3784 (N_3784,N_761,N_3525);
xnor U3785 (N_3785,N_2968,N_1806);
xnor U3786 (N_3786,N_3215,N_72);
or U3787 (N_3787,N_115,N_3050);
or U3788 (N_3788,N_3745,N_3422);
or U3789 (N_3789,N_3288,N_3747);
and U3790 (N_3790,In_3911,N_1365);
nor U3791 (N_3791,N_3556,N_2932);
nand U3792 (N_3792,N_3286,In_3908);
nand U3793 (N_3793,N_3456,N_2717);
xor U3794 (N_3794,N_560,N_2733);
and U3795 (N_3795,N_2463,N_2342);
xor U3796 (N_3796,N_2312,N_3662);
and U3797 (N_3797,N_3585,In_4834);
or U3798 (N_3798,N_2864,In_424);
nor U3799 (N_3799,N_2470,N_1858);
nand U3800 (N_3800,N_2447,N_3731);
nor U3801 (N_3801,In_3772,N_3064);
xor U3802 (N_3802,In_2750,N_1803);
nor U3803 (N_3803,N_3330,N_3601);
and U3804 (N_3804,N_265,N_3708);
and U3805 (N_3805,N_3529,N_3557);
xnor U3806 (N_3806,N_1294,N_1155);
or U3807 (N_3807,N_2752,N_3631);
nand U3808 (N_3808,N_1559,N_1752);
nand U3809 (N_3809,N_3138,N_2183);
nand U3810 (N_3810,N_3653,N_1064);
and U3811 (N_3811,N_3099,In_872);
and U3812 (N_3812,N_1501,N_2606);
nor U3813 (N_3813,N_3697,In_4808);
and U3814 (N_3814,N_3124,N_3197);
nor U3815 (N_3815,N_2825,N_326);
and U3816 (N_3816,In_2049,N_2693);
nor U3817 (N_3817,N_2594,N_2309);
xor U3818 (N_3818,N_2441,N_3048);
xnor U3819 (N_3819,In_936,N_3540);
xnor U3820 (N_3820,In_4081,N_3415);
nor U3821 (N_3821,N_2237,N_2947);
and U3822 (N_3822,In_2506,N_2274);
xnor U3823 (N_3823,N_3264,N_1369);
and U3824 (N_3824,N_3537,N_3683);
xor U3825 (N_3825,N_1399,N_2261);
or U3826 (N_3826,In_2082,N_2148);
xnor U3827 (N_3827,N_2763,N_1156);
nand U3828 (N_3828,N_3550,N_3386);
nor U3829 (N_3829,In_1004,N_3664);
and U3830 (N_3830,In_4233,In_2819);
nor U3831 (N_3831,N_3333,N_1790);
nor U3832 (N_3832,N_2137,N_2368);
xnor U3833 (N_3833,N_2328,N_2620);
nand U3834 (N_3834,N_2135,N_3575);
nor U3835 (N_3835,N_3533,N_301);
and U3836 (N_3836,N_3729,N_3738);
xor U3837 (N_3837,N_3000,N_2387);
xnor U3838 (N_3838,In_593,N_518);
nand U3839 (N_3839,N_3446,In_2622);
xor U3840 (N_3840,N_3656,N_3039);
or U3841 (N_3841,In_3727,N_3154);
nand U3842 (N_3842,N_3163,In_2927);
nor U3843 (N_3843,N_3433,In_3253);
or U3844 (N_3844,In_2933,N_2728);
nor U3845 (N_3845,N_3498,N_1545);
or U3846 (N_3846,N_1976,N_3746);
nor U3847 (N_3847,N_3484,In_3044);
or U3848 (N_3848,In_3037,N_3526);
nor U3849 (N_3849,In_1430,In_2307);
and U3850 (N_3850,N_3100,N_3420);
nand U3851 (N_3851,N_3449,In_1598);
xnor U3852 (N_3852,N_1615,N_3004);
xnor U3853 (N_3853,N_3040,N_3239);
xor U3854 (N_3854,N_2959,In_486);
nor U3855 (N_3855,N_2179,N_3612);
nor U3856 (N_3856,In_914,N_1927);
and U3857 (N_3857,N_3487,N_2079);
and U3858 (N_3858,In_2815,In_232);
or U3859 (N_3859,N_3573,In_1981);
nor U3860 (N_3860,N_3478,N_1401);
and U3861 (N_3861,In_4210,N_3032);
xor U3862 (N_3862,N_3444,N_3348);
or U3863 (N_3863,N_2670,N_3393);
xnor U3864 (N_3864,N_2830,In_3971);
xor U3865 (N_3865,N_3590,N_3654);
xnor U3866 (N_3866,In_3167,N_3072);
xnor U3867 (N_3867,N_2882,In_428);
nand U3868 (N_3868,N_3251,N_170);
nand U3869 (N_3869,N_2226,In_260);
nor U3870 (N_3870,N_2141,N_3167);
or U3871 (N_3871,In_1963,N_3615);
nor U3872 (N_3872,In_2064,N_3431);
or U3873 (N_3873,N_731,In_1548);
nor U3874 (N_3874,N_3321,N_3326);
and U3875 (N_3875,In_2736,N_2433);
or U3876 (N_3876,In_151,N_2865);
and U3877 (N_3877,N_3684,N_3740);
nand U3878 (N_3878,In_2888,N_2709);
or U3879 (N_3879,N_1598,N_3445);
xnor U3880 (N_3880,N_1198,N_3467);
or U3881 (N_3881,In_2958,N_1824);
or U3882 (N_3882,N_3598,N_1537);
and U3883 (N_3883,N_3430,N_3158);
nand U3884 (N_3884,N_3735,N_3584);
or U3885 (N_3885,N_3076,N_2431);
and U3886 (N_3886,N_2727,N_2364);
nor U3887 (N_3887,N_3469,N_3454);
and U3888 (N_3888,N_3543,In_602);
xor U3889 (N_3889,N_3207,N_3670);
and U3890 (N_3890,N_3102,N_3357);
nand U3891 (N_3891,N_1480,N_3028);
nor U3892 (N_3892,N_2841,N_3453);
xnor U3893 (N_3893,In_1488,In_253);
and U3894 (N_3894,In_3067,N_2650);
and U3895 (N_3895,N_2549,N_3301);
or U3896 (N_3896,N_1811,N_2741);
nand U3897 (N_3897,N_2521,N_2990);
xnor U3898 (N_3898,In_2375,In_3160);
nand U3899 (N_3899,N_2722,In_663);
xor U3900 (N_3900,N_3450,N_3551);
or U3901 (N_3901,N_3688,In_1023);
nand U3902 (N_3902,N_3734,N_2508);
and U3903 (N_3903,N_2408,N_1291);
xor U3904 (N_3904,N_2901,N_2903);
and U3905 (N_3905,In_3414,N_1913);
nand U3906 (N_3906,In_2762,N_613);
xor U3907 (N_3907,N_3667,N_3150);
nand U3908 (N_3908,In_4188,N_2955);
nor U3909 (N_3909,N_2803,N_2636);
or U3910 (N_3910,N_3622,N_1822);
nor U3911 (N_3911,In_758,N_3295);
nand U3912 (N_3912,In_1689,N_1175);
xnor U3913 (N_3913,In_1885,In_1119);
xnor U3914 (N_3914,N_3250,N_2578);
and U3915 (N_3915,N_3109,N_3675);
and U3916 (N_3916,N_116,N_2232);
and U3917 (N_3917,N_3685,N_3698);
nor U3918 (N_3918,N_3439,N_3328);
nand U3919 (N_3919,N_1596,N_3365);
xor U3920 (N_3920,In_1284,In_2021);
nand U3921 (N_3921,N_2409,N_1830);
and U3922 (N_3922,N_3403,N_3436);
or U3923 (N_3923,N_3476,N_2600);
and U3924 (N_3924,N_1105,N_3730);
nand U3925 (N_3925,N_3504,N_1036);
nor U3926 (N_3926,N_3644,N_3659);
and U3927 (N_3927,N_3680,N_2889);
or U3928 (N_3928,N_2979,N_3652);
nor U3929 (N_3929,N_1492,N_1952);
xor U3930 (N_3930,N_3732,N_3212);
nor U3931 (N_3931,N_3058,N_3669);
nand U3932 (N_3932,In_2293,In_513);
or U3933 (N_3933,N_2056,N_248);
or U3934 (N_3934,N_3600,In_1716);
xnor U3935 (N_3935,N_2245,N_3466);
nor U3936 (N_3936,N_1987,N_3214);
or U3937 (N_3937,N_457,N_3218);
nand U3938 (N_3938,N_3630,N_1676);
nor U3939 (N_3939,N_3682,N_1632);
or U3940 (N_3940,N_2502,In_1966);
or U3941 (N_3941,In_4362,N_3539);
nor U3942 (N_3942,N_1227,N_2658);
and U3943 (N_3943,N_2299,In_265);
nor U3944 (N_3944,N_404,In_3661);
xnor U3945 (N_3945,N_2886,In_1125);
or U3946 (N_3946,In_846,N_1877);
or U3947 (N_3947,N_2688,N_3103);
or U3948 (N_3948,In_1549,In_2207);
and U3949 (N_3949,N_2972,N_2504);
and U3950 (N_3950,In_1408,In_4652);
nand U3951 (N_3951,N_3553,In_2449);
or U3952 (N_3952,In_337,N_2893);
xnor U3953 (N_3953,N_2999,N_2455);
or U3954 (N_3954,In_3797,N_2490);
or U3955 (N_3955,N_3628,N_3090);
nand U3956 (N_3956,N_3082,N_2866);
or U3957 (N_3957,N_2427,In_3573);
nand U3958 (N_3958,N_2291,N_3299);
xnor U3959 (N_3959,N_993,In_3773);
nor U3960 (N_3960,N_3419,N_3180);
nand U3961 (N_3961,N_2821,In_4611);
and U3962 (N_3962,In_3563,N_2856);
xor U3963 (N_3963,In_2817,In_2409);
xnor U3964 (N_3964,In_2236,N_3503);
xnor U3965 (N_3965,N_3648,N_3302);
nor U3966 (N_3966,N_3019,N_3562);
or U3967 (N_3967,N_3364,N_3340);
nand U3968 (N_3968,N_2867,N_3571);
or U3969 (N_3969,N_1099,In_3769);
nand U3970 (N_3970,In_1964,N_3468);
nor U3971 (N_3971,N_3136,In_3078);
and U3972 (N_3972,N_119,N_3629);
and U3973 (N_3973,N_512,In_1882);
or U3974 (N_3974,N_3610,N_2209);
or U3975 (N_3975,N_3170,N_2734);
nor U3976 (N_3976,In_2222,N_3704);
nand U3977 (N_3977,N_424,N_3351);
nand U3978 (N_3978,In_925,In_4503);
nor U3979 (N_3979,N_1981,In_3127);
or U3980 (N_3980,N_3692,In_4512);
or U3981 (N_3981,N_3520,N_1826);
or U3982 (N_3982,N_3710,N_3131);
xor U3983 (N_3983,N_3377,N_3307);
nor U3984 (N_3984,N_2870,N_3741);
and U3985 (N_3985,In_4063,N_1832);
or U3986 (N_3986,In_4959,N_2746);
nor U3987 (N_3987,In_1534,N_2742);
or U3988 (N_3988,N_3527,N_3204);
xnor U3989 (N_3989,N_2480,N_3651);
nor U3990 (N_3990,N_3238,N_3308);
nor U3991 (N_3991,In_450,N_3513);
nand U3992 (N_3992,N_3289,N_3192);
and U3993 (N_3993,N_1603,N_2884);
and U3994 (N_3994,N_3638,N_2843);
and U3995 (N_3995,N_3721,N_3356);
and U3996 (N_3996,N_1555,In_2928);
xnor U3997 (N_3997,N_1932,N_3530);
or U3998 (N_3998,In_1274,In_3302);
nor U3999 (N_3999,In_3359,N_3566);
nor U4000 (N_4000,N_3716,N_3711);
nor U4001 (N_4001,N_3947,N_3392);
or U4002 (N_4002,N_3998,N_2685);
nor U4003 (N_4003,N_3416,In_2430);
or U4004 (N_4004,N_3193,N_2106);
xnor U4005 (N_4005,N_3826,N_3661);
or U4006 (N_4006,N_3785,N_3208);
nand U4007 (N_4007,N_3223,N_3398);
nor U4008 (N_4008,N_2124,N_3913);
nor U4009 (N_4009,N_255,N_3376);
xnor U4010 (N_4010,N_2511,N_2731);
and U4011 (N_4011,N_3975,In_3378);
and U4012 (N_4012,N_3719,N_3860);
nor U4013 (N_4013,In_3912,N_3854);
and U4014 (N_4014,In_4015,N_3763);
nand U4015 (N_4015,N_2055,N_2832);
nor U4016 (N_4016,N_2906,N_2697);
and U4017 (N_4017,In_3075,In_4326);
nor U4018 (N_4018,N_3865,N_3781);
and U4019 (N_4019,N_2666,N_3679);
xnor U4020 (N_4020,N_2844,N_2754);
nand U4021 (N_4021,N_3750,In_4999);
nand U4022 (N_4022,N_3296,N_1115);
xnor U4023 (N_4023,N_3905,N_3791);
and U4024 (N_4024,N_2711,N_3512);
xor U4025 (N_4025,N_3727,N_3899);
nor U4026 (N_4026,In_2871,N_3786);
xor U4027 (N_4027,N_3953,N_1833);
xor U4028 (N_4028,N_3852,N_3620);
and U4029 (N_4029,N_3185,In_2030);
xnor U4030 (N_4030,N_3126,N_1461);
xnor U4031 (N_4031,N_949,N_3971);
nand U4032 (N_4032,N_3819,N_3896);
nor U4033 (N_4033,N_2965,N_2446);
xnor U4034 (N_4034,N_3770,N_3985);
or U4035 (N_4035,N_2943,N_2971);
nor U4036 (N_4036,N_3458,N_3867);
nor U4037 (N_4037,N_3148,N_3455);
nor U4038 (N_4038,N_3043,N_3800);
or U4039 (N_4039,N_3924,N_3339);
xnor U4040 (N_4040,In_3474,N_3567);
and U4041 (N_4041,N_1581,N_3771);
xnor U4042 (N_4042,N_3510,N_3338);
nand U4043 (N_4043,N_1871,In_2616);
or U4044 (N_4044,In_3013,In_2894);
nor U4045 (N_4045,N_3929,N_120);
nand U4046 (N_4046,N_3228,N_3609);
nand U4047 (N_4047,N_264,N_3666);
nand U4048 (N_4048,N_3616,N_2477);
or U4049 (N_4049,N_1051,N_3756);
and U4050 (N_4050,N_3806,N_3774);
or U4051 (N_4051,In_2672,N_3303);
nand U4052 (N_4052,N_3912,In_266);
or U4053 (N_4053,N_3816,N_3502);
xor U4054 (N_4054,N_3877,N_2586);
nand U4055 (N_4055,N_3932,N_1959);
or U4056 (N_4056,N_3650,N_3546);
nor U4057 (N_4057,N_3804,N_3911);
or U4058 (N_4058,In_4856,N_3948);
nand U4059 (N_4059,In_2893,N_3421);
and U4060 (N_4060,N_3373,N_3663);
and U4061 (N_4061,N_3936,N_3026);
xor U4062 (N_4062,N_3424,N_2951);
nor U4063 (N_4063,N_3964,N_3665);
or U4064 (N_4064,N_2219,In_4727);
and U4065 (N_4065,N_3888,N_3277);
or U4066 (N_4066,N_2465,In_774);
nor U4067 (N_4067,N_2684,N_2307);
and U4068 (N_4068,N_3946,N_2869);
nand U4069 (N_4069,In_631,N_1231);
nand U4070 (N_4070,N_3972,N_3970);
or U4071 (N_4071,In_2938,N_3849);
nand U4072 (N_4072,N_643,N_3313);
xnor U4073 (N_4073,N_3260,N_1636);
nor U4074 (N_4074,N_2966,N_2168);
and U4075 (N_4075,N_3891,N_3488);
nand U4076 (N_4076,N_3893,N_3694);
nand U4077 (N_4077,N_3262,N_3801);
nor U4078 (N_4078,N_2211,N_1828);
xnor U4079 (N_4079,N_3751,N_1113);
nand U4080 (N_4080,N_714,N_3830);
xor U4081 (N_4081,N_3718,N_3276);
or U4082 (N_4082,N_3400,N_3634);
or U4083 (N_4083,N_1382,N_3625);
and U4084 (N_4084,N_3815,N_3495);
nor U4085 (N_4085,N_3833,N_971);
and U4086 (N_4086,N_1050,N_3011);
nand U4087 (N_4087,N_2320,N_3853);
or U4088 (N_4088,N_3805,N_3894);
nor U4089 (N_4089,N_3459,In_4850);
nor U4090 (N_4090,N_3592,N_3908);
nand U4091 (N_4091,N_1607,N_3676);
or U4092 (N_4092,In_1280,N_2787);
xnor U4093 (N_4093,N_3824,N_3465);
nor U4094 (N_4094,N_1892,N_3882);
nand U4095 (N_4095,N_3544,N_3937);
and U4096 (N_4096,N_890,N_2669);
and U4097 (N_4097,N_390,N_2766);
nor U4098 (N_4098,In_2259,In_1557);
and U4099 (N_4099,N_3817,N_790);
nor U4100 (N_4100,N_3358,In_1361);
nor U4101 (N_4101,N_3792,N_3950);
or U4102 (N_4102,In_727,N_427);
nand U4103 (N_4103,N_3397,N_2356);
xnor U4104 (N_4104,In_127,N_3831);
or U4105 (N_4105,N_3880,N_3569);
xor U4106 (N_4106,N_3524,N_3020);
nand U4107 (N_4107,N_3754,N_3368);
xnor U4108 (N_4108,N_2556,N_3607);
nor U4109 (N_4109,N_2491,In_2749);
nor U4110 (N_4110,N_3935,N_2797);
xor U4111 (N_4111,N_3968,N_483);
nand U4112 (N_4112,N_1755,N_3722);
or U4113 (N_4113,N_1955,N_444);
or U4114 (N_4114,N_3505,N_3956);
or U4115 (N_4115,N_3139,N_3933);
nand U4116 (N_4116,N_3969,In_3321);
and U4117 (N_4117,N_1200,N_3013);
and U4118 (N_4118,N_3532,N_3921);
or U4119 (N_4119,N_3752,N_3982);
or U4120 (N_4120,N_2174,N_3823);
xnor U4121 (N_4121,N_2519,N_3157);
nand U4122 (N_4122,N_1886,N_2139);
and U4123 (N_4123,N_3096,N_1353);
and U4124 (N_4124,N_3611,N_3989);
xor U4125 (N_4125,In_1944,N_3152);
nand U4126 (N_4126,N_3645,N_3978);
and U4127 (N_4127,In_1664,N_3673);
or U4128 (N_4128,N_3885,N_3973);
nand U4129 (N_4129,In_2257,In_3716);
nor U4130 (N_4130,N_3900,N_3983);
xor U4131 (N_4131,N_3827,N_3690);
nand U4132 (N_4132,N_3962,In_1892);
and U4133 (N_4133,N_827,N_2579);
and U4134 (N_4134,In_1278,N_3720);
nand U4135 (N_4135,N_3235,N_3383);
nor U4136 (N_4136,N_2680,In_3948);
nor U4137 (N_4137,N_3739,N_2493);
or U4138 (N_4138,N_3067,N_2887);
nand U4139 (N_4139,N_3926,In_1812);
and U4140 (N_4140,N_3790,N_3374);
and U4141 (N_4141,N_3712,N_3545);
xnor U4142 (N_4142,N_1071,N_3033);
xnor U4143 (N_4143,N_3534,N_3382);
or U4144 (N_4144,N_3749,N_3618);
nor U4145 (N_4145,N_3681,N_3828);
nand U4146 (N_4146,N_2009,N_298);
nor U4147 (N_4147,N_3065,N_3266);
nor U4148 (N_4148,N_3797,N_3576);
nor U4149 (N_4149,N_3346,In_2079);
nand U4150 (N_4150,N_2126,N_3347);
xor U4151 (N_4151,In_3182,In_4410);
and U4152 (N_4152,N_3273,In_945);
nand U4153 (N_4153,N_3787,N_3778);
xor U4154 (N_4154,N_3390,In_3265);
nor U4155 (N_4155,N_3977,In_2754);
or U4156 (N_4156,N_2896,N_3372);
and U4157 (N_4157,N_2316,N_3270);
xnor U4158 (N_4158,N_3285,N_1993);
nand U4159 (N_4159,N_2806,N_1041);
xnor U4160 (N_4160,N_3563,N_3070);
nand U4161 (N_4161,N_3162,In_1264);
nor U4162 (N_4162,N_3760,N_3918);
and U4163 (N_4163,N_1248,N_2522);
and U4164 (N_4164,N_3999,N_2982);
nor U4165 (N_4165,N_2518,N_3335);
xnor U4166 (N_4166,N_929,N_3706);
nor U4167 (N_4167,N_3427,In_3762);
and U4168 (N_4168,N_2363,In_1461);
xor U4169 (N_4169,N_2327,N_3602);
xor U4170 (N_4170,In_4799,N_3876);
or U4171 (N_4171,N_3516,In_2788);
nor U4172 (N_4172,In_4536,N_3736);
and U4173 (N_4173,N_3125,N_3265);
or U4174 (N_4174,N_3794,N_3137);
xor U4175 (N_4175,N_3572,In_863);
nand U4176 (N_4176,N_3840,N_3247);
or U4177 (N_4177,N_3940,N_3254);
and U4178 (N_4178,N_3564,N_1619);
nor U4179 (N_4179,In_4464,In_1316);
nor U4180 (N_4180,N_3930,In_4195);
nand U4181 (N_4181,N_2571,N_1088);
nand U4182 (N_4182,N_2890,N_3901);
nor U4183 (N_4183,In_4587,N_831);
and U4184 (N_4184,N_2297,In_3269);
and U4185 (N_4185,N_2412,N_970);
or U4186 (N_4186,N_3642,N_1917);
xor U4187 (N_4187,N_3892,N_3294);
or U4188 (N_4188,N_1881,N_3429);
nor U4189 (N_4189,N_1069,N_3069);
or U4190 (N_4190,N_1810,N_2789);
or U4191 (N_4191,N_1711,N_3726);
or U4192 (N_4192,N_3870,N_3388);
and U4193 (N_4193,In_3102,N_3775);
or U4194 (N_4194,N_3443,N_233);
or U4195 (N_4195,N_3757,N_2573);
or U4196 (N_4196,N_2275,N_2641);
xnor U4197 (N_4197,N_2822,N_3588);
nor U4198 (N_4198,N_3003,N_343);
and U4199 (N_4199,N_3845,N_3107);
nor U4200 (N_4200,N_2705,N_3219);
nor U4201 (N_4201,N_3761,N_3869);
and U4202 (N_4202,N_3910,N_3574);
or U4203 (N_4203,In_3538,N_2842);
nor U4204 (N_4204,In_2883,N_1883);
xnor U4205 (N_4205,N_2712,N_3737);
nor U4206 (N_4206,N_3110,N_2286);
nand U4207 (N_4207,N_3379,N_3635);
nand U4208 (N_4208,N_1276,In_643);
xor U4209 (N_4209,N_110,In_830);
xor U4210 (N_4210,N_3639,N_1739);
or U4211 (N_4211,N_2831,N_3281);
and U4212 (N_4212,N_2462,N_3897);
and U4213 (N_4213,N_2084,N_3965);
nand U4214 (N_4214,N_3511,N_2253);
and U4215 (N_4215,N_2941,N_1821);
and U4216 (N_4216,N_3733,In_3440);
nor U4217 (N_4217,In_3353,N_3007);
and U4218 (N_4218,In_3497,N_869);
and U4219 (N_4219,In_3464,In_2967);
nand U4220 (N_4220,N_2777,N_3141);
nor U4221 (N_4221,N_3624,N_3604);
nand U4222 (N_4222,N_3471,N_3902);
and U4223 (N_4223,N_3232,N_3886);
or U4224 (N_4224,In_4145,In_1769);
xnor U4225 (N_4225,N_1281,N_3808);
xor U4226 (N_4226,N_1130,N_3278);
nand U4227 (N_4227,N_3874,In_3566);
xnor U4228 (N_4228,N_799,N_13);
nand U4229 (N_4229,N_3568,N_1635);
xor U4230 (N_4230,N_3098,In_461);
xor U4231 (N_4231,N_3599,N_87);
and U4232 (N_4232,In_1928,N_2716);
or U4233 (N_4233,N_1984,N_2264);
nand U4234 (N_4234,N_2621,N_2543);
xnor U4235 (N_4235,N_3234,N_1513);
or U4236 (N_4236,N_3988,N_2397);
xnor U4237 (N_4237,N_421,In_3221);
nand U4238 (N_4238,N_3856,N_3198);
xor U4239 (N_4239,N_3859,In_3510);
and U4240 (N_4240,N_3767,N_3820);
xor U4241 (N_4241,N_3784,N_3773);
nand U4242 (N_4242,N_3941,N_3895);
nand U4243 (N_4243,N_2461,N_3759);
or U4244 (N_4244,N_2469,N_3724);
xnor U4245 (N_4245,N_3779,N_3660);
and U4246 (N_4246,N_3916,N_3818);
xnor U4247 (N_4247,N_3906,N_3821);
nor U4248 (N_4248,N_835,N_3623);
or U4249 (N_4249,N_3637,N_3814);
nor U4250 (N_4250,N_3955,N_3674);
nor U4251 (N_4251,N_4245,N_3258);
xor U4252 (N_4252,N_2196,N_3409);
xor U4253 (N_4253,N_3961,N_3705);
nor U4254 (N_4254,In_4511,N_3810);
xor U4255 (N_4255,N_4196,N_4244);
nor U4256 (N_4256,N_3188,N_3837);
nor U4257 (N_4257,N_3851,N_4111);
nor U4258 (N_4258,N_4002,In_2095);
xor U4259 (N_4259,N_3279,N_4210);
or U4260 (N_4260,N_2584,N_3871);
xor U4261 (N_4261,N_4243,N_1422);
or U4262 (N_4262,N_3515,N_3490);
and U4263 (N_4263,In_2038,N_2001);
nand U4264 (N_4264,In_2490,N_3838);
nand U4265 (N_4265,N_4107,N_3485);
and U4266 (N_4266,N_3015,N_3994);
nor U4267 (N_4267,N_3945,N_4167);
nor U4268 (N_4268,N_3508,N_3306);
and U4269 (N_4269,N_1761,N_4033);
nand U4270 (N_4270,N_873,N_3160);
or U4271 (N_4271,N_4089,N_1813);
and U4272 (N_4272,N_4074,In_117);
nor U4273 (N_4273,N_2269,N_3559);
or U4274 (N_4274,N_4077,N_4224);
and U4275 (N_4275,N_3312,N_3500);
nand U4276 (N_4276,N_3687,N_4104);
nor U4277 (N_4277,N_3617,In_3937);
xnor U4278 (N_4278,N_4072,N_4075);
nand U4279 (N_4279,N_4133,N_4202);
and U4280 (N_4280,N_3016,N_4218);
nand U4281 (N_4281,N_2753,N_3668);
and U4282 (N_4282,N_3586,N_3327);
or U4283 (N_4283,N_4031,N_4180);
or U4284 (N_4284,N_3887,In_948);
nand U4285 (N_4285,N_3552,N_3879);
nor U4286 (N_4286,N_4005,N_973);
and U4287 (N_4287,N_4053,N_4145);
xor U4288 (N_4288,N_4010,N_4050);
xor U4289 (N_4289,N_3772,N_3812);
xor U4290 (N_4290,N_3031,N_3858);
or U4291 (N_4291,N_4149,N_1719);
nand U4292 (N_4292,N_3621,N_3825);
or U4293 (N_4293,N_4222,N_2241);
nand U4294 (N_4294,N_4115,N_3560);
or U4295 (N_4295,N_4082,N_3848);
and U4296 (N_4296,N_4187,N_4161);
and U4297 (N_4297,N_2720,In_95);
xnor U4298 (N_4298,In_1475,N_85);
nand U4299 (N_4299,In_1057,N_3714);
xor U4300 (N_4300,N_4169,N_3725);
nand U4301 (N_4301,N_3864,N_2767);
nor U4302 (N_4302,N_3178,N_3834);
or U4303 (N_4303,N_3451,N_4143);
or U4304 (N_4304,N_3796,N_4141);
xor U4305 (N_4305,N_3802,N_4012);
nor U4306 (N_4306,N_4013,N_3021);
nor U4307 (N_4307,N_4153,N_4108);
nor U4308 (N_4308,N_3993,N_4027);
nor U4309 (N_4309,N_3378,N_4015);
xor U4310 (N_4310,N_3613,N_594);
and U4311 (N_4311,N_4123,In_2225);
xnor U4312 (N_4312,N_3060,N_2695);
or U4313 (N_4313,N_3140,N_3872);
xnor U4314 (N_4314,N_4212,N_2961);
or U4315 (N_4315,N_1933,In_3851);
nor U4316 (N_4316,N_3658,N_3996);
nor U4317 (N_4317,N_3919,N_3934);
xnor U4318 (N_4318,N_4201,In_4665);
and U4319 (N_4319,N_3813,In_3825);
or U4320 (N_4320,N_4207,In_1691);
nand U4321 (N_4321,N_4247,N_3012);
nor U4322 (N_4322,N_3768,N_4231);
nand U4323 (N_4323,N_3531,N_3541);
nor U4324 (N_4324,N_2539,N_1499);
xor U4325 (N_4325,N_3287,N_3976);
xor U4326 (N_4326,N_4152,N_3855);
or U4327 (N_4327,N_3881,N_3700);
and U4328 (N_4328,N_3678,In_1589);
xnor U4329 (N_4329,N_4188,N_1260);
nand U4330 (N_4330,N_4030,N_4094);
nor U4331 (N_4331,N_3769,N_4131);
nor U4332 (N_4332,N_3071,In_1286);
xor U4333 (N_4333,N_2935,N_3389);
and U4334 (N_4334,N_3846,In_3282);
nand U4335 (N_4335,N_3555,N_3780);
nand U4336 (N_4336,N_3873,N_4175);
nand U4337 (N_4337,N_4211,N_3997);
nand U4338 (N_4338,N_3408,N_3960);
nand U4339 (N_4339,N_3857,N_2776);
nand U4340 (N_4340,In_3309,In_1235);
nor U4341 (N_4341,N_3649,N_1054);
xor U4342 (N_4342,N_3261,N_3728);
nor U4343 (N_4343,N_4019,N_4116);
nor U4344 (N_4344,N_2454,In_1643);
nor U4345 (N_4345,N_3558,N_3271);
or U4346 (N_4346,N_3702,N_4138);
nor U4347 (N_4347,In_2042,N_1139);
nor U4348 (N_4348,In_1288,N_3519);
and U4349 (N_4349,N_3438,N_4093);
xor U4350 (N_4350,N_3799,N_4037);
nand U4351 (N_4351,N_4217,In_1750);
nand U4352 (N_4352,N_4226,N_3795);
xor U4353 (N_4353,N_3974,N_4197);
nand U4354 (N_4354,In_1563,N_4129);
or U4355 (N_4355,N_3925,N_3889);
and U4356 (N_4356,N_4199,N_1572);
xor U4357 (N_4357,N_2088,N_2557);
xnor U4358 (N_4358,In_2946,N_4214);
and U4359 (N_4359,N_4183,N_3514);
or U4360 (N_4360,In_3392,N_3672);
nor U4361 (N_4361,N_9,N_3939);
or U4362 (N_4362,N_2970,N_4213);
xnor U4363 (N_4363,N_3709,N_4192);
or U4364 (N_4364,N_2682,N_3230);
or U4365 (N_4365,N_3183,N_4008);
xnor U4366 (N_4366,N_4163,N_4184);
nand U4367 (N_4367,N_4101,N_3951);
or U4368 (N_4368,N_3715,In_3615);
and U4369 (N_4369,N_4102,N_3822);
xor U4370 (N_4370,N_3984,N_3890);
and U4371 (N_4371,N_3432,N_3923);
xnor U4372 (N_4372,N_3765,N_4092);
nand U4373 (N_4373,N_4024,In_747);
nor U4374 (N_4374,N_2476,N_4110);
xor U4375 (N_4375,N_3943,In_4085);
or U4376 (N_4376,N_4018,N_1340);
xor U4377 (N_4377,N_2846,N_4173);
nor U4378 (N_4378,N_4181,N_4017);
xor U4379 (N_4379,N_3863,N_4109);
nand U4380 (N_4380,N_2715,N_3367);
nand U4381 (N_4381,N_4087,N_4204);
and U4382 (N_4382,N_3336,N_4228);
or U4383 (N_4383,N_1939,In_3514);
nor U4384 (N_4384,N_3542,N_547);
or U4385 (N_4385,N_4172,In_3942);
nor U4386 (N_4386,N_3807,N_3334);
and U4387 (N_4387,In_1040,N_2288);
nor U4388 (N_4388,N_883,N_4157);
and U4389 (N_4389,N_4240,In_2632);
nand U4390 (N_4390,N_4233,N_2142);
nor U4391 (N_4391,In_1972,N_2820);
nand U4392 (N_4392,N_3457,N_4190);
and U4393 (N_4393,N_3371,N_4047);
or U4394 (N_4394,N_3963,N_2259);
or U4395 (N_4395,N_4126,N_1498);
nor U4396 (N_4396,N_757,N_3696);
and U4397 (N_4397,N_2529,N_3928);
nor U4398 (N_4398,N_3120,N_4071);
xor U4399 (N_4399,N_4043,N_4156);
nor U4400 (N_4400,N_4191,N_3699);
nand U4401 (N_4401,N_818,N_3832);
xnor U4402 (N_4402,N_1854,N_4219);
or U4403 (N_4403,N_3753,N_3497);
xor U4404 (N_4404,In_1743,N_4113);
xor U4405 (N_4405,N_877,N_4230);
xor U4406 (N_4406,N_3583,In_3730);
nand U4407 (N_4407,N_1485,N_2976);
xor U4408 (N_4408,N_4195,N_4070);
nand U4409 (N_4409,N_3636,N_3633);
nand U4410 (N_4410,N_3297,N_4080);
or U4411 (N_4411,N_3341,N_3842);
and U4412 (N_4412,N_3593,N_4147);
or U4413 (N_4413,N_2755,N_4114);
nor U4414 (N_4414,N_3764,N_3957);
and U4415 (N_4415,N_4068,N_4121);
nor U4416 (N_4416,N_3522,N_3104);
xnor U4417 (N_4417,N_3755,N_840);
or U4418 (N_4418,N_3655,N_3835);
nor U4419 (N_4419,N_2768,N_4215);
or U4420 (N_4420,N_2989,N_3944);
xor U4421 (N_4421,In_819,N_1588);
or U4422 (N_4422,N_3844,N_3300);
or U4423 (N_4423,N_3591,N_1882);
or U4424 (N_4424,N_4160,N_3494);
nor U4425 (N_4425,N_4176,N_4132);
or U4426 (N_4426,N_2930,N_4165);
and U4427 (N_4427,N_3594,N_4038);
nand U4428 (N_4428,N_4146,N_4248);
nand U4429 (N_4429,N_4136,N_4054);
or U4430 (N_4430,N_1610,N_4016);
xnor U4431 (N_4431,N_3322,N_4249);
or U4432 (N_4432,N_3904,N_3345);
nor U4433 (N_4433,In_2984,N_4032);
or U4434 (N_4434,N_3723,N_3987);
or U4435 (N_4435,N_3967,N_3548);
nand U4436 (N_4436,In_4225,N_3713);
and U4437 (N_4437,N_3561,N_1736);
nor U4438 (N_4438,N_1699,N_4223);
xor U4439 (N_4439,N_4118,N_3861);
or U4440 (N_4440,N_196,In_3007);
nor U4441 (N_4441,In_195,N_3862);
nor U4442 (N_4442,N_1085,N_4021);
xnor U4443 (N_4443,N_2057,N_2495);
or U4444 (N_4444,In_3064,N_2987);
nor U4445 (N_4445,N_4225,N_4220);
nand U4446 (N_4446,N_3798,N_2824);
xor U4447 (N_4447,N_1728,N_4229);
and U4448 (N_4448,N_4242,N_3811);
nor U4449 (N_4449,N_3353,In_3089);
or U4450 (N_4450,N_3954,N_4091);
nor U4451 (N_4451,In_3284,N_4142);
nor U4452 (N_4452,N_3493,N_3748);
xor U4453 (N_4453,N_4186,N_4059);
nand U4454 (N_4454,N_3405,N_3579);
xor U4455 (N_4455,N_2376,N_3147);
and U4456 (N_4456,N_3362,N_2032);
nor U4457 (N_4457,N_3587,In_1440);
and U4458 (N_4458,N_3742,N_3528);
nor U4459 (N_4459,N_4079,N_3305);
nand U4460 (N_4460,N_4127,N_4023);
and U4461 (N_4461,N_3836,N_2063);
nand U4462 (N_4462,N_4064,N_4200);
xnor U4463 (N_4463,N_3707,N_3547);
and U4464 (N_4464,N_3875,N_4083);
or U4465 (N_4465,N_3605,N_3619);
or U4466 (N_4466,N_1638,N_4097);
and U4467 (N_4467,N_1764,In_1905);
and U4468 (N_4468,N_3536,N_4189);
xor U4469 (N_4469,N_3758,N_3473);
and U4470 (N_4470,In_3882,N_4099);
and U4471 (N_4471,N_4168,N_3627);
or U4472 (N_4472,In_1575,N_4103);
or U4473 (N_4473,N_4216,N_3884);
or U4474 (N_4474,N_3632,N_4177);
nand U4475 (N_4475,N_3920,N_4178);
nand U4476 (N_4476,N_2653,N_4117);
xor U4477 (N_4477,N_3788,N_4105);
nor U4478 (N_4478,In_346,N_3782);
and U4479 (N_4479,N_3309,N_4193);
nand U4480 (N_4480,N_4159,N_2769);
nand U4481 (N_4481,N_4001,N_3387);
nand U4482 (N_4482,N_2939,N_3268);
xnor U4483 (N_4483,N_4124,N_4198);
nor U4484 (N_4484,N_3626,N_563);
xor U4485 (N_4485,N_3907,N_4206);
nor U4486 (N_4486,N_3931,N_4048);
and U4487 (N_4487,N_2729,N_3922);
xnor U4488 (N_4488,N_4166,N_3657);
and U4489 (N_4489,N_2661,In_2477);
or U4490 (N_4490,N_4006,N_1618);
nand U4491 (N_4491,N_1698,In_1873);
or U4492 (N_4492,N_4085,N_4234);
nor U4493 (N_4493,N_2206,N_4150);
and U4494 (N_4494,N_3981,In_1886);
nand U4495 (N_4495,N_1121,N_527);
and U4496 (N_4496,N_4020,N_4046);
or U4497 (N_4497,N_3917,N_3992);
and U4498 (N_4498,N_4236,N_2058);
nand U4499 (N_4499,N_4063,N_4022);
or U4500 (N_4500,N_4269,N_4261);
and U4501 (N_4501,N_4493,N_4360);
and U4502 (N_4502,In_2124,N_4443);
or U4503 (N_4503,N_4235,In_4338);
nor U4504 (N_4504,N_4339,N_4460);
or U4505 (N_4505,N_4291,N_4462);
xor U4506 (N_4506,N_4406,N_4473);
nand U4507 (N_4507,N_4492,N_4058);
or U4508 (N_4508,N_4039,N_4425);
and U4509 (N_4509,N_4076,N_4065);
or U4510 (N_4510,N_4349,N_3995);
nor U4511 (N_4511,N_4441,N_4487);
and U4512 (N_4512,N_4351,In_4913);
xor U4513 (N_4513,N_4467,N_4363);
nand U4514 (N_4514,N_3695,N_4403);
and U4515 (N_4515,N_3517,N_4140);
nand U4516 (N_4516,N_1272,In_4963);
and U4517 (N_4517,N_3766,N_4447);
nand U4518 (N_4518,N_4250,N_4232);
nand U4519 (N_4519,N_4432,N_4321);
nor U4520 (N_4520,N_3641,N_4237);
and U4521 (N_4521,N_4098,N_4426);
nand U4522 (N_4522,N_4292,N_4424);
nor U4523 (N_4523,N_4313,N_4434);
nor U4524 (N_4524,N_3578,N_4011);
xor U4525 (N_4525,N_1082,N_4128);
xnor U4526 (N_4526,N_4182,N_4411);
nor U4527 (N_4527,N_4325,N_4276);
nand U4528 (N_4528,N_3990,N_4435);
and U4529 (N_4529,N_4045,N_4328);
and U4530 (N_4530,N_126,N_4372);
nand U4531 (N_4531,N_4284,N_4084);
or U4532 (N_4532,N_4439,N_3640);
nor U4533 (N_4533,N_4436,N_4446);
and U4534 (N_4534,N_4170,N_4049);
and U4535 (N_4535,N_3878,N_4055);
nand U4536 (N_4536,N_4307,In_757);
or U4537 (N_4537,N_4451,N_4297);
or U4538 (N_4538,N_4371,N_3461);
nand U4539 (N_4539,N_2640,N_3647);
nor U4540 (N_4540,N_3538,N_4352);
nand U4541 (N_4541,N_4334,N_4489);
nand U4542 (N_4542,N_997,N_3116);
or U4543 (N_4543,N_4450,N_4042);
and U4544 (N_4544,N_3298,N_4060);
and U4545 (N_4545,N_4026,N_4322);
or U4546 (N_4546,N_3717,N_4278);
nand U4547 (N_4547,N_4442,N_3047);
nand U4548 (N_4548,N_4366,N_1957);
and U4549 (N_4549,N_3190,N_2868);
and U4550 (N_4550,N_4100,N_4056);
nand U4551 (N_4551,N_3898,N_2258);
nor U4552 (N_4552,N_4482,N_3958);
xor U4553 (N_4553,N_4329,N_4295);
and U4554 (N_4554,N_4078,N_4380);
nor U4555 (N_4555,N_4429,N_3359);
or U4556 (N_4556,N_4381,N_4412);
nor U4557 (N_4557,N_3041,N_4499);
nand U4558 (N_4558,N_4401,N_4452);
or U4559 (N_4559,N_4014,N_4384);
or U4560 (N_4560,N_3437,N_4388);
and U4561 (N_4561,N_4088,N_4000);
nor U4562 (N_4562,N_4281,N_4377);
or U4563 (N_4563,N_4479,N_3507);
or U4564 (N_4564,N_3366,N_3452);
and U4565 (N_4565,N_4290,N_2314);
nand U4566 (N_4566,N_1887,N_4469);
nand U4567 (N_4567,N_4470,N_4305);
and U4568 (N_4568,N_4258,N_4044);
nand U4569 (N_4569,N_4497,N_4268);
nand U4570 (N_4570,N_4028,N_4270);
and U4571 (N_4571,N_4433,N_1973);
and U4572 (N_4572,N_4194,N_3506);
and U4573 (N_4573,N_4311,N_4040);
xor U4574 (N_4574,N_4326,N_3691);
or U4575 (N_4575,In_2794,N_3868);
xnor U4576 (N_4576,N_4151,N_4481);
nor U4577 (N_4577,N_4367,N_4337);
nand U4578 (N_4578,N_3809,N_4246);
and U4579 (N_4579,N_4428,N_4393);
nand U4580 (N_4580,N_4414,N_4356);
xnor U4581 (N_4581,N_4241,N_2646);
nor U4582 (N_4582,N_4413,N_4343);
xnor U4583 (N_4583,N_3689,N_4346);
and U4584 (N_4584,N_4125,N_4304);
nor U4585 (N_4585,N_2771,N_4364);
and U4586 (N_4586,N_4239,N_3949);
nand U4587 (N_4587,N_4359,N_4437);
and U4588 (N_4588,N_4468,N_4154);
xnor U4589 (N_4589,N_3847,N_4330);
nor U4590 (N_4590,N_4361,N_3521);
and U4591 (N_4591,N_4288,N_4301);
and U4592 (N_4592,N_4081,N_4309);
nor U4593 (N_4593,N_4490,N_4327);
and U4594 (N_4594,N_4410,N_4251);
nor U4595 (N_4595,N_3577,N_4383);
xor U4596 (N_4596,N_4035,In_3258);
or U4597 (N_4597,N_4324,N_3938);
or U4598 (N_4598,N_3883,N_4262);
nand U4599 (N_4599,N_2484,N_4185);
nor U4600 (N_4600,N_4134,N_4474);
xor U4601 (N_4601,N_3991,N_4112);
and U4602 (N_4602,N_3226,N_3518);
nor U4603 (N_4603,N_4061,N_3776);
nor U4604 (N_4604,N_4302,N_4277);
xor U4605 (N_4605,N_2185,N_4294);
nand U4606 (N_4606,N_4095,N_4421);
and U4607 (N_4607,N_1202,In_2847);
nor U4608 (N_4608,N_3501,N_4280);
nor U4609 (N_4609,N_4208,N_2809);
nor U4610 (N_4610,N_4415,N_4358);
and U4611 (N_4611,N_3829,N_4209);
and U4612 (N_4612,N_4296,In_3413);
xor U4613 (N_4613,N_4405,N_4137);
nor U4614 (N_4614,In_3049,N_4392);
nand U4615 (N_4615,N_4041,N_4454);
xor U4616 (N_4616,N_4357,N_2639);
xor U4617 (N_4617,N_3175,N_4472);
nand U4618 (N_4618,N_4488,N_1909);
nand U4619 (N_4619,N_4106,N_4263);
nand U4620 (N_4620,N_4275,N_3986);
nor U4621 (N_4621,N_3059,N_4404);
nor U4622 (N_4622,N_4260,N_4362);
xnor U4623 (N_4623,N_4162,N_3686);
xor U4624 (N_4624,N_4314,N_4130);
and U4625 (N_4625,N_3196,N_4350);
xnor U4626 (N_4626,N_4254,N_4320);
nor U4627 (N_4627,N_793,N_4034);
nor U4628 (N_4628,N_4402,N_4485);
and U4629 (N_4629,N_4221,N_4455);
nor U4630 (N_4630,N_4480,N_3290);
and U4631 (N_4631,N_4003,N_4096);
xor U4632 (N_4632,N_4466,N_3701);
nor U4633 (N_4633,N_4494,N_3803);
nor U4634 (N_4634,N_4158,N_4312);
or U4635 (N_4635,N_4344,N_3979);
xor U4636 (N_4636,N_3643,N_4438);
or U4637 (N_4637,N_4310,N_4491);
nor U4638 (N_4638,N_3927,N_3839);
nor U4639 (N_4639,N_4459,N_4345);
xor U4640 (N_4640,N_3603,In_4239);
nor U4641 (N_4641,In_477,N_4120);
nand U4642 (N_4642,N_4338,N_3909);
nor U4643 (N_4643,N_4341,N_4257);
and U4644 (N_4644,N_4007,N_4256);
nand U4645 (N_4645,N_4308,N_2905);
and U4646 (N_4646,N_2358,N_3866);
nor U4647 (N_4647,N_4203,N_4375);
nand U4648 (N_4648,N_4395,N_4398);
xnor U4649 (N_4649,N_3176,In_955);
xnor U4650 (N_4650,N_3793,N_4259);
xnor U4651 (N_4651,N_3608,N_3081);
nand U4652 (N_4652,N_4287,N_3942);
or U4653 (N_4653,N_4486,N_4449);
nand U4654 (N_4654,N_4478,N_4394);
xnor U4655 (N_4655,In_3323,N_2332);
and U4656 (N_4656,N_4135,N_614);
nand U4657 (N_4657,N_4317,N_4144);
nand U4658 (N_4658,N_4399,N_4052);
or U4659 (N_4659,N_4306,N_4205);
or U4660 (N_4660,N_3703,N_3762);
or U4661 (N_4661,N_4417,In_2779);
or U4662 (N_4662,N_2602,N_4348);
and U4663 (N_4663,N_4029,N_4456);
and U4664 (N_4664,N_4390,N_3850);
nand U4665 (N_4665,N_4086,N_3523);
nor U4666 (N_4666,N_4036,N_401);
xor U4667 (N_4667,N_4369,N_3646);
nand U4668 (N_4668,N_4289,N_4273);
nand U4669 (N_4669,N_3486,N_509);
or U4670 (N_4670,N_4387,N_3903);
and U4671 (N_4671,N_4293,In_2735);
or U4672 (N_4672,N_3677,N_4385);
or U4673 (N_4673,N_4286,N_4386);
nand U4674 (N_4674,N_2994,N_4354);
nand U4675 (N_4675,N_4448,N_1473);
or U4676 (N_4676,N_4391,N_4420);
nor U4677 (N_4677,N_4431,N_4471);
or U4678 (N_4678,N_3318,N_2301);
nand U4679 (N_4679,N_4331,N_4368);
or U4680 (N_4680,N_4342,N_2916);
or U4681 (N_4681,N_4440,N_4416);
nand U4682 (N_4682,N_4332,N_4463);
nor U4683 (N_4683,N_4066,N_4067);
xnor U4684 (N_4684,N_3606,N_4316);
or U4685 (N_4685,N_4266,N_4155);
or U4686 (N_4686,N_3959,N_4255);
xor U4687 (N_4687,N_3404,N_2355);
nor U4688 (N_4688,N_3582,N_3477);
nand U4689 (N_4689,N_4378,N_3509);
and U4690 (N_4690,N_3914,N_3173);
xnor U4691 (N_4691,N_2336,In_269);
xor U4692 (N_4692,N_4253,N_4457);
nor U4693 (N_4693,N_4227,N_4009);
nor U4694 (N_4694,N_4353,N_3952);
nand U4695 (N_4695,N_4148,N_4444);
nand U4696 (N_4696,N_4453,N_4427);
or U4697 (N_4697,N_4119,N_4419);
xor U4698 (N_4698,N_867,N_4279);
nand U4699 (N_4699,In_769,N_3980);
nand U4700 (N_4700,N_3841,N_4238);
or U4701 (N_4701,N_4318,N_4355);
nor U4702 (N_4702,N_4458,N_2161);
or U4703 (N_4703,N_2701,N_3001);
and U4704 (N_4704,N_3252,N_4335);
nor U4705 (N_4705,N_4122,N_3915);
nor U4706 (N_4706,N_4090,N_4336);
xor U4707 (N_4707,N_4252,N_4483);
nor U4708 (N_4708,N_3789,N_4445);
nand U4709 (N_4709,N_4423,N_2362);
and U4710 (N_4710,N_4340,N_733);
nand U4711 (N_4711,N_4315,N_4464);
or U4712 (N_4712,N_4139,N_4073);
nand U4713 (N_4713,N_4396,N_2323);
and U4714 (N_4714,N_4282,N_4051);
nor U4715 (N_4715,N_2974,N_4495);
nand U4716 (N_4716,N_4303,N_4498);
nand U4717 (N_4717,N_4267,N_4283);
or U4718 (N_4718,N_4004,N_4274);
nor U4719 (N_4719,N_4461,N_4300);
nor U4720 (N_4720,N_2845,N_4418);
xnor U4721 (N_4721,N_3783,N_4379);
nand U4722 (N_4722,N_2458,N_4069);
and U4723 (N_4723,N_4422,N_2203);
xor U4724 (N_4724,N_4179,N_4496);
nand U4725 (N_4725,N_4347,N_4370);
nor U4726 (N_4726,N_4382,N_4264);
nand U4727 (N_4727,N_3966,N_4409);
or U4728 (N_4728,N_3227,N_4365);
nand U4729 (N_4729,N_4407,N_4299);
or U4730 (N_4730,N_4298,N_4265);
xor U4731 (N_4731,N_4408,N_4174);
nand U4732 (N_4732,N_4272,N_4475);
or U4733 (N_4733,N_4057,N_3843);
nand U4734 (N_4734,N_4484,N_4476);
or U4735 (N_4735,N_658,N_4374);
nor U4736 (N_4736,N_4400,N_4062);
nor U4737 (N_4737,N_1749,N_3597);
xor U4738 (N_4738,N_4171,N_2924);
xor U4739 (N_4739,In_2027,N_3777);
xor U4740 (N_4740,N_4271,N_3221);
or U4741 (N_4741,N_4025,In_3715);
nand U4742 (N_4742,N_4373,In_1932);
nor U4743 (N_4743,N_4376,N_4397);
xor U4744 (N_4744,N_4465,N_4430);
nand U4745 (N_4745,N_4319,N_4389);
or U4746 (N_4746,N_3407,N_4323);
xnor U4747 (N_4747,N_2897,N_4164);
xnor U4748 (N_4748,N_4333,N_4477);
xnor U4749 (N_4749,In_4461,N_4285);
xor U4750 (N_4750,N_4727,N_4612);
and U4751 (N_4751,N_4615,N_4636);
nand U4752 (N_4752,N_4563,N_4577);
or U4753 (N_4753,N_4582,N_4676);
xnor U4754 (N_4754,N_4541,N_4620);
or U4755 (N_4755,N_4672,N_4721);
xor U4756 (N_4756,N_4540,N_4702);
and U4757 (N_4757,N_4746,N_4630);
nor U4758 (N_4758,N_4629,N_4644);
xnor U4759 (N_4759,N_4737,N_4710);
nor U4760 (N_4760,N_4678,N_4679);
nand U4761 (N_4761,N_4673,N_4575);
nor U4762 (N_4762,N_4616,N_4628);
or U4763 (N_4763,N_4581,N_4525);
nor U4764 (N_4764,N_4553,N_4514);
nand U4765 (N_4765,N_4505,N_4684);
nor U4766 (N_4766,N_4548,N_4655);
and U4767 (N_4767,N_4669,N_4635);
and U4768 (N_4768,N_4583,N_4667);
or U4769 (N_4769,N_4743,N_4736);
xor U4770 (N_4770,N_4572,N_4698);
nor U4771 (N_4771,N_4560,N_4645);
or U4772 (N_4772,N_4703,N_4731);
and U4773 (N_4773,N_4738,N_4518);
nor U4774 (N_4774,N_4535,N_4585);
nand U4775 (N_4775,N_4653,N_4506);
nor U4776 (N_4776,N_4566,N_4602);
nor U4777 (N_4777,N_4555,N_4634);
nor U4778 (N_4778,N_4646,N_4617);
and U4779 (N_4779,N_4697,N_4732);
nand U4780 (N_4780,N_4539,N_4683);
nand U4781 (N_4781,N_4536,N_4633);
xor U4782 (N_4782,N_4614,N_4709);
nor U4783 (N_4783,N_4537,N_4598);
nand U4784 (N_4784,N_4526,N_4632);
nand U4785 (N_4785,N_4508,N_4650);
xor U4786 (N_4786,N_4661,N_4608);
nor U4787 (N_4787,N_4547,N_4619);
or U4788 (N_4788,N_4512,N_4649);
or U4789 (N_4789,N_4741,N_4519);
and U4790 (N_4790,N_4686,N_4701);
nand U4791 (N_4791,N_4704,N_4681);
xor U4792 (N_4792,N_4517,N_4692);
xnor U4793 (N_4793,N_4613,N_4603);
nand U4794 (N_4794,N_4663,N_4543);
xnor U4795 (N_4795,N_4747,N_4516);
xor U4796 (N_4796,N_4670,N_4597);
or U4797 (N_4797,N_4570,N_4587);
or U4798 (N_4798,N_4627,N_4622);
or U4799 (N_4799,N_4618,N_4579);
nand U4800 (N_4800,N_4651,N_4596);
or U4801 (N_4801,N_4641,N_4658);
and U4802 (N_4802,N_4594,N_4599);
nand U4803 (N_4803,N_4550,N_4730);
xor U4804 (N_4804,N_4677,N_4690);
nand U4805 (N_4805,N_4545,N_4657);
nor U4806 (N_4806,N_4546,N_4665);
xor U4807 (N_4807,N_4664,N_4718);
and U4808 (N_4808,N_4523,N_4584);
nor U4809 (N_4809,N_4674,N_4705);
xnor U4810 (N_4810,N_4662,N_4515);
or U4811 (N_4811,N_4590,N_4564);
xnor U4812 (N_4812,N_4671,N_4502);
xor U4813 (N_4813,N_4666,N_4643);
or U4814 (N_4814,N_4625,N_4648);
nand U4815 (N_4815,N_4503,N_4691);
nor U4816 (N_4816,N_4578,N_4529);
xor U4817 (N_4817,N_4700,N_4513);
nor U4818 (N_4818,N_4609,N_4726);
xor U4819 (N_4819,N_4593,N_4680);
nor U4820 (N_4820,N_4652,N_4600);
xor U4821 (N_4821,N_4722,N_4561);
and U4822 (N_4822,N_4574,N_4682);
nand U4823 (N_4823,N_4562,N_4527);
xor U4824 (N_4824,N_4688,N_4626);
xnor U4825 (N_4825,N_4554,N_4610);
or U4826 (N_4826,N_4604,N_4501);
nor U4827 (N_4827,N_4693,N_4511);
and U4828 (N_4828,N_4735,N_4713);
or U4829 (N_4829,N_4591,N_4638);
nand U4830 (N_4830,N_4500,N_4708);
nand U4831 (N_4831,N_4685,N_4606);
or U4832 (N_4832,N_4723,N_4605);
or U4833 (N_4833,N_4687,N_4534);
and U4834 (N_4834,N_4568,N_4571);
nand U4835 (N_4835,N_4725,N_4601);
and U4836 (N_4836,N_4711,N_4734);
or U4837 (N_4837,N_4538,N_4706);
nand U4838 (N_4838,N_4558,N_4694);
and U4839 (N_4839,N_4668,N_4717);
xor U4840 (N_4840,N_4699,N_4637);
nand U4841 (N_4841,N_4507,N_4559);
or U4842 (N_4842,N_4524,N_4544);
xor U4843 (N_4843,N_4696,N_4504);
nor U4844 (N_4844,N_4576,N_4552);
nor U4845 (N_4845,N_4531,N_4689);
nor U4846 (N_4846,N_4586,N_4509);
nand U4847 (N_4847,N_4528,N_4660);
nand U4848 (N_4848,N_4647,N_4588);
xnor U4849 (N_4849,N_4530,N_4532);
nor U4850 (N_4850,N_4733,N_4556);
and U4851 (N_4851,N_4569,N_4719);
xnor U4852 (N_4852,N_4712,N_4520);
or U4853 (N_4853,N_4551,N_4549);
nor U4854 (N_4854,N_4567,N_4695);
nor U4855 (N_4855,N_4522,N_4714);
or U4856 (N_4856,N_4749,N_4744);
nand U4857 (N_4857,N_4621,N_4707);
and U4858 (N_4858,N_4624,N_4595);
xor U4859 (N_4859,N_4589,N_4748);
and U4860 (N_4860,N_4724,N_4716);
xnor U4861 (N_4861,N_4729,N_4623);
and U4862 (N_4862,N_4510,N_4742);
nand U4863 (N_4863,N_4521,N_4745);
nor U4864 (N_4864,N_4533,N_4580);
and U4865 (N_4865,N_4715,N_4740);
or U4866 (N_4866,N_4542,N_4739);
or U4867 (N_4867,N_4639,N_4607);
nor U4868 (N_4868,N_4565,N_4631);
or U4869 (N_4869,N_4720,N_4728);
and U4870 (N_4870,N_4656,N_4642);
nand U4871 (N_4871,N_4654,N_4675);
and U4872 (N_4872,N_4592,N_4573);
and U4873 (N_4873,N_4659,N_4611);
xnor U4874 (N_4874,N_4640,N_4557);
nor U4875 (N_4875,N_4603,N_4676);
and U4876 (N_4876,N_4621,N_4598);
and U4877 (N_4877,N_4558,N_4567);
and U4878 (N_4878,N_4585,N_4717);
nand U4879 (N_4879,N_4502,N_4596);
xnor U4880 (N_4880,N_4560,N_4598);
nand U4881 (N_4881,N_4722,N_4721);
or U4882 (N_4882,N_4613,N_4506);
xnor U4883 (N_4883,N_4711,N_4739);
or U4884 (N_4884,N_4670,N_4745);
or U4885 (N_4885,N_4550,N_4578);
nor U4886 (N_4886,N_4544,N_4703);
and U4887 (N_4887,N_4606,N_4687);
nand U4888 (N_4888,N_4702,N_4734);
and U4889 (N_4889,N_4705,N_4733);
or U4890 (N_4890,N_4701,N_4544);
xnor U4891 (N_4891,N_4622,N_4656);
nor U4892 (N_4892,N_4523,N_4625);
or U4893 (N_4893,N_4685,N_4628);
xor U4894 (N_4894,N_4639,N_4556);
nor U4895 (N_4895,N_4679,N_4552);
nand U4896 (N_4896,N_4693,N_4590);
xor U4897 (N_4897,N_4648,N_4549);
or U4898 (N_4898,N_4588,N_4714);
and U4899 (N_4899,N_4630,N_4678);
xor U4900 (N_4900,N_4534,N_4667);
nand U4901 (N_4901,N_4518,N_4618);
nand U4902 (N_4902,N_4657,N_4600);
xnor U4903 (N_4903,N_4507,N_4629);
and U4904 (N_4904,N_4581,N_4542);
nand U4905 (N_4905,N_4634,N_4608);
or U4906 (N_4906,N_4643,N_4727);
and U4907 (N_4907,N_4738,N_4571);
xor U4908 (N_4908,N_4683,N_4630);
xnor U4909 (N_4909,N_4604,N_4578);
nor U4910 (N_4910,N_4633,N_4671);
nand U4911 (N_4911,N_4683,N_4720);
nand U4912 (N_4912,N_4661,N_4606);
nor U4913 (N_4913,N_4597,N_4687);
or U4914 (N_4914,N_4501,N_4598);
nand U4915 (N_4915,N_4672,N_4604);
or U4916 (N_4916,N_4673,N_4657);
xor U4917 (N_4917,N_4567,N_4688);
nand U4918 (N_4918,N_4689,N_4702);
nor U4919 (N_4919,N_4575,N_4594);
or U4920 (N_4920,N_4605,N_4628);
xnor U4921 (N_4921,N_4676,N_4664);
nor U4922 (N_4922,N_4559,N_4605);
or U4923 (N_4923,N_4571,N_4642);
or U4924 (N_4924,N_4598,N_4684);
and U4925 (N_4925,N_4741,N_4706);
nand U4926 (N_4926,N_4523,N_4599);
nand U4927 (N_4927,N_4564,N_4603);
nand U4928 (N_4928,N_4666,N_4614);
nand U4929 (N_4929,N_4544,N_4649);
nor U4930 (N_4930,N_4690,N_4673);
or U4931 (N_4931,N_4642,N_4507);
or U4932 (N_4932,N_4543,N_4573);
xnor U4933 (N_4933,N_4658,N_4594);
or U4934 (N_4934,N_4720,N_4542);
nor U4935 (N_4935,N_4691,N_4523);
and U4936 (N_4936,N_4674,N_4524);
or U4937 (N_4937,N_4567,N_4575);
nand U4938 (N_4938,N_4717,N_4563);
and U4939 (N_4939,N_4629,N_4721);
and U4940 (N_4940,N_4707,N_4516);
and U4941 (N_4941,N_4583,N_4727);
and U4942 (N_4942,N_4692,N_4715);
nand U4943 (N_4943,N_4594,N_4651);
and U4944 (N_4944,N_4698,N_4716);
xnor U4945 (N_4945,N_4720,N_4686);
nor U4946 (N_4946,N_4637,N_4672);
nand U4947 (N_4947,N_4585,N_4681);
xor U4948 (N_4948,N_4746,N_4514);
nor U4949 (N_4949,N_4663,N_4719);
nor U4950 (N_4950,N_4550,N_4649);
and U4951 (N_4951,N_4741,N_4717);
nor U4952 (N_4952,N_4651,N_4562);
xnor U4953 (N_4953,N_4500,N_4609);
and U4954 (N_4954,N_4658,N_4710);
xnor U4955 (N_4955,N_4540,N_4512);
xnor U4956 (N_4956,N_4659,N_4594);
xnor U4957 (N_4957,N_4736,N_4516);
nor U4958 (N_4958,N_4700,N_4736);
or U4959 (N_4959,N_4733,N_4708);
and U4960 (N_4960,N_4666,N_4746);
and U4961 (N_4961,N_4675,N_4749);
nor U4962 (N_4962,N_4535,N_4575);
or U4963 (N_4963,N_4699,N_4745);
and U4964 (N_4964,N_4653,N_4513);
nand U4965 (N_4965,N_4596,N_4511);
xnor U4966 (N_4966,N_4639,N_4550);
nor U4967 (N_4967,N_4593,N_4702);
or U4968 (N_4968,N_4504,N_4589);
xor U4969 (N_4969,N_4700,N_4699);
xnor U4970 (N_4970,N_4566,N_4505);
xnor U4971 (N_4971,N_4706,N_4675);
xnor U4972 (N_4972,N_4564,N_4589);
nor U4973 (N_4973,N_4534,N_4539);
nor U4974 (N_4974,N_4500,N_4734);
and U4975 (N_4975,N_4609,N_4664);
nand U4976 (N_4976,N_4542,N_4749);
nand U4977 (N_4977,N_4558,N_4555);
nor U4978 (N_4978,N_4635,N_4506);
nor U4979 (N_4979,N_4653,N_4744);
or U4980 (N_4980,N_4641,N_4726);
nor U4981 (N_4981,N_4610,N_4502);
nor U4982 (N_4982,N_4744,N_4630);
or U4983 (N_4983,N_4511,N_4502);
xor U4984 (N_4984,N_4675,N_4717);
xnor U4985 (N_4985,N_4609,N_4622);
or U4986 (N_4986,N_4518,N_4516);
xnor U4987 (N_4987,N_4681,N_4684);
and U4988 (N_4988,N_4639,N_4516);
nand U4989 (N_4989,N_4614,N_4668);
nor U4990 (N_4990,N_4644,N_4717);
or U4991 (N_4991,N_4660,N_4521);
or U4992 (N_4992,N_4730,N_4633);
and U4993 (N_4993,N_4599,N_4537);
xnor U4994 (N_4994,N_4563,N_4705);
xnor U4995 (N_4995,N_4637,N_4629);
and U4996 (N_4996,N_4705,N_4515);
and U4997 (N_4997,N_4598,N_4719);
nor U4998 (N_4998,N_4524,N_4505);
nand U4999 (N_4999,N_4540,N_4560);
or U5000 (N_5000,N_4884,N_4874);
and U5001 (N_5001,N_4825,N_4821);
nor U5002 (N_5002,N_4794,N_4954);
xor U5003 (N_5003,N_4799,N_4784);
xor U5004 (N_5004,N_4993,N_4869);
or U5005 (N_5005,N_4816,N_4945);
and U5006 (N_5006,N_4877,N_4774);
and U5007 (N_5007,N_4786,N_4820);
nor U5008 (N_5008,N_4873,N_4887);
and U5009 (N_5009,N_4757,N_4853);
and U5010 (N_5010,N_4771,N_4787);
or U5011 (N_5011,N_4909,N_4833);
or U5012 (N_5012,N_4751,N_4768);
and U5013 (N_5013,N_4906,N_4889);
nor U5014 (N_5014,N_4900,N_4929);
nor U5015 (N_5015,N_4978,N_4922);
nand U5016 (N_5016,N_4994,N_4948);
nor U5017 (N_5017,N_4933,N_4987);
and U5018 (N_5018,N_4932,N_4903);
nand U5019 (N_5019,N_4805,N_4928);
and U5020 (N_5020,N_4923,N_4913);
xnor U5021 (N_5021,N_4898,N_4844);
nand U5022 (N_5022,N_4990,N_4983);
or U5023 (N_5023,N_4755,N_4885);
xnor U5024 (N_5024,N_4819,N_4812);
and U5025 (N_5025,N_4785,N_4826);
xor U5026 (N_5026,N_4813,N_4952);
nor U5027 (N_5027,N_4750,N_4902);
xnor U5028 (N_5028,N_4829,N_4959);
nor U5029 (N_5029,N_4895,N_4924);
xor U5030 (N_5030,N_4807,N_4958);
xnor U5031 (N_5031,N_4834,N_4839);
nand U5032 (N_5032,N_4998,N_4846);
xnor U5033 (N_5033,N_4946,N_4880);
or U5034 (N_5034,N_4966,N_4775);
nor U5035 (N_5035,N_4767,N_4836);
and U5036 (N_5036,N_4843,N_4861);
nand U5037 (N_5037,N_4942,N_4917);
or U5038 (N_5038,N_4970,N_4875);
nand U5039 (N_5039,N_4842,N_4972);
or U5040 (N_5040,N_4817,N_4968);
and U5041 (N_5041,N_4862,N_4940);
nor U5042 (N_5042,N_4852,N_4883);
and U5043 (N_5043,N_4871,N_4851);
and U5044 (N_5044,N_4879,N_4863);
or U5045 (N_5045,N_4988,N_4753);
nand U5046 (N_5046,N_4802,N_4960);
nor U5047 (N_5047,N_4865,N_4927);
nand U5048 (N_5048,N_4882,N_4769);
xor U5049 (N_5049,N_4788,N_4758);
nand U5050 (N_5050,N_4752,N_4763);
or U5051 (N_5051,N_4806,N_4838);
nor U5052 (N_5052,N_4860,N_4891);
nand U5053 (N_5053,N_4830,N_4803);
xnor U5054 (N_5054,N_4809,N_4951);
or U5055 (N_5055,N_4992,N_4956);
and U5056 (N_5056,N_4849,N_4930);
nor U5057 (N_5057,N_4881,N_4893);
nand U5058 (N_5058,N_4811,N_4872);
nor U5059 (N_5059,N_4938,N_4984);
and U5060 (N_5060,N_4770,N_4981);
or U5061 (N_5061,N_4965,N_4814);
xnor U5062 (N_5062,N_4778,N_4798);
or U5063 (N_5063,N_4975,N_4756);
or U5064 (N_5064,N_4762,N_4989);
nor U5065 (N_5065,N_4991,N_4907);
or U5066 (N_5066,N_4947,N_4766);
nor U5067 (N_5067,N_4870,N_4760);
nor U5068 (N_5068,N_4916,N_4973);
and U5069 (N_5069,N_4776,N_4901);
and U5070 (N_5070,N_4919,N_4997);
and U5071 (N_5071,N_4828,N_4854);
and U5072 (N_5072,N_4921,N_4824);
or U5073 (N_5073,N_4912,N_4772);
nand U5074 (N_5074,N_4980,N_4969);
xnor U5075 (N_5075,N_4831,N_4858);
xor U5076 (N_5076,N_4804,N_4962);
xor U5077 (N_5077,N_4995,N_4855);
xnor U5078 (N_5078,N_4935,N_4761);
nor U5079 (N_5079,N_4795,N_4979);
or U5080 (N_5080,N_4827,N_4890);
or U5081 (N_5081,N_4796,N_4868);
and U5082 (N_5082,N_4944,N_4949);
xnor U5083 (N_5083,N_4850,N_4777);
nand U5084 (N_5084,N_4985,N_4801);
or U5085 (N_5085,N_4996,N_4918);
nand U5086 (N_5086,N_4892,N_4925);
xnor U5087 (N_5087,N_4792,N_4876);
xor U5088 (N_5088,N_4967,N_4971);
nor U5089 (N_5089,N_4931,N_4832);
xor U5090 (N_5090,N_4790,N_4976);
nand U5091 (N_5091,N_4964,N_4905);
xnor U5092 (N_5092,N_4797,N_4859);
nand U5093 (N_5093,N_4754,N_4939);
nand U5094 (N_5094,N_4974,N_4982);
and U5095 (N_5095,N_4793,N_4963);
nor U5096 (N_5096,N_4941,N_4800);
and U5097 (N_5097,N_4822,N_4910);
or U5098 (N_5098,N_4781,N_4866);
or U5099 (N_5099,N_4765,N_4955);
xor U5100 (N_5100,N_4837,N_4911);
xnor U5101 (N_5101,N_4789,N_4920);
nand U5102 (N_5102,N_4914,N_4897);
or U5103 (N_5103,N_4864,N_4791);
and U5104 (N_5104,N_4953,N_4904);
xnor U5105 (N_5105,N_4810,N_4857);
xor U5106 (N_5106,N_4950,N_4961);
or U5107 (N_5107,N_4908,N_4759);
or U5108 (N_5108,N_4818,N_4823);
or U5109 (N_5109,N_4856,N_4808);
xor U5110 (N_5110,N_4845,N_4888);
and U5111 (N_5111,N_4934,N_4783);
nand U5112 (N_5112,N_4899,N_4894);
and U5113 (N_5113,N_4841,N_4848);
nand U5114 (N_5114,N_4936,N_4926);
or U5115 (N_5115,N_4878,N_4773);
nor U5116 (N_5116,N_4779,N_4867);
or U5117 (N_5117,N_4896,N_4957);
or U5118 (N_5118,N_4915,N_4782);
and U5119 (N_5119,N_4999,N_4986);
and U5120 (N_5120,N_4886,N_4937);
or U5121 (N_5121,N_4815,N_4847);
xnor U5122 (N_5122,N_4943,N_4977);
xor U5123 (N_5123,N_4764,N_4835);
xnor U5124 (N_5124,N_4780,N_4840);
or U5125 (N_5125,N_4937,N_4905);
nand U5126 (N_5126,N_4936,N_4801);
xnor U5127 (N_5127,N_4827,N_4809);
or U5128 (N_5128,N_4989,N_4953);
nand U5129 (N_5129,N_4788,N_4967);
or U5130 (N_5130,N_4844,N_4908);
and U5131 (N_5131,N_4755,N_4883);
nor U5132 (N_5132,N_4900,N_4918);
nand U5133 (N_5133,N_4852,N_4857);
nor U5134 (N_5134,N_4755,N_4794);
nand U5135 (N_5135,N_4880,N_4902);
or U5136 (N_5136,N_4956,N_4929);
and U5137 (N_5137,N_4847,N_4785);
nand U5138 (N_5138,N_4783,N_4810);
xor U5139 (N_5139,N_4928,N_4964);
nor U5140 (N_5140,N_4954,N_4802);
nand U5141 (N_5141,N_4792,N_4977);
xor U5142 (N_5142,N_4926,N_4805);
nand U5143 (N_5143,N_4985,N_4999);
xnor U5144 (N_5144,N_4989,N_4969);
nor U5145 (N_5145,N_4883,N_4906);
nor U5146 (N_5146,N_4884,N_4795);
or U5147 (N_5147,N_4951,N_4841);
xor U5148 (N_5148,N_4793,N_4751);
nor U5149 (N_5149,N_4943,N_4964);
and U5150 (N_5150,N_4860,N_4798);
xnor U5151 (N_5151,N_4945,N_4993);
nor U5152 (N_5152,N_4866,N_4821);
nor U5153 (N_5153,N_4788,N_4970);
nor U5154 (N_5154,N_4992,N_4833);
nor U5155 (N_5155,N_4999,N_4779);
and U5156 (N_5156,N_4857,N_4926);
or U5157 (N_5157,N_4984,N_4763);
nand U5158 (N_5158,N_4960,N_4984);
or U5159 (N_5159,N_4953,N_4790);
xor U5160 (N_5160,N_4822,N_4924);
nor U5161 (N_5161,N_4969,N_4929);
and U5162 (N_5162,N_4896,N_4816);
and U5163 (N_5163,N_4789,N_4770);
nand U5164 (N_5164,N_4858,N_4967);
xor U5165 (N_5165,N_4869,N_4945);
xor U5166 (N_5166,N_4849,N_4931);
xnor U5167 (N_5167,N_4812,N_4850);
nand U5168 (N_5168,N_4938,N_4751);
and U5169 (N_5169,N_4837,N_4792);
or U5170 (N_5170,N_4886,N_4905);
xor U5171 (N_5171,N_4825,N_4971);
or U5172 (N_5172,N_4805,N_4980);
nand U5173 (N_5173,N_4992,N_4834);
xor U5174 (N_5174,N_4867,N_4798);
nand U5175 (N_5175,N_4754,N_4869);
or U5176 (N_5176,N_4782,N_4887);
or U5177 (N_5177,N_4986,N_4870);
nand U5178 (N_5178,N_4888,N_4943);
nand U5179 (N_5179,N_4817,N_4871);
and U5180 (N_5180,N_4932,N_4818);
nor U5181 (N_5181,N_4861,N_4784);
nor U5182 (N_5182,N_4835,N_4932);
or U5183 (N_5183,N_4977,N_4772);
or U5184 (N_5184,N_4870,N_4901);
xnor U5185 (N_5185,N_4884,N_4767);
and U5186 (N_5186,N_4782,N_4898);
and U5187 (N_5187,N_4979,N_4897);
nand U5188 (N_5188,N_4999,N_4947);
nand U5189 (N_5189,N_4964,N_4779);
xnor U5190 (N_5190,N_4970,N_4989);
and U5191 (N_5191,N_4884,N_4938);
xnor U5192 (N_5192,N_4750,N_4899);
nor U5193 (N_5193,N_4881,N_4795);
or U5194 (N_5194,N_4848,N_4859);
nor U5195 (N_5195,N_4823,N_4925);
or U5196 (N_5196,N_4803,N_4974);
nand U5197 (N_5197,N_4856,N_4939);
or U5198 (N_5198,N_4774,N_4860);
and U5199 (N_5199,N_4882,N_4764);
nand U5200 (N_5200,N_4805,N_4825);
nand U5201 (N_5201,N_4779,N_4983);
and U5202 (N_5202,N_4855,N_4988);
xor U5203 (N_5203,N_4838,N_4792);
or U5204 (N_5204,N_4914,N_4942);
nor U5205 (N_5205,N_4919,N_4937);
xnor U5206 (N_5206,N_4839,N_4779);
or U5207 (N_5207,N_4754,N_4877);
xor U5208 (N_5208,N_4892,N_4941);
and U5209 (N_5209,N_4909,N_4988);
nand U5210 (N_5210,N_4929,N_4954);
nor U5211 (N_5211,N_4796,N_4849);
or U5212 (N_5212,N_4956,N_4918);
xor U5213 (N_5213,N_4756,N_4906);
nor U5214 (N_5214,N_4931,N_4755);
xor U5215 (N_5215,N_4932,N_4881);
or U5216 (N_5216,N_4840,N_4978);
or U5217 (N_5217,N_4830,N_4860);
or U5218 (N_5218,N_4959,N_4926);
nor U5219 (N_5219,N_4936,N_4827);
nor U5220 (N_5220,N_4984,N_4858);
and U5221 (N_5221,N_4873,N_4985);
and U5222 (N_5222,N_4800,N_4829);
and U5223 (N_5223,N_4993,N_4874);
nor U5224 (N_5224,N_4846,N_4915);
nor U5225 (N_5225,N_4816,N_4828);
or U5226 (N_5226,N_4796,N_4882);
xor U5227 (N_5227,N_4872,N_4914);
nor U5228 (N_5228,N_4806,N_4797);
nand U5229 (N_5229,N_4774,N_4834);
and U5230 (N_5230,N_4754,N_4862);
nor U5231 (N_5231,N_4831,N_4990);
xnor U5232 (N_5232,N_4916,N_4807);
nor U5233 (N_5233,N_4901,N_4859);
and U5234 (N_5234,N_4936,N_4811);
nor U5235 (N_5235,N_4855,N_4876);
nand U5236 (N_5236,N_4885,N_4785);
or U5237 (N_5237,N_4918,N_4968);
xor U5238 (N_5238,N_4797,N_4794);
nor U5239 (N_5239,N_4862,N_4792);
nor U5240 (N_5240,N_4933,N_4830);
or U5241 (N_5241,N_4915,N_4767);
or U5242 (N_5242,N_4937,N_4847);
and U5243 (N_5243,N_4881,N_4885);
nor U5244 (N_5244,N_4869,N_4757);
nand U5245 (N_5245,N_4896,N_4925);
or U5246 (N_5246,N_4924,N_4870);
and U5247 (N_5247,N_4974,N_4781);
or U5248 (N_5248,N_4935,N_4973);
xor U5249 (N_5249,N_4890,N_4776);
nand U5250 (N_5250,N_5031,N_5144);
nand U5251 (N_5251,N_5126,N_5046);
or U5252 (N_5252,N_5245,N_5184);
nand U5253 (N_5253,N_5098,N_5217);
nor U5254 (N_5254,N_5199,N_5226);
and U5255 (N_5255,N_5118,N_5124);
and U5256 (N_5256,N_5102,N_5053);
xnor U5257 (N_5257,N_5151,N_5248);
or U5258 (N_5258,N_5106,N_5224);
and U5259 (N_5259,N_5092,N_5074);
nor U5260 (N_5260,N_5197,N_5081);
or U5261 (N_5261,N_5166,N_5119);
and U5262 (N_5262,N_5146,N_5041);
nand U5263 (N_5263,N_5194,N_5061);
or U5264 (N_5264,N_5138,N_5085);
nor U5265 (N_5265,N_5228,N_5071);
nor U5266 (N_5266,N_5082,N_5060);
nor U5267 (N_5267,N_5019,N_5153);
nor U5268 (N_5268,N_5243,N_5103);
and U5269 (N_5269,N_5037,N_5149);
nand U5270 (N_5270,N_5120,N_5008);
nor U5271 (N_5271,N_5180,N_5208);
xor U5272 (N_5272,N_5001,N_5070);
and U5273 (N_5273,N_5003,N_5158);
or U5274 (N_5274,N_5054,N_5203);
and U5275 (N_5275,N_5067,N_5006);
or U5276 (N_5276,N_5056,N_5175);
and U5277 (N_5277,N_5177,N_5160);
nand U5278 (N_5278,N_5219,N_5017);
and U5279 (N_5279,N_5117,N_5131);
nand U5280 (N_5280,N_5134,N_5209);
nand U5281 (N_5281,N_5018,N_5049);
xnor U5282 (N_5282,N_5140,N_5167);
and U5283 (N_5283,N_5002,N_5097);
and U5284 (N_5284,N_5240,N_5246);
nand U5285 (N_5285,N_5173,N_5005);
nor U5286 (N_5286,N_5236,N_5139);
nand U5287 (N_5287,N_5135,N_5183);
and U5288 (N_5288,N_5030,N_5028);
nand U5289 (N_5289,N_5057,N_5155);
nor U5290 (N_5290,N_5221,N_5068);
and U5291 (N_5291,N_5244,N_5233);
nor U5292 (N_5292,N_5052,N_5156);
nor U5293 (N_5293,N_5210,N_5215);
or U5294 (N_5294,N_5076,N_5211);
nor U5295 (N_5295,N_5036,N_5190);
nor U5296 (N_5296,N_5200,N_5004);
nor U5297 (N_5297,N_5172,N_5242);
nand U5298 (N_5298,N_5050,N_5170);
nor U5299 (N_5299,N_5114,N_5062);
and U5300 (N_5300,N_5168,N_5162);
nor U5301 (N_5301,N_5132,N_5058);
or U5302 (N_5302,N_5064,N_5129);
xor U5303 (N_5303,N_5145,N_5109);
nand U5304 (N_5304,N_5013,N_5047);
nand U5305 (N_5305,N_5027,N_5011);
or U5306 (N_5306,N_5086,N_5009);
or U5307 (N_5307,N_5234,N_5029);
or U5308 (N_5308,N_5195,N_5218);
nor U5309 (N_5309,N_5178,N_5164);
nand U5310 (N_5310,N_5213,N_5142);
nand U5311 (N_5311,N_5077,N_5084);
nand U5312 (N_5312,N_5137,N_5038);
nand U5313 (N_5313,N_5043,N_5113);
nand U5314 (N_5314,N_5127,N_5187);
nand U5315 (N_5315,N_5022,N_5089);
xor U5316 (N_5316,N_5032,N_5035);
nor U5317 (N_5317,N_5222,N_5059);
nand U5318 (N_5318,N_5096,N_5010);
xor U5319 (N_5319,N_5093,N_5107);
nor U5320 (N_5320,N_5148,N_5110);
nor U5321 (N_5321,N_5101,N_5034);
and U5322 (N_5322,N_5090,N_5189);
or U5323 (N_5323,N_5133,N_5123);
or U5324 (N_5324,N_5014,N_5238);
nand U5325 (N_5325,N_5078,N_5185);
or U5326 (N_5326,N_5202,N_5136);
nor U5327 (N_5327,N_5212,N_5021);
and U5328 (N_5328,N_5020,N_5108);
or U5329 (N_5329,N_5044,N_5048);
and U5330 (N_5330,N_5186,N_5191);
and U5331 (N_5331,N_5176,N_5141);
nor U5332 (N_5332,N_5179,N_5051);
xnor U5333 (N_5333,N_5111,N_5235);
and U5334 (N_5334,N_5066,N_5165);
or U5335 (N_5335,N_5122,N_5152);
nand U5336 (N_5336,N_5237,N_5104);
and U5337 (N_5337,N_5055,N_5094);
xnor U5338 (N_5338,N_5116,N_5042);
xor U5339 (N_5339,N_5040,N_5024);
xnor U5340 (N_5340,N_5161,N_5225);
or U5341 (N_5341,N_5112,N_5174);
nand U5342 (N_5342,N_5039,N_5000);
and U5343 (N_5343,N_5227,N_5025);
or U5344 (N_5344,N_5007,N_5087);
or U5345 (N_5345,N_5157,N_5171);
nand U5346 (N_5346,N_5181,N_5150);
xnor U5347 (N_5347,N_5163,N_5045);
xnor U5348 (N_5348,N_5100,N_5154);
nor U5349 (N_5349,N_5080,N_5249);
nor U5350 (N_5350,N_5205,N_5201);
or U5351 (N_5351,N_5083,N_5230);
nor U5352 (N_5352,N_5220,N_5073);
nand U5353 (N_5353,N_5015,N_5072);
or U5354 (N_5354,N_5069,N_5128);
or U5355 (N_5355,N_5247,N_5099);
or U5356 (N_5356,N_5206,N_5091);
or U5357 (N_5357,N_5204,N_5130);
nand U5358 (N_5358,N_5214,N_5033);
or U5359 (N_5359,N_5147,N_5231);
or U5360 (N_5360,N_5159,N_5182);
xnor U5361 (N_5361,N_5216,N_5088);
nor U5362 (N_5362,N_5198,N_5115);
nor U5363 (N_5363,N_5193,N_5012);
and U5364 (N_5364,N_5105,N_5143);
xor U5365 (N_5365,N_5079,N_5192);
nor U5366 (N_5366,N_5065,N_5095);
nand U5367 (N_5367,N_5196,N_5232);
nor U5368 (N_5368,N_5063,N_5169);
and U5369 (N_5369,N_5121,N_5241);
or U5370 (N_5370,N_5016,N_5023);
nand U5371 (N_5371,N_5229,N_5125);
nand U5372 (N_5372,N_5188,N_5223);
nand U5373 (N_5373,N_5239,N_5075);
and U5374 (N_5374,N_5207,N_5026);
nor U5375 (N_5375,N_5055,N_5211);
xnor U5376 (N_5376,N_5135,N_5186);
or U5377 (N_5377,N_5057,N_5196);
or U5378 (N_5378,N_5165,N_5079);
and U5379 (N_5379,N_5032,N_5241);
or U5380 (N_5380,N_5177,N_5080);
xor U5381 (N_5381,N_5014,N_5108);
and U5382 (N_5382,N_5240,N_5247);
nor U5383 (N_5383,N_5211,N_5092);
and U5384 (N_5384,N_5104,N_5059);
nor U5385 (N_5385,N_5195,N_5041);
and U5386 (N_5386,N_5173,N_5047);
nand U5387 (N_5387,N_5209,N_5175);
nand U5388 (N_5388,N_5075,N_5036);
and U5389 (N_5389,N_5177,N_5207);
and U5390 (N_5390,N_5129,N_5232);
nand U5391 (N_5391,N_5114,N_5028);
nand U5392 (N_5392,N_5168,N_5236);
xnor U5393 (N_5393,N_5231,N_5238);
nand U5394 (N_5394,N_5112,N_5003);
nand U5395 (N_5395,N_5232,N_5109);
nor U5396 (N_5396,N_5146,N_5153);
and U5397 (N_5397,N_5199,N_5229);
and U5398 (N_5398,N_5128,N_5105);
nand U5399 (N_5399,N_5225,N_5070);
nor U5400 (N_5400,N_5076,N_5056);
or U5401 (N_5401,N_5099,N_5052);
and U5402 (N_5402,N_5108,N_5242);
nor U5403 (N_5403,N_5026,N_5149);
or U5404 (N_5404,N_5165,N_5222);
xor U5405 (N_5405,N_5057,N_5246);
xor U5406 (N_5406,N_5126,N_5201);
xnor U5407 (N_5407,N_5056,N_5155);
or U5408 (N_5408,N_5177,N_5014);
nand U5409 (N_5409,N_5226,N_5175);
nor U5410 (N_5410,N_5088,N_5013);
nand U5411 (N_5411,N_5229,N_5001);
and U5412 (N_5412,N_5119,N_5201);
nor U5413 (N_5413,N_5040,N_5041);
and U5414 (N_5414,N_5065,N_5003);
and U5415 (N_5415,N_5040,N_5208);
xnor U5416 (N_5416,N_5135,N_5188);
nor U5417 (N_5417,N_5129,N_5013);
xor U5418 (N_5418,N_5006,N_5175);
or U5419 (N_5419,N_5012,N_5197);
nor U5420 (N_5420,N_5213,N_5170);
nand U5421 (N_5421,N_5232,N_5244);
nand U5422 (N_5422,N_5054,N_5002);
nor U5423 (N_5423,N_5054,N_5223);
xnor U5424 (N_5424,N_5022,N_5076);
and U5425 (N_5425,N_5241,N_5073);
xnor U5426 (N_5426,N_5215,N_5140);
or U5427 (N_5427,N_5044,N_5154);
xor U5428 (N_5428,N_5215,N_5051);
xor U5429 (N_5429,N_5138,N_5162);
nand U5430 (N_5430,N_5046,N_5012);
nand U5431 (N_5431,N_5029,N_5149);
nor U5432 (N_5432,N_5109,N_5000);
or U5433 (N_5433,N_5009,N_5214);
xor U5434 (N_5434,N_5078,N_5065);
and U5435 (N_5435,N_5230,N_5001);
or U5436 (N_5436,N_5075,N_5234);
and U5437 (N_5437,N_5117,N_5160);
or U5438 (N_5438,N_5041,N_5239);
nor U5439 (N_5439,N_5044,N_5194);
nand U5440 (N_5440,N_5035,N_5127);
nand U5441 (N_5441,N_5133,N_5075);
or U5442 (N_5442,N_5014,N_5208);
and U5443 (N_5443,N_5038,N_5141);
nand U5444 (N_5444,N_5146,N_5142);
nand U5445 (N_5445,N_5027,N_5016);
xor U5446 (N_5446,N_5188,N_5125);
nor U5447 (N_5447,N_5226,N_5239);
xnor U5448 (N_5448,N_5072,N_5018);
nor U5449 (N_5449,N_5067,N_5002);
nor U5450 (N_5450,N_5064,N_5011);
nor U5451 (N_5451,N_5109,N_5014);
nand U5452 (N_5452,N_5080,N_5105);
xor U5453 (N_5453,N_5120,N_5172);
xor U5454 (N_5454,N_5033,N_5043);
or U5455 (N_5455,N_5239,N_5163);
nor U5456 (N_5456,N_5219,N_5190);
xor U5457 (N_5457,N_5041,N_5100);
nand U5458 (N_5458,N_5094,N_5173);
and U5459 (N_5459,N_5003,N_5101);
or U5460 (N_5460,N_5101,N_5082);
nand U5461 (N_5461,N_5241,N_5172);
nor U5462 (N_5462,N_5038,N_5013);
and U5463 (N_5463,N_5205,N_5109);
xor U5464 (N_5464,N_5161,N_5239);
nor U5465 (N_5465,N_5053,N_5164);
nand U5466 (N_5466,N_5116,N_5107);
or U5467 (N_5467,N_5181,N_5160);
and U5468 (N_5468,N_5178,N_5148);
xnor U5469 (N_5469,N_5033,N_5186);
and U5470 (N_5470,N_5151,N_5014);
nor U5471 (N_5471,N_5176,N_5206);
and U5472 (N_5472,N_5200,N_5117);
xnor U5473 (N_5473,N_5181,N_5231);
and U5474 (N_5474,N_5098,N_5029);
nor U5475 (N_5475,N_5022,N_5101);
and U5476 (N_5476,N_5032,N_5188);
nor U5477 (N_5477,N_5044,N_5024);
nand U5478 (N_5478,N_5046,N_5063);
xor U5479 (N_5479,N_5085,N_5239);
nor U5480 (N_5480,N_5091,N_5234);
xnor U5481 (N_5481,N_5182,N_5215);
and U5482 (N_5482,N_5218,N_5157);
or U5483 (N_5483,N_5226,N_5014);
xor U5484 (N_5484,N_5111,N_5230);
and U5485 (N_5485,N_5110,N_5182);
or U5486 (N_5486,N_5238,N_5026);
and U5487 (N_5487,N_5117,N_5158);
xnor U5488 (N_5488,N_5060,N_5026);
nand U5489 (N_5489,N_5097,N_5088);
xnor U5490 (N_5490,N_5094,N_5157);
xnor U5491 (N_5491,N_5000,N_5185);
nor U5492 (N_5492,N_5015,N_5154);
nor U5493 (N_5493,N_5117,N_5017);
nor U5494 (N_5494,N_5082,N_5085);
or U5495 (N_5495,N_5209,N_5130);
or U5496 (N_5496,N_5049,N_5143);
and U5497 (N_5497,N_5188,N_5119);
nor U5498 (N_5498,N_5242,N_5110);
xor U5499 (N_5499,N_5064,N_5244);
xnor U5500 (N_5500,N_5490,N_5372);
xor U5501 (N_5501,N_5459,N_5401);
nor U5502 (N_5502,N_5368,N_5434);
xor U5503 (N_5503,N_5413,N_5478);
or U5504 (N_5504,N_5393,N_5255);
or U5505 (N_5505,N_5306,N_5251);
nor U5506 (N_5506,N_5287,N_5286);
or U5507 (N_5507,N_5273,N_5353);
nor U5508 (N_5508,N_5440,N_5317);
nor U5509 (N_5509,N_5430,N_5428);
nand U5510 (N_5510,N_5263,N_5330);
xor U5511 (N_5511,N_5480,N_5270);
or U5512 (N_5512,N_5378,N_5408);
xnor U5513 (N_5513,N_5448,N_5371);
and U5514 (N_5514,N_5276,N_5265);
xor U5515 (N_5515,N_5380,N_5322);
nand U5516 (N_5516,N_5320,N_5376);
nor U5517 (N_5517,N_5453,N_5477);
or U5518 (N_5518,N_5429,N_5405);
or U5519 (N_5519,N_5302,N_5410);
and U5520 (N_5520,N_5421,N_5484);
xnor U5521 (N_5521,N_5321,N_5483);
nor U5522 (N_5522,N_5388,N_5467);
nand U5523 (N_5523,N_5274,N_5419);
nand U5524 (N_5524,N_5495,N_5374);
and U5525 (N_5525,N_5444,N_5327);
and U5526 (N_5526,N_5402,N_5316);
nand U5527 (N_5527,N_5310,N_5325);
nand U5528 (N_5528,N_5397,N_5358);
nor U5529 (N_5529,N_5272,N_5344);
and U5530 (N_5530,N_5418,N_5454);
xnor U5531 (N_5531,N_5257,N_5349);
and U5532 (N_5532,N_5267,N_5319);
xnor U5533 (N_5533,N_5357,N_5362);
nand U5534 (N_5534,N_5291,N_5400);
and U5535 (N_5535,N_5447,N_5346);
nor U5536 (N_5536,N_5392,N_5443);
xor U5537 (N_5537,N_5307,N_5343);
or U5538 (N_5538,N_5394,N_5498);
xor U5539 (N_5539,N_5445,N_5363);
xor U5540 (N_5540,N_5354,N_5422);
and U5541 (N_5541,N_5347,N_5297);
and U5542 (N_5542,N_5461,N_5414);
nand U5543 (N_5543,N_5377,N_5342);
nand U5544 (N_5544,N_5333,N_5281);
nand U5545 (N_5545,N_5389,N_5278);
nand U5546 (N_5546,N_5465,N_5390);
nand U5547 (N_5547,N_5289,N_5488);
or U5548 (N_5548,N_5283,N_5260);
or U5549 (N_5549,N_5350,N_5335);
nor U5550 (N_5550,N_5258,N_5370);
xnor U5551 (N_5551,N_5387,N_5271);
and U5552 (N_5552,N_5455,N_5412);
and U5553 (N_5553,N_5315,N_5373);
nand U5554 (N_5554,N_5279,N_5472);
and U5555 (N_5555,N_5337,N_5326);
nand U5556 (N_5556,N_5303,N_5417);
and U5557 (N_5557,N_5441,N_5460);
nor U5558 (N_5558,N_5314,N_5464);
and U5559 (N_5559,N_5288,N_5407);
or U5560 (N_5560,N_5481,N_5313);
and U5561 (N_5561,N_5427,N_5463);
nor U5562 (N_5562,N_5379,N_5375);
xor U5563 (N_5563,N_5384,N_5295);
and U5564 (N_5564,N_5442,N_5339);
or U5565 (N_5565,N_5446,N_5449);
and U5566 (N_5566,N_5280,N_5311);
xnor U5567 (N_5567,N_5491,N_5499);
nor U5568 (N_5568,N_5294,N_5256);
and U5569 (N_5569,N_5452,N_5406);
nor U5570 (N_5570,N_5391,N_5367);
or U5571 (N_5571,N_5360,N_5494);
nor U5572 (N_5572,N_5431,N_5398);
xnor U5573 (N_5573,N_5356,N_5298);
nand U5574 (N_5574,N_5415,N_5275);
nor U5575 (N_5575,N_5309,N_5476);
or U5576 (N_5576,N_5424,N_5404);
and U5577 (N_5577,N_5469,N_5497);
nor U5578 (N_5578,N_5355,N_5340);
nor U5579 (N_5579,N_5290,N_5277);
or U5580 (N_5580,N_5336,N_5474);
or U5581 (N_5581,N_5475,N_5383);
and U5582 (N_5582,N_5423,N_5433);
xnor U5583 (N_5583,N_5436,N_5334);
nor U5584 (N_5584,N_5284,N_5359);
xor U5585 (N_5585,N_5438,N_5351);
and U5586 (N_5586,N_5411,N_5471);
xnor U5587 (N_5587,N_5299,N_5261);
or U5588 (N_5588,N_5312,N_5403);
or U5589 (N_5589,N_5262,N_5493);
or U5590 (N_5590,N_5352,N_5338);
nor U5591 (N_5591,N_5268,N_5470);
or U5592 (N_5592,N_5269,N_5492);
or U5593 (N_5593,N_5426,N_5396);
nand U5594 (N_5594,N_5425,N_5259);
and U5595 (N_5595,N_5292,N_5485);
xnor U5596 (N_5596,N_5264,N_5348);
xor U5597 (N_5597,N_5496,N_5381);
and U5598 (N_5598,N_5486,N_5324);
xor U5599 (N_5599,N_5318,N_5399);
nor U5600 (N_5600,N_5473,N_5487);
xnor U5601 (N_5601,N_5304,N_5439);
nand U5602 (N_5602,N_5432,N_5254);
or U5603 (N_5603,N_5466,N_5285);
xnor U5604 (N_5604,N_5462,N_5468);
xor U5605 (N_5605,N_5409,N_5345);
xor U5606 (N_5606,N_5361,N_5332);
or U5607 (N_5607,N_5458,N_5308);
xnor U5608 (N_5608,N_5386,N_5305);
and U5609 (N_5609,N_5253,N_5369);
nor U5610 (N_5610,N_5420,N_5385);
nor U5611 (N_5611,N_5328,N_5331);
and U5612 (N_5612,N_5329,N_5456);
nand U5613 (N_5613,N_5450,N_5252);
or U5614 (N_5614,N_5364,N_5323);
xor U5615 (N_5615,N_5451,N_5296);
nand U5616 (N_5616,N_5365,N_5437);
nand U5617 (N_5617,N_5479,N_5300);
nor U5618 (N_5618,N_5416,N_5341);
nor U5619 (N_5619,N_5395,N_5382);
nor U5620 (N_5620,N_5435,N_5366);
xnor U5621 (N_5621,N_5301,N_5266);
or U5622 (N_5622,N_5489,N_5250);
nand U5623 (N_5623,N_5482,N_5282);
or U5624 (N_5624,N_5457,N_5293);
and U5625 (N_5625,N_5377,N_5319);
nor U5626 (N_5626,N_5361,N_5345);
xnor U5627 (N_5627,N_5463,N_5284);
or U5628 (N_5628,N_5455,N_5370);
nand U5629 (N_5629,N_5420,N_5462);
xnor U5630 (N_5630,N_5392,N_5251);
nand U5631 (N_5631,N_5362,N_5416);
nor U5632 (N_5632,N_5463,N_5436);
nor U5633 (N_5633,N_5393,N_5420);
and U5634 (N_5634,N_5426,N_5488);
and U5635 (N_5635,N_5260,N_5342);
nand U5636 (N_5636,N_5316,N_5326);
nand U5637 (N_5637,N_5488,N_5276);
or U5638 (N_5638,N_5403,N_5287);
xor U5639 (N_5639,N_5398,N_5256);
nor U5640 (N_5640,N_5302,N_5380);
nand U5641 (N_5641,N_5335,N_5355);
nand U5642 (N_5642,N_5452,N_5474);
nand U5643 (N_5643,N_5339,N_5446);
xnor U5644 (N_5644,N_5389,N_5470);
xor U5645 (N_5645,N_5337,N_5458);
or U5646 (N_5646,N_5432,N_5314);
nor U5647 (N_5647,N_5263,N_5375);
xnor U5648 (N_5648,N_5369,N_5260);
nor U5649 (N_5649,N_5390,N_5314);
nor U5650 (N_5650,N_5381,N_5403);
and U5651 (N_5651,N_5312,N_5453);
xnor U5652 (N_5652,N_5298,N_5447);
and U5653 (N_5653,N_5320,N_5462);
and U5654 (N_5654,N_5442,N_5462);
nand U5655 (N_5655,N_5436,N_5424);
nor U5656 (N_5656,N_5487,N_5434);
and U5657 (N_5657,N_5327,N_5277);
nand U5658 (N_5658,N_5277,N_5379);
and U5659 (N_5659,N_5381,N_5270);
xor U5660 (N_5660,N_5302,N_5281);
xor U5661 (N_5661,N_5412,N_5442);
xnor U5662 (N_5662,N_5315,N_5471);
and U5663 (N_5663,N_5410,N_5495);
and U5664 (N_5664,N_5394,N_5299);
and U5665 (N_5665,N_5423,N_5475);
or U5666 (N_5666,N_5255,N_5458);
nor U5667 (N_5667,N_5384,N_5495);
xnor U5668 (N_5668,N_5273,N_5433);
nor U5669 (N_5669,N_5337,N_5493);
nand U5670 (N_5670,N_5294,N_5479);
and U5671 (N_5671,N_5455,N_5422);
or U5672 (N_5672,N_5477,N_5473);
and U5673 (N_5673,N_5418,N_5311);
nor U5674 (N_5674,N_5351,N_5289);
xnor U5675 (N_5675,N_5429,N_5418);
nor U5676 (N_5676,N_5358,N_5445);
xor U5677 (N_5677,N_5429,N_5254);
and U5678 (N_5678,N_5326,N_5333);
or U5679 (N_5679,N_5261,N_5384);
or U5680 (N_5680,N_5444,N_5259);
nor U5681 (N_5681,N_5354,N_5402);
or U5682 (N_5682,N_5437,N_5366);
or U5683 (N_5683,N_5483,N_5490);
xnor U5684 (N_5684,N_5446,N_5322);
xnor U5685 (N_5685,N_5265,N_5394);
nor U5686 (N_5686,N_5426,N_5314);
and U5687 (N_5687,N_5440,N_5271);
xnor U5688 (N_5688,N_5389,N_5370);
xnor U5689 (N_5689,N_5408,N_5361);
or U5690 (N_5690,N_5264,N_5292);
xnor U5691 (N_5691,N_5378,N_5279);
or U5692 (N_5692,N_5254,N_5442);
nor U5693 (N_5693,N_5291,N_5425);
xor U5694 (N_5694,N_5372,N_5368);
or U5695 (N_5695,N_5265,N_5378);
nand U5696 (N_5696,N_5323,N_5336);
xor U5697 (N_5697,N_5253,N_5409);
xor U5698 (N_5698,N_5279,N_5411);
nand U5699 (N_5699,N_5450,N_5270);
nor U5700 (N_5700,N_5481,N_5316);
xor U5701 (N_5701,N_5375,N_5451);
and U5702 (N_5702,N_5277,N_5424);
nor U5703 (N_5703,N_5469,N_5258);
nand U5704 (N_5704,N_5392,N_5452);
or U5705 (N_5705,N_5258,N_5448);
or U5706 (N_5706,N_5328,N_5304);
nor U5707 (N_5707,N_5267,N_5386);
xor U5708 (N_5708,N_5253,N_5314);
xor U5709 (N_5709,N_5491,N_5298);
xnor U5710 (N_5710,N_5430,N_5342);
xnor U5711 (N_5711,N_5373,N_5395);
nor U5712 (N_5712,N_5308,N_5424);
or U5713 (N_5713,N_5450,N_5421);
nor U5714 (N_5714,N_5497,N_5393);
nor U5715 (N_5715,N_5490,N_5277);
nand U5716 (N_5716,N_5381,N_5298);
and U5717 (N_5717,N_5479,N_5487);
nor U5718 (N_5718,N_5376,N_5497);
xor U5719 (N_5719,N_5347,N_5321);
and U5720 (N_5720,N_5453,N_5348);
xnor U5721 (N_5721,N_5366,N_5423);
and U5722 (N_5722,N_5310,N_5347);
nand U5723 (N_5723,N_5499,N_5476);
nand U5724 (N_5724,N_5487,N_5312);
xor U5725 (N_5725,N_5254,N_5335);
or U5726 (N_5726,N_5427,N_5488);
xor U5727 (N_5727,N_5333,N_5368);
nand U5728 (N_5728,N_5339,N_5275);
nand U5729 (N_5729,N_5323,N_5280);
nor U5730 (N_5730,N_5460,N_5261);
or U5731 (N_5731,N_5255,N_5405);
and U5732 (N_5732,N_5318,N_5326);
or U5733 (N_5733,N_5432,N_5280);
and U5734 (N_5734,N_5366,N_5341);
and U5735 (N_5735,N_5446,N_5288);
and U5736 (N_5736,N_5435,N_5252);
or U5737 (N_5737,N_5342,N_5467);
nor U5738 (N_5738,N_5329,N_5420);
and U5739 (N_5739,N_5479,N_5459);
nand U5740 (N_5740,N_5305,N_5331);
xnor U5741 (N_5741,N_5395,N_5282);
xnor U5742 (N_5742,N_5466,N_5390);
nand U5743 (N_5743,N_5333,N_5263);
nor U5744 (N_5744,N_5452,N_5300);
xor U5745 (N_5745,N_5276,N_5402);
nand U5746 (N_5746,N_5333,N_5301);
or U5747 (N_5747,N_5357,N_5266);
and U5748 (N_5748,N_5429,N_5362);
and U5749 (N_5749,N_5488,N_5414);
or U5750 (N_5750,N_5642,N_5509);
nand U5751 (N_5751,N_5553,N_5731);
or U5752 (N_5752,N_5571,N_5663);
or U5753 (N_5753,N_5564,N_5609);
or U5754 (N_5754,N_5681,N_5607);
xor U5755 (N_5755,N_5540,N_5631);
nor U5756 (N_5756,N_5620,N_5599);
nand U5757 (N_5757,N_5649,N_5547);
and U5758 (N_5758,N_5656,N_5630);
xnor U5759 (N_5759,N_5559,N_5736);
or U5760 (N_5760,N_5622,N_5661);
and U5761 (N_5761,N_5659,N_5598);
nor U5762 (N_5762,N_5670,N_5569);
nand U5763 (N_5763,N_5733,N_5601);
nand U5764 (N_5764,N_5636,N_5665);
or U5765 (N_5765,N_5572,N_5512);
nor U5766 (N_5766,N_5685,N_5701);
and U5767 (N_5767,N_5632,N_5695);
nand U5768 (N_5768,N_5710,N_5618);
and U5769 (N_5769,N_5527,N_5592);
and U5770 (N_5770,N_5530,N_5662);
nand U5771 (N_5771,N_5664,N_5591);
nand U5772 (N_5772,N_5696,N_5721);
nor U5773 (N_5773,N_5674,N_5623);
xnor U5774 (N_5774,N_5600,N_5605);
nor U5775 (N_5775,N_5680,N_5703);
xnor U5776 (N_5776,N_5725,N_5699);
nand U5777 (N_5777,N_5708,N_5737);
or U5778 (N_5778,N_5522,N_5525);
and U5779 (N_5779,N_5686,N_5619);
or U5780 (N_5780,N_5552,N_5705);
and U5781 (N_5781,N_5560,N_5746);
nand U5782 (N_5782,N_5551,N_5612);
nand U5783 (N_5783,N_5748,N_5719);
or U5784 (N_5784,N_5727,N_5742);
nor U5785 (N_5785,N_5640,N_5513);
nand U5786 (N_5786,N_5570,N_5644);
and U5787 (N_5787,N_5712,N_5694);
xnor U5788 (N_5788,N_5668,N_5637);
and U5789 (N_5789,N_5543,N_5720);
or U5790 (N_5790,N_5741,N_5698);
xnor U5791 (N_5791,N_5511,N_5517);
and U5792 (N_5792,N_5690,N_5743);
and U5793 (N_5793,N_5647,N_5518);
nand U5794 (N_5794,N_5507,N_5654);
nor U5795 (N_5795,N_5613,N_5740);
xnor U5796 (N_5796,N_5526,N_5616);
nor U5797 (N_5797,N_5519,N_5542);
nand U5798 (N_5798,N_5505,N_5716);
or U5799 (N_5799,N_5538,N_5745);
xnor U5800 (N_5800,N_5626,N_5679);
nand U5801 (N_5801,N_5568,N_5523);
nand U5802 (N_5802,N_5545,N_5625);
nand U5803 (N_5803,N_5653,N_5520);
and U5804 (N_5804,N_5557,N_5735);
or U5805 (N_5805,N_5531,N_5641);
nand U5806 (N_5806,N_5728,N_5606);
and U5807 (N_5807,N_5580,N_5726);
nor U5808 (N_5808,N_5677,N_5702);
xor U5809 (N_5809,N_5666,N_5718);
xor U5810 (N_5810,N_5567,N_5658);
or U5811 (N_5811,N_5574,N_5585);
or U5812 (N_5812,N_5627,N_5575);
nor U5813 (N_5813,N_5500,N_5660);
or U5814 (N_5814,N_5744,N_5717);
and U5815 (N_5815,N_5675,N_5562);
or U5816 (N_5816,N_5515,N_5713);
and U5817 (N_5817,N_5628,N_5577);
and U5818 (N_5818,N_5581,N_5688);
and U5819 (N_5819,N_5617,N_5534);
and U5820 (N_5820,N_5673,N_5730);
nand U5821 (N_5821,N_5589,N_5536);
nand U5822 (N_5822,N_5638,N_5693);
nor U5823 (N_5823,N_5724,N_5516);
xnor U5824 (N_5824,N_5593,N_5529);
nor U5825 (N_5825,N_5706,N_5715);
nand U5826 (N_5826,N_5624,N_5588);
or U5827 (N_5827,N_5602,N_5645);
xnor U5828 (N_5828,N_5503,N_5597);
nor U5829 (N_5829,N_5683,N_5554);
nand U5830 (N_5830,N_5639,N_5603);
xor U5831 (N_5831,N_5711,N_5539);
and U5832 (N_5832,N_5544,N_5573);
nor U5833 (N_5833,N_5650,N_5729);
xnor U5834 (N_5834,N_5667,N_5652);
and U5835 (N_5835,N_5687,N_5689);
or U5836 (N_5836,N_5749,N_5556);
and U5837 (N_5837,N_5535,N_5566);
or U5838 (N_5838,N_5651,N_5576);
nand U5839 (N_5839,N_5524,N_5546);
xor U5840 (N_5840,N_5697,N_5594);
xnor U5841 (N_5841,N_5610,N_5558);
nand U5842 (N_5842,N_5508,N_5587);
nor U5843 (N_5843,N_5528,N_5604);
and U5844 (N_5844,N_5583,N_5676);
xnor U5845 (N_5845,N_5709,N_5596);
nand U5846 (N_5846,N_5504,N_5747);
or U5847 (N_5847,N_5657,N_5502);
nor U5848 (N_5848,N_5579,N_5646);
nor U5849 (N_5849,N_5578,N_5700);
nand U5850 (N_5850,N_5672,N_5608);
nor U5851 (N_5851,N_5648,N_5506);
or U5852 (N_5852,N_5738,N_5561);
nand U5853 (N_5853,N_5582,N_5643);
xor U5854 (N_5854,N_5684,N_5521);
xor U5855 (N_5855,N_5590,N_5707);
xor U5856 (N_5856,N_5537,N_5514);
and U5857 (N_5857,N_5669,N_5739);
nor U5858 (N_5858,N_5532,N_5533);
and U5859 (N_5859,N_5722,N_5615);
nor U5860 (N_5860,N_5614,N_5678);
nor U5861 (N_5861,N_5734,N_5565);
nor U5862 (N_5862,N_5563,N_5714);
and U5863 (N_5863,N_5548,N_5584);
or U5864 (N_5864,N_5541,N_5671);
nor U5865 (N_5865,N_5629,N_5691);
xor U5866 (N_5866,N_5692,N_5611);
and U5867 (N_5867,N_5655,N_5634);
or U5868 (N_5868,N_5510,N_5595);
nor U5869 (N_5869,N_5682,N_5635);
xnor U5870 (N_5870,N_5633,N_5501);
nand U5871 (N_5871,N_5586,N_5723);
or U5872 (N_5872,N_5549,N_5555);
xnor U5873 (N_5873,N_5621,N_5732);
or U5874 (N_5874,N_5704,N_5550);
or U5875 (N_5875,N_5521,N_5733);
xnor U5876 (N_5876,N_5745,N_5534);
nand U5877 (N_5877,N_5738,N_5669);
and U5878 (N_5878,N_5512,N_5641);
and U5879 (N_5879,N_5636,N_5744);
nor U5880 (N_5880,N_5516,N_5709);
xnor U5881 (N_5881,N_5523,N_5550);
nor U5882 (N_5882,N_5634,N_5742);
or U5883 (N_5883,N_5679,N_5737);
and U5884 (N_5884,N_5536,N_5645);
or U5885 (N_5885,N_5556,N_5721);
nor U5886 (N_5886,N_5718,N_5542);
nand U5887 (N_5887,N_5674,N_5562);
nor U5888 (N_5888,N_5548,N_5653);
xnor U5889 (N_5889,N_5585,N_5532);
xor U5890 (N_5890,N_5569,N_5533);
or U5891 (N_5891,N_5743,N_5612);
or U5892 (N_5892,N_5622,N_5663);
nor U5893 (N_5893,N_5686,N_5650);
and U5894 (N_5894,N_5504,N_5609);
and U5895 (N_5895,N_5636,N_5693);
and U5896 (N_5896,N_5709,N_5674);
xor U5897 (N_5897,N_5671,N_5675);
and U5898 (N_5898,N_5599,N_5708);
nand U5899 (N_5899,N_5665,N_5739);
nor U5900 (N_5900,N_5600,N_5644);
xor U5901 (N_5901,N_5703,N_5748);
nand U5902 (N_5902,N_5665,N_5584);
xor U5903 (N_5903,N_5747,N_5567);
or U5904 (N_5904,N_5719,N_5706);
nor U5905 (N_5905,N_5696,N_5727);
or U5906 (N_5906,N_5620,N_5748);
nand U5907 (N_5907,N_5696,N_5739);
xnor U5908 (N_5908,N_5601,N_5648);
xnor U5909 (N_5909,N_5561,N_5667);
xnor U5910 (N_5910,N_5578,N_5666);
nor U5911 (N_5911,N_5606,N_5627);
and U5912 (N_5912,N_5596,N_5647);
nand U5913 (N_5913,N_5731,N_5741);
or U5914 (N_5914,N_5533,N_5642);
nand U5915 (N_5915,N_5618,N_5517);
nand U5916 (N_5916,N_5731,N_5567);
nor U5917 (N_5917,N_5571,N_5502);
nor U5918 (N_5918,N_5602,N_5617);
xnor U5919 (N_5919,N_5554,N_5531);
xnor U5920 (N_5920,N_5579,N_5534);
and U5921 (N_5921,N_5627,N_5513);
or U5922 (N_5922,N_5588,N_5649);
nor U5923 (N_5923,N_5565,N_5558);
and U5924 (N_5924,N_5704,N_5748);
nand U5925 (N_5925,N_5662,N_5668);
nor U5926 (N_5926,N_5717,N_5627);
or U5927 (N_5927,N_5515,N_5516);
nand U5928 (N_5928,N_5637,N_5618);
xor U5929 (N_5929,N_5600,N_5574);
or U5930 (N_5930,N_5706,N_5627);
nand U5931 (N_5931,N_5660,N_5637);
nand U5932 (N_5932,N_5696,N_5638);
and U5933 (N_5933,N_5688,N_5744);
xnor U5934 (N_5934,N_5563,N_5575);
and U5935 (N_5935,N_5675,N_5531);
nor U5936 (N_5936,N_5518,N_5500);
xor U5937 (N_5937,N_5698,N_5613);
xor U5938 (N_5938,N_5685,N_5617);
or U5939 (N_5939,N_5572,N_5676);
nor U5940 (N_5940,N_5743,N_5510);
nand U5941 (N_5941,N_5626,N_5513);
and U5942 (N_5942,N_5644,N_5734);
or U5943 (N_5943,N_5601,N_5564);
and U5944 (N_5944,N_5578,N_5516);
or U5945 (N_5945,N_5660,N_5749);
nor U5946 (N_5946,N_5731,N_5530);
nand U5947 (N_5947,N_5574,N_5580);
and U5948 (N_5948,N_5541,N_5690);
nor U5949 (N_5949,N_5731,N_5582);
or U5950 (N_5950,N_5742,N_5565);
and U5951 (N_5951,N_5607,N_5635);
nor U5952 (N_5952,N_5630,N_5595);
or U5953 (N_5953,N_5735,N_5733);
or U5954 (N_5954,N_5657,N_5527);
and U5955 (N_5955,N_5623,N_5658);
and U5956 (N_5956,N_5635,N_5711);
nor U5957 (N_5957,N_5642,N_5579);
and U5958 (N_5958,N_5564,N_5649);
or U5959 (N_5959,N_5564,N_5673);
and U5960 (N_5960,N_5636,N_5707);
nor U5961 (N_5961,N_5748,N_5557);
xnor U5962 (N_5962,N_5628,N_5569);
nor U5963 (N_5963,N_5668,N_5575);
and U5964 (N_5964,N_5602,N_5547);
xor U5965 (N_5965,N_5501,N_5655);
nand U5966 (N_5966,N_5565,N_5501);
nand U5967 (N_5967,N_5571,N_5632);
xor U5968 (N_5968,N_5631,N_5515);
or U5969 (N_5969,N_5533,N_5695);
nor U5970 (N_5970,N_5718,N_5654);
and U5971 (N_5971,N_5617,N_5618);
and U5972 (N_5972,N_5532,N_5690);
nand U5973 (N_5973,N_5533,N_5614);
and U5974 (N_5974,N_5691,N_5728);
nor U5975 (N_5975,N_5733,N_5531);
nor U5976 (N_5976,N_5517,N_5625);
and U5977 (N_5977,N_5585,N_5534);
nand U5978 (N_5978,N_5691,N_5683);
xor U5979 (N_5979,N_5516,N_5737);
and U5980 (N_5980,N_5650,N_5677);
or U5981 (N_5981,N_5563,N_5600);
xor U5982 (N_5982,N_5502,N_5558);
or U5983 (N_5983,N_5689,N_5672);
and U5984 (N_5984,N_5528,N_5650);
nor U5985 (N_5985,N_5622,N_5600);
or U5986 (N_5986,N_5647,N_5694);
xnor U5987 (N_5987,N_5740,N_5691);
nor U5988 (N_5988,N_5614,N_5667);
nor U5989 (N_5989,N_5611,N_5735);
and U5990 (N_5990,N_5666,N_5625);
nand U5991 (N_5991,N_5715,N_5632);
or U5992 (N_5992,N_5569,N_5501);
nor U5993 (N_5993,N_5501,N_5621);
xor U5994 (N_5994,N_5626,N_5562);
nor U5995 (N_5995,N_5569,N_5506);
nor U5996 (N_5996,N_5659,N_5622);
and U5997 (N_5997,N_5709,N_5665);
or U5998 (N_5998,N_5503,N_5519);
or U5999 (N_5999,N_5643,N_5524);
or U6000 (N_6000,N_5833,N_5961);
nor U6001 (N_6001,N_5827,N_5960);
or U6002 (N_6002,N_5798,N_5926);
nor U6003 (N_6003,N_5794,N_5896);
xnor U6004 (N_6004,N_5964,N_5879);
or U6005 (N_6005,N_5868,N_5840);
or U6006 (N_6006,N_5807,N_5908);
and U6007 (N_6007,N_5828,N_5788);
or U6008 (N_6008,N_5915,N_5950);
xnor U6009 (N_6009,N_5822,N_5989);
and U6010 (N_6010,N_5824,N_5885);
xnor U6011 (N_6011,N_5831,N_5957);
xnor U6012 (N_6012,N_5948,N_5771);
and U6013 (N_6013,N_5834,N_5913);
or U6014 (N_6014,N_5803,N_5965);
nand U6015 (N_6015,N_5953,N_5871);
and U6016 (N_6016,N_5778,N_5990);
or U6017 (N_6017,N_5867,N_5914);
nand U6018 (N_6018,N_5789,N_5889);
xor U6019 (N_6019,N_5755,N_5762);
xor U6020 (N_6020,N_5882,N_5893);
nand U6021 (N_6021,N_5761,N_5928);
xnor U6022 (N_6022,N_5826,N_5797);
nor U6023 (N_6023,N_5765,N_5825);
xnor U6024 (N_6024,N_5808,N_5864);
nand U6025 (N_6025,N_5901,N_5830);
nor U6026 (N_6026,N_5924,N_5897);
and U6027 (N_6027,N_5891,N_5818);
nand U6028 (N_6028,N_5810,N_5854);
or U6029 (N_6029,N_5955,N_5836);
nor U6030 (N_6030,N_5768,N_5941);
nand U6031 (N_6031,N_5860,N_5995);
or U6032 (N_6032,N_5877,N_5863);
nor U6033 (N_6033,N_5951,N_5911);
and U6034 (N_6034,N_5750,N_5925);
xor U6035 (N_6035,N_5876,N_5967);
xor U6036 (N_6036,N_5886,N_5918);
and U6037 (N_6037,N_5804,N_5982);
or U6038 (N_6038,N_5958,N_5983);
or U6039 (N_6039,N_5784,N_5875);
nand U6040 (N_6040,N_5754,N_5832);
xor U6041 (N_6041,N_5992,N_5796);
and U6042 (N_6042,N_5841,N_5974);
or U6043 (N_6043,N_5997,N_5870);
or U6044 (N_6044,N_5900,N_5846);
nand U6045 (N_6045,N_5999,N_5902);
xor U6046 (N_6046,N_5776,N_5934);
xnor U6047 (N_6047,N_5952,N_5777);
or U6048 (N_6048,N_5976,N_5767);
or U6049 (N_6049,N_5869,N_5963);
and U6050 (N_6050,N_5987,N_5790);
nand U6051 (N_6051,N_5862,N_5922);
xnor U6052 (N_6052,N_5843,N_5758);
nand U6053 (N_6053,N_5785,N_5763);
xor U6054 (N_6054,N_5786,N_5929);
or U6055 (N_6055,N_5919,N_5799);
and U6056 (N_6056,N_5814,N_5975);
nor U6057 (N_6057,N_5887,N_5773);
xor U6058 (N_6058,N_5971,N_5966);
nand U6059 (N_6059,N_5943,N_5793);
and U6060 (N_6060,N_5993,N_5783);
xnor U6061 (N_6061,N_5935,N_5903);
nor U6062 (N_6062,N_5861,N_5855);
or U6063 (N_6063,N_5930,N_5751);
xor U6064 (N_6064,N_5851,N_5844);
nor U6065 (N_6065,N_5968,N_5984);
nor U6066 (N_6066,N_5812,N_5959);
xor U6067 (N_6067,N_5760,N_5837);
nand U6068 (N_6068,N_5939,N_5811);
and U6069 (N_6069,N_5838,N_5865);
xor U6070 (N_6070,N_5916,N_5931);
nor U6071 (N_6071,N_5806,N_5949);
nor U6072 (N_6072,N_5970,N_5848);
or U6073 (N_6073,N_5756,N_5782);
xor U6074 (N_6074,N_5892,N_5772);
nand U6075 (N_6075,N_5849,N_5937);
nand U6076 (N_6076,N_5839,N_5859);
nand U6077 (N_6077,N_5847,N_5759);
xor U6078 (N_6078,N_5853,N_5819);
xnor U6079 (N_6079,N_5775,N_5998);
and U6080 (N_6080,N_5947,N_5856);
or U6081 (N_6081,N_5991,N_5969);
and U6082 (N_6082,N_5821,N_5907);
nor U6083 (N_6083,N_5820,N_5816);
xnor U6084 (N_6084,N_5920,N_5766);
nor U6085 (N_6085,N_5800,N_5986);
xor U6086 (N_6086,N_5905,N_5792);
and U6087 (N_6087,N_5757,N_5904);
nor U6088 (N_6088,N_5888,N_5954);
nor U6089 (N_6089,N_5752,N_5942);
or U6090 (N_6090,N_5835,N_5764);
xor U6091 (N_6091,N_5972,N_5753);
nand U6092 (N_6092,N_5874,N_5917);
xor U6093 (N_6093,N_5817,N_5933);
nor U6094 (N_6094,N_5912,N_5858);
or U6095 (N_6095,N_5894,N_5770);
and U6096 (N_6096,N_5779,N_5805);
nand U6097 (N_6097,N_5890,N_5923);
or U6098 (N_6098,N_5781,N_5988);
nand U6099 (N_6099,N_5994,N_5980);
or U6100 (N_6100,N_5787,N_5866);
or U6101 (N_6101,N_5873,N_5791);
xnor U6102 (N_6102,N_5944,N_5978);
xnor U6103 (N_6103,N_5884,N_5979);
and U6104 (N_6104,N_5815,N_5850);
nand U6105 (N_6105,N_5977,N_5940);
xnor U6106 (N_6106,N_5956,N_5880);
or U6107 (N_6107,N_5938,N_5932);
and U6108 (N_6108,N_5899,N_5909);
nand U6109 (N_6109,N_5945,N_5829);
and U6110 (N_6110,N_5823,N_5946);
nor U6111 (N_6111,N_5985,N_5906);
xnor U6112 (N_6112,N_5883,N_5878);
xor U6113 (N_6113,N_5981,N_5962);
or U6114 (N_6114,N_5780,N_5910);
nand U6115 (N_6115,N_5898,N_5895);
xnor U6116 (N_6116,N_5845,N_5842);
xnor U6117 (N_6117,N_5973,N_5921);
xnor U6118 (N_6118,N_5801,N_5852);
nand U6119 (N_6119,N_5809,N_5813);
and U6120 (N_6120,N_5795,N_5872);
xor U6121 (N_6121,N_5774,N_5927);
and U6122 (N_6122,N_5936,N_5996);
and U6123 (N_6123,N_5802,N_5769);
nor U6124 (N_6124,N_5881,N_5857);
nor U6125 (N_6125,N_5982,N_5782);
and U6126 (N_6126,N_5757,N_5818);
and U6127 (N_6127,N_5944,N_5766);
nor U6128 (N_6128,N_5851,N_5905);
xnor U6129 (N_6129,N_5759,N_5851);
and U6130 (N_6130,N_5817,N_5833);
nand U6131 (N_6131,N_5986,N_5861);
and U6132 (N_6132,N_5957,N_5807);
or U6133 (N_6133,N_5875,N_5764);
or U6134 (N_6134,N_5900,N_5947);
nand U6135 (N_6135,N_5870,N_5782);
nand U6136 (N_6136,N_5768,N_5790);
or U6137 (N_6137,N_5888,N_5821);
and U6138 (N_6138,N_5781,N_5766);
nor U6139 (N_6139,N_5898,N_5992);
or U6140 (N_6140,N_5885,N_5756);
nor U6141 (N_6141,N_5995,N_5895);
or U6142 (N_6142,N_5976,N_5788);
xnor U6143 (N_6143,N_5868,N_5917);
nand U6144 (N_6144,N_5853,N_5856);
xnor U6145 (N_6145,N_5765,N_5794);
xnor U6146 (N_6146,N_5872,N_5820);
nand U6147 (N_6147,N_5764,N_5896);
nand U6148 (N_6148,N_5871,N_5806);
and U6149 (N_6149,N_5836,N_5811);
nor U6150 (N_6150,N_5809,N_5996);
nor U6151 (N_6151,N_5775,N_5919);
nor U6152 (N_6152,N_5831,N_5778);
nand U6153 (N_6153,N_5882,N_5939);
nand U6154 (N_6154,N_5908,N_5819);
xnor U6155 (N_6155,N_5851,N_5798);
xnor U6156 (N_6156,N_5771,N_5790);
or U6157 (N_6157,N_5981,N_5951);
nand U6158 (N_6158,N_5877,N_5953);
and U6159 (N_6159,N_5867,N_5885);
and U6160 (N_6160,N_5785,N_5891);
and U6161 (N_6161,N_5768,N_5924);
or U6162 (N_6162,N_5966,N_5989);
and U6163 (N_6163,N_5750,N_5927);
nand U6164 (N_6164,N_5919,N_5961);
or U6165 (N_6165,N_5859,N_5868);
or U6166 (N_6166,N_5875,N_5935);
or U6167 (N_6167,N_5989,N_5958);
and U6168 (N_6168,N_5897,N_5797);
or U6169 (N_6169,N_5810,N_5929);
and U6170 (N_6170,N_5950,N_5982);
nor U6171 (N_6171,N_5944,N_5801);
nor U6172 (N_6172,N_5804,N_5840);
xnor U6173 (N_6173,N_5808,N_5901);
nor U6174 (N_6174,N_5806,N_5969);
nand U6175 (N_6175,N_5808,N_5989);
and U6176 (N_6176,N_5912,N_5951);
or U6177 (N_6177,N_5940,N_5933);
nor U6178 (N_6178,N_5760,N_5751);
and U6179 (N_6179,N_5931,N_5767);
or U6180 (N_6180,N_5772,N_5782);
and U6181 (N_6181,N_5800,N_5983);
nor U6182 (N_6182,N_5884,N_5770);
nand U6183 (N_6183,N_5942,N_5963);
xor U6184 (N_6184,N_5877,N_5856);
xnor U6185 (N_6185,N_5800,N_5804);
xnor U6186 (N_6186,N_5779,N_5914);
xnor U6187 (N_6187,N_5956,N_5895);
or U6188 (N_6188,N_5943,N_5957);
and U6189 (N_6189,N_5788,N_5897);
nor U6190 (N_6190,N_5880,N_5756);
or U6191 (N_6191,N_5942,N_5960);
xor U6192 (N_6192,N_5799,N_5792);
and U6193 (N_6193,N_5827,N_5794);
and U6194 (N_6194,N_5904,N_5809);
and U6195 (N_6195,N_5895,N_5801);
xnor U6196 (N_6196,N_5900,N_5774);
and U6197 (N_6197,N_5955,N_5968);
and U6198 (N_6198,N_5801,N_5837);
or U6199 (N_6199,N_5998,N_5855);
or U6200 (N_6200,N_5920,N_5850);
and U6201 (N_6201,N_5855,N_5979);
or U6202 (N_6202,N_5991,N_5947);
nor U6203 (N_6203,N_5990,N_5915);
xnor U6204 (N_6204,N_5852,N_5849);
nor U6205 (N_6205,N_5753,N_5965);
xor U6206 (N_6206,N_5823,N_5752);
nor U6207 (N_6207,N_5775,N_5932);
xnor U6208 (N_6208,N_5975,N_5877);
or U6209 (N_6209,N_5903,N_5898);
nor U6210 (N_6210,N_5790,N_5900);
and U6211 (N_6211,N_5972,N_5854);
xor U6212 (N_6212,N_5973,N_5996);
and U6213 (N_6213,N_5773,N_5892);
nand U6214 (N_6214,N_5925,N_5903);
xor U6215 (N_6215,N_5913,N_5794);
nand U6216 (N_6216,N_5802,N_5915);
xnor U6217 (N_6217,N_5802,N_5816);
nand U6218 (N_6218,N_5982,N_5893);
xor U6219 (N_6219,N_5805,N_5794);
or U6220 (N_6220,N_5793,N_5900);
or U6221 (N_6221,N_5950,N_5951);
nand U6222 (N_6222,N_5760,N_5936);
xor U6223 (N_6223,N_5755,N_5750);
nand U6224 (N_6224,N_5943,N_5932);
and U6225 (N_6225,N_5920,N_5915);
and U6226 (N_6226,N_5977,N_5884);
nand U6227 (N_6227,N_5758,N_5958);
nor U6228 (N_6228,N_5846,N_5953);
or U6229 (N_6229,N_5760,N_5985);
nor U6230 (N_6230,N_5935,N_5787);
xnor U6231 (N_6231,N_5771,N_5926);
nand U6232 (N_6232,N_5883,N_5961);
or U6233 (N_6233,N_5767,N_5773);
nand U6234 (N_6234,N_5795,N_5890);
nor U6235 (N_6235,N_5812,N_5753);
and U6236 (N_6236,N_5828,N_5882);
or U6237 (N_6237,N_5799,N_5939);
and U6238 (N_6238,N_5916,N_5993);
nand U6239 (N_6239,N_5882,N_5958);
or U6240 (N_6240,N_5814,N_5777);
nand U6241 (N_6241,N_5947,N_5925);
nand U6242 (N_6242,N_5975,N_5960);
nand U6243 (N_6243,N_5862,N_5812);
xor U6244 (N_6244,N_5787,N_5902);
or U6245 (N_6245,N_5923,N_5807);
nand U6246 (N_6246,N_5888,N_5794);
and U6247 (N_6247,N_5873,N_5802);
or U6248 (N_6248,N_5846,N_5793);
and U6249 (N_6249,N_5942,N_5781);
or U6250 (N_6250,N_6127,N_6240);
or U6251 (N_6251,N_6070,N_6122);
and U6252 (N_6252,N_6158,N_6106);
and U6253 (N_6253,N_6123,N_6237);
nor U6254 (N_6254,N_6246,N_6110);
nand U6255 (N_6255,N_6193,N_6002);
and U6256 (N_6256,N_6149,N_6133);
nand U6257 (N_6257,N_6040,N_6215);
or U6258 (N_6258,N_6170,N_6155);
or U6259 (N_6259,N_6136,N_6147);
or U6260 (N_6260,N_6128,N_6053);
and U6261 (N_6261,N_6081,N_6164);
and U6262 (N_6262,N_6118,N_6238);
and U6263 (N_6263,N_6068,N_6163);
nand U6264 (N_6264,N_6066,N_6161);
and U6265 (N_6265,N_6013,N_6176);
nor U6266 (N_6266,N_6172,N_6138);
and U6267 (N_6267,N_6220,N_6219);
and U6268 (N_6268,N_6005,N_6047);
nor U6269 (N_6269,N_6062,N_6055);
and U6270 (N_6270,N_6025,N_6229);
nor U6271 (N_6271,N_6049,N_6144);
nand U6272 (N_6272,N_6096,N_6145);
nor U6273 (N_6273,N_6212,N_6042);
nor U6274 (N_6274,N_6208,N_6109);
or U6275 (N_6275,N_6031,N_6200);
nand U6276 (N_6276,N_6190,N_6232);
or U6277 (N_6277,N_6023,N_6192);
nor U6278 (N_6278,N_6157,N_6179);
xnor U6279 (N_6279,N_6035,N_6195);
xor U6280 (N_6280,N_6223,N_6084);
or U6281 (N_6281,N_6079,N_6146);
and U6282 (N_6282,N_6159,N_6218);
nand U6283 (N_6283,N_6078,N_6196);
nor U6284 (N_6284,N_6236,N_6225);
xnor U6285 (N_6285,N_6139,N_6117);
nor U6286 (N_6286,N_6069,N_6168);
and U6287 (N_6287,N_6227,N_6071);
and U6288 (N_6288,N_6050,N_6124);
nor U6289 (N_6289,N_6171,N_6051);
nand U6290 (N_6290,N_6248,N_6156);
and U6291 (N_6291,N_6173,N_6082);
or U6292 (N_6292,N_6222,N_6119);
or U6293 (N_6293,N_6043,N_6113);
and U6294 (N_6294,N_6152,N_6150);
and U6295 (N_6295,N_6239,N_6142);
nor U6296 (N_6296,N_6107,N_6014);
nand U6297 (N_6297,N_6009,N_6131);
nand U6298 (N_6298,N_6210,N_6092);
nand U6299 (N_6299,N_6036,N_6003);
xnor U6300 (N_6300,N_6094,N_6116);
nand U6301 (N_6301,N_6089,N_6058);
or U6302 (N_6302,N_6194,N_6045);
xnor U6303 (N_6303,N_6126,N_6008);
nand U6304 (N_6304,N_6199,N_6201);
or U6305 (N_6305,N_6143,N_6244);
nor U6306 (N_6306,N_6102,N_6216);
nor U6307 (N_6307,N_6234,N_6203);
and U6308 (N_6308,N_6108,N_6099);
nand U6309 (N_6309,N_6182,N_6028);
xor U6310 (N_6310,N_6174,N_6075);
or U6311 (N_6311,N_6076,N_6016);
nor U6312 (N_6312,N_6154,N_6022);
or U6313 (N_6313,N_6024,N_6202);
nor U6314 (N_6314,N_6186,N_6226);
and U6315 (N_6315,N_6129,N_6006);
and U6316 (N_6316,N_6130,N_6034);
nand U6317 (N_6317,N_6011,N_6233);
nor U6318 (N_6318,N_6048,N_6015);
xor U6319 (N_6319,N_6057,N_6000);
and U6320 (N_6320,N_6169,N_6114);
xor U6321 (N_6321,N_6032,N_6181);
nor U6322 (N_6322,N_6039,N_6166);
or U6323 (N_6323,N_6019,N_6178);
and U6324 (N_6324,N_6044,N_6197);
xnor U6325 (N_6325,N_6067,N_6162);
xnor U6326 (N_6326,N_6007,N_6137);
nand U6327 (N_6327,N_6101,N_6148);
nand U6328 (N_6328,N_6141,N_6091);
or U6329 (N_6329,N_6018,N_6213);
nand U6330 (N_6330,N_6121,N_6065);
xor U6331 (N_6331,N_6090,N_6249);
nor U6332 (N_6332,N_6242,N_6105);
xnor U6333 (N_6333,N_6231,N_6061);
nor U6334 (N_6334,N_6093,N_6205);
nand U6335 (N_6335,N_6017,N_6206);
or U6336 (N_6336,N_6098,N_6010);
or U6337 (N_6337,N_6020,N_6054);
xor U6338 (N_6338,N_6247,N_6088);
nor U6339 (N_6339,N_6103,N_6185);
nand U6340 (N_6340,N_6080,N_6207);
xor U6341 (N_6341,N_6132,N_6027);
or U6342 (N_6342,N_6060,N_6187);
xor U6343 (N_6343,N_6063,N_6073);
nand U6344 (N_6344,N_6104,N_6064);
nor U6345 (N_6345,N_6224,N_6097);
or U6346 (N_6346,N_6086,N_6217);
xnor U6347 (N_6347,N_6189,N_6111);
and U6348 (N_6348,N_6134,N_6112);
or U6349 (N_6349,N_6165,N_6140);
or U6350 (N_6350,N_6026,N_6211);
nor U6351 (N_6351,N_6085,N_6183);
xor U6352 (N_6352,N_6241,N_6184);
and U6353 (N_6353,N_6243,N_6021);
nor U6354 (N_6354,N_6072,N_6160);
nand U6355 (N_6355,N_6030,N_6214);
or U6356 (N_6356,N_6230,N_6052);
and U6357 (N_6357,N_6221,N_6175);
xnor U6358 (N_6358,N_6245,N_6115);
nor U6359 (N_6359,N_6188,N_6125);
nand U6360 (N_6360,N_6059,N_6180);
or U6361 (N_6361,N_6191,N_6135);
xnor U6362 (N_6362,N_6012,N_6100);
or U6363 (N_6363,N_6153,N_6177);
nand U6364 (N_6364,N_6204,N_6235);
and U6365 (N_6365,N_6083,N_6004);
and U6366 (N_6366,N_6041,N_6001);
nand U6367 (N_6367,N_6056,N_6087);
xor U6368 (N_6368,N_6077,N_6046);
xor U6369 (N_6369,N_6038,N_6033);
and U6370 (N_6370,N_6095,N_6167);
and U6371 (N_6371,N_6228,N_6198);
and U6372 (N_6372,N_6209,N_6120);
or U6373 (N_6373,N_6037,N_6151);
nand U6374 (N_6374,N_6074,N_6029);
nor U6375 (N_6375,N_6083,N_6021);
or U6376 (N_6376,N_6241,N_6068);
xnor U6377 (N_6377,N_6135,N_6147);
or U6378 (N_6378,N_6118,N_6224);
nand U6379 (N_6379,N_6014,N_6229);
nand U6380 (N_6380,N_6152,N_6001);
nor U6381 (N_6381,N_6083,N_6163);
or U6382 (N_6382,N_6071,N_6001);
xor U6383 (N_6383,N_6115,N_6184);
and U6384 (N_6384,N_6226,N_6080);
or U6385 (N_6385,N_6200,N_6131);
or U6386 (N_6386,N_6191,N_6107);
nand U6387 (N_6387,N_6204,N_6209);
and U6388 (N_6388,N_6032,N_6154);
xnor U6389 (N_6389,N_6167,N_6140);
and U6390 (N_6390,N_6161,N_6228);
nand U6391 (N_6391,N_6053,N_6015);
xor U6392 (N_6392,N_6123,N_6248);
or U6393 (N_6393,N_6248,N_6174);
nand U6394 (N_6394,N_6114,N_6096);
and U6395 (N_6395,N_6022,N_6095);
xnor U6396 (N_6396,N_6105,N_6010);
or U6397 (N_6397,N_6238,N_6150);
and U6398 (N_6398,N_6188,N_6046);
and U6399 (N_6399,N_6151,N_6020);
xor U6400 (N_6400,N_6017,N_6102);
and U6401 (N_6401,N_6122,N_6148);
xnor U6402 (N_6402,N_6211,N_6150);
nand U6403 (N_6403,N_6228,N_6159);
and U6404 (N_6404,N_6233,N_6183);
xor U6405 (N_6405,N_6071,N_6239);
nor U6406 (N_6406,N_6064,N_6248);
nor U6407 (N_6407,N_6190,N_6165);
nand U6408 (N_6408,N_6194,N_6208);
and U6409 (N_6409,N_6130,N_6206);
xnor U6410 (N_6410,N_6006,N_6170);
or U6411 (N_6411,N_6058,N_6217);
nor U6412 (N_6412,N_6153,N_6183);
nand U6413 (N_6413,N_6114,N_6218);
or U6414 (N_6414,N_6100,N_6025);
and U6415 (N_6415,N_6068,N_6015);
nand U6416 (N_6416,N_6235,N_6055);
xor U6417 (N_6417,N_6086,N_6249);
and U6418 (N_6418,N_6020,N_6012);
nor U6419 (N_6419,N_6067,N_6113);
or U6420 (N_6420,N_6008,N_6229);
nand U6421 (N_6421,N_6203,N_6135);
nand U6422 (N_6422,N_6089,N_6068);
or U6423 (N_6423,N_6145,N_6174);
nor U6424 (N_6424,N_6052,N_6108);
nand U6425 (N_6425,N_6063,N_6168);
or U6426 (N_6426,N_6014,N_6122);
xor U6427 (N_6427,N_6121,N_6213);
or U6428 (N_6428,N_6146,N_6125);
nand U6429 (N_6429,N_6244,N_6167);
and U6430 (N_6430,N_6024,N_6034);
or U6431 (N_6431,N_6238,N_6077);
nor U6432 (N_6432,N_6142,N_6044);
nand U6433 (N_6433,N_6081,N_6178);
and U6434 (N_6434,N_6101,N_6131);
or U6435 (N_6435,N_6140,N_6128);
nor U6436 (N_6436,N_6193,N_6149);
or U6437 (N_6437,N_6012,N_6071);
nand U6438 (N_6438,N_6036,N_6239);
xnor U6439 (N_6439,N_6216,N_6142);
nand U6440 (N_6440,N_6151,N_6051);
and U6441 (N_6441,N_6113,N_6237);
nand U6442 (N_6442,N_6111,N_6169);
and U6443 (N_6443,N_6156,N_6043);
xor U6444 (N_6444,N_6019,N_6114);
and U6445 (N_6445,N_6074,N_6042);
nor U6446 (N_6446,N_6088,N_6011);
nor U6447 (N_6447,N_6206,N_6209);
xor U6448 (N_6448,N_6122,N_6117);
nand U6449 (N_6449,N_6020,N_6185);
xnor U6450 (N_6450,N_6212,N_6002);
nor U6451 (N_6451,N_6123,N_6091);
xor U6452 (N_6452,N_6082,N_6193);
or U6453 (N_6453,N_6204,N_6172);
xnor U6454 (N_6454,N_6115,N_6193);
and U6455 (N_6455,N_6093,N_6192);
nor U6456 (N_6456,N_6180,N_6230);
or U6457 (N_6457,N_6016,N_6182);
and U6458 (N_6458,N_6157,N_6222);
and U6459 (N_6459,N_6148,N_6092);
and U6460 (N_6460,N_6066,N_6214);
and U6461 (N_6461,N_6165,N_6136);
nor U6462 (N_6462,N_6118,N_6173);
nor U6463 (N_6463,N_6158,N_6149);
nor U6464 (N_6464,N_6224,N_6203);
xnor U6465 (N_6465,N_6246,N_6195);
nor U6466 (N_6466,N_6237,N_6053);
and U6467 (N_6467,N_6145,N_6042);
and U6468 (N_6468,N_6192,N_6055);
and U6469 (N_6469,N_6229,N_6248);
or U6470 (N_6470,N_6218,N_6134);
xor U6471 (N_6471,N_6208,N_6068);
and U6472 (N_6472,N_6221,N_6166);
nand U6473 (N_6473,N_6086,N_6234);
or U6474 (N_6474,N_6170,N_6148);
and U6475 (N_6475,N_6125,N_6156);
xor U6476 (N_6476,N_6031,N_6113);
nand U6477 (N_6477,N_6057,N_6106);
and U6478 (N_6478,N_6103,N_6232);
nor U6479 (N_6479,N_6051,N_6011);
and U6480 (N_6480,N_6110,N_6217);
nor U6481 (N_6481,N_6144,N_6040);
or U6482 (N_6482,N_6079,N_6222);
xor U6483 (N_6483,N_6229,N_6141);
and U6484 (N_6484,N_6003,N_6170);
and U6485 (N_6485,N_6098,N_6156);
nand U6486 (N_6486,N_6077,N_6009);
or U6487 (N_6487,N_6203,N_6198);
nand U6488 (N_6488,N_6207,N_6055);
nor U6489 (N_6489,N_6227,N_6015);
xnor U6490 (N_6490,N_6043,N_6129);
and U6491 (N_6491,N_6190,N_6111);
nor U6492 (N_6492,N_6206,N_6029);
xnor U6493 (N_6493,N_6187,N_6061);
nand U6494 (N_6494,N_6083,N_6008);
nor U6495 (N_6495,N_6038,N_6157);
and U6496 (N_6496,N_6087,N_6205);
or U6497 (N_6497,N_6122,N_6030);
and U6498 (N_6498,N_6164,N_6235);
nand U6499 (N_6499,N_6001,N_6101);
nand U6500 (N_6500,N_6284,N_6390);
nor U6501 (N_6501,N_6453,N_6342);
nor U6502 (N_6502,N_6369,N_6444);
xnor U6503 (N_6503,N_6330,N_6278);
or U6504 (N_6504,N_6340,N_6266);
and U6505 (N_6505,N_6480,N_6384);
nand U6506 (N_6506,N_6479,N_6419);
nor U6507 (N_6507,N_6304,N_6485);
nand U6508 (N_6508,N_6375,N_6397);
nand U6509 (N_6509,N_6407,N_6422);
xnor U6510 (N_6510,N_6337,N_6403);
nor U6511 (N_6511,N_6484,N_6400);
and U6512 (N_6512,N_6425,N_6416);
xor U6513 (N_6513,N_6296,N_6410);
xor U6514 (N_6514,N_6260,N_6309);
or U6515 (N_6515,N_6362,N_6415);
or U6516 (N_6516,N_6414,N_6336);
nand U6517 (N_6517,N_6273,N_6412);
or U6518 (N_6518,N_6282,N_6382);
and U6519 (N_6519,N_6316,N_6460);
xnor U6520 (N_6520,N_6344,N_6314);
and U6521 (N_6521,N_6417,N_6276);
or U6522 (N_6522,N_6264,N_6277);
and U6523 (N_6523,N_6457,N_6478);
nand U6524 (N_6524,N_6379,N_6312);
and U6525 (N_6525,N_6474,N_6321);
nor U6526 (N_6526,N_6315,N_6499);
or U6527 (N_6527,N_6476,N_6353);
or U6528 (N_6528,N_6385,N_6424);
nand U6529 (N_6529,N_6324,N_6274);
and U6530 (N_6530,N_6402,N_6252);
xor U6531 (N_6531,N_6463,N_6395);
or U6532 (N_6532,N_6438,N_6448);
xor U6533 (N_6533,N_6263,N_6470);
nor U6534 (N_6534,N_6280,N_6387);
nand U6535 (N_6535,N_6318,N_6398);
nand U6536 (N_6536,N_6350,N_6446);
nor U6537 (N_6537,N_6366,N_6386);
xnor U6538 (N_6538,N_6449,N_6396);
and U6539 (N_6539,N_6404,N_6394);
nor U6540 (N_6540,N_6334,N_6421);
or U6541 (N_6541,N_6360,N_6466);
and U6542 (N_6542,N_6465,N_6311);
and U6543 (N_6543,N_6468,N_6301);
or U6544 (N_6544,N_6496,N_6456);
or U6545 (N_6545,N_6347,N_6488);
nand U6546 (N_6546,N_6430,N_6335);
xor U6547 (N_6547,N_6307,N_6391);
or U6548 (N_6548,N_6420,N_6493);
xnor U6549 (N_6549,N_6310,N_6423);
xor U6550 (N_6550,N_6303,N_6445);
nor U6551 (N_6551,N_6472,N_6408);
xnor U6552 (N_6552,N_6329,N_6254);
or U6553 (N_6553,N_6464,N_6434);
nor U6554 (N_6554,N_6482,N_6367);
and U6555 (N_6555,N_6346,N_6442);
or U6556 (N_6556,N_6487,N_6295);
xor U6557 (N_6557,N_6343,N_6411);
or U6558 (N_6558,N_6495,N_6293);
nand U6559 (N_6559,N_6306,N_6376);
and U6560 (N_6560,N_6297,N_6327);
nor U6561 (N_6561,N_6418,N_6257);
and U6562 (N_6562,N_6298,N_6462);
and U6563 (N_6563,N_6497,N_6440);
or U6564 (N_6564,N_6255,N_6270);
or U6565 (N_6565,N_6291,N_6331);
nand U6566 (N_6566,N_6355,N_6299);
and U6567 (N_6567,N_6392,N_6409);
nor U6568 (N_6568,N_6380,N_6313);
nand U6569 (N_6569,N_6377,N_6427);
nor U6570 (N_6570,N_6486,N_6426);
xnor U6571 (N_6571,N_6439,N_6326);
nor U6572 (N_6572,N_6250,N_6477);
nand U6573 (N_6573,N_6429,N_6364);
xor U6574 (N_6574,N_6428,N_6268);
nand U6575 (N_6575,N_6262,N_6374);
xnor U6576 (N_6576,N_6498,N_6283);
xnor U6577 (N_6577,N_6437,N_6305);
or U6578 (N_6578,N_6467,N_6454);
nor U6579 (N_6579,N_6272,N_6302);
nand U6580 (N_6580,N_6450,N_6265);
and U6581 (N_6581,N_6461,N_6363);
nand U6582 (N_6582,N_6333,N_6361);
or U6583 (N_6583,N_6368,N_6287);
nor U6584 (N_6584,N_6251,N_6458);
nor U6585 (N_6585,N_6253,N_6459);
xnor U6586 (N_6586,N_6483,N_6443);
and U6587 (N_6587,N_6383,N_6317);
nor U6588 (N_6588,N_6341,N_6288);
nor U6589 (N_6589,N_6285,N_6351);
or U6590 (N_6590,N_6256,N_6381);
and U6591 (N_6591,N_6399,N_6371);
nand U6592 (N_6592,N_6332,N_6328);
or U6593 (N_6593,N_6389,N_6432);
nand U6594 (N_6594,N_6469,N_6365);
xor U6595 (N_6595,N_6373,N_6441);
nor U6596 (N_6596,N_6357,N_6473);
and U6597 (N_6597,N_6300,N_6406);
nand U6598 (N_6598,N_6294,N_6352);
nor U6599 (N_6599,N_6359,N_6271);
nor U6600 (N_6600,N_6281,N_6322);
xnor U6601 (N_6601,N_6378,N_6475);
and U6602 (N_6602,N_6492,N_6491);
nand U6603 (N_6603,N_6435,N_6258);
xnor U6604 (N_6604,N_6481,N_6490);
nand U6605 (N_6605,N_6323,N_6289);
nand U6606 (N_6606,N_6471,N_6405);
and U6607 (N_6607,N_6356,N_6279);
xnor U6608 (N_6608,N_6290,N_6269);
or U6609 (N_6609,N_6372,N_6286);
nor U6610 (N_6610,N_6308,N_6358);
and U6611 (N_6611,N_6354,N_6455);
and U6612 (N_6612,N_6261,N_6348);
and U6613 (N_6613,N_6401,N_6292);
and U6614 (N_6614,N_6393,N_6259);
and U6615 (N_6615,N_6320,N_6275);
xnor U6616 (N_6616,N_6433,N_6267);
nor U6617 (N_6617,N_6489,N_6451);
or U6618 (N_6618,N_6345,N_6319);
nor U6619 (N_6619,N_6338,N_6447);
nor U6620 (N_6620,N_6431,N_6370);
or U6621 (N_6621,N_6325,N_6339);
xnor U6622 (N_6622,N_6436,N_6413);
or U6623 (N_6623,N_6388,N_6452);
nor U6624 (N_6624,N_6494,N_6349);
xor U6625 (N_6625,N_6379,N_6367);
nand U6626 (N_6626,N_6295,N_6491);
and U6627 (N_6627,N_6475,N_6278);
nand U6628 (N_6628,N_6445,N_6414);
nand U6629 (N_6629,N_6333,N_6260);
and U6630 (N_6630,N_6391,N_6471);
or U6631 (N_6631,N_6330,N_6456);
and U6632 (N_6632,N_6350,N_6415);
nor U6633 (N_6633,N_6486,N_6380);
nor U6634 (N_6634,N_6367,N_6497);
or U6635 (N_6635,N_6328,N_6304);
or U6636 (N_6636,N_6330,N_6311);
xnor U6637 (N_6637,N_6315,N_6343);
or U6638 (N_6638,N_6316,N_6313);
nor U6639 (N_6639,N_6379,N_6365);
and U6640 (N_6640,N_6390,N_6440);
nand U6641 (N_6641,N_6297,N_6272);
xnor U6642 (N_6642,N_6305,N_6415);
and U6643 (N_6643,N_6399,N_6429);
or U6644 (N_6644,N_6447,N_6484);
and U6645 (N_6645,N_6399,N_6433);
nand U6646 (N_6646,N_6386,N_6442);
and U6647 (N_6647,N_6269,N_6489);
or U6648 (N_6648,N_6302,N_6441);
nand U6649 (N_6649,N_6479,N_6496);
and U6650 (N_6650,N_6263,N_6315);
nor U6651 (N_6651,N_6498,N_6477);
and U6652 (N_6652,N_6454,N_6452);
xor U6653 (N_6653,N_6325,N_6491);
xor U6654 (N_6654,N_6297,N_6373);
and U6655 (N_6655,N_6291,N_6305);
xnor U6656 (N_6656,N_6336,N_6388);
nand U6657 (N_6657,N_6356,N_6403);
and U6658 (N_6658,N_6391,N_6481);
and U6659 (N_6659,N_6429,N_6390);
and U6660 (N_6660,N_6418,N_6323);
nor U6661 (N_6661,N_6407,N_6498);
xor U6662 (N_6662,N_6331,N_6420);
nor U6663 (N_6663,N_6482,N_6274);
nand U6664 (N_6664,N_6467,N_6344);
and U6665 (N_6665,N_6413,N_6334);
nand U6666 (N_6666,N_6281,N_6354);
nor U6667 (N_6667,N_6358,N_6368);
nand U6668 (N_6668,N_6487,N_6358);
nor U6669 (N_6669,N_6445,N_6476);
nor U6670 (N_6670,N_6365,N_6329);
xor U6671 (N_6671,N_6458,N_6310);
or U6672 (N_6672,N_6441,N_6399);
nand U6673 (N_6673,N_6419,N_6318);
and U6674 (N_6674,N_6496,N_6499);
or U6675 (N_6675,N_6293,N_6320);
xor U6676 (N_6676,N_6288,N_6475);
or U6677 (N_6677,N_6329,N_6343);
or U6678 (N_6678,N_6251,N_6479);
xnor U6679 (N_6679,N_6371,N_6251);
and U6680 (N_6680,N_6331,N_6377);
and U6681 (N_6681,N_6264,N_6289);
nand U6682 (N_6682,N_6393,N_6366);
or U6683 (N_6683,N_6442,N_6380);
xor U6684 (N_6684,N_6496,N_6339);
xor U6685 (N_6685,N_6473,N_6489);
xor U6686 (N_6686,N_6439,N_6397);
xnor U6687 (N_6687,N_6291,N_6416);
nand U6688 (N_6688,N_6283,N_6472);
and U6689 (N_6689,N_6330,N_6424);
and U6690 (N_6690,N_6317,N_6377);
xor U6691 (N_6691,N_6444,N_6366);
nor U6692 (N_6692,N_6355,N_6366);
xor U6693 (N_6693,N_6348,N_6317);
nand U6694 (N_6694,N_6360,N_6426);
nand U6695 (N_6695,N_6476,N_6338);
nand U6696 (N_6696,N_6487,N_6481);
nand U6697 (N_6697,N_6478,N_6293);
xor U6698 (N_6698,N_6294,N_6355);
or U6699 (N_6699,N_6277,N_6396);
nor U6700 (N_6700,N_6435,N_6401);
or U6701 (N_6701,N_6295,N_6370);
xnor U6702 (N_6702,N_6449,N_6429);
nand U6703 (N_6703,N_6275,N_6489);
or U6704 (N_6704,N_6425,N_6319);
xor U6705 (N_6705,N_6305,N_6304);
nor U6706 (N_6706,N_6356,N_6348);
nor U6707 (N_6707,N_6360,N_6300);
nor U6708 (N_6708,N_6262,N_6304);
nand U6709 (N_6709,N_6319,N_6476);
or U6710 (N_6710,N_6462,N_6378);
xor U6711 (N_6711,N_6306,N_6302);
nor U6712 (N_6712,N_6493,N_6494);
or U6713 (N_6713,N_6432,N_6342);
or U6714 (N_6714,N_6334,N_6357);
or U6715 (N_6715,N_6412,N_6253);
xnor U6716 (N_6716,N_6269,N_6306);
or U6717 (N_6717,N_6276,N_6401);
nor U6718 (N_6718,N_6256,N_6401);
or U6719 (N_6719,N_6366,N_6443);
and U6720 (N_6720,N_6438,N_6292);
nor U6721 (N_6721,N_6290,N_6488);
xor U6722 (N_6722,N_6325,N_6312);
or U6723 (N_6723,N_6326,N_6254);
xnor U6724 (N_6724,N_6399,N_6330);
or U6725 (N_6725,N_6460,N_6328);
and U6726 (N_6726,N_6272,N_6258);
nand U6727 (N_6727,N_6347,N_6324);
xor U6728 (N_6728,N_6409,N_6270);
and U6729 (N_6729,N_6452,N_6409);
nand U6730 (N_6730,N_6339,N_6380);
xor U6731 (N_6731,N_6325,N_6475);
xnor U6732 (N_6732,N_6275,N_6253);
nand U6733 (N_6733,N_6425,N_6265);
xnor U6734 (N_6734,N_6312,N_6283);
or U6735 (N_6735,N_6324,N_6371);
and U6736 (N_6736,N_6415,N_6375);
and U6737 (N_6737,N_6358,N_6336);
and U6738 (N_6738,N_6424,N_6332);
nor U6739 (N_6739,N_6432,N_6329);
nand U6740 (N_6740,N_6491,N_6355);
xor U6741 (N_6741,N_6356,N_6338);
and U6742 (N_6742,N_6339,N_6315);
nand U6743 (N_6743,N_6445,N_6392);
nand U6744 (N_6744,N_6337,N_6408);
or U6745 (N_6745,N_6372,N_6430);
or U6746 (N_6746,N_6308,N_6264);
and U6747 (N_6747,N_6480,N_6334);
or U6748 (N_6748,N_6468,N_6397);
nand U6749 (N_6749,N_6253,N_6487);
and U6750 (N_6750,N_6593,N_6693);
xnor U6751 (N_6751,N_6543,N_6579);
and U6752 (N_6752,N_6659,N_6747);
and U6753 (N_6753,N_6565,N_6596);
and U6754 (N_6754,N_6511,N_6712);
nor U6755 (N_6755,N_6550,N_6518);
and U6756 (N_6756,N_6594,N_6674);
xor U6757 (N_6757,N_6698,N_6616);
or U6758 (N_6758,N_6651,N_6525);
nor U6759 (N_6759,N_6542,N_6634);
or U6760 (N_6760,N_6691,N_6728);
xnor U6761 (N_6761,N_6605,N_6715);
xnor U6762 (N_6762,N_6602,N_6512);
and U6763 (N_6763,N_6576,N_6531);
or U6764 (N_6764,N_6636,N_6666);
and U6765 (N_6765,N_6647,N_6718);
nor U6766 (N_6766,N_6574,N_6668);
and U6767 (N_6767,N_6702,N_6696);
and U6768 (N_6768,N_6617,N_6721);
xor U6769 (N_6769,N_6713,N_6716);
xnor U6770 (N_6770,N_6645,N_6708);
xor U6771 (N_6771,N_6719,N_6506);
nand U6772 (N_6772,N_6569,N_6629);
nor U6773 (N_6773,N_6709,N_6606);
xor U6774 (N_6774,N_6673,N_6717);
xnor U6775 (N_6775,N_6692,N_6662);
or U6776 (N_6776,N_6678,N_6580);
or U6777 (N_6777,N_6515,N_6612);
nand U6778 (N_6778,N_6639,N_6735);
or U6779 (N_6779,N_6567,N_6526);
xnor U6780 (N_6780,N_6738,N_6746);
xnor U6781 (N_6781,N_6592,N_6701);
or U6782 (N_6782,N_6649,N_6503);
xor U6783 (N_6783,N_6581,N_6749);
nor U6784 (N_6784,N_6578,N_6736);
nor U6785 (N_6785,N_6615,N_6614);
or U6786 (N_6786,N_6502,N_6588);
xnor U6787 (N_6787,N_6732,N_6711);
nand U6788 (N_6788,N_6589,N_6663);
nor U6789 (N_6789,N_6740,N_6539);
and U6790 (N_6790,N_6532,N_6670);
xor U6791 (N_6791,N_6573,N_6563);
xor U6792 (N_6792,N_6650,N_6582);
xor U6793 (N_6793,N_6695,N_6655);
and U6794 (N_6794,N_6609,N_6611);
nand U6795 (N_6795,N_6600,N_6687);
nand U6796 (N_6796,N_6646,N_6680);
xnor U6797 (N_6797,N_6590,N_6720);
nor U6798 (N_6798,N_6724,N_6560);
or U6799 (N_6799,N_6704,N_6552);
xor U6800 (N_6800,N_6585,N_6599);
nand U6801 (N_6801,N_6684,N_6640);
nor U6802 (N_6802,N_6501,N_6509);
nand U6803 (N_6803,N_6648,N_6570);
nor U6804 (N_6804,N_6672,N_6683);
and U6805 (N_6805,N_6730,N_6627);
xnor U6806 (N_6806,N_6628,N_6558);
xnor U6807 (N_6807,N_6729,N_6726);
and U6808 (N_6808,N_6598,N_6507);
nand U6809 (N_6809,N_6556,N_6528);
nand U6810 (N_6810,N_6633,N_6621);
nor U6811 (N_6811,N_6530,N_6522);
or U6812 (N_6812,N_6562,N_6685);
and U6813 (N_6813,N_6748,N_6632);
xnor U6814 (N_6814,N_6660,N_6745);
nand U6815 (N_6815,N_6638,N_6608);
and U6816 (N_6816,N_6519,N_6737);
or U6817 (N_6817,N_6547,N_6658);
or U6818 (N_6818,N_6675,N_6669);
or U6819 (N_6819,N_6641,N_6535);
nand U6820 (N_6820,N_6623,N_6686);
nor U6821 (N_6821,N_6619,N_6557);
nor U6822 (N_6822,N_6723,N_6707);
nor U6823 (N_6823,N_6591,N_6546);
and U6824 (N_6824,N_6739,N_6554);
xnor U6825 (N_6825,N_6653,N_6555);
and U6826 (N_6826,N_6700,N_6742);
and U6827 (N_6827,N_6635,N_6610);
or U6828 (N_6828,N_6601,N_6607);
nor U6829 (N_6829,N_6652,N_6553);
nand U6830 (N_6830,N_6731,N_6677);
xor U6831 (N_6831,N_6620,N_6624);
nor U6832 (N_6832,N_6604,N_6706);
and U6833 (N_6833,N_6699,N_6521);
nor U6834 (N_6834,N_6710,N_6540);
nand U6835 (N_6835,N_6741,N_6622);
nand U6836 (N_6836,N_6637,N_6688);
nand U6837 (N_6837,N_6527,N_6541);
and U6838 (N_6838,N_6597,N_6679);
nor U6839 (N_6839,N_6642,N_6661);
nand U6840 (N_6840,N_6537,N_6545);
and U6841 (N_6841,N_6544,N_6743);
or U6842 (N_6842,N_6566,N_6603);
nor U6843 (N_6843,N_6523,N_6689);
xor U6844 (N_6844,N_6690,N_6705);
or U6845 (N_6845,N_6551,N_6534);
and U6846 (N_6846,N_6734,N_6571);
or U6847 (N_6847,N_6657,N_6618);
xor U6848 (N_6848,N_6664,N_6714);
nand U6849 (N_6849,N_6722,N_6514);
or U6850 (N_6850,N_6725,N_6529);
xor U6851 (N_6851,N_6548,N_6665);
or U6852 (N_6852,N_6694,N_6671);
nor U6853 (N_6853,N_6744,N_6549);
nor U6854 (N_6854,N_6500,N_6625);
nand U6855 (N_6855,N_6654,N_6533);
nand U6856 (N_6856,N_6667,N_6626);
nand U6857 (N_6857,N_6656,N_6733);
nand U6858 (N_6858,N_6676,N_6587);
or U6859 (N_6859,N_6697,N_6630);
nand U6860 (N_6860,N_6524,N_6564);
or U6861 (N_6861,N_6510,N_6572);
and U6862 (N_6862,N_6727,N_6538);
or U6863 (N_6863,N_6631,N_6577);
nor U6864 (N_6864,N_6682,N_6536);
xor U6865 (N_6865,N_6584,N_6681);
or U6866 (N_6866,N_6586,N_6513);
or U6867 (N_6867,N_6517,N_6559);
and U6868 (N_6868,N_6643,N_6568);
nor U6869 (N_6869,N_6583,N_6644);
and U6870 (N_6870,N_6520,N_6504);
xor U6871 (N_6871,N_6561,N_6575);
or U6872 (N_6872,N_6508,N_6703);
nor U6873 (N_6873,N_6595,N_6505);
nand U6874 (N_6874,N_6516,N_6613);
nand U6875 (N_6875,N_6542,N_6545);
xor U6876 (N_6876,N_6598,N_6673);
or U6877 (N_6877,N_6687,N_6663);
or U6878 (N_6878,N_6614,N_6506);
nand U6879 (N_6879,N_6695,N_6505);
and U6880 (N_6880,N_6707,N_6506);
and U6881 (N_6881,N_6673,N_6728);
nor U6882 (N_6882,N_6599,N_6718);
nand U6883 (N_6883,N_6534,N_6688);
nor U6884 (N_6884,N_6557,N_6710);
xnor U6885 (N_6885,N_6684,N_6529);
and U6886 (N_6886,N_6551,N_6597);
xor U6887 (N_6887,N_6623,N_6502);
nand U6888 (N_6888,N_6670,N_6604);
nand U6889 (N_6889,N_6688,N_6570);
and U6890 (N_6890,N_6720,N_6608);
nand U6891 (N_6891,N_6628,N_6568);
and U6892 (N_6892,N_6584,N_6724);
nor U6893 (N_6893,N_6640,N_6507);
nor U6894 (N_6894,N_6560,N_6641);
nand U6895 (N_6895,N_6686,N_6512);
xnor U6896 (N_6896,N_6723,N_6546);
nor U6897 (N_6897,N_6729,N_6707);
and U6898 (N_6898,N_6619,N_6715);
or U6899 (N_6899,N_6685,N_6620);
nor U6900 (N_6900,N_6618,N_6519);
xor U6901 (N_6901,N_6708,N_6531);
xnor U6902 (N_6902,N_6632,N_6527);
and U6903 (N_6903,N_6679,N_6502);
nor U6904 (N_6904,N_6519,N_6735);
nor U6905 (N_6905,N_6674,N_6734);
nand U6906 (N_6906,N_6697,N_6511);
or U6907 (N_6907,N_6538,N_6500);
xnor U6908 (N_6908,N_6528,N_6548);
nand U6909 (N_6909,N_6589,N_6669);
and U6910 (N_6910,N_6699,N_6643);
or U6911 (N_6911,N_6742,N_6683);
nand U6912 (N_6912,N_6631,N_6694);
or U6913 (N_6913,N_6693,N_6542);
nor U6914 (N_6914,N_6526,N_6736);
nand U6915 (N_6915,N_6718,N_6531);
xor U6916 (N_6916,N_6646,N_6725);
or U6917 (N_6917,N_6589,N_6654);
or U6918 (N_6918,N_6673,N_6721);
xnor U6919 (N_6919,N_6679,N_6503);
xor U6920 (N_6920,N_6606,N_6695);
xor U6921 (N_6921,N_6554,N_6714);
and U6922 (N_6922,N_6534,N_6651);
xor U6923 (N_6923,N_6573,N_6507);
nor U6924 (N_6924,N_6734,N_6687);
nand U6925 (N_6925,N_6738,N_6589);
nand U6926 (N_6926,N_6599,N_6614);
nor U6927 (N_6927,N_6578,N_6608);
and U6928 (N_6928,N_6729,N_6737);
nand U6929 (N_6929,N_6691,N_6550);
and U6930 (N_6930,N_6736,N_6523);
and U6931 (N_6931,N_6741,N_6675);
or U6932 (N_6932,N_6657,N_6583);
or U6933 (N_6933,N_6559,N_6700);
xnor U6934 (N_6934,N_6634,N_6698);
nor U6935 (N_6935,N_6646,N_6536);
and U6936 (N_6936,N_6530,N_6598);
or U6937 (N_6937,N_6695,N_6568);
or U6938 (N_6938,N_6558,N_6570);
xnor U6939 (N_6939,N_6691,N_6651);
and U6940 (N_6940,N_6692,N_6608);
nor U6941 (N_6941,N_6615,N_6625);
nand U6942 (N_6942,N_6554,N_6579);
nand U6943 (N_6943,N_6742,N_6662);
nor U6944 (N_6944,N_6508,N_6707);
nand U6945 (N_6945,N_6594,N_6676);
nand U6946 (N_6946,N_6524,N_6556);
nor U6947 (N_6947,N_6613,N_6702);
or U6948 (N_6948,N_6724,N_6602);
nand U6949 (N_6949,N_6716,N_6673);
or U6950 (N_6950,N_6529,N_6514);
and U6951 (N_6951,N_6680,N_6707);
nand U6952 (N_6952,N_6674,N_6618);
and U6953 (N_6953,N_6559,N_6614);
or U6954 (N_6954,N_6640,N_6741);
or U6955 (N_6955,N_6527,N_6579);
or U6956 (N_6956,N_6718,N_6536);
or U6957 (N_6957,N_6677,N_6556);
nand U6958 (N_6958,N_6726,N_6714);
and U6959 (N_6959,N_6587,N_6714);
or U6960 (N_6960,N_6582,N_6567);
nor U6961 (N_6961,N_6520,N_6527);
xor U6962 (N_6962,N_6668,N_6634);
and U6963 (N_6963,N_6565,N_6609);
nand U6964 (N_6964,N_6555,N_6722);
or U6965 (N_6965,N_6616,N_6510);
nand U6966 (N_6966,N_6626,N_6582);
xnor U6967 (N_6967,N_6715,N_6508);
xnor U6968 (N_6968,N_6652,N_6732);
nor U6969 (N_6969,N_6529,N_6574);
nor U6970 (N_6970,N_6520,N_6559);
nand U6971 (N_6971,N_6669,N_6727);
or U6972 (N_6972,N_6627,N_6621);
nand U6973 (N_6973,N_6722,N_6613);
nor U6974 (N_6974,N_6524,N_6555);
xor U6975 (N_6975,N_6585,N_6744);
or U6976 (N_6976,N_6733,N_6727);
nand U6977 (N_6977,N_6634,N_6525);
nor U6978 (N_6978,N_6684,N_6678);
xnor U6979 (N_6979,N_6537,N_6530);
nand U6980 (N_6980,N_6554,N_6537);
or U6981 (N_6981,N_6688,N_6645);
xnor U6982 (N_6982,N_6547,N_6529);
xnor U6983 (N_6983,N_6684,N_6722);
and U6984 (N_6984,N_6685,N_6606);
nor U6985 (N_6985,N_6749,N_6500);
nor U6986 (N_6986,N_6525,N_6561);
or U6987 (N_6987,N_6693,N_6615);
and U6988 (N_6988,N_6693,N_6523);
or U6989 (N_6989,N_6623,N_6708);
nor U6990 (N_6990,N_6596,N_6560);
or U6991 (N_6991,N_6524,N_6687);
or U6992 (N_6992,N_6524,N_6720);
nor U6993 (N_6993,N_6626,N_6705);
nand U6994 (N_6994,N_6541,N_6701);
nor U6995 (N_6995,N_6607,N_6585);
xnor U6996 (N_6996,N_6582,N_6608);
nor U6997 (N_6997,N_6575,N_6626);
and U6998 (N_6998,N_6703,N_6526);
nor U6999 (N_6999,N_6666,N_6566);
xnor U7000 (N_7000,N_6845,N_6832);
nand U7001 (N_7001,N_6991,N_6978);
or U7002 (N_7002,N_6848,N_6955);
nor U7003 (N_7003,N_6807,N_6916);
nor U7004 (N_7004,N_6925,N_6990);
xor U7005 (N_7005,N_6939,N_6843);
and U7006 (N_7006,N_6881,N_6893);
nand U7007 (N_7007,N_6970,N_6971);
or U7008 (N_7008,N_6915,N_6953);
and U7009 (N_7009,N_6918,N_6873);
nand U7010 (N_7010,N_6750,N_6894);
or U7011 (N_7011,N_6917,N_6757);
xor U7012 (N_7012,N_6865,N_6907);
and U7013 (N_7013,N_6968,N_6982);
nand U7014 (N_7014,N_6803,N_6836);
and U7015 (N_7015,N_6884,N_6853);
and U7016 (N_7016,N_6801,N_6919);
xnor U7017 (N_7017,N_6872,N_6776);
and U7018 (N_7018,N_6805,N_6863);
and U7019 (N_7019,N_6870,N_6995);
xor U7020 (N_7020,N_6963,N_6756);
xor U7021 (N_7021,N_6794,N_6828);
or U7022 (N_7022,N_6935,N_6902);
xor U7023 (N_7023,N_6986,N_6823);
and U7024 (N_7024,N_6886,N_6849);
or U7025 (N_7025,N_6979,N_6974);
nor U7026 (N_7026,N_6854,N_6842);
and U7027 (N_7027,N_6763,N_6834);
and U7028 (N_7028,N_6829,N_6969);
and U7029 (N_7029,N_6835,N_6856);
and U7030 (N_7030,N_6754,N_6795);
and U7031 (N_7031,N_6879,N_6771);
and U7032 (N_7032,N_6851,N_6952);
or U7033 (N_7033,N_6777,N_6793);
xor U7034 (N_7034,N_6764,N_6784);
nor U7035 (N_7035,N_6831,N_6948);
nand U7036 (N_7036,N_6781,N_6958);
and U7037 (N_7037,N_6812,N_6800);
nand U7038 (N_7038,N_6837,N_6909);
nor U7039 (N_7039,N_6810,N_6941);
nor U7040 (N_7040,N_6906,N_6956);
or U7041 (N_7041,N_6871,N_6821);
and U7042 (N_7042,N_6840,N_6896);
nand U7043 (N_7043,N_6804,N_6944);
nand U7044 (N_7044,N_6892,N_6921);
and U7045 (N_7045,N_6996,N_6949);
nor U7046 (N_7046,N_6799,N_6911);
or U7047 (N_7047,N_6838,N_6857);
or U7048 (N_7048,N_6796,N_6772);
nor U7049 (N_7049,N_6993,N_6768);
nand U7050 (N_7050,N_6761,N_6975);
nor U7051 (N_7051,N_6850,N_6816);
nor U7052 (N_7052,N_6903,N_6876);
and U7053 (N_7053,N_6959,N_6759);
nand U7054 (N_7054,N_6976,N_6938);
and U7055 (N_7055,N_6887,N_6822);
nand U7056 (N_7056,N_6890,N_6895);
nand U7057 (N_7057,N_6862,N_6913);
xnor U7058 (N_7058,N_6806,N_6847);
or U7059 (N_7059,N_6880,N_6813);
or U7060 (N_7060,N_6904,N_6932);
nor U7061 (N_7061,N_6785,N_6942);
nor U7062 (N_7062,N_6770,N_6830);
nor U7063 (N_7063,N_6965,N_6927);
nand U7064 (N_7064,N_6751,N_6769);
xnor U7065 (N_7065,N_6888,N_6923);
or U7066 (N_7066,N_6758,N_6877);
or U7067 (N_7067,N_6934,N_6966);
nor U7068 (N_7068,N_6852,N_6885);
xor U7069 (N_7069,N_6767,N_6824);
xnor U7070 (N_7070,N_6814,N_6826);
nand U7071 (N_7071,N_6914,N_6954);
nor U7072 (N_7072,N_6908,N_6753);
and U7073 (N_7073,N_6878,N_6928);
xor U7074 (N_7074,N_6827,N_6985);
nor U7075 (N_7075,N_6773,N_6868);
nand U7076 (N_7076,N_6957,N_6988);
or U7077 (N_7077,N_6861,N_6855);
xor U7078 (N_7078,N_6946,N_6980);
and U7079 (N_7079,N_6936,N_6792);
nor U7080 (N_7080,N_6866,N_6931);
or U7081 (N_7081,N_6839,N_6947);
or U7082 (N_7082,N_6820,N_6858);
nor U7083 (N_7083,N_6790,N_6897);
xor U7084 (N_7084,N_6818,N_6950);
and U7085 (N_7085,N_6867,N_6984);
nor U7086 (N_7086,N_6844,N_6994);
nor U7087 (N_7087,N_6798,N_6926);
and U7088 (N_7088,N_6869,N_6983);
or U7089 (N_7089,N_6815,N_6766);
nand U7090 (N_7090,N_6780,N_6752);
or U7091 (N_7091,N_6951,N_6783);
nand U7092 (N_7092,N_6841,N_6762);
and U7093 (N_7093,N_6981,N_6987);
or U7094 (N_7094,N_6802,N_6977);
xnor U7095 (N_7095,N_6960,N_6972);
and U7096 (N_7096,N_6874,N_6898);
or U7097 (N_7097,N_6791,N_6901);
or U7098 (N_7098,N_6775,N_6962);
xnor U7099 (N_7099,N_6833,N_6809);
nor U7100 (N_7100,N_6900,N_6961);
and U7101 (N_7101,N_6786,N_6899);
or U7102 (N_7102,N_6864,N_6910);
or U7103 (N_7103,N_6787,N_6825);
nand U7104 (N_7104,N_6933,N_6967);
xnor U7105 (N_7105,N_6782,N_6859);
or U7106 (N_7106,N_6883,N_6905);
or U7107 (N_7107,N_6797,N_6891);
nand U7108 (N_7108,N_6929,N_6973);
nand U7109 (N_7109,N_6779,N_6964);
nor U7110 (N_7110,N_6889,N_6819);
xnor U7111 (N_7111,N_6760,N_6937);
nand U7112 (N_7112,N_6989,N_6924);
or U7113 (N_7113,N_6940,N_6808);
nand U7114 (N_7114,N_6774,N_6778);
and U7115 (N_7115,N_6999,N_6930);
or U7116 (N_7116,N_6998,N_6922);
or U7117 (N_7117,N_6860,N_6992);
nor U7118 (N_7118,N_6882,N_6755);
and U7119 (N_7119,N_6945,N_6789);
nand U7120 (N_7120,N_6997,N_6846);
or U7121 (N_7121,N_6912,N_6943);
and U7122 (N_7122,N_6788,N_6920);
nor U7123 (N_7123,N_6875,N_6811);
and U7124 (N_7124,N_6765,N_6817);
xnor U7125 (N_7125,N_6920,N_6877);
nand U7126 (N_7126,N_6995,N_6970);
and U7127 (N_7127,N_6849,N_6774);
or U7128 (N_7128,N_6956,N_6877);
xor U7129 (N_7129,N_6860,N_6753);
and U7130 (N_7130,N_6800,N_6955);
or U7131 (N_7131,N_6750,N_6816);
or U7132 (N_7132,N_6785,N_6972);
xnor U7133 (N_7133,N_6894,N_6988);
xor U7134 (N_7134,N_6933,N_6872);
or U7135 (N_7135,N_6764,N_6896);
nor U7136 (N_7136,N_6841,N_6940);
or U7137 (N_7137,N_6956,N_6939);
nand U7138 (N_7138,N_6804,N_6937);
and U7139 (N_7139,N_6889,N_6845);
or U7140 (N_7140,N_6964,N_6772);
nand U7141 (N_7141,N_6992,N_6789);
and U7142 (N_7142,N_6924,N_6829);
and U7143 (N_7143,N_6924,N_6785);
nor U7144 (N_7144,N_6931,N_6954);
nand U7145 (N_7145,N_6976,N_6842);
or U7146 (N_7146,N_6761,N_6823);
and U7147 (N_7147,N_6896,N_6794);
nor U7148 (N_7148,N_6877,N_6897);
and U7149 (N_7149,N_6777,N_6969);
or U7150 (N_7150,N_6774,N_6856);
nor U7151 (N_7151,N_6836,N_6787);
and U7152 (N_7152,N_6988,N_6763);
and U7153 (N_7153,N_6842,N_6999);
or U7154 (N_7154,N_6991,N_6976);
nand U7155 (N_7155,N_6854,N_6961);
or U7156 (N_7156,N_6790,N_6889);
xnor U7157 (N_7157,N_6897,N_6951);
nor U7158 (N_7158,N_6778,N_6958);
or U7159 (N_7159,N_6760,N_6837);
nor U7160 (N_7160,N_6855,N_6876);
nor U7161 (N_7161,N_6778,N_6768);
nand U7162 (N_7162,N_6883,N_6752);
xnor U7163 (N_7163,N_6833,N_6860);
nand U7164 (N_7164,N_6818,N_6843);
or U7165 (N_7165,N_6783,N_6912);
or U7166 (N_7166,N_6876,N_6895);
xnor U7167 (N_7167,N_6798,N_6818);
or U7168 (N_7168,N_6904,N_6859);
and U7169 (N_7169,N_6826,N_6848);
xor U7170 (N_7170,N_6886,N_6880);
xnor U7171 (N_7171,N_6895,N_6990);
nor U7172 (N_7172,N_6973,N_6907);
nor U7173 (N_7173,N_6808,N_6775);
and U7174 (N_7174,N_6957,N_6965);
or U7175 (N_7175,N_6762,N_6912);
nor U7176 (N_7176,N_6770,N_6852);
nor U7177 (N_7177,N_6892,N_6805);
nand U7178 (N_7178,N_6892,N_6934);
or U7179 (N_7179,N_6866,N_6904);
xor U7180 (N_7180,N_6783,N_6892);
nor U7181 (N_7181,N_6925,N_6839);
nor U7182 (N_7182,N_6920,N_6870);
or U7183 (N_7183,N_6796,N_6803);
and U7184 (N_7184,N_6836,N_6924);
nand U7185 (N_7185,N_6769,N_6827);
and U7186 (N_7186,N_6835,N_6911);
and U7187 (N_7187,N_6798,N_6929);
nand U7188 (N_7188,N_6870,N_6768);
xnor U7189 (N_7189,N_6933,N_6880);
nand U7190 (N_7190,N_6909,N_6997);
nor U7191 (N_7191,N_6930,N_6964);
and U7192 (N_7192,N_6978,N_6810);
or U7193 (N_7193,N_6956,N_6871);
or U7194 (N_7194,N_6767,N_6860);
nand U7195 (N_7195,N_6995,N_6865);
xnor U7196 (N_7196,N_6785,N_6879);
or U7197 (N_7197,N_6758,N_6822);
xor U7198 (N_7198,N_6854,N_6987);
and U7199 (N_7199,N_6760,N_6947);
nand U7200 (N_7200,N_6781,N_6873);
nand U7201 (N_7201,N_6902,N_6982);
nand U7202 (N_7202,N_6933,N_6766);
and U7203 (N_7203,N_6871,N_6750);
nand U7204 (N_7204,N_6972,N_6833);
nor U7205 (N_7205,N_6873,N_6877);
nand U7206 (N_7206,N_6968,N_6753);
xor U7207 (N_7207,N_6848,N_6908);
and U7208 (N_7208,N_6800,N_6934);
or U7209 (N_7209,N_6932,N_6883);
nand U7210 (N_7210,N_6987,N_6767);
xnor U7211 (N_7211,N_6772,N_6775);
and U7212 (N_7212,N_6917,N_6909);
nand U7213 (N_7213,N_6978,N_6844);
nor U7214 (N_7214,N_6941,N_6789);
or U7215 (N_7215,N_6765,N_6796);
or U7216 (N_7216,N_6945,N_6795);
nor U7217 (N_7217,N_6854,N_6979);
and U7218 (N_7218,N_6990,N_6832);
nand U7219 (N_7219,N_6844,N_6842);
or U7220 (N_7220,N_6966,N_6919);
nor U7221 (N_7221,N_6819,N_6962);
nor U7222 (N_7222,N_6935,N_6792);
nand U7223 (N_7223,N_6927,N_6964);
or U7224 (N_7224,N_6767,N_6966);
and U7225 (N_7225,N_6944,N_6795);
nor U7226 (N_7226,N_6980,N_6782);
or U7227 (N_7227,N_6788,N_6951);
xnor U7228 (N_7228,N_6873,N_6795);
xnor U7229 (N_7229,N_6760,N_6889);
or U7230 (N_7230,N_6846,N_6871);
nor U7231 (N_7231,N_6752,N_6948);
nor U7232 (N_7232,N_6752,N_6921);
nor U7233 (N_7233,N_6964,N_6807);
and U7234 (N_7234,N_6936,N_6766);
or U7235 (N_7235,N_6827,N_6779);
nor U7236 (N_7236,N_6961,N_6893);
or U7237 (N_7237,N_6852,N_6984);
nor U7238 (N_7238,N_6821,N_6927);
nand U7239 (N_7239,N_6981,N_6971);
nor U7240 (N_7240,N_6974,N_6775);
and U7241 (N_7241,N_6988,N_6978);
nand U7242 (N_7242,N_6914,N_6865);
nand U7243 (N_7243,N_6802,N_6823);
xnor U7244 (N_7244,N_6764,N_6972);
xor U7245 (N_7245,N_6806,N_6919);
and U7246 (N_7246,N_6818,N_6809);
xnor U7247 (N_7247,N_6979,N_6990);
xor U7248 (N_7248,N_6750,N_6930);
and U7249 (N_7249,N_6828,N_6965);
or U7250 (N_7250,N_7048,N_7199);
nand U7251 (N_7251,N_7124,N_7022);
nor U7252 (N_7252,N_7079,N_7036);
xor U7253 (N_7253,N_7189,N_7192);
nand U7254 (N_7254,N_7059,N_7066);
xnor U7255 (N_7255,N_7216,N_7068);
and U7256 (N_7256,N_7032,N_7152);
and U7257 (N_7257,N_7226,N_7146);
nor U7258 (N_7258,N_7098,N_7134);
or U7259 (N_7259,N_7183,N_7221);
nand U7260 (N_7260,N_7116,N_7111);
nand U7261 (N_7261,N_7043,N_7172);
xor U7262 (N_7262,N_7013,N_7207);
nand U7263 (N_7263,N_7218,N_7180);
or U7264 (N_7264,N_7144,N_7074);
and U7265 (N_7265,N_7108,N_7246);
nand U7266 (N_7266,N_7039,N_7009);
xor U7267 (N_7267,N_7031,N_7075);
and U7268 (N_7268,N_7064,N_7001);
and U7269 (N_7269,N_7167,N_7018);
and U7270 (N_7270,N_7087,N_7030);
and U7271 (N_7271,N_7238,N_7085);
or U7272 (N_7272,N_7091,N_7149);
nor U7273 (N_7273,N_7093,N_7140);
or U7274 (N_7274,N_7073,N_7110);
nand U7275 (N_7275,N_7159,N_7233);
nand U7276 (N_7276,N_7200,N_7065);
nor U7277 (N_7277,N_7240,N_7109);
or U7278 (N_7278,N_7229,N_7025);
or U7279 (N_7279,N_7176,N_7129);
and U7280 (N_7280,N_7014,N_7042);
xnor U7281 (N_7281,N_7128,N_7212);
nor U7282 (N_7282,N_7104,N_7205);
nor U7283 (N_7283,N_7024,N_7041);
nor U7284 (N_7284,N_7148,N_7099);
nor U7285 (N_7285,N_7121,N_7114);
xnor U7286 (N_7286,N_7203,N_7228);
nand U7287 (N_7287,N_7217,N_7070);
nor U7288 (N_7288,N_7100,N_7188);
nor U7289 (N_7289,N_7053,N_7056);
nand U7290 (N_7290,N_7225,N_7008);
or U7291 (N_7291,N_7224,N_7236);
xor U7292 (N_7292,N_7135,N_7165);
nor U7293 (N_7293,N_7050,N_7164);
nand U7294 (N_7294,N_7173,N_7137);
and U7295 (N_7295,N_7231,N_7220);
nand U7296 (N_7296,N_7047,N_7069);
xor U7297 (N_7297,N_7011,N_7143);
or U7298 (N_7298,N_7150,N_7182);
nor U7299 (N_7299,N_7016,N_7208);
nand U7300 (N_7300,N_7198,N_7211);
or U7301 (N_7301,N_7219,N_7177);
or U7302 (N_7302,N_7132,N_7045);
nand U7303 (N_7303,N_7082,N_7058);
nor U7304 (N_7304,N_7141,N_7103);
nor U7305 (N_7305,N_7202,N_7044);
or U7306 (N_7306,N_7102,N_7094);
nand U7307 (N_7307,N_7125,N_7184);
nor U7308 (N_7308,N_7088,N_7245);
and U7309 (N_7309,N_7197,N_7154);
or U7310 (N_7310,N_7239,N_7005);
nand U7311 (N_7311,N_7092,N_7247);
and U7312 (N_7312,N_7210,N_7115);
and U7313 (N_7313,N_7223,N_7248);
nor U7314 (N_7314,N_7190,N_7195);
or U7315 (N_7315,N_7118,N_7232);
nor U7316 (N_7316,N_7076,N_7027);
or U7317 (N_7317,N_7123,N_7168);
and U7318 (N_7318,N_7158,N_7117);
and U7319 (N_7319,N_7185,N_7107);
xnor U7320 (N_7320,N_7175,N_7193);
xnor U7321 (N_7321,N_7206,N_7153);
and U7322 (N_7322,N_7089,N_7051);
xnor U7323 (N_7323,N_7007,N_7170);
and U7324 (N_7324,N_7057,N_7105);
or U7325 (N_7325,N_7122,N_7215);
nor U7326 (N_7326,N_7162,N_7020);
or U7327 (N_7327,N_7004,N_7234);
xnor U7328 (N_7328,N_7080,N_7151);
nand U7329 (N_7329,N_7242,N_7213);
nand U7330 (N_7330,N_7244,N_7026);
or U7331 (N_7331,N_7230,N_7201);
and U7332 (N_7332,N_7133,N_7040);
or U7333 (N_7333,N_7037,N_7097);
xor U7334 (N_7334,N_7196,N_7034);
nand U7335 (N_7335,N_7010,N_7178);
nor U7336 (N_7336,N_7171,N_7084);
and U7337 (N_7337,N_7002,N_7077);
or U7338 (N_7338,N_7072,N_7157);
nand U7339 (N_7339,N_7033,N_7209);
xor U7340 (N_7340,N_7191,N_7046);
xor U7341 (N_7341,N_7187,N_7023);
nor U7342 (N_7342,N_7090,N_7081);
or U7343 (N_7343,N_7106,N_7155);
xnor U7344 (N_7344,N_7235,N_7028);
xor U7345 (N_7345,N_7126,N_7127);
and U7346 (N_7346,N_7038,N_7078);
or U7347 (N_7347,N_7054,N_7119);
nand U7348 (N_7348,N_7169,N_7156);
xnor U7349 (N_7349,N_7147,N_7035);
or U7350 (N_7350,N_7083,N_7136);
nand U7351 (N_7351,N_7071,N_7095);
nand U7352 (N_7352,N_7055,N_7179);
xnor U7353 (N_7353,N_7000,N_7241);
or U7354 (N_7354,N_7222,N_7142);
nor U7355 (N_7355,N_7130,N_7112);
and U7356 (N_7356,N_7249,N_7161);
xor U7357 (N_7357,N_7015,N_7194);
nand U7358 (N_7358,N_7139,N_7060);
xnor U7359 (N_7359,N_7243,N_7062);
nand U7360 (N_7360,N_7166,N_7186);
or U7361 (N_7361,N_7086,N_7029);
xnor U7362 (N_7362,N_7204,N_7174);
nor U7363 (N_7363,N_7138,N_7237);
nor U7364 (N_7364,N_7019,N_7163);
or U7365 (N_7365,N_7131,N_7006);
xnor U7366 (N_7366,N_7063,N_7120);
and U7367 (N_7367,N_7003,N_7181);
xor U7368 (N_7368,N_7145,N_7101);
nor U7369 (N_7369,N_7061,N_7160);
nand U7370 (N_7370,N_7096,N_7021);
and U7371 (N_7371,N_7227,N_7049);
xor U7372 (N_7372,N_7214,N_7067);
and U7373 (N_7373,N_7017,N_7052);
nand U7374 (N_7374,N_7012,N_7113);
and U7375 (N_7375,N_7008,N_7211);
nor U7376 (N_7376,N_7181,N_7182);
nand U7377 (N_7377,N_7039,N_7208);
and U7378 (N_7378,N_7033,N_7171);
nand U7379 (N_7379,N_7052,N_7200);
nand U7380 (N_7380,N_7178,N_7102);
or U7381 (N_7381,N_7143,N_7191);
nand U7382 (N_7382,N_7061,N_7032);
and U7383 (N_7383,N_7235,N_7157);
and U7384 (N_7384,N_7042,N_7180);
xnor U7385 (N_7385,N_7137,N_7177);
xnor U7386 (N_7386,N_7067,N_7164);
nand U7387 (N_7387,N_7095,N_7101);
or U7388 (N_7388,N_7231,N_7137);
nor U7389 (N_7389,N_7127,N_7230);
or U7390 (N_7390,N_7068,N_7243);
nand U7391 (N_7391,N_7048,N_7121);
nor U7392 (N_7392,N_7140,N_7202);
nor U7393 (N_7393,N_7200,N_7132);
or U7394 (N_7394,N_7002,N_7075);
and U7395 (N_7395,N_7140,N_7007);
nor U7396 (N_7396,N_7198,N_7027);
nor U7397 (N_7397,N_7065,N_7052);
nand U7398 (N_7398,N_7169,N_7249);
or U7399 (N_7399,N_7049,N_7120);
and U7400 (N_7400,N_7101,N_7226);
or U7401 (N_7401,N_7076,N_7216);
xor U7402 (N_7402,N_7204,N_7127);
xor U7403 (N_7403,N_7173,N_7005);
and U7404 (N_7404,N_7135,N_7203);
xnor U7405 (N_7405,N_7153,N_7125);
or U7406 (N_7406,N_7199,N_7109);
nand U7407 (N_7407,N_7080,N_7009);
nand U7408 (N_7408,N_7009,N_7036);
or U7409 (N_7409,N_7000,N_7185);
nor U7410 (N_7410,N_7046,N_7209);
or U7411 (N_7411,N_7247,N_7220);
xnor U7412 (N_7412,N_7234,N_7124);
xnor U7413 (N_7413,N_7149,N_7077);
nand U7414 (N_7414,N_7170,N_7235);
or U7415 (N_7415,N_7125,N_7162);
nor U7416 (N_7416,N_7233,N_7014);
and U7417 (N_7417,N_7053,N_7115);
nand U7418 (N_7418,N_7129,N_7011);
nand U7419 (N_7419,N_7239,N_7175);
and U7420 (N_7420,N_7025,N_7022);
nand U7421 (N_7421,N_7243,N_7233);
nand U7422 (N_7422,N_7176,N_7139);
or U7423 (N_7423,N_7094,N_7236);
nor U7424 (N_7424,N_7141,N_7206);
or U7425 (N_7425,N_7184,N_7136);
or U7426 (N_7426,N_7228,N_7219);
nor U7427 (N_7427,N_7131,N_7223);
or U7428 (N_7428,N_7005,N_7054);
nand U7429 (N_7429,N_7245,N_7091);
and U7430 (N_7430,N_7043,N_7001);
or U7431 (N_7431,N_7046,N_7240);
or U7432 (N_7432,N_7078,N_7014);
nand U7433 (N_7433,N_7127,N_7062);
nor U7434 (N_7434,N_7203,N_7176);
or U7435 (N_7435,N_7188,N_7010);
nor U7436 (N_7436,N_7028,N_7159);
and U7437 (N_7437,N_7022,N_7108);
nand U7438 (N_7438,N_7196,N_7190);
or U7439 (N_7439,N_7047,N_7010);
nor U7440 (N_7440,N_7235,N_7041);
and U7441 (N_7441,N_7021,N_7099);
and U7442 (N_7442,N_7134,N_7240);
xor U7443 (N_7443,N_7117,N_7193);
and U7444 (N_7444,N_7185,N_7023);
nor U7445 (N_7445,N_7175,N_7176);
xor U7446 (N_7446,N_7215,N_7110);
nand U7447 (N_7447,N_7073,N_7120);
and U7448 (N_7448,N_7173,N_7228);
nand U7449 (N_7449,N_7207,N_7015);
or U7450 (N_7450,N_7123,N_7239);
xor U7451 (N_7451,N_7080,N_7240);
or U7452 (N_7452,N_7136,N_7089);
nor U7453 (N_7453,N_7232,N_7048);
nand U7454 (N_7454,N_7214,N_7001);
or U7455 (N_7455,N_7040,N_7024);
nor U7456 (N_7456,N_7083,N_7114);
nand U7457 (N_7457,N_7029,N_7207);
and U7458 (N_7458,N_7039,N_7061);
xnor U7459 (N_7459,N_7135,N_7034);
xor U7460 (N_7460,N_7244,N_7136);
or U7461 (N_7461,N_7029,N_7122);
nor U7462 (N_7462,N_7168,N_7189);
nand U7463 (N_7463,N_7055,N_7241);
and U7464 (N_7464,N_7075,N_7052);
nor U7465 (N_7465,N_7112,N_7146);
nand U7466 (N_7466,N_7216,N_7247);
and U7467 (N_7467,N_7051,N_7210);
xor U7468 (N_7468,N_7015,N_7161);
xnor U7469 (N_7469,N_7154,N_7043);
or U7470 (N_7470,N_7120,N_7060);
nand U7471 (N_7471,N_7038,N_7221);
nand U7472 (N_7472,N_7232,N_7219);
and U7473 (N_7473,N_7063,N_7161);
nand U7474 (N_7474,N_7152,N_7147);
nand U7475 (N_7475,N_7061,N_7053);
or U7476 (N_7476,N_7232,N_7167);
and U7477 (N_7477,N_7084,N_7007);
or U7478 (N_7478,N_7097,N_7074);
xnor U7479 (N_7479,N_7132,N_7093);
nand U7480 (N_7480,N_7096,N_7036);
and U7481 (N_7481,N_7146,N_7006);
or U7482 (N_7482,N_7133,N_7093);
nand U7483 (N_7483,N_7194,N_7150);
or U7484 (N_7484,N_7210,N_7202);
or U7485 (N_7485,N_7107,N_7023);
nand U7486 (N_7486,N_7214,N_7000);
and U7487 (N_7487,N_7055,N_7142);
and U7488 (N_7488,N_7128,N_7244);
xor U7489 (N_7489,N_7080,N_7208);
and U7490 (N_7490,N_7246,N_7107);
xor U7491 (N_7491,N_7080,N_7105);
nor U7492 (N_7492,N_7177,N_7135);
nand U7493 (N_7493,N_7133,N_7105);
nor U7494 (N_7494,N_7221,N_7176);
nand U7495 (N_7495,N_7173,N_7219);
or U7496 (N_7496,N_7027,N_7151);
xor U7497 (N_7497,N_7228,N_7049);
or U7498 (N_7498,N_7136,N_7013);
xor U7499 (N_7499,N_7030,N_7080);
xnor U7500 (N_7500,N_7275,N_7421);
or U7501 (N_7501,N_7318,N_7471);
xnor U7502 (N_7502,N_7309,N_7356);
nor U7503 (N_7503,N_7448,N_7419);
nor U7504 (N_7504,N_7317,N_7447);
or U7505 (N_7505,N_7369,N_7461);
nand U7506 (N_7506,N_7385,N_7282);
nor U7507 (N_7507,N_7340,N_7303);
nand U7508 (N_7508,N_7284,N_7281);
nand U7509 (N_7509,N_7298,N_7494);
and U7510 (N_7510,N_7406,N_7417);
and U7511 (N_7511,N_7366,N_7405);
and U7512 (N_7512,N_7264,N_7364);
nor U7513 (N_7513,N_7467,N_7423);
nand U7514 (N_7514,N_7381,N_7386);
nor U7515 (N_7515,N_7465,N_7397);
and U7516 (N_7516,N_7491,N_7472);
xnor U7517 (N_7517,N_7258,N_7322);
nor U7518 (N_7518,N_7291,N_7443);
nor U7519 (N_7519,N_7262,N_7367);
or U7520 (N_7520,N_7348,N_7300);
xnor U7521 (N_7521,N_7251,N_7352);
nor U7522 (N_7522,N_7365,N_7402);
and U7523 (N_7523,N_7350,N_7452);
nand U7524 (N_7524,N_7445,N_7329);
and U7525 (N_7525,N_7325,N_7279);
and U7526 (N_7526,N_7328,N_7389);
nand U7527 (N_7527,N_7437,N_7408);
xnor U7528 (N_7528,N_7285,N_7411);
nand U7529 (N_7529,N_7260,N_7272);
nor U7530 (N_7530,N_7478,N_7439);
nand U7531 (N_7531,N_7430,N_7359);
nor U7532 (N_7532,N_7353,N_7254);
and U7533 (N_7533,N_7458,N_7480);
nand U7534 (N_7534,N_7259,N_7257);
xor U7535 (N_7535,N_7357,N_7349);
xnor U7536 (N_7536,N_7312,N_7400);
nand U7537 (N_7537,N_7473,N_7296);
nand U7538 (N_7538,N_7360,N_7487);
xnor U7539 (N_7539,N_7392,N_7307);
nor U7540 (N_7540,N_7354,N_7435);
and U7541 (N_7541,N_7370,N_7475);
and U7542 (N_7542,N_7394,N_7489);
nor U7543 (N_7543,N_7396,N_7306);
xor U7544 (N_7544,N_7433,N_7265);
and U7545 (N_7545,N_7483,N_7278);
nand U7546 (N_7546,N_7399,N_7401);
or U7547 (N_7547,N_7256,N_7498);
nand U7548 (N_7548,N_7302,N_7476);
and U7549 (N_7549,N_7334,N_7269);
and U7550 (N_7550,N_7431,N_7362);
nand U7551 (N_7551,N_7455,N_7299);
or U7552 (N_7552,N_7315,N_7422);
nor U7553 (N_7553,N_7323,N_7468);
and U7554 (N_7554,N_7355,N_7444);
or U7555 (N_7555,N_7384,N_7415);
nand U7556 (N_7556,N_7333,N_7407);
nand U7557 (N_7557,N_7286,N_7324);
nor U7558 (N_7558,N_7441,N_7288);
and U7559 (N_7559,N_7482,N_7289);
nor U7560 (N_7560,N_7297,N_7273);
and U7561 (N_7561,N_7363,N_7438);
nor U7562 (N_7562,N_7409,N_7398);
or U7563 (N_7563,N_7450,N_7492);
or U7564 (N_7564,N_7379,N_7280);
nand U7565 (N_7565,N_7342,N_7267);
nor U7566 (N_7566,N_7429,N_7294);
nand U7567 (N_7567,N_7375,N_7404);
xor U7568 (N_7568,N_7388,N_7368);
xnor U7569 (N_7569,N_7477,N_7341);
or U7570 (N_7570,N_7481,N_7464);
xnor U7571 (N_7571,N_7361,N_7283);
nor U7572 (N_7572,N_7451,N_7466);
xor U7573 (N_7573,N_7321,N_7330);
xor U7574 (N_7574,N_7446,N_7270);
nand U7575 (N_7575,N_7380,N_7486);
nor U7576 (N_7576,N_7474,N_7311);
nor U7577 (N_7577,N_7308,N_7484);
and U7578 (N_7578,N_7428,N_7319);
or U7579 (N_7579,N_7292,N_7449);
or U7580 (N_7580,N_7337,N_7346);
xor U7581 (N_7581,N_7343,N_7436);
or U7582 (N_7582,N_7347,N_7295);
nand U7583 (N_7583,N_7456,N_7331);
nor U7584 (N_7584,N_7310,N_7424);
nor U7585 (N_7585,N_7412,N_7326);
xor U7586 (N_7586,N_7304,N_7268);
nor U7587 (N_7587,N_7377,N_7293);
xnor U7588 (N_7588,N_7263,N_7387);
nor U7589 (N_7589,N_7344,N_7332);
nand U7590 (N_7590,N_7252,N_7493);
nand U7591 (N_7591,N_7414,N_7338);
and U7592 (N_7592,N_7434,N_7425);
nor U7593 (N_7593,N_7371,N_7479);
xor U7594 (N_7594,N_7305,N_7327);
xnor U7595 (N_7595,N_7314,N_7255);
or U7596 (N_7596,N_7490,N_7287);
and U7597 (N_7597,N_7393,N_7403);
xnor U7598 (N_7598,N_7442,N_7470);
nor U7599 (N_7599,N_7276,N_7460);
and U7600 (N_7600,N_7373,N_7410);
xor U7601 (N_7601,N_7358,N_7374);
nand U7602 (N_7602,N_7463,N_7301);
nor U7603 (N_7603,N_7336,N_7469);
nor U7604 (N_7604,N_7496,N_7457);
xnor U7605 (N_7605,N_7432,N_7376);
xor U7606 (N_7606,N_7420,N_7426);
and U7607 (N_7607,N_7271,N_7495);
nor U7608 (N_7608,N_7391,N_7413);
and U7609 (N_7609,N_7378,N_7382);
or U7610 (N_7610,N_7488,N_7497);
xnor U7611 (N_7611,N_7313,N_7454);
nor U7612 (N_7612,N_7253,N_7499);
xor U7613 (N_7613,N_7345,N_7316);
nand U7614 (N_7614,N_7277,N_7339);
and U7615 (N_7615,N_7290,N_7383);
xor U7616 (N_7616,N_7418,N_7335);
xor U7617 (N_7617,N_7351,N_7427);
nor U7618 (N_7618,N_7459,N_7485);
and U7619 (N_7619,N_7462,N_7416);
nand U7620 (N_7620,N_7395,N_7453);
xnor U7621 (N_7621,N_7390,N_7266);
xor U7622 (N_7622,N_7250,N_7440);
nor U7623 (N_7623,N_7320,N_7274);
nor U7624 (N_7624,N_7261,N_7372);
or U7625 (N_7625,N_7308,N_7372);
and U7626 (N_7626,N_7327,N_7310);
xnor U7627 (N_7627,N_7287,N_7400);
and U7628 (N_7628,N_7360,N_7319);
or U7629 (N_7629,N_7340,N_7260);
and U7630 (N_7630,N_7265,N_7360);
nand U7631 (N_7631,N_7262,N_7308);
and U7632 (N_7632,N_7263,N_7408);
or U7633 (N_7633,N_7318,N_7411);
nand U7634 (N_7634,N_7390,N_7289);
or U7635 (N_7635,N_7286,N_7426);
nand U7636 (N_7636,N_7267,N_7376);
xnor U7637 (N_7637,N_7332,N_7301);
nor U7638 (N_7638,N_7348,N_7386);
xor U7639 (N_7639,N_7291,N_7408);
nor U7640 (N_7640,N_7265,N_7473);
and U7641 (N_7641,N_7275,N_7440);
nand U7642 (N_7642,N_7305,N_7483);
nand U7643 (N_7643,N_7475,N_7310);
and U7644 (N_7644,N_7489,N_7260);
xnor U7645 (N_7645,N_7433,N_7275);
nand U7646 (N_7646,N_7491,N_7424);
nand U7647 (N_7647,N_7387,N_7302);
nor U7648 (N_7648,N_7372,N_7401);
and U7649 (N_7649,N_7442,N_7345);
nand U7650 (N_7650,N_7339,N_7390);
xnor U7651 (N_7651,N_7286,N_7277);
or U7652 (N_7652,N_7322,N_7391);
or U7653 (N_7653,N_7264,N_7381);
xor U7654 (N_7654,N_7268,N_7447);
nor U7655 (N_7655,N_7381,N_7277);
nand U7656 (N_7656,N_7409,N_7461);
nor U7657 (N_7657,N_7307,N_7484);
xor U7658 (N_7658,N_7272,N_7346);
or U7659 (N_7659,N_7374,N_7267);
xnor U7660 (N_7660,N_7406,N_7294);
nand U7661 (N_7661,N_7302,N_7288);
and U7662 (N_7662,N_7401,N_7313);
xnor U7663 (N_7663,N_7480,N_7451);
nor U7664 (N_7664,N_7340,N_7496);
nand U7665 (N_7665,N_7483,N_7306);
nand U7666 (N_7666,N_7460,N_7424);
nand U7667 (N_7667,N_7478,N_7414);
and U7668 (N_7668,N_7475,N_7446);
nor U7669 (N_7669,N_7447,N_7402);
and U7670 (N_7670,N_7355,N_7259);
and U7671 (N_7671,N_7274,N_7427);
nor U7672 (N_7672,N_7411,N_7457);
nand U7673 (N_7673,N_7493,N_7451);
and U7674 (N_7674,N_7474,N_7476);
nand U7675 (N_7675,N_7271,N_7288);
or U7676 (N_7676,N_7387,N_7343);
xor U7677 (N_7677,N_7393,N_7315);
nor U7678 (N_7678,N_7404,N_7368);
and U7679 (N_7679,N_7271,N_7356);
xnor U7680 (N_7680,N_7337,N_7265);
nor U7681 (N_7681,N_7488,N_7366);
xor U7682 (N_7682,N_7406,N_7480);
xnor U7683 (N_7683,N_7299,N_7268);
and U7684 (N_7684,N_7348,N_7313);
xnor U7685 (N_7685,N_7256,N_7334);
or U7686 (N_7686,N_7331,N_7327);
and U7687 (N_7687,N_7407,N_7457);
and U7688 (N_7688,N_7396,N_7376);
or U7689 (N_7689,N_7453,N_7318);
or U7690 (N_7690,N_7492,N_7302);
xor U7691 (N_7691,N_7434,N_7419);
and U7692 (N_7692,N_7260,N_7313);
and U7693 (N_7693,N_7492,N_7257);
and U7694 (N_7694,N_7363,N_7429);
and U7695 (N_7695,N_7389,N_7304);
or U7696 (N_7696,N_7441,N_7463);
nand U7697 (N_7697,N_7258,N_7430);
or U7698 (N_7698,N_7424,N_7329);
xnor U7699 (N_7699,N_7487,N_7251);
and U7700 (N_7700,N_7327,N_7490);
xor U7701 (N_7701,N_7271,N_7452);
nor U7702 (N_7702,N_7263,N_7405);
or U7703 (N_7703,N_7407,N_7494);
nor U7704 (N_7704,N_7319,N_7251);
and U7705 (N_7705,N_7379,N_7483);
xor U7706 (N_7706,N_7381,N_7461);
xnor U7707 (N_7707,N_7418,N_7433);
or U7708 (N_7708,N_7310,N_7402);
nor U7709 (N_7709,N_7293,N_7263);
nor U7710 (N_7710,N_7250,N_7260);
nand U7711 (N_7711,N_7490,N_7414);
nor U7712 (N_7712,N_7365,N_7261);
or U7713 (N_7713,N_7462,N_7472);
and U7714 (N_7714,N_7376,N_7472);
nand U7715 (N_7715,N_7487,N_7315);
xor U7716 (N_7716,N_7419,N_7483);
xnor U7717 (N_7717,N_7307,N_7285);
nand U7718 (N_7718,N_7378,N_7362);
and U7719 (N_7719,N_7360,N_7345);
nor U7720 (N_7720,N_7363,N_7277);
and U7721 (N_7721,N_7373,N_7254);
and U7722 (N_7722,N_7357,N_7385);
or U7723 (N_7723,N_7407,N_7307);
nand U7724 (N_7724,N_7458,N_7433);
nor U7725 (N_7725,N_7403,N_7443);
nor U7726 (N_7726,N_7272,N_7342);
nor U7727 (N_7727,N_7252,N_7311);
or U7728 (N_7728,N_7265,N_7427);
and U7729 (N_7729,N_7489,N_7480);
or U7730 (N_7730,N_7461,N_7336);
nor U7731 (N_7731,N_7370,N_7324);
xnor U7732 (N_7732,N_7424,N_7295);
xnor U7733 (N_7733,N_7339,N_7358);
or U7734 (N_7734,N_7357,N_7450);
xnor U7735 (N_7735,N_7305,N_7313);
nand U7736 (N_7736,N_7413,N_7308);
and U7737 (N_7737,N_7384,N_7323);
xnor U7738 (N_7738,N_7415,N_7282);
nor U7739 (N_7739,N_7337,N_7441);
and U7740 (N_7740,N_7342,N_7476);
or U7741 (N_7741,N_7395,N_7485);
and U7742 (N_7742,N_7287,N_7444);
nor U7743 (N_7743,N_7403,N_7468);
nand U7744 (N_7744,N_7421,N_7419);
nor U7745 (N_7745,N_7417,N_7329);
xnor U7746 (N_7746,N_7293,N_7360);
nand U7747 (N_7747,N_7339,N_7486);
or U7748 (N_7748,N_7397,N_7346);
xnor U7749 (N_7749,N_7476,N_7482);
and U7750 (N_7750,N_7616,N_7543);
nor U7751 (N_7751,N_7737,N_7548);
nor U7752 (N_7752,N_7563,N_7549);
nand U7753 (N_7753,N_7671,N_7514);
nand U7754 (N_7754,N_7683,N_7556);
nand U7755 (N_7755,N_7668,N_7732);
nor U7756 (N_7756,N_7555,N_7697);
or U7757 (N_7757,N_7526,N_7680);
xnor U7758 (N_7758,N_7505,N_7622);
xnor U7759 (N_7759,N_7714,N_7586);
or U7760 (N_7760,N_7702,N_7538);
nor U7761 (N_7761,N_7627,N_7749);
nor U7762 (N_7762,N_7710,N_7676);
nor U7763 (N_7763,N_7547,N_7695);
or U7764 (N_7764,N_7648,N_7582);
and U7765 (N_7765,N_7635,N_7643);
nor U7766 (N_7766,N_7621,N_7561);
nor U7767 (N_7767,N_7507,N_7504);
xor U7768 (N_7768,N_7532,N_7649);
xnor U7769 (N_7769,N_7735,N_7742);
nand U7770 (N_7770,N_7642,N_7607);
xor U7771 (N_7771,N_7740,N_7747);
xor U7772 (N_7772,N_7545,N_7730);
and U7773 (N_7773,N_7592,N_7550);
nor U7774 (N_7774,N_7728,N_7654);
nand U7775 (N_7775,N_7723,N_7738);
nand U7776 (N_7776,N_7693,N_7703);
xnor U7777 (N_7777,N_7587,N_7694);
nor U7778 (N_7778,N_7717,N_7523);
and U7779 (N_7779,N_7571,N_7589);
and U7780 (N_7780,N_7594,N_7533);
nor U7781 (N_7781,N_7713,N_7729);
nor U7782 (N_7782,N_7577,N_7708);
nor U7783 (N_7783,N_7591,N_7516);
and U7784 (N_7784,N_7739,N_7600);
nand U7785 (N_7785,N_7559,N_7660);
xnor U7786 (N_7786,N_7520,N_7701);
nand U7787 (N_7787,N_7630,N_7704);
or U7788 (N_7788,N_7678,N_7634);
nor U7789 (N_7789,N_7528,N_7527);
xnor U7790 (N_7790,N_7509,N_7593);
nor U7791 (N_7791,N_7576,N_7597);
xnor U7792 (N_7792,N_7652,N_7707);
nand U7793 (N_7793,N_7614,N_7746);
and U7794 (N_7794,N_7689,N_7610);
or U7795 (N_7795,N_7584,N_7684);
or U7796 (N_7796,N_7631,N_7640);
and U7797 (N_7797,N_7570,N_7688);
nor U7798 (N_7798,N_7724,N_7595);
or U7799 (N_7799,N_7691,N_7679);
nor U7800 (N_7800,N_7674,N_7588);
nand U7801 (N_7801,N_7639,N_7568);
or U7802 (N_7802,N_7733,N_7743);
and U7803 (N_7803,N_7657,N_7675);
or U7804 (N_7804,N_7522,N_7603);
nor U7805 (N_7805,N_7531,N_7551);
or U7806 (N_7806,N_7727,N_7651);
nand U7807 (N_7807,N_7655,N_7682);
and U7808 (N_7808,N_7517,N_7669);
or U7809 (N_7809,N_7530,N_7578);
xor U7810 (N_7810,N_7511,N_7557);
nand U7811 (N_7811,N_7629,N_7656);
and U7812 (N_7812,N_7672,N_7725);
or U7813 (N_7813,N_7513,N_7540);
nand U7814 (N_7814,N_7687,N_7662);
nor U7815 (N_7815,N_7506,N_7685);
nor U7816 (N_7816,N_7647,N_7501);
xor U7817 (N_7817,N_7529,N_7510);
and U7818 (N_7818,N_7598,N_7542);
nand U7819 (N_7819,N_7736,N_7663);
or U7820 (N_7820,N_7508,N_7638);
nand U7821 (N_7821,N_7601,N_7536);
and U7822 (N_7822,N_7625,N_7612);
nor U7823 (N_7823,N_7572,N_7661);
xor U7824 (N_7824,N_7515,N_7650);
xnor U7825 (N_7825,N_7623,N_7681);
and U7826 (N_7826,N_7718,N_7580);
nor U7827 (N_7827,N_7521,N_7604);
nand U7828 (N_7828,N_7562,N_7575);
nand U7829 (N_7829,N_7569,N_7664);
nor U7830 (N_7830,N_7565,N_7525);
xnor U7831 (N_7831,N_7537,N_7636);
and U7832 (N_7832,N_7573,N_7615);
or U7833 (N_7833,N_7644,N_7626);
and U7834 (N_7834,N_7566,N_7558);
nor U7835 (N_7835,N_7722,N_7609);
and U7836 (N_7836,N_7734,N_7641);
nand U7837 (N_7837,N_7605,N_7599);
xor U7838 (N_7838,N_7602,N_7744);
nand U7839 (N_7839,N_7706,N_7741);
nand U7840 (N_7840,N_7590,N_7709);
nor U7841 (N_7841,N_7686,N_7535);
and U7842 (N_7842,N_7618,N_7645);
or U7843 (N_7843,N_7711,N_7726);
nand U7844 (N_7844,N_7617,N_7628);
xnor U7845 (N_7845,N_7692,N_7715);
and U7846 (N_7846,N_7585,N_7519);
nor U7847 (N_7847,N_7611,N_7544);
nor U7848 (N_7848,N_7721,N_7698);
nand U7849 (N_7849,N_7564,N_7574);
nor U7850 (N_7850,N_7665,N_7658);
nand U7851 (N_7851,N_7620,N_7502);
and U7852 (N_7852,N_7552,N_7524);
or U7853 (N_7853,N_7606,N_7699);
or U7854 (N_7854,N_7716,N_7646);
nor U7855 (N_7855,N_7745,N_7541);
nor U7856 (N_7856,N_7690,N_7705);
and U7857 (N_7857,N_7613,N_7512);
nand U7858 (N_7858,N_7719,N_7554);
or U7859 (N_7859,N_7581,N_7696);
xnor U7860 (N_7860,N_7659,N_7700);
and U7861 (N_7861,N_7637,N_7633);
xnor U7862 (N_7862,N_7503,N_7677);
xnor U7863 (N_7863,N_7567,N_7653);
or U7864 (N_7864,N_7560,N_7712);
or U7865 (N_7865,N_7632,N_7596);
xnor U7866 (N_7866,N_7539,N_7500);
xnor U7867 (N_7867,N_7553,N_7667);
nor U7868 (N_7868,N_7670,N_7534);
and U7869 (N_7869,N_7608,N_7731);
xnor U7870 (N_7870,N_7579,N_7546);
xor U7871 (N_7871,N_7673,N_7619);
and U7872 (N_7872,N_7666,N_7624);
and U7873 (N_7873,N_7748,N_7720);
or U7874 (N_7874,N_7583,N_7518);
or U7875 (N_7875,N_7620,N_7534);
nand U7876 (N_7876,N_7512,N_7516);
nand U7877 (N_7877,N_7508,N_7528);
and U7878 (N_7878,N_7504,N_7685);
xor U7879 (N_7879,N_7602,N_7746);
nor U7880 (N_7880,N_7587,N_7723);
or U7881 (N_7881,N_7520,N_7527);
or U7882 (N_7882,N_7582,N_7711);
nor U7883 (N_7883,N_7623,N_7527);
nor U7884 (N_7884,N_7647,N_7693);
nand U7885 (N_7885,N_7744,N_7670);
nor U7886 (N_7886,N_7626,N_7586);
nor U7887 (N_7887,N_7557,N_7504);
nand U7888 (N_7888,N_7656,N_7717);
xor U7889 (N_7889,N_7730,N_7646);
or U7890 (N_7890,N_7742,N_7644);
xnor U7891 (N_7891,N_7646,N_7569);
and U7892 (N_7892,N_7573,N_7671);
nand U7893 (N_7893,N_7651,N_7712);
nand U7894 (N_7894,N_7724,N_7534);
and U7895 (N_7895,N_7541,N_7657);
nand U7896 (N_7896,N_7607,N_7514);
or U7897 (N_7897,N_7628,N_7698);
and U7898 (N_7898,N_7544,N_7540);
nand U7899 (N_7899,N_7636,N_7565);
nand U7900 (N_7900,N_7661,N_7651);
nand U7901 (N_7901,N_7609,N_7613);
nor U7902 (N_7902,N_7729,N_7730);
nand U7903 (N_7903,N_7658,N_7629);
nor U7904 (N_7904,N_7653,N_7731);
or U7905 (N_7905,N_7732,N_7659);
nand U7906 (N_7906,N_7642,N_7561);
xor U7907 (N_7907,N_7697,N_7556);
and U7908 (N_7908,N_7716,N_7567);
or U7909 (N_7909,N_7720,N_7693);
nand U7910 (N_7910,N_7616,N_7612);
or U7911 (N_7911,N_7583,N_7727);
nand U7912 (N_7912,N_7687,N_7532);
or U7913 (N_7913,N_7607,N_7736);
or U7914 (N_7914,N_7702,N_7696);
xor U7915 (N_7915,N_7659,N_7569);
nand U7916 (N_7916,N_7718,N_7586);
xor U7917 (N_7917,N_7554,N_7652);
and U7918 (N_7918,N_7569,N_7729);
and U7919 (N_7919,N_7706,N_7703);
xnor U7920 (N_7920,N_7716,N_7545);
nand U7921 (N_7921,N_7573,N_7682);
xnor U7922 (N_7922,N_7601,N_7619);
and U7923 (N_7923,N_7678,N_7706);
nand U7924 (N_7924,N_7585,N_7659);
nand U7925 (N_7925,N_7632,N_7575);
or U7926 (N_7926,N_7708,N_7522);
xnor U7927 (N_7927,N_7713,N_7644);
nand U7928 (N_7928,N_7660,N_7574);
xnor U7929 (N_7929,N_7618,N_7577);
xnor U7930 (N_7930,N_7684,N_7729);
or U7931 (N_7931,N_7694,N_7522);
xnor U7932 (N_7932,N_7647,N_7524);
xor U7933 (N_7933,N_7624,N_7512);
nor U7934 (N_7934,N_7722,N_7731);
nor U7935 (N_7935,N_7583,N_7668);
nand U7936 (N_7936,N_7650,N_7513);
or U7937 (N_7937,N_7595,N_7691);
nand U7938 (N_7938,N_7723,N_7658);
xor U7939 (N_7939,N_7687,N_7673);
or U7940 (N_7940,N_7686,N_7726);
nand U7941 (N_7941,N_7700,N_7500);
xnor U7942 (N_7942,N_7549,N_7686);
and U7943 (N_7943,N_7635,N_7600);
or U7944 (N_7944,N_7628,N_7624);
and U7945 (N_7945,N_7555,N_7621);
nor U7946 (N_7946,N_7705,N_7666);
and U7947 (N_7947,N_7658,N_7632);
and U7948 (N_7948,N_7723,N_7581);
nand U7949 (N_7949,N_7662,N_7712);
nand U7950 (N_7950,N_7701,N_7606);
and U7951 (N_7951,N_7716,N_7692);
nor U7952 (N_7952,N_7744,N_7707);
nor U7953 (N_7953,N_7610,N_7730);
xnor U7954 (N_7954,N_7630,N_7532);
nor U7955 (N_7955,N_7667,N_7696);
and U7956 (N_7956,N_7556,N_7646);
and U7957 (N_7957,N_7676,N_7735);
xor U7958 (N_7958,N_7733,N_7645);
xnor U7959 (N_7959,N_7600,N_7506);
and U7960 (N_7960,N_7698,N_7730);
or U7961 (N_7961,N_7691,N_7600);
nand U7962 (N_7962,N_7680,N_7667);
nor U7963 (N_7963,N_7704,N_7690);
or U7964 (N_7964,N_7739,N_7714);
or U7965 (N_7965,N_7691,N_7731);
and U7966 (N_7966,N_7690,N_7551);
xnor U7967 (N_7967,N_7739,N_7564);
or U7968 (N_7968,N_7625,N_7737);
nor U7969 (N_7969,N_7708,N_7599);
and U7970 (N_7970,N_7529,N_7639);
or U7971 (N_7971,N_7726,N_7684);
nor U7972 (N_7972,N_7608,N_7717);
nand U7973 (N_7973,N_7616,N_7631);
nor U7974 (N_7974,N_7667,N_7559);
nand U7975 (N_7975,N_7698,N_7654);
and U7976 (N_7976,N_7655,N_7673);
nor U7977 (N_7977,N_7595,N_7507);
and U7978 (N_7978,N_7741,N_7634);
or U7979 (N_7979,N_7662,N_7670);
and U7980 (N_7980,N_7653,N_7639);
and U7981 (N_7981,N_7651,N_7730);
nor U7982 (N_7982,N_7704,N_7550);
xor U7983 (N_7983,N_7539,N_7515);
or U7984 (N_7984,N_7632,N_7673);
or U7985 (N_7985,N_7598,N_7603);
xor U7986 (N_7986,N_7550,N_7504);
or U7987 (N_7987,N_7712,N_7666);
nor U7988 (N_7988,N_7673,N_7645);
xor U7989 (N_7989,N_7577,N_7711);
xor U7990 (N_7990,N_7633,N_7678);
or U7991 (N_7991,N_7704,N_7726);
xnor U7992 (N_7992,N_7667,N_7652);
nor U7993 (N_7993,N_7563,N_7709);
nand U7994 (N_7994,N_7542,N_7658);
nand U7995 (N_7995,N_7595,N_7744);
nand U7996 (N_7996,N_7731,N_7515);
nor U7997 (N_7997,N_7544,N_7691);
nor U7998 (N_7998,N_7513,N_7528);
xor U7999 (N_7999,N_7566,N_7581);
xnor U8000 (N_8000,N_7899,N_7765);
or U8001 (N_8001,N_7945,N_7872);
or U8002 (N_8002,N_7982,N_7770);
or U8003 (N_8003,N_7835,N_7892);
nor U8004 (N_8004,N_7957,N_7831);
xnor U8005 (N_8005,N_7924,N_7841);
or U8006 (N_8006,N_7869,N_7907);
and U8007 (N_8007,N_7875,N_7920);
and U8008 (N_8008,N_7828,N_7790);
and U8009 (N_8009,N_7874,N_7755);
or U8010 (N_8010,N_7884,N_7888);
or U8011 (N_8011,N_7805,N_7904);
or U8012 (N_8012,N_7783,N_7999);
nand U8013 (N_8013,N_7962,N_7819);
or U8014 (N_8014,N_7991,N_7974);
xnor U8015 (N_8015,N_7840,N_7824);
nand U8016 (N_8016,N_7967,N_7791);
nand U8017 (N_8017,N_7988,N_7970);
nand U8018 (N_8018,N_7911,N_7782);
nor U8019 (N_8019,N_7871,N_7804);
nand U8020 (N_8020,N_7906,N_7788);
nand U8021 (N_8021,N_7898,N_7981);
nand U8022 (N_8022,N_7969,N_7921);
nand U8023 (N_8023,N_7860,N_7849);
and U8024 (N_8024,N_7777,N_7958);
xor U8025 (N_8025,N_7811,N_7933);
and U8026 (N_8026,N_7881,N_7918);
nand U8027 (N_8027,N_7803,N_7758);
xnor U8028 (N_8028,N_7902,N_7767);
nand U8029 (N_8029,N_7887,N_7810);
xor U8030 (N_8030,N_7822,N_7823);
xnor U8031 (N_8031,N_7814,N_7968);
and U8032 (N_8032,N_7943,N_7785);
nor U8033 (N_8033,N_7975,N_7763);
nor U8034 (N_8034,N_7926,N_7961);
nand U8035 (N_8035,N_7858,N_7886);
and U8036 (N_8036,N_7838,N_7784);
and U8037 (N_8037,N_7751,N_7890);
nand U8038 (N_8038,N_7854,N_7995);
xor U8039 (N_8039,N_7844,N_7948);
xnor U8040 (N_8040,N_7864,N_7793);
nor U8041 (N_8041,N_7885,N_7990);
or U8042 (N_8042,N_7753,N_7868);
xor U8043 (N_8043,N_7913,N_7837);
nand U8044 (N_8044,N_7927,N_7774);
or U8045 (N_8045,N_7772,N_7891);
or U8046 (N_8046,N_7759,N_7994);
xnor U8047 (N_8047,N_7873,N_7825);
nand U8048 (N_8048,N_7798,N_7951);
xnor U8049 (N_8049,N_7878,N_7925);
xnor U8050 (N_8050,N_7937,N_7983);
xor U8051 (N_8051,N_7909,N_7847);
nor U8052 (N_8052,N_7768,N_7977);
nand U8053 (N_8053,N_7773,N_7795);
or U8054 (N_8054,N_7963,N_7832);
xor U8055 (N_8055,N_7752,N_7972);
xnor U8056 (N_8056,N_7861,N_7857);
and U8057 (N_8057,N_7778,N_7809);
xnor U8058 (N_8058,N_7802,N_7946);
nand U8059 (N_8059,N_7756,N_7940);
or U8060 (N_8060,N_7930,N_7956);
and U8061 (N_8061,N_7905,N_7931);
or U8062 (N_8062,N_7808,N_7980);
and U8063 (N_8063,N_7914,N_7944);
nand U8064 (N_8064,N_7764,N_7880);
nor U8065 (N_8065,N_7923,N_7859);
nand U8066 (N_8066,N_7922,N_7987);
nor U8067 (N_8067,N_7820,N_7757);
or U8068 (N_8068,N_7817,N_7966);
xnor U8069 (N_8069,N_7992,N_7973);
nand U8070 (N_8070,N_7863,N_7776);
xor U8071 (N_8071,N_7794,N_7797);
xor U8072 (N_8072,N_7807,N_7912);
nor U8073 (N_8073,N_7771,N_7762);
xor U8074 (N_8074,N_7750,N_7845);
nand U8075 (N_8075,N_7928,N_7953);
and U8076 (N_8076,N_7754,N_7998);
nor U8077 (N_8077,N_7787,N_7942);
xnor U8078 (N_8078,N_7894,N_7896);
nor U8079 (N_8079,N_7936,N_7893);
or U8080 (N_8080,N_7939,N_7851);
and U8081 (N_8081,N_7766,N_7979);
nor U8082 (N_8082,N_7976,N_7935);
nor U8083 (N_8083,N_7842,N_7865);
nand U8084 (N_8084,N_7852,N_7836);
xor U8085 (N_8085,N_7846,N_7908);
nor U8086 (N_8086,N_7760,N_7806);
and U8087 (N_8087,N_7826,N_7917);
and U8088 (N_8088,N_7866,N_7781);
xor U8089 (N_8089,N_7816,N_7870);
nor U8090 (N_8090,N_7895,N_7856);
nor U8091 (N_8091,N_7883,N_7993);
xnor U8092 (N_8092,N_7789,N_7862);
or U8093 (N_8093,N_7949,N_7929);
nand U8094 (N_8094,N_7834,N_7761);
or U8095 (N_8095,N_7916,N_7952);
nor U8096 (N_8096,N_7978,N_7986);
xor U8097 (N_8097,N_7964,N_7959);
nand U8098 (N_8098,N_7934,N_7950);
nand U8099 (N_8099,N_7855,N_7843);
or U8100 (N_8100,N_7996,N_7786);
or U8101 (N_8101,N_7780,N_7897);
nand U8102 (N_8102,N_7901,N_7812);
xnor U8103 (N_8103,N_7867,N_7919);
and U8104 (N_8104,N_7900,N_7839);
and U8105 (N_8105,N_7938,N_7889);
and U8106 (N_8106,N_7960,N_7779);
and U8107 (N_8107,N_7821,N_7954);
xnor U8108 (N_8108,N_7829,N_7876);
nor U8109 (N_8109,N_7903,N_7915);
xnor U8110 (N_8110,N_7932,N_7853);
nand U8111 (N_8111,N_7792,N_7965);
and U8112 (N_8112,N_7955,N_7799);
and U8113 (N_8113,N_7910,N_7989);
xor U8114 (N_8114,N_7769,N_7941);
or U8115 (N_8115,N_7985,N_7947);
nor U8116 (N_8116,N_7850,N_7830);
nand U8117 (N_8117,N_7848,N_7833);
xnor U8118 (N_8118,N_7775,N_7800);
and U8119 (N_8119,N_7984,N_7815);
nor U8120 (N_8120,N_7796,N_7827);
xnor U8121 (N_8121,N_7882,N_7813);
or U8122 (N_8122,N_7877,N_7879);
and U8123 (N_8123,N_7971,N_7997);
or U8124 (N_8124,N_7818,N_7801);
nand U8125 (N_8125,N_7902,N_7997);
xor U8126 (N_8126,N_7801,N_7870);
and U8127 (N_8127,N_7881,N_7833);
nand U8128 (N_8128,N_7980,N_7947);
xnor U8129 (N_8129,N_7933,N_7754);
and U8130 (N_8130,N_7829,N_7825);
xnor U8131 (N_8131,N_7911,N_7825);
xor U8132 (N_8132,N_7762,N_7839);
nor U8133 (N_8133,N_7896,N_7801);
nor U8134 (N_8134,N_7799,N_7872);
xor U8135 (N_8135,N_7825,N_7877);
and U8136 (N_8136,N_7759,N_7960);
and U8137 (N_8137,N_7819,N_7806);
and U8138 (N_8138,N_7819,N_7794);
and U8139 (N_8139,N_7906,N_7763);
nand U8140 (N_8140,N_7908,N_7826);
and U8141 (N_8141,N_7845,N_7900);
and U8142 (N_8142,N_7936,N_7869);
nand U8143 (N_8143,N_7921,N_7964);
nand U8144 (N_8144,N_7832,N_7750);
and U8145 (N_8145,N_7908,N_7898);
and U8146 (N_8146,N_7931,N_7844);
and U8147 (N_8147,N_7981,N_7804);
nor U8148 (N_8148,N_7772,N_7862);
xnor U8149 (N_8149,N_7991,N_7832);
and U8150 (N_8150,N_7991,N_7951);
or U8151 (N_8151,N_7801,N_7763);
and U8152 (N_8152,N_7810,N_7920);
or U8153 (N_8153,N_7984,N_7972);
nor U8154 (N_8154,N_7952,N_7890);
nand U8155 (N_8155,N_7818,N_7969);
nand U8156 (N_8156,N_7909,N_7897);
xnor U8157 (N_8157,N_7790,N_7822);
or U8158 (N_8158,N_7828,N_7882);
nor U8159 (N_8159,N_7997,N_7789);
nand U8160 (N_8160,N_7845,N_7753);
and U8161 (N_8161,N_7954,N_7935);
and U8162 (N_8162,N_7960,N_7767);
xnor U8163 (N_8163,N_7938,N_7826);
nand U8164 (N_8164,N_7998,N_7928);
and U8165 (N_8165,N_7829,N_7901);
nand U8166 (N_8166,N_7788,N_7959);
xnor U8167 (N_8167,N_7980,N_7796);
xnor U8168 (N_8168,N_7948,N_7838);
nand U8169 (N_8169,N_7941,N_7798);
or U8170 (N_8170,N_7984,N_7848);
xnor U8171 (N_8171,N_7962,N_7760);
or U8172 (N_8172,N_7899,N_7891);
nor U8173 (N_8173,N_7968,N_7764);
or U8174 (N_8174,N_7912,N_7896);
nor U8175 (N_8175,N_7777,N_7791);
xor U8176 (N_8176,N_7802,N_7824);
xnor U8177 (N_8177,N_7933,N_7859);
nor U8178 (N_8178,N_7954,N_7970);
xnor U8179 (N_8179,N_7840,N_7852);
or U8180 (N_8180,N_7937,N_7876);
nand U8181 (N_8181,N_7904,N_7802);
nand U8182 (N_8182,N_7902,N_7930);
and U8183 (N_8183,N_7961,N_7934);
and U8184 (N_8184,N_7831,N_7886);
and U8185 (N_8185,N_7870,N_7848);
xor U8186 (N_8186,N_7992,N_7928);
nand U8187 (N_8187,N_7968,N_7793);
nor U8188 (N_8188,N_7932,N_7957);
nand U8189 (N_8189,N_7815,N_7993);
or U8190 (N_8190,N_7989,N_7938);
xnor U8191 (N_8191,N_7845,N_7799);
nor U8192 (N_8192,N_7876,N_7839);
nand U8193 (N_8193,N_7782,N_7846);
xor U8194 (N_8194,N_7981,N_7767);
or U8195 (N_8195,N_7757,N_7848);
or U8196 (N_8196,N_7805,N_7865);
xnor U8197 (N_8197,N_7975,N_7882);
or U8198 (N_8198,N_7915,N_7919);
xnor U8199 (N_8199,N_7918,N_7775);
or U8200 (N_8200,N_7791,N_7906);
nand U8201 (N_8201,N_7962,N_7782);
and U8202 (N_8202,N_7767,N_7918);
nand U8203 (N_8203,N_7932,N_7820);
or U8204 (N_8204,N_7926,N_7884);
xor U8205 (N_8205,N_7872,N_7816);
nand U8206 (N_8206,N_7982,N_7828);
or U8207 (N_8207,N_7960,N_7984);
and U8208 (N_8208,N_7802,N_7968);
and U8209 (N_8209,N_7943,N_7877);
nand U8210 (N_8210,N_7910,N_7914);
or U8211 (N_8211,N_7841,N_7928);
xor U8212 (N_8212,N_7833,N_7774);
nand U8213 (N_8213,N_7905,N_7753);
nor U8214 (N_8214,N_7773,N_7770);
nor U8215 (N_8215,N_7789,N_7949);
and U8216 (N_8216,N_7963,N_7997);
nand U8217 (N_8217,N_7794,N_7791);
xor U8218 (N_8218,N_7850,N_7762);
nand U8219 (N_8219,N_7841,N_7769);
nand U8220 (N_8220,N_7966,N_7928);
and U8221 (N_8221,N_7974,N_7948);
nand U8222 (N_8222,N_7799,N_7930);
xor U8223 (N_8223,N_7996,N_7929);
nor U8224 (N_8224,N_7955,N_7782);
nand U8225 (N_8225,N_7931,N_7956);
xor U8226 (N_8226,N_7897,N_7768);
nor U8227 (N_8227,N_7837,N_7936);
nor U8228 (N_8228,N_7792,N_7781);
and U8229 (N_8229,N_7976,N_7760);
and U8230 (N_8230,N_7961,N_7959);
and U8231 (N_8231,N_7899,N_7869);
nor U8232 (N_8232,N_7930,N_7977);
xor U8233 (N_8233,N_7806,N_7763);
xnor U8234 (N_8234,N_7893,N_7933);
nand U8235 (N_8235,N_7755,N_7885);
nor U8236 (N_8236,N_7967,N_7812);
and U8237 (N_8237,N_7816,N_7973);
nor U8238 (N_8238,N_7969,N_7821);
xnor U8239 (N_8239,N_7789,N_7843);
xor U8240 (N_8240,N_7789,N_7965);
xnor U8241 (N_8241,N_7756,N_7859);
xor U8242 (N_8242,N_7768,N_7988);
and U8243 (N_8243,N_7878,N_7852);
nand U8244 (N_8244,N_7782,N_7900);
nand U8245 (N_8245,N_7766,N_7775);
xor U8246 (N_8246,N_7763,N_7978);
xor U8247 (N_8247,N_7764,N_7843);
and U8248 (N_8248,N_7958,N_7929);
nor U8249 (N_8249,N_7757,N_7756);
xnor U8250 (N_8250,N_8228,N_8188);
nor U8251 (N_8251,N_8242,N_8244);
or U8252 (N_8252,N_8074,N_8180);
and U8253 (N_8253,N_8078,N_8010);
or U8254 (N_8254,N_8235,N_8050);
xor U8255 (N_8255,N_8229,N_8088);
xnor U8256 (N_8256,N_8239,N_8012);
nand U8257 (N_8257,N_8245,N_8029);
xnor U8258 (N_8258,N_8182,N_8051);
or U8259 (N_8259,N_8001,N_8038);
xnor U8260 (N_8260,N_8045,N_8137);
xnor U8261 (N_8261,N_8062,N_8067);
nand U8262 (N_8262,N_8119,N_8141);
nor U8263 (N_8263,N_8020,N_8130);
or U8264 (N_8264,N_8087,N_8168);
xnor U8265 (N_8265,N_8146,N_8004);
nand U8266 (N_8266,N_8128,N_8124);
nand U8267 (N_8267,N_8200,N_8063);
nand U8268 (N_8268,N_8216,N_8083);
xor U8269 (N_8269,N_8129,N_8201);
xor U8270 (N_8270,N_8014,N_8054);
or U8271 (N_8271,N_8175,N_8032);
nor U8272 (N_8272,N_8060,N_8121);
nor U8273 (N_8273,N_8003,N_8217);
xor U8274 (N_8274,N_8034,N_8234);
nor U8275 (N_8275,N_8036,N_8084);
and U8276 (N_8276,N_8043,N_8006);
nand U8277 (N_8277,N_8132,N_8222);
xnor U8278 (N_8278,N_8184,N_8098);
and U8279 (N_8279,N_8136,N_8196);
xnor U8280 (N_8280,N_8225,N_8172);
or U8281 (N_8281,N_8241,N_8199);
nor U8282 (N_8282,N_8071,N_8076);
nand U8283 (N_8283,N_8169,N_8072);
xnor U8284 (N_8284,N_8171,N_8191);
nor U8285 (N_8285,N_8024,N_8149);
or U8286 (N_8286,N_8185,N_8125);
nor U8287 (N_8287,N_8215,N_8041);
and U8288 (N_8288,N_8138,N_8077);
and U8289 (N_8289,N_8070,N_8114);
xor U8290 (N_8290,N_8106,N_8120);
xor U8291 (N_8291,N_8056,N_8019);
nor U8292 (N_8292,N_8008,N_8194);
and U8293 (N_8293,N_8118,N_8123);
or U8294 (N_8294,N_8190,N_8248);
or U8295 (N_8295,N_8107,N_8101);
and U8296 (N_8296,N_8142,N_8179);
and U8297 (N_8297,N_8047,N_8150);
xnor U8298 (N_8298,N_8134,N_8237);
and U8299 (N_8299,N_8233,N_8213);
or U8300 (N_8300,N_8156,N_8195);
nor U8301 (N_8301,N_8207,N_8000);
nand U8302 (N_8302,N_8193,N_8144);
nand U8303 (N_8303,N_8174,N_8218);
xor U8304 (N_8304,N_8173,N_8040);
nand U8305 (N_8305,N_8075,N_8057);
or U8306 (N_8306,N_8249,N_8203);
xnor U8307 (N_8307,N_8095,N_8015);
or U8308 (N_8308,N_8048,N_8011);
nor U8309 (N_8309,N_8122,N_8031);
or U8310 (N_8310,N_8167,N_8065);
nand U8311 (N_8311,N_8105,N_8025);
or U8312 (N_8312,N_8178,N_8037);
nor U8313 (N_8313,N_8064,N_8127);
nor U8314 (N_8314,N_8018,N_8022);
or U8315 (N_8315,N_8177,N_8210);
xor U8316 (N_8316,N_8214,N_8086);
and U8317 (N_8317,N_8186,N_8163);
or U8318 (N_8318,N_8027,N_8104);
or U8319 (N_8319,N_8073,N_8230);
nand U8320 (N_8320,N_8231,N_8209);
nand U8321 (N_8321,N_8165,N_8108);
nand U8322 (N_8322,N_8079,N_8017);
nand U8323 (N_8323,N_8223,N_8133);
and U8324 (N_8324,N_8154,N_8147);
nand U8325 (N_8325,N_8059,N_8166);
and U8326 (N_8326,N_8189,N_8139);
and U8327 (N_8327,N_8109,N_8126);
and U8328 (N_8328,N_8091,N_8205);
nor U8329 (N_8329,N_8159,N_8090);
xnor U8330 (N_8330,N_8145,N_8198);
nor U8331 (N_8331,N_8042,N_8092);
nand U8332 (N_8332,N_8009,N_8227);
xnor U8333 (N_8333,N_8023,N_8080);
and U8334 (N_8334,N_8183,N_8208);
nand U8335 (N_8335,N_8033,N_8030);
xnor U8336 (N_8336,N_8096,N_8102);
nand U8337 (N_8337,N_8143,N_8164);
nor U8338 (N_8338,N_8093,N_8116);
nor U8339 (N_8339,N_8204,N_8002);
or U8340 (N_8340,N_8247,N_8066);
or U8341 (N_8341,N_8240,N_8021);
xnor U8342 (N_8342,N_8148,N_8155);
and U8343 (N_8343,N_8158,N_8243);
and U8344 (N_8344,N_8206,N_8028);
xnor U8345 (N_8345,N_8151,N_8152);
xnor U8346 (N_8346,N_8046,N_8157);
nor U8347 (N_8347,N_8140,N_8085);
or U8348 (N_8348,N_8005,N_8007);
xnor U8349 (N_8349,N_8100,N_8115);
or U8350 (N_8350,N_8112,N_8238);
and U8351 (N_8351,N_8068,N_8232);
or U8352 (N_8352,N_8170,N_8013);
nand U8353 (N_8353,N_8246,N_8160);
nor U8354 (N_8354,N_8176,N_8181);
nor U8355 (N_8355,N_8153,N_8192);
xor U8356 (N_8356,N_8081,N_8058);
nand U8357 (N_8357,N_8049,N_8039);
and U8358 (N_8358,N_8224,N_8221);
xor U8359 (N_8359,N_8055,N_8111);
or U8360 (N_8360,N_8131,N_8035);
nor U8361 (N_8361,N_8082,N_8061);
and U8362 (N_8362,N_8103,N_8211);
xnor U8363 (N_8363,N_8161,N_8212);
xnor U8364 (N_8364,N_8197,N_8089);
nor U8365 (N_8365,N_8162,N_8044);
nand U8366 (N_8366,N_8187,N_8016);
nand U8367 (N_8367,N_8117,N_8053);
xnor U8368 (N_8368,N_8094,N_8202);
xnor U8369 (N_8369,N_8219,N_8135);
xnor U8370 (N_8370,N_8052,N_8220);
nand U8371 (N_8371,N_8226,N_8069);
nand U8372 (N_8372,N_8236,N_8110);
and U8373 (N_8373,N_8026,N_8113);
xnor U8374 (N_8374,N_8099,N_8097);
or U8375 (N_8375,N_8058,N_8084);
nand U8376 (N_8376,N_8132,N_8061);
xnor U8377 (N_8377,N_8133,N_8020);
xnor U8378 (N_8378,N_8118,N_8162);
and U8379 (N_8379,N_8135,N_8152);
and U8380 (N_8380,N_8047,N_8009);
xnor U8381 (N_8381,N_8147,N_8242);
xnor U8382 (N_8382,N_8225,N_8113);
or U8383 (N_8383,N_8038,N_8091);
nor U8384 (N_8384,N_8028,N_8129);
nor U8385 (N_8385,N_8201,N_8245);
or U8386 (N_8386,N_8037,N_8195);
xor U8387 (N_8387,N_8054,N_8170);
or U8388 (N_8388,N_8156,N_8031);
and U8389 (N_8389,N_8215,N_8108);
nand U8390 (N_8390,N_8165,N_8215);
xor U8391 (N_8391,N_8030,N_8015);
and U8392 (N_8392,N_8226,N_8002);
nor U8393 (N_8393,N_8230,N_8052);
xnor U8394 (N_8394,N_8042,N_8172);
nand U8395 (N_8395,N_8076,N_8011);
or U8396 (N_8396,N_8234,N_8123);
nor U8397 (N_8397,N_8075,N_8113);
nand U8398 (N_8398,N_8241,N_8202);
or U8399 (N_8399,N_8056,N_8129);
nand U8400 (N_8400,N_8224,N_8151);
or U8401 (N_8401,N_8241,N_8110);
or U8402 (N_8402,N_8230,N_8032);
xor U8403 (N_8403,N_8160,N_8079);
and U8404 (N_8404,N_8049,N_8184);
and U8405 (N_8405,N_8113,N_8060);
or U8406 (N_8406,N_8180,N_8090);
and U8407 (N_8407,N_8043,N_8157);
or U8408 (N_8408,N_8115,N_8125);
nand U8409 (N_8409,N_8186,N_8087);
and U8410 (N_8410,N_8053,N_8191);
xor U8411 (N_8411,N_8138,N_8192);
and U8412 (N_8412,N_8114,N_8028);
and U8413 (N_8413,N_8119,N_8015);
nor U8414 (N_8414,N_8008,N_8109);
nand U8415 (N_8415,N_8078,N_8221);
nand U8416 (N_8416,N_8020,N_8228);
or U8417 (N_8417,N_8015,N_8201);
nand U8418 (N_8418,N_8220,N_8071);
nand U8419 (N_8419,N_8060,N_8207);
or U8420 (N_8420,N_8188,N_8077);
and U8421 (N_8421,N_8087,N_8152);
xnor U8422 (N_8422,N_8233,N_8090);
xnor U8423 (N_8423,N_8181,N_8035);
or U8424 (N_8424,N_8241,N_8112);
nor U8425 (N_8425,N_8020,N_8189);
and U8426 (N_8426,N_8156,N_8173);
nor U8427 (N_8427,N_8187,N_8149);
nand U8428 (N_8428,N_8247,N_8089);
xnor U8429 (N_8429,N_8100,N_8049);
xnor U8430 (N_8430,N_8035,N_8165);
xor U8431 (N_8431,N_8135,N_8025);
and U8432 (N_8432,N_8033,N_8014);
nor U8433 (N_8433,N_8133,N_8038);
xnor U8434 (N_8434,N_8047,N_8180);
nor U8435 (N_8435,N_8239,N_8090);
and U8436 (N_8436,N_8173,N_8239);
xnor U8437 (N_8437,N_8120,N_8027);
xnor U8438 (N_8438,N_8155,N_8018);
nor U8439 (N_8439,N_8085,N_8222);
nand U8440 (N_8440,N_8122,N_8132);
nor U8441 (N_8441,N_8217,N_8202);
nand U8442 (N_8442,N_8075,N_8055);
xor U8443 (N_8443,N_8006,N_8169);
or U8444 (N_8444,N_8023,N_8028);
or U8445 (N_8445,N_8244,N_8249);
nor U8446 (N_8446,N_8119,N_8159);
xnor U8447 (N_8447,N_8205,N_8084);
and U8448 (N_8448,N_8078,N_8175);
xnor U8449 (N_8449,N_8057,N_8109);
and U8450 (N_8450,N_8210,N_8048);
xor U8451 (N_8451,N_8081,N_8138);
nor U8452 (N_8452,N_8115,N_8249);
nand U8453 (N_8453,N_8235,N_8216);
xnor U8454 (N_8454,N_8134,N_8191);
and U8455 (N_8455,N_8088,N_8041);
xnor U8456 (N_8456,N_8043,N_8183);
nor U8457 (N_8457,N_8036,N_8079);
or U8458 (N_8458,N_8104,N_8021);
and U8459 (N_8459,N_8147,N_8013);
and U8460 (N_8460,N_8213,N_8146);
and U8461 (N_8461,N_8042,N_8088);
nor U8462 (N_8462,N_8137,N_8231);
nor U8463 (N_8463,N_8041,N_8015);
nor U8464 (N_8464,N_8232,N_8080);
nand U8465 (N_8465,N_8216,N_8073);
nand U8466 (N_8466,N_8085,N_8167);
and U8467 (N_8467,N_8243,N_8155);
xnor U8468 (N_8468,N_8150,N_8192);
nand U8469 (N_8469,N_8030,N_8040);
and U8470 (N_8470,N_8165,N_8141);
nor U8471 (N_8471,N_8020,N_8005);
nand U8472 (N_8472,N_8018,N_8071);
xor U8473 (N_8473,N_8146,N_8244);
xnor U8474 (N_8474,N_8196,N_8138);
or U8475 (N_8475,N_8194,N_8248);
nor U8476 (N_8476,N_8169,N_8019);
xnor U8477 (N_8477,N_8240,N_8159);
and U8478 (N_8478,N_8074,N_8097);
nor U8479 (N_8479,N_8011,N_8030);
nor U8480 (N_8480,N_8063,N_8098);
xnor U8481 (N_8481,N_8191,N_8212);
nand U8482 (N_8482,N_8223,N_8106);
nor U8483 (N_8483,N_8096,N_8115);
and U8484 (N_8484,N_8101,N_8029);
or U8485 (N_8485,N_8228,N_8187);
and U8486 (N_8486,N_8045,N_8125);
xnor U8487 (N_8487,N_8090,N_8162);
or U8488 (N_8488,N_8235,N_8133);
or U8489 (N_8489,N_8106,N_8221);
xor U8490 (N_8490,N_8014,N_8155);
xor U8491 (N_8491,N_8117,N_8086);
nand U8492 (N_8492,N_8048,N_8022);
and U8493 (N_8493,N_8019,N_8079);
nor U8494 (N_8494,N_8057,N_8000);
nor U8495 (N_8495,N_8106,N_8171);
or U8496 (N_8496,N_8012,N_8110);
nor U8497 (N_8497,N_8151,N_8145);
or U8498 (N_8498,N_8164,N_8121);
or U8499 (N_8499,N_8026,N_8220);
xor U8500 (N_8500,N_8250,N_8253);
or U8501 (N_8501,N_8283,N_8369);
and U8502 (N_8502,N_8440,N_8328);
and U8503 (N_8503,N_8384,N_8436);
and U8504 (N_8504,N_8399,N_8289);
and U8505 (N_8505,N_8290,N_8373);
and U8506 (N_8506,N_8458,N_8464);
and U8507 (N_8507,N_8450,N_8404);
xor U8508 (N_8508,N_8459,N_8262);
or U8509 (N_8509,N_8340,N_8318);
xor U8510 (N_8510,N_8371,N_8461);
xnor U8511 (N_8511,N_8447,N_8357);
and U8512 (N_8512,N_8286,N_8346);
nor U8513 (N_8513,N_8417,N_8396);
nand U8514 (N_8514,N_8493,N_8266);
and U8515 (N_8515,N_8293,N_8301);
xor U8516 (N_8516,N_8356,N_8261);
or U8517 (N_8517,N_8398,N_8383);
nor U8518 (N_8518,N_8496,N_8341);
nand U8519 (N_8519,N_8326,N_8263);
and U8520 (N_8520,N_8403,N_8278);
nand U8521 (N_8521,N_8377,N_8457);
or U8522 (N_8522,N_8470,N_8315);
and U8523 (N_8523,N_8406,N_8338);
xnor U8524 (N_8524,N_8255,N_8280);
xnor U8525 (N_8525,N_8479,N_8355);
and U8526 (N_8526,N_8478,N_8305);
xnor U8527 (N_8527,N_8390,N_8313);
and U8528 (N_8528,N_8385,N_8425);
and U8529 (N_8529,N_8325,N_8468);
or U8530 (N_8530,N_8499,N_8471);
xnor U8531 (N_8531,N_8343,N_8473);
xnor U8532 (N_8532,N_8310,N_8448);
nor U8533 (N_8533,N_8484,N_8257);
and U8534 (N_8534,N_8363,N_8292);
or U8535 (N_8535,N_8296,N_8317);
or U8536 (N_8536,N_8455,N_8364);
or U8537 (N_8537,N_8433,N_8347);
nor U8538 (N_8538,N_8467,N_8462);
nand U8539 (N_8539,N_8392,N_8449);
or U8540 (N_8540,N_8432,N_8402);
and U8541 (N_8541,N_8258,N_8331);
and U8542 (N_8542,N_8451,N_8276);
and U8543 (N_8543,N_8423,N_8434);
nor U8544 (N_8544,N_8274,N_8490);
and U8545 (N_8545,N_8372,N_8441);
nor U8546 (N_8546,N_8422,N_8316);
and U8547 (N_8547,N_8264,N_8345);
nor U8548 (N_8548,N_8307,N_8486);
or U8549 (N_8549,N_8379,N_8285);
and U8550 (N_8550,N_8472,N_8270);
and U8551 (N_8551,N_8284,N_8495);
nand U8552 (N_8552,N_8420,N_8424);
xnor U8553 (N_8553,N_8498,N_8311);
nand U8554 (N_8554,N_8275,N_8314);
xnor U8555 (N_8555,N_8446,N_8438);
xnor U8556 (N_8556,N_8352,N_8351);
xnor U8557 (N_8557,N_8342,N_8251);
nor U8558 (N_8558,N_8330,N_8463);
nor U8559 (N_8559,N_8329,N_8295);
or U8560 (N_8560,N_8456,N_8437);
or U8561 (N_8561,N_8271,N_8312);
nand U8562 (N_8562,N_8485,N_8254);
nand U8563 (N_8563,N_8435,N_8322);
xor U8564 (N_8564,N_8426,N_8297);
nand U8565 (N_8565,N_8260,N_8308);
nor U8566 (N_8566,N_8302,N_8411);
nand U8567 (N_8567,N_8413,N_8487);
nand U8568 (N_8568,N_8454,N_8494);
and U8569 (N_8569,N_8335,N_8367);
and U8570 (N_8570,N_8349,N_8475);
nor U8571 (N_8571,N_8469,N_8419);
nor U8572 (N_8572,N_8272,N_8460);
xor U8573 (N_8573,N_8304,N_8334);
nand U8574 (N_8574,N_8418,N_8482);
xnor U8575 (N_8575,N_8442,N_8353);
nor U8576 (N_8576,N_8393,N_8386);
nor U8577 (N_8577,N_8430,N_8474);
nand U8578 (N_8578,N_8374,N_8282);
xnor U8579 (N_8579,N_8465,N_8332);
xor U8580 (N_8580,N_8412,N_8466);
nor U8581 (N_8581,N_8376,N_8256);
nor U8582 (N_8582,N_8439,N_8327);
nor U8583 (N_8583,N_8344,N_8303);
nand U8584 (N_8584,N_8323,N_8281);
and U8585 (N_8585,N_8294,N_8333);
nor U8586 (N_8586,N_8480,N_8336);
and U8587 (N_8587,N_8387,N_8259);
nand U8588 (N_8588,N_8299,N_8319);
xor U8589 (N_8589,N_8415,N_8416);
xor U8590 (N_8590,N_8414,N_8429);
or U8591 (N_8591,N_8277,N_8300);
nor U8592 (N_8592,N_8348,N_8324);
or U8593 (N_8593,N_8444,N_8267);
nor U8594 (N_8594,N_8408,N_8269);
and U8595 (N_8595,N_8443,N_8358);
or U8596 (N_8596,N_8394,N_8400);
nor U8597 (N_8597,N_8361,N_8375);
or U8598 (N_8598,N_8427,N_8306);
and U8599 (N_8599,N_8350,N_8291);
xor U8600 (N_8600,N_8339,N_8483);
xnor U8601 (N_8601,N_8407,N_8431);
and U8602 (N_8602,N_8477,N_8320);
xnor U8603 (N_8603,N_8481,N_8288);
nand U8604 (N_8604,N_8382,N_8287);
xor U8605 (N_8605,N_8410,N_8359);
xnor U8606 (N_8606,N_8497,N_8362);
xor U8607 (N_8607,N_8368,N_8378);
and U8608 (N_8608,N_8445,N_8405);
or U8609 (N_8609,N_8252,N_8365);
xor U8610 (N_8610,N_8279,N_8492);
nor U8611 (N_8611,N_8491,N_8452);
and U8612 (N_8612,N_8421,N_8453);
and U8613 (N_8613,N_8273,N_8476);
and U8614 (N_8614,N_8409,N_8389);
xnor U8615 (N_8615,N_8370,N_8397);
nand U8616 (N_8616,N_8395,N_8309);
xor U8617 (N_8617,N_8381,N_8488);
xnor U8618 (N_8618,N_8388,N_8401);
xnor U8619 (N_8619,N_8428,N_8268);
nor U8620 (N_8620,N_8298,N_8354);
or U8621 (N_8621,N_8391,N_8337);
xor U8622 (N_8622,N_8321,N_8380);
or U8623 (N_8623,N_8366,N_8489);
nand U8624 (N_8624,N_8360,N_8265);
or U8625 (N_8625,N_8377,N_8494);
xor U8626 (N_8626,N_8255,N_8275);
xor U8627 (N_8627,N_8318,N_8307);
or U8628 (N_8628,N_8398,N_8323);
and U8629 (N_8629,N_8270,N_8404);
xor U8630 (N_8630,N_8476,N_8409);
and U8631 (N_8631,N_8309,N_8252);
or U8632 (N_8632,N_8433,N_8294);
and U8633 (N_8633,N_8288,N_8342);
or U8634 (N_8634,N_8362,N_8421);
or U8635 (N_8635,N_8383,N_8257);
nand U8636 (N_8636,N_8252,N_8314);
xor U8637 (N_8637,N_8307,N_8434);
or U8638 (N_8638,N_8471,N_8321);
nor U8639 (N_8639,N_8382,N_8360);
nand U8640 (N_8640,N_8275,N_8448);
and U8641 (N_8641,N_8469,N_8372);
nor U8642 (N_8642,N_8288,N_8304);
nor U8643 (N_8643,N_8469,N_8322);
nor U8644 (N_8644,N_8345,N_8313);
xor U8645 (N_8645,N_8456,N_8288);
xor U8646 (N_8646,N_8386,N_8320);
nand U8647 (N_8647,N_8430,N_8256);
xnor U8648 (N_8648,N_8414,N_8280);
or U8649 (N_8649,N_8296,N_8442);
nand U8650 (N_8650,N_8309,N_8383);
xor U8651 (N_8651,N_8416,N_8457);
and U8652 (N_8652,N_8446,N_8352);
nand U8653 (N_8653,N_8379,N_8281);
nor U8654 (N_8654,N_8301,N_8477);
xor U8655 (N_8655,N_8387,N_8365);
or U8656 (N_8656,N_8429,N_8390);
and U8657 (N_8657,N_8433,N_8349);
nand U8658 (N_8658,N_8437,N_8274);
nor U8659 (N_8659,N_8324,N_8428);
and U8660 (N_8660,N_8321,N_8350);
or U8661 (N_8661,N_8343,N_8273);
xnor U8662 (N_8662,N_8379,N_8443);
xor U8663 (N_8663,N_8252,N_8301);
and U8664 (N_8664,N_8386,N_8343);
or U8665 (N_8665,N_8425,N_8369);
and U8666 (N_8666,N_8397,N_8452);
xor U8667 (N_8667,N_8471,N_8445);
nand U8668 (N_8668,N_8402,N_8466);
nand U8669 (N_8669,N_8257,N_8498);
or U8670 (N_8670,N_8476,N_8368);
nand U8671 (N_8671,N_8448,N_8427);
xor U8672 (N_8672,N_8250,N_8479);
nand U8673 (N_8673,N_8299,N_8414);
and U8674 (N_8674,N_8296,N_8470);
nor U8675 (N_8675,N_8430,N_8257);
xor U8676 (N_8676,N_8300,N_8427);
or U8677 (N_8677,N_8261,N_8264);
and U8678 (N_8678,N_8264,N_8349);
nand U8679 (N_8679,N_8268,N_8498);
nand U8680 (N_8680,N_8269,N_8416);
or U8681 (N_8681,N_8309,N_8455);
or U8682 (N_8682,N_8355,N_8343);
xor U8683 (N_8683,N_8375,N_8479);
xnor U8684 (N_8684,N_8409,N_8452);
xnor U8685 (N_8685,N_8464,N_8421);
and U8686 (N_8686,N_8317,N_8300);
nor U8687 (N_8687,N_8330,N_8312);
nand U8688 (N_8688,N_8496,N_8382);
nor U8689 (N_8689,N_8497,N_8351);
or U8690 (N_8690,N_8493,N_8380);
nand U8691 (N_8691,N_8283,N_8345);
nand U8692 (N_8692,N_8370,N_8361);
and U8693 (N_8693,N_8471,N_8416);
and U8694 (N_8694,N_8426,N_8251);
nand U8695 (N_8695,N_8497,N_8405);
xnor U8696 (N_8696,N_8356,N_8460);
nor U8697 (N_8697,N_8259,N_8358);
xnor U8698 (N_8698,N_8289,N_8450);
nand U8699 (N_8699,N_8369,N_8287);
nor U8700 (N_8700,N_8354,N_8482);
xor U8701 (N_8701,N_8402,N_8407);
or U8702 (N_8702,N_8403,N_8482);
nor U8703 (N_8703,N_8401,N_8472);
and U8704 (N_8704,N_8417,N_8391);
xnor U8705 (N_8705,N_8455,N_8486);
xnor U8706 (N_8706,N_8467,N_8495);
nand U8707 (N_8707,N_8405,N_8296);
and U8708 (N_8708,N_8272,N_8413);
nand U8709 (N_8709,N_8333,N_8445);
nand U8710 (N_8710,N_8444,N_8472);
or U8711 (N_8711,N_8303,N_8257);
or U8712 (N_8712,N_8292,N_8301);
nor U8713 (N_8713,N_8315,N_8371);
and U8714 (N_8714,N_8268,N_8488);
nor U8715 (N_8715,N_8414,N_8423);
nor U8716 (N_8716,N_8489,N_8325);
or U8717 (N_8717,N_8446,N_8310);
xnor U8718 (N_8718,N_8435,N_8471);
nor U8719 (N_8719,N_8410,N_8485);
xnor U8720 (N_8720,N_8309,N_8467);
and U8721 (N_8721,N_8440,N_8391);
nor U8722 (N_8722,N_8275,N_8326);
and U8723 (N_8723,N_8459,N_8347);
or U8724 (N_8724,N_8422,N_8327);
nand U8725 (N_8725,N_8473,N_8394);
and U8726 (N_8726,N_8415,N_8344);
nor U8727 (N_8727,N_8457,N_8310);
nand U8728 (N_8728,N_8416,N_8317);
xor U8729 (N_8729,N_8416,N_8321);
or U8730 (N_8730,N_8271,N_8359);
or U8731 (N_8731,N_8423,N_8362);
and U8732 (N_8732,N_8321,N_8406);
and U8733 (N_8733,N_8263,N_8365);
xnor U8734 (N_8734,N_8272,N_8270);
or U8735 (N_8735,N_8464,N_8325);
or U8736 (N_8736,N_8293,N_8373);
nor U8737 (N_8737,N_8366,N_8450);
or U8738 (N_8738,N_8341,N_8474);
and U8739 (N_8739,N_8379,N_8355);
nand U8740 (N_8740,N_8466,N_8497);
and U8741 (N_8741,N_8300,N_8297);
nand U8742 (N_8742,N_8426,N_8267);
nand U8743 (N_8743,N_8458,N_8280);
nor U8744 (N_8744,N_8418,N_8385);
or U8745 (N_8745,N_8352,N_8395);
nand U8746 (N_8746,N_8463,N_8472);
xor U8747 (N_8747,N_8289,N_8407);
xor U8748 (N_8748,N_8299,N_8281);
xnor U8749 (N_8749,N_8277,N_8258);
or U8750 (N_8750,N_8592,N_8501);
nand U8751 (N_8751,N_8560,N_8661);
or U8752 (N_8752,N_8637,N_8660);
nor U8753 (N_8753,N_8503,N_8509);
xor U8754 (N_8754,N_8571,N_8574);
nor U8755 (N_8755,N_8718,N_8628);
and U8756 (N_8756,N_8566,N_8720);
or U8757 (N_8757,N_8506,N_8572);
and U8758 (N_8758,N_8589,N_8519);
xor U8759 (N_8759,N_8645,N_8740);
nand U8760 (N_8760,N_8601,N_8714);
nor U8761 (N_8761,N_8694,N_8521);
or U8762 (N_8762,N_8692,N_8688);
nor U8763 (N_8763,N_8553,N_8681);
nor U8764 (N_8764,N_8656,N_8596);
or U8765 (N_8765,N_8626,N_8742);
or U8766 (N_8766,N_8723,N_8726);
and U8767 (N_8767,N_8543,N_8607);
and U8768 (N_8768,N_8559,N_8582);
xor U8769 (N_8769,N_8548,N_8747);
nor U8770 (N_8770,N_8530,N_8642);
or U8771 (N_8771,N_8508,N_8616);
nand U8772 (N_8772,N_8654,N_8513);
and U8773 (N_8773,N_8665,N_8526);
and U8774 (N_8774,N_8746,N_8691);
or U8775 (N_8775,N_8536,N_8672);
or U8776 (N_8776,N_8658,N_8563);
nand U8777 (N_8777,N_8732,N_8625);
xor U8778 (N_8778,N_8611,N_8550);
xnor U8779 (N_8779,N_8738,N_8593);
xor U8780 (N_8780,N_8554,N_8523);
nand U8781 (N_8781,N_8657,N_8734);
or U8782 (N_8782,N_8729,N_8659);
xnor U8783 (N_8783,N_8520,N_8619);
nor U8784 (N_8784,N_8635,N_8664);
nand U8785 (N_8785,N_8675,N_8748);
nor U8786 (N_8786,N_8695,N_8666);
nand U8787 (N_8787,N_8594,N_8533);
xor U8788 (N_8788,N_8562,N_8545);
and U8789 (N_8789,N_8663,N_8606);
or U8790 (N_8790,N_8680,N_8623);
nor U8791 (N_8791,N_8522,N_8615);
nand U8792 (N_8792,N_8557,N_8683);
and U8793 (N_8793,N_8669,N_8540);
or U8794 (N_8794,N_8622,N_8547);
and U8795 (N_8795,N_8577,N_8573);
nor U8796 (N_8796,N_8518,N_8649);
nor U8797 (N_8797,N_8673,N_8597);
or U8798 (N_8798,N_8648,N_8724);
or U8799 (N_8799,N_8525,N_8638);
nor U8800 (N_8800,N_8705,N_8627);
nand U8801 (N_8801,N_8655,N_8689);
or U8802 (N_8802,N_8668,N_8507);
and U8803 (N_8803,N_8579,N_8538);
nor U8804 (N_8804,N_8618,N_8568);
and U8805 (N_8805,N_8633,N_8708);
xor U8806 (N_8806,N_8532,N_8736);
and U8807 (N_8807,N_8544,N_8730);
and U8808 (N_8808,N_8502,N_8721);
and U8809 (N_8809,N_8735,N_8690);
and U8810 (N_8810,N_8725,N_8727);
xor U8811 (N_8811,N_8583,N_8650);
nand U8812 (N_8812,N_8700,N_8693);
nor U8813 (N_8813,N_8512,N_8684);
xnor U8814 (N_8814,N_8702,N_8514);
and U8815 (N_8815,N_8555,N_8676);
or U8816 (N_8816,N_8524,N_8713);
nor U8817 (N_8817,N_8617,N_8576);
nand U8818 (N_8818,N_8586,N_8609);
nor U8819 (N_8819,N_8529,N_8677);
nand U8820 (N_8820,N_8652,N_8717);
nor U8821 (N_8821,N_8632,N_8667);
and U8822 (N_8822,N_8542,N_8670);
nand U8823 (N_8823,N_8612,N_8614);
xor U8824 (N_8824,N_8636,N_8564);
or U8825 (N_8825,N_8682,N_8674);
nor U8826 (N_8826,N_8551,N_8510);
or U8827 (N_8827,N_8546,N_8696);
xnor U8828 (N_8828,N_8706,N_8699);
nand U8829 (N_8829,N_8745,N_8644);
or U8830 (N_8830,N_8527,N_8539);
xor U8831 (N_8831,N_8578,N_8653);
or U8832 (N_8832,N_8517,N_8712);
or U8833 (N_8833,N_8603,N_8600);
nor U8834 (N_8834,N_8709,N_8504);
xnor U8835 (N_8835,N_8516,N_8588);
nand U8836 (N_8836,N_8584,N_8534);
nand U8837 (N_8837,N_8741,N_8646);
or U8838 (N_8838,N_8575,N_8549);
or U8839 (N_8839,N_8737,N_8686);
or U8840 (N_8840,N_8505,N_8580);
or U8841 (N_8841,N_8608,N_8685);
and U8842 (N_8842,N_8641,N_8744);
nand U8843 (N_8843,N_8613,N_8552);
or U8844 (N_8844,N_8634,N_8590);
xnor U8845 (N_8845,N_8610,N_8624);
nor U8846 (N_8846,N_8581,N_8733);
and U8847 (N_8847,N_8567,N_8561);
nor U8848 (N_8848,N_8698,N_8569);
nand U8849 (N_8849,N_8621,N_8556);
xor U8850 (N_8850,N_8749,N_8558);
nor U8851 (N_8851,N_8715,N_8679);
or U8852 (N_8852,N_8604,N_8701);
and U8853 (N_8853,N_8697,N_8647);
nor U8854 (N_8854,N_8639,N_8687);
or U8855 (N_8855,N_8528,N_8620);
nand U8856 (N_8856,N_8711,N_8731);
and U8857 (N_8857,N_8541,N_8598);
nor U8858 (N_8858,N_8631,N_8511);
and U8859 (N_8859,N_8591,N_8739);
nand U8860 (N_8860,N_8535,N_8662);
xor U8861 (N_8861,N_8703,N_8678);
nor U8862 (N_8862,N_8531,N_8537);
xnor U8863 (N_8863,N_8500,N_8719);
nand U8864 (N_8864,N_8587,N_8565);
xor U8865 (N_8865,N_8595,N_8722);
nor U8866 (N_8866,N_8570,N_8629);
nor U8867 (N_8867,N_8630,N_8643);
xnor U8868 (N_8868,N_8605,N_8651);
nand U8869 (N_8869,N_8602,N_8743);
xor U8870 (N_8870,N_8599,N_8585);
or U8871 (N_8871,N_8704,N_8728);
or U8872 (N_8872,N_8671,N_8716);
and U8873 (N_8873,N_8640,N_8515);
and U8874 (N_8874,N_8710,N_8707);
nor U8875 (N_8875,N_8625,N_8584);
nand U8876 (N_8876,N_8677,N_8639);
xnor U8877 (N_8877,N_8532,N_8668);
and U8878 (N_8878,N_8546,N_8683);
nand U8879 (N_8879,N_8623,N_8722);
nand U8880 (N_8880,N_8532,N_8519);
or U8881 (N_8881,N_8648,N_8560);
or U8882 (N_8882,N_8666,N_8528);
xor U8883 (N_8883,N_8669,N_8666);
nor U8884 (N_8884,N_8535,N_8677);
and U8885 (N_8885,N_8670,N_8621);
or U8886 (N_8886,N_8522,N_8563);
nand U8887 (N_8887,N_8550,N_8749);
nor U8888 (N_8888,N_8650,N_8688);
and U8889 (N_8889,N_8710,N_8660);
xor U8890 (N_8890,N_8672,N_8735);
or U8891 (N_8891,N_8519,N_8593);
or U8892 (N_8892,N_8584,N_8611);
and U8893 (N_8893,N_8727,N_8544);
or U8894 (N_8894,N_8532,N_8650);
nand U8895 (N_8895,N_8698,N_8692);
and U8896 (N_8896,N_8573,N_8743);
or U8897 (N_8897,N_8515,N_8550);
xnor U8898 (N_8898,N_8527,N_8723);
or U8899 (N_8899,N_8618,N_8671);
xnor U8900 (N_8900,N_8538,N_8657);
or U8901 (N_8901,N_8715,N_8578);
and U8902 (N_8902,N_8723,N_8645);
and U8903 (N_8903,N_8646,N_8598);
nand U8904 (N_8904,N_8663,N_8670);
xnor U8905 (N_8905,N_8715,N_8648);
xor U8906 (N_8906,N_8520,N_8680);
nand U8907 (N_8907,N_8671,N_8628);
or U8908 (N_8908,N_8621,N_8674);
xor U8909 (N_8909,N_8613,N_8577);
and U8910 (N_8910,N_8592,N_8507);
nor U8911 (N_8911,N_8658,N_8687);
xnor U8912 (N_8912,N_8729,N_8658);
nand U8913 (N_8913,N_8579,N_8513);
or U8914 (N_8914,N_8548,N_8709);
nand U8915 (N_8915,N_8667,N_8704);
nor U8916 (N_8916,N_8667,N_8739);
nor U8917 (N_8917,N_8667,N_8671);
nand U8918 (N_8918,N_8600,N_8580);
xor U8919 (N_8919,N_8551,N_8558);
and U8920 (N_8920,N_8708,N_8651);
nor U8921 (N_8921,N_8562,N_8691);
nor U8922 (N_8922,N_8565,N_8555);
or U8923 (N_8923,N_8710,N_8583);
or U8924 (N_8924,N_8542,N_8590);
xor U8925 (N_8925,N_8718,N_8621);
xor U8926 (N_8926,N_8713,N_8733);
and U8927 (N_8927,N_8706,N_8657);
nor U8928 (N_8928,N_8732,N_8692);
nand U8929 (N_8929,N_8719,N_8537);
nand U8930 (N_8930,N_8589,N_8510);
and U8931 (N_8931,N_8606,N_8554);
or U8932 (N_8932,N_8563,N_8592);
nand U8933 (N_8933,N_8628,N_8604);
nor U8934 (N_8934,N_8651,N_8719);
nand U8935 (N_8935,N_8517,N_8505);
nor U8936 (N_8936,N_8659,N_8693);
nand U8937 (N_8937,N_8736,N_8675);
xor U8938 (N_8938,N_8653,N_8571);
nand U8939 (N_8939,N_8545,N_8529);
nor U8940 (N_8940,N_8698,N_8736);
and U8941 (N_8941,N_8657,N_8675);
or U8942 (N_8942,N_8723,N_8601);
nor U8943 (N_8943,N_8543,N_8730);
and U8944 (N_8944,N_8696,N_8727);
or U8945 (N_8945,N_8617,N_8600);
and U8946 (N_8946,N_8668,N_8649);
nand U8947 (N_8947,N_8571,N_8735);
and U8948 (N_8948,N_8526,N_8530);
and U8949 (N_8949,N_8739,N_8641);
nor U8950 (N_8950,N_8511,N_8634);
xor U8951 (N_8951,N_8615,N_8562);
nor U8952 (N_8952,N_8687,N_8517);
nand U8953 (N_8953,N_8649,N_8662);
xor U8954 (N_8954,N_8679,N_8555);
and U8955 (N_8955,N_8615,N_8620);
nand U8956 (N_8956,N_8650,N_8640);
nand U8957 (N_8957,N_8644,N_8642);
nand U8958 (N_8958,N_8591,N_8690);
and U8959 (N_8959,N_8703,N_8631);
nor U8960 (N_8960,N_8571,N_8741);
and U8961 (N_8961,N_8702,N_8573);
nand U8962 (N_8962,N_8606,N_8647);
and U8963 (N_8963,N_8559,N_8625);
or U8964 (N_8964,N_8644,N_8681);
or U8965 (N_8965,N_8734,N_8600);
nor U8966 (N_8966,N_8584,N_8515);
and U8967 (N_8967,N_8612,N_8545);
nand U8968 (N_8968,N_8694,N_8564);
nor U8969 (N_8969,N_8674,N_8566);
and U8970 (N_8970,N_8691,N_8636);
nor U8971 (N_8971,N_8691,N_8686);
nand U8972 (N_8972,N_8684,N_8617);
nand U8973 (N_8973,N_8729,N_8521);
nor U8974 (N_8974,N_8546,N_8569);
and U8975 (N_8975,N_8738,N_8588);
or U8976 (N_8976,N_8570,N_8694);
nor U8977 (N_8977,N_8643,N_8590);
and U8978 (N_8978,N_8643,N_8684);
and U8979 (N_8979,N_8644,N_8542);
xnor U8980 (N_8980,N_8746,N_8621);
and U8981 (N_8981,N_8607,N_8685);
and U8982 (N_8982,N_8674,N_8651);
nor U8983 (N_8983,N_8525,N_8532);
or U8984 (N_8984,N_8716,N_8679);
nand U8985 (N_8985,N_8570,N_8659);
nor U8986 (N_8986,N_8533,N_8643);
xor U8987 (N_8987,N_8715,N_8556);
or U8988 (N_8988,N_8732,N_8709);
and U8989 (N_8989,N_8654,N_8663);
xnor U8990 (N_8990,N_8737,N_8610);
nand U8991 (N_8991,N_8540,N_8618);
and U8992 (N_8992,N_8674,N_8696);
nand U8993 (N_8993,N_8518,N_8553);
nand U8994 (N_8994,N_8521,N_8618);
xnor U8995 (N_8995,N_8702,N_8534);
xor U8996 (N_8996,N_8546,N_8667);
or U8997 (N_8997,N_8730,N_8618);
nand U8998 (N_8998,N_8554,N_8549);
nand U8999 (N_8999,N_8685,N_8671);
and U9000 (N_9000,N_8983,N_8769);
and U9001 (N_9001,N_8944,N_8807);
or U9002 (N_9002,N_8949,N_8818);
and U9003 (N_9003,N_8956,N_8923);
xnor U9004 (N_9004,N_8768,N_8839);
nor U9005 (N_9005,N_8950,N_8872);
xor U9006 (N_9006,N_8777,N_8867);
or U9007 (N_9007,N_8780,N_8759);
nor U9008 (N_9008,N_8912,N_8767);
and U9009 (N_9009,N_8922,N_8958);
and U9010 (N_9010,N_8760,N_8813);
xor U9011 (N_9011,N_8786,N_8809);
or U9012 (N_9012,N_8810,N_8954);
and U9013 (N_9013,N_8888,N_8842);
xor U9014 (N_9014,N_8990,N_8996);
nand U9015 (N_9015,N_8795,N_8981);
and U9016 (N_9016,N_8880,N_8801);
and U9017 (N_9017,N_8857,N_8840);
or U9018 (N_9018,N_8982,N_8925);
and U9019 (N_9019,N_8750,N_8911);
xnor U9020 (N_9020,N_8800,N_8783);
and U9021 (N_9021,N_8788,N_8995);
nor U9022 (N_9022,N_8785,N_8793);
xor U9023 (N_9023,N_8751,N_8881);
nor U9024 (N_9024,N_8805,N_8917);
or U9025 (N_9025,N_8782,N_8851);
xnor U9026 (N_9026,N_8992,N_8860);
or U9027 (N_9027,N_8862,N_8919);
xnor U9028 (N_9028,N_8892,N_8808);
xor U9029 (N_9029,N_8987,N_8787);
or U9030 (N_9030,N_8850,N_8963);
or U9031 (N_9031,N_8943,N_8914);
or U9032 (N_9032,N_8988,N_8827);
xnor U9033 (N_9033,N_8927,N_8924);
nand U9034 (N_9034,N_8967,N_8804);
nor U9035 (N_9035,N_8855,N_8965);
nor U9036 (N_9036,N_8883,N_8898);
or U9037 (N_9037,N_8904,N_8823);
and U9038 (N_9038,N_8970,N_8999);
or U9039 (N_9039,N_8941,N_8802);
and U9040 (N_9040,N_8754,N_8779);
xnor U9041 (N_9041,N_8935,N_8928);
xor U9042 (N_9042,N_8994,N_8895);
nor U9043 (N_9043,N_8920,N_8790);
nand U9044 (N_9044,N_8846,N_8910);
nand U9045 (N_9045,N_8775,N_8984);
and U9046 (N_9046,N_8887,N_8953);
nor U9047 (N_9047,N_8766,N_8765);
nand U9048 (N_9048,N_8930,N_8781);
nor U9049 (N_9049,N_8896,N_8908);
nand U9050 (N_9050,N_8833,N_8761);
nand U9051 (N_9051,N_8791,N_8980);
nor U9052 (N_9052,N_8755,N_8957);
and U9053 (N_9053,N_8960,N_8964);
xor U9054 (N_9054,N_8752,N_8939);
nand U9055 (N_9055,N_8838,N_8794);
xor U9056 (N_9056,N_8985,N_8929);
nor U9057 (N_9057,N_8799,N_8962);
nand U9058 (N_9058,N_8797,N_8843);
nor U9059 (N_9059,N_8918,N_8905);
or U9060 (N_9060,N_8770,N_8875);
and U9061 (N_9061,N_8861,N_8758);
nand U9062 (N_9062,N_8945,N_8946);
nand U9063 (N_9063,N_8977,N_8834);
or U9064 (N_9064,N_8913,N_8991);
nor U9065 (N_9065,N_8772,N_8968);
nand U9066 (N_9066,N_8948,N_8829);
nand U9067 (N_9067,N_8899,N_8778);
xnor U9068 (N_9068,N_8792,N_8932);
nor U9069 (N_9069,N_8821,N_8885);
or U9070 (N_9070,N_8940,N_8884);
and U9071 (N_9071,N_8878,N_8877);
xnor U9072 (N_9072,N_8831,N_8921);
and U9073 (N_9073,N_8803,N_8784);
nand U9074 (N_9074,N_8820,N_8952);
nand U9075 (N_9075,N_8825,N_8891);
or U9076 (N_9076,N_8974,N_8856);
nor U9077 (N_9077,N_8816,N_8893);
nor U9078 (N_9078,N_8889,N_8894);
or U9079 (N_9079,N_8973,N_8906);
nor U9080 (N_9080,N_8830,N_8832);
nor U9081 (N_9081,N_8947,N_8835);
or U9082 (N_9082,N_8886,N_8771);
nand U9083 (N_9083,N_8972,N_8763);
nor U9084 (N_9084,N_8931,N_8882);
nand U9085 (N_9085,N_8955,N_8847);
nor U9086 (N_9086,N_8819,N_8853);
or U9087 (N_9087,N_8938,N_8890);
xor U9088 (N_9088,N_8774,N_8773);
xor U9089 (N_9089,N_8969,N_8849);
or U9090 (N_9090,N_8854,N_8826);
nor U9091 (N_9091,N_8874,N_8815);
nor U9092 (N_9092,N_8997,N_8993);
and U9093 (N_9093,N_8812,N_8836);
nand U9094 (N_9094,N_8822,N_8814);
nand U9095 (N_9095,N_8986,N_8789);
or U9096 (N_9096,N_8907,N_8909);
and U9097 (N_9097,N_8897,N_8806);
or U9098 (N_9098,N_8959,N_8870);
and U9099 (N_9099,N_8811,N_8876);
xor U9100 (N_9100,N_8824,N_8976);
nand U9101 (N_9101,N_8844,N_8848);
nand U9102 (N_9102,N_8873,N_8753);
and U9103 (N_9103,N_8762,N_8926);
and U9104 (N_9104,N_8852,N_8915);
or U9105 (N_9105,N_8858,N_8978);
and U9106 (N_9106,N_8859,N_8756);
nand U9107 (N_9107,N_8868,N_8966);
nand U9108 (N_9108,N_8845,N_8879);
and U9109 (N_9109,N_8776,N_8869);
and U9110 (N_9110,N_8934,N_8901);
nand U9111 (N_9111,N_8841,N_8864);
and U9112 (N_9112,N_8817,N_8951);
xnor U9113 (N_9113,N_8961,N_8933);
nor U9114 (N_9114,N_8900,N_8916);
nor U9115 (N_9115,N_8903,N_8998);
and U9116 (N_9116,N_8837,N_8989);
nor U9117 (N_9117,N_8971,N_8937);
xnor U9118 (N_9118,N_8902,N_8979);
and U9119 (N_9119,N_8757,N_8975);
and U9120 (N_9120,N_8866,N_8796);
nand U9121 (N_9121,N_8871,N_8798);
nand U9122 (N_9122,N_8764,N_8828);
or U9123 (N_9123,N_8936,N_8863);
nand U9124 (N_9124,N_8942,N_8865);
and U9125 (N_9125,N_8893,N_8814);
or U9126 (N_9126,N_8943,N_8775);
xor U9127 (N_9127,N_8785,N_8999);
nor U9128 (N_9128,N_8993,N_8777);
nand U9129 (N_9129,N_8801,N_8860);
xnor U9130 (N_9130,N_8826,N_8802);
or U9131 (N_9131,N_8843,N_8799);
nor U9132 (N_9132,N_8772,N_8851);
and U9133 (N_9133,N_8820,N_8982);
and U9134 (N_9134,N_8843,N_8825);
or U9135 (N_9135,N_8928,N_8978);
nand U9136 (N_9136,N_8956,N_8915);
nand U9137 (N_9137,N_8958,N_8855);
or U9138 (N_9138,N_8933,N_8981);
xnor U9139 (N_9139,N_8810,N_8796);
and U9140 (N_9140,N_8966,N_8846);
nor U9141 (N_9141,N_8842,N_8900);
or U9142 (N_9142,N_8866,N_8893);
nor U9143 (N_9143,N_8843,N_8769);
and U9144 (N_9144,N_8898,N_8962);
nor U9145 (N_9145,N_8857,N_8987);
nor U9146 (N_9146,N_8769,N_8857);
and U9147 (N_9147,N_8904,N_8869);
nand U9148 (N_9148,N_8987,N_8869);
xnor U9149 (N_9149,N_8888,N_8795);
nor U9150 (N_9150,N_8844,N_8983);
or U9151 (N_9151,N_8972,N_8939);
nand U9152 (N_9152,N_8783,N_8999);
nor U9153 (N_9153,N_8812,N_8879);
and U9154 (N_9154,N_8802,N_8831);
and U9155 (N_9155,N_8784,N_8852);
or U9156 (N_9156,N_8950,N_8874);
nor U9157 (N_9157,N_8762,N_8855);
nand U9158 (N_9158,N_8846,N_8760);
nor U9159 (N_9159,N_8951,N_8762);
xor U9160 (N_9160,N_8756,N_8813);
nand U9161 (N_9161,N_8911,N_8994);
and U9162 (N_9162,N_8851,N_8872);
or U9163 (N_9163,N_8773,N_8958);
xnor U9164 (N_9164,N_8815,N_8993);
and U9165 (N_9165,N_8972,N_8988);
and U9166 (N_9166,N_8949,N_8908);
or U9167 (N_9167,N_8963,N_8881);
nand U9168 (N_9168,N_8830,N_8946);
xnor U9169 (N_9169,N_8906,N_8797);
xnor U9170 (N_9170,N_8910,N_8933);
or U9171 (N_9171,N_8751,N_8780);
and U9172 (N_9172,N_8958,N_8856);
xor U9173 (N_9173,N_8869,N_8977);
nor U9174 (N_9174,N_8932,N_8869);
or U9175 (N_9175,N_8802,N_8780);
nand U9176 (N_9176,N_8925,N_8864);
xnor U9177 (N_9177,N_8965,N_8778);
nor U9178 (N_9178,N_8754,N_8859);
xor U9179 (N_9179,N_8854,N_8859);
nor U9180 (N_9180,N_8880,N_8881);
and U9181 (N_9181,N_8771,N_8815);
nor U9182 (N_9182,N_8970,N_8803);
xor U9183 (N_9183,N_8841,N_8876);
nor U9184 (N_9184,N_8757,N_8913);
nand U9185 (N_9185,N_8777,N_8792);
nor U9186 (N_9186,N_8845,N_8818);
and U9187 (N_9187,N_8762,N_8756);
or U9188 (N_9188,N_8932,N_8789);
xor U9189 (N_9189,N_8757,N_8825);
and U9190 (N_9190,N_8768,N_8908);
xnor U9191 (N_9191,N_8799,N_8906);
xor U9192 (N_9192,N_8863,N_8805);
nor U9193 (N_9193,N_8923,N_8809);
nor U9194 (N_9194,N_8773,N_8930);
and U9195 (N_9195,N_8885,N_8759);
nand U9196 (N_9196,N_8800,N_8770);
and U9197 (N_9197,N_8926,N_8903);
nor U9198 (N_9198,N_8902,N_8898);
or U9199 (N_9199,N_8957,N_8971);
and U9200 (N_9200,N_8798,N_8982);
xor U9201 (N_9201,N_8762,N_8966);
or U9202 (N_9202,N_8830,N_8819);
xor U9203 (N_9203,N_8910,N_8875);
and U9204 (N_9204,N_8891,N_8841);
nor U9205 (N_9205,N_8797,N_8800);
nor U9206 (N_9206,N_8917,N_8904);
xor U9207 (N_9207,N_8798,N_8931);
or U9208 (N_9208,N_8861,N_8815);
or U9209 (N_9209,N_8978,N_8851);
and U9210 (N_9210,N_8817,N_8757);
or U9211 (N_9211,N_8989,N_8948);
xnor U9212 (N_9212,N_8837,N_8993);
or U9213 (N_9213,N_8765,N_8964);
nand U9214 (N_9214,N_8928,N_8949);
nor U9215 (N_9215,N_8941,N_8758);
xnor U9216 (N_9216,N_8992,N_8949);
xor U9217 (N_9217,N_8982,N_8879);
nand U9218 (N_9218,N_8982,N_8906);
or U9219 (N_9219,N_8970,N_8790);
xnor U9220 (N_9220,N_8865,N_8856);
or U9221 (N_9221,N_8995,N_8888);
nor U9222 (N_9222,N_8943,N_8913);
or U9223 (N_9223,N_8782,N_8911);
or U9224 (N_9224,N_8992,N_8921);
or U9225 (N_9225,N_8840,N_8795);
nand U9226 (N_9226,N_8980,N_8960);
xnor U9227 (N_9227,N_8954,N_8793);
and U9228 (N_9228,N_8768,N_8919);
nor U9229 (N_9229,N_8769,N_8761);
xor U9230 (N_9230,N_8914,N_8981);
or U9231 (N_9231,N_8903,N_8929);
xnor U9232 (N_9232,N_8843,N_8946);
and U9233 (N_9233,N_8813,N_8750);
or U9234 (N_9234,N_8835,N_8857);
nand U9235 (N_9235,N_8856,N_8828);
nor U9236 (N_9236,N_8821,N_8819);
or U9237 (N_9237,N_8769,N_8874);
or U9238 (N_9238,N_8802,N_8926);
nor U9239 (N_9239,N_8774,N_8972);
or U9240 (N_9240,N_8799,N_8805);
nor U9241 (N_9241,N_8980,N_8790);
and U9242 (N_9242,N_8860,N_8966);
nand U9243 (N_9243,N_8863,N_8760);
or U9244 (N_9244,N_8899,N_8866);
nor U9245 (N_9245,N_8893,N_8943);
xor U9246 (N_9246,N_8759,N_8917);
nand U9247 (N_9247,N_8872,N_8917);
xor U9248 (N_9248,N_8850,N_8973);
and U9249 (N_9249,N_8988,N_8791);
xor U9250 (N_9250,N_9213,N_9000);
xnor U9251 (N_9251,N_9092,N_9078);
or U9252 (N_9252,N_9105,N_9192);
xnor U9253 (N_9253,N_9153,N_9248);
nor U9254 (N_9254,N_9208,N_9154);
and U9255 (N_9255,N_9028,N_9061);
and U9256 (N_9256,N_9062,N_9172);
and U9257 (N_9257,N_9225,N_9064);
nand U9258 (N_9258,N_9017,N_9196);
or U9259 (N_9259,N_9195,N_9115);
or U9260 (N_9260,N_9226,N_9119);
nand U9261 (N_9261,N_9096,N_9100);
nor U9262 (N_9262,N_9194,N_9025);
or U9263 (N_9263,N_9075,N_9109);
nand U9264 (N_9264,N_9134,N_9233);
and U9265 (N_9265,N_9131,N_9110);
nor U9266 (N_9266,N_9050,N_9164);
nand U9267 (N_9267,N_9007,N_9161);
or U9268 (N_9268,N_9139,N_9016);
xnor U9269 (N_9269,N_9051,N_9166);
nor U9270 (N_9270,N_9169,N_9060);
or U9271 (N_9271,N_9173,N_9106);
or U9272 (N_9272,N_9136,N_9066);
xnor U9273 (N_9273,N_9206,N_9217);
xnor U9274 (N_9274,N_9155,N_9053);
or U9275 (N_9275,N_9239,N_9203);
nor U9276 (N_9276,N_9093,N_9207);
xor U9277 (N_9277,N_9212,N_9118);
xnor U9278 (N_9278,N_9104,N_9114);
nor U9279 (N_9279,N_9214,N_9210);
and U9280 (N_9280,N_9170,N_9179);
and U9281 (N_9281,N_9032,N_9009);
nand U9282 (N_9282,N_9188,N_9037);
and U9283 (N_9283,N_9163,N_9123);
and U9284 (N_9284,N_9059,N_9073);
or U9285 (N_9285,N_9090,N_9211);
nand U9286 (N_9286,N_9095,N_9112);
and U9287 (N_9287,N_9113,N_9247);
nor U9288 (N_9288,N_9005,N_9027);
and U9289 (N_9289,N_9116,N_9083);
xnor U9290 (N_9290,N_9237,N_9184);
nand U9291 (N_9291,N_9038,N_9145);
or U9292 (N_9292,N_9220,N_9071);
or U9293 (N_9293,N_9130,N_9117);
nand U9294 (N_9294,N_9080,N_9129);
or U9295 (N_9295,N_9156,N_9224);
and U9296 (N_9296,N_9185,N_9209);
or U9297 (N_9297,N_9054,N_9168);
nor U9298 (N_9298,N_9198,N_9019);
nor U9299 (N_9299,N_9193,N_9033);
and U9300 (N_9300,N_9199,N_9178);
or U9301 (N_9301,N_9036,N_9165);
nand U9302 (N_9302,N_9200,N_9243);
nand U9303 (N_9303,N_9121,N_9102);
and U9304 (N_9304,N_9138,N_9085);
nand U9305 (N_9305,N_9079,N_9055);
nand U9306 (N_9306,N_9142,N_9159);
or U9307 (N_9307,N_9152,N_9058);
nand U9308 (N_9308,N_9035,N_9187);
xor U9309 (N_9309,N_9158,N_9120);
and U9310 (N_9310,N_9218,N_9204);
and U9311 (N_9311,N_9230,N_9127);
or U9312 (N_9312,N_9070,N_9146);
nand U9313 (N_9313,N_9081,N_9189);
nand U9314 (N_9314,N_9018,N_9183);
nor U9315 (N_9315,N_9008,N_9175);
and U9316 (N_9316,N_9103,N_9011);
and U9317 (N_9317,N_9176,N_9144);
or U9318 (N_9318,N_9098,N_9021);
and U9319 (N_9319,N_9240,N_9219);
xnor U9320 (N_9320,N_9097,N_9167);
xnor U9321 (N_9321,N_9235,N_9141);
or U9322 (N_9322,N_9034,N_9132);
nor U9323 (N_9323,N_9125,N_9012);
or U9324 (N_9324,N_9186,N_9133);
nand U9325 (N_9325,N_9040,N_9014);
or U9326 (N_9326,N_9190,N_9249);
nand U9327 (N_9327,N_9020,N_9089);
and U9328 (N_9328,N_9088,N_9216);
xor U9329 (N_9329,N_9108,N_9221);
or U9330 (N_9330,N_9010,N_9047);
nor U9331 (N_9331,N_9162,N_9222);
nor U9332 (N_9332,N_9041,N_9236);
nor U9333 (N_9333,N_9234,N_9024);
nor U9334 (N_9334,N_9245,N_9094);
xor U9335 (N_9335,N_9191,N_9084);
or U9336 (N_9336,N_9231,N_9140);
nand U9337 (N_9337,N_9148,N_9023);
and U9338 (N_9338,N_9029,N_9002);
and U9339 (N_9339,N_9241,N_9077);
and U9340 (N_9340,N_9147,N_9128);
nor U9341 (N_9341,N_9150,N_9045);
xor U9342 (N_9342,N_9068,N_9074);
nand U9343 (N_9343,N_9101,N_9030);
nand U9344 (N_9344,N_9151,N_9202);
or U9345 (N_9345,N_9087,N_9067);
and U9346 (N_9346,N_9076,N_9082);
xor U9347 (N_9347,N_9232,N_9022);
or U9348 (N_9348,N_9143,N_9039);
xnor U9349 (N_9349,N_9065,N_9174);
or U9350 (N_9350,N_9244,N_9046);
nand U9351 (N_9351,N_9063,N_9056);
nand U9352 (N_9352,N_9099,N_9135);
xnor U9353 (N_9353,N_9026,N_9171);
nand U9354 (N_9354,N_9003,N_9013);
nand U9355 (N_9355,N_9107,N_9057);
nand U9356 (N_9356,N_9048,N_9052);
nor U9357 (N_9357,N_9086,N_9006);
or U9358 (N_9358,N_9205,N_9091);
nor U9359 (N_9359,N_9160,N_9197);
nand U9360 (N_9360,N_9238,N_9215);
nor U9361 (N_9361,N_9069,N_9228);
and U9362 (N_9362,N_9044,N_9031);
nor U9363 (N_9363,N_9015,N_9111);
xnor U9364 (N_9364,N_9124,N_9242);
and U9365 (N_9365,N_9004,N_9072);
and U9366 (N_9366,N_9137,N_9122);
nand U9367 (N_9367,N_9227,N_9043);
nor U9368 (N_9368,N_9201,N_9177);
xnor U9369 (N_9369,N_9180,N_9001);
nor U9370 (N_9370,N_9246,N_9126);
and U9371 (N_9371,N_9042,N_9149);
and U9372 (N_9372,N_9157,N_9229);
xnor U9373 (N_9373,N_9182,N_9181);
nor U9374 (N_9374,N_9049,N_9223);
or U9375 (N_9375,N_9018,N_9235);
or U9376 (N_9376,N_9207,N_9024);
and U9377 (N_9377,N_9163,N_9166);
and U9378 (N_9378,N_9214,N_9021);
and U9379 (N_9379,N_9245,N_9040);
xor U9380 (N_9380,N_9059,N_9144);
and U9381 (N_9381,N_9204,N_9116);
nand U9382 (N_9382,N_9009,N_9080);
nor U9383 (N_9383,N_9175,N_9037);
nor U9384 (N_9384,N_9082,N_9179);
nor U9385 (N_9385,N_9146,N_9245);
or U9386 (N_9386,N_9059,N_9180);
nand U9387 (N_9387,N_9066,N_9192);
xnor U9388 (N_9388,N_9177,N_9188);
and U9389 (N_9389,N_9219,N_9168);
nor U9390 (N_9390,N_9125,N_9164);
and U9391 (N_9391,N_9215,N_9166);
xor U9392 (N_9392,N_9188,N_9089);
nand U9393 (N_9393,N_9075,N_9091);
xnor U9394 (N_9394,N_9243,N_9122);
nor U9395 (N_9395,N_9245,N_9219);
or U9396 (N_9396,N_9123,N_9227);
nor U9397 (N_9397,N_9155,N_9236);
xor U9398 (N_9398,N_9015,N_9227);
xnor U9399 (N_9399,N_9097,N_9226);
or U9400 (N_9400,N_9228,N_9094);
or U9401 (N_9401,N_9089,N_9073);
and U9402 (N_9402,N_9235,N_9224);
or U9403 (N_9403,N_9245,N_9226);
and U9404 (N_9404,N_9162,N_9233);
nand U9405 (N_9405,N_9005,N_9163);
and U9406 (N_9406,N_9150,N_9051);
or U9407 (N_9407,N_9215,N_9059);
xor U9408 (N_9408,N_9073,N_9102);
and U9409 (N_9409,N_9105,N_9138);
nand U9410 (N_9410,N_9222,N_9232);
nand U9411 (N_9411,N_9073,N_9123);
or U9412 (N_9412,N_9103,N_9244);
or U9413 (N_9413,N_9205,N_9212);
nand U9414 (N_9414,N_9066,N_9196);
or U9415 (N_9415,N_9138,N_9214);
nor U9416 (N_9416,N_9189,N_9002);
xor U9417 (N_9417,N_9220,N_9078);
or U9418 (N_9418,N_9092,N_9145);
or U9419 (N_9419,N_9169,N_9053);
nor U9420 (N_9420,N_9012,N_9185);
or U9421 (N_9421,N_9039,N_9207);
nand U9422 (N_9422,N_9150,N_9064);
nor U9423 (N_9423,N_9002,N_9077);
nand U9424 (N_9424,N_9087,N_9197);
nor U9425 (N_9425,N_9109,N_9082);
nor U9426 (N_9426,N_9100,N_9119);
nor U9427 (N_9427,N_9084,N_9183);
xnor U9428 (N_9428,N_9239,N_9063);
nor U9429 (N_9429,N_9178,N_9233);
or U9430 (N_9430,N_9062,N_9039);
or U9431 (N_9431,N_9167,N_9111);
or U9432 (N_9432,N_9127,N_9006);
nor U9433 (N_9433,N_9032,N_9173);
xnor U9434 (N_9434,N_9185,N_9221);
nor U9435 (N_9435,N_9115,N_9176);
nand U9436 (N_9436,N_9085,N_9233);
and U9437 (N_9437,N_9182,N_9012);
nor U9438 (N_9438,N_9155,N_9054);
or U9439 (N_9439,N_9220,N_9190);
nand U9440 (N_9440,N_9010,N_9046);
nand U9441 (N_9441,N_9177,N_9079);
or U9442 (N_9442,N_9201,N_9068);
nor U9443 (N_9443,N_9162,N_9163);
nor U9444 (N_9444,N_9180,N_9023);
and U9445 (N_9445,N_9080,N_9065);
and U9446 (N_9446,N_9239,N_9044);
xnor U9447 (N_9447,N_9079,N_9160);
and U9448 (N_9448,N_9199,N_9172);
nand U9449 (N_9449,N_9072,N_9049);
nor U9450 (N_9450,N_9110,N_9042);
and U9451 (N_9451,N_9114,N_9087);
or U9452 (N_9452,N_9021,N_9238);
xnor U9453 (N_9453,N_9018,N_9186);
xor U9454 (N_9454,N_9111,N_9054);
xnor U9455 (N_9455,N_9204,N_9232);
or U9456 (N_9456,N_9229,N_9028);
and U9457 (N_9457,N_9143,N_9092);
xnor U9458 (N_9458,N_9202,N_9170);
xnor U9459 (N_9459,N_9169,N_9164);
xnor U9460 (N_9460,N_9169,N_9055);
and U9461 (N_9461,N_9247,N_9181);
and U9462 (N_9462,N_9116,N_9131);
nand U9463 (N_9463,N_9145,N_9048);
nor U9464 (N_9464,N_9024,N_9030);
xnor U9465 (N_9465,N_9200,N_9233);
or U9466 (N_9466,N_9067,N_9153);
nor U9467 (N_9467,N_9117,N_9137);
or U9468 (N_9468,N_9141,N_9077);
and U9469 (N_9469,N_9120,N_9008);
or U9470 (N_9470,N_9245,N_9182);
and U9471 (N_9471,N_9196,N_9170);
xnor U9472 (N_9472,N_9185,N_9237);
and U9473 (N_9473,N_9132,N_9218);
nor U9474 (N_9474,N_9139,N_9239);
nand U9475 (N_9475,N_9183,N_9158);
and U9476 (N_9476,N_9087,N_9110);
and U9477 (N_9477,N_9046,N_9111);
nand U9478 (N_9478,N_9095,N_9074);
or U9479 (N_9479,N_9237,N_9212);
or U9480 (N_9480,N_9160,N_9238);
nand U9481 (N_9481,N_9056,N_9050);
nor U9482 (N_9482,N_9176,N_9073);
nand U9483 (N_9483,N_9180,N_9214);
xnor U9484 (N_9484,N_9062,N_9099);
and U9485 (N_9485,N_9179,N_9143);
or U9486 (N_9486,N_9178,N_9066);
xor U9487 (N_9487,N_9219,N_9204);
xnor U9488 (N_9488,N_9202,N_9023);
and U9489 (N_9489,N_9107,N_9202);
nor U9490 (N_9490,N_9237,N_9151);
nor U9491 (N_9491,N_9110,N_9199);
and U9492 (N_9492,N_9204,N_9214);
xor U9493 (N_9493,N_9078,N_9038);
xnor U9494 (N_9494,N_9126,N_9161);
or U9495 (N_9495,N_9106,N_9118);
xnor U9496 (N_9496,N_9170,N_9017);
nor U9497 (N_9497,N_9097,N_9098);
nor U9498 (N_9498,N_9035,N_9186);
nor U9499 (N_9499,N_9142,N_9091);
nand U9500 (N_9500,N_9364,N_9472);
nor U9501 (N_9501,N_9256,N_9488);
xor U9502 (N_9502,N_9459,N_9419);
or U9503 (N_9503,N_9464,N_9293);
and U9504 (N_9504,N_9453,N_9455);
or U9505 (N_9505,N_9297,N_9397);
xor U9506 (N_9506,N_9416,N_9351);
nand U9507 (N_9507,N_9435,N_9374);
or U9508 (N_9508,N_9285,N_9302);
nor U9509 (N_9509,N_9360,N_9252);
and U9510 (N_9510,N_9375,N_9441);
nor U9511 (N_9511,N_9279,N_9482);
xnor U9512 (N_9512,N_9429,N_9295);
or U9513 (N_9513,N_9440,N_9315);
nor U9514 (N_9514,N_9267,N_9340);
nor U9515 (N_9515,N_9296,N_9257);
or U9516 (N_9516,N_9475,N_9437);
nor U9517 (N_9517,N_9373,N_9409);
nor U9518 (N_9518,N_9423,N_9408);
nand U9519 (N_9519,N_9269,N_9286);
nor U9520 (N_9520,N_9299,N_9304);
and U9521 (N_9521,N_9449,N_9291);
nor U9522 (N_9522,N_9460,N_9294);
or U9523 (N_9523,N_9354,N_9319);
and U9524 (N_9524,N_9368,N_9344);
xnor U9525 (N_9525,N_9276,N_9413);
or U9526 (N_9526,N_9468,N_9260);
xor U9527 (N_9527,N_9425,N_9405);
xnor U9528 (N_9528,N_9311,N_9384);
xor U9529 (N_9529,N_9390,N_9357);
and U9530 (N_9530,N_9277,N_9387);
nand U9531 (N_9531,N_9376,N_9301);
nand U9532 (N_9532,N_9446,N_9289);
or U9533 (N_9533,N_9379,N_9424);
xnor U9534 (N_9534,N_9473,N_9402);
or U9535 (N_9535,N_9489,N_9485);
nand U9536 (N_9536,N_9454,N_9303);
and U9537 (N_9537,N_9307,N_9491);
and U9538 (N_9538,N_9263,N_9271);
and U9539 (N_9539,N_9268,N_9395);
xor U9540 (N_9540,N_9382,N_9380);
and U9541 (N_9541,N_9461,N_9363);
nand U9542 (N_9542,N_9439,N_9262);
or U9543 (N_9543,N_9420,N_9261);
nor U9544 (N_9544,N_9258,N_9280);
xor U9545 (N_9545,N_9457,N_9329);
or U9546 (N_9546,N_9490,N_9350);
xnor U9547 (N_9547,N_9392,N_9284);
nor U9548 (N_9548,N_9345,N_9412);
nor U9549 (N_9549,N_9452,N_9337);
and U9550 (N_9550,N_9332,N_9254);
nor U9551 (N_9551,N_9442,N_9481);
and U9552 (N_9552,N_9275,N_9386);
xor U9553 (N_9553,N_9391,N_9253);
or U9554 (N_9554,N_9436,N_9445);
or U9555 (N_9555,N_9336,N_9342);
nor U9556 (N_9556,N_9317,N_9410);
xnor U9557 (N_9557,N_9355,N_9444);
nor U9558 (N_9558,N_9343,N_9400);
or U9559 (N_9559,N_9306,N_9465);
nor U9560 (N_9560,N_9333,N_9298);
or U9561 (N_9561,N_9270,N_9484);
xnor U9562 (N_9562,N_9292,N_9418);
or U9563 (N_9563,N_9347,N_9300);
and U9564 (N_9564,N_9366,N_9407);
and U9565 (N_9565,N_9266,N_9448);
xor U9566 (N_9566,N_9398,N_9492);
nand U9567 (N_9567,N_9471,N_9281);
nand U9568 (N_9568,N_9352,N_9338);
and U9569 (N_9569,N_9255,N_9499);
xnor U9570 (N_9570,N_9341,N_9381);
xor U9571 (N_9571,N_9426,N_9288);
nand U9572 (N_9572,N_9378,N_9399);
or U9573 (N_9573,N_9493,N_9325);
nor U9574 (N_9574,N_9272,N_9334);
nand U9575 (N_9575,N_9483,N_9335);
or U9576 (N_9576,N_9434,N_9316);
and U9577 (N_9577,N_9458,N_9327);
nor U9578 (N_9578,N_9406,N_9273);
or U9579 (N_9579,N_9466,N_9312);
nand U9580 (N_9580,N_9462,N_9328);
nor U9581 (N_9581,N_9428,N_9290);
and U9582 (N_9582,N_9496,N_9305);
or U9583 (N_9583,N_9371,N_9264);
and U9584 (N_9584,N_9498,N_9411);
or U9585 (N_9585,N_9330,N_9438);
or U9586 (N_9586,N_9393,N_9287);
nor U9587 (N_9587,N_9283,N_9323);
nor U9588 (N_9588,N_9365,N_9361);
nor U9589 (N_9589,N_9470,N_9433);
or U9590 (N_9590,N_9321,N_9309);
and U9591 (N_9591,N_9396,N_9478);
and U9592 (N_9592,N_9310,N_9414);
nor U9593 (N_9593,N_9486,N_9372);
nor U9594 (N_9594,N_9265,N_9259);
or U9595 (N_9595,N_9487,N_9404);
xnor U9596 (N_9596,N_9403,N_9450);
and U9597 (N_9597,N_9313,N_9431);
nand U9598 (N_9598,N_9251,N_9417);
nand U9599 (N_9599,N_9421,N_9349);
nor U9600 (N_9600,N_9427,N_9389);
and U9601 (N_9601,N_9331,N_9274);
nor U9602 (N_9602,N_9385,N_9476);
xnor U9603 (N_9603,N_9477,N_9447);
and U9604 (N_9604,N_9339,N_9497);
xnor U9605 (N_9605,N_9479,N_9278);
and U9606 (N_9606,N_9443,N_9358);
nor U9607 (N_9607,N_9432,N_9324);
nor U9608 (N_9608,N_9370,N_9430);
nand U9609 (N_9609,N_9422,N_9467);
or U9610 (N_9610,N_9367,N_9415);
nand U9611 (N_9611,N_9353,N_9282);
nand U9612 (N_9612,N_9394,N_9348);
nor U9613 (N_9613,N_9474,N_9494);
xor U9614 (N_9614,N_9346,N_9362);
nand U9615 (N_9615,N_9469,N_9456);
and U9616 (N_9616,N_9495,N_9359);
xnor U9617 (N_9617,N_9388,N_9320);
and U9618 (N_9618,N_9377,N_9308);
nor U9619 (N_9619,N_9383,N_9451);
nand U9620 (N_9620,N_9463,N_9322);
and U9621 (N_9621,N_9369,N_9314);
and U9622 (N_9622,N_9326,N_9401);
xnor U9623 (N_9623,N_9250,N_9480);
or U9624 (N_9624,N_9356,N_9318);
and U9625 (N_9625,N_9320,N_9281);
or U9626 (N_9626,N_9353,N_9446);
nand U9627 (N_9627,N_9391,N_9322);
or U9628 (N_9628,N_9332,N_9309);
xor U9629 (N_9629,N_9292,N_9410);
xor U9630 (N_9630,N_9368,N_9493);
xor U9631 (N_9631,N_9343,N_9305);
and U9632 (N_9632,N_9363,N_9488);
or U9633 (N_9633,N_9406,N_9476);
and U9634 (N_9634,N_9267,N_9297);
and U9635 (N_9635,N_9259,N_9281);
xor U9636 (N_9636,N_9353,N_9283);
xor U9637 (N_9637,N_9335,N_9267);
or U9638 (N_9638,N_9327,N_9280);
xor U9639 (N_9639,N_9299,N_9442);
nor U9640 (N_9640,N_9445,N_9312);
nand U9641 (N_9641,N_9432,N_9319);
and U9642 (N_9642,N_9344,N_9260);
and U9643 (N_9643,N_9477,N_9432);
and U9644 (N_9644,N_9364,N_9496);
or U9645 (N_9645,N_9322,N_9332);
and U9646 (N_9646,N_9428,N_9496);
nor U9647 (N_9647,N_9498,N_9353);
or U9648 (N_9648,N_9441,N_9279);
nand U9649 (N_9649,N_9430,N_9424);
nand U9650 (N_9650,N_9420,N_9412);
and U9651 (N_9651,N_9273,N_9350);
or U9652 (N_9652,N_9350,N_9254);
nand U9653 (N_9653,N_9455,N_9252);
nand U9654 (N_9654,N_9297,N_9340);
or U9655 (N_9655,N_9252,N_9414);
and U9656 (N_9656,N_9321,N_9320);
or U9657 (N_9657,N_9267,N_9461);
xnor U9658 (N_9658,N_9477,N_9278);
nand U9659 (N_9659,N_9305,N_9361);
nor U9660 (N_9660,N_9406,N_9465);
nand U9661 (N_9661,N_9403,N_9319);
and U9662 (N_9662,N_9362,N_9364);
or U9663 (N_9663,N_9470,N_9442);
and U9664 (N_9664,N_9438,N_9396);
nor U9665 (N_9665,N_9342,N_9433);
xnor U9666 (N_9666,N_9275,N_9277);
xor U9667 (N_9667,N_9297,N_9453);
nand U9668 (N_9668,N_9320,N_9429);
xor U9669 (N_9669,N_9333,N_9334);
and U9670 (N_9670,N_9383,N_9467);
or U9671 (N_9671,N_9378,N_9481);
nand U9672 (N_9672,N_9362,N_9402);
or U9673 (N_9673,N_9334,N_9297);
nor U9674 (N_9674,N_9463,N_9383);
nand U9675 (N_9675,N_9341,N_9347);
nor U9676 (N_9676,N_9440,N_9345);
xnor U9677 (N_9677,N_9463,N_9350);
and U9678 (N_9678,N_9281,N_9274);
or U9679 (N_9679,N_9412,N_9343);
xor U9680 (N_9680,N_9482,N_9309);
nand U9681 (N_9681,N_9399,N_9250);
and U9682 (N_9682,N_9351,N_9461);
nand U9683 (N_9683,N_9392,N_9358);
nand U9684 (N_9684,N_9383,N_9398);
xnor U9685 (N_9685,N_9459,N_9343);
and U9686 (N_9686,N_9450,N_9257);
or U9687 (N_9687,N_9480,N_9432);
or U9688 (N_9688,N_9339,N_9444);
and U9689 (N_9689,N_9429,N_9416);
nand U9690 (N_9690,N_9432,N_9277);
or U9691 (N_9691,N_9272,N_9256);
nand U9692 (N_9692,N_9407,N_9295);
or U9693 (N_9693,N_9282,N_9478);
and U9694 (N_9694,N_9460,N_9448);
and U9695 (N_9695,N_9423,N_9472);
nand U9696 (N_9696,N_9448,N_9366);
nor U9697 (N_9697,N_9298,N_9348);
nand U9698 (N_9698,N_9474,N_9451);
and U9699 (N_9699,N_9265,N_9434);
xnor U9700 (N_9700,N_9339,N_9416);
and U9701 (N_9701,N_9324,N_9329);
nor U9702 (N_9702,N_9415,N_9498);
nor U9703 (N_9703,N_9354,N_9295);
and U9704 (N_9704,N_9369,N_9265);
xor U9705 (N_9705,N_9269,N_9338);
nand U9706 (N_9706,N_9307,N_9457);
xnor U9707 (N_9707,N_9478,N_9462);
nand U9708 (N_9708,N_9324,N_9304);
nor U9709 (N_9709,N_9306,N_9493);
xnor U9710 (N_9710,N_9276,N_9363);
nand U9711 (N_9711,N_9415,N_9478);
nand U9712 (N_9712,N_9430,N_9497);
xor U9713 (N_9713,N_9436,N_9318);
or U9714 (N_9714,N_9430,N_9321);
xor U9715 (N_9715,N_9498,N_9369);
and U9716 (N_9716,N_9433,N_9372);
xnor U9717 (N_9717,N_9415,N_9491);
nor U9718 (N_9718,N_9443,N_9364);
nand U9719 (N_9719,N_9293,N_9409);
nand U9720 (N_9720,N_9342,N_9386);
nand U9721 (N_9721,N_9375,N_9341);
or U9722 (N_9722,N_9341,N_9471);
or U9723 (N_9723,N_9443,N_9254);
and U9724 (N_9724,N_9369,N_9358);
nand U9725 (N_9725,N_9362,N_9394);
nand U9726 (N_9726,N_9391,N_9274);
xor U9727 (N_9727,N_9429,N_9297);
nor U9728 (N_9728,N_9265,N_9430);
xor U9729 (N_9729,N_9491,N_9355);
xor U9730 (N_9730,N_9471,N_9492);
xnor U9731 (N_9731,N_9292,N_9330);
xor U9732 (N_9732,N_9283,N_9394);
nand U9733 (N_9733,N_9306,N_9492);
nand U9734 (N_9734,N_9356,N_9363);
and U9735 (N_9735,N_9479,N_9424);
or U9736 (N_9736,N_9369,N_9334);
or U9737 (N_9737,N_9316,N_9400);
xnor U9738 (N_9738,N_9467,N_9386);
nand U9739 (N_9739,N_9352,N_9335);
nand U9740 (N_9740,N_9440,N_9308);
and U9741 (N_9741,N_9394,N_9250);
nand U9742 (N_9742,N_9459,N_9482);
or U9743 (N_9743,N_9415,N_9406);
or U9744 (N_9744,N_9293,N_9259);
xnor U9745 (N_9745,N_9340,N_9271);
nor U9746 (N_9746,N_9315,N_9346);
xnor U9747 (N_9747,N_9269,N_9444);
and U9748 (N_9748,N_9414,N_9330);
nor U9749 (N_9749,N_9397,N_9372);
nor U9750 (N_9750,N_9670,N_9692);
and U9751 (N_9751,N_9699,N_9620);
nand U9752 (N_9752,N_9700,N_9702);
nand U9753 (N_9753,N_9701,N_9735);
nor U9754 (N_9754,N_9551,N_9707);
nand U9755 (N_9755,N_9723,N_9527);
nor U9756 (N_9756,N_9681,N_9673);
and U9757 (N_9757,N_9609,N_9617);
or U9758 (N_9758,N_9598,N_9561);
nand U9759 (N_9759,N_9520,N_9526);
nor U9760 (N_9760,N_9649,N_9662);
and U9761 (N_9761,N_9508,N_9656);
nand U9762 (N_9762,N_9563,N_9559);
xnor U9763 (N_9763,N_9522,N_9680);
nor U9764 (N_9764,N_9713,N_9646);
nand U9765 (N_9765,N_9556,N_9507);
nor U9766 (N_9766,N_9584,N_9577);
or U9767 (N_9767,N_9570,N_9585);
nor U9768 (N_9768,N_9568,N_9652);
xnor U9769 (N_9769,N_9572,N_9709);
or U9770 (N_9770,N_9521,N_9573);
nor U9771 (N_9771,N_9612,N_9583);
or U9772 (N_9772,N_9546,N_9616);
and U9773 (N_9773,N_9606,N_9574);
and U9774 (N_9774,N_9621,N_9553);
nand U9775 (N_9775,N_9655,N_9630);
xnor U9776 (N_9776,N_9664,N_9675);
xnor U9777 (N_9777,N_9710,N_9679);
xor U9778 (N_9778,N_9727,N_9725);
xnor U9779 (N_9779,N_9562,N_9684);
nand U9780 (N_9780,N_9566,N_9668);
nor U9781 (N_9781,N_9537,N_9637);
and U9782 (N_9782,N_9635,N_9629);
and U9783 (N_9783,N_9558,N_9678);
xnor U9784 (N_9784,N_9535,N_9665);
or U9785 (N_9785,N_9571,N_9627);
or U9786 (N_9786,N_9614,N_9696);
nor U9787 (N_9787,N_9595,N_9632);
and U9788 (N_9788,N_9506,N_9517);
and U9789 (N_9789,N_9607,N_9683);
nor U9790 (N_9790,N_9599,N_9624);
or U9791 (N_9791,N_9738,N_9720);
nand U9792 (N_9792,N_9643,N_9667);
or U9793 (N_9793,N_9653,N_9545);
nand U9794 (N_9794,N_9660,N_9687);
and U9795 (N_9795,N_9705,N_9671);
nand U9796 (N_9796,N_9704,N_9540);
nor U9797 (N_9797,N_9512,N_9596);
or U9798 (N_9798,N_9676,N_9525);
xor U9799 (N_9799,N_9576,N_9730);
and U9800 (N_9800,N_9682,N_9590);
xor U9801 (N_9801,N_9743,N_9511);
and U9802 (N_9802,N_9581,N_9603);
and U9803 (N_9803,N_9533,N_9600);
and U9804 (N_9804,N_9569,N_9711);
xor U9805 (N_9805,N_9605,N_9549);
and U9806 (N_9806,N_9501,N_9721);
nor U9807 (N_9807,N_9714,N_9661);
and U9808 (N_9808,N_9726,N_9633);
nor U9809 (N_9809,N_9748,N_9552);
and U9810 (N_9810,N_9503,N_9604);
xor U9811 (N_9811,N_9706,N_9523);
xnor U9812 (N_9812,N_9728,N_9610);
xnor U9813 (N_9813,N_9504,N_9638);
and U9814 (N_9814,N_9644,N_9641);
nor U9815 (N_9815,N_9593,N_9509);
or U9816 (N_9816,N_9640,N_9529);
xor U9817 (N_9817,N_9745,N_9623);
and U9818 (N_9818,N_9611,N_9686);
and U9819 (N_9819,N_9597,N_9669);
nand U9820 (N_9820,N_9685,N_9651);
nor U9821 (N_9821,N_9531,N_9650);
nand U9822 (N_9822,N_9544,N_9659);
nor U9823 (N_9823,N_9532,N_9708);
xor U9824 (N_9824,N_9719,N_9642);
nand U9825 (N_9825,N_9582,N_9602);
xnor U9826 (N_9826,N_9625,N_9524);
nor U9827 (N_9827,N_9515,N_9548);
nor U9828 (N_9828,N_9541,N_9674);
or U9829 (N_9829,N_9542,N_9550);
nor U9830 (N_9830,N_9575,N_9618);
nor U9831 (N_9831,N_9695,N_9736);
or U9832 (N_9832,N_9663,N_9619);
nor U9833 (N_9833,N_9626,N_9564);
nand U9834 (N_9834,N_9615,N_9694);
xnor U9835 (N_9835,N_9703,N_9510);
nand U9836 (N_9836,N_9737,N_9534);
xnor U9837 (N_9837,N_9565,N_9519);
or U9838 (N_9838,N_9631,N_9739);
and U9839 (N_9839,N_9693,N_9555);
and U9840 (N_9840,N_9744,N_9654);
xor U9841 (N_9841,N_9732,N_9689);
xnor U9842 (N_9842,N_9500,N_9592);
nand U9843 (N_9843,N_9567,N_9698);
xnor U9844 (N_9844,N_9724,N_9536);
nand U9845 (N_9845,N_9691,N_9677);
nand U9846 (N_9846,N_9749,N_9560);
xnor U9847 (N_9847,N_9746,N_9733);
nor U9848 (N_9848,N_9608,N_9505);
nand U9849 (N_9849,N_9530,N_9578);
nor U9850 (N_9850,N_9591,N_9718);
xnor U9851 (N_9851,N_9613,N_9741);
or U9852 (N_9852,N_9715,N_9740);
or U9853 (N_9853,N_9658,N_9729);
nand U9854 (N_9854,N_9697,N_9717);
and U9855 (N_9855,N_9657,N_9648);
xor U9856 (N_9856,N_9543,N_9538);
xor U9857 (N_9857,N_9587,N_9636);
or U9858 (N_9858,N_9645,N_9716);
xor U9859 (N_9859,N_9589,N_9690);
or U9860 (N_9860,N_9672,N_9539);
or U9861 (N_9861,N_9514,N_9622);
and U9862 (N_9862,N_9518,N_9502);
nand U9863 (N_9863,N_9747,N_9666);
and U9864 (N_9864,N_9588,N_9722);
nand U9865 (N_9865,N_9554,N_9639);
xor U9866 (N_9866,N_9557,N_9601);
or U9867 (N_9867,N_9547,N_9731);
nor U9868 (N_9868,N_9688,N_9594);
or U9869 (N_9869,N_9742,N_9516);
or U9870 (N_9870,N_9579,N_9513);
xnor U9871 (N_9871,N_9734,N_9628);
nand U9872 (N_9872,N_9647,N_9634);
nor U9873 (N_9873,N_9586,N_9528);
and U9874 (N_9874,N_9712,N_9580);
nand U9875 (N_9875,N_9616,N_9645);
xor U9876 (N_9876,N_9560,N_9518);
xor U9877 (N_9877,N_9547,N_9538);
or U9878 (N_9878,N_9612,N_9571);
and U9879 (N_9879,N_9531,N_9658);
xor U9880 (N_9880,N_9624,N_9744);
xor U9881 (N_9881,N_9659,N_9593);
or U9882 (N_9882,N_9585,N_9547);
or U9883 (N_9883,N_9669,N_9651);
xnor U9884 (N_9884,N_9732,N_9707);
xor U9885 (N_9885,N_9508,N_9749);
and U9886 (N_9886,N_9500,N_9615);
nand U9887 (N_9887,N_9527,N_9627);
nand U9888 (N_9888,N_9615,N_9692);
and U9889 (N_9889,N_9615,N_9565);
xnor U9890 (N_9890,N_9712,N_9690);
nor U9891 (N_9891,N_9565,N_9673);
nor U9892 (N_9892,N_9651,N_9668);
nor U9893 (N_9893,N_9639,N_9642);
nor U9894 (N_9894,N_9737,N_9562);
or U9895 (N_9895,N_9644,N_9672);
xnor U9896 (N_9896,N_9543,N_9502);
and U9897 (N_9897,N_9619,N_9675);
nand U9898 (N_9898,N_9679,N_9695);
nand U9899 (N_9899,N_9551,N_9738);
xor U9900 (N_9900,N_9627,N_9556);
and U9901 (N_9901,N_9598,N_9747);
nor U9902 (N_9902,N_9546,N_9596);
xnor U9903 (N_9903,N_9539,N_9537);
and U9904 (N_9904,N_9743,N_9540);
and U9905 (N_9905,N_9514,N_9538);
nor U9906 (N_9906,N_9540,N_9589);
xor U9907 (N_9907,N_9619,N_9561);
and U9908 (N_9908,N_9665,N_9561);
nor U9909 (N_9909,N_9624,N_9534);
xnor U9910 (N_9910,N_9548,N_9675);
nand U9911 (N_9911,N_9539,N_9690);
nand U9912 (N_9912,N_9739,N_9614);
nor U9913 (N_9913,N_9723,N_9558);
nand U9914 (N_9914,N_9541,N_9551);
nand U9915 (N_9915,N_9587,N_9596);
nor U9916 (N_9916,N_9574,N_9721);
or U9917 (N_9917,N_9670,N_9700);
nor U9918 (N_9918,N_9645,N_9692);
or U9919 (N_9919,N_9659,N_9529);
or U9920 (N_9920,N_9700,N_9711);
nor U9921 (N_9921,N_9578,N_9681);
xnor U9922 (N_9922,N_9530,N_9580);
xnor U9923 (N_9923,N_9505,N_9502);
or U9924 (N_9924,N_9700,N_9503);
or U9925 (N_9925,N_9707,N_9557);
or U9926 (N_9926,N_9686,N_9730);
and U9927 (N_9927,N_9550,N_9673);
or U9928 (N_9928,N_9726,N_9677);
nor U9929 (N_9929,N_9682,N_9537);
nand U9930 (N_9930,N_9631,N_9593);
xnor U9931 (N_9931,N_9708,N_9723);
xnor U9932 (N_9932,N_9580,N_9698);
and U9933 (N_9933,N_9518,N_9658);
nand U9934 (N_9934,N_9706,N_9571);
nand U9935 (N_9935,N_9682,N_9651);
and U9936 (N_9936,N_9557,N_9510);
xnor U9937 (N_9937,N_9737,N_9636);
nor U9938 (N_9938,N_9563,N_9737);
or U9939 (N_9939,N_9563,N_9691);
and U9940 (N_9940,N_9571,N_9548);
xnor U9941 (N_9941,N_9633,N_9664);
nand U9942 (N_9942,N_9548,N_9607);
nand U9943 (N_9943,N_9730,N_9704);
nand U9944 (N_9944,N_9625,N_9504);
nor U9945 (N_9945,N_9616,N_9558);
nor U9946 (N_9946,N_9597,N_9646);
and U9947 (N_9947,N_9706,N_9594);
xor U9948 (N_9948,N_9564,N_9704);
or U9949 (N_9949,N_9568,N_9686);
nor U9950 (N_9950,N_9507,N_9554);
xnor U9951 (N_9951,N_9596,N_9628);
nor U9952 (N_9952,N_9641,N_9576);
xnor U9953 (N_9953,N_9534,N_9566);
nand U9954 (N_9954,N_9693,N_9548);
or U9955 (N_9955,N_9568,N_9694);
xor U9956 (N_9956,N_9549,N_9668);
or U9957 (N_9957,N_9514,N_9746);
nor U9958 (N_9958,N_9708,N_9628);
or U9959 (N_9959,N_9633,N_9690);
and U9960 (N_9960,N_9714,N_9623);
nand U9961 (N_9961,N_9599,N_9649);
or U9962 (N_9962,N_9513,N_9503);
or U9963 (N_9963,N_9679,N_9749);
nor U9964 (N_9964,N_9538,N_9739);
or U9965 (N_9965,N_9716,N_9647);
and U9966 (N_9966,N_9710,N_9661);
and U9967 (N_9967,N_9583,N_9741);
nor U9968 (N_9968,N_9724,N_9563);
xor U9969 (N_9969,N_9640,N_9596);
nand U9970 (N_9970,N_9735,N_9597);
or U9971 (N_9971,N_9647,N_9568);
xor U9972 (N_9972,N_9618,N_9592);
xnor U9973 (N_9973,N_9557,N_9705);
or U9974 (N_9974,N_9567,N_9710);
nand U9975 (N_9975,N_9736,N_9524);
nor U9976 (N_9976,N_9737,N_9590);
xor U9977 (N_9977,N_9501,N_9669);
or U9978 (N_9978,N_9600,N_9721);
nand U9979 (N_9979,N_9724,N_9557);
and U9980 (N_9980,N_9658,N_9513);
xnor U9981 (N_9981,N_9648,N_9728);
nand U9982 (N_9982,N_9741,N_9564);
xnor U9983 (N_9983,N_9625,N_9714);
nor U9984 (N_9984,N_9743,N_9576);
nand U9985 (N_9985,N_9666,N_9634);
xor U9986 (N_9986,N_9724,N_9700);
xnor U9987 (N_9987,N_9625,N_9669);
or U9988 (N_9988,N_9744,N_9587);
nor U9989 (N_9989,N_9664,N_9748);
nor U9990 (N_9990,N_9728,N_9678);
and U9991 (N_9991,N_9690,N_9513);
xnor U9992 (N_9992,N_9571,N_9654);
or U9993 (N_9993,N_9579,N_9647);
nand U9994 (N_9994,N_9630,N_9578);
nand U9995 (N_9995,N_9707,N_9500);
or U9996 (N_9996,N_9528,N_9517);
or U9997 (N_9997,N_9673,N_9652);
xnor U9998 (N_9998,N_9633,N_9655);
and U9999 (N_9999,N_9617,N_9615);
and U10000 (N_10000,N_9975,N_9900);
or U10001 (N_10001,N_9800,N_9830);
nand U10002 (N_10002,N_9783,N_9942);
or U10003 (N_10003,N_9853,N_9798);
nor U10004 (N_10004,N_9922,N_9931);
nand U10005 (N_10005,N_9791,N_9823);
xnor U10006 (N_10006,N_9768,N_9905);
xnor U10007 (N_10007,N_9896,N_9805);
nor U10008 (N_10008,N_9985,N_9822);
and U10009 (N_10009,N_9818,N_9976);
or U10010 (N_10010,N_9839,N_9821);
or U10011 (N_10011,N_9842,N_9879);
nand U10012 (N_10012,N_9772,N_9781);
and U10013 (N_10013,N_9849,N_9915);
xor U10014 (N_10014,N_9943,N_9968);
nand U10015 (N_10015,N_9996,N_9950);
or U10016 (N_10016,N_9825,N_9856);
or U10017 (N_10017,N_9992,N_9803);
and U10018 (N_10018,N_9859,N_9832);
or U10019 (N_10019,N_9850,N_9851);
nor U10020 (N_10020,N_9995,N_9979);
and U10021 (N_10021,N_9928,N_9901);
nand U10022 (N_10022,N_9993,N_9758);
nor U10023 (N_10023,N_9785,N_9880);
or U10024 (N_10024,N_9898,N_9776);
xnor U10025 (N_10025,N_9903,N_9873);
and U10026 (N_10026,N_9764,N_9933);
nor U10027 (N_10027,N_9906,N_9918);
or U10028 (N_10028,N_9925,N_9835);
and U10029 (N_10029,N_9956,N_9869);
and U10030 (N_10030,N_9899,N_9760);
or U10031 (N_10031,N_9801,N_9940);
nor U10032 (N_10032,N_9930,N_9824);
and U10033 (N_10033,N_9809,N_9989);
and U10034 (N_10034,N_9755,N_9957);
or U10035 (N_10035,N_9965,N_9958);
and U10036 (N_10036,N_9794,N_9828);
and U10037 (N_10037,N_9819,N_9786);
and U10038 (N_10038,N_9977,N_9883);
nand U10039 (N_10039,N_9787,N_9862);
nor U10040 (N_10040,N_9868,N_9757);
and U10041 (N_10041,N_9953,N_9890);
or U10042 (N_10042,N_9891,N_9987);
nor U10043 (N_10043,N_9813,N_9827);
nor U10044 (N_10044,N_9877,N_9848);
or U10045 (N_10045,N_9967,N_9959);
xor U10046 (N_10046,N_9756,N_9904);
and U10047 (N_10047,N_9952,N_9889);
and U10048 (N_10048,N_9780,N_9852);
nand U10049 (N_10049,N_9875,N_9867);
or U10050 (N_10050,N_9806,N_9847);
nand U10051 (N_10051,N_9971,N_9866);
nor U10052 (N_10052,N_9913,N_9796);
nor U10053 (N_10053,N_9834,N_9944);
nand U10054 (N_10054,N_9750,N_9935);
or U10055 (N_10055,N_9961,N_9797);
or U10056 (N_10056,N_9765,N_9921);
nand U10057 (N_10057,N_9964,N_9988);
nand U10058 (N_10058,N_9861,N_9841);
nand U10059 (N_10059,N_9816,N_9990);
nand U10060 (N_10060,N_9924,N_9811);
or U10061 (N_10061,N_9936,N_9826);
and U10062 (N_10062,N_9810,N_9878);
nand U10063 (N_10063,N_9802,N_9897);
nand U10064 (N_10064,N_9972,N_9920);
nor U10065 (N_10065,N_9991,N_9955);
and U10066 (N_10066,N_9888,N_9884);
or U10067 (N_10067,N_9941,N_9970);
or U10068 (N_10068,N_9881,N_9751);
or U10069 (N_10069,N_9817,N_9939);
nand U10070 (N_10070,N_9934,N_9857);
nor U10071 (N_10071,N_9767,N_9912);
and U10072 (N_10072,N_9982,N_9998);
nand U10073 (N_10073,N_9763,N_9782);
nand U10074 (N_10074,N_9840,N_9895);
or U10075 (N_10075,N_9854,N_9871);
nor U10076 (N_10076,N_9790,N_9784);
or U10077 (N_10077,N_9844,N_9814);
nor U10078 (N_10078,N_9812,N_9752);
xnor U10079 (N_10079,N_9815,N_9799);
and U10080 (N_10080,N_9984,N_9773);
xnor U10081 (N_10081,N_9914,N_9999);
xor U10082 (N_10082,N_9948,N_9973);
nand U10083 (N_10083,N_9917,N_9769);
nand U10084 (N_10084,N_9874,N_9908);
or U10085 (N_10085,N_9980,N_9754);
and U10086 (N_10086,N_9932,N_9882);
nor U10087 (N_10087,N_9845,N_9929);
nand U10088 (N_10088,N_9909,N_9937);
or U10089 (N_10089,N_9926,N_9774);
nand U10090 (N_10090,N_9770,N_9762);
and U10091 (N_10091,N_9870,N_9978);
nand U10092 (N_10092,N_9795,N_9833);
nand U10093 (N_10093,N_9789,N_9969);
and U10094 (N_10094,N_9876,N_9893);
nand U10095 (N_10095,N_9872,N_9907);
nand U10096 (N_10096,N_9892,N_9986);
nand U10097 (N_10097,N_9886,N_9885);
nand U10098 (N_10098,N_9804,N_9902);
or U10099 (N_10099,N_9927,N_9983);
nor U10100 (N_10100,N_9792,N_9974);
nor U10101 (N_10101,N_9759,N_9766);
nor U10102 (N_10102,N_9836,N_9949);
nor U10103 (N_10103,N_9793,N_9831);
nand U10104 (N_10104,N_9963,N_9788);
nor U10105 (N_10105,N_9981,N_9946);
nand U10106 (N_10106,N_9808,N_9843);
or U10107 (N_10107,N_9954,N_9938);
nor U10108 (N_10108,N_9863,N_9775);
nor U10109 (N_10109,N_9771,N_9829);
xor U10110 (N_10110,N_9947,N_9887);
nand U10111 (N_10111,N_9807,N_9858);
nor U10112 (N_10112,N_9864,N_9910);
nor U10113 (N_10113,N_9997,N_9923);
nand U10114 (N_10114,N_9837,N_9960);
and U10115 (N_10115,N_9945,N_9951);
and U10116 (N_10116,N_9778,N_9894);
or U10117 (N_10117,N_9962,N_9966);
xor U10118 (N_10118,N_9865,N_9779);
or U10119 (N_10119,N_9753,N_9860);
or U10120 (N_10120,N_9919,N_9994);
nor U10121 (N_10121,N_9820,N_9838);
xor U10122 (N_10122,N_9911,N_9761);
nor U10123 (N_10123,N_9916,N_9846);
xnor U10124 (N_10124,N_9777,N_9855);
nand U10125 (N_10125,N_9897,N_9805);
xnor U10126 (N_10126,N_9986,N_9932);
and U10127 (N_10127,N_9960,N_9829);
nor U10128 (N_10128,N_9942,N_9992);
nand U10129 (N_10129,N_9768,N_9774);
nand U10130 (N_10130,N_9917,N_9882);
nand U10131 (N_10131,N_9822,N_9867);
nand U10132 (N_10132,N_9758,N_9985);
or U10133 (N_10133,N_9756,N_9873);
xnor U10134 (N_10134,N_9922,N_9804);
or U10135 (N_10135,N_9796,N_9811);
xnor U10136 (N_10136,N_9776,N_9904);
nand U10137 (N_10137,N_9826,N_9776);
or U10138 (N_10138,N_9922,N_9994);
nand U10139 (N_10139,N_9935,N_9823);
xor U10140 (N_10140,N_9965,N_9978);
nand U10141 (N_10141,N_9832,N_9908);
or U10142 (N_10142,N_9926,N_9930);
nand U10143 (N_10143,N_9834,N_9783);
nor U10144 (N_10144,N_9995,N_9885);
or U10145 (N_10145,N_9793,N_9997);
and U10146 (N_10146,N_9756,N_9796);
nor U10147 (N_10147,N_9832,N_9757);
nand U10148 (N_10148,N_9934,N_9941);
nand U10149 (N_10149,N_9897,N_9933);
xnor U10150 (N_10150,N_9942,N_9911);
xor U10151 (N_10151,N_9965,N_9773);
nor U10152 (N_10152,N_9769,N_9834);
nor U10153 (N_10153,N_9934,N_9980);
nand U10154 (N_10154,N_9793,N_9836);
or U10155 (N_10155,N_9974,N_9991);
xnor U10156 (N_10156,N_9868,N_9932);
nand U10157 (N_10157,N_9800,N_9978);
xnor U10158 (N_10158,N_9982,N_9835);
nand U10159 (N_10159,N_9873,N_9823);
and U10160 (N_10160,N_9936,N_9751);
and U10161 (N_10161,N_9844,N_9875);
or U10162 (N_10162,N_9864,N_9841);
or U10163 (N_10163,N_9907,N_9987);
nand U10164 (N_10164,N_9937,N_9842);
nand U10165 (N_10165,N_9981,N_9986);
nor U10166 (N_10166,N_9853,N_9875);
xor U10167 (N_10167,N_9804,N_9886);
and U10168 (N_10168,N_9781,N_9965);
xor U10169 (N_10169,N_9863,N_9956);
nand U10170 (N_10170,N_9938,N_9906);
and U10171 (N_10171,N_9796,N_9878);
nor U10172 (N_10172,N_9953,N_9810);
and U10173 (N_10173,N_9867,N_9908);
and U10174 (N_10174,N_9774,N_9862);
nor U10175 (N_10175,N_9968,N_9965);
or U10176 (N_10176,N_9869,N_9912);
nor U10177 (N_10177,N_9751,N_9951);
nor U10178 (N_10178,N_9818,N_9912);
nand U10179 (N_10179,N_9888,N_9832);
xnor U10180 (N_10180,N_9964,N_9933);
or U10181 (N_10181,N_9813,N_9910);
xor U10182 (N_10182,N_9945,N_9941);
nor U10183 (N_10183,N_9883,N_9830);
and U10184 (N_10184,N_9860,N_9799);
nor U10185 (N_10185,N_9829,N_9775);
nand U10186 (N_10186,N_9878,N_9801);
nand U10187 (N_10187,N_9864,N_9827);
nand U10188 (N_10188,N_9918,N_9796);
nand U10189 (N_10189,N_9994,N_9996);
or U10190 (N_10190,N_9850,N_9907);
or U10191 (N_10191,N_9794,N_9872);
and U10192 (N_10192,N_9808,N_9856);
and U10193 (N_10193,N_9908,N_9757);
nand U10194 (N_10194,N_9848,N_9928);
nand U10195 (N_10195,N_9939,N_9886);
nand U10196 (N_10196,N_9895,N_9876);
and U10197 (N_10197,N_9830,N_9925);
nand U10198 (N_10198,N_9929,N_9853);
and U10199 (N_10199,N_9916,N_9874);
xor U10200 (N_10200,N_9821,N_9762);
nand U10201 (N_10201,N_9917,N_9874);
nor U10202 (N_10202,N_9829,N_9894);
xor U10203 (N_10203,N_9839,N_9769);
xnor U10204 (N_10204,N_9791,N_9960);
nor U10205 (N_10205,N_9784,N_9764);
xnor U10206 (N_10206,N_9914,N_9808);
and U10207 (N_10207,N_9972,N_9937);
and U10208 (N_10208,N_9835,N_9856);
and U10209 (N_10209,N_9871,N_9831);
and U10210 (N_10210,N_9936,N_9832);
nor U10211 (N_10211,N_9948,N_9852);
nand U10212 (N_10212,N_9878,N_9852);
nand U10213 (N_10213,N_9943,N_9963);
and U10214 (N_10214,N_9904,N_9956);
or U10215 (N_10215,N_9929,N_9944);
and U10216 (N_10216,N_9924,N_9777);
nor U10217 (N_10217,N_9781,N_9932);
and U10218 (N_10218,N_9911,N_9764);
nand U10219 (N_10219,N_9973,N_9852);
nand U10220 (N_10220,N_9826,N_9841);
and U10221 (N_10221,N_9766,N_9924);
and U10222 (N_10222,N_9992,N_9896);
nand U10223 (N_10223,N_9793,N_9906);
nand U10224 (N_10224,N_9757,N_9849);
or U10225 (N_10225,N_9792,N_9910);
nand U10226 (N_10226,N_9821,N_9785);
nand U10227 (N_10227,N_9853,N_9841);
or U10228 (N_10228,N_9796,N_9769);
xor U10229 (N_10229,N_9811,N_9931);
nor U10230 (N_10230,N_9763,N_9976);
nand U10231 (N_10231,N_9994,N_9975);
or U10232 (N_10232,N_9870,N_9769);
and U10233 (N_10233,N_9944,N_9911);
or U10234 (N_10234,N_9890,N_9815);
xnor U10235 (N_10235,N_9836,N_9897);
and U10236 (N_10236,N_9824,N_9951);
and U10237 (N_10237,N_9936,N_9790);
xor U10238 (N_10238,N_9807,N_9790);
xnor U10239 (N_10239,N_9899,N_9801);
nor U10240 (N_10240,N_9884,N_9774);
or U10241 (N_10241,N_9936,N_9812);
nor U10242 (N_10242,N_9995,N_9852);
nor U10243 (N_10243,N_9961,N_9811);
nand U10244 (N_10244,N_9840,N_9832);
or U10245 (N_10245,N_9985,N_9778);
and U10246 (N_10246,N_9752,N_9836);
nor U10247 (N_10247,N_9771,N_9822);
nor U10248 (N_10248,N_9892,N_9915);
and U10249 (N_10249,N_9849,N_9780);
and U10250 (N_10250,N_10077,N_10090);
nor U10251 (N_10251,N_10022,N_10123);
or U10252 (N_10252,N_10147,N_10110);
or U10253 (N_10253,N_10025,N_10176);
nor U10254 (N_10254,N_10130,N_10157);
nand U10255 (N_10255,N_10126,N_10214);
nor U10256 (N_10256,N_10146,N_10236);
nand U10257 (N_10257,N_10012,N_10032);
or U10258 (N_10258,N_10225,N_10233);
xnor U10259 (N_10259,N_10000,N_10241);
nor U10260 (N_10260,N_10072,N_10155);
xnor U10261 (N_10261,N_10149,N_10196);
and U10262 (N_10262,N_10228,N_10240);
nor U10263 (N_10263,N_10198,N_10001);
nand U10264 (N_10264,N_10019,N_10230);
nor U10265 (N_10265,N_10222,N_10009);
nor U10266 (N_10266,N_10010,N_10002);
and U10267 (N_10267,N_10144,N_10112);
and U10268 (N_10268,N_10177,N_10114);
nand U10269 (N_10269,N_10165,N_10101);
nand U10270 (N_10270,N_10104,N_10053);
xnor U10271 (N_10271,N_10178,N_10029);
xor U10272 (N_10272,N_10172,N_10079);
and U10273 (N_10273,N_10096,N_10071);
and U10274 (N_10274,N_10073,N_10068);
nor U10275 (N_10275,N_10092,N_10189);
or U10276 (N_10276,N_10095,N_10105);
or U10277 (N_10277,N_10132,N_10201);
or U10278 (N_10278,N_10014,N_10224);
xnor U10279 (N_10279,N_10119,N_10135);
or U10280 (N_10280,N_10218,N_10148);
or U10281 (N_10281,N_10041,N_10024);
nand U10282 (N_10282,N_10160,N_10020);
and U10283 (N_10283,N_10106,N_10061);
or U10284 (N_10284,N_10211,N_10212);
and U10285 (N_10285,N_10182,N_10205);
or U10286 (N_10286,N_10063,N_10044);
xnor U10287 (N_10287,N_10006,N_10150);
xor U10288 (N_10288,N_10076,N_10199);
and U10289 (N_10289,N_10028,N_10107);
nand U10290 (N_10290,N_10158,N_10109);
nand U10291 (N_10291,N_10216,N_10015);
nor U10292 (N_10292,N_10220,N_10026);
or U10293 (N_10293,N_10181,N_10129);
and U10294 (N_10294,N_10229,N_10121);
and U10295 (N_10295,N_10200,N_10103);
and U10296 (N_10296,N_10081,N_10162);
nor U10297 (N_10297,N_10088,N_10007);
nor U10298 (N_10298,N_10069,N_10179);
xor U10299 (N_10299,N_10238,N_10049);
and U10300 (N_10300,N_10141,N_10192);
nand U10301 (N_10301,N_10037,N_10004);
or U10302 (N_10302,N_10169,N_10183);
nor U10303 (N_10303,N_10204,N_10011);
xnor U10304 (N_10304,N_10208,N_10223);
xor U10305 (N_10305,N_10075,N_10074);
xor U10306 (N_10306,N_10239,N_10050);
or U10307 (N_10307,N_10067,N_10046);
xnor U10308 (N_10308,N_10133,N_10221);
xor U10309 (N_10309,N_10153,N_10131);
xor U10310 (N_10310,N_10138,N_10246);
nand U10311 (N_10311,N_10168,N_10226);
nand U10312 (N_10312,N_10108,N_10186);
nor U10313 (N_10313,N_10066,N_10091);
nand U10314 (N_10314,N_10042,N_10070);
nand U10315 (N_10315,N_10152,N_10234);
or U10316 (N_10316,N_10062,N_10060);
nor U10317 (N_10317,N_10143,N_10188);
xnor U10318 (N_10318,N_10030,N_10111);
nand U10319 (N_10319,N_10086,N_10163);
nand U10320 (N_10320,N_10247,N_10191);
and U10321 (N_10321,N_10159,N_10016);
or U10322 (N_10322,N_10083,N_10115);
and U10323 (N_10323,N_10033,N_10235);
nor U10324 (N_10324,N_10118,N_10059);
or U10325 (N_10325,N_10097,N_10173);
nand U10326 (N_10326,N_10185,N_10171);
nand U10327 (N_10327,N_10054,N_10156);
and U10328 (N_10328,N_10139,N_10055);
and U10329 (N_10329,N_10021,N_10151);
nand U10330 (N_10330,N_10098,N_10248);
xnor U10331 (N_10331,N_10134,N_10213);
and U10332 (N_10332,N_10142,N_10122);
and U10333 (N_10333,N_10195,N_10210);
and U10334 (N_10334,N_10102,N_10035);
xnor U10335 (N_10335,N_10080,N_10045);
xor U10336 (N_10336,N_10005,N_10018);
or U10337 (N_10337,N_10064,N_10244);
or U10338 (N_10338,N_10057,N_10167);
and U10339 (N_10339,N_10215,N_10125);
nand U10340 (N_10340,N_10166,N_10154);
nand U10341 (N_10341,N_10023,N_10180);
xor U10342 (N_10342,N_10082,N_10113);
xnor U10343 (N_10343,N_10137,N_10232);
and U10344 (N_10344,N_10043,N_10227);
xor U10345 (N_10345,N_10056,N_10194);
or U10346 (N_10346,N_10031,N_10193);
xnor U10347 (N_10347,N_10231,N_10128);
and U10348 (N_10348,N_10116,N_10017);
xor U10349 (N_10349,N_10085,N_10175);
nor U10350 (N_10350,N_10209,N_10003);
xor U10351 (N_10351,N_10197,N_10202);
nor U10352 (N_10352,N_10219,N_10084);
and U10353 (N_10353,N_10038,N_10093);
or U10354 (N_10354,N_10013,N_10243);
nand U10355 (N_10355,N_10052,N_10034);
nand U10356 (N_10356,N_10065,N_10161);
or U10357 (N_10357,N_10207,N_10140);
and U10358 (N_10358,N_10184,N_10136);
xnor U10359 (N_10359,N_10242,N_10124);
nor U10360 (N_10360,N_10087,N_10145);
nor U10361 (N_10361,N_10078,N_10036);
nor U10362 (N_10362,N_10217,N_10245);
xnor U10363 (N_10363,N_10174,N_10094);
xnor U10364 (N_10364,N_10100,N_10039);
or U10365 (N_10365,N_10237,N_10040);
and U10366 (N_10366,N_10190,N_10164);
nor U10367 (N_10367,N_10047,N_10117);
nand U10368 (N_10368,N_10048,N_10120);
nor U10369 (N_10369,N_10027,N_10203);
or U10370 (N_10370,N_10099,N_10187);
nor U10371 (N_10371,N_10089,N_10249);
or U10372 (N_10372,N_10127,N_10206);
nand U10373 (N_10373,N_10170,N_10008);
and U10374 (N_10374,N_10058,N_10051);
nand U10375 (N_10375,N_10057,N_10137);
xor U10376 (N_10376,N_10169,N_10241);
nor U10377 (N_10377,N_10021,N_10168);
or U10378 (N_10378,N_10049,N_10215);
xnor U10379 (N_10379,N_10022,N_10061);
or U10380 (N_10380,N_10211,N_10224);
or U10381 (N_10381,N_10156,N_10196);
nor U10382 (N_10382,N_10231,N_10020);
and U10383 (N_10383,N_10084,N_10023);
nand U10384 (N_10384,N_10143,N_10070);
nand U10385 (N_10385,N_10004,N_10194);
and U10386 (N_10386,N_10170,N_10010);
nor U10387 (N_10387,N_10041,N_10114);
xnor U10388 (N_10388,N_10188,N_10097);
xnor U10389 (N_10389,N_10125,N_10226);
xor U10390 (N_10390,N_10054,N_10171);
nor U10391 (N_10391,N_10242,N_10072);
and U10392 (N_10392,N_10106,N_10133);
and U10393 (N_10393,N_10234,N_10225);
or U10394 (N_10394,N_10009,N_10132);
and U10395 (N_10395,N_10067,N_10122);
and U10396 (N_10396,N_10057,N_10232);
nand U10397 (N_10397,N_10129,N_10235);
xor U10398 (N_10398,N_10223,N_10176);
and U10399 (N_10399,N_10242,N_10118);
or U10400 (N_10400,N_10209,N_10049);
nor U10401 (N_10401,N_10240,N_10176);
nor U10402 (N_10402,N_10117,N_10036);
or U10403 (N_10403,N_10247,N_10039);
nand U10404 (N_10404,N_10010,N_10067);
nor U10405 (N_10405,N_10015,N_10166);
xnor U10406 (N_10406,N_10084,N_10176);
or U10407 (N_10407,N_10128,N_10117);
and U10408 (N_10408,N_10243,N_10127);
nor U10409 (N_10409,N_10020,N_10039);
and U10410 (N_10410,N_10064,N_10106);
or U10411 (N_10411,N_10150,N_10212);
nand U10412 (N_10412,N_10136,N_10201);
nand U10413 (N_10413,N_10144,N_10106);
and U10414 (N_10414,N_10160,N_10242);
nand U10415 (N_10415,N_10122,N_10108);
or U10416 (N_10416,N_10221,N_10243);
xnor U10417 (N_10417,N_10186,N_10110);
or U10418 (N_10418,N_10161,N_10157);
or U10419 (N_10419,N_10004,N_10249);
nor U10420 (N_10420,N_10126,N_10003);
xnor U10421 (N_10421,N_10138,N_10065);
nor U10422 (N_10422,N_10111,N_10221);
and U10423 (N_10423,N_10111,N_10171);
nor U10424 (N_10424,N_10099,N_10191);
xor U10425 (N_10425,N_10230,N_10011);
nor U10426 (N_10426,N_10241,N_10117);
or U10427 (N_10427,N_10012,N_10163);
and U10428 (N_10428,N_10099,N_10008);
and U10429 (N_10429,N_10018,N_10085);
and U10430 (N_10430,N_10084,N_10099);
and U10431 (N_10431,N_10132,N_10219);
and U10432 (N_10432,N_10168,N_10130);
nand U10433 (N_10433,N_10140,N_10002);
nor U10434 (N_10434,N_10158,N_10080);
or U10435 (N_10435,N_10043,N_10155);
nand U10436 (N_10436,N_10050,N_10217);
and U10437 (N_10437,N_10105,N_10161);
nor U10438 (N_10438,N_10164,N_10236);
or U10439 (N_10439,N_10034,N_10030);
nor U10440 (N_10440,N_10145,N_10125);
nand U10441 (N_10441,N_10077,N_10007);
nand U10442 (N_10442,N_10211,N_10166);
xor U10443 (N_10443,N_10234,N_10098);
nor U10444 (N_10444,N_10042,N_10220);
xnor U10445 (N_10445,N_10200,N_10048);
nand U10446 (N_10446,N_10238,N_10187);
and U10447 (N_10447,N_10215,N_10236);
xor U10448 (N_10448,N_10142,N_10204);
or U10449 (N_10449,N_10120,N_10193);
xnor U10450 (N_10450,N_10243,N_10199);
or U10451 (N_10451,N_10049,N_10072);
xor U10452 (N_10452,N_10159,N_10028);
xnor U10453 (N_10453,N_10006,N_10112);
xor U10454 (N_10454,N_10163,N_10168);
nor U10455 (N_10455,N_10180,N_10209);
nand U10456 (N_10456,N_10123,N_10040);
xor U10457 (N_10457,N_10145,N_10001);
or U10458 (N_10458,N_10128,N_10043);
and U10459 (N_10459,N_10116,N_10075);
nor U10460 (N_10460,N_10153,N_10037);
nand U10461 (N_10461,N_10138,N_10195);
nand U10462 (N_10462,N_10031,N_10196);
nand U10463 (N_10463,N_10093,N_10125);
nand U10464 (N_10464,N_10032,N_10067);
nand U10465 (N_10465,N_10181,N_10183);
or U10466 (N_10466,N_10073,N_10152);
or U10467 (N_10467,N_10107,N_10088);
and U10468 (N_10468,N_10205,N_10186);
xnor U10469 (N_10469,N_10021,N_10220);
nand U10470 (N_10470,N_10238,N_10108);
nor U10471 (N_10471,N_10233,N_10245);
xnor U10472 (N_10472,N_10021,N_10125);
and U10473 (N_10473,N_10230,N_10233);
and U10474 (N_10474,N_10081,N_10159);
xor U10475 (N_10475,N_10037,N_10073);
nor U10476 (N_10476,N_10226,N_10053);
xnor U10477 (N_10477,N_10003,N_10152);
nand U10478 (N_10478,N_10050,N_10123);
and U10479 (N_10479,N_10067,N_10157);
and U10480 (N_10480,N_10038,N_10148);
nand U10481 (N_10481,N_10237,N_10052);
xnor U10482 (N_10482,N_10062,N_10235);
and U10483 (N_10483,N_10234,N_10224);
xnor U10484 (N_10484,N_10191,N_10246);
nor U10485 (N_10485,N_10032,N_10112);
and U10486 (N_10486,N_10111,N_10193);
nor U10487 (N_10487,N_10171,N_10133);
or U10488 (N_10488,N_10088,N_10009);
nand U10489 (N_10489,N_10101,N_10074);
or U10490 (N_10490,N_10221,N_10101);
and U10491 (N_10491,N_10096,N_10188);
xnor U10492 (N_10492,N_10175,N_10233);
and U10493 (N_10493,N_10030,N_10141);
nor U10494 (N_10494,N_10016,N_10127);
xnor U10495 (N_10495,N_10035,N_10027);
or U10496 (N_10496,N_10008,N_10048);
xor U10497 (N_10497,N_10243,N_10226);
xor U10498 (N_10498,N_10220,N_10001);
and U10499 (N_10499,N_10006,N_10186);
nor U10500 (N_10500,N_10436,N_10439);
xnor U10501 (N_10501,N_10313,N_10354);
xnor U10502 (N_10502,N_10386,N_10307);
nor U10503 (N_10503,N_10331,N_10359);
nand U10504 (N_10504,N_10365,N_10356);
nand U10505 (N_10505,N_10312,N_10486);
and U10506 (N_10506,N_10363,N_10333);
or U10507 (N_10507,N_10300,N_10367);
or U10508 (N_10508,N_10343,N_10492);
and U10509 (N_10509,N_10444,N_10419);
nor U10510 (N_10510,N_10472,N_10303);
nor U10511 (N_10511,N_10376,N_10299);
and U10512 (N_10512,N_10301,N_10268);
xnor U10513 (N_10513,N_10403,N_10498);
xor U10514 (N_10514,N_10291,N_10379);
nor U10515 (N_10515,N_10271,N_10448);
or U10516 (N_10516,N_10273,N_10325);
xor U10517 (N_10517,N_10450,N_10378);
or U10518 (N_10518,N_10382,N_10362);
nand U10519 (N_10519,N_10267,N_10321);
and U10520 (N_10520,N_10457,N_10285);
and U10521 (N_10521,N_10428,N_10259);
nor U10522 (N_10522,N_10329,N_10318);
and U10523 (N_10523,N_10425,N_10401);
nor U10524 (N_10524,N_10264,N_10395);
or U10525 (N_10525,N_10319,N_10347);
or U10526 (N_10526,N_10274,N_10293);
nor U10527 (N_10527,N_10396,N_10353);
nor U10528 (N_10528,N_10371,N_10421);
nand U10529 (N_10529,N_10465,N_10314);
or U10530 (N_10530,N_10435,N_10361);
or U10531 (N_10531,N_10449,N_10494);
nor U10532 (N_10532,N_10466,N_10281);
and U10533 (N_10533,N_10487,N_10430);
nor U10534 (N_10534,N_10337,N_10459);
nor U10535 (N_10535,N_10404,N_10263);
nor U10536 (N_10536,N_10284,N_10276);
xnor U10537 (N_10537,N_10411,N_10364);
and U10538 (N_10538,N_10324,N_10289);
xnor U10539 (N_10539,N_10406,N_10261);
nand U10540 (N_10540,N_10458,N_10352);
nand U10541 (N_10541,N_10255,N_10456);
xor U10542 (N_10542,N_10477,N_10470);
or U10543 (N_10543,N_10310,N_10393);
nor U10544 (N_10544,N_10429,N_10489);
and U10545 (N_10545,N_10366,N_10311);
and U10546 (N_10546,N_10417,N_10455);
nand U10547 (N_10547,N_10265,N_10344);
xnor U10548 (N_10548,N_10335,N_10341);
xor U10549 (N_10549,N_10290,N_10295);
and U10550 (N_10550,N_10283,N_10479);
nor U10551 (N_10551,N_10407,N_10409);
nor U10552 (N_10552,N_10345,N_10447);
and U10553 (N_10553,N_10340,N_10254);
and U10554 (N_10554,N_10413,N_10277);
or U10555 (N_10555,N_10297,N_10309);
nand U10556 (N_10556,N_10278,N_10256);
xnor U10557 (N_10557,N_10330,N_10391);
xor U10558 (N_10558,N_10420,N_10397);
nor U10559 (N_10559,N_10402,N_10262);
and U10560 (N_10560,N_10424,N_10322);
and U10561 (N_10561,N_10334,N_10306);
and U10562 (N_10562,N_10369,N_10380);
or U10563 (N_10563,N_10302,N_10328);
xnor U10564 (N_10564,N_10480,N_10394);
xnor U10565 (N_10565,N_10412,N_10390);
and U10566 (N_10566,N_10499,N_10279);
or U10567 (N_10567,N_10317,N_10304);
nor U10568 (N_10568,N_10440,N_10437);
xnor U10569 (N_10569,N_10443,N_10408);
xor U10570 (N_10570,N_10422,N_10308);
xor U10571 (N_10571,N_10383,N_10346);
nor U10572 (N_10572,N_10358,N_10451);
or U10573 (N_10573,N_10296,N_10280);
xor U10574 (N_10574,N_10462,N_10305);
or U10575 (N_10575,N_10389,N_10453);
nor U10576 (N_10576,N_10342,N_10253);
and U10577 (N_10577,N_10475,N_10468);
and U10578 (N_10578,N_10415,N_10372);
nand U10579 (N_10579,N_10438,N_10463);
nand U10580 (N_10580,N_10288,N_10351);
and U10581 (N_10581,N_10461,N_10484);
and U10582 (N_10582,N_10410,N_10442);
nor U10583 (N_10583,N_10482,N_10478);
and U10584 (N_10584,N_10483,N_10323);
or U10585 (N_10585,N_10473,N_10441);
and U10586 (N_10586,N_10286,N_10399);
or U10587 (N_10587,N_10320,N_10460);
or U10588 (N_10588,N_10282,N_10474);
xor U10589 (N_10589,N_10427,N_10381);
nand U10590 (N_10590,N_10467,N_10418);
or U10591 (N_10591,N_10400,N_10495);
nand U10592 (N_10592,N_10452,N_10497);
or U10593 (N_10593,N_10339,N_10433);
xor U10594 (N_10594,N_10454,N_10388);
nor U10595 (N_10595,N_10292,N_10387);
or U10596 (N_10596,N_10370,N_10485);
nor U10597 (N_10597,N_10385,N_10338);
xnor U10598 (N_10598,N_10348,N_10490);
or U10599 (N_10599,N_10252,N_10392);
nor U10600 (N_10600,N_10272,N_10446);
nand U10601 (N_10601,N_10464,N_10287);
nor U10602 (N_10602,N_10373,N_10332);
xnor U10603 (N_10603,N_10298,N_10368);
xor U10604 (N_10604,N_10416,N_10336);
xor U10605 (N_10605,N_10349,N_10469);
and U10606 (N_10606,N_10257,N_10405);
xnor U10607 (N_10607,N_10496,N_10426);
xnor U10608 (N_10608,N_10476,N_10258);
and U10609 (N_10609,N_10350,N_10384);
nand U10610 (N_10610,N_10270,N_10260);
nor U10611 (N_10611,N_10471,N_10445);
xor U10612 (N_10612,N_10250,N_10326);
xor U10613 (N_10613,N_10481,N_10315);
nor U10614 (N_10614,N_10431,N_10375);
nand U10615 (N_10615,N_10269,N_10355);
nand U10616 (N_10616,N_10294,N_10414);
and U10617 (N_10617,N_10491,N_10275);
and U10618 (N_10618,N_10327,N_10357);
nand U10619 (N_10619,N_10398,N_10251);
and U10620 (N_10620,N_10423,N_10374);
xnor U10621 (N_10621,N_10493,N_10434);
or U10622 (N_10622,N_10266,N_10377);
nor U10623 (N_10623,N_10360,N_10488);
xnor U10624 (N_10624,N_10432,N_10316);
xnor U10625 (N_10625,N_10310,N_10499);
nand U10626 (N_10626,N_10400,N_10488);
xnor U10627 (N_10627,N_10499,N_10263);
xor U10628 (N_10628,N_10453,N_10376);
nor U10629 (N_10629,N_10417,N_10329);
and U10630 (N_10630,N_10262,N_10284);
and U10631 (N_10631,N_10318,N_10341);
nor U10632 (N_10632,N_10480,N_10427);
and U10633 (N_10633,N_10265,N_10402);
nand U10634 (N_10634,N_10498,N_10375);
xor U10635 (N_10635,N_10322,N_10457);
nor U10636 (N_10636,N_10431,N_10395);
or U10637 (N_10637,N_10341,N_10382);
and U10638 (N_10638,N_10458,N_10408);
nand U10639 (N_10639,N_10319,N_10438);
or U10640 (N_10640,N_10363,N_10402);
and U10641 (N_10641,N_10275,N_10367);
or U10642 (N_10642,N_10427,N_10252);
or U10643 (N_10643,N_10420,N_10427);
and U10644 (N_10644,N_10490,N_10496);
and U10645 (N_10645,N_10274,N_10423);
xnor U10646 (N_10646,N_10435,N_10323);
nand U10647 (N_10647,N_10250,N_10484);
or U10648 (N_10648,N_10314,N_10458);
nor U10649 (N_10649,N_10253,N_10387);
nand U10650 (N_10650,N_10440,N_10272);
nand U10651 (N_10651,N_10289,N_10426);
nand U10652 (N_10652,N_10488,N_10273);
and U10653 (N_10653,N_10438,N_10451);
xnor U10654 (N_10654,N_10291,N_10310);
nor U10655 (N_10655,N_10434,N_10273);
nand U10656 (N_10656,N_10281,N_10311);
nand U10657 (N_10657,N_10435,N_10458);
nor U10658 (N_10658,N_10282,N_10444);
nand U10659 (N_10659,N_10365,N_10362);
xor U10660 (N_10660,N_10321,N_10368);
or U10661 (N_10661,N_10322,N_10463);
xor U10662 (N_10662,N_10274,N_10329);
or U10663 (N_10663,N_10433,N_10360);
and U10664 (N_10664,N_10393,N_10341);
nor U10665 (N_10665,N_10351,N_10354);
nor U10666 (N_10666,N_10363,N_10259);
or U10667 (N_10667,N_10285,N_10293);
and U10668 (N_10668,N_10284,N_10482);
and U10669 (N_10669,N_10381,N_10401);
xnor U10670 (N_10670,N_10288,N_10313);
xnor U10671 (N_10671,N_10290,N_10469);
and U10672 (N_10672,N_10262,N_10302);
or U10673 (N_10673,N_10278,N_10367);
nor U10674 (N_10674,N_10313,N_10255);
or U10675 (N_10675,N_10327,N_10423);
nand U10676 (N_10676,N_10358,N_10268);
and U10677 (N_10677,N_10329,N_10309);
or U10678 (N_10678,N_10466,N_10378);
and U10679 (N_10679,N_10454,N_10499);
and U10680 (N_10680,N_10357,N_10308);
or U10681 (N_10681,N_10292,N_10441);
nor U10682 (N_10682,N_10371,N_10403);
and U10683 (N_10683,N_10341,N_10365);
nand U10684 (N_10684,N_10477,N_10454);
nor U10685 (N_10685,N_10392,N_10398);
nand U10686 (N_10686,N_10459,N_10350);
nand U10687 (N_10687,N_10365,N_10252);
nor U10688 (N_10688,N_10274,N_10389);
nor U10689 (N_10689,N_10433,N_10464);
or U10690 (N_10690,N_10443,N_10390);
nor U10691 (N_10691,N_10297,N_10416);
or U10692 (N_10692,N_10436,N_10403);
nand U10693 (N_10693,N_10401,N_10308);
and U10694 (N_10694,N_10488,N_10482);
and U10695 (N_10695,N_10365,N_10401);
nand U10696 (N_10696,N_10482,N_10271);
xor U10697 (N_10697,N_10304,N_10295);
or U10698 (N_10698,N_10448,N_10277);
and U10699 (N_10699,N_10450,N_10479);
xnor U10700 (N_10700,N_10396,N_10496);
xor U10701 (N_10701,N_10430,N_10471);
nand U10702 (N_10702,N_10420,N_10387);
and U10703 (N_10703,N_10419,N_10384);
nor U10704 (N_10704,N_10423,N_10440);
xnor U10705 (N_10705,N_10449,N_10454);
or U10706 (N_10706,N_10437,N_10456);
or U10707 (N_10707,N_10438,N_10297);
nor U10708 (N_10708,N_10408,N_10260);
nand U10709 (N_10709,N_10389,N_10385);
and U10710 (N_10710,N_10273,N_10440);
or U10711 (N_10711,N_10416,N_10413);
or U10712 (N_10712,N_10271,N_10351);
nand U10713 (N_10713,N_10450,N_10404);
and U10714 (N_10714,N_10419,N_10481);
nand U10715 (N_10715,N_10282,N_10377);
nor U10716 (N_10716,N_10386,N_10495);
and U10717 (N_10717,N_10468,N_10402);
and U10718 (N_10718,N_10268,N_10363);
nor U10719 (N_10719,N_10453,N_10362);
and U10720 (N_10720,N_10419,N_10322);
or U10721 (N_10721,N_10289,N_10451);
xnor U10722 (N_10722,N_10372,N_10376);
nor U10723 (N_10723,N_10463,N_10367);
or U10724 (N_10724,N_10435,N_10459);
or U10725 (N_10725,N_10383,N_10365);
and U10726 (N_10726,N_10350,N_10386);
xnor U10727 (N_10727,N_10478,N_10450);
or U10728 (N_10728,N_10404,N_10259);
nand U10729 (N_10729,N_10308,N_10483);
or U10730 (N_10730,N_10424,N_10388);
or U10731 (N_10731,N_10454,N_10456);
nand U10732 (N_10732,N_10381,N_10336);
and U10733 (N_10733,N_10271,N_10415);
or U10734 (N_10734,N_10271,N_10467);
and U10735 (N_10735,N_10250,N_10313);
or U10736 (N_10736,N_10315,N_10452);
and U10737 (N_10737,N_10461,N_10431);
nor U10738 (N_10738,N_10340,N_10319);
nor U10739 (N_10739,N_10378,N_10325);
and U10740 (N_10740,N_10331,N_10274);
or U10741 (N_10741,N_10452,N_10345);
nand U10742 (N_10742,N_10420,N_10428);
xor U10743 (N_10743,N_10349,N_10352);
and U10744 (N_10744,N_10327,N_10338);
nand U10745 (N_10745,N_10411,N_10313);
and U10746 (N_10746,N_10454,N_10336);
nor U10747 (N_10747,N_10314,N_10255);
or U10748 (N_10748,N_10430,N_10251);
xor U10749 (N_10749,N_10395,N_10272);
and U10750 (N_10750,N_10617,N_10523);
nand U10751 (N_10751,N_10736,N_10661);
and U10752 (N_10752,N_10651,N_10627);
nand U10753 (N_10753,N_10587,N_10606);
nand U10754 (N_10754,N_10598,N_10748);
or U10755 (N_10755,N_10577,N_10637);
and U10756 (N_10756,N_10695,N_10729);
nand U10757 (N_10757,N_10520,N_10526);
nand U10758 (N_10758,N_10723,N_10713);
or U10759 (N_10759,N_10676,N_10559);
and U10760 (N_10760,N_10660,N_10508);
and U10761 (N_10761,N_10571,N_10739);
or U10762 (N_10762,N_10538,N_10721);
nor U10763 (N_10763,N_10543,N_10730);
nor U10764 (N_10764,N_10649,N_10532);
xnor U10765 (N_10765,N_10528,N_10529);
and U10766 (N_10766,N_10607,N_10689);
nor U10767 (N_10767,N_10634,N_10547);
or U10768 (N_10768,N_10553,N_10568);
or U10769 (N_10769,N_10671,N_10658);
or U10770 (N_10770,N_10515,N_10597);
nor U10771 (N_10771,N_10717,N_10708);
nand U10772 (N_10772,N_10635,N_10629);
nor U10773 (N_10773,N_10584,N_10690);
nor U10774 (N_10774,N_10534,N_10565);
xor U10775 (N_10775,N_10657,N_10745);
and U10776 (N_10776,N_10731,N_10561);
nor U10777 (N_10777,N_10572,N_10623);
or U10778 (N_10778,N_10616,N_10602);
nor U10779 (N_10779,N_10593,N_10533);
nor U10780 (N_10780,N_10664,N_10514);
nand U10781 (N_10781,N_10503,N_10720);
nor U10782 (N_10782,N_10619,N_10611);
nand U10783 (N_10783,N_10662,N_10679);
nand U10784 (N_10784,N_10700,N_10556);
xnor U10785 (N_10785,N_10567,N_10653);
nand U10786 (N_10786,N_10531,N_10574);
xor U10787 (N_10787,N_10507,N_10677);
and U10788 (N_10788,N_10636,N_10734);
nand U10789 (N_10789,N_10663,N_10699);
nor U10790 (N_10790,N_10537,N_10579);
xor U10791 (N_10791,N_10749,N_10554);
and U10792 (N_10792,N_10605,N_10702);
nand U10793 (N_10793,N_10578,N_10674);
nor U10794 (N_10794,N_10640,N_10545);
xnor U10795 (N_10795,N_10518,N_10673);
and U10796 (N_10796,N_10557,N_10610);
or U10797 (N_10797,N_10712,N_10551);
and U10798 (N_10798,N_10624,N_10599);
nand U10799 (N_10799,N_10678,N_10737);
or U10800 (N_10800,N_10550,N_10648);
nor U10801 (N_10801,N_10686,N_10724);
nand U10802 (N_10802,N_10659,N_10718);
or U10803 (N_10803,N_10735,N_10600);
nor U10804 (N_10804,N_10536,N_10522);
or U10805 (N_10805,N_10524,N_10590);
nand U10806 (N_10806,N_10620,N_10705);
nand U10807 (N_10807,N_10668,N_10741);
nand U10808 (N_10808,N_10563,N_10552);
and U10809 (N_10809,N_10628,N_10687);
or U10810 (N_10810,N_10513,N_10680);
xnor U10811 (N_10811,N_10516,N_10615);
or U10812 (N_10812,N_10525,N_10733);
and U10813 (N_10813,N_10633,N_10509);
and U10814 (N_10814,N_10530,N_10746);
xnor U10815 (N_10815,N_10594,N_10697);
nand U10816 (N_10816,N_10585,N_10639);
nand U10817 (N_10817,N_10609,N_10544);
nand U10818 (N_10818,N_10696,N_10645);
xor U10819 (N_10819,N_10728,N_10747);
xor U10820 (N_10820,N_10710,N_10719);
nand U10821 (N_10821,N_10519,N_10738);
or U10822 (N_10822,N_10506,N_10641);
or U10823 (N_10823,N_10670,N_10706);
and U10824 (N_10824,N_10669,N_10698);
nor U10825 (N_10825,N_10727,N_10682);
or U10826 (N_10826,N_10622,N_10707);
nand U10827 (N_10827,N_10573,N_10608);
or U10828 (N_10828,N_10715,N_10586);
nand U10829 (N_10829,N_10596,N_10643);
or U10830 (N_10830,N_10672,N_10591);
nor U10831 (N_10831,N_10694,N_10638);
xor U10832 (N_10832,N_10541,N_10539);
xnor U10833 (N_10833,N_10501,N_10742);
xnor U10834 (N_10834,N_10564,N_10691);
xnor U10835 (N_10835,N_10502,N_10511);
nor U10836 (N_10836,N_10632,N_10684);
nor U10837 (N_10837,N_10601,N_10740);
xor U10838 (N_10838,N_10667,N_10744);
nor U10839 (N_10839,N_10681,N_10630);
or U10840 (N_10840,N_10644,N_10535);
xor U10841 (N_10841,N_10583,N_10560);
nor U10842 (N_10842,N_10711,N_10562);
nor U10843 (N_10843,N_10592,N_10625);
nor U10844 (N_10844,N_10692,N_10549);
nor U10845 (N_10845,N_10714,N_10704);
xnor U10846 (N_10846,N_10626,N_10569);
xnor U10847 (N_10847,N_10703,N_10618);
or U10848 (N_10848,N_10546,N_10576);
or U10849 (N_10849,N_10575,N_10656);
or U10850 (N_10850,N_10621,N_10588);
and U10851 (N_10851,N_10716,N_10566);
and U10852 (N_10852,N_10517,N_10650);
nand U10853 (N_10853,N_10654,N_10504);
xnor U10854 (N_10854,N_10521,N_10614);
nor U10855 (N_10855,N_10505,N_10647);
and U10856 (N_10856,N_10725,N_10722);
nor U10857 (N_10857,N_10683,N_10675);
nand U10858 (N_10858,N_10510,N_10512);
nor U10859 (N_10859,N_10580,N_10732);
or U10860 (N_10860,N_10743,N_10688);
xor U10861 (N_10861,N_10570,N_10642);
nor U10862 (N_10862,N_10666,N_10693);
and U10863 (N_10863,N_10685,N_10603);
and U10864 (N_10864,N_10581,N_10604);
xnor U10865 (N_10865,N_10527,N_10540);
nor U10866 (N_10866,N_10612,N_10665);
and U10867 (N_10867,N_10652,N_10655);
or U10868 (N_10868,N_10613,N_10726);
nand U10869 (N_10869,N_10701,N_10558);
or U10870 (N_10870,N_10646,N_10500);
nand U10871 (N_10871,N_10548,N_10631);
nand U10872 (N_10872,N_10595,N_10555);
and U10873 (N_10873,N_10709,N_10589);
or U10874 (N_10874,N_10542,N_10582);
and U10875 (N_10875,N_10614,N_10655);
nor U10876 (N_10876,N_10521,N_10623);
or U10877 (N_10877,N_10611,N_10513);
or U10878 (N_10878,N_10625,N_10516);
or U10879 (N_10879,N_10732,N_10632);
xnor U10880 (N_10880,N_10585,N_10713);
and U10881 (N_10881,N_10738,N_10552);
xor U10882 (N_10882,N_10537,N_10630);
xor U10883 (N_10883,N_10560,N_10657);
nor U10884 (N_10884,N_10598,N_10648);
and U10885 (N_10885,N_10682,N_10508);
nand U10886 (N_10886,N_10521,N_10600);
nor U10887 (N_10887,N_10603,N_10690);
and U10888 (N_10888,N_10541,N_10609);
and U10889 (N_10889,N_10591,N_10643);
and U10890 (N_10890,N_10608,N_10562);
or U10891 (N_10891,N_10653,N_10635);
or U10892 (N_10892,N_10582,N_10603);
nor U10893 (N_10893,N_10512,N_10557);
and U10894 (N_10894,N_10518,N_10534);
nor U10895 (N_10895,N_10711,N_10638);
nand U10896 (N_10896,N_10672,N_10732);
or U10897 (N_10897,N_10710,N_10542);
nand U10898 (N_10898,N_10737,N_10502);
or U10899 (N_10899,N_10633,N_10643);
and U10900 (N_10900,N_10590,N_10615);
nor U10901 (N_10901,N_10723,N_10624);
and U10902 (N_10902,N_10559,N_10551);
nand U10903 (N_10903,N_10565,N_10529);
nor U10904 (N_10904,N_10610,N_10626);
and U10905 (N_10905,N_10688,N_10650);
nand U10906 (N_10906,N_10568,N_10694);
nor U10907 (N_10907,N_10674,N_10607);
nor U10908 (N_10908,N_10631,N_10602);
nor U10909 (N_10909,N_10626,N_10585);
nor U10910 (N_10910,N_10698,N_10664);
nor U10911 (N_10911,N_10718,N_10707);
xnor U10912 (N_10912,N_10513,N_10700);
nor U10913 (N_10913,N_10729,N_10748);
or U10914 (N_10914,N_10715,N_10520);
and U10915 (N_10915,N_10735,N_10506);
or U10916 (N_10916,N_10711,N_10550);
nor U10917 (N_10917,N_10614,N_10549);
or U10918 (N_10918,N_10581,N_10692);
and U10919 (N_10919,N_10557,N_10712);
or U10920 (N_10920,N_10597,N_10745);
or U10921 (N_10921,N_10628,N_10542);
nand U10922 (N_10922,N_10691,N_10507);
or U10923 (N_10923,N_10570,N_10718);
nor U10924 (N_10924,N_10659,N_10559);
and U10925 (N_10925,N_10648,N_10627);
xnor U10926 (N_10926,N_10636,N_10516);
nor U10927 (N_10927,N_10655,N_10738);
and U10928 (N_10928,N_10522,N_10572);
nand U10929 (N_10929,N_10508,N_10633);
nand U10930 (N_10930,N_10685,N_10513);
and U10931 (N_10931,N_10579,N_10682);
xor U10932 (N_10932,N_10683,N_10672);
and U10933 (N_10933,N_10640,N_10514);
or U10934 (N_10934,N_10509,N_10527);
or U10935 (N_10935,N_10723,N_10651);
xor U10936 (N_10936,N_10555,N_10515);
nand U10937 (N_10937,N_10654,N_10671);
and U10938 (N_10938,N_10732,N_10638);
and U10939 (N_10939,N_10603,N_10647);
nor U10940 (N_10940,N_10587,N_10512);
or U10941 (N_10941,N_10693,N_10504);
nor U10942 (N_10942,N_10709,N_10627);
xor U10943 (N_10943,N_10715,N_10664);
or U10944 (N_10944,N_10647,N_10604);
and U10945 (N_10945,N_10594,N_10573);
nand U10946 (N_10946,N_10624,N_10654);
nor U10947 (N_10947,N_10672,N_10737);
nor U10948 (N_10948,N_10600,N_10554);
nor U10949 (N_10949,N_10610,N_10579);
xnor U10950 (N_10950,N_10687,N_10510);
nand U10951 (N_10951,N_10532,N_10712);
xnor U10952 (N_10952,N_10518,N_10537);
or U10953 (N_10953,N_10630,N_10506);
nor U10954 (N_10954,N_10721,N_10659);
nand U10955 (N_10955,N_10721,N_10528);
xor U10956 (N_10956,N_10738,N_10747);
and U10957 (N_10957,N_10611,N_10530);
xor U10958 (N_10958,N_10532,N_10527);
nand U10959 (N_10959,N_10532,N_10663);
xnor U10960 (N_10960,N_10663,N_10534);
xnor U10961 (N_10961,N_10593,N_10581);
or U10962 (N_10962,N_10746,N_10624);
xor U10963 (N_10963,N_10714,N_10613);
or U10964 (N_10964,N_10642,N_10527);
nand U10965 (N_10965,N_10564,N_10719);
nor U10966 (N_10966,N_10618,N_10640);
or U10967 (N_10967,N_10595,N_10678);
nand U10968 (N_10968,N_10522,N_10579);
or U10969 (N_10969,N_10588,N_10678);
and U10970 (N_10970,N_10669,N_10660);
or U10971 (N_10971,N_10729,N_10643);
nand U10972 (N_10972,N_10592,N_10516);
nor U10973 (N_10973,N_10640,N_10733);
or U10974 (N_10974,N_10732,N_10533);
nor U10975 (N_10975,N_10617,N_10522);
nor U10976 (N_10976,N_10543,N_10668);
or U10977 (N_10977,N_10580,N_10671);
nor U10978 (N_10978,N_10662,N_10574);
xnor U10979 (N_10979,N_10542,N_10525);
nand U10980 (N_10980,N_10619,N_10530);
nor U10981 (N_10981,N_10712,N_10578);
nor U10982 (N_10982,N_10683,N_10574);
nor U10983 (N_10983,N_10735,N_10620);
or U10984 (N_10984,N_10639,N_10743);
xnor U10985 (N_10985,N_10703,N_10631);
nor U10986 (N_10986,N_10630,N_10584);
xor U10987 (N_10987,N_10535,N_10655);
or U10988 (N_10988,N_10725,N_10543);
nand U10989 (N_10989,N_10611,N_10684);
nand U10990 (N_10990,N_10675,N_10633);
or U10991 (N_10991,N_10540,N_10565);
nor U10992 (N_10992,N_10705,N_10561);
or U10993 (N_10993,N_10512,N_10742);
nand U10994 (N_10994,N_10717,N_10556);
xnor U10995 (N_10995,N_10689,N_10540);
xnor U10996 (N_10996,N_10735,N_10736);
or U10997 (N_10997,N_10707,N_10591);
and U10998 (N_10998,N_10549,N_10664);
xor U10999 (N_10999,N_10616,N_10558);
nor U11000 (N_11000,N_10944,N_10770);
and U11001 (N_11001,N_10939,N_10879);
nor U11002 (N_11002,N_10885,N_10765);
nor U11003 (N_11003,N_10900,N_10966);
nor U11004 (N_11004,N_10799,N_10921);
and U11005 (N_11005,N_10769,N_10842);
xor U11006 (N_11006,N_10898,N_10903);
or U11007 (N_11007,N_10923,N_10912);
and U11008 (N_11008,N_10779,N_10946);
and U11009 (N_11009,N_10959,N_10845);
or U11010 (N_11010,N_10777,N_10920);
nand U11011 (N_11011,N_10774,N_10865);
or U11012 (N_11012,N_10801,N_10907);
xor U11013 (N_11013,N_10975,N_10827);
xnor U11014 (N_11014,N_10823,N_10994);
or U11015 (N_11015,N_10965,N_10943);
nand U11016 (N_11016,N_10895,N_10928);
nor U11017 (N_11017,N_10844,N_10876);
or U11018 (N_11018,N_10970,N_10983);
and U11019 (N_11019,N_10955,N_10889);
and U11020 (N_11020,N_10767,N_10961);
nand U11021 (N_11021,N_10836,N_10753);
nor U11022 (N_11022,N_10820,N_10817);
nand U11023 (N_11023,N_10870,N_10888);
nor U11024 (N_11024,N_10978,N_10853);
nand U11025 (N_11025,N_10788,N_10843);
or U11026 (N_11026,N_10868,N_10867);
nand U11027 (N_11027,N_10794,N_10951);
nand U11028 (N_11028,N_10996,N_10755);
nor U11029 (N_11029,N_10851,N_10809);
xor U11030 (N_11030,N_10798,N_10783);
nand U11031 (N_11031,N_10887,N_10785);
nand U11032 (N_11032,N_10913,N_10942);
and U11033 (N_11033,N_10778,N_10856);
or U11034 (N_11034,N_10986,N_10969);
xnor U11035 (N_11035,N_10873,N_10808);
nor U11036 (N_11036,N_10901,N_10968);
xnor U11037 (N_11037,N_10987,N_10859);
or U11038 (N_11038,N_10833,N_10752);
or U11039 (N_11039,N_10991,N_10750);
and U11040 (N_11040,N_10791,N_10818);
or U11041 (N_11041,N_10981,N_10758);
and U11042 (N_11042,N_10926,N_10771);
and U11043 (N_11043,N_10953,N_10916);
and U11044 (N_11044,N_10947,N_10899);
nor U11045 (N_11045,N_10945,N_10977);
or U11046 (N_11046,N_10906,N_10908);
nor U11047 (N_11047,N_10919,N_10979);
and U11048 (N_11048,N_10917,N_10963);
xor U11049 (N_11049,N_10890,N_10999);
nand U11050 (N_11050,N_10782,N_10918);
nand U11051 (N_11051,N_10967,N_10762);
nand U11052 (N_11052,N_10846,N_10992);
nor U11053 (N_11053,N_10790,N_10909);
or U11054 (N_11054,N_10819,N_10993);
nor U11055 (N_11055,N_10948,N_10829);
nand U11056 (N_11056,N_10830,N_10828);
or U11057 (N_11057,N_10897,N_10858);
xnor U11058 (N_11058,N_10998,N_10850);
xor U11059 (N_11059,N_10924,N_10795);
xnor U11060 (N_11060,N_10973,N_10780);
xnor U11061 (N_11061,N_10796,N_10892);
or U11062 (N_11062,N_10766,N_10922);
xor U11063 (N_11063,N_10800,N_10935);
and U11064 (N_11064,N_10880,N_10826);
nor U11065 (N_11065,N_10840,N_10960);
and U11066 (N_11066,N_10927,N_10754);
nand U11067 (N_11067,N_10952,N_10806);
nor U11068 (N_11068,N_10756,N_10849);
nor U11069 (N_11069,N_10982,N_10934);
nor U11070 (N_11070,N_10886,N_10792);
nand U11071 (N_11071,N_10757,N_10929);
or U11072 (N_11072,N_10980,N_10878);
or U11073 (N_11073,N_10989,N_10874);
and U11074 (N_11074,N_10882,N_10976);
and U11075 (N_11075,N_10835,N_10797);
xnor U11076 (N_11076,N_10787,N_10915);
nor U11077 (N_11077,N_10995,N_10781);
xnor U11078 (N_11078,N_10875,N_10932);
nand U11079 (N_11079,N_10894,N_10825);
or U11080 (N_11080,N_10805,N_10848);
xor U11081 (N_11081,N_10904,N_10861);
or U11082 (N_11082,N_10764,N_10881);
or U11083 (N_11083,N_10810,N_10854);
or U11084 (N_11084,N_10807,N_10786);
xnor U11085 (N_11085,N_10855,N_10925);
xor U11086 (N_11086,N_10841,N_10896);
or U11087 (N_11087,N_10814,N_10883);
nand U11088 (N_11088,N_10871,N_10831);
xnor U11089 (N_11089,N_10941,N_10893);
xor U11090 (N_11090,N_10937,N_10776);
nand U11091 (N_11091,N_10933,N_10803);
and U11092 (N_11092,N_10872,N_10911);
and U11093 (N_11093,N_10950,N_10860);
and U11094 (N_11094,N_10839,N_10822);
or U11095 (N_11095,N_10866,N_10768);
nand U11096 (N_11096,N_10763,N_10834);
or U11097 (N_11097,N_10949,N_10954);
or U11098 (N_11098,N_10832,N_10812);
nor U11099 (N_11099,N_10793,N_10789);
xor U11100 (N_11100,N_10761,N_10773);
nand U11101 (N_11101,N_10902,N_10804);
or U11102 (N_11102,N_10940,N_10772);
nor U11103 (N_11103,N_10884,N_10962);
nand U11104 (N_11104,N_10852,N_10964);
and U11105 (N_11105,N_10936,N_10930);
xnor U11106 (N_11106,N_10863,N_10821);
nand U11107 (N_11107,N_10985,N_10997);
nor U11108 (N_11108,N_10784,N_10971);
and U11109 (N_11109,N_10811,N_10984);
and U11110 (N_11110,N_10972,N_10760);
nand U11111 (N_11111,N_10824,N_10905);
nand U11112 (N_11112,N_10990,N_10813);
nor U11113 (N_11113,N_10869,N_10857);
nor U11114 (N_11114,N_10837,N_10838);
nor U11115 (N_11115,N_10862,N_10891);
and U11116 (N_11116,N_10938,N_10914);
xor U11117 (N_11117,N_10910,N_10816);
xor U11118 (N_11118,N_10974,N_10958);
and U11119 (N_11119,N_10864,N_10957);
nand U11120 (N_11120,N_10956,N_10877);
and U11121 (N_11121,N_10988,N_10751);
nand U11122 (N_11122,N_10847,N_10759);
xnor U11123 (N_11123,N_10802,N_10931);
nor U11124 (N_11124,N_10775,N_10815);
nor U11125 (N_11125,N_10888,N_10914);
or U11126 (N_11126,N_10882,N_10823);
xor U11127 (N_11127,N_10807,N_10949);
nor U11128 (N_11128,N_10907,N_10971);
xnor U11129 (N_11129,N_10792,N_10993);
or U11130 (N_11130,N_10988,N_10882);
or U11131 (N_11131,N_10945,N_10980);
xor U11132 (N_11132,N_10947,N_10858);
and U11133 (N_11133,N_10851,N_10760);
or U11134 (N_11134,N_10888,N_10968);
xor U11135 (N_11135,N_10830,N_10835);
nor U11136 (N_11136,N_10848,N_10925);
nor U11137 (N_11137,N_10835,N_10810);
nand U11138 (N_11138,N_10955,N_10942);
or U11139 (N_11139,N_10796,N_10881);
xor U11140 (N_11140,N_10963,N_10956);
and U11141 (N_11141,N_10776,N_10984);
and U11142 (N_11142,N_10830,N_10991);
and U11143 (N_11143,N_10990,N_10786);
and U11144 (N_11144,N_10966,N_10954);
xnor U11145 (N_11145,N_10752,N_10949);
nand U11146 (N_11146,N_10867,N_10820);
xor U11147 (N_11147,N_10781,N_10829);
or U11148 (N_11148,N_10773,N_10809);
and U11149 (N_11149,N_10937,N_10822);
xnor U11150 (N_11150,N_10914,N_10864);
xnor U11151 (N_11151,N_10783,N_10761);
xnor U11152 (N_11152,N_10787,N_10792);
and U11153 (N_11153,N_10858,N_10993);
nor U11154 (N_11154,N_10819,N_10822);
nand U11155 (N_11155,N_10983,N_10789);
nand U11156 (N_11156,N_10829,N_10889);
nand U11157 (N_11157,N_10806,N_10834);
and U11158 (N_11158,N_10849,N_10750);
nand U11159 (N_11159,N_10867,N_10924);
xnor U11160 (N_11160,N_10845,N_10902);
xnor U11161 (N_11161,N_10836,N_10763);
xnor U11162 (N_11162,N_10811,N_10875);
xor U11163 (N_11163,N_10867,N_10926);
xor U11164 (N_11164,N_10964,N_10966);
nand U11165 (N_11165,N_10946,N_10798);
nor U11166 (N_11166,N_10822,N_10885);
and U11167 (N_11167,N_10834,N_10835);
and U11168 (N_11168,N_10958,N_10790);
and U11169 (N_11169,N_10977,N_10810);
nand U11170 (N_11170,N_10996,N_10807);
and U11171 (N_11171,N_10846,N_10927);
xor U11172 (N_11172,N_10921,N_10996);
xnor U11173 (N_11173,N_10773,N_10894);
xor U11174 (N_11174,N_10866,N_10788);
nand U11175 (N_11175,N_10751,N_10959);
and U11176 (N_11176,N_10763,N_10824);
nand U11177 (N_11177,N_10782,N_10767);
and U11178 (N_11178,N_10888,N_10957);
and U11179 (N_11179,N_10857,N_10909);
xor U11180 (N_11180,N_10991,N_10842);
and U11181 (N_11181,N_10776,N_10958);
nand U11182 (N_11182,N_10988,N_10834);
nand U11183 (N_11183,N_10783,N_10919);
nand U11184 (N_11184,N_10939,N_10830);
nand U11185 (N_11185,N_10923,N_10818);
xnor U11186 (N_11186,N_10780,N_10773);
nor U11187 (N_11187,N_10910,N_10870);
nor U11188 (N_11188,N_10977,N_10875);
nor U11189 (N_11189,N_10940,N_10866);
and U11190 (N_11190,N_10813,N_10770);
nor U11191 (N_11191,N_10875,N_10819);
nor U11192 (N_11192,N_10872,N_10899);
nor U11193 (N_11193,N_10911,N_10897);
nor U11194 (N_11194,N_10921,N_10830);
xnor U11195 (N_11195,N_10846,N_10854);
and U11196 (N_11196,N_10864,N_10787);
nand U11197 (N_11197,N_10750,N_10760);
xnor U11198 (N_11198,N_10774,N_10914);
and U11199 (N_11199,N_10801,N_10997);
or U11200 (N_11200,N_10830,N_10818);
or U11201 (N_11201,N_10913,N_10827);
nor U11202 (N_11202,N_10793,N_10766);
or U11203 (N_11203,N_10782,N_10931);
or U11204 (N_11204,N_10843,N_10854);
and U11205 (N_11205,N_10908,N_10980);
and U11206 (N_11206,N_10983,N_10877);
nor U11207 (N_11207,N_10760,N_10804);
nor U11208 (N_11208,N_10903,N_10858);
xor U11209 (N_11209,N_10925,N_10868);
and U11210 (N_11210,N_10805,N_10901);
or U11211 (N_11211,N_10819,N_10797);
or U11212 (N_11212,N_10857,N_10880);
or U11213 (N_11213,N_10977,N_10772);
nand U11214 (N_11214,N_10760,N_10770);
nand U11215 (N_11215,N_10810,N_10862);
and U11216 (N_11216,N_10943,N_10950);
or U11217 (N_11217,N_10858,N_10899);
nand U11218 (N_11218,N_10950,N_10835);
nand U11219 (N_11219,N_10983,N_10917);
nor U11220 (N_11220,N_10900,N_10878);
nand U11221 (N_11221,N_10876,N_10903);
and U11222 (N_11222,N_10956,N_10827);
xnor U11223 (N_11223,N_10786,N_10936);
and U11224 (N_11224,N_10767,N_10969);
nand U11225 (N_11225,N_10806,N_10893);
nor U11226 (N_11226,N_10891,N_10900);
nand U11227 (N_11227,N_10992,N_10854);
nor U11228 (N_11228,N_10799,N_10800);
or U11229 (N_11229,N_10821,N_10804);
xnor U11230 (N_11230,N_10973,N_10920);
and U11231 (N_11231,N_10829,N_10980);
nor U11232 (N_11232,N_10759,N_10957);
xnor U11233 (N_11233,N_10866,N_10750);
and U11234 (N_11234,N_10835,N_10771);
or U11235 (N_11235,N_10897,N_10855);
and U11236 (N_11236,N_10783,N_10947);
or U11237 (N_11237,N_10905,N_10852);
xor U11238 (N_11238,N_10810,N_10971);
or U11239 (N_11239,N_10975,N_10892);
nor U11240 (N_11240,N_10823,N_10752);
nor U11241 (N_11241,N_10893,N_10998);
xor U11242 (N_11242,N_10781,N_10898);
or U11243 (N_11243,N_10974,N_10881);
xnor U11244 (N_11244,N_10755,N_10951);
nor U11245 (N_11245,N_10945,N_10878);
and U11246 (N_11246,N_10930,N_10858);
or U11247 (N_11247,N_10766,N_10977);
or U11248 (N_11248,N_10900,N_10775);
nand U11249 (N_11249,N_10958,N_10758);
nand U11250 (N_11250,N_11230,N_11117);
nand U11251 (N_11251,N_11052,N_11217);
and U11252 (N_11252,N_11008,N_11192);
nand U11253 (N_11253,N_11019,N_11003);
and U11254 (N_11254,N_11134,N_11059);
and U11255 (N_11255,N_11051,N_11076);
and U11256 (N_11256,N_11246,N_11058);
and U11257 (N_11257,N_11164,N_11079);
or U11258 (N_11258,N_11032,N_11185);
xnor U11259 (N_11259,N_11025,N_11173);
nor U11260 (N_11260,N_11114,N_11238);
and U11261 (N_11261,N_11021,N_11043);
xor U11262 (N_11262,N_11140,N_11099);
or U11263 (N_11263,N_11026,N_11163);
nor U11264 (N_11264,N_11147,N_11012);
nor U11265 (N_11265,N_11011,N_11017);
nand U11266 (N_11266,N_11207,N_11095);
and U11267 (N_11267,N_11063,N_11159);
nor U11268 (N_11268,N_11161,N_11139);
or U11269 (N_11269,N_11036,N_11202);
and U11270 (N_11270,N_11082,N_11240);
nor U11271 (N_11271,N_11123,N_11160);
xnor U11272 (N_11272,N_11199,N_11215);
or U11273 (N_11273,N_11141,N_11183);
nor U11274 (N_11274,N_11234,N_11085);
xnor U11275 (N_11275,N_11064,N_11239);
nor U11276 (N_11276,N_11006,N_11055);
or U11277 (N_11277,N_11062,N_11169);
xor U11278 (N_11278,N_11113,N_11096);
nor U11279 (N_11279,N_11050,N_11224);
nand U11280 (N_11280,N_11108,N_11195);
xor U11281 (N_11281,N_11177,N_11142);
nand U11282 (N_11282,N_11233,N_11110);
xnor U11283 (N_11283,N_11129,N_11150);
and U11284 (N_11284,N_11037,N_11024);
nor U11285 (N_11285,N_11124,N_11033);
xnor U11286 (N_11286,N_11188,N_11228);
and U11287 (N_11287,N_11198,N_11039);
or U11288 (N_11288,N_11148,N_11105);
nand U11289 (N_11289,N_11145,N_11023);
or U11290 (N_11290,N_11083,N_11162);
nor U11291 (N_11291,N_11004,N_11226);
nor U11292 (N_11292,N_11002,N_11181);
and U11293 (N_11293,N_11212,N_11216);
and U11294 (N_11294,N_11049,N_11102);
or U11295 (N_11295,N_11093,N_11107);
xnor U11296 (N_11296,N_11167,N_11081);
nand U11297 (N_11297,N_11087,N_11007);
or U11298 (N_11298,N_11047,N_11194);
xor U11299 (N_11299,N_11090,N_11205);
nand U11300 (N_11300,N_11018,N_11186);
nand U11301 (N_11301,N_11094,N_11061);
nor U11302 (N_11302,N_11133,N_11184);
or U11303 (N_11303,N_11190,N_11193);
or U11304 (N_11304,N_11080,N_11112);
xor U11305 (N_11305,N_11098,N_11213);
nor U11306 (N_11306,N_11241,N_11187);
xnor U11307 (N_11307,N_11221,N_11034);
nor U11308 (N_11308,N_11203,N_11040);
xnor U11309 (N_11309,N_11088,N_11211);
and U11310 (N_11310,N_11072,N_11128);
nand U11311 (N_11311,N_11138,N_11237);
or U11312 (N_11312,N_11172,N_11156);
nor U11313 (N_11313,N_11057,N_11120);
and U11314 (N_11314,N_11200,N_11014);
nor U11315 (N_11315,N_11009,N_11158);
or U11316 (N_11316,N_11231,N_11175);
or U11317 (N_11317,N_11097,N_11091);
and U11318 (N_11318,N_11191,N_11196);
xor U11319 (N_11319,N_11127,N_11044);
nand U11320 (N_11320,N_11001,N_11146);
or U11321 (N_11321,N_11243,N_11220);
xnor U11322 (N_11322,N_11125,N_11131);
and U11323 (N_11323,N_11029,N_11111);
or U11324 (N_11324,N_11078,N_11013);
and U11325 (N_11325,N_11104,N_11168);
and U11326 (N_11326,N_11242,N_11121);
xnor U11327 (N_11327,N_11101,N_11130);
or U11328 (N_11328,N_11126,N_11042);
xnor U11329 (N_11329,N_11074,N_11070);
xor U11330 (N_11330,N_11092,N_11236);
nor U11331 (N_11331,N_11000,N_11119);
nor U11332 (N_11332,N_11046,N_11149);
or U11333 (N_11333,N_11218,N_11115);
nand U11334 (N_11334,N_11045,N_11075);
and U11335 (N_11335,N_11077,N_11144);
xnor U11336 (N_11336,N_11068,N_11084);
xnor U11337 (N_11337,N_11152,N_11176);
nand U11338 (N_11338,N_11151,N_11005);
xnor U11339 (N_11339,N_11219,N_11071);
xnor U11340 (N_11340,N_11030,N_11031);
xor U11341 (N_11341,N_11015,N_11041);
and U11342 (N_11342,N_11229,N_11214);
xor U11343 (N_11343,N_11106,N_11225);
nor U11344 (N_11344,N_11054,N_11206);
and U11345 (N_11345,N_11065,N_11069);
nor U11346 (N_11346,N_11089,N_11244);
nor U11347 (N_11347,N_11100,N_11201);
nand U11348 (N_11348,N_11245,N_11155);
and U11349 (N_11349,N_11248,N_11016);
and U11350 (N_11350,N_11235,N_11022);
nor U11351 (N_11351,N_11182,N_11189);
nor U11352 (N_11352,N_11053,N_11027);
xnor U11353 (N_11353,N_11086,N_11143);
nor U11354 (N_11354,N_11048,N_11171);
or U11355 (N_11355,N_11180,N_11122);
nand U11356 (N_11356,N_11067,N_11208);
nor U11357 (N_11357,N_11179,N_11247);
xnor U11358 (N_11358,N_11010,N_11056);
nor U11359 (N_11359,N_11165,N_11109);
nor U11360 (N_11360,N_11210,N_11222);
xor U11361 (N_11361,N_11157,N_11116);
nor U11362 (N_11362,N_11204,N_11132);
nor U11363 (N_11363,N_11223,N_11035);
and U11364 (N_11364,N_11197,N_11170);
nor U11365 (N_11365,N_11232,N_11174);
or U11366 (N_11366,N_11178,N_11154);
xnor U11367 (N_11367,N_11136,N_11135);
nor U11368 (N_11368,N_11103,N_11118);
and U11369 (N_11369,N_11066,N_11073);
xor U11370 (N_11370,N_11249,N_11227);
or U11371 (N_11371,N_11137,N_11153);
or U11372 (N_11372,N_11028,N_11060);
and U11373 (N_11373,N_11166,N_11038);
nor U11374 (N_11374,N_11209,N_11020);
or U11375 (N_11375,N_11222,N_11118);
and U11376 (N_11376,N_11105,N_11104);
xor U11377 (N_11377,N_11186,N_11236);
nor U11378 (N_11378,N_11079,N_11048);
nor U11379 (N_11379,N_11119,N_11220);
nand U11380 (N_11380,N_11038,N_11049);
nand U11381 (N_11381,N_11005,N_11135);
nor U11382 (N_11382,N_11170,N_11225);
nand U11383 (N_11383,N_11214,N_11143);
xor U11384 (N_11384,N_11040,N_11244);
or U11385 (N_11385,N_11217,N_11028);
and U11386 (N_11386,N_11143,N_11072);
or U11387 (N_11387,N_11247,N_11181);
and U11388 (N_11388,N_11079,N_11180);
nand U11389 (N_11389,N_11163,N_11228);
and U11390 (N_11390,N_11055,N_11225);
nand U11391 (N_11391,N_11015,N_11134);
xnor U11392 (N_11392,N_11048,N_11006);
nand U11393 (N_11393,N_11238,N_11240);
nor U11394 (N_11394,N_11153,N_11071);
xor U11395 (N_11395,N_11065,N_11202);
xnor U11396 (N_11396,N_11036,N_11245);
and U11397 (N_11397,N_11033,N_11067);
or U11398 (N_11398,N_11169,N_11113);
nor U11399 (N_11399,N_11121,N_11168);
or U11400 (N_11400,N_11079,N_11158);
nor U11401 (N_11401,N_11078,N_11092);
or U11402 (N_11402,N_11072,N_11090);
nand U11403 (N_11403,N_11102,N_11197);
nor U11404 (N_11404,N_11089,N_11079);
and U11405 (N_11405,N_11126,N_11137);
or U11406 (N_11406,N_11209,N_11234);
nor U11407 (N_11407,N_11188,N_11200);
nor U11408 (N_11408,N_11198,N_11052);
and U11409 (N_11409,N_11198,N_11030);
nor U11410 (N_11410,N_11181,N_11115);
nand U11411 (N_11411,N_11111,N_11241);
xor U11412 (N_11412,N_11113,N_11035);
xnor U11413 (N_11413,N_11120,N_11060);
nand U11414 (N_11414,N_11220,N_11160);
xnor U11415 (N_11415,N_11214,N_11171);
xor U11416 (N_11416,N_11244,N_11134);
and U11417 (N_11417,N_11086,N_11007);
nor U11418 (N_11418,N_11010,N_11050);
and U11419 (N_11419,N_11121,N_11195);
nand U11420 (N_11420,N_11185,N_11050);
nor U11421 (N_11421,N_11118,N_11053);
nand U11422 (N_11422,N_11168,N_11053);
or U11423 (N_11423,N_11069,N_11212);
and U11424 (N_11424,N_11072,N_11189);
and U11425 (N_11425,N_11186,N_11076);
or U11426 (N_11426,N_11106,N_11058);
nand U11427 (N_11427,N_11116,N_11214);
nand U11428 (N_11428,N_11113,N_11043);
nand U11429 (N_11429,N_11021,N_11003);
nor U11430 (N_11430,N_11187,N_11022);
nand U11431 (N_11431,N_11185,N_11119);
nand U11432 (N_11432,N_11030,N_11117);
xnor U11433 (N_11433,N_11244,N_11202);
nor U11434 (N_11434,N_11064,N_11246);
nand U11435 (N_11435,N_11237,N_11108);
xor U11436 (N_11436,N_11148,N_11109);
or U11437 (N_11437,N_11168,N_11092);
or U11438 (N_11438,N_11230,N_11139);
nand U11439 (N_11439,N_11129,N_11002);
nor U11440 (N_11440,N_11126,N_11221);
xnor U11441 (N_11441,N_11204,N_11040);
nor U11442 (N_11442,N_11111,N_11000);
nor U11443 (N_11443,N_11019,N_11181);
nand U11444 (N_11444,N_11015,N_11096);
nor U11445 (N_11445,N_11197,N_11149);
nor U11446 (N_11446,N_11193,N_11128);
or U11447 (N_11447,N_11202,N_11173);
nor U11448 (N_11448,N_11158,N_11108);
or U11449 (N_11449,N_11039,N_11229);
and U11450 (N_11450,N_11221,N_11042);
nor U11451 (N_11451,N_11041,N_11052);
nand U11452 (N_11452,N_11087,N_11131);
and U11453 (N_11453,N_11210,N_11204);
nor U11454 (N_11454,N_11052,N_11188);
nor U11455 (N_11455,N_11038,N_11100);
and U11456 (N_11456,N_11133,N_11099);
nor U11457 (N_11457,N_11223,N_11099);
or U11458 (N_11458,N_11026,N_11102);
and U11459 (N_11459,N_11099,N_11176);
and U11460 (N_11460,N_11171,N_11123);
xnor U11461 (N_11461,N_11120,N_11064);
nand U11462 (N_11462,N_11144,N_11082);
nand U11463 (N_11463,N_11054,N_11039);
and U11464 (N_11464,N_11170,N_11059);
nand U11465 (N_11465,N_11123,N_11241);
nand U11466 (N_11466,N_11198,N_11076);
nor U11467 (N_11467,N_11192,N_11101);
nor U11468 (N_11468,N_11232,N_11059);
nand U11469 (N_11469,N_11216,N_11073);
and U11470 (N_11470,N_11095,N_11150);
nand U11471 (N_11471,N_11129,N_11201);
nor U11472 (N_11472,N_11121,N_11170);
xor U11473 (N_11473,N_11061,N_11229);
nand U11474 (N_11474,N_11056,N_11162);
nand U11475 (N_11475,N_11156,N_11192);
or U11476 (N_11476,N_11102,N_11235);
or U11477 (N_11477,N_11077,N_11171);
nand U11478 (N_11478,N_11238,N_11092);
and U11479 (N_11479,N_11186,N_11022);
or U11480 (N_11480,N_11125,N_11146);
nand U11481 (N_11481,N_11093,N_11083);
or U11482 (N_11482,N_11115,N_11201);
or U11483 (N_11483,N_11127,N_11075);
or U11484 (N_11484,N_11046,N_11204);
xnor U11485 (N_11485,N_11048,N_11128);
nor U11486 (N_11486,N_11087,N_11228);
nor U11487 (N_11487,N_11087,N_11160);
and U11488 (N_11488,N_11019,N_11066);
nand U11489 (N_11489,N_11081,N_11050);
nor U11490 (N_11490,N_11052,N_11189);
xor U11491 (N_11491,N_11190,N_11069);
nand U11492 (N_11492,N_11243,N_11150);
xor U11493 (N_11493,N_11002,N_11176);
xor U11494 (N_11494,N_11114,N_11203);
and U11495 (N_11495,N_11104,N_11154);
nor U11496 (N_11496,N_11196,N_11167);
xnor U11497 (N_11497,N_11214,N_11164);
nor U11498 (N_11498,N_11236,N_11045);
and U11499 (N_11499,N_11043,N_11057);
xor U11500 (N_11500,N_11401,N_11441);
nand U11501 (N_11501,N_11464,N_11412);
and U11502 (N_11502,N_11272,N_11348);
or U11503 (N_11503,N_11434,N_11334);
or U11504 (N_11504,N_11450,N_11446);
nand U11505 (N_11505,N_11492,N_11495);
xor U11506 (N_11506,N_11268,N_11435);
nand U11507 (N_11507,N_11312,N_11380);
and U11508 (N_11508,N_11447,N_11389);
or U11509 (N_11509,N_11384,N_11275);
xnor U11510 (N_11510,N_11433,N_11449);
and U11511 (N_11511,N_11487,N_11358);
and U11512 (N_11512,N_11440,N_11349);
nor U11513 (N_11513,N_11338,N_11354);
nand U11514 (N_11514,N_11273,N_11254);
nand U11515 (N_11515,N_11282,N_11372);
and U11516 (N_11516,N_11451,N_11415);
nor U11517 (N_11517,N_11497,N_11267);
nand U11518 (N_11518,N_11473,N_11363);
xnor U11519 (N_11519,N_11336,N_11365);
nand U11520 (N_11520,N_11416,N_11394);
and U11521 (N_11521,N_11253,N_11430);
xnor U11522 (N_11522,N_11343,N_11357);
and U11523 (N_11523,N_11321,N_11340);
nor U11524 (N_11524,N_11327,N_11477);
or U11525 (N_11525,N_11499,N_11310);
or U11526 (N_11526,N_11454,N_11437);
or U11527 (N_11527,N_11373,N_11261);
nand U11528 (N_11528,N_11291,N_11298);
xor U11529 (N_11529,N_11421,N_11364);
nor U11530 (N_11530,N_11426,N_11342);
or U11531 (N_11531,N_11279,N_11257);
nand U11532 (N_11532,N_11323,N_11324);
and U11533 (N_11533,N_11470,N_11370);
and U11534 (N_11534,N_11475,N_11280);
and U11535 (N_11535,N_11431,N_11306);
or U11536 (N_11536,N_11453,N_11406);
nor U11537 (N_11537,N_11423,N_11381);
and U11538 (N_11538,N_11307,N_11424);
nand U11539 (N_11539,N_11420,N_11258);
or U11540 (N_11540,N_11395,N_11445);
xor U11541 (N_11541,N_11404,N_11271);
xnor U11542 (N_11542,N_11391,N_11469);
nor U11543 (N_11543,N_11317,N_11320);
or U11544 (N_11544,N_11376,N_11480);
xnor U11545 (N_11545,N_11374,N_11403);
nor U11546 (N_11546,N_11304,N_11408);
nor U11547 (N_11547,N_11368,N_11297);
or U11548 (N_11548,N_11344,N_11333);
and U11549 (N_11549,N_11439,N_11418);
nor U11550 (N_11550,N_11377,N_11493);
nor U11551 (N_11551,N_11322,N_11300);
nand U11552 (N_11552,N_11484,N_11331);
nor U11553 (N_11553,N_11432,N_11386);
xor U11554 (N_11554,N_11417,N_11498);
and U11555 (N_11555,N_11491,N_11255);
xnor U11556 (N_11556,N_11335,N_11330);
and U11557 (N_11557,N_11325,N_11438);
nand U11558 (N_11558,N_11353,N_11339);
and U11559 (N_11559,N_11296,N_11371);
nand U11560 (N_11560,N_11458,N_11251);
nor U11561 (N_11561,N_11410,N_11481);
xor U11562 (N_11562,N_11276,N_11465);
nor U11563 (N_11563,N_11337,N_11318);
xnor U11564 (N_11564,N_11482,N_11490);
nand U11565 (N_11565,N_11341,N_11387);
nand U11566 (N_11566,N_11382,N_11379);
and U11567 (N_11567,N_11313,N_11428);
and U11568 (N_11568,N_11478,N_11274);
nor U11569 (N_11569,N_11488,N_11355);
nand U11570 (N_11570,N_11471,N_11396);
nand U11571 (N_11571,N_11350,N_11311);
nor U11572 (N_11572,N_11463,N_11278);
xor U11573 (N_11573,N_11346,N_11448);
or U11574 (N_11574,N_11444,N_11486);
nor U11575 (N_11575,N_11294,N_11316);
xnor U11576 (N_11576,N_11356,N_11496);
nand U11577 (N_11577,N_11263,N_11411);
xnor U11578 (N_11578,N_11460,N_11302);
or U11579 (N_11579,N_11351,N_11256);
nand U11580 (N_11580,N_11284,N_11378);
and U11581 (N_11581,N_11277,N_11369);
or U11582 (N_11582,N_11398,N_11301);
and U11583 (N_11583,N_11436,N_11328);
or U11584 (N_11584,N_11388,N_11283);
and U11585 (N_11585,N_11452,N_11375);
and U11586 (N_11586,N_11314,N_11390);
nand U11587 (N_11587,N_11457,N_11414);
nor U11588 (N_11588,N_11329,N_11269);
xnor U11589 (N_11589,N_11494,N_11285);
nand U11590 (N_11590,N_11270,N_11466);
nand U11591 (N_11591,N_11286,N_11472);
or U11592 (N_11592,N_11459,N_11289);
and U11593 (N_11593,N_11303,N_11299);
and U11594 (N_11594,N_11399,N_11397);
or U11595 (N_11595,N_11308,N_11326);
nand U11596 (N_11596,N_11467,N_11315);
and U11597 (N_11597,N_11292,N_11405);
nor U11598 (N_11598,N_11392,N_11468);
xnor U11599 (N_11599,N_11345,N_11383);
nand U11600 (N_11600,N_11360,N_11385);
nand U11601 (N_11601,N_11309,N_11367);
or U11602 (N_11602,N_11455,N_11264);
or U11603 (N_11603,N_11402,N_11352);
xnor U11604 (N_11604,N_11347,N_11474);
and U11605 (N_11605,N_11462,N_11295);
and U11606 (N_11606,N_11250,N_11425);
xnor U11607 (N_11607,N_11476,N_11266);
xnor U11608 (N_11608,N_11332,N_11422);
xnor U11609 (N_11609,N_11479,N_11259);
nand U11610 (N_11610,N_11400,N_11413);
or U11611 (N_11611,N_11489,N_11442);
nand U11612 (N_11612,N_11265,N_11485);
nor U11613 (N_11613,N_11359,N_11419);
or U11614 (N_11614,N_11456,N_11461);
and U11615 (N_11615,N_11287,N_11305);
nor U11616 (N_11616,N_11288,N_11293);
and U11617 (N_11617,N_11443,N_11483);
or U11618 (N_11618,N_11429,N_11409);
nand U11619 (N_11619,N_11362,N_11427);
nand U11620 (N_11620,N_11319,N_11252);
and U11621 (N_11621,N_11290,N_11262);
nor U11622 (N_11622,N_11407,N_11361);
and U11623 (N_11623,N_11393,N_11260);
and U11624 (N_11624,N_11281,N_11366);
nand U11625 (N_11625,N_11416,N_11268);
or U11626 (N_11626,N_11280,N_11422);
xnor U11627 (N_11627,N_11493,N_11266);
nand U11628 (N_11628,N_11357,N_11478);
or U11629 (N_11629,N_11293,N_11330);
nand U11630 (N_11630,N_11264,N_11346);
xor U11631 (N_11631,N_11466,N_11382);
nand U11632 (N_11632,N_11432,N_11339);
nand U11633 (N_11633,N_11303,N_11267);
xor U11634 (N_11634,N_11360,N_11318);
xnor U11635 (N_11635,N_11450,N_11301);
and U11636 (N_11636,N_11359,N_11444);
and U11637 (N_11637,N_11489,N_11418);
nor U11638 (N_11638,N_11353,N_11275);
and U11639 (N_11639,N_11294,N_11355);
xor U11640 (N_11640,N_11317,N_11440);
or U11641 (N_11641,N_11489,N_11322);
nand U11642 (N_11642,N_11250,N_11306);
nand U11643 (N_11643,N_11377,N_11296);
xor U11644 (N_11644,N_11461,N_11487);
nor U11645 (N_11645,N_11258,N_11346);
nand U11646 (N_11646,N_11309,N_11478);
xor U11647 (N_11647,N_11447,N_11450);
nand U11648 (N_11648,N_11342,N_11394);
xnor U11649 (N_11649,N_11296,N_11427);
nor U11650 (N_11650,N_11473,N_11377);
or U11651 (N_11651,N_11360,N_11461);
or U11652 (N_11652,N_11290,N_11475);
or U11653 (N_11653,N_11320,N_11403);
nand U11654 (N_11654,N_11252,N_11351);
or U11655 (N_11655,N_11454,N_11389);
nand U11656 (N_11656,N_11297,N_11447);
or U11657 (N_11657,N_11292,N_11484);
and U11658 (N_11658,N_11481,N_11490);
xnor U11659 (N_11659,N_11373,N_11311);
xor U11660 (N_11660,N_11401,N_11428);
and U11661 (N_11661,N_11434,N_11480);
and U11662 (N_11662,N_11463,N_11348);
and U11663 (N_11663,N_11424,N_11403);
nor U11664 (N_11664,N_11483,N_11313);
xor U11665 (N_11665,N_11261,N_11332);
nor U11666 (N_11666,N_11384,N_11496);
and U11667 (N_11667,N_11328,N_11420);
nor U11668 (N_11668,N_11409,N_11425);
nor U11669 (N_11669,N_11267,N_11332);
or U11670 (N_11670,N_11357,N_11327);
nand U11671 (N_11671,N_11314,N_11274);
nor U11672 (N_11672,N_11433,N_11382);
or U11673 (N_11673,N_11438,N_11297);
or U11674 (N_11674,N_11365,N_11383);
and U11675 (N_11675,N_11319,N_11378);
nor U11676 (N_11676,N_11432,N_11337);
and U11677 (N_11677,N_11426,N_11347);
xnor U11678 (N_11678,N_11454,N_11488);
xor U11679 (N_11679,N_11428,N_11379);
or U11680 (N_11680,N_11294,N_11468);
nor U11681 (N_11681,N_11453,N_11345);
xor U11682 (N_11682,N_11273,N_11348);
xnor U11683 (N_11683,N_11454,N_11411);
or U11684 (N_11684,N_11265,N_11443);
and U11685 (N_11685,N_11330,N_11403);
nor U11686 (N_11686,N_11475,N_11303);
nand U11687 (N_11687,N_11414,N_11469);
nand U11688 (N_11688,N_11337,N_11397);
xnor U11689 (N_11689,N_11310,N_11485);
and U11690 (N_11690,N_11370,N_11430);
or U11691 (N_11691,N_11310,N_11261);
or U11692 (N_11692,N_11413,N_11316);
xor U11693 (N_11693,N_11408,N_11303);
nand U11694 (N_11694,N_11334,N_11481);
xnor U11695 (N_11695,N_11491,N_11429);
or U11696 (N_11696,N_11460,N_11264);
and U11697 (N_11697,N_11357,N_11313);
nor U11698 (N_11698,N_11349,N_11341);
and U11699 (N_11699,N_11297,N_11401);
nand U11700 (N_11700,N_11313,N_11307);
or U11701 (N_11701,N_11273,N_11377);
nor U11702 (N_11702,N_11455,N_11284);
nand U11703 (N_11703,N_11479,N_11466);
nor U11704 (N_11704,N_11486,N_11287);
or U11705 (N_11705,N_11343,N_11282);
xor U11706 (N_11706,N_11349,N_11276);
nand U11707 (N_11707,N_11407,N_11386);
xor U11708 (N_11708,N_11401,N_11426);
and U11709 (N_11709,N_11325,N_11268);
nor U11710 (N_11710,N_11443,N_11399);
or U11711 (N_11711,N_11275,N_11413);
nor U11712 (N_11712,N_11372,N_11375);
or U11713 (N_11713,N_11343,N_11488);
or U11714 (N_11714,N_11451,N_11396);
and U11715 (N_11715,N_11497,N_11380);
nor U11716 (N_11716,N_11474,N_11468);
nand U11717 (N_11717,N_11277,N_11269);
or U11718 (N_11718,N_11272,N_11356);
and U11719 (N_11719,N_11474,N_11423);
and U11720 (N_11720,N_11416,N_11495);
or U11721 (N_11721,N_11436,N_11350);
nand U11722 (N_11722,N_11380,N_11313);
xor U11723 (N_11723,N_11262,N_11353);
xnor U11724 (N_11724,N_11448,N_11357);
nand U11725 (N_11725,N_11466,N_11423);
nand U11726 (N_11726,N_11375,N_11382);
and U11727 (N_11727,N_11492,N_11416);
nor U11728 (N_11728,N_11338,N_11401);
xnor U11729 (N_11729,N_11382,N_11384);
xor U11730 (N_11730,N_11314,N_11252);
or U11731 (N_11731,N_11311,N_11392);
xor U11732 (N_11732,N_11267,N_11384);
nor U11733 (N_11733,N_11333,N_11337);
or U11734 (N_11734,N_11419,N_11477);
and U11735 (N_11735,N_11303,N_11427);
nor U11736 (N_11736,N_11364,N_11256);
or U11737 (N_11737,N_11302,N_11462);
nor U11738 (N_11738,N_11492,N_11479);
and U11739 (N_11739,N_11388,N_11290);
nor U11740 (N_11740,N_11281,N_11258);
nand U11741 (N_11741,N_11340,N_11293);
or U11742 (N_11742,N_11336,N_11327);
xor U11743 (N_11743,N_11325,N_11477);
xor U11744 (N_11744,N_11319,N_11315);
nand U11745 (N_11745,N_11326,N_11426);
nor U11746 (N_11746,N_11361,N_11455);
or U11747 (N_11747,N_11344,N_11471);
and U11748 (N_11748,N_11282,N_11263);
or U11749 (N_11749,N_11429,N_11455);
and U11750 (N_11750,N_11632,N_11594);
xnor U11751 (N_11751,N_11748,N_11580);
nand U11752 (N_11752,N_11615,N_11633);
and U11753 (N_11753,N_11686,N_11502);
xor U11754 (N_11754,N_11742,N_11567);
nor U11755 (N_11755,N_11735,N_11500);
nand U11756 (N_11756,N_11668,N_11576);
or U11757 (N_11757,N_11690,N_11639);
and U11758 (N_11758,N_11643,N_11609);
and U11759 (N_11759,N_11699,N_11739);
xor U11760 (N_11760,N_11610,N_11710);
nor U11761 (N_11761,N_11661,N_11571);
or U11762 (N_11762,N_11674,N_11600);
and U11763 (N_11763,N_11722,N_11716);
or U11764 (N_11764,N_11707,N_11520);
nand U11765 (N_11765,N_11590,N_11582);
xor U11766 (N_11766,N_11721,N_11746);
nor U11767 (N_11767,N_11676,N_11630);
and U11768 (N_11768,N_11635,N_11522);
and U11769 (N_11769,N_11715,N_11547);
nor U11770 (N_11770,N_11568,N_11551);
nand U11771 (N_11771,N_11507,N_11664);
nand U11772 (N_11772,N_11538,N_11548);
or U11773 (N_11773,N_11618,N_11526);
nand U11774 (N_11774,N_11670,N_11720);
nor U11775 (N_11775,N_11585,N_11569);
xnor U11776 (N_11776,N_11671,N_11693);
nand U11777 (N_11777,N_11588,N_11577);
nand U11778 (N_11778,N_11684,N_11705);
and U11779 (N_11779,N_11613,N_11692);
nor U11780 (N_11780,N_11597,N_11599);
nor U11781 (N_11781,N_11659,N_11738);
xor U11782 (N_11782,N_11648,N_11589);
and U11783 (N_11783,N_11637,N_11730);
xnor U11784 (N_11784,N_11719,N_11662);
nor U11785 (N_11785,N_11549,N_11640);
nand U11786 (N_11786,N_11687,N_11681);
nor U11787 (N_11787,N_11697,N_11559);
and U11788 (N_11788,N_11679,N_11701);
nand U11789 (N_11789,N_11745,N_11677);
or U11790 (N_11790,N_11698,N_11629);
xor U11791 (N_11791,N_11656,N_11503);
nand U11792 (N_11792,N_11654,N_11660);
nor U11793 (N_11793,N_11527,N_11572);
xor U11794 (N_11794,N_11657,N_11561);
nand U11795 (N_11795,N_11505,N_11624);
nor U11796 (N_11796,N_11734,N_11712);
nor U11797 (N_11797,N_11528,N_11563);
and U11798 (N_11798,N_11510,N_11573);
xor U11799 (N_11799,N_11592,N_11553);
xnor U11800 (N_11800,N_11675,N_11727);
and U11801 (N_11801,N_11516,N_11606);
nor U11802 (N_11802,N_11669,N_11509);
and U11803 (N_11803,N_11542,N_11519);
nor U11804 (N_11804,N_11608,N_11747);
or U11805 (N_11805,N_11565,N_11733);
or U11806 (N_11806,N_11541,N_11560);
nand U11807 (N_11807,N_11501,N_11703);
xnor U11808 (N_11808,N_11512,N_11546);
xnor U11809 (N_11809,N_11605,N_11696);
nand U11810 (N_11810,N_11658,N_11612);
nor U11811 (N_11811,N_11614,N_11749);
and U11812 (N_11812,N_11566,N_11685);
xor U11813 (N_11813,N_11530,N_11517);
nand U11814 (N_11814,N_11673,N_11623);
and U11815 (N_11815,N_11591,N_11544);
xor U11816 (N_11816,N_11653,N_11650);
or U11817 (N_11817,N_11732,N_11557);
and U11818 (N_11818,N_11678,N_11700);
xnor U11819 (N_11819,N_11578,N_11575);
or U11820 (N_11820,N_11718,N_11593);
nand U11821 (N_11821,N_11598,N_11724);
nor U11822 (N_11822,N_11731,N_11555);
or U11823 (N_11823,N_11634,N_11627);
nand U11824 (N_11824,N_11611,N_11725);
nor U11825 (N_11825,N_11655,N_11583);
and U11826 (N_11826,N_11711,N_11694);
nor U11827 (N_11827,N_11683,N_11704);
xor U11828 (N_11828,N_11743,N_11601);
nand U11829 (N_11829,N_11619,N_11642);
or U11830 (N_11830,N_11728,N_11532);
or U11831 (N_11831,N_11558,N_11562);
or U11832 (N_11832,N_11645,N_11666);
nor U11833 (N_11833,N_11688,N_11596);
and U11834 (N_11834,N_11550,N_11570);
xor U11835 (N_11835,N_11511,N_11523);
or U11836 (N_11836,N_11514,N_11531);
nor U11837 (N_11837,N_11604,N_11741);
and U11838 (N_11838,N_11536,N_11525);
or U11839 (N_11839,N_11702,N_11652);
or U11840 (N_11840,N_11672,N_11628);
nand U11841 (N_11841,N_11641,N_11524);
nand U11842 (N_11842,N_11506,N_11513);
xnor U11843 (N_11843,N_11744,N_11736);
or U11844 (N_11844,N_11706,N_11626);
xnor U11845 (N_11845,N_11584,N_11587);
or U11846 (N_11846,N_11621,N_11545);
nand U11847 (N_11847,N_11717,N_11726);
and U11848 (N_11848,N_11616,N_11554);
nor U11849 (N_11849,N_11595,N_11665);
nor U11850 (N_11850,N_11708,N_11689);
xor U11851 (N_11851,N_11740,N_11508);
nand U11852 (N_11852,N_11713,N_11714);
and U11853 (N_11853,N_11607,N_11521);
and U11854 (N_11854,N_11540,N_11518);
or U11855 (N_11855,N_11556,N_11667);
nand U11856 (N_11856,N_11533,N_11603);
and U11857 (N_11857,N_11620,N_11504);
and U11858 (N_11858,N_11602,N_11638);
or U11859 (N_11859,N_11695,N_11539);
nand U11860 (N_11860,N_11574,N_11586);
or U11861 (N_11861,N_11564,N_11691);
nor U11862 (N_11862,N_11663,N_11631);
nand U11863 (N_11863,N_11649,N_11625);
or U11864 (N_11864,N_11617,N_11581);
xor U11865 (N_11865,N_11543,N_11682);
nand U11866 (N_11866,N_11529,N_11579);
xnor U11867 (N_11867,N_11729,N_11709);
nand U11868 (N_11868,N_11636,N_11622);
xor U11869 (N_11869,N_11644,N_11534);
or U11870 (N_11870,N_11651,N_11535);
xnor U11871 (N_11871,N_11680,N_11723);
xnor U11872 (N_11872,N_11537,N_11647);
nor U11873 (N_11873,N_11646,N_11515);
and U11874 (N_11874,N_11737,N_11552);
or U11875 (N_11875,N_11574,N_11511);
xnor U11876 (N_11876,N_11668,N_11714);
xnor U11877 (N_11877,N_11682,N_11692);
xor U11878 (N_11878,N_11749,N_11531);
nand U11879 (N_11879,N_11535,N_11632);
nand U11880 (N_11880,N_11622,N_11682);
and U11881 (N_11881,N_11666,N_11722);
nor U11882 (N_11882,N_11562,N_11665);
or U11883 (N_11883,N_11603,N_11559);
nor U11884 (N_11884,N_11657,N_11731);
or U11885 (N_11885,N_11714,N_11685);
xnor U11886 (N_11886,N_11643,N_11618);
or U11887 (N_11887,N_11606,N_11508);
or U11888 (N_11888,N_11696,N_11531);
nor U11889 (N_11889,N_11557,N_11538);
and U11890 (N_11890,N_11715,N_11746);
nor U11891 (N_11891,N_11567,N_11552);
and U11892 (N_11892,N_11565,N_11734);
nand U11893 (N_11893,N_11553,N_11600);
nor U11894 (N_11894,N_11723,N_11707);
xnor U11895 (N_11895,N_11533,N_11571);
nand U11896 (N_11896,N_11585,N_11713);
or U11897 (N_11897,N_11506,N_11640);
nor U11898 (N_11898,N_11503,N_11575);
and U11899 (N_11899,N_11748,N_11724);
nor U11900 (N_11900,N_11690,N_11702);
nand U11901 (N_11901,N_11711,N_11712);
and U11902 (N_11902,N_11564,N_11622);
nand U11903 (N_11903,N_11576,N_11718);
or U11904 (N_11904,N_11504,N_11741);
and U11905 (N_11905,N_11522,N_11746);
nor U11906 (N_11906,N_11668,N_11558);
xor U11907 (N_11907,N_11726,N_11515);
and U11908 (N_11908,N_11671,N_11591);
or U11909 (N_11909,N_11615,N_11723);
nor U11910 (N_11910,N_11606,N_11511);
nand U11911 (N_11911,N_11538,N_11716);
or U11912 (N_11912,N_11572,N_11519);
xor U11913 (N_11913,N_11608,N_11576);
xor U11914 (N_11914,N_11602,N_11731);
and U11915 (N_11915,N_11668,N_11632);
nor U11916 (N_11916,N_11624,N_11575);
and U11917 (N_11917,N_11726,N_11678);
nor U11918 (N_11918,N_11629,N_11562);
nor U11919 (N_11919,N_11647,N_11519);
or U11920 (N_11920,N_11746,N_11612);
or U11921 (N_11921,N_11569,N_11529);
or U11922 (N_11922,N_11552,N_11649);
and U11923 (N_11923,N_11732,N_11689);
or U11924 (N_11924,N_11722,N_11522);
xor U11925 (N_11925,N_11569,N_11543);
xnor U11926 (N_11926,N_11667,N_11640);
nand U11927 (N_11927,N_11714,N_11575);
nand U11928 (N_11928,N_11733,N_11626);
or U11929 (N_11929,N_11619,N_11675);
and U11930 (N_11930,N_11682,N_11646);
or U11931 (N_11931,N_11693,N_11638);
xnor U11932 (N_11932,N_11585,N_11556);
and U11933 (N_11933,N_11666,N_11512);
or U11934 (N_11934,N_11678,N_11613);
xor U11935 (N_11935,N_11706,N_11643);
or U11936 (N_11936,N_11524,N_11630);
nor U11937 (N_11937,N_11564,N_11696);
or U11938 (N_11938,N_11650,N_11708);
or U11939 (N_11939,N_11643,N_11563);
or U11940 (N_11940,N_11640,N_11588);
or U11941 (N_11941,N_11713,N_11610);
or U11942 (N_11942,N_11569,N_11527);
and U11943 (N_11943,N_11683,N_11533);
and U11944 (N_11944,N_11747,N_11560);
nand U11945 (N_11945,N_11692,N_11596);
and U11946 (N_11946,N_11712,N_11614);
xnor U11947 (N_11947,N_11746,N_11652);
nand U11948 (N_11948,N_11680,N_11554);
nand U11949 (N_11949,N_11688,N_11605);
and U11950 (N_11950,N_11578,N_11652);
xor U11951 (N_11951,N_11603,N_11690);
or U11952 (N_11952,N_11506,N_11673);
nor U11953 (N_11953,N_11660,N_11665);
and U11954 (N_11954,N_11511,N_11636);
xor U11955 (N_11955,N_11726,N_11554);
xnor U11956 (N_11956,N_11640,N_11673);
nand U11957 (N_11957,N_11574,N_11680);
or U11958 (N_11958,N_11651,N_11567);
or U11959 (N_11959,N_11565,N_11538);
nand U11960 (N_11960,N_11511,N_11562);
and U11961 (N_11961,N_11591,N_11532);
and U11962 (N_11962,N_11518,N_11565);
nor U11963 (N_11963,N_11568,N_11734);
xor U11964 (N_11964,N_11724,N_11658);
and U11965 (N_11965,N_11657,N_11694);
nand U11966 (N_11966,N_11608,N_11659);
or U11967 (N_11967,N_11655,N_11596);
nor U11968 (N_11968,N_11602,N_11627);
nor U11969 (N_11969,N_11538,N_11568);
nor U11970 (N_11970,N_11745,N_11511);
xnor U11971 (N_11971,N_11672,N_11747);
nand U11972 (N_11972,N_11537,N_11653);
and U11973 (N_11973,N_11657,N_11668);
xor U11974 (N_11974,N_11634,N_11671);
or U11975 (N_11975,N_11555,N_11620);
xor U11976 (N_11976,N_11704,N_11741);
xnor U11977 (N_11977,N_11598,N_11635);
or U11978 (N_11978,N_11615,N_11631);
and U11979 (N_11979,N_11560,N_11513);
xnor U11980 (N_11980,N_11594,N_11515);
xor U11981 (N_11981,N_11551,N_11630);
or U11982 (N_11982,N_11537,N_11628);
nor U11983 (N_11983,N_11575,N_11744);
or U11984 (N_11984,N_11606,N_11527);
nand U11985 (N_11985,N_11522,N_11578);
nand U11986 (N_11986,N_11646,N_11617);
xor U11987 (N_11987,N_11557,N_11718);
and U11988 (N_11988,N_11548,N_11736);
nand U11989 (N_11989,N_11567,N_11700);
nand U11990 (N_11990,N_11597,N_11620);
or U11991 (N_11991,N_11586,N_11584);
nand U11992 (N_11992,N_11699,N_11558);
nand U11993 (N_11993,N_11555,N_11621);
nand U11994 (N_11994,N_11688,N_11630);
xor U11995 (N_11995,N_11563,N_11662);
xor U11996 (N_11996,N_11514,N_11740);
nor U11997 (N_11997,N_11610,N_11597);
xnor U11998 (N_11998,N_11563,N_11589);
or U11999 (N_11999,N_11700,N_11737);
and U12000 (N_12000,N_11964,N_11760);
nor U12001 (N_12001,N_11866,N_11784);
or U12002 (N_12002,N_11805,N_11811);
nand U12003 (N_12003,N_11820,N_11899);
xor U12004 (N_12004,N_11864,N_11799);
or U12005 (N_12005,N_11840,N_11813);
nor U12006 (N_12006,N_11795,N_11900);
nor U12007 (N_12007,N_11817,N_11780);
nand U12008 (N_12008,N_11877,N_11983);
xnor U12009 (N_12009,N_11855,N_11940);
nor U12010 (N_12010,N_11844,N_11908);
nor U12011 (N_12011,N_11829,N_11783);
xor U12012 (N_12012,N_11876,N_11965);
and U12013 (N_12013,N_11819,N_11985);
and U12014 (N_12014,N_11788,N_11991);
nand U12015 (N_12015,N_11972,N_11987);
xor U12016 (N_12016,N_11845,N_11935);
nand U12017 (N_12017,N_11766,N_11892);
and U12018 (N_12018,N_11994,N_11849);
nor U12019 (N_12019,N_11753,N_11936);
xor U12020 (N_12020,N_11816,N_11762);
or U12021 (N_12021,N_11993,N_11938);
xor U12022 (N_12022,N_11898,N_11761);
or U12023 (N_12023,N_11778,N_11773);
or U12024 (N_12024,N_11856,N_11997);
xor U12025 (N_12025,N_11958,N_11962);
xor U12026 (N_12026,N_11974,N_11794);
and U12027 (N_12027,N_11868,N_11986);
xnor U12028 (N_12028,N_11843,N_11836);
nand U12029 (N_12029,N_11809,N_11968);
or U12030 (N_12030,N_11905,N_11869);
and U12031 (N_12031,N_11919,N_11850);
nand U12032 (N_12032,N_11888,N_11966);
nand U12033 (N_12033,N_11975,N_11981);
and U12034 (N_12034,N_11859,N_11901);
nor U12035 (N_12035,N_11772,N_11918);
or U12036 (N_12036,N_11890,N_11990);
nor U12037 (N_12037,N_11906,N_11752);
xor U12038 (N_12038,N_11846,N_11977);
nand U12039 (N_12039,N_11954,N_11973);
xnor U12040 (N_12040,N_11942,N_11848);
and U12041 (N_12041,N_11959,N_11910);
nand U12042 (N_12042,N_11924,N_11804);
and U12043 (N_12043,N_11808,N_11912);
or U12044 (N_12044,N_11758,N_11777);
nor U12045 (N_12045,N_11948,N_11909);
xor U12046 (N_12046,N_11812,N_11923);
xnor U12047 (N_12047,N_11814,N_11828);
or U12048 (N_12048,N_11832,N_11872);
or U12049 (N_12049,N_11945,N_11771);
xor U12050 (N_12050,N_11895,N_11992);
nor U12051 (N_12051,N_11956,N_11765);
nor U12052 (N_12052,N_11838,N_11767);
and U12053 (N_12053,N_11893,N_11914);
xnor U12054 (N_12054,N_11837,N_11928);
and U12055 (N_12055,N_11786,N_11917);
nor U12056 (N_12056,N_11759,N_11827);
or U12057 (N_12057,N_11854,N_11878);
or U12058 (N_12058,N_11963,N_11807);
nor U12059 (N_12059,N_11881,N_11800);
nor U12060 (N_12060,N_11770,N_11999);
nand U12061 (N_12061,N_11861,N_11961);
nor U12062 (N_12062,N_11781,N_11949);
or U12063 (N_12063,N_11875,N_11955);
and U12064 (N_12064,N_11915,N_11857);
nor U12065 (N_12065,N_11852,N_11998);
nor U12066 (N_12066,N_11889,N_11835);
and U12067 (N_12067,N_11996,N_11871);
nor U12068 (N_12068,N_11950,N_11957);
or U12069 (N_12069,N_11894,N_11775);
xor U12070 (N_12070,N_11769,N_11885);
or U12071 (N_12071,N_11870,N_11879);
and U12072 (N_12072,N_11984,N_11793);
xor U12073 (N_12073,N_11853,N_11937);
xor U12074 (N_12074,N_11947,N_11930);
and U12075 (N_12075,N_11929,N_11904);
and U12076 (N_12076,N_11863,N_11941);
or U12077 (N_12077,N_11790,N_11865);
and U12078 (N_12078,N_11971,N_11810);
nand U12079 (N_12079,N_11916,N_11982);
xnor U12080 (N_12080,N_11862,N_11939);
and U12081 (N_12081,N_11911,N_11860);
xnor U12082 (N_12082,N_11883,N_11874);
or U12083 (N_12083,N_11851,N_11821);
or U12084 (N_12084,N_11755,N_11933);
nor U12085 (N_12085,N_11751,N_11970);
nor U12086 (N_12086,N_11884,N_11989);
or U12087 (N_12087,N_11822,N_11951);
nor U12088 (N_12088,N_11921,N_11927);
xor U12089 (N_12089,N_11903,N_11802);
and U12090 (N_12090,N_11953,N_11979);
and U12091 (N_12091,N_11797,N_11934);
xor U12092 (N_12092,N_11980,N_11787);
or U12093 (N_12093,N_11831,N_11842);
nor U12094 (N_12094,N_11926,N_11995);
and U12095 (N_12095,N_11858,N_11932);
or U12096 (N_12096,N_11768,N_11833);
xnor U12097 (N_12097,N_11823,N_11750);
xor U12098 (N_12098,N_11976,N_11887);
or U12099 (N_12099,N_11922,N_11969);
or U12100 (N_12100,N_11789,N_11824);
nand U12101 (N_12101,N_11902,N_11764);
and U12102 (N_12102,N_11931,N_11798);
or U12103 (N_12103,N_11782,N_11886);
nand U12104 (N_12104,N_11776,N_11774);
nand U12105 (N_12105,N_11960,N_11880);
and U12106 (N_12106,N_11891,N_11978);
nand U12107 (N_12107,N_11830,N_11847);
nand U12108 (N_12108,N_11803,N_11867);
and U12109 (N_12109,N_11841,N_11897);
xor U12110 (N_12110,N_11825,N_11754);
or U12111 (N_12111,N_11815,N_11925);
nand U12112 (N_12112,N_11967,N_11907);
and U12113 (N_12113,N_11796,N_11920);
xnor U12114 (N_12114,N_11801,N_11952);
xor U12115 (N_12115,N_11896,N_11763);
nand U12116 (N_12116,N_11943,N_11779);
xnor U12117 (N_12117,N_11818,N_11946);
and U12118 (N_12118,N_11834,N_11785);
nand U12119 (N_12119,N_11839,N_11913);
or U12120 (N_12120,N_11988,N_11944);
nand U12121 (N_12121,N_11806,N_11792);
xor U12122 (N_12122,N_11826,N_11882);
nor U12123 (N_12123,N_11791,N_11757);
nand U12124 (N_12124,N_11756,N_11873);
nand U12125 (N_12125,N_11980,N_11872);
nand U12126 (N_12126,N_11771,N_11895);
nand U12127 (N_12127,N_11777,N_11905);
nand U12128 (N_12128,N_11882,N_11808);
nand U12129 (N_12129,N_11966,N_11822);
nand U12130 (N_12130,N_11965,N_11885);
or U12131 (N_12131,N_11951,N_11859);
nor U12132 (N_12132,N_11886,N_11801);
nor U12133 (N_12133,N_11830,N_11870);
xor U12134 (N_12134,N_11867,N_11816);
nor U12135 (N_12135,N_11786,N_11889);
nor U12136 (N_12136,N_11846,N_11911);
or U12137 (N_12137,N_11945,N_11823);
nand U12138 (N_12138,N_11942,N_11916);
or U12139 (N_12139,N_11988,N_11863);
nand U12140 (N_12140,N_11855,N_11906);
or U12141 (N_12141,N_11818,N_11798);
xnor U12142 (N_12142,N_11924,N_11923);
nor U12143 (N_12143,N_11756,N_11792);
or U12144 (N_12144,N_11889,N_11914);
or U12145 (N_12145,N_11983,N_11879);
nor U12146 (N_12146,N_11877,N_11848);
or U12147 (N_12147,N_11986,N_11983);
and U12148 (N_12148,N_11961,N_11986);
or U12149 (N_12149,N_11754,N_11870);
or U12150 (N_12150,N_11908,N_11918);
or U12151 (N_12151,N_11780,N_11956);
or U12152 (N_12152,N_11990,N_11991);
nor U12153 (N_12153,N_11960,N_11884);
or U12154 (N_12154,N_11969,N_11871);
or U12155 (N_12155,N_11810,N_11832);
and U12156 (N_12156,N_11928,N_11859);
nand U12157 (N_12157,N_11752,N_11793);
nor U12158 (N_12158,N_11801,N_11993);
xnor U12159 (N_12159,N_11826,N_11874);
xor U12160 (N_12160,N_11820,N_11849);
nor U12161 (N_12161,N_11760,N_11961);
xor U12162 (N_12162,N_11951,N_11883);
nor U12163 (N_12163,N_11826,N_11787);
and U12164 (N_12164,N_11990,N_11912);
xnor U12165 (N_12165,N_11764,N_11803);
and U12166 (N_12166,N_11815,N_11999);
nand U12167 (N_12167,N_11809,N_11806);
nand U12168 (N_12168,N_11892,N_11773);
nand U12169 (N_12169,N_11751,N_11949);
and U12170 (N_12170,N_11788,N_11780);
and U12171 (N_12171,N_11948,N_11940);
xnor U12172 (N_12172,N_11797,N_11912);
nand U12173 (N_12173,N_11949,N_11759);
nor U12174 (N_12174,N_11788,N_11899);
nand U12175 (N_12175,N_11929,N_11752);
nand U12176 (N_12176,N_11978,N_11911);
and U12177 (N_12177,N_11945,N_11982);
xor U12178 (N_12178,N_11942,N_11762);
nor U12179 (N_12179,N_11772,N_11982);
nor U12180 (N_12180,N_11882,N_11757);
nand U12181 (N_12181,N_11879,N_11981);
xnor U12182 (N_12182,N_11892,N_11761);
or U12183 (N_12183,N_11844,N_11853);
nor U12184 (N_12184,N_11919,N_11963);
nand U12185 (N_12185,N_11868,N_11907);
and U12186 (N_12186,N_11907,N_11844);
nand U12187 (N_12187,N_11851,N_11832);
and U12188 (N_12188,N_11807,N_11992);
nor U12189 (N_12189,N_11837,N_11915);
xnor U12190 (N_12190,N_11889,N_11761);
and U12191 (N_12191,N_11831,N_11913);
xnor U12192 (N_12192,N_11961,N_11801);
xnor U12193 (N_12193,N_11838,N_11868);
or U12194 (N_12194,N_11969,N_11762);
or U12195 (N_12195,N_11903,N_11832);
nor U12196 (N_12196,N_11943,N_11973);
nand U12197 (N_12197,N_11998,N_11850);
and U12198 (N_12198,N_11868,N_11860);
and U12199 (N_12199,N_11833,N_11904);
or U12200 (N_12200,N_11936,N_11918);
or U12201 (N_12201,N_11937,N_11952);
or U12202 (N_12202,N_11959,N_11844);
nand U12203 (N_12203,N_11811,N_11761);
xnor U12204 (N_12204,N_11831,N_11808);
and U12205 (N_12205,N_11878,N_11927);
xnor U12206 (N_12206,N_11973,N_11858);
nand U12207 (N_12207,N_11766,N_11845);
or U12208 (N_12208,N_11977,N_11844);
xor U12209 (N_12209,N_11981,N_11803);
and U12210 (N_12210,N_11892,N_11938);
or U12211 (N_12211,N_11867,N_11826);
xnor U12212 (N_12212,N_11997,N_11984);
nand U12213 (N_12213,N_11882,N_11803);
xnor U12214 (N_12214,N_11976,N_11869);
nand U12215 (N_12215,N_11788,N_11864);
and U12216 (N_12216,N_11913,N_11990);
xor U12217 (N_12217,N_11964,N_11986);
or U12218 (N_12218,N_11796,N_11887);
and U12219 (N_12219,N_11861,N_11958);
nor U12220 (N_12220,N_11772,N_11991);
nand U12221 (N_12221,N_11823,N_11847);
xnor U12222 (N_12222,N_11884,N_11857);
nand U12223 (N_12223,N_11964,N_11994);
xnor U12224 (N_12224,N_11761,N_11978);
nand U12225 (N_12225,N_11895,N_11813);
xor U12226 (N_12226,N_11790,N_11905);
nand U12227 (N_12227,N_11866,N_11792);
nor U12228 (N_12228,N_11832,N_11815);
nor U12229 (N_12229,N_11750,N_11981);
or U12230 (N_12230,N_11750,N_11932);
xor U12231 (N_12231,N_11863,N_11816);
or U12232 (N_12232,N_11777,N_11782);
and U12233 (N_12233,N_11803,N_11997);
or U12234 (N_12234,N_11912,N_11907);
nor U12235 (N_12235,N_11792,N_11978);
xor U12236 (N_12236,N_11847,N_11906);
or U12237 (N_12237,N_11812,N_11819);
or U12238 (N_12238,N_11998,N_11838);
nor U12239 (N_12239,N_11766,N_11800);
and U12240 (N_12240,N_11943,N_11942);
nor U12241 (N_12241,N_11984,N_11921);
nand U12242 (N_12242,N_11830,N_11781);
nand U12243 (N_12243,N_11927,N_11946);
nor U12244 (N_12244,N_11851,N_11868);
xor U12245 (N_12245,N_11936,N_11980);
nand U12246 (N_12246,N_11855,N_11807);
nor U12247 (N_12247,N_11873,N_11968);
and U12248 (N_12248,N_11772,N_11761);
or U12249 (N_12249,N_11956,N_11861);
or U12250 (N_12250,N_12128,N_12002);
and U12251 (N_12251,N_12109,N_12066);
and U12252 (N_12252,N_12052,N_12126);
and U12253 (N_12253,N_12000,N_12203);
xnor U12254 (N_12254,N_12168,N_12057);
xnor U12255 (N_12255,N_12046,N_12217);
and U12256 (N_12256,N_12174,N_12032);
nand U12257 (N_12257,N_12170,N_12195);
or U12258 (N_12258,N_12073,N_12020);
xor U12259 (N_12259,N_12103,N_12224);
xor U12260 (N_12260,N_12024,N_12165);
nor U12261 (N_12261,N_12177,N_12064);
and U12262 (N_12262,N_12065,N_12081);
xnor U12263 (N_12263,N_12121,N_12102);
nor U12264 (N_12264,N_12127,N_12218);
xnor U12265 (N_12265,N_12184,N_12058);
nor U12266 (N_12266,N_12245,N_12225);
xnor U12267 (N_12267,N_12162,N_12036);
or U12268 (N_12268,N_12160,N_12139);
nand U12269 (N_12269,N_12227,N_12012);
xnor U12270 (N_12270,N_12172,N_12242);
and U12271 (N_12271,N_12043,N_12230);
nand U12272 (N_12272,N_12232,N_12241);
or U12273 (N_12273,N_12204,N_12180);
and U12274 (N_12274,N_12053,N_12238);
or U12275 (N_12275,N_12205,N_12220);
and U12276 (N_12276,N_12152,N_12117);
or U12277 (N_12277,N_12106,N_12236);
nor U12278 (N_12278,N_12200,N_12068);
and U12279 (N_12279,N_12097,N_12096);
nor U12280 (N_12280,N_12156,N_12215);
xor U12281 (N_12281,N_12202,N_12069);
nor U12282 (N_12282,N_12147,N_12100);
and U12283 (N_12283,N_12044,N_12019);
nor U12284 (N_12284,N_12209,N_12243);
nor U12285 (N_12285,N_12076,N_12182);
nand U12286 (N_12286,N_12189,N_12023);
and U12287 (N_12287,N_12146,N_12059);
nor U12288 (N_12288,N_12110,N_12016);
and U12289 (N_12289,N_12143,N_12158);
or U12290 (N_12290,N_12025,N_12042);
and U12291 (N_12291,N_12211,N_12003);
xor U12292 (N_12292,N_12239,N_12027);
or U12293 (N_12293,N_12055,N_12134);
xor U12294 (N_12294,N_12092,N_12108);
and U12295 (N_12295,N_12045,N_12163);
nor U12296 (N_12296,N_12122,N_12192);
nor U12297 (N_12297,N_12034,N_12240);
and U12298 (N_12298,N_12178,N_12071);
nand U12299 (N_12299,N_12190,N_12228);
nand U12300 (N_12300,N_12233,N_12087);
nand U12301 (N_12301,N_12001,N_12007);
or U12302 (N_12302,N_12048,N_12226);
nand U12303 (N_12303,N_12051,N_12207);
nand U12304 (N_12304,N_12054,N_12155);
and U12305 (N_12305,N_12145,N_12026);
and U12306 (N_12306,N_12061,N_12235);
xor U12307 (N_12307,N_12093,N_12095);
nand U12308 (N_12308,N_12231,N_12196);
or U12309 (N_12309,N_12077,N_12098);
nand U12310 (N_12310,N_12033,N_12104);
or U12311 (N_12311,N_12244,N_12086);
and U12312 (N_12312,N_12116,N_12056);
and U12313 (N_12313,N_12094,N_12216);
and U12314 (N_12314,N_12010,N_12210);
and U12315 (N_12315,N_12130,N_12229);
nor U12316 (N_12316,N_12072,N_12080);
or U12317 (N_12317,N_12187,N_12037);
nor U12318 (N_12318,N_12213,N_12021);
xor U12319 (N_12319,N_12142,N_12006);
nand U12320 (N_12320,N_12132,N_12079);
nor U12321 (N_12321,N_12137,N_12169);
nor U12322 (N_12322,N_12176,N_12136);
or U12323 (N_12323,N_12017,N_12031);
xor U12324 (N_12324,N_12113,N_12223);
xnor U12325 (N_12325,N_12085,N_12140);
nor U12326 (N_12326,N_12246,N_12171);
and U12327 (N_12327,N_12015,N_12035);
or U12328 (N_12328,N_12039,N_12214);
nand U12329 (N_12329,N_12135,N_12050);
and U12330 (N_12330,N_12199,N_12179);
and U12331 (N_12331,N_12074,N_12167);
nor U12332 (N_12332,N_12193,N_12107);
and U12333 (N_12333,N_12183,N_12125);
xnor U12334 (N_12334,N_12049,N_12201);
or U12335 (N_12335,N_12157,N_12151);
nor U12336 (N_12336,N_12159,N_12191);
nand U12337 (N_12337,N_12060,N_12181);
or U12338 (N_12338,N_12101,N_12018);
nor U12339 (N_12339,N_12197,N_12091);
or U12340 (N_12340,N_12247,N_12028);
nor U12341 (N_12341,N_12112,N_12022);
nand U12342 (N_12342,N_12148,N_12186);
nor U12343 (N_12343,N_12185,N_12198);
xor U12344 (N_12344,N_12208,N_12038);
nand U12345 (N_12345,N_12138,N_12150);
nor U12346 (N_12346,N_12014,N_12206);
nor U12347 (N_12347,N_12029,N_12118);
nor U12348 (N_12348,N_12188,N_12248);
or U12349 (N_12349,N_12131,N_12030);
nand U12350 (N_12350,N_12008,N_12222);
xor U12351 (N_12351,N_12133,N_12089);
nand U12352 (N_12352,N_12175,N_12141);
nand U12353 (N_12353,N_12153,N_12237);
nor U12354 (N_12354,N_12164,N_12090);
xor U12355 (N_12355,N_12154,N_12005);
nand U12356 (N_12356,N_12041,N_12166);
and U12357 (N_12357,N_12249,N_12013);
nor U12358 (N_12358,N_12004,N_12083);
and U12359 (N_12359,N_12120,N_12123);
xnor U12360 (N_12360,N_12070,N_12084);
xnor U12361 (N_12361,N_12119,N_12234);
or U12362 (N_12362,N_12219,N_12062);
and U12363 (N_12363,N_12078,N_12212);
xor U12364 (N_12364,N_12173,N_12009);
nand U12365 (N_12365,N_12111,N_12149);
nand U12366 (N_12366,N_12088,N_12063);
nor U12367 (N_12367,N_12047,N_12124);
xnor U12368 (N_12368,N_12144,N_12099);
or U12369 (N_12369,N_12114,N_12075);
or U12370 (N_12370,N_12221,N_12040);
or U12371 (N_12371,N_12115,N_12105);
nor U12372 (N_12372,N_12194,N_12161);
xor U12373 (N_12373,N_12129,N_12067);
nor U12374 (N_12374,N_12082,N_12011);
and U12375 (N_12375,N_12166,N_12159);
nor U12376 (N_12376,N_12148,N_12244);
or U12377 (N_12377,N_12040,N_12138);
xor U12378 (N_12378,N_12088,N_12079);
and U12379 (N_12379,N_12218,N_12132);
or U12380 (N_12380,N_12000,N_12129);
xnor U12381 (N_12381,N_12086,N_12077);
xor U12382 (N_12382,N_12245,N_12044);
nor U12383 (N_12383,N_12134,N_12057);
and U12384 (N_12384,N_12036,N_12096);
or U12385 (N_12385,N_12113,N_12243);
xnor U12386 (N_12386,N_12065,N_12103);
nand U12387 (N_12387,N_12087,N_12145);
or U12388 (N_12388,N_12121,N_12010);
nor U12389 (N_12389,N_12115,N_12143);
or U12390 (N_12390,N_12033,N_12010);
and U12391 (N_12391,N_12070,N_12164);
nand U12392 (N_12392,N_12158,N_12184);
xor U12393 (N_12393,N_12176,N_12130);
and U12394 (N_12394,N_12164,N_12206);
or U12395 (N_12395,N_12186,N_12125);
and U12396 (N_12396,N_12207,N_12009);
nand U12397 (N_12397,N_12015,N_12041);
nor U12398 (N_12398,N_12106,N_12083);
and U12399 (N_12399,N_12098,N_12032);
nand U12400 (N_12400,N_12027,N_12220);
xnor U12401 (N_12401,N_12133,N_12014);
nor U12402 (N_12402,N_12094,N_12013);
nand U12403 (N_12403,N_12186,N_12036);
xnor U12404 (N_12404,N_12179,N_12226);
xor U12405 (N_12405,N_12026,N_12222);
and U12406 (N_12406,N_12225,N_12173);
nor U12407 (N_12407,N_12164,N_12177);
or U12408 (N_12408,N_12136,N_12054);
or U12409 (N_12409,N_12136,N_12153);
nor U12410 (N_12410,N_12086,N_12092);
nor U12411 (N_12411,N_12116,N_12106);
or U12412 (N_12412,N_12041,N_12151);
or U12413 (N_12413,N_12028,N_12205);
xor U12414 (N_12414,N_12113,N_12234);
xor U12415 (N_12415,N_12188,N_12005);
xnor U12416 (N_12416,N_12130,N_12076);
nor U12417 (N_12417,N_12145,N_12081);
and U12418 (N_12418,N_12083,N_12171);
or U12419 (N_12419,N_12014,N_12043);
xor U12420 (N_12420,N_12082,N_12046);
xor U12421 (N_12421,N_12190,N_12048);
nand U12422 (N_12422,N_12005,N_12234);
nand U12423 (N_12423,N_12143,N_12058);
xor U12424 (N_12424,N_12068,N_12070);
or U12425 (N_12425,N_12057,N_12092);
nor U12426 (N_12426,N_12063,N_12066);
and U12427 (N_12427,N_12192,N_12130);
nor U12428 (N_12428,N_12097,N_12021);
nand U12429 (N_12429,N_12048,N_12150);
xor U12430 (N_12430,N_12068,N_12236);
or U12431 (N_12431,N_12133,N_12119);
nor U12432 (N_12432,N_12034,N_12173);
nor U12433 (N_12433,N_12231,N_12245);
nor U12434 (N_12434,N_12075,N_12152);
xor U12435 (N_12435,N_12135,N_12059);
nor U12436 (N_12436,N_12188,N_12136);
nor U12437 (N_12437,N_12156,N_12243);
nor U12438 (N_12438,N_12095,N_12162);
and U12439 (N_12439,N_12197,N_12193);
xnor U12440 (N_12440,N_12004,N_12154);
and U12441 (N_12441,N_12002,N_12029);
or U12442 (N_12442,N_12124,N_12154);
nor U12443 (N_12443,N_12203,N_12103);
nor U12444 (N_12444,N_12217,N_12220);
nor U12445 (N_12445,N_12055,N_12049);
nand U12446 (N_12446,N_12147,N_12155);
and U12447 (N_12447,N_12019,N_12176);
nor U12448 (N_12448,N_12060,N_12081);
xnor U12449 (N_12449,N_12221,N_12192);
nor U12450 (N_12450,N_12035,N_12198);
and U12451 (N_12451,N_12096,N_12232);
or U12452 (N_12452,N_12103,N_12166);
nor U12453 (N_12453,N_12143,N_12129);
xnor U12454 (N_12454,N_12201,N_12228);
nor U12455 (N_12455,N_12195,N_12030);
nand U12456 (N_12456,N_12007,N_12095);
and U12457 (N_12457,N_12171,N_12206);
nand U12458 (N_12458,N_12121,N_12056);
and U12459 (N_12459,N_12116,N_12203);
nor U12460 (N_12460,N_12096,N_12200);
nor U12461 (N_12461,N_12163,N_12206);
xor U12462 (N_12462,N_12199,N_12153);
xnor U12463 (N_12463,N_12242,N_12115);
xnor U12464 (N_12464,N_12194,N_12062);
nand U12465 (N_12465,N_12232,N_12182);
or U12466 (N_12466,N_12022,N_12198);
xnor U12467 (N_12467,N_12120,N_12078);
xnor U12468 (N_12468,N_12002,N_12165);
and U12469 (N_12469,N_12075,N_12164);
xor U12470 (N_12470,N_12170,N_12234);
or U12471 (N_12471,N_12177,N_12008);
or U12472 (N_12472,N_12091,N_12107);
nand U12473 (N_12473,N_12132,N_12171);
xnor U12474 (N_12474,N_12150,N_12050);
nor U12475 (N_12475,N_12245,N_12014);
xor U12476 (N_12476,N_12090,N_12148);
nor U12477 (N_12477,N_12085,N_12103);
nand U12478 (N_12478,N_12223,N_12241);
or U12479 (N_12479,N_12215,N_12003);
or U12480 (N_12480,N_12036,N_12243);
or U12481 (N_12481,N_12168,N_12160);
nor U12482 (N_12482,N_12161,N_12074);
or U12483 (N_12483,N_12140,N_12173);
xor U12484 (N_12484,N_12181,N_12230);
nand U12485 (N_12485,N_12244,N_12157);
nand U12486 (N_12486,N_12075,N_12176);
and U12487 (N_12487,N_12200,N_12197);
nand U12488 (N_12488,N_12235,N_12134);
or U12489 (N_12489,N_12010,N_12093);
or U12490 (N_12490,N_12197,N_12087);
or U12491 (N_12491,N_12137,N_12006);
nand U12492 (N_12492,N_12166,N_12171);
nand U12493 (N_12493,N_12178,N_12091);
xor U12494 (N_12494,N_12135,N_12123);
nor U12495 (N_12495,N_12078,N_12119);
nor U12496 (N_12496,N_12159,N_12185);
and U12497 (N_12497,N_12010,N_12217);
xor U12498 (N_12498,N_12215,N_12241);
xnor U12499 (N_12499,N_12224,N_12128);
nor U12500 (N_12500,N_12342,N_12286);
or U12501 (N_12501,N_12421,N_12258);
and U12502 (N_12502,N_12344,N_12436);
xor U12503 (N_12503,N_12423,N_12400);
nor U12504 (N_12504,N_12255,N_12386);
and U12505 (N_12505,N_12497,N_12406);
or U12506 (N_12506,N_12431,N_12388);
nand U12507 (N_12507,N_12446,N_12324);
xnor U12508 (N_12508,N_12323,N_12458);
xnor U12509 (N_12509,N_12276,N_12280);
xor U12510 (N_12510,N_12496,N_12483);
nand U12511 (N_12511,N_12385,N_12326);
or U12512 (N_12512,N_12393,N_12405);
xor U12513 (N_12513,N_12461,N_12440);
and U12514 (N_12514,N_12335,N_12430);
xnor U12515 (N_12515,N_12456,N_12384);
nor U12516 (N_12516,N_12447,N_12357);
or U12517 (N_12517,N_12443,N_12266);
xnor U12518 (N_12518,N_12398,N_12460);
nor U12519 (N_12519,N_12304,N_12473);
nor U12520 (N_12520,N_12284,N_12265);
or U12521 (N_12521,N_12377,N_12451);
and U12522 (N_12522,N_12292,N_12309);
and U12523 (N_12523,N_12469,N_12271);
and U12524 (N_12524,N_12261,N_12389);
xor U12525 (N_12525,N_12364,N_12395);
or U12526 (N_12526,N_12471,N_12404);
nand U12527 (N_12527,N_12345,N_12362);
and U12528 (N_12528,N_12359,N_12348);
and U12529 (N_12529,N_12274,N_12422);
nand U12530 (N_12530,N_12257,N_12272);
and U12531 (N_12531,N_12489,N_12254);
nor U12532 (N_12532,N_12347,N_12498);
or U12533 (N_12533,N_12313,N_12339);
nand U12534 (N_12534,N_12307,N_12275);
nand U12535 (N_12535,N_12330,N_12399);
xnor U12536 (N_12536,N_12334,N_12415);
and U12537 (N_12537,N_12267,N_12486);
xnor U12538 (N_12538,N_12301,N_12351);
nor U12539 (N_12539,N_12371,N_12290);
nand U12540 (N_12540,N_12441,N_12478);
nand U12541 (N_12541,N_12303,N_12297);
nor U12542 (N_12542,N_12358,N_12369);
or U12543 (N_12543,N_12472,N_12302);
or U12544 (N_12544,N_12321,N_12310);
nand U12545 (N_12545,N_12419,N_12437);
xnor U12546 (N_12546,N_12352,N_12413);
and U12547 (N_12547,N_12374,N_12448);
xor U12548 (N_12548,N_12317,N_12314);
nand U12549 (N_12549,N_12312,N_12477);
nand U12550 (N_12550,N_12452,N_12349);
nor U12551 (N_12551,N_12495,N_12277);
or U12552 (N_12552,N_12328,N_12288);
and U12553 (N_12553,N_12337,N_12403);
and U12554 (N_12554,N_12269,N_12382);
nand U12555 (N_12555,N_12391,N_12465);
xor U12556 (N_12556,N_12341,N_12432);
nor U12557 (N_12557,N_12412,N_12468);
or U12558 (N_12558,N_12285,N_12372);
or U12559 (N_12559,N_12250,N_12340);
nor U12560 (N_12560,N_12463,N_12390);
or U12561 (N_12561,N_12363,N_12361);
or U12562 (N_12562,N_12418,N_12373);
or U12563 (N_12563,N_12260,N_12289);
xnor U12564 (N_12564,N_12376,N_12444);
xor U12565 (N_12565,N_12273,N_12279);
nor U12566 (N_12566,N_12488,N_12474);
nor U12567 (N_12567,N_12350,N_12333);
xnor U12568 (N_12568,N_12467,N_12427);
xnor U12569 (N_12569,N_12428,N_12375);
xnor U12570 (N_12570,N_12380,N_12439);
xnor U12571 (N_12571,N_12353,N_12480);
and U12572 (N_12572,N_12453,N_12424);
nand U12573 (N_12573,N_12251,N_12490);
nand U12574 (N_12574,N_12356,N_12379);
nand U12575 (N_12575,N_12354,N_12378);
or U12576 (N_12576,N_12466,N_12476);
xor U12577 (N_12577,N_12367,N_12336);
or U12578 (N_12578,N_12252,N_12387);
nand U12579 (N_12579,N_12318,N_12368);
nor U12580 (N_12580,N_12397,N_12487);
or U12581 (N_12581,N_12283,N_12355);
and U12582 (N_12582,N_12396,N_12365);
xnor U12583 (N_12583,N_12455,N_12256);
or U12584 (N_12584,N_12479,N_12270);
or U12585 (N_12585,N_12401,N_12499);
and U12586 (N_12586,N_12492,N_12278);
nor U12587 (N_12587,N_12433,N_12485);
nor U12588 (N_12588,N_12484,N_12268);
xnor U12589 (N_12589,N_12416,N_12296);
or U12590 (N_12590,N_12253,N_12294);
xnor U12591 (N_12591,N_12315,N_12408);
nand U12592 (N_12592,N_12470,N_12482);
or U12593 (N_12593,N_12299,N_12402);
nand U12594 (N_12594,N_12327,N_12481);
xor U12595 (N_12595,N_12491,N_12305);
xnor U12596 (N_12596,N_12407,N_12287);
or U12597 (N_12597,N_12425,N_12329);
nor U12598 (N_12598,N_12346,N_12311);
xor U12599 (N_12599,N_12464,N_12282);
xnor U12600 (N_12600,N_12410,N_12259);
xnor U12601 (N_12601,N_12392,N_12445);
or U12602 (N_12602,N_12264,N_12438);
nand U12603 (N_12603,N_12475,N_12414);
or U12604 (N_12604,N_12370,N_12429);
xnor U12605 (N_12605,N_12316,N_12435);
nand U12606 (N_12606,N_12426,N_12291);
xor U12607 (N_12607,N_12322,N_12308);
xnor U12608 (N_12608,N_12381,N_12262);
or U12609 (N_12609,N_12434,N_12411);
xor U12610 (N_12610,N_12331,N_12332);
nor U12611 (N_12611,N_12366,N_12281);
or U12612 (N_12612,N_12306,N_12442);
xor U12613 (N_12613,N_12449,N_12494);
or U12614 (N_12614,N_12462,N_12457);
xnor U12615 (N_12615,N_12298,N_12409);
nand U12616 (N_12616,N_12320,N_12417);
and U12617 (N_12617,N_12459,N_12360);
nor U12618 (N_12618,N_12454,N_12295);
and U12619 (N_12619,N_12394,N_12383);
nor U12620 (N_12620,N_12325,N_12293);
nand U12621 (N_12621,N_12300,N_12343);
or U12622 (N_12622,N_12450,N_12493);
or U12623 (N_12623,N_12319,N_12420);
nor U12624 (N_12624,N_12263,N_12338);
xor U12625 (N_12625,N_12278,N_12450);
nand U12626 (N_12626,N_12396,N_12448);
or U12627 (N_12627,N_12263,N_12406);
nand U12628 (N_12628,N_12444,N_12400);
and U12629 (N_12629,N_12296,N_12457);
or U12630 (N_12630,N_12296,N_12311);
nand U12631 (N_12631,N_12393,N_12277);
nor U12632 (N_12632,N_12453,N_12486);
nor U12633 (N_12633,N_12456,N_12472);
nor U12634 (N_12634,N_12400,N_12307);
nand U12635 (N_12635,N_12364,N_12381);
or U12636 (N_12636,N_12461,N_12474);
xnor U12637 (N_12637,N_12257,N_12367);
and U12638 (N_12638,N_12331,N_12366);
nand U12639 (N_12639,N_12395,N_12366);
nand U12640 (N_12640,N_12498,N_12368);
and U12641 (N_12641,N_12431,N_12460);
xnor U12642 (N_12642,N_12433,N_12442);
xor U12643 (N_12643,N_12297,N_12320);
nor U12644 (N_12644,N_12498,N_12471);
nor U12645 (N_12645,N_12479,N_12391);
nand U12646 (N_12646,N_12440,N_12294);
nand U12647 (N_12647,N_12327,N_12331);
nand U12648 (N_12648,N_12434,N_12327);
nand U12649 (N_12649,N_12353,N_12338);
nand U12650 (N_12650,N_12466,N_12373);
nor U12651 (N_12651,N_12365,N_12398);
xnor U12652 (N_12652,N_12483,N_12404);
or U12653 (N_12653,N_12423,N_12386);
nand U12654 (N_12654,N_12373,N_12456);
xnor U12655 (N_12655,N_12471,N_12446);
nand U12656 (N_12656,N_12409,N_12301);
and U12657 (N_12657,N_12493,N_12318);
xor U12658 (N_12658,N_12318,N_12396);
nor U12659 (N_12659,N_12441,N_12469);
xnor U12660 (N_12660,N_12342,N_12469);
xor U12661 (N_12661,N_12473,N_12441);
nor U12662 (N_12662,N_12297,N_12428);
xor U12663 (N_12663,N_12269,N_12432);
nor U12664 (N_12664,N_12279,N_12448);
nand U12665 (N_12665,N_12336,N_12463);
nor U12666 (N_12666,N_12404,N_12252);
nand U12667 (N_12667,N_12395,N_12396);
xor U12668 (N_12668,N_12250,N_12409);
and U12669 (N_12669,N_12405,N_12388);
and U12670 (N_12670,N_12434,N_12308);
xnor U12671 (N_12671,N_12445,N_12337);
or U12672 (N_12672,N_12255,N_12442);
xor U12673 (N_12673,N_12403,N_12420);
nor U12674 (N_12674,N_12454,N_12307);
nand U12675 (N_12675,N_12487,N_12442);
and U12676 (N_12676,N_12465,N_12314);
or U12677 (N_12677,N_12362,N_12412);
nand U12678 (N_12678,N_12486,N_12292);
nand U12679 (N_12679,N_12347,N_12373);
xnor U12680 (N_12680,N_12397,N_12392);
nand U12681 (N_12681,N_12484,N_12460);
or U12682 (N_12682,N_12385,N_12393);
nor U12683 (N_12683,N_12312,N_12483);
xnor U12684 (N_12684,N_12499,N_12430);
or U12685 (N_12685,N_12350,N_12482);
xnor U12686 (N_12686,N_12410,N_12348);
nand U12687 (N_12687,N_12254,N_12318);
or U12688 (N_12688,N_12289,N_12384);
xnor U12689 (N_12689,N_12445,N_12301);
nor U12690 (N_12690,N_12392,N_12464);
nor U12691 (N_12691,N_12456,N_12391);
nand U12692 (N_12692,N_12352,N_12271);
xor U12693 (N_12693,N_12364,N_12445);
and U12694 (N_12694,N_12437,N_12465);
and U12695 (N_12695,N_12407,N_12401);
nor U12696 (N_12696,N_12252,N_12472);
nand U12697 (N_12697,N_12407,N_12316);
nor U12698 (N_12698,N_12399,N_12315);
xor U12699 (N_12699,N_12482,N_12326);
nand U12700 (N_12700,N_12334,N_12393);
nor U12701 (N_12701,N_12259,N_12430);
nor U12702 (N_12702,N_12311,N_12382);
and U12703 (N_12703,N_12338,N_12261);
xnor U12704 (N_12704,N_12440,N_12316);
or U12705 (N_12705,N_12426,N_12448);
or U12706 (N_12706,N_12491,N_12385);
and U12707 (N_12707,N_12300,N_12256);
or U12708 (N_12708,N_12450,N_12265);
xnor U12709 (N_12709,N_12467,N_12294);
nor U12710 (N_12710,N_12316,N_12289);
and U12711 (N_12711,N_12477,N_12280);
xnor U12712 (N_12712,N_12281,N_12440);
xor U12713 (N_12713,N_12474,N_12425);
nor U12714 (N_12714,N_12476,N_12497);
and U12715 (N_12715,N_12402,N_12488);
xnor U12716 (N_12716,N_12311,N_12270);
or U12717 (N_12717,N_12433,N_12367);
nor U12718 (N_12718,N_12355,N_12378);
and U12719 (N_12719,N_12336,N_12473);
nand U12720 (N_12720,N_12368,N_12327);
xnor U12721 (N_12721,N_12390,N_12414);
nor U12722 (N_12722,N_12301,N_12276);
nand U12723 (N_12723,N_12493,N_12292);
and U12724 (N_12724,N_12498,N_12279);
or U12725 (N_12725,N_12497,N_12496);
xnor U12726 (N_12726,N_12364,N_12377);
nor U12727 (N_12727,N_12494,N_12409);
nor U12728 (N_12728,N_12308,N_12407);
or U12729 (N_12729,N_12303,N_12253);
or U12730 (N_12730,N_12492,N_12399);
or U12731 (N_12731,N_12418,N_12316);
nor U12732 (N_12732,N_12458,N_12356);
xor U12733 (N_12733,N_12423,N_12390);
and U12734 (N_12734,N_12446,N_12477);
xnor U12735 (N_12735,N_12398,N_12395);
nor U12736 (N_12736,N_12294,N_12349);
nand U12737 (N_12737,N_12388,N_12463);
or U12738 (N_12738,N_12305,N_12288);
and U12739 (N_12739,N_12450,N_12262);
and U12740 (N_12740,N_12301,N_12284);
and U12741 (N_12741,N_12446,N_12280);
nor U12742 (N_12742,N_12363,N_12395);
and U12743 (N_12743,N_12305,N_12308);
nand U12744 (N_12744,N_12316,N_12286);
and U12745 (N_12745,N_12252,N_12306);
nor U12746 (N_12746,N_12391,N_12476);
nand U12747 (N_12747,N_12295,N_12466);
or U12748 (N_12748,N_12320,N_12354);
xnor U12749 (N_12749,N_12425,N_12385);
and U12750 (N_12750,N_12685,N_12573);
or U12751 (N_12751,N_12716,N_12734);
xnor U12752 (N_12752,N_12540,N_12706);
or U12753 (N_12753,N_12641,N_12747);
xor U12754 (N_12754,N_12568,N_12661);
nor U12755 (N_12755,N_12567,N_12727);
or U12756 (N_12756,N_12707,N_12749);
and U12757 (N_12757,N_12596,N_12587);
and U12758 (N_12758,N_12735,N_12742);
nor U12759 (N_12759,N_12569,N_12691);
and U12760 (N_12760,N_12631,N_12558);
nor U12761 (N_12761,N_12740,N_12636);
nand U12762 (N_12762,N_12659,N_12705);
nor U12763 (N_12763,N_12578,N_12741);
nor U12764 (N_12764,N_12511,N_12724);
xnor U12765 (N_12765,N_12680,N_12515);
nor U12766 (N_12766,N_12585,N_12621);
nor U12767 (N_12767,N_12512,N_12736);
and U12768 (N_12768,N_12637,N_12652);
and U12769 (N_12769,N_12729,N_12725);
nor U12770 (N_12770,N_12551,N_12719);
xnor U12771 (N_12771,N_12528,N_12732);
and U12772 (N_12772,N_12582,N_12581);
and U12773 (N_12773,N_12586,N_12699);
nor U12774 (N_12774,N_12660,N_12522);
or U12775 (N_12775,N_12575,N_12550);
xnor U12776 (N_12776,N_12632,N_12628);
nand U12777 (N_12777,N_12686,N_12730);
or U12778 (N_12778,N_12650,N_12698);
and U12779 (N_12779,N_12668,N_12542);
or U12780 (N_12780,N_12526,N_12745);
nand U12781 (N_12781,N_12547,N_12503);
nand U12782 (N_12782,N_12545,N_12604);
and U12783 (N_12783,N_12692,N_12700);
or U12784 (N_12784,N_12651,N_12605);
and U12785 (N_12785,N_12669,N_12502);
and U12786 (N_12786,N_12667,N_12748);
nand U12787 (N_12787,N_12524,N_12639);
nand U12788 (N_12788,N_12623,N_12607);
xor U12789 (N_12789,N_12633,N_12688);
or U12790 (N_12790,N_12554,N_12520);
and U12791 (N_12791,N_12629,N_12555);
and U12792 (N_12792,N_12689,N_12563);
nand U12793 (N_12793,N_12562,N_12721);
xnor U12794 (N_12794,N_12588,N_12715);
and U12795 (N_12795,N_12674,N_12525);
or U12796 (N_12796,N_12609,N_12549);
nand U12797 (N_12797,N_12658,N_12703);
or U12798 (N_12798,N_12600,N_12720);
nand U12799 (N_12799,N_12744,N_12509);
or U12800 (N_12800,N_12717,N_12572);
nand U12801 (N_12801,N_12574,N_12655);
nand U12802 (N_12802,N_12625,N_12595);
or U12803 (N_12803,N_12684,N_12532);
nand U12804 (N_12804,N_12694,N_12533);
nor U12805 (N_12805,N_12696,N_12530);
nand U12806 (N_12806,N_12675,N_12709);
xnor U12807 (N_12807,N_12556,N_12708);
and U12808 (N_12808,N_12593,N_12552);
and U12809 (N_12809,N_12682,N_12634);
nor U12810 (N_12810,N_12597,N_12642);
nand U12811 (N_12811,N_12601,N_12571);
and U12812 (N_12812,N_12678,N_12619);
xor U12813 (N_12813,N_12670,N_12687);
xor U12814 (N_12814,N_12535,N_12591);
or U12815 (N_12815,N_12612,N_12598);
nand U12816 (N_12816,N_12713,N_12677);
or U12817 (N_12817,N_12516,N_12695);
xor U12818 (N_12818,N_12614,N_12743);
xnor U12819 (N_12819,N_12589,N_12505);
and U12820 (N_12820,N_12643,N_12671);
nand U12821 (N_12821,N_12590,N_12594);
xnor U12822 (N_12822,N_12676,N_12646);
or U12823 (N_12823,N_12517,N_12656);
and U12824 (N_12824,N_12583,N_12733);
nor U12825 (N_12825,N_12622,N_12662);
nand U12826 (N_12826,N_12647,N_12560);
nand U12827 (N_12827,N_12506,N_12663);
and U12828 (N_12828,N_12504,N_12538);
nand U12829 (N_12829,N_12599,N_12710);
nand U12830 (N_12830,N_12559,N_12579);
nor U12831 (N_12831,N_12544,N_12536);
nor U12832 (N_12832,N_12518,N_12508);
xor U12833 (N_12833,N_12712,N_12626);
or U12834 (N_12834,N_12738,N_12565);
or U12835 (N_12835,N_12697,N_12640);
nand U12836 (N_12836,N_12543,N_12739);
nand U12837 (N_12837,N_12722,N_12714);
nand U12838 (N_12838,N_12531,N_12611);
nor U12839 (N_12839,N_12566,N_12548);
nand U12840 (N_12840,N_12702,N_12534);
nand U12841 (N_12841,N_12657,N_12666);
nand U12842 (N_12842,N_12693,N_12606);
or U12843 (N_12843,N_12602,N_12653);
nor U12844 (N_12844,N_12513,N_12701);
nand U12845 (N_12845,N_12673,N_12603);
nand U12846 (N_12846,N_12672,N_12557);
or U12847 (N_12847,N_12523,N_12737);
nor U12848 (N_12848,N_12564,N_12570);
and U12849 (N_12849,N_12718,N_12507);
nand U12850 (N_12850,N_12500,N_12746);
nor U12851 (N_12851,N_12608,N_12519);
or U12852 (N_12852,N_12615,N_12521);
nor U12853 (N_12853,N_12537,N_12630);
nor U12854 (N_12854,N_12649,N_12627);
nand U12855 (N_12855,N_12610,N_12561);
or U12856 (N_12856,N_12635,N_12577);
nand U12857 (N_12857,N_12711,N_12683);
or U12858 (N_12858,N_12546,N_12728);
nand U12859 (N_12859,N_12541,N_12592);
or U12860 (N_12860,N_12731,N_12529);
or U12861 (N_12861,N_12723,N_12624);
nand U12862 (N_12862,N_12580,N_12501);
nor U12863 (N_12863,N_12664,N_12613);
xnor U12864 (N_12864,N_12553,N_12620);
and U12865 (N_12865,N_12648,N_12704);
nand U12866 (N_12866,N_12576,N_12681);
nand U12867 (N_12867,N_12514,N_12527);
nand U12868 (N_12868,N_12618,N_12539);
and U12869 (N_12869,N_12665,N_12584);
or U12870 (N_12870,N_12616,N_12617);
and U12871 (N_12871,N_12654,N_12638);
and U12872 (N_12872,N_12690,N_12510);
and U12873 (N_12873,N_12679,N_12644);
or U12874 (N_12874,N_12645,N_12726);
xor U12875 (N_12875,N_12563,N_12709);
nor U12876 (N_12876,N_12517,N_12682);
and U12877 (N_12877,N_12542,N_12742);
xor U12878 (N_12878,N_12663,N_12537);
nand U12879 (N_12879,N_12617,N_12598);
xnor U12880 (N_12880,N_12683,N_12639);
nor U12881 (N_12881,N_12556,N_12572);
nor U12882 (N_12882,N_12738,N_12694);
nor U12883 (N_12883,N_12503,N_12664);
or U12884 (N_12884,N_12595,N_12582);
nand U12885 (N_12885,N_12516,N_12558);
nand U12886 (N_12886,N_12535,N_12684);
and U12887 (N_12887,N_12688,N_12603);
and U12888 (N_12888,N_12687,N_12646);
or U12889 (N_12889,N_12711,N_12529);
nand U12890 (N_12890,N_12620,N_12581);
nand U12891 (N_12891,N_12587,N_12577);
nand U12892 (N_12892,N_12536,N_12693);
nor U12893 (N_12893,N_12618,N_12696);
or U12894 (N_12894,N_12648,N_12585);
nor U12895 (N_12895,N_12519,N_12742);
or U12896 (N_12896,N_12717,N_12570);
nor U12897 (N_12897,N_12692,N_12576);
or U12898 (N_12898,N_12542,N_12559);
or U12899 (N_12899,N_12665,N_12581);
nand U12900 (N_12900,N_12546,N_12720);
xor U12901 (N_12901,N_12693,N_12707);
or U12902 (N_12902,N_12571,N_12732);
nor U12903 (N_12903,N_12655,N_12562);
or U12904 (N_12904,N_12578,N_12744);
and U12905 (N_12905,N_12681,N_12717);
nand U12906 (N_12906,N_12526,N_12614);
and U12907 (N_12907,N_12623,N_12721);
or U12908 (N_12908,N_12600,N_12508);
and U12909 (N_12909,N_12571,N_12572);
nor U12910 (N_12910,N_12689,N_12680);
nand U12911 (N_12911,N_12518,N_12640);
nand U12912 (N_12912,N_12728,N_12505);
xnor U12913 (N_12913,N_12535,N_12714);
xor U12914 (N_12914,N_12749,N_12571);
and U12915 (N_12915,N_12519,N_12614);
nand U12916 (N_12916,N_12587,N_12645);
xnor U12917 (N_12917,N_12616,N_12675);
and U12918 (N_12918,N_12682,N_12692);
and U12919 (N_12919,N_12562,N_12733);
or U12920 (N_12920,N_12649,N_12609);
or U12921 (N_12921,N_12524,N_12516);
or U12922 (N_12922,N_12531,N_12633);
xor U12923 (N_12923,N_12532,N_12601);
or U12924 (N_12924,N_12535,N_12741);
xnor U12925 (N_12925,N_12710,N_12729);
xnor U12926 (N_12926,N_12713,N_12721);
and U12927 (N_12927,N_12636,N_12630);
nor U12928 (N_12928,N_12603,N_12660);
nor U12929 (N_12929,N_12610,N_12707);
or U12930 (N_12930,N_12705,N_12625);
and U12931 (N_12931,N_12532,N_12716);
and U12932 (N_12932,N_12663,N_12694);
or U12933 (N_12933,N_12668,N_12581);
xor U12934 (N_12934,N_12736,N_12582);
and U12935 (N_12935,N_12679,N_12704);
nor U12936 (N_12936,N_12548,N_12622);
nor U12937 (N_12937,N_12619,N_12695);
nor U12938 (N_12938,N_12694,N_12675);
xnor U12939 (N_12939,N_12741,N_12530);
nand U12940 (N_12940,N_12678,N_12561);
nand U12941 (N_12941,N_12689,N_12567);
nand U12942 (N_12942,N_12622,N_12603);
or U12943 (N_12943,N_12516,N_12707);
or U12944 (N_12944,N_12565,N_12743);
xor U12945 (N_12945,N_12568,N_12564);
nor U12946 (N_12946,N_12699,N_12600);
nand U12947 (N_12947,N_12602,N_12746);
or U12948 (N_12948,N_12616,N_12679);
nor U12949 (N_12949,N_12525,N_12677);
or U12950 (N_12950,N_12554,N_12668);
and U12951 (N_12951,N_12542,N_12566);
or U12952 (N_12952,N_12582,N_12647);
nand U12953 (N_12953,N_12520,N_12637);
or U12954 (N_12954,N_12724,N_12685);
and U12955 (N_12955,N_12588,N_12697);
xnor U12956 (N_12956,N_12605,N_12703);
and U12957 (N_12957,N_12507,N_12695);
xnor U12958 (N_12958,N_12626,N_12639);
xor U12959 (N_12959,N_12748,N_12725);
nand U12960 (N_12960,N_12699,N_12623);
xnor U12961 (N_12961,N_12516,N_12607);
or U12962 (N_12962,N_12606,N_12626);
or U12963 (N_12963,N_12529,N_12627);
and U12964 (N_12964,N_12510,N_12725);
and U12965 (N_12965,N_12576,N_12728);
or U12966 (N_12966,N_12585,N_12642);
xor U12967 (N_12967,N_12720,N_12677);
nand U12968 (N_12968,N_12699,N_12705);
or U12969 (N_12969,N_12562,N_12568);
and U12970 (N_12970,N_12729,N_12558);
nor U12971 (N_12971,N_12535,N_12747);
or U12972 (N_12972,N_12581,N_12670);
or U12973 (N_12973,N_12732,N_12560);
nor U12974 (N_12974,N_12549,N_12641);
nor U12975 (N_12975,N_12654,N_12675);
xor U12976 (N_12976,N_12672,N_12590);
or U12977 (N_12977,N_12572,N_12545);
nand U12978 (N_12978,N_12571,N_12644);
nor U12979 (N_12979,N_12536,N_12509);
and U12980 (N_12980,N_12623,N_12537);
and U12981 (N_12981,N_12749,N_12676);
and U12982 (N_12982,N_12588,N_12501);
and U12983 (N_12983,N_12503,N_12663);
nor U12984 (N_12984,N_12716,N_12675);
or U12985 (N_12985,N_12730,N_12720);
or U12986 (N_12986,N_12647,N_12705);
or U12987 (N_12987,N_12701,N_12563);
and U12988 (N_12988,N_12617,N_12558);
nand U12989 (N_12989,N_12686,N_12647);
xor U12990 (N_12990,N_12664,N_12597);
nand U12991 (N_12991,N_12719,N_12673);
or U12992 (N_12992,N_12695,N_12675);
or U12993 (N_12993,N_12629,N_12682);
and U12994 (N_12994,N_12694,N_12529);
nor U12995 (N_12995,N_12601,N_12580);
nor U12996 (N_12996,N_12503,N_12728);
and U12997 (N_12997,N_12692,N_12555);
xnor U12998 (N_12998,N_12714,N_12740);
nand U12999 (N_12999,N_12632,N_12520);
nor U13000 (N_13000,N_12774,N_12823);
nand U13001 (N_13001,N_12845,N_12846);
nand U13002 (N_13002,N_12946,N_12772);
nand U13003 (N_13003,N_12789,N_12922);
or U13004 (N_13004,N_12999,N_12764);
nor U13005 (N_13005,N_12954,N_12861);
or U13006 (N_13006,N_12941,N_12935);
nor U13007 (N_13007,N_12785,N_12803);
nor U13008 (N_13008,N_12997,N_12948);
xnor U13009 (N_13009,N_12925,N_12841);
and U13010 (N_13010,N_12876,N_12753);
nor U13011 (N_13011,N_12996,N_12831);
and U13012 (N_13012,N_12920,N_12796);
and U13013 (N_13013,N_12908,N_12942);
nor U13014 (N_13014,N_12938,N_12856);
nor U13015 (N_13015,N_12965,N_12927);
and U13016 (N_13016,N_12873,N_12889);
or U13017 (N_13017,N_12888,N_12833);
or U13018 (N_13018,N_12982,N_12821);
nor U13019 (N_13019,N_12991,N_12896);
or U13020 (N_13020,N_12912,N_12877);
and U13021 (N_13021,N_12787,N_12816);
or U13022 (N_13022,N_12924,N_12783);
and U13023 (N_13023,N_12763,N_12869);
nor U13024 (N_13024,N_12824,N_12849);
nor U13025 (N_13025,N_12932,N_12865);
or U13026 (N_13026,N_12778,N_12830);
and U13027 (N_13027,N_12759,N_12780);
or U13028 (N_13028,N_12978,N_12804);
and U13029 (N_13029,N_12878,N_12874);
nor U13030 (N_13030,N_12945,N_12981);
xor U13031 (N_13031,N_12819,N_12977);
or U13032 (N_13032,N_12769,N_12779);
xor U13033 (N_13033,N_12984,N_12893);
nand U13034 (N_13034,N_12926,N_12989);
nand U13035 (N_13035,N_12798,N_12884);
nor U13036 (N_13036,N_12975,N_12799);
or U13037 (N_13037,N_12868,N_12959);
xnor U13038 (N_13038,N_12901,N_12903);
xor U13039 (N_13039,N_12966,N_12914);
or U13040 (N_13040,N_12825,N_12788);
or U13041 (N_13041,N_12900,N_12971);
and U13042 (N_13042,N_12757,N_12930);
nand U13043 (N_13043,N_12771,N_12910);
xnor U13044 (N_13044,N_12974,N_12921);
or U13045 (N_13045,N_12963,N_12775);
nor U13046 (N_13046,N_12832,N_12871);
and U13047 (N_13047,N_12915,N_12943);
and U13048 (N_13048,N_12793,N_12863);
and U13049 (N_13049,N_12766,N_12969);
nor U13050 (N_13050,N_12762,N_12907);
and U13051 (N_13051,N_12847,N_12962);
nor U13052 (N_13052,N_12794,N_12990);
nor U13053 (N_13053,N_12891,N_12752);
xnor U13054 (N_13054,N_12813,N_12802);
or U13055 (N_13055,N_12906,N_12844);
nand U13056 (N_13056,N_12870,N_12812);
nand U13057 (N_13057,N_12980,N_12987);
nand U13058 (N_13058,N_12947,N_12857);
and U13059 (N_13059,N_12756,N_12795);
nor U13060 (N_13060,N_12809,N_12854);
nand U13061 (N_13061,N_12904,N_12820);
or U13062 (N_13062,N_12867,N_12911);
or U13063 (N_13063,N_12973,N_12970);
xnor U13064 (N_13064,N_12807,N_12968);
and U13065 (N_13065,N_12808,N_12894);
and U13066 (N_13066,N_12883,N_12827);
nor U13067 (N_13067,N_12767,N_12750);
and U13068 (N_13068,N_12957,N_12781);
or U13069 (N_13069,N_12862,N_12885);
nand U13070 (N_13070,N_12995,N_12951);
and U13071 (N_13071,N_12864,N_12958);
xor U13072 (N_13072,N_12770,N_12953);
nor U13073 (N_13073,N_12934,N_12838);
and U13074 (N_13074,N_12853,N_12994);
nand U13075 (N_13075,N_12950,N_12758);
nand U13076 (N_13076,N_12851,N_12837);
nor U13077 (N_13077,N_12944,N_12782);
xnor U13078 (N_13078,N_12986,N_12992);
nor U13079 (N_13079,N_12751,N_12937);
and U13080 (N_13080,N_12826,N_12879);
nor U13081 (N_13081,N_12834,N_12828);
and U13082 (N_13082,N_12866,N_12899);
nand U13083 (N_13083,N_12939,N_12858);
xnor U13084 (N_13084,N_12761,N_12792);
and U13085 (N_13085,N_12817,N_12790);
nor U13086 (N_13086,N_12805,N_12786);
nor U13087 (N_13087,N_12880,N_12859);
nor U13088 (N_13088,N_12765,N_12822);
nor U13089 (N_13089,N_12760,N_12902);
nor U13090 (N_13090,N_12988,N_12860);
nor U13091 (N_13091,N_12754,N_12895);
and U13092 (N_13092,N_12852,N_12843);
xor U13093 (N_13093,N_12940,N_12773);
or U13094 (N_13094,N_12886,N_12836);
xnor U13095 (N_13095,N_12918,N_12848);
and U13096 (N_13096,N_12777,N_12875);
or U13097 (N_13097,N_12979,N_12964);
xnor U13098 (N_13098,N_12897,N_12829);
xnor U13099 (N_13099,N_12976,N_12815);
xnor U13100 (N_13100,N_12872,N_12797);
or U13101 (N_13101,N_12919,N_12993);
nor U13102 (N_13102,N_12917,N_12967);
nor U13103 (N_13103,N_12983,N_12791);
nor U13104 (N_13104,N_12985,N_12913);
nor U13105 (N_13105,N_12936,N_12928);
nor U13106 (N_13106,N_12929,N_12855);
nand U13107 (N_13107,N_12961,N_12890);
and U13108 (N_13108,N_12818,N_12835);
and U13109 (N_13109,N_12810,N_12839);
or U13110 (N_13110,N_12882,N_12801);
xnor U13111 (N_13111,N_12881,N_12850);
xor U13112 (N_13112,N_12905,N_12800);
or U13113 (N_13113,N_12776,N_12811);
or U13114 (N_13114,N_12949,N_12923);
or U13115 (N_13115,N_12842,N_12887);
nor U13116 (N_13116,N_12933,N_12806);
or U13117 (N_13117,N_12784,N_12814);
nor U13118 (N_13118,N_12952,N_12892);
nand U13119 (N_13119,N_12998,N_12956);
nor U13120 (N_13120,N_12916,N_12960);
or U13121 (N_13121,N_12955,N_12972);
xnor U13122 (N_13122,N_12909,N_12768);
or U13123 (N_13123,N_12755,N_12898);
xor U13124 (N_13124,N_12931,N_12840);
xor U13125 (N_13125,N_12966,N_12761);
xor U13126 (N_13126,N_12823,N_12994);
nand U13127 (N_13127,N_12817,N_12918);
nor U13128 (N_13128,N_12956,N_12794);
xnor U13129 (N_13129,N_12983,N_12802);
and U13130 (N_13130,N_12789,N_12822);
or U13131 (N_13131,N_12834,N_12969);
or U13132 (N_13132,N_12966,N_12970);
nor U13133 (N_13133,N_12789,N_12896);
and U13134 (N_13134,N_12987,N_12944);
or U13135 (N_13135,N_12764,N_12926);
xor U13136 (N_13136,N_12937,N_12834);
or U13137 (N_13137,N_12991,N_12888);
or U13138 (N_13138,N_12952,N_12857);
and U13139 (N_13139,N_12773,N_12786);
and U13140 (N_13140,N_12926,N_12849);
nor U13141 (N_13141,N_12948,N_12970);
nor U13142 (N_13142,N_12772,N_12851);
nand U13143 (N_13143,N_12773,N_12937);
nor U13144 (N_13144,N_12867,N_12899);
nand U13145 (N_13145,N_12890,N_12963);
nor U13146 (N_13146,N_12841,N_12975);
xnor U13147 (N_13147,N_12836,N_12927);
xnor U13148 (N_13148,N_12930,N_12825);
and U13149 (N_13149,N_12840,N_12751);
nand U13150 (N_13150,N_12768,N_12794);
xnor U13151 (N_13151,N_12865,N_12770);
and U13152 (N_13152,N_12779,N_12997);
nor U13153 (N_13153,N_12752,N_12818);
and U13154 (N_13154,N_12750,N_12995);
xor U13155 (N_13155,N_12893,N_12858);
nand U13156 (N_13156,N_12935,N_12831);
nand U13157 (N_13157,N_12872,N_12760);
xnor U13158 (N_13158,N_12921,N_12836);
and U13159 (N_13159,N_12893,N_12787);
nor U13160 (N_13160,N_12913,N_12912);
xor U13161 (N_13161,N_12825,N_12877);
nor U13162 (N_13162,N_12901,N_12822);
nand U13163 (N_13163,N_12751,N_12825);
nor U13164 (N_13164,N_12812,N_12817);
nand U13165 (N_13165,N_12955,N_12998);
nor U13166 (N_13166,N_12772,N_12967);
xnor U13167 (N_13167,N_12967,N_12946);
and U13168 (N_13168,N_12874,N_12796);
and U13169 (N_13169,N_12866,N_12884);
nor U13170 (N_13170,N_12894,N_12913);
nor U13171 (N_13171,N_12842,N_12991);
nor U13172 (N_13172,N_12801,N_12773);
or U13173 (N_13173,N_12767,N_12809);
and U13174 (N_13174,N_12883,N_12971);
or U13175 (N_13175,N_12837,N_12936);
or U13176 (N_13176,N_12811,N_12792);
nand U13177 (N_13177,N_12990,N_12893);
or U13178 (N_13178,N_12980,N_12856);
or U13179 (N_13179,N_12980,N_12966);
xor U13180 (N_13180,N_12966,N_12855);
and U13181 (N_13181,N_12841,N_12900);
nand U13182 (N_13182,N_12946,N_12755);
or U13183 (N_13183,N_12926,N_12899);
nand U13184 (N_13184,N_12756,N_12831);
xor U13185 (N_13185,N_12755,N_12947);
or U13186 (N_13186,N_12871,N_12913);
or U13187 (N_13187,N_12880,N_12877);
and U13188 (N_13188,N_12801,N_12972);
nor U13189 (N_13189,N_12891,N_12825);
and U13190 (N_13190,N_12890,N_12921);
and U13191 (N_13191,N_12968,N_12951);
xnor U13192 (N_13192,N_12851,N_12836);
or U13193 (N_13193,N_12903,N_12959);
nor U13194 (N_13194,N_12839,N_12780);
or U13195 (N_13195,N_12841,N_12867);
nor U13196 (N_13196,N_12845,N_12873);
nor U13197 (N_13197,N_12860,N_12961);
and U13198 (N_13198,N_12903,N_12893);
nor U13199 (N_13199,N_12996,N_12859);
nand U13200 (N_13200,N_12937,N_12939);
or U13201 (N_13201,N_12953,N_12834);
nand U13202 (N_13202,N_12927,N_12772);
and U13203 (N_13203,N_12864,N_12899);
nand U13204 (N_13204,N_12944,N_12868);
and U13205 (N_13205,N_12770,N_12990);
nor U13206 (N_13206,N_12979,N_12928);
xnor U13207 (N_13207,N_12920,N_12919);
nand U13208 (N_13208,N_12892,N_12942);
nand U13209 (N_13209,N_12890,N_12974);
nor U13210 (N_13210,N_12895,N_12923);
and U13211 (N_13211,N_12993,N_12851);
or U13212 (N_13212,N_12986,N_12950);
or U13213 (N_13213,N_12756,N_12763);
nand U13214 (N_13214,N_12930,N_12956);
and U13215 (N_13215,N_12754,N_12982);
nor U13216 (N_13216,N_12984,N_12993);
nor U13217 (N_13217,N_12919,N_12860);
xnor U13218 (N_13218,N_12794,N_12878);
nand U13219 (N_13219,N_12949,N_12927);
xnor U13220 (N_13220,N_12943,N_12840);
and U13221 (N_13221,N_12881,N_12782);
or U13222 (N_13222,N_12842,N_12852);
xor U13223 (N_13223,N_12852,N_12992);
xnor U13224 (N_13224,N_12847,N_12882);
or U13225 (N_13225,N_12938,N_12949);
nand U13226 (N_13226,N_12861,N_12766);
nor U13227 (N_13227,N_12995,N_12943);
nor U13228 (N_13228,N_12909,N_12791);
nor U13229 (N_13229,N_12758,N_12978);
nand U13230 (N_13230,N_12919,N_12858);
and U13231 (N_13231,N_12787,N_12891);
and U13232 (N_13232,N_12771,N_12757);
xor U13233 (N_13233,N_12919,N_12837);
nor U13234 (N_13234,N_12803,N_12832);
nand U13235 (N_13235,N_12927,N_12943);
nor U13236 (N_13236,N_12846,N_12917);
nor U13237 (N_13237,N_12964,N_12798);
and U13238 (N_13238,N_12881,N_12929);
nor U13239 (N_13239,N_12856,N_12994);
or U13240 (N_13240,N_12997,N_12892);
nand U13241 (N_13241,N_12901,N_12963);
xnor U13242 (N_13242,N_12768,N_12828);
nor U13243 (N_13243,N_12788,N_12969);
and U13244 (N_13244,N_12873,N_12954);
nor U13245 (N_13245,N_12862,N_12760);
nand U13246 (N_13246,N_12754,N_12752);
xor U13247 (N_13247,N_12804,N_12945);
nand U13248 (N_13248,N_12950,N_12771);
nor U13249 (N_13249,N_12774,N_12933);
nand U13250 (N_13250,N_13135,N_13175);
xnor U13251 (N_13251,N_13109,N_13116);
or U13252 (N_13252,N_13023,N_13231);
xor U13253 (N_13253,N_13245,N_13075);
nor U13254 (N_13254,N_13129,N_13153);
nor U13255 (N_13255,N_13131,N_13022);
or U13256 (N_13256,N_13025,N_13078);
or U13257 (N_13257,N_13030,N_13236);
xnor U13258 (N_13258,N_13125,N_13076);
nor U13259 (N_13259,N_13120,N_13107);
and U13260 (N_13260,N_13056,N_13148);
nand U13261 (N_13261,N_13203,N_13186);
xnor U13262 (N_13262,N_13096,N_13095);
nor U13263 (N_13263,N_13014,N_13185);
nand U13264 (N_13264,N_13062,N_13234);
and U13265 (N_13265,N_13141,N_13071);
xnor U13266 (N_13266,N_13220,N_13092);
nor U13267 (N_13267,N_13146,N_13003);
xor U13268 (N_13268,N_13222,N_13080);
nand U13269 (N_13269,N_13027,N_13201);
nand U13270 (N_13270,N_13207,N_13167);
nor U13271 (N_13271,N_13211,N_13124);
nand U13272 (N_13272,N_13055,N_13205);
xor U13273 (N_13273,N_13101,N_13232);
nor U13274 (N_13274,N_13145,N_13065);
nor U13275 (N_13275,N_13108,N_13090);
xor U13276 (N_13276,N_13039,N_13020);
nand U13277 (N_13277,N_13190,N_13048);
and U13278 (N_13278,N_13173,N_13158);
and U13279 (N_13279,N_13210,N_13011);
xor U13280 (N_13280,N_13053,N_13100);
nor U13281 (N_13281,N_13017,N_13215);
xor U13282 (N_13282,N_13157,N_13021);
nor U13283 (N_13283,N_13209,N_13128);
or U13284 (N_13284,N_13156,N_13196);
or U13285 (N_13285,N_13226,N_13034);
nand U13286 (N_13286,N_13008,N_13244);
or U13287 (N_13287,N_13192,N_13106);
nand U13288 (N_13288,N_13189,N_13174);
nand U13289 (N_13289,N_13044,N_13067);
xor U13290 (N_13290,N_13200,N_13235);
nor U13291 (N_13291,N_13068,N_13041);
or U13292 (N_13292,N_13038,N_13180);
nand U13293 (N_13293,N_13103,N_13084);
xnor U13294 (N_13294,N_13249,N_13091);
nor U13295 (N_13295,N_13197,N_13006);
and U13296 (N_13296,N_13227,N_13152);
or U13297 (N_13297,N_13111,N_13233);
and U13298 (N_13298,N_13051,N_13015);
nand U13299 (N_13299,N_13079,N_13182);
nand U13300 (N_13300,N_13213,N_13198);
nand U13301 (N_13301,N_13136,N_13043);
nand U13302 (N_13302,N_13168,N_13126);
xor U13303 (N_13303,N_13072,N_13086);
xnor U13304 (N_13304,N_13113,N_13242);
and U13305 (N_13305,N_13112,N_13105);
nor U13306 (N_13306,N_13133,N_13149);
or U13307 (N_13307,N_13144,N_13214);
or U13308 (N_13308,N_13165,N_13001);
nand U13309 (N_13309,N_13024,N_13195);
or U13310 (N_13310,N_13117,N_13224);
and U13311 (N_13311,N_13052,N_13206);
nor U13312 (N_13312,N_13121,N_13247);
nor U13313 (N_13313,N_13238,N_13179);
nand U13314 (N_13314,N_13114,N_13187);
or U13315 (N_13315,N_13164,N_13202);
or U13316 (N_13316,N_13002,N_13037);
xor U13317 (N_13317,N_13005,N_13177);
nand U13318 (N_13318,N_13139,N_13069);
and U13319 (N_13319,N_13013,N_13031);
nand U13320 (N_13320,N_13059,N_13089);
nand U13321 (N_13321,N_13243,N_13240);
nand U13322 (N_13322,N_13223,N_13188);
nor U13323 (N_13323,N_13077,N_13176);
xnor U13324 (N_13324,N_13221,N_13082);
or U13325 (N_13325,N_13110,N_13150);
nor U13326 (N_13326,N_13087,N_13217);
and U13327 (N_13327,N_13000,N_13183);
xor U13328 (N_13328,N_13035,N_13193);
or U13329 (N_13329,N_13248,N_13191);
and U13330 (N_13330,N_13032,N_13098);
nand U13331 (N_13331,N_13219,N_13147);
xor U13332 (N_13332,N_13061,N_13119);
and U13333 (N_13333,N_13163,N_13130);
and U13334 (N_13334,N_13064,N_13058);
and U13335 (N_13335,N_13134,N_13042);
and U13336 (N_13336,N_13073,N_13143);
nand U13337 (N_13337,N_13070,N_13012);
nor U13338 (N_13338,N_13208,N_13166);
nor U13339 (N_13339,N_13159,N_13097);
or U13340 (N_13340,N_13004,N_13122);
nand U13341 (N_13341,N_13026,N_13118);
xnor U13342 (N_13342,N_13046,N_13140);
or U13343 (N_13343,N_13194,N_13178);
nor U13344 (N_13344,N_13230,N_13169);
xor U13345 (N_13345,N_13029,N_13010);
nand U13346 (N_13346,N_13016,N_13019);
and U13347 (N_13347,N_13216,N_13172);
and U13348 (N_13348,N_13239,N_13184);
and U13349 (N_13349,N_13047,N_13241);
nor U13350 (N_13350,N_13094,N_13054);
xor U13351 (N_13351,N_13151,N_13154);
and U13352 (N_13352,N_13028,N_13063);
and U13353 (N_13353,N_13142,N_13161);
nand U13354 (N_13354,N_13137,N_13160);
and U13355 (N_13355,N_13040,N_13225);
nand U13356 (N_13356,N_13066,N_13049);
and U13357 (N_13357,N_13199,N_13033);
xor U13358 (N_13358,N_13212,N_13057);
nand U13359 (N_13359,N_13060,N_13132);
xnor U13360 (N_13360,N_13018,N_13155);
and U13361 (N_13361,N_13009,N_13204);
xor U13362 (N_13362,N_13036,N_13074);
xor U13363 (N_13363,N_13088,N_13218);
xor U13364 (N_13364,N_13050,N_13083);
or U13365 (N_13365,N_13099,N_13102);
xnor U13366 (N_13366,N_13123,N_13115);
and U13367 (N_13367,N_13170,N_13229);
xnor U13368 (N_13368,N_13228,N_13138);
nor U13369 (N_13369,N_13171,N_13162);
and U13370 (N_13370,N_13045,N_13081);
nand U13371 (N_13371,N_13237,N_13246);
or U13372 (N_13372,N_13007,N_13127);
nand U13373 (N_13373,N_13085,N_13104);
xnor U13374 (N_13374,N_13181,N_13093);
and U13375 (N_13375,N_13117,N_13193);
or U13376 (N_13376,N_13119,N_13080);
nor U13377 (N_13377,N_13120,N_13117);
xor U13378 (N_13378,N_13041,N_13248);
nand U13379 (N_13379,N_13104,N_13122);
xor U13380 (N_13380,N_13148,N_13088);
or U13381 (N_13381,N_13225,N_13070);
or U13382 (N_13382,N_13208,N_13074);
nor U13383 (N_13383,N_13234,N_13203);
nand U13384 (N_13384,N_13120,N_13238);
xnor U13385 (N_13385,N_13144,N_13207);
and U13386 (N_13386,N_13110,N_13059);
and U13387 (N_13387,N_13058,N_13202);
nand U13388 (N_13388,N_13036,N_13054);
nor U13389 (N_13389,N_13189,N_13127);
xnor U13390 (N_13390,N_13151,N_13073);
xor U13391 (N_13391,N_13181,N_13061);
nand U13392 (N_13392,N_13095,N_13083);
nand U13393 (N_13393,N_13019,N_13052);
and U13394 (N_13394,N_13134,N_13076);
xor U13395 (N_13395,N_13169,N_13105);
nand U13396 (N_13396,N_13019,N_13155);
or U13397 (N_13397,N_13087,N_13054);
xor U13398 (N_13398,N_13151,N_13157);
nand U13399 (N_13399,N_13203,N_13148);
and U13400 (N_13400,N_13225,N_13160);
and U13401 (N_13401,N_13243,N_13091);
nand U13402 (N_13402,N_13085,N_13163);
xor U13403 (N_13403,N_13003,N_13038);
nand U13404 (N_13404,N_13137,N_13195);
nor U13405 (N_13405,N_13019,N_13159);
nand U13406 (N_13406,N_13036,N_13151);
or U13407 (N_13407,N_13038,N_13223);
xnor U13408 (N_13408,N_13057,N_13071);
nor U13409 (N_13409,N_13025,N_13169);
nor U13410 (N_13410,N_13032,N_13149);
xnor U13411 (N_13411,N_13174,N_13106);
nand U13412 (N_13412,N_13207,N_13046);
xor U13413 (N_13413,N_13041,N_13237);
or U13414 (N_13414,N_13123,N_13106);
xnor U13415 (N_13415,N_13125,N_13011);
nand U13416 (N_13416,N_13239,N_13006);
nor U13417 (N_13417,N_13052,N_13069);
or U13418 (N_13418,N_13227,N_13145);
or U13419 (N_13419,N_13033,N_13146);
nor U13420 (N_13420,N_13023,N_13142);
xor U13421 (N_13421,N_13154,N_13008);
nor U13422 (N_13422,N_13125,N_13073);
and U13423 (N_13423,N_13185,N_13160);
xor U13424 (N_13424,N_13109,N_13216);
or U13425 (N_13425,N_13047,N_13167);
nand U13426 (N_13426,N_13144,N_13244);
xor U13427 (N_13427,N_13042,N_13036);
or U13428 (N_13428,N_13182,N_13017);
xor U13429 (N_13429,N_13106,N_13067);
or U13430 (N_13430,N_13003,N_13197);
xor U13431 (N_13431,N_13143,N_13103);
and U13432 (N_13432,N_13135,N_13219);
nand U13433 (N_13433,N_13174,N_13066);
nor U13434 (N_13434,N_13123,N_13029);
or U13435 (N_13435,N_13166,N_13028);
and U13436 (N_13436,N_13100,N_13086);
or U13437 (N_13437,N_13010,N_13239);
xor U13438 (N_13438,N_13245,N_13242);
nand U13439 (N_13439,N_13195,N_13071);
xor U13440 (N_13440,N_13159,N_13055);
nand U13441 (N_13441,N_13094,N_13114);
nor U13442 (N_13442,N_13085,N_13212);
nand U13443 (N_13443,N_13116,N_13135);
xnor U13444 (N_13444,N_13071,N_13136);
xnor U13445 (N_13445,N_13110,N_13210);
xnor U13446 (N_13446,N_13046,N_13172);
xor U13447 (N_13447,N_13093,N_13038);
or U13448 (N_13448,N_13007,N_13170);
or U13449 (N_13449,N_13154,N_13199);
and U13450 (N_13450,N_13073,N_13225);
and U13451 (N_13451,N_13109,N_13162);
and U13452 (N_13452,N_13197,N_13172);
xor U13453 (N_13453,N_13041,N_13147);
nand U13454 (N_13454,N_13144,N_13100);
nand U13455 (N_13455,N_13119,N_13179);
xor U13456 (N_13456,N_13207,N_13051);
nand U13457 (N_13457,N_13210,N_13012);
nor U13458 (N_13458,N_13243,N_13136);
xor U13459 (N_13459,N_13140,N_13031);
or U13460 (N_13460,N_13231,N_13217);
and U13461 (N_13461,N_13031,N_13167);
nor U13462 (N_13462,N_13215,N_13053);
and U13463 (N_13463,N_13211,N_13207);
nand U13464 (N_13464,N_13002,N_13232);
or U13465 (N_13465,N_13229,N_13009);
nand U13466 (N_13466,N_13101,N_13237);
xnor U13467 (N_13467,N_13176,N_13076);
and U13468 (N_13468,N_13188,N_13144);
and U13469 (N_13469,N_13045,N_13132);
nor U13470 (N_13470,N_13119,N_13185);
and U13471 (N_13471,N_13136,N_13127);
xnor U13472 (N_13472,N_13204,N_13071);
nor U13473 (N_13473,N_13063,N_13108);
nand U13474 (N_13474,N_13196,N_13232);
or U13475 (N_13475,N_13197,N_13027);
or U13476 (N_13476,N_13154,N_13112);
and U13477 (N_13477,N_13097,N_13236);
or U13478 (N_13478,N_13245,N_13090);
or U13479 (N_13479,N_13032,N_13078);
or U13480 (N_13480,N_13178,N_13043);
or U13481 (N_13481,N_13170,N_13096);
and U13482 (N_13482,N_13009,N_13169);
and U13483 (N_13483,N_13242,N_13032);
xnor U13484 (N_13484,N_13007,N_13033);
or U13485 (N_13485,N_13085,N_13146);
and U13486 (N_13486,N_13016,N_13092);
nand U13487 (N_13487,N_13029,N_13036);
nor U13488 (N_13488,N_13068,N_13174);
xor U13489 (N_13489,N_13155,N_13233);
xor U13490 (N_13490,N_13133,N_13016);
nand U13491 (N_13491,N_13111,N_13226);
xor U13492 (N_13492,N_13081,N_13220);
xor U13493 (N_13493,N_13171,N_13247);
or U13494 (N_13494,N_13042,N_13214);
and U13495 (N_13495,N_13010,N_13191);
nand U13496 (N_13496,N_13071,N_13109);
nor U13497 (N_13497,N_13126,N_13045);
xor U13498 (N_13498,N_13051,N_13122);
nand U13499 (N_13499,N_13035,N_13223);
or U13500 (N_13500,N_13370,N_13467);
xor U13501 (N_13501,N_13390,N_13379);
and U13502 (N_13502,N_13431,N_13327);
nand U13503 (N_13503,N_13301,N_13291);
nor U13504 (N_13504,N_13374,N_13385);
nand U13505 (N_13505,N_13356,N_13286);
or U13506 (N_13506,N_13324,N_13300);
and U13507 (N_13507,N_13391,N_13416);
nor U13508 (N_13508,N_13285,N_13277);
nand U13509 (N_13509,N_13456,N_13446);
and U13510 (N_13510,N_13478,N_13273);
and U13511 (N_13511,N_13399,N_13290);
nand U13512 (N_13512,N_13339,N_13357);
xnor U13513 (N_13513,N_13373,N_13426);
xor U13514 (N_13514,N_13263,N_13303);
and U13515 (N_13515,N_13365,N_13352);
and U13516 (N_13516,N_13322,N_13316);
and U13517 (N_13517,N_13423,N_13477);
xnor U13518 (N_13518,N_13372,N_13296);
or U13519 (N_13519,N_13360,N_13441);
nor U13520 (N_13520,N_13461,N_13338);
or U13521 (N_13521,N_13480,N_13418);
or U13522 (N_13522,N_13438,N_13491);
nor U13523 (N_13523,N_13450,N_13464);
or U13524 (N_13524,N_13264,N_13350);
and U13525 (N_13525,N_13326,N_13499);
nor U13526 (N_13526,N_13334,N_13255);
and U13527 (N_13527,N_13451,N_13346);
xor U13528 (N_13528,N_13295,N_13443);
and U13529 (N_13529,N_13279,N_13458);
nor U13530 (N_13530,N_13332,N_13254);
or U13531 (N_13531,N_13258,N_13293);
and U13532 (N_13532,N_13323,N_13311);
nand U13533 (N_13533,N_13319,N_13473);
xor U13534 (N_13534,N_13363,N_13309);
nand U13535 (N_13535,N_13427,N_13275);
or U13536 (N_13536,N_13392,N_13433);
or U13537 (N_13537,N_13381,N_13417);
xor U13538 (N_13538,N_13410,N_13487);
or U13539 (N_13539,N_13449,N_13278);
nor U13540 (N_13540,N_13272,N_13409);
and U13541 (N_13541,N_13483,N_13497);
or U13542 (N_13542,N_13469,N_13287);
nor U13543 (N_13543,N_13261,N_13305);
or U13544 (N_13544,N_13369,N_13412);
xnor U13545 (N_13545,N_13345,N_13453);
nand U13546 (N_13546,N_13414,N_13289);
nor U13547 (N_13547,N_13398,N_13269);
xor U13548 (N_13548,N_13342,N_13362);
nor U13549 (N_13549,N_13407,N_13270);
and U13550 (N_13550,N_13479,N_13328);
or U13551 (N_13551,N_13354,N_13468);
nand U13552 (N_13552,N_13424,N_13492);
and U13553 (N_13553,N_13382,N_13406);
nor U13554 (N_13554,N_13383,N_13494);
nand U13555 (N_13555,N_13429,N_13436);
or U13556 (N_13556,N_13358,N_13318);
and U13557 (N_13557,N_13386,N_13434);
nand U13558 (N_13558,N_13475,N_13283);
nor U13559 (N_13559,N_13395,N_13257);
nand U13560 (N_13560,N_13280,N_13337);
nand U13561 (N_13561,N_13353,N_13420);
nor U13562 (N_13562,N_13481,N_13294);
xnor U13563 (N_13563,N_13276,N_13355);
or U13564 (N_13564,N_13260,N_13447);
nor U13565 (N_13565,N_13298,N_13321);
nor U13566 (N_13566,N_13393,N_13401);
and U13567 (N_13567,N_13419,N_13344);
or U13568 (N_13568,N_13425,N_13387);
and U13569 (N_13569,N_13366,N_13484);
nor U13570 (N_13570,N_13320,N_13333);
nor U13571 (N_13571,N_13306,N_13282);
and U13572 (N_13572,N_13304,N_13371);
or U13573 (N_13573,N_13396,N_13375);
nand U13574 (N_13574,N_13400,N_13380);
and U13575 (N_13575,N_13347,N_13329);
and U13576 (N_13576,N_13428,N_13348);
or U13577 (N_13577,N_13266,N_13368);
nand U13578 (N_13578,N_13251,N_13466);
nand U13579 (N_13579,N_13343,N_13459);
or U13580 (N_13580,N_13476,N_13376);
and U13581 (N_13581,N_13377,N_13367);
or U13582 (N_13582,N_13361,N_13435);
nor U13583 (N_13583,N_13486,N_13397);
nand U13584 (N_13584,N_13335,N_13474);
xor U13585 (N_13585,N_13307,N_13485);
nor U13586 (N_13586,N_13364,N_13378);
or U13587 (N_13587,N_13310,N_13405);
and U13588 (N_13588,N_13454,N_13463);
xor U13589 (N_13589,N_13432,N_13482);
nand U13590 (N_13590,N_13336,N_13292);
nor U13591 (N_13591,N_13471,N_13402);
xnor U13592 (N_13592,N_13422,N_13267);
or U13593 (N_13593,N_13288,N_13314);
and U13594 (N_13594,N_13325,N_13351);
nand U13595 (N_13595,N_13445,N_13496);
and U13596 (N_13596,N_13302,N_13340);
nand U13597 (N_13597,N_13262,N_13384);
nand U13598 (N_13598,N_13488,N_13317);
or U13599 (N_13599,N_13349,N_13452);
or U13600 (N_13600,N_13448,N_13330);
nand U13601 (N_13601,N_13250,N_13495);
or U13602 (N_13602,N_13498,N_13388);
and U13603 (N_13603,N_13256,N_13470);
nand U13604 (N_13604,N_13489,N_13439);
or U13605 (N_13605,N_13284,N_13415);
and U13606 (N_13606,N_13389,N_13404);
nand U13607 (N_13607,N_13271,N_13465);
xor U13608 (N_13608,N_13253,N_13297);
nor U13609 (N_13609,N_13493,N_13394);
nand U13610 (N_13610,N_13315,N_13460);
nor U13611 (N_13611,N_13413,N_13265);
nand U13612 (N_13612,N_13313,N_13259);
and U13613 (N_13613,N_13472,N_13455);
nand U13614 (N_13614,N_13359,N_13444);
and U13615 (N_13615,N_13440,N_13341);
nand U13616 (N_13616,N_13411,N_13252);
and U13617 (N_13617,N_13430,N_13442);
xor U13618 (N_13618,N_13331,N_13490);
nor U13619 (N_13619,N_13457,N_13308);
xor U13620 (N_13620,N_13274,N_13421);
nand U13621 (N_13621,N_13437,N_13462);
nand U13622 (N_13622,N_13408,N_13299);
or U13623 (N_13623,N_13403,N_13281);
and U13624 (N_13624,N_13268,N_13312);
and U13625 (N_13625,N_13399,N_13394);
nor U13626 (N_13626,N_13492,N_13394);
or U13627 (N_13627,N_13479,N_13426);
nor U13628 (N_13628,N_13330,N_13251);
and U13629 (N_13629,N_13437,N_13324);
xnor U13630 (N_13630,N_13354,N_13486);
nand U13631 (N_13631,N_13334,N_13395);
nand U13632 (N_13632,N_13350,N_13341);
nand U13633 (N_13633,N_13478,N_13348);
xnor U13634 (N_13634,N_13313,N_13318);
nor U13635 (N_13635,N_13369,N_13410);
nand U13636 (N_13636,N_13476,N_13303);
and U13637 (N_13637,N_13425,N_13327);
and U13638 (N_13638,N_13486,N_13403);
or U13639 (N_13639,N_13463,N_13336);
and U13640 (N_13640,N_13421,N_13322);
nand U13641 (N_13641,N_13332,N_13250);
nor U13642 (N_13642,N_13374,N_13384);
xnor U13643 (N_13643,N_13449,N_13257);
and U13644 (N_13644,N_13451,N_13418);
or U13645 (N_13645,N_13349,N_13445);
and U13646 (N_13646,N_13268,N_13427);
and U13647 (N_13647,N_13489,N_13471);
xnor U13648 (N_13648,N_13481,N_13478);
or U13649 (N_13649,N_13390,N_13349);
or U13650 (N_13650,N_13491,N_13412);
nor U13651 (N_13651,N_13289,N_13420);
nand U13652 (N_13652,N_13431,N_13277);
nand U13653 (N_13653,N_13286,N_13440);
nor U13654 (N_13654,N_13354,N_13406);
xnor U13655 (N_13655,N_13394,N_13489);
nor U13656 (N_13656,N_13428,N_13250);
nand U13657 (N_13657,N_13311,N_13482);
nand U13658 (N_13658,N_13383,N_13450);
nor U13659 (N_13659,N_13381,N_13252);
nor U13660 (N_13660,N_13447,N_13412);
and U13661 (N_13661,N_13251,N_13366);
xnor U13662 (N_13662,N_13267,N_13324);
nand U13663 (N_13663,N_13289,N_13421);
or U13664 (N_13664,N_13307,N_13399);
nor U13665 (N_13665,N_13496,N_13337);
nor U13666 (N_13666,N_13494,N_13322);
nor U13667 (N_13667,N_13448,N_13381);
nand U13668 (N_13668,N_13492,N_13455);
nor U13669 (N_13669,N_13269,N_13294);
xnor U13670 (N_13670,N_13393,N_13360);
nor U13671 (N_13671,N_13451,N_13462);
xnor U13672 (N_13672,N_13362,N_13453);
and U13673 (N_13673,N_13266,N_13467);
or U13674 (N_13674,N_13295,N_13486);
xnor U13675 (N_13675,N_13357,N_13427);
and U13676 (N_13676,N_13399,N_13344);
and U13677 (N_13677,N_13265,N_13274);
and U13678 (N_13678,N_13334,N_13328);
or U13679 (N_13679,N_13351,N_13379);
nor U13680 (N_13680,N_13342,N_13448);
and U13681 (N_13681,N_13322,N_13324);
and U13682 (N_13682,N_13325,N_13430);
and U13683 (N_13683,N_13488,N_13333);
or U13684 (N_13684,N_13450,N_13254);
and U13685 (N_13685,N_13293,N_13427);
nor U13686 (N_13686,N_13321,N_13402);
and U13687 (N_13687,N_13355,N_13489);
nand U13688 (N_13688,N_13281,N_13298);
or U13689 (N_13689,N_13260,N_13348);
and U13690 (N_13690,N_13260,N_13254);
xor U13691 (N_13691,N_13398,N_13343);
or U13692 (N_13692,N_13374,N_13341);
xnor U13693 (N_13693,N_13341,N_13491);
or U13694 (N_13694,N_13279,N_13356);
xnor U13695 (N_13695,N_13489,N_13397);
nand U13696 (N_13696,N_13494,N_13289);
or U13697 (N_13697,N_13348,N_13389);
and U13698 (N_13698,N_13285,N_13443);
xnor U13699 (N_13699,N_13445,N_13278);
nand U13700 (N_13700,N_13447,N_13278);
nor U13701 (N_13701,N_13270,N_13382);
xor U13702 (N_13702,N_13416,N_13423);
nor U13703 (N_13703,N_13486,N_13326);
and U13704 (N_13704,N_13318,N_13314);
nand U13705 (N_13705,N_13473,N_13360);
nand U13706 (N_13706,N_13479,N_13312);
nor U13707 (N_13707,N_13443,N_13288);
xor U13708 (N_13708,N_13263,N_13379);
nor U13709 (N_13709,N_13272,N_13496);
nand U13710 (N_13710,N_13358,N_13441);
nand U13711 (N_13711,N_13347,N_13350);
nand U13712 (N_13712,N_13250,N_13331);
nand U13713 (N_13713,N_13447,N_13318);
nand U13714 (N_13714,N_13384,N_13312);
nor U13715 (N_13715,N_13405,N_13465);
xnor U13716 (N_13716,N_13424,N_13475);
xor U13717 (N_13717,N_13340,N_13441);
nor U13718 (N_13718,N_13428,N_13359);
nor U13719 (N_13719,N_13412,N_13406);
xnor U13720 (N_13720,N_13369,N_13494);
nor U13721 (N_13721,N_13450,N_13430);
nand U13722 (N_13722,N_13253,N_13322);
nor U13723 (N_13723,N_13286,N_13353);
and U13724 (N_13724,N_13333,N_13337);
nand U13725 (N_13725,N_13456,N_13315);
and U13726 (N_13726,N_13269,N_13251);
or U13727 (N_13727,N_13311,N_13439);
xnor U13728 (N_13728,N_13467,N_13433);
or U13729 (N_13729,N_13428,N_13270);
and U13730 (N_13730,N_13478,N_13253);
nor U13731 (N_13731,N_13478,N_13460);
nor U13732 (N_13732,N_13338,N_13426);
xnor U13733 (N_13733,N_13463,N_13488);
nand U13734 (N_13734,N_13362,N_13262);
or U13735 (N_13735,N_13345,N_13485);
nand U13736 (N_13736,N_13288,N_13345);
and U13737 (N_13737,N_13469,N_13435);
xnor U13738 (N_13738,N_13495,N_13499);
and U13739 (N_13739,N_13381,N_13298);
nor U13740 (N_13740,N_13406,N_13272);
xor U13741 (N_13741,N_13451,N_13274);
or U13742 (N_13742,N_13473,N_13460);
or U13743 (N_13743,N_13377,N_13397);
nor U13744 (N_13744,N_13434,N_13476);
nand U13745 (N_13745,N_13436,N_13409);
nor U13746 (N_13746,N_13317,N_13348);
xnor U13747 (N_13747,N_13490,N_13475);
nand U13748 (N_13748,N_13290,N_13364);
or U13749 (N_13749,N_13297,N_13258);
or U13750 (N_13750,N_13547,N_13558);
xnor U13751 (N_13751,N_13665,N_13514);
xor U13752 (N_13752,N_13653,N_13604);
and U13753 (N_13753,N_13701,N_13629);
and U13754 (N_13754,N_13656,N_13601);
and U13755 (N_13755,N_13615,N_13559);
xnor U13756 (N_13756,N_13612,N_13677);
or U13757 (N_13757,N_13694,N_13556);
nand U13758 (N_13758,N_13692,N_13678);
or U13759 (N_13759,N_13614,N_13647);
nor U13760 (N_13760,N_13589,N_13606);
nand U13761 (N_13761,N_13509,N_13680);
and U13762 (N_13762,N_13603,N_13578);
xor U13763 (N_13763,N_13628,N_13633);
nor U13764 (N_13764,N_13587,N_13535);
xnor U13765 (N_13765,N_13654,N_13505);
nand U13766 (N_13766,N_13609,N_13700);
nand U13767 (N_13767,N_13643,N_13516);
xor U13768 (N_13768,N_13607,N_13693);
nand U13769 (N_13769,N_13690,N_13721);
and U13770 (N_13770,N_13662,N_13573);
and U13771 (N_13771,N_13675,N_13687);
xnor U13772 (N_13772,N_13741,N_13548);
or U13773 (N_13773,N_13746,N_13507);
nand U13774 (N_13774,N_13672,N_13722);
or U13775 (N_13775,N_13704,N_13709);
nor U13776 (N_13776,N_13626,N_13733);
nand U13777 (N_13777,N_13616,N_13510);
nand U13778 (N_13778,N_13745,N_13584);
or U13779 (N_13779,N_13632,N_13728);
nor U13780 (N_13780,N_13664,N_13568);
nor U13781 (N_13781,N_13511,N_13641);
nand U13782 (N_13782,N_13667,N_13699);
nor U13783 (N_13783,N_13705,N_13506);
nor U13784 (N_13784,N_13540,N_13726);
xor U13785 (N_13785,N_13503,N_13537);
and U13786 (N_13786,N_13658,N_13543);
xor U13787 (N_13787,N_13621,N_13706);
and U13788 (N_13788,N_13521,N_13608);
nor U13789 (N_13789,N_13524,N_13689);
xor U13790 (N_13790,N_13613,N_13671);
and U13791 (N_13791,N_13669,N_13736);
nand U13792 (N_13792,N_13594,N_13528);
xor U13793 (N_13793,N_13517,N_13552);
and U13794 (N_13794,N_13534,N_13597);
xnor U13795 (N_13795,N_13649,N_13622);
or U13796 (N_13796,N_13707,N_13673);
and U13797 (N_13797,N_13637,N_13523);
nor U13798 (N_13798,N_13554,N_13661);
and U13799 (N_13799,N_13681,N_13576);
nor U13800 (N_13800,N_13512,N_13644);
nor U13801 (N_13801,N_13522,N_13611);
xor U13802 (N_13802,N_13651,N_13686);
or U13803 (N_13803,N_13623,N_13570);
and U13804 (N_13804,N_13740,N_13545);
or U13805 (N_13805,N_13749,N_13716);
nor U13806 (N_13806,N_13638,N_13504);
or U13807 (N_13807,N_13725,N_13565);
nor U13808 (N_13808,N_13555,N_13526);
nand U13809 (N_13809,N_13571,N_13569);
nand U13810 (N_13810,N_13581,N_13640);
or U13811 (N_13811,N_13557,N_13739);
xnor U13812 (N_13812,N_13583,N_13718);
nor U13813 (N_13813,N_13525,N_13702);
nand U13814 (N_13814,N_13530,N_13560);
nand U13815 (N_13815,N_13592,N_13684);
nand U13816 (N_13816,N_13634,N_13600);
xor U13817 (N_13817,N_13588,N_13742);
and U13818 (N_13818,N_13659,N_13635);
or U13819 (N_13819,N_13636,N_13602);
nor U13820 (N_13820,N_13546,N_13532);
or U13821 (N_13821,N_13579,N_13657);
xnor U13822 (N_13822,N_13610,N_13691);
or U13823 (N_13823,N_13748,N_13500);
xnor U13824 (N_13824,N_13561,N_13563);
nor U13825 (N_13825,N_13679,N_13685);
and U13826 (N_13826,N_13599,N_13668);
or U13827 (N_13827,N_13648,N_13715);
or U13828 (N_13828,N_13660,N_13703);
nor U13829 (N_13829,N_13712,N_13591);
and U13830 (N_13830,N_13541,N_13708);
and U13831 (N_13831,N_13566,N_13713);
and U13832 (N_13832,N_13627,N_13596);
nand U13833 (N_13833,N_13574,N_13572);
nand U13834 (N_13834,N_13670,N_13618);
xor U13835 (N_13835,N_13595,N_13551);
xnor U13836 (N_13836,N_13585,N_13717);
and U13837 (N_13837,N_13593,N_13743);
and U13838 (N_13838,N_13732,N_13564);
nand U13839 (N_13839,N_13734,N_13682);
and U13840 (N_13840,N_13630,N_13646);
and U13841 (N_13841,N_13586,N_13536);
xor U13842 (N_13842,N_13655,N_13695);
nor U13843 (N_13843,N_13711,N_13650);
or U13844 (N_13844,N_13619,N_13723);
xor U13845 (N_13845,N_13549,N_13518);
xnor U13846 (N_13846,N_13533,N_13519);
nor U13847 (N_13847,N_13501,N_13744);
nor U13848 (N_13848,N_13538,N_13631);
or U13849 (N_13849,N_13575,N_13624);
or U13850 (N_13850,N_13735,N_13508);
xor U13851 (N_13851,N_13710,N_13683);
or U13852 (N_13852,N_13727,N_13730);
nand U13853 (N_13853,N_13663,N_13531);
or U13854 (N_13854,N_13513,N_13747);
nand U13855 (N_13855,N_13729,N_13676);
xnor U13856 (N_13856,N_13639,N_13645);
nand U13857 (N_13857,N_13515,N_13590);
or U13858 (N_13858,N_13605,N_13580);
and U13859 (N_13859,N_13724,N_13620);
and U13860 (N_13860,N_13698,N_13617);
or U13861 (N_13861,N_13688,N_13553);
xor U13862 (N_13862,N_13544,N_13529);
or U13863 (N_13863,N_13567,N_13502);
nand U13864 (N_13864,N_13625,N_13720);
or U13865 (N_13865,N_13527,N_13697);
xor U13866 (N_13866,N_13738,N_13737);
nor U13867 (N_13867,N_13562,N_13542);
nor U13868 (N_13868,N_13582,N_13550);
xnor U13869 (N_13869,N_13714,N_13652);
and U13870 (N_13870,N_13539,N_13731);
or U13871 (N_13871,N_13520,N_13674);
and U13872 (N_13872,N_13642,N_13719);
nand U13873 (N_13873,N_13598,N_13666);
and U13874 (N_13874,N_13577,N_13696);
nand U13875 (N_13875,N_13633,N_13651);
nor U13876 (N_13876,N_13512,N_13636);
nor U13877 (N_13877,N_13613,N_13550);
xor U13878 (N_13878,N_13529,N_13658);
xor U13879 (N_13879,N_13730,N_13512);
nand U13880 (N_13880,N_13728,N_13605);
or U13881 (N_13881,N_13528,N_13648);
and U13882 (N_13882,N_13738,N_13717);
and U13883 (N_13883,N_13618,N_13667);
nand U13884 (N_13884,N_13712,N_13658);
and U13885 (N_13885,N_13686,N_13500);
and U13886 (N_13886,N_13653,N_13623);
xnor U13887 (N_13887,N_13525,N_13633);
nand U13888 (N_13888,N_13627,N_13615);
nor U13889 (N_13889,N_13564,N_13674);
nor U13890 (N_13890,N_13665,N_13683);
nor U13891 (N_13891,N_13646,N_13544);
xnor U13892 (N_13892,N_13598,N_13605);
nor U13893 (N_13893,N_13507,N_13588);
nor U13894 (N_13894,N_13531,N_13611);
or U13895 (N_13895,N_13617,N_13563);
or U13896 (N_13896,N_13646,N_13703);
nor U13897 (N_13897,N_13703,N_13689);
xnor U13898 (N_13898,N_13579,N_13503);
xnor U13899 (N_13899,N_13586,N_13681);
nor U13900 (N_13900,N_13722,N_13513);
or U13901 (N_13901,N_13716,N_13556);
xor U13902 (N_13902,N_13611,N_13744);
xnor U13903 (N_13903,N_13749,N_13556);
nor U13904 (N_13904,N_13652,N_13579);
xnor U13905 (N_13905,N_13606,N_13593);
nor U13906 (N_13906,N_13603,N_13697);
and U13907 (N_13907,N_13667,N_13563);
nor U13908 (N_13908,N_13670,N_13595);
and U13909 (N_13909,N_13549,N_13714);
xor U13910 (N_13910,N_13721,N_13719);
nor U13911 (N_13911,N_13623,N_13631);
and U13912 (N_13912,N_13516,N_13735);
nor U13913 (N_13913,N_13727,N_13553);
nor U13914 (N_13914,N_13523,N_13731);
or U13915 (N_13915,N_13611,N_13677);
and U13916 (N_13916,N_13603,N_13724);
and U13917 (N_13917,N_13700,N_13747);
nor U13918 (N_13918,N_13666,N_13639);
and U13919 (N_13919,N_13652,N_13514);
xor U13920 (N_13920,N_13637,N_13584);
xnor U13921 (N_13921,N_13740,N_13592);
nand U13922 (N_13922,N_13676,N_13675);
nand U13923 (N_13923,N_13748,N_13557);
and U13924 (N_13924,N_13563,N_13682);
nand U13925 (N_13925,N_13550,N_13596);
xor U13926 (N_13926,N_13668,N_13593);
nor U13927 (N_13927,N_13578,N_13566);
nand U13928 (N_13928,N_13604,N_13731);
nand U13929 (N_13929,N_13702,N_13514);
xor U13930 (N_13930,N_13643,N_13659);
nand U13931 (N_13931,N_13664,N_13611);
nor U13932 (N_13932,N_13529,N_13684);
nand U13933 (N_13933,N_13610,N_13617);
and U13934 (N_13934,N_13583,N_13743);
nand U13935 (N_13935,N_13650,N_13733);
and U13936 (N_13936,N_13710,N_13549);
or U13937 (N_13937,N_13737,N_13668);
nand U13938 (N_13938,N_13708,N_13662);
or U13939 (N_13939,N_13733,N_13672);
or U13940 (N_13940,N_13649,N_13653);
nor U13941 (N_13941,N_13715,N_13552);
and U13942 (N_13942,N_13743,N_13671);
and U13943 (N_13943,N_13546,N_13561);
and U13944 (N_13944,N_13648,N_13533);
and U13945 (N_13945,N_13672,N_13669);
nor U13946 (N_13946,N_13503,N_13748);
or U13947 (N_13947,N_13607,N_13649);
nand U13948 (N_13948,N_13670,N_13570);
and U13949 (N_13949,N_13683,N_13652);
and U13950 (N_13950,N_13701,N_13709);
nand U13951 (N_13951,N_13620,N_13686);
and U13952 (N_13952,N_13749,N_13511);
xnor U13953 (N_13953,N_13667,N_13555);
nand U13954 (N_13954,N_13707,N_13553);
nor U13955 (N_13955,N_13557,N_13592);
and U13956 (N_13956,N_13545,N_13695);
and U13957 (N_13957,N_13515,N_13724);
and U13958 (N_13958,N_13649,N_13611);
or U13959 (N_13959,N_13573,N_13623);
and U13960 (N_13960,N_13654,N_13561);
nor U13961 (N_13961,N_13722,N_13675);
and U13962 (N_13962,N_13700,N_13710);
nor U13963 (N_13963,N_13666,N_13596);
nand U13964 (N_13964,N_13516,N_13582);
or U13965 (N_13965,N_13655,N_13661);
and U13966 (N_13966,N_13509,N_13728);
nand U13967 (N_13967,N_13658,N_13577);
nand U13968 (N_13968,N_13741,N_13603);
xnor U13969 (N_13969,N_13638,N_13511);
or U13970 (N_13970,N_13743,N_13737);
nand U13971 (N_13971,N_13707,N_13711);
nor U13972 (N_13972,N_13658,N_13734);
nor U13973 (N_13973,N_13614,N_13584);
nand U13974 (N_13974,N_13664,N_13676);
nor U13975 (N_13975,N_13735,N_13547);
or U13976 (N_13976,N_13546,N_13515);
nand U13977 (N_13977,N_13582,N_13662);
nor U13978 (N_13978,N_13532,N_13735);
nand U13979 (N_13979,N_13701,N_13744);
or U13980 (N_13980,N_13588,N_13719);
nor U13981 (N_13981,N_13516,N_13511);
xor U13982 (N_13982,N_13749,N_13740);
or U13983 (N_13983,N_13545,N_13705);
nor U13984 (N_13984,N_13621,N_13540);
nand U13985 (N_13985,N_13628,N_13723);
or U13986 (N_13986,N_13654,N_13713);
nand U13987 (N_13987,N_13691,N_13529);
nor U13988 (N_13988,N_13550,N_13566);
and U13989 (N_13989,N_13734,N_13659);
and U13990 (N_13990,N_13710,N_13682);
nor U13991 (N_13991,N_13666,N_13632);
nand U13992 (N_13992,N_13612,N_13641);
or U13993 (N_13993,N_13565,N_13701);
xnor U13994 (N_13994,N_13669,N_13650);
xor U13995 (N_13995,N_13678,N_13689);
and U13996 (N_13996,N_13558,N_13613);
and U13997 (N_13997,N_13634,N_13512);
xor U13998 (N_13998,N_13725,N_13569);
or U13999 (N_13999,N_13524,N_13579);
xor U14000 (N_14000,N_13803,N_13919);
and U14001 (N_14001,N_13780,N_13886);
xnor U14002 (N_14002,N_13892,N_13767);
nor U14003 (N_14003,N_13963,N_13914);
xnor U14004 (N_14004,N_13847,N_13883);
nor U14005 (N_14005,N_13943,N_13861);
nand U14006 (N_14006,N_13974,N_13960);
or U14007 (N_14007,N_13990,N_13876);
and U14008 (N_14008,N_13811,N_13750);
or U14009 (N_14009,N_13879,N_13796);
or U14010 (N_14010,N_13875,N_13901);
nand U14011 (N_14011,N_13928,N_13944);
nor U14012 (N_14012,N_13957,N_13762);
nor U14013 (N_14013,N_13830,N_13893);
and U14014 (N_14014,N_13826,N_13786);
or U14015 (N_14015,N_13797,N_13999);
nand U14016 (N_14016,N_13833,N_13848);
xor U14017 (N_14017,N_13906,N_13840);
nand U14018 (N_14018,N_13801,N_13831);
nand U14019 (N_14019,N_13806,N_13955);
nor U14020 (N_14020,N_13761,N_13985);
nand U14021 (N_14021,N_13968,N_13857);
or U14022 (N_14022,N_13766,N_13822);
nand U14023 (N_14023,N_13937,N_13846);
xnor U14024 (N_14024,N_13874,N_13975);
or U14025 (N_14025,N_13828,N_13878);
xnor U14026 (N_14026,N_13757,N_13946);
and U14027 (N_14027,N_13983,N_13866);
nand U14028 (N_14028,N_13841,N_13864);
or U14029 (N_14029,N_13933,N_13823);
nand U14030 (N_14030,N_13877,N_13821);
nand U14031 (N_14031,N_13979,N_13896);
nor U14032 (N_14032,N_13954,N_13941);
and U14033 (N_14033,N_13865,N_13768);
xor U14034 (N_14034,N_13987,N_13973);
or U14035 (N_14035,N_13977,N_13887);
or U14036 (N_14036,N_13770,N_13966);
or U14037 (N_14037,N_13905,N_13882);
xnor U14038 (N_14038,N_13751,N_13777);
and U14039 (N_14039,N_13899,N_13863);
xor U14040 (N_14040,N_13935,N_13781);
or U14041 (N_14041,N_13785,N_13853);
nor U14042 (N_14042,N_13862,N_13858);
nand U14043 (N_14043,N_13981,N_13754);
xnor U14044 (N_14044,N_13769,N_13995);
and U14045 (N_14045,N_13918,N_13965);
nor U14046 (N_14046,N_13889,N_13792);
and U14047 (N_14047,N_13800,N_13917);
xor U14048 (N_14048,N_13779,N_13815);
nand U14049 (N_14049,N_13939,N_13911);
nor U14050 (N_14050,N_13895,N_13772);
nand U14051 (N_14051,N_13756,N_13812);
nor U14052 (N_14052,N_13898,N_13798);
or U14053 (N_14053,N_13788,N_13787);
and U14054 (N_14054,N_13904,N_13989);
xor U14055 (N_14055,N_13993,N_13764);
nand U14056 (N_14056,N_13805,N_13802);
nand U14057 (N_14057,N_13890,N_13845);
nand U14058 (N_14058,N_13967,N_13940);
or U14059 (N_14059,N_13991,N_13956);
nor U14060 (N_14060,N_13818,N_13799);
and U14061 (N_14061,N_13888,N_13851);
xor U14062 (N_14062,N_13884,N_13854);
nand U14063 (N_14063,N_13948,N_13825);
nor U14064 (N_14064,N_13832,N_13843);
nand U14065 (N_14065,N_13871,N_13922);
or U14066 (N_14066,N_13894,N_13872);
xor U14067 (N_14067,N_13813,N_13932);
nand U14068 (N_14068,N_13870,N_13763);
nor U14069 (N_14069,N_13789,N_13807);
nor U14070 (N_14070,N_13902,N_13951);
and U14071 (N_14071,N_13827,N_13984);
or U14072 (N_14072,N_13774,N_13867);
nand U14073 (N_14073,N_13753,N_13916);
nand U14074 (N_14074,N_13820,N_13850);
and U14075 (N_14075,N_13844,N_13793);
or U14076 (N_14076,N_13924,N_13880);
xor U14077 (N_14077,N_13783,N_13929);
nand U14078 (N_14078,N_13997,N_13931);
nand U14079 (N_14079,N_13834,N_13810);
or U14080 (N_14080,N_13936,N_13791);
nand U14081 (N_14081,N_13860,N_13868);
or U14082 (N_14082,N_13925,N_13869);
and U14083 (N_14083,N_13838,N_13961);
xnor U14084 (N_14084,N_13920,N_13942);
and U14085 (N_14085,N_13817,N_13913);
nand U14086 (N_14086,N_13923,N_13809);
nand U14087 (N_14087,N_13775,N_13819);
and U14088 (N_14088,N_13962,N_13824);
nor U14089 (N_14089,N_13814,N_13926);
or U14090 (N_14090,N_13778,N_13760);
nand U14091 (N_14091,N_13910,N_13915);
xor U14092 (N_14092,N_13835,N_13976);
xnor U14093 (N_14093,N_13994,N_13856);
xnor U14094 (N_14094,N_13837,N_13934);
or U14095 (N_14095,N_13849,N_13836);
and U14096 (N_14096,N_13765,N_13852);
and U14097 (N_14097,N_13912,N_13839);
nand U14098 (N_14098,N_13759,N_13959);
or U14099 (N_14099,N_13903,N_13776);
and U14100 (N_14100,N_13804,N_13752);
nand U14101 (N_14101,N_13930,N_13784);
xnor U14102 (N_14102,N_13908,N_13972);
or U14103 (N_14103,N_13859,N_13921);
nand U14104 (N_14104,N_13873,N_13900);
or U14105 (N_14105,N_13945,N_13927);
or U14106 (N_14106,N_13808,N_13982);
nand U14107 (N_14107,N_13988,N_13795);
nand U14108 (N_14108,N_13953,N_13950);
nand U14109 (N_14109,N_13816,N_13790);
and U14110 (N_14110,N_13971,N_13771);
or U14111 (N_14111,N_13938,N_13986);
and U14112 (N_14112,N_13794,N_13996);
xor U14113 (N_14113,N_13881,N_13949);
xnor U14114 (N_14114,N_13969,N_13978);
or U14115 (N_14115,N_13885,N_13964);
xor U14116 (N_14116,N_13842,N_13897);
and U14117 (N_14117,N_13952,N_13907);
nand U14118 (N_14118,N_13773,N_13782);
xor U14119 (N_14119,N_13998,N_13970);
and U14120 (N_14120,N_13891,N_13909);
nor U14121 (N_14121,N_13980,N_13947);
nor U14122 (N_14122,N_13855,N_13829);
or U14123 (N_14123,N_13755,N_13992);
or U14124 (N_14124,N_13758,N_13958);
xnor U14125 (N_14125,N_13810,N_13827);
nand U14126 (N_14126,N_13804,N_13859);
xnor U14127 (N_14127,N_13771,N_13885);
and U14128 (N_14128,N_13800,N_13795);
xnor U14129 (N_14129,N_13894,N_13811);
or U14130 (N_14130,N_13814,N_13896);
nor U14131 (N_14131,N_13880,N_13850);
nand U14132 (N_14132,N_13844,N_13871);
or U14133 (N_14133,N_13808,N_13761);
xnor U14134 (N_14134,N_13932,N_13819);
nand U14135 (N_14135,N_13947,N_13972);
nand U14136 (N_14136,N_13891,N_13916);
xor U14137 (N_14137,N_13810,N_13980);
and U14138 (N_14138,N_13910,N_13837);
nand U14139 (N_14139,N_13956,N_13754);
nand U14140 (N_14140,N_13835,N_13920);
or U14141 (N_14141,N_13928,N_13832);
nor U14142 (N_14142,N_13940,N_13799);
nand U14143 (N_14143,N_13822,N_13754);
or U14144 (N_14144,N_13852,N_13782);
or U14145 (N_14145,N_13861,N_13958);
xor U14146 (N_14146,N_13798,N_13968);
and U14147 (N_14147,N_13956,N_13964);
nand U14148 (N_14148,N_13763,N_13966);
nand U14149 (N_14149,N_13979,N_13772);
nor U14150 (N_14150,N_13836,N_13858);
and U14151 (N_14151,N_13800,N_13756);
or U14152 (N_14152,N_13779,N_13887);
xor U14153 (N_14153,N_13964,N_13783);
nand U14154 (N_14154,N_13937,N_13938);
xnor U14155 (N_14155,N_13805,N_13927);
nand U14156 (N_14156,N_13795,N_13871);
nor U14157 (N_14157,N_13990,N_13968);
nand U14158 (N_14158,N_13856,N_13878);
and U14159 (N_14159,N_13977,N_13907);
and U14160 (N_14160,N_13958,N_13842);
nand U14161 (N_14161,N_13815,N_13842);
nor U14162 (N_14162,N_13910,N_13974);
xnor U14163 (N_14163,N_13827,N_13903);
or U14164 (N_14164,N_13963,N_13954);
nand U14165 (N_14165,N_13983,N_13994);
and U14166 (N_14166,N_13919,N_13985);
or U14167 (N_14167,N_13848,N_13838);
nand U14168 (N_14168,N_13801,N_13946);
nor U14169 (N_14169,N_13900,N_13980);
and U14170 (N_14170,N_13808,N_13900);
nor U14171 (N_14171,N_13901,N_13844);
and U14172 (N_14172,N_13998,N_13982);
xnor U14173 (N_14173,N_13937,N_13956);
or U14174 (N_14174,N_13979,N_13856);
or U14175 (N_14175,N_13851,N_13893);
nor U14176 (N_14176,N_13813,N_13946);
or U14177 (N_14177,N_13955,N_13898);
and U14178 (N_14178,N_13763,N_13845);
nand U14179 (N_14179,N_13997,N_13921);
nand U14180 (N_14180,N_13787,N_13952);
nor U14181 (N_14181,N_13757,N_13926);
and U14182 (N_14182,N_13839,N_13944);
or U14183 (N_14183,N_13925,N_13911);
nand U14184 (N_14184,N_13843,N_13914);
or U14185 (N_14185,N_13880,N_13838);
xor U14186 (N_14186,N_13803,N_13768);
nor U14187 (N_14187,N_13893,N_13888);
and U14188 (N_14188,N_13868,N_13965);
and U14189 (N_14189,N_13779,N_13974);
xor U14190 (N_14190,N_13906,N_13929);
xor U14191 (N_14191,N_13797,N_13750);
xnor U14192 (N_14192,N_13953,N_13940);
nor U14193 (N_14193,N_13975,N_13837);
nor U14194 (N_14194,N_13755,N_13881);
or U14195 (N_14195,N_13953,N_13978);
or U14196 (N_14196,N_13921,N_13891);
or U14197 (N_14197,N_13973,N_13955);
nand U14198 (N_14198,N_13928,N_13927);
and U14199 (N_14199,N_13882,N_13896);
nand U14200 (N_14200,N_13841,N_13768);
nand U14201 (N_14201,N_13865,N_13918);
or U14202 (N_14202,N_13772,N_13752);
nand U14203 (N_14203,N_13945,N_13950);
xor U14204 (N_14204,N_13755,N_13861);
and U14205 (N_14205,N_13924,N_13810);
nor U14206 (N_14206,N_13777,N_13950);
or U14207 (N_14207,N_13889,N_13996);
and U14208 (N_14208,N_13926,N_13942);
nand U14209 (N_14209,N_13772,N_13941);
xor U14210 (N_14210,N_13911,N_13783);
xnor U14211 (N_14211,N_13949,N_13893);
and U14212 (N_14212,N_13852,N_13814);
nand U14213 (N_14213,N_13791,N_13842);
and U14214 (N_14214,N_13988,N_13797);
xnor U14215 (N_14215,N_13918,N_13814);
or U14216 (N_14216,N_13850,N_13815);
or U14217 (N_14217,N_13953,N_13824);
nor U14218 (N_14218,N_13890,N_13999);
nor U14219 (N_14219,N_13836,N_13818);
nand U14220 (N_14220,N_13908,N_13798);
nor U14221 (N_14221,N_13865,N_13871);
nor U14222 (N_14222,N_13856,N_13906);
xnor U14223 (N_14223,N_13999,N_13937);
and U14224 (N_14224,N_13756,N_13856);
or U14225 (N_14225,N_13809,N_13770);
and U14226 (N_14226,N_13874,N_13806);
nor U14227 (N_14227,N_13755,N_13849);
or U14228 (N_14228,N_13752,N_13825);
nor U14229 (N_14229,N_13859,N_13931);
or U14230 (N_14230,N_13984,N_13828);
xnor U14231 (N_14231,N_13804,N_13941);
and U14232 (N_14232,N_13818,N_13890);
xnor U14233 (N_14233,N_13905,N_13791);
nand U14234 (N_14234,N_13846,N_13955);
and U14235 (N_14235,N_13815,N_13760);
and U14236 (N_14236,N_13946,N_13878);
or U14237 (N_14237,N_13848,N_13863);
nor U14238 (N_14238,N_13751,N_13864);
and U14239 (N_14239,N_13794,N_13862);
nand U14240 (N_14240,N_13900,N_13861);
nand U14241 (N_14241,N_13817,N_13886);
or U14242 (N_14242,N_13763,N_13872);
or U14243 (N_14243,N_13980,N_13921);
or U14244 (N_14244,N_13900,N_13765);
xnor U14245 (N_14245,N_13933,N_13976);
xnor U14246 (N_14246,N_13985,N_13791);
nor U14247 (N_14247,N_13830,N_13945);
nor U14248 (N_14248,N_13771,N_13905);
nand U14249 (N_14249,N_13794,N_13942);
or U14250 (N_14250,N_14141,N_14180);
or U14251 (N_14251,N_14234,N_14037);
nand U14252 (N_14252,N_14010,N_14096);
nor U14253 (N_14253,N_14082,N_14212);
xor U14254 (N_14254,N_14056,N_14106);
or U14255 (N_14255,N_14189,N_14199);
or U14256 (N_14256,N_14134,N_14057);
xnor U14257 (N_14257,N_14066,N_14247);
nand U14258 (N_14258,N_14140,N_14148);
nor U14259 (N_14259,N_14014,N_14008);
or U14260 (N_14260,N_14110,N_14088);
and U14261 (N_14261,N_14054,N_14155);
nor U14262 (N_14262,N_14249,N_14003);
xnor U14263 (N_14263,N_14025,N_14102);
or U14264 (N_14264,N_14211,N_14092);
xor U14265 (N_14265,N_14004,N_14103);
nand U14266 (N_14266,N_14118,N_14062);
and U14267 (N_14267,N_14204,N_14233);
or U14268 (N_14268,N_14237,N_14001);
xnor U14269 (N_14269,N_14201,N_14151);
xor U14270 (N_14270,N_14187,N_14031);
nor U14271 (N_14271,N_14162,N_14229);
and U14272 (N_14272,N_14217,N_14084);
and U14273 (N_14273,N_14123,N_14013);
or U14274 (N_14274,N_14173,N_14163);
xor U14275 (N_14275,N_14072,N_14024);
or U14276 (N_14276,N_14090,N_14152);
and U14277 (N_14277,N_14169,N_14100);
nand U14278 (N_14278,N_14073,N_14042);
xnor U14279 (N_14279,N_14193,N_14006);
xor U14280 (N_14280,N_14114,N_14023);
and U14281 (N_14281,N_14130,N_14133);
xor U14282 (N_14282,N_14190,N_14105);
and U14283 (N_14283,N_14016,N_14227);
and U14284 (N_14284,N_14074,N_14104);
xor U14285 (N_14285,N_14149,N_14039);
xnor U14286 (N_14286,N_14135,N_14243);
nand U14287 (N_14287,N_14112,N_14051);
and U14288 (N_14288,N_14172,N_14012);
nor U14289 (N_14289,N_14144,N_14132);
or U14290 (N_14290,N_14245,N_14027);
nand U14291 (N_14291,N_14099,N_14226);
and U14292 (N_14292,N_14126,N_14108);
and U14293 (N_14293,N_14115,N_14041);
and U14294 (N_14294,N_14160,N_14116);
or U14295 (N_14295,N_14098,N_14026);
nand U14296 (N_14296,N_14195,N_14036);
and U14297 (N_14297,N_14040,N_14223);
and U14298 (N_14298,N_14030,N_14079);
xnor U14299 (N_14299,N_14166,N_14034);
nand U14300 (N_14300,N_14033,N_14181);
or U14301 (N_14301,N_14081,N_14136);
or U14302 (N_14302,N_14121,N_14224);
nor U14303 (N_14303,N_14047,N_14119);
xnor U14304 (N_14304,N_14182,N_14202);
nor U14305 (N_14305,N_14046,N_14240);
and U14306 (N_14306,N_14188,N_14053);
xor U14307 (N_14307,N_14021,N_14083);
nor U14308 (N_14308,N_14035,N_14060);
and U14309 (N_14309,N_14007,N_14129);
or U14310 (N_14310,N_14145,N_14045);
or U14311 (N_14311,N_14177,N_14097);
or U14312 (N_14312,N_14048,N_14065);
xnor U14313 (N_14313,N_14131,N_14020);
and U14314 (N_14314,N_14002,N_14186);
and U14315 (N_14315,N_14159,N_14069);
or U14316 (N_14316,N_14101,N_14207);
nor U14317 (N_14317,N_14158,N_14168);
and U14318 (N_14318,N_14218,N_14117);
nor U14319 (N_14319,N_14128,N_14086);
and U14320 (N_14320,N_14009,N_14091);
xor U14321 (N_14321,N_14248,N_14167);
nand U14322 (N_14322,N_14078,N_14064);
nand U14323 (N_14323,N_14153,N_14070);
and U14324 (N_14324,N_14228,N_14044);
nor U14325 (N_14325,N_14179,N_14208);
and U14326 (N_14326,N_14067,N_14242);
xnor U14327 (N_14327,N_14170,N_14244);
nand U14328 (N_14328,N_14137,N_14171);
nand U14329 (N_14329,N_14176,N_14210);
and U14330 (N_14330,N_14184,N_14087);
xor U14331 (N_14331,N_14213,N_14221);
xnor U14332 (N_14332,N_14220,N_14018);
nor U14333 (N_14333,N_14235,N_14209);
nand U14334 (N_14334,N_14185,N_14038);
nand U14335 (N_14335,N_14178,N_14068);
nor U14336 (N_14336,N_14236,N_14146);
nor U14337 (N_14337,N_14198,N_14094);
nand U14338 (N_14338,N_14015,N_14093);
or U14339 (N_14339,N_14022,N_14058);
nor U14340 (N_14340,N_14120,N_14143);
and U14341 (N_14341,N_14241,N_14192);
nor U14342 (N_14342,N_14230,N_14183);
and U14343 (N_14343,N_14032,N_14174);
xor U14344 (N_14344,N_14216,N_14175);
and U14345 (N_14345,N_14138,N_14246);
xnor U14346 (N_14346,N_14222,N_14127);
nor U14347 (N_14347,N_14239,N_14111);
or U14348 (N_14348,N_14109,N_14019);
and U14349 (N_14349,N_14028,N_14075);
nand U14350 (N_14350,N_14011,N_14238);
and U14351 (N_14351,N_14164,N_14206);
and U14352 (N_14352,N_14156,N_14005);
and U14353 (N_14353,N_14071,N_14165);
and U14354 (N_14354,N_14203,N_14017);
or U14355 (N_14355,N_14139,N_14077);
or U14356 (N_14356,N_14050,N_14063);
nor U14357 (N_14357,N_14194,N_14154);
and U14358 (N_14358,N_14076,N_14049);
xor U14359 (N_14359,N_14232,N_14142);
or U14360 (N_14360,N_14000,N_14113);
and U14361 (N_14361,N_14225,N_14061);
and U14362 (N_14362,N_14052,N_14059);
and U14363 (N_14363,N_14200,N_14089);
or U14364 (N_14364,N_14125,N_14043);
or U14365 (N_14365,N_14161,N_14085);
nor U14366 (N_14366,N_14214,N_14095);
nand U14367 (N_14367,N_14196,N_14231);
and U14368 (N_14368,N_14124,N_14122);
and U14369 (N_14369,N_14157,N_14205);
nor U14370 (N_14370,N_14197,N_14219);
nor U14371 (N_14371,N_14147,N_14107);
nor U14372 (N_14372,N_14191,N_14080);
xnor U14373 (N_14373,N_14055,N_14150);
and U14374 (N_14374,N_14215,N_14029);
nand U14375 (N_14375,N_14203,N_14092);
or U14376 (N_14376,N_14208,N_14134);
or U14377 (N_14377,N_14034,N_14106);
xor U14378 (N_14378,N_14241,N_14079);
nand U14379 (N_14379,N_14045,N_14151);
and U14380 (N_14380,N_14176,N_14147);
or U14381 (N_14381,N_14174,N_14056);
and U14382 (N_14382,N_14064,N_14004);
or U14383 (N_14383,N_14024,N_14184);
nor U14384 (N_14384,N_14193,N_14194);
or U14385 (N_14385,N_14142,N_14006);
or U14386 (N_14386,N_14119,N_14127);
nand U14387 (N_14387,N_14227,N_14010);
nor U14388 (N_14388,N_14061,N_14008);
xnor U14389 (N_14389,N_14197,N_14169);
and U14390 (N_14390,N_14246,N_14129);
or U14391 (N_14391,N_14155,N_14038);
and U14392 (N_14392,N_14226,N_14076);
nand U14393 (N_14393,N_14117,N_14017);
or U14394 (N_14394,N_14236,N_14031);
nand U14395 (N_14395,N_14239,N_14006);
nor U14396 (N_14396,N_14223,N_14210);
and U14397 (N_14397,N_14100,N_14216);
nor U14398 (N_14398,N_14041,N_14054);
or U14399 (N_14399,N_14178,N_14193);
nor U14400 (N_14400,N_14174,N_14241);
and U14401 (N_14401,N_14189,N_14125);
and U14402 (N_14402,N_14158,N_14019);
or U14403 (N_14403,N_14003,N_14107);
and U14404 (N_14404,N_14025,N_14203);
nand U14405 (N_14405,N_14088,N_14213);
xnor U14406 (N_14406,N_14127,N_14141);
and U14407 (N_14407,N_14177,N_14176);
or U14408 (N_14408,N_14220,N_14234);
or U14409 (N_14409,N_14091,N_14192);
nor U14410 (N_14410,N_14022,N_14115);
nand U14411 (N_14411,N_14226,N_14149);
xor U14412 (N_14412,N_14225,N_14011);
or U14413 (N_14413,N_14202,N_14115);
or U14414 (N_14414,N_14231,N_14107);
nor U14415 (N_14415,N_14230,N_14231);
nor U14416 (N_14416,N_14071,N_14218);
xor U14417 (N_14417,N_14147,N_14196);
nand U14418 (N_14418,N_14218,N_14225);
nor U14419 (N_14419,N_14088,N_14051);
nor U14420 (N_14420,N_14172,N_14031);
and U14421 (N_14421,N_14155,N_14051);
xnor U14422 (N_14422,N_14243,N_14174);
nor U14423 (N_14423,N_14057,N_14148);
nor U14424 (N_14424,N_14011,N_14219);
nand U14425 (N_14425,N_14115,N_14174);
xnor U14426 (N_14426,N_14045,N_14089);
and U14427 (N_14427,N_14105,N_14044);
nor U14428 (N_14428,N_14176,N_14168);
nand U14429 (N_14429,N_14042,N_14005);
xnor U14430 (N_14430,N_14091,N_14124);
or U14431 (N_14431,N_14001,N_14042);
nor U14432 (N_14432,N_14056,N_14067);
and U14433 (N_14433,N_14224,N_14099);
or U14434 (N_14434,N_14062,N_14087);
nand U14435 (N_14435,N_14021,N_14085);
and U14436 (N_14436,N_14046,N_14142);
xor U14437 (N_14437,N_14237,N_14224);
xor U14438 (N_14438,N_14145,N_14086);
nor U14439 (N_14439,N_14204,N_14201);
xor U14440 (N_14440,N_14039,N_14214);
nor U14441 (N_14441,N_14072,N_14147);
and U14442 (N_14442,N_14125,N_14009);
and U14443 (N_14443,N_14209,N_14236);
xnor U14444 (N_14444,N_14216,N_14065);
xor U14445 (N_14445,N_14053,N_14112);
and U14446 (N_14446,N_14144,N_14099);
nor U14447 (N_14447,N_14234,N_14058);
xor U14448 (N_14448,N_14031,N_14141);
and U14449 (N_14449,N_14001,N_14174);
and U14450 (N_14450,N_14111,N_14123);
and U14451 (N_14451,N_14218,N_14186);
or U14452 (N_14452,N_14026,N_14129);
xor U14453 (N_14453,N_14080,N_14083);
nor U14454 (N_14454,N_14093,N_14043);
xor U14455 (N_14455,N_14198,N_14080);
xnor U14456 (N_14456,N_14206,N_14107);
or U14457 (N_14457,N_14142,N_14180);
xnor U14458 (N_14458,N_14182,N_14015);
and U14459 (N_14459,N_14233,N_14111);
or U14460 (N_14460,N_14135,N_14010);
and U14461 (N_14461,N_14085,N_14235);
or U14462 (N_14462,N_14018,N_14123);
xor U14463 (N_14463,N_14246,N_14196);
nand U14464 (N_14464,N_14059,N_14196);
xnor U14465 (N_14465,N_14021,N_14126);
nand U14466 (N_14466,N_14211,N_14126);
and U14467 (N_14467,N_14157,N_14041);
xnor U14468 (N_14468,N_14222,N_14173);
or U14469 (N_14469,N_14018,N_14163);
xnor U14470 (N_14470,N_14220,N_14052);
xnor U14471 (N_14471,N_14137,N_14121);
xnor U14472 (N_14472,N_14044,N_14021);
or U14473 (N_14473,N_14042,N_14238);
and U14474 (N_14474,N_14226,N_14072);
nor U14475 (N_14475,N_14108,N_14017);
nor U14476 (N_14476,N_14213,N_14045);
or U14477 (N_14477,N_14042,N_14044);
xnor U14478 (N_14478,N_14095,N_14100);
nor U14479 (N_14479,N_14166,N_14225);
xor U14480 (N_14480,N_14159,N_14103);
xnor U14481 (N_14481,N_14248,N_14022);
xnor U14482 (N_14482,N_14131,N_14184);
nand U14483 (N_14483,N_14019,N_14247);
xnor U14484 (N_14484,N_14151,N_14005);
xnor U14485 (N_14485,N_14007,N_14154);
or U14486 (N_14486,N_14130,N_14151);
nand U14487 (N_14487,N_14094,N_14108);
nor U14488 (N_14488,N_14109,N_14081);
nand U14489 (N_14489,N_14085,N_14106);
or U14490 (N_14490,N_14213,N_14046);
or U14491 (N_14491,N_14132,N_14060);
or U14492 (N_14492,N_14221,N_14126);
nand U14493 (N_14493,N_14032,N_14150);
and U14494 (N_14494,N_14210,N_14087);
xnor U14495 (N_14495,N_14196,N_14079);
nand U14496 (N_14496,N_14018,N_14019);
nor U14497 (N_14497,N_14133,N_14110);
xnor U14498 (N_14498,N_14161,N_14187);
or U14499 (N_14499,N_14202,N_14007);
or U14500 (N_14500,N_14407,N_14293);
and U14501 (N_14501,N_14297,N_14290);
xnor U14502 (N_14502,N_14366,N_14393);
nand U14503 (N_14503,N_14443,N_14333);
or U14504 (N_14504,N_14343,N_14310);
xnor U14505 (N_14505,N_14433,N_14405);
xnor U14506 (N_14506,N_14312,N_14431);
and U14507 (N_14507,N_14497,N_14378);
and U14508 (N_14508,N_14449,N_14499);
nor U14509 (N_14509,N_14417,N_14390);
and U14510 (N_14510,N_14464,N_14353);
or U14511 (N_14511,N_14493,N_14352);
nor U14512 (N_14512,N_14380,N_14482);
nand U14513 (N_14513,N_14489,N_14439);
and U14514 (N_14514,N_14256,N_14325);
xor U14515 (N_14515,N_14280,N_14294);
and U14516 (N_14516,N_14438,N_14252);
xor U14517 (N_14517,N_14484,N_14316);
xnor U14518 (N_14518,N_14286,N_14479);
and U14519 (N_14519,N_14428,N_14491);
or U14520 (N_14520,N_14460,N_14445);
or U14521 (N_14521,N_14367,N_14328);
nor U14522 (N_14522,N_14391,N_14269);
nor U14523 (N_14523,N_14329,N_14301);
nor U14524 (N_14524,N_14476,N_14319);
or U14525 (N_14525,N_14307,N_14488);
nand U14526 (N_14526,N_14336,N_14300);
xor U14527 (N_14527,N_14330,N_14478);
xnor U14528 (N_14528,N_14250,N_14372);
xnor U14529 (N_14529,N_14322,N_14348);
nor U14530 (N_14530,N_14485,N_14399);
nor U14531 (N_14531,N_14344,N_14317);
nand U14532 (N_14532,N_14442,N_14462);
and U14533 (N_14533,N_14412,N_14483);
nand U14534 (N_14534,N_14292,N_14456);
nor U14535 (N_14535,N_14427,N_14283);
nor U14536 (N_14536,N_14468,N_14435);
nand U14537 (N_14537,N_14263,N_14459);
xor U14538 (N_14538,N_14327,N_14262);
nor U14539 (N_14539,N_14376,N_14425);
xnor U14540 (N_14540,N_14430,N_14289);
or U14541 (N_14541,N_14345,N_14311);
or U14542 (N_14542,N_14447,N_14466);
and U14543 (N_14543,N_14326,N_14382);
xor U14544 (N_14544,N_14415,N_14429);
or U14545 (N_14545,N_14303,N_14346);
nand U14546 (N_14546,N_14287,N_14259);
nand U14547 (N_14547,N_14419,N_14337);
or U14548 (N_14548,N_14323,N_14272);
and U14549 (N_14549,N_14444,N_14260);
nand U14550 (N_14550,N_14349,N_14281);
or U14551 (N_14551,N_14291,N_14395);
nor U14552 (N_14552,N_14432,N_14461);
nor U14553 (N_14553,N_14304,N_14341);
nand U14554 (N_14554,N_14457,N_14318);
or U14555 (N_14555,N_14254,N_14475);
xor U14556 (N_14556,N_14487,N_14267);
or U14557 (N_14557,N_14371,N_14356);
or U14558 (N_14558,N_14387,N_14373);
xnor U14559 (N_14559,N_14320,N_14480);
nand U14560 (N_14560,N_14278,N_14458);
and U14561 (N_14561,N_14408,N_14298);
nor U14562 (N_14562,N_14473,N_14418);
nor U14563 (N_14563,N_14455,N_14261);
or U14564 (N_14564,N_14406,N_14369);
nand U14565 (N_14565,N_14306,N_14340);
nor U14566 (N_14566,N_14490,N_14446);
xnor U14567 (N_14567,N_14339,N_14463);
and U14568 (N_14568,N_14386,N_14251);
and U14569 (N_14569,N_14315,N_14299);
nor U14570 (N_14570,N_14355,N_14365);
or U14571 (N_14571,N_14381,N_14383);
nor U14572 (N_14572,N_14441,N_14270);
or U14573 (N_14573,N_14389,N_14398);
or U14574 (N_14574,N_14358,N_14454);
or U14575 (N_14575,N_14375,N_14305);
nand U14576 (N_14576,N_14402,N_14354);
and U14577 (N_14577,N_14275,N_14440);
and U14578 (N_14578,N_14410,N_14266);
or U14579 (N_14579,N_14268,N_14332);
and U14580 (N_14580,N_14423,N_14401);
nor U14581 (N_14581,N_14351,N_14424);
xnor U14582 (N_14582,N_14359,N_14481);
and U14583 (N_14583,N_14388,N_14452);
and U14584 (N_14584,N_14295,N_14416);
or U14585 (N_14585,N_14363,N_14364);
and U14586 (N_14586,N_14265,N_14360);
xor U14587 (N_14587,N_14374,N_14400);
nor U14588 (N_14588,N_14421,N_14394);
or U14589 (N_14589,N_14321,N_14377);
nor U14590 (N_14590,N_14296,N_14477);
nand U14591 (N_14591,N_14471,N_14282);
nand U14592 (N_14592,N_14302,N_14436);
nor U14593 (N_14593,N_14350,N_14335);
or U14594 (N_14594,N_14411,N_14469);
nor U14595 (N_14595,N_14308,N_14486);
or U14596 (N_14596,N_14370,N_14409);
nand U14597 (N_14597,N_14494,N_14496);
nand U14598 (N_14598,N_14279,N_14347);
nand U14599 (N_14599,N_14420,N_14277);
xor U14600 (N_14600,N_14334,N_14396);
nand U14601 (N_14601,N_14313,N_14379);
nand U14602 (N_14602,N_14255,N_14368);
nand U14603 (N_14603,N_14338,N_14495);
or U14604 (N_14604,N_14273,N_14288);
and U14605 (N_14605,N_14253,N_14414);
nand U14606 (N_14606,N_14397,N_14448);
xor U14607 (N_14607,N_14492,N_14271);
nor U14608 (N_14608,N_14472,N_14470);
xor U14609 (N_14609,N_14403,N_14274);
or U14610 (N_14610,N_14276,N_14264);
and U14611 (N_14611,N_14392,N_14309);
nor U14612 (N_14612,N_14314,N_14437);
nor U14613 (N_14613,N_14404,N_14467);
or U14614 (N_14614,N_14331,N_14422);
nand U14615 (N_14615,N_14385,N_14384);
and U14616 (N_14616,N_14451,N_14426);
nand U14617 (N_14617,N_14284,N_14434);
or U14618 (N_14618,N_14361,N_14474);
nor U14619 (N_14619,N_14285,N_14450);
nand U14620 (N_14620,N_14465,N_14324);
and U14621 (N_14621,N_14453,N_14257);
nand U14622 (N_14622,N_14498,N_14413);
nand U14623 (N_14623,N_14342,N_14362);
or U14624 (N_14624,N_14357,N_14258);
xor U14625 (N_14625,N_14294,N_14364);
nor U14626 (N_14626,N_14367,N_14342);
nand U14627 (N_14627,N_14314,N_14466);
xnor U14628 (N_14628,N_14461,N_14418);
or U14629 (N_14629,N_14265,N_14296);
nand U14630 (N_14630,N_14444,N_14411);
nand U14631 (N_14631,N_14461,N_14316);
nor U14632 (N_14632,N_14295,N_14435);
nor U14633 (N_14633,N_14301,N_14403);
or U14634 (N_14634,N_14400,N_14356);
xnor U14635 (N_14635,N_14406,N_14414);
or U14636 (N_14636,N_14377,N_14350);
nor U14637 (N_14637,N_14421,N_14455);
or U14638 (N_14638,N_14298,N_14274);
xor U14639 (N_14639,N_14382,N_14273);
nand U14640 (N_14640,N_14273,N_14293);
nor U14641 (N_14641,N_14369,N_14253);
nor U14642 (N_14642,N_14278,N_14345);
and U14643 (N_14643,N_14424,N_14491);
nor U14644 (N_14644,N_14470,N_14440);
and U14645 (N_14645,N_14302,N_14274);
nand U14646 (N_14646,N_14421,N_14372);
nand U14647 (N_14647,N_14271,N_14441);
nor U14648 (N_14648,N_14443,N_14409);
and U14649 (N_14649,N_14482,N_14352);
xor U14650 (N_14650,N_14333,N_14335);
xnor U14651 (N_14651,N_14386,N_14309);
nand U14652 (N_14652,N_14405,N_14313);
nand U14653 (N_14653,N_14344,N_14364);
xnor U14654 (N_14654,N_14469,N_14325);
or U14655 (N_14655,N_14316,N_14270);
nand U14656 (N_14656,N_14365,N_14314);
xor U14657 (N_14657,N_14397,N_14382);
or U14658 (N_14658,N_14349,N_14272);
or U14659 (N_14659,N_14302,N_14399);
nor U14660 (N_14660,N_14465,N_14303);
or U14661 (N_14661,N_14295,N_14262);
nand U14662 (N_14662,N_14279,N_14411);
nor U14663 (N_14663,N_14266,N_14329);
nor U14664 (N_14664,N_14422,N_14377);
xor U14665 (N_14665,N_14310,N_14403);
nand U14666 (N_14666,N_14457,N_14401);
nor U14667 (N_14667,N_14421,N_14325);
nor U14668 (N_14668,N_14459,N_14381);
or U14669 (N_14669,N_14402,N_14376);
nor U14670 (N_14670,N_14376,N_14270);
nand U14671 (N_14671,N_14408,N_14345);
nand U14672 (N_14672,N_14310,N_14493);
or U14673 (N_14673,N_14344,N_14352);
nand U14674 (N_14674,N_14303,N_14268);
xor U14675 (N_14675,N_14473,N_14268);
and U14676 (N_14676,N_14383,N_14446);
or U14677 (N_14677,N_14484,N_14459);
nand U14678 (N_14678,N_14495,N_14478);
and U14679 (N_14679,N_14336,N_14431);
or U14680 (N_14680,N_14304,N_14463);
or U14681 (N_14681,N_14432,N_14330);
nand U14682 (N_14682,N_14286,N_14474);
or U14683 (N_14683,N_14483,N_14487);
or U14684 (N_14684,N_14446,N_14465);
nand U14685 (N_14685,N_14458,N_14305);
nor U14686 (N_14686,N_14439,N_14478);
xnor U14687 (N_14687,N_14288,N_14480);
nand U14688 (N_14688,N_14389,N_14481);
xnor U14689 (N_14689,N_14390,N_14384);
and U14690 (N_14690,N_14270,N_14406);
nor U14691 (N_14691,N_14382,N_14340);
nor U14692 (N_14692,N_14258,N_14431);
or U14693 (N_14693,N_14353,N_14458);
and U14694 (N_14694,N_14443,N_14365);
and U14695 (N_14695,N_14494,N_14325);
xnor U14696 (N_14696,N_14429,N_14327);
xnor U14697 (N_14697,N_14311,N_14269);
xor U14698 (N_14698,N_14389,N_14361);
and U14699 (N_14699,N_14386,N_14440);
and U14700 (N_14700,N_14449,N_14420);
or U14701 (N_14701,N_14456,N_14435);
xor U14702 (N_14702,N_14496,N_14252);
nand U14703 (N_14703,N_14453,N_14436);
nand U14704 (N_14704,N_14427,N_14282);
xor U14705 (N_14705,N_14483,N_14451);
and U14706 (N_14706,N_14453,N_14334);
nor U14707 (N_14707,N_14384,N_14363);
nor U14708 (N_14708,N_14456,N_14325);
nor U14709 (N_14709,N_14338,N_14374);
nor U14710 (N_14710,N_14446,N_14469);
nor U14711 (N_14711,N_14321,N_14491);
and U14712 (N_14712,N_14256,N_14499);
or U14713 (N_14713,N_14425,N_14282);
nor U14714 (N_14714,N_14388,N_14334);
nor U14715 (N_14715,N_14400,N_14263);
nor U14716 (N_14716,N_14307,N_14408);
nand U14717 (N_14717,N_14407,N_14341);
and U14718 (N_14718,N_14417,N_14278);
nor U14719 (N_14719,N_14343,N_14294);
xor U14720 (N_14720,N_14475,N_14322);
nor U14721 (N_14721,N_14403,N_14459);
nand U14722 (N_14722,N_14451,N_14261);
or U14723 (N_14723,N_14292,N_14256);
nand U14724 (N_14724,N_14485,N_14266);
nor U14725 (N_14725,N_14309,N_14462);
nor U14726 (N_14726,N_14372,N_14447);
nand U14727 (N_14727,N_14316,N_14382);
nor U14728 (N_14728,N_14268,N_14438);
nand U14729 (N_14729,N_14409,N_14420);
xor U14730 (N_14730,N_14333,N_14250);
nand U14731 (N_14731,N_14379,N_14272);
nand U14732 (N_14732,N_14352,N_14439);
and U14733 (N_14733,N_14320,N_14255);
xnor U14734 (N_14734,N_14429,N_14411);
and U14735 (N_14735,N_14288,N_14423);
and U14736 (N_14736,N_14449,N_14442);
or U14737 (N_14737,N_14282,N_14360);
xor U14738 (N_14738,N_14385,N_14375);
and U14739 (N_14739,N_14366,N_14253);
nor U14740 (N_14740,N_14378,N_14434);
nor U14741 (N_14741,N_14413,N_14252);
xor U14742 (N_14742,N_14352,N_14447);
nor U14743 (N_14743,N_14281,N_14420);
nor U14744 (N_14744,N_14268,N_14355);
nor U14745 (N_14745,N_14253,N_14349);
nor U14746 (N_14746,N_14397,N_14340);
nand U14747 (N_14747,N_14270,N_14437);
and U14748 (N_14748,N_14348,N_14460);
nand U14749 (N_14749,N_14430,N_14278);
and U14750 (N_14750,N_14638,N_14647);
nand U14751 (N_14751,N_14701,N_14548);
xnor U14752 (N_14752,N_14578,N_14737);
and U14753 (N_14753,N_14740,N_14553);
nand U14754 (N_14754,N_14608,N_14529);
and U14755 (N_14755,N_14663,N_14625);
nand U14756 (N_14756,N_14585,N_14695);
and U14757 (N_14757,N_14590,N_14557);
xnor U14758 (N_14758,N_14530,N_14576);
nand U14759 (N_14759,N_14653,N_14639);
or U14760 (N_14760,N_14565,N_14513);
nand U14761 (N_14761,N_14501,N_14635);
or U14762 (N_14762,N_14615,N_14672);
or U14763 (N_14763,N_14729,N_14743);
or U14764 (N_14764,N_14609,N_14711);
xnor U14765 (N_14765,N_14602,N_14561);
or U14766 (N_14766,N_14598,N_14623);
nor U14767 (N_14767,N_14500,N_14721);
nand U14768 (N_14768,N_14610,N_14707);
and U14769 (N_14769,N_14744,N_14675);
and U14770 (N_14770,N_14633,N_14533);
nor U14771 (N_14771,N_14569,N_14535);
xor U14772 (N_14772,N_14730,N_14634);
or U14773 (N_14773,N_14525,N_14521);
or U14774 (N_14774,N_14660,N_14505);
nand U14775 (N_14775,N_14732,N_14550);
xnor U14776 (N_14776,N_14607,N_14617);
nand U14777 (N_14777,N_14583,N_14523);
or U14778 (N_14778,N_14592,N_14571);
nand U14779 (N_14779,N_14657,N_14670);
nand U14780 (N_14780,N_14596,N_14502);
nand U14781 (N_14781,N_14567,N_14741);
nor U14782 (N_14782,N_14518,N_14616);
and U14783 (N_14783,N_14549,N_14570);
and U14784 (N_14784,N_14629,N_14747);
and U14785 (N_14785,N_14659,N_14555);
nand U14786 (N_14786,N_14506,N_14587);
and U14787 (N_14787,N_14690,N_14710);
or U14788 (N_14788,N_14726,N_14686);
and U14789 (N_14789,N_14536,N_14544);
or U14790 (N_14790,N_14692,N_14630);
and U14791 (N_14791,N_14717,N_14621);
or U14792 (N_14792,N_14594,N_14719);
or U14793 (N_14793,N_14709,N_14539);
or U14794 (N_14794,N_14574,N_14545);
nor U14795 (N_14795,N_14632,N_14515);
and U14796 (N_14796,N_14626,N_14679);
nor U14797 (N_14797,N_14705,N_14595);
xnor U14798 (N_14798,N_14712,N_14508);
or U14799 (N_14799,N_14517,N_14674);
or U14800 (N_14800,N_14559,N_14563);
nand U14801 (N_14801,N_14601,N_14714);
xnor U14802 (N_14802,N_14669,N_14661);
or U14803 (N_14803,N_14667,N_14727);
or U14804 (N_14804,N_14586,N_14580);
nand U14805 (N_14805,N_14572,N_14560);
xnor U14806 (N_14806,N_14636,N_14694);
and U14807 (N_14807,N_14599,N_14614);
and U14808 (N_14808,N_14734,N_14564);
xnor U14809 (N_14809,N_14573,N_14650);
or U14810 (N_14810,N_14748,N_14738);
or U14811 (N_14811,N_14620,N_14579);
nand U14812 (N_14812,N_14666,N_14678);
nor U14813 (N_14813,N_14520,N_14648);
nand U14814 (N_14814,N_14558,N_14628);
nand U14815 (N_14815,N_14507,N_14649);
or U14816 (N_14816,N_14644,N_14685);
nor U14817 (N_14817,N_14673,N_14627);
nand U14818 (N_14818,N_14688,N_14514);
xor U14819 (N_14819,N_14683,N_14677);
nor U14820 (N_14820,N_14668,N_14640);
or U14821 (N_14821,N_14687,N_14735);
or U14822 (N_14822,N_14728,N_14597);
xor U14823 (N_14823,N_14691,N_14624);
xor U14824 (N_14824,N_14656,N_14566);
xor U14825 (N_14825,N_14618,N_14604);
nor U14826 (N_14826,N_14724,N_14551);
or U14827 (N_14827,N_14509,N_14611);
xnor U14828 (N_14828,N_14682,N_14642);
or U14829 (N_14829,N_14708,N_14736);
nor U14830 (N_14830,N_14622,N_14681);
nor U14831 (N_14831,N_14531,N_14749);
xor U14832 (N_14832,N_14613,N_14619);
nand U14833 (N_14833,N_14511,N_14704);
nor U14834 (N_14834,N_14742,N_14699);
xor U14835 (N_14835,N_14698,N_14541);
nand U14836 (N_14836,N_14603,N_14713);
and U14837 (N_14837,N_14655,N_14503);
nor U14838 (N_14838,N_14588,N_14577);
or U14839 (N_14839,N_14662,N_14593);
and U14840 (N_14840,N_14733,N_14582);
or U14841 (N_14841,N_14562,N_14589);
xor U14842 (N_14842,N_14532,N_14702);
or U14843 (N_14843,N_14676,N_14546);
xor U14844 (N_14844,N_14720,N_14697);
and U14845 (N_14845,N_14700,N_14645);
and U14846 (N_14846,N_14654,N_14554);
xor U14847 (N_14847,N_14581,N_14684);
xor U14848 (N_14848,N_14725,N_14680);
or U14849 (N_14849,N_14542,N_14665);
nor U14850 (N_14850,N_14600,N_14703);
nand U14851 (N_14851,N_14658,N_14540);
nor U14852 (N_14852,N_14556,N_14537);
nor U14853 (N_14853,N_14671,N_14664);
nand U14854 (N_14854,N_14519,N_14693);
or U14855 (N_14855,N_14731,N_14696);
or U14856 (N_14856,N_14716,N_14516);
xnor U14857 (N_14857,N_14528,N_14522);
xor U14858 (N_14858,N_14591,N_14510);
nor U14859 (N_14859,N_14512,N_14534);
and U14860 (N_14860,N_14526,N_14739);
and U14861 (N_14861,N_14723,N_14652);
nand U14862 (N_14862,N_14641,N_14643);
and U14863 (N_14863,N_14606,N_14575);
nand U14864 (N_14864,N_14746,N_14538);
nor U14865 (N_14865,N_14547,N_14745);
nor U14866 (N_14866,N_14718,N_14706);
nand U14867 (N_14867,N_14722,N_14568);
or U14868 (N_14868,N_14552,N_14605);
and U14869 (N_14869,N_14637,N_14631);
nor U14870 (N_14870,N_14527,N_14689);
nor U14871 (N_14871,N_14524,N_14584);
xor U14872 (N_14872,N_14715,N_14504);
or U14873 (N_14873,N_14543,N_14646);
nand U14874 (N_14874,N_14651,N_14612);
nand U14875 (N_14875,N_14585,N_14587);
or U14876 (N_14876,N_14538,N_14645);
or U14877 (N_14877,N_14586,N_14700);
nand U14878 (N_14878,N_14604,N_14718);
xnor U14879 (N_14879,N_14526,N_14536);
nor U14880 (N_14880,N_14736,N_14682);
xor U14881 (N_14881,N_14693,N_14583);
nand U14882 (N_14882,N_14500,N_14632);
and U14883 (N_14883,N_14661,N_14747);
or U14884 (N_14884,N_14536,N_14705);
xor U14885 (N_14885,N_14636,N_14523);
xnor U14886 (N_14886,N_14523,N_14616);
nor U14887 (N_14887,N_14664,N_14674);
nor U14888 (N_14888,N_14552,N_14596);
nor U14889 (N_14889,N_14535,N_14644);
or U14890 (N_14890,N_14678,N_14614);
nand U14891 (N_14891,N_14598,N_14520);
nand U14892 (N_14892,N_14730,N_14502);
nand U14893 (N_14893,N_14657,N_14674);
and U14894 (N_14894,N_14666,N_14524);
nor U14895 (N_14895,N_14627,N_14511);
or U14896 (N_14896,N_14696,N_14673);
nor U14897 (N_14897,N_14522,N_14700);
nand U14898 (N_14898,N_14608,N_14594);
nand U14899 (N_14899,N_14727,N_14500);
or U14900 (N_14900,N_14530,N_14532);
or U14901 (N_14901,N_14733,N_14609);
nand U14902 (N_14902,N_14650,N_14724);
nor U14903 (N_14903,N_14502,N_14604);
nand U14904 (N_14904,N_14512,N_14506);
or U14905 (N_14905,N_14662,N_14649);
nor U14906 (N_14906,N_14744,N_14690);
xnor U14907 (N_14907,N_14725,N_14709);
nor U14908 (N_14908,N_14717,N_14548);
or U14909 (N_14909,N_14731,N_14736);
and U14910 (N_14910,N_14717,N_14564);
xor U14911 (N_14911,N_14650,N_14545);
and U14912 (N_14912,N_14644,N_14513);
and U14913 (N_14913,N_14506,N_14649);
and U14914 (N_14914,N_14558,N_14644);
xor U14915 (N_14915,N_14623,N_14693);
nand U14916 (N_14916,N_14685,N_14672);
or U14917 (N_14917,N_14539,N_14519);
xnor U14918 (N_14918,N_14694,N_14590);
nand U14919 (N_14919,N_14695,N_14708);
nor U14920 (N_14920,N_14611,N_14534);
nand U14921 (N_14921,N_14528,N_14521);
and U14922 (N_14922,N_14604,N_14591);
xor U14923 (N_14923,N_14708,N_14697);
or U14924 (N_14924,N_14677,N_14648);
and U14925 (N_14925,N_14518,N_14640);
nand U14926 (N_14926,N_14682,N_14537);
and U14927 (N_14927,N_14526,N_14521);
nand U14928 (N_14928,N_14552,N_14553);
or U14929 (N_14929,N_14680,N_14562);
nor U14930 (N_14930,N_14695,N_14502);
nor U14931 (N_14931,N_14707,N_14615);
or U14932 (N_14932,N_14682,N_14711);
nor U14933 (N_14933,N_14726,N_14599);
or U14934 (N_14934,N_14693,N_14717);
nor U14935 (N_14935,N_14705,N_14720);
xnor U14936 (N_14936,N_14619,N_14636);
nand U14937 (N_14937,N_14662,N_14639);
nand U14938 (N_14938,N_14679,N_14515);
and U14939 (N_14939,N_14531,N_14723);
and U14940 (N_14940,N_14646,N_14558);
or U14941 (N_14941,N_14508,N_14613);
nor U14942 (N_14942,N_14734,N_14593);
nor U14943 (N_14943,N_14560,N_14599);
and U14944 (N_14944,N_14532,N_14619);
and U14945 (N_14945,N_14744,N_14595);
or U14946 (N_14946,N_14517,N_14565);
xor U14947 (N_14947,N_14542,N_14622);
and U14948 (N_14948,N_14723,N_14749);
nor U14949 (N_14949,N_14739,N_14710);
xnor U14950 (N_14950,N_14518,N_14650);
or U14951 (N_14951,N_14743,N_14553);
and U14952 (N_14952,N_14692,N_14609);
nand U14953 (N_14953,N_14675,N_14503);
nor U14954 (N_14954,N_14622,N_14513);
or U14955 (N_14955,N_14736,N_14603);
nor U14956 (N_14956,N_14636,N_14527);
or U14957 (N_14957,N_14581,N_14638);
and U14958 (N_14958,N_14632,N_14722);
xnor U14959 (N_14959,N_14611,N_14733);
nor U14960 (N_14960,N_14641,N_14527);
and U14961 (N_14961,N_14514,N_14546);
xnor U14962 (N_14962,N_14538,N_14590);
or U14963 (N_14963,N_14689,N_14531);
xor U14964 (N_14964,N_14742,N_14706);
xor U14965 (N_14965,N_14730,N_14544);
nor U14966 (N_14966,N_14541,N_14596);
xor U14967 (N_14967,N_14609,N_14641);
and U14968 (N_14968,N_14675,N_14548);
and U14969 (N_14969,N_14592,N_14521);
xnor U14970 (N_14970,N_14728,N_14570);
and U14971 (N_14971,N_14537,N_14601);
and U14972 (N_14972,N_14586,N_14726);
nand U14973 (N_14973,N_14748,N_14593);
xor U14974 (N_14974,N_14559,N_14690);
nand U14975 (N_14975,N_14512,N_14721);
nand U14976 (N_14976,N_14538,N_14741);
xor U14977 (N_14977,N_14553,N_14679);
xnor U14978 (N_14978,N_14692,N_14601);
xor U14979 (N_14979,N_14570,N_14652);
or U14980 (N_14980,N_14714,N_14571);
xor U14981 (N_14981,N_14727,N_14587);
nor U14982 (N_14982,N_14660,N_14639);
xnor U14983 (N_14983,N_14661,N_14706);
or U14984 (N_14984,N_14741,N_14705);
nand U14985 (N_14985,N_14700,N_14746);
nand U14986 (N_14986,N_14604,N_14549);
or U14987 (N_14987,N_14609,N_14732);
or U14988 (N_14988,N_14504,N_14566);
nand U14989 (N_14989,N_14738,N_14570);
and U14990 (N_14990,N_14604,N_14715);
nor U14991 (N_14991,N_14709,N_14528);
or U14992 (N_14992,N_14615,N_14556);
nand U14993 (N_14993,N_14650,N_14556);
nor U14994 (N_14994,N_14748,N_14658);
nand U14995 (N_14995,N_14590,N_14512);
nor U14996 (N_14996,N_14611,N_14500);
nor U14997 (N_14997,N_14510,N_14669);
nor U14998 (N_14998,N_14742,N_14737);
xor U14999 (N_14999,N_14556,N_14656);
xor U15000 (N_15000,N_14940,N_14991);
and U15001 (N_15001,N_14766,N_14828);
xnor U15002 (N_15002,N_14826,N_14820);
and U15003 (N_15003,N_14767,N_14960);
nor U15004 (N_15004,N_14895,N_14778);
xor U15005 (N_15005,N_14953,N_14894);
and U15006 (N_15006,N_14760,N_14815);
xnor U15007 (N_15007,N_14857,N_14817);
xnor U15008 (N_15008,N_14876,N_14919);
and U15009 (N_15009,N_14784,N_14984);
nand U15010 (N_15010,N_14750,N_14887);
nor U15011 (N_15011,N_14798,N_14934);
or U15012 (N_15012,N_14783,N_14850);
nand U15013 (N_15013,N_14928,N_14755);
xor U15014 (N_15014,N_14906,N_14879);
nor U15015 (N_15015,N_14931,N_14914);
and U15016 (N_15016,N_14909,N_14987);
or U15017 (N_15017,N_14859,N_14901);
nand U15018 (N_15018,N_14967,N_14849);
xnor U15019 (N_15019,N_14846,N_14830);
nand U15020 (N_15020,N_14860,N_14863);
or U15021 (N_15021,N_14908,N_14795);
and U15022 (N_15022,N_14982,N_14754);
xor U15023 (N_15023,N_14855,N_14833);
xnor U15024 (N_15024,N_14911,N_14980);
xor U15025 (N_15025,N_14912,N_14814);
or U15026 (N_15026,N_14944,N_14804);
and U15027 (N_15027,N_14831,N_14852);
nand U15028 (N_15028,N_14832,N_14966);
and U15029 (N_15029,N_14756,N_14921);
or U15030 (N_15030,N_14816,N_14769);
or U15031 (N_15031,N_14922,N_14770);
and U15032 (N_15032,N_14839,N_14883);
nand U15033 (N_15033,N_14990,N_14842);
and U15034 (N_15034,N_14862,N_14868);
and U15035 (N_15035,N_14943,N_14896);
nor U15036 (N_15036,N_14905,N_14771);
or U15037 (N_15037,N_14904,N_14822);
nand U15038 (N_15038,N_14981,N_14913);
nand U15039 (N_15039,N_14818,N_14992);
nor U15040 (N_15040,N_14873,N_14989);
and U15041 (N_15041,N_14971,N_14875);
nor U15042 (N_15042,N_14979,N_14917);
xor U15043 (N_15043,N_14927,N_14877);
xnor U15044 (N_15044,N_14886,N_14916);
and U15045 (N_15045,N_14952,N_14891);
nand U15046 (N_15046,N_14761,N_14938);
or U15047 (N_15047,N_14794,N_14793);
and U15048 (N_15048,N_14976,N_14752);
and U15049 (N_15049,N_14777,N_14958);
xnor U15050 (N_15050,N_14929,N_14805);
nor U15051 (N_15051,N_14969,N_14856);
xor U15052 (N_15052,N_14785,N_14951);
or U15053 (N_15053,N_14851,N_14866);
nand U15054 (N_15054,N_14803,N_14763);
xor U15055 (N_15055,N_14834,N_14937);
xor U15056 (N_15056,N_14897,N_14829);
nor U15057 (N_15057,N_14759,N_14955);
nand U15058 (N_15058,N_14776,N_14843);
or U15059 (N_15059,N_14933,N_14995);
nand U15060 (N_15060,N_14930,N_14978);
nand U15061 (N_15061,N_14920,N_14764);
or U15062 (N_15062,N_14810,N_14800);
nand U15063 (N_15063,N_14848,N_14959);
xnor U15064 (N_15064,N_14926,N_14792);
nor U15065 (N_15065,N_14972,N_14884);
nand U15066 (N_15066,N_14854,N_14789);
nor U15067 (N_15067,N_14935,N_14941);
xnor U15068 (N_15068,N_14903,N_14924);
and U15069 (N_15069,N_14998,N_14880);
or U15070 (N_15070,N_14845,N_14946);
nand U15071 (N_15071,N_14964,N_14945);
nand U15072 (N_15072,N_14821,N_14762);
xor U15073 (N_15073,N_14819,N_14807);
xor U15074 (N_15074,N_14915,N_14988);
or U15075 (N_15075,N_14888,N_14806);
nand U15076 (N_15076,N_14936,N_14753);
nor U15077 (N_15077,N_14882,N_14965);
nor U15078 (N_15078,N_14932,N_14977);
xor U15079 (N_15079,N_14768,N_14892);
nand U15080 (N_15080,N_14962,N_14837);
nand U15081 (N_15081,N_14782,N_14900);
nand U15082 (N_15082,N_14994,N_14786);
or U15083 (N_15083,N_14775,N_14847);
nor U15084 (N_15084,N_14881,N_14864);
or U15085 (N_15085,N_14893,N_14779);
xnor U15086 (N_15086,N_14918,N_14996);
or U15087 (N_15087,N_14954,N_14899);
and U15088 (N_15088,N_14950,N_14885);
and U15089 (N_15089,N_14808,N_14898);
nor U15090 (N_15090,N_14802,N_14948);
or U15091 (N_15091,N_14986,N_14983);
or U15092 (N_15092,N_14809,N_14751);
xor U15093 (N_15093,N_14907,N_14773);
nand U15094 (N_15094,N_14844,N_14811);
nand U15095 (N_15095,N_14925,N_14957);
xnor U15096 (N_15096,N_14947,N_14942);
nor U15097 (N_15097,N_14801,N_14780);
and U15098 (N_15098,N_14824,N_14867);
nor U15099 (N_15099,N_14865,N_14796);
and U15100 (N_15100,N_14889,N_14825);
nand U15101 (N_15101,N_14974,N_14853);
and U15102 (N_15102,N_14788,N_14787);
xor U15103 (N_15103,N_14997,N_14812);
nand U15104 (N_15104,N_14823,N_14874);
xor U15105 (N_15105,N_14975,N_14758);
nor U15106 (N_15106,N_14871,N_14999);
and U15107 (N_15107,N_14968,N_14993);
nand U15108 (N_15108,N_14949,N_14791);
nor U15109 (N_15109,N_14910,N_14838);
or U15110 (N_15110,N_14790,N_14970);
xnor U15111 (N_15111,N_14939,N_14878);
nand U15112 (N_15112,N_14813,N_14840);
nor U15113 (N_15113,N_14923,N_14890);
nor U15114 (N_15114,N_14869,N_14870);
nand U15115 (N_15115,N_14872,N_14858);
nand U15116 (N_15116,N_14781,N_14836);
or U15117 (N_15117,N_14772,N_14956);
or U15118 (N_15118,N_14765,N_14973);
and U15119 (N_15119,N_14985,N_14799);
xnor U15120 (N_15120,N_14835,N_14757);
nand U15121 (N_15121,N_14861,N_14774);
xnor U15122 (N_15122,N_14841,N_14797);
nand U15123 (N_15123,N_14827,N_14902);
or U15124 (N_15124,N_14963,N_14961);
nand U15125 (N_15125,N_14841,N_14848);
xor U15126 (N_15126,N_14927,N_14798);
nand U15127 (N_15127,N_14994,N_14984);
and U15128 (N_15128,N_14842,N_14872);
nor U15129 (N_15129,N_14771,N_14976);
or U15130 (N_15130,N_14889,N_14955);
or U15131 (N_15131,N_14853,N_14772);
xor U15132 (N_15132,N_14851,N_14971);
nor U15133 (N_15133,N_14878,N_14999);
nor U15134 (N_15134,N_14928,N_14831);
nand U15135 (N_15135,N_14757,N_14922);
nand U15136 (N_15136,N_14895,N_14913);
xor U15137 (N_15137,N_14942,N_14796);
nor U15138 (N_15138,N_14959,N_14935);
nor U15139 (N_15139,N_14987,N_14935);
nand U15140 (N_15140,N_14762,N_14843);
and U15141 (N_15141,N_14776,N_14855);
xnor U15142 (N_15142,N_14894,N_14917);
and U15143 (N_15143,N_14856,N_14948);
and U15144 (N_15144,N_14770,N_14979);
xor U15145 (N_15145,N_14964,N_14985);
nand U15146 (N_15146,N_14938,N_14847);
nand U15147 (N_15147,N_14837,N_14752);
nor U15148 (N_15148,N_14812,N_14909);
nand U15149 (N_15149,N_14931,N_14869);
nand U15150 (N_15150,N_14868,N_14824);
and U15151 (N_15151,N_14756,N_14822);
nand U15152 (N_15152,N_14782,N_14854);
nor U15153 (N_15153,N_14882,N_14917);
nor U15154 (N_15154,N_14818,N_14895);
or U15155 (N_15155,N_14895,N_14928);
nand U15156 (N_15156,N_14822,N_14858);
nor U15157 (N_15157,N_14927,N_14780);
nor U15158 (N_15158,N_14862,N_14974);
nor U15159 (N_15159,N_14902,N_14994);
nor U15160 (N_15160,N_14757,N_14806);
and U15161 (N_15161,N_14805,N_14855);
nor U15162 (N_15162,N_14897,N_14809);
xor U15163 (N_15163,N_14916,N_14901);
nand U15164 (N_15164,N_14894,N_14819);
and U15165 (N_15165,N_14820,N_14867);
or U15166 (N_15166,N_14778,N_14764);
or U15167 (N_15167,N_14845,N_14931);
xor U15168 (N_15168,N_14909,N_14824);
nor U15169 (N_15169,N_14869,N_14751);
and U15170 (N_15170,N_14787,N_14786);
xor U15171 (N_15171,N_14911,N_14832);
nor U15172 (N_15172,N_14818,N_14839);
xnor U15173 (N_15173,N_14988,N_14846);
and U15174 (N_15174,N_14987,N_14778);
nand U15175 (N_15175,N_14836,N_14882);
xor U15176 (N_15176,N_14958,N_14886);
or U15177 (N_15177,N_14952,N_14896);
nand U15178 (N_15178,N_14921,N_14765);
nand U15179 (N_15179,N_14825,N_14789);
or U15180 (N_15180,N_14757,N_14911);
xor U15181 (N_15181,N_14789,N_14956);
nand U15182 (N_15182,N_14946,N_14788);
or U15183 (N_15183,N_14929,N_14837);
nand U15184 (N_15184,N_14776,N_14938);
nand U15185 (N_15185,N_14950,N_14907);
and U15186 (N_15186,N_14967,N_14909);
and U15187 (N_15187,N_14940,N_14793);
or U15188 (N_15188,N_14935,N_14769);
nor U15189 (N_15189,N_14981,N_14817);
or U15190 (N_15190,N_14960,N_14894);
nand U15191 (N_15191,N_14806,N_14892);
nand U15192 (N_15192,N_14972,N_14800);
or U15193 (N_15193,N_14761,N_14933);
nand U15194 (N_15194,N_14911,N_14768);
nor U15195 (N_15195,N_14780,N_14942);
nor U15196 (N_15196,N_14863,N_14876);
or U15197 (N_15197,N_14880,N_14866);
nor U15198 (N_15198,N_14968,N_14857);
and U15199 (N_15199,N_14964,N_14857);
nor U15200 (N_15200,N_14929,N_14788);
nand U15201 (N_15201,N_14776,N_14753);
xor U15202 (N_15202,N_14910,N_14985);
nand U15203 (N_15203,N_14961,N_14934);
nand U15204 (N_15204,N_14842,N_14903);
xnor U15205 (N_15205,N_14784,N_14799);
nor U15206 (N_15206,N_14791,N_14939);
nand U15207 (N_15207,N_14806,N_14765);
xor U15208 (N_15208,N_14896,N_14779);
nand U15209 (N_15209,N_14841,N_14778);
nor U15210 (N_15210,N_14801,N_14913);
nand U15211 (N_15211,N_14960,N_14931);
xnor U15212 (N_15212,N_14906,N_14848);
and U15213 (N_15213,N_14772,N_14854);
nand U15214 (N_15214,N_14891,N_14833);
or U15215 (N_15215,N_14882,N_14991);
xor U15216 (N_15216,N_14812,N_14980);
xor U15217 (N_15217,N_14911,N_14845);
or U15218 (N_15218,N_14999,N_14799);
and U15219 (N_15219,N_14920,N_14977);
and U15220 (N_15220,N_14776,N_14927);
or U15221 (N_15221,N_14805,N_14815);
nor U15222 (N_15222,N_14915,N_14930);
nand U15223 (N_15223,N_14986,N_14775);
nand U15224 (N_15224,N_14932,N_14844);
or U15225 (N_15225,N_14941,N_14978);
nor U15226 (N_15226,N_14888,N_14869);
xor U15227 (N_15227,N_14966,N_14827);
nor U15228 (N_15228,N_14771,N_14896);
nand U15229 (N_15229,N_14837,N_14755);
or U15230 (N_15230,N_14777,N_14834);
nor U15231 (N_15231,N_14773,N_14868);
nand U15232 (N_15232,N_14899,N_14752);
nor U15233 (N_15233,N_14867,N_14810);
nand U15234 (N_15234,N_14899,N_14916);
xnor U15235 (N_15235,N_14885,N_14828);
nand U15236 (N_15236,N_14824,N_14765);
nor U15237 (N_15237,N_14770,N_14859);
and U15238 (N_15238,N_14890,N_14962);
nor U15239 (N_15239,N_14796,N_14937);
and U15240 (N_15240,N_14946,N_14979);
or U15241 (N_15241,N_14814,N_14864);
nand U15242 (N_15242,N_14877,N_14942);
nand U15243 (N_15243,N_14775,N_14773);
xor U15244 (N_15244,N_14864,N_14910);
and U15245 (N_15245,N_14960,N_14884);
and U15246 (N_15246,N_14821,N_14961);
nand U15247 (N_15247,N_14826,N_14917);
and U15248 (N_15248,N_14965,N_14950);
or U15249 (N_15249,N_14840,N_14971);
or U15250 (N_15250,N_15216,N_15223);
or U15251 (N_15251,N_15039,N_15117);
nand U15252 (N_15252,N_15221,N_15029);
and U15253 (N_15253,N_15175,N_15178);
xor U15254 (N_15254,N_15053,N_15046);
or U15255 (N_15255,N_15222,N_15112);
and U15256 (N_15256,N_15094,N_15086);
or U15257 (N_15257,N_15027,N_15061);
and U15258 (N_15258,N_15241,N_15113);
and U15259 (N_15259,N_15049,N_15203);
nor U15260 (N_15260,N_15197,N_15167);
and U15261 (N_15261,N_15065,N_15147);
xor U15262 (N_15262,N_15108,N_15236);
xor U15263 (N_15263,N_15083,N_15028);
and U15264 (N_15264,N_15063,N_15023);
nor U15265 (N_15265,N_15201,N_15106);
nand U15266 (N_15266,N_15180,N_15124);
xor U15267 (N_15267,N_15032,N_15107);
or U15268 (N_15268,N_15099,N_15170);
or U15269 (N_15269,N_15037,N_15096);
nand U15270 (N_15270,N_15205,N_15013);
xnor U15271 (N_15271,N_15076,N_15231);
and U15272 (N_15272,N_15152,N_15213);
nor U15273 (N_15273,N_15082,N_15142);
xnor U15274 (N_15274,N_15204,N_15101);
xor U15275 (N_15275,N_15200,N_15026);
and U15276 (N_15276,N_15169,N_15234);
nor U15277 (N_15277,N_15041,N_15121);
xnor U15278 (N_15278,N_15186,N_15244);
xnor U15279 (N_15279,N_15220,N_15055);
or U15280 (N_15280,N_15181,N_15034);
nand U15281 (N_15281,N_15102,N_15016);
nand U15282 (N_15282,N_15182,N_15093);
nor U15283 (N_15283,N_15163,N_15162);
or U15284 (N_15284,N_15062,N_15024);
and U15285 (N_15285,N_15010,N_15044);
nand U15286 (N_15286,N_15144,N_15068);
and U15287 (N_15287,N_15080,N_15136);
xor U15288 (N_15288,N_15095,N_15226);
nand U15289 (N_15289,N_15059,N_15211);
and U15290 (N_15290,N_15020,N_15155);
nor U15291 (N_15291,N_15171,N_15189);
nand U15292 (N_15292,N_15057,N_15176);
or U15293 (N_15293,N_15100,N_15103);
nand U15294 (N_15294,N_15067,N_15038);
and U15295 (N_15295,N_15237,N_15151);
xor U15296 (N_15296,N_15021,N_15025);
nor U15297 (N_15297,N_15130,N_15156);
and U15298 (N_15298,N_15173,N_15132);
nand U15299 (N_15299,N_15116,N_15247);
xnor U15300 (N_15300,N_15225,N_15122);
nand U15301 (N_15301,N_15232,N_15000);
or U15302 (N_15302,N_15177,N_15126);
nor U15303 (N_15303,N_15030,N_15114);
and U15304 (N_15304,N_15207,N_15085);
or U15305 (N_15305,N_15127,N_15192);
or U15306 (N_15306,N_15139,N_15091);
or U15307 (N_15307,N_15157,N_15002);
xnor U15308 (N_15308,N_15092,N_15145);
or U15309 (N_15309,N_15081,N_15185);
xnor U15310 (N_15310,N_15078,N_15218);
and U15311 (N_15311,N_15131,N_15150);
and U15312 (N_15312,N_15123,N_15184);
and U15313 (N_15313,N_15054,N_15249);
nand U15314 (N_15314,N_15210,N_15235);
and U15315 (N_15315,N_15153,N_15073);
nor U15316 (N_15316,N_15109,N_15069);
xnor U15317 (N_15317,N_15036,N_15051);
and U15318 (N_15318,N_15140,N_15209);
nand U15319 (N_15319,N_15005,N_15008);
nor U15320 (N_15320,N_15042,N_15227);
and U15321 (N_15321,N_15017,N_15164);
or U15322 (N_15322,N_15168,N_15084);
nor U15323 (N_15323,N_15007,N_15208);
or U15324 (N_15324,N_15075,N_15001);
or U15325 (N_15325,N_15072,N_15159);
nand U15326 (N_15326,N_15110,N_15154);
nor U15327 (N_15327,N_15228,N_15187);
nor U15328 (N_15328,N_15012,N_15141);
xor U15329 (N_15329,N_15148,N_15104);
and U15330 (N_15330,N_15089,N_15233);
nor U15331 (N_15331,N_15011,N_15158);
xnor U15332 (N_15332,N_15190,N_15242);
nor U15333 (N_15333,N_15120,N_15060);
and U15334 (N_15334,N_15217,N_15058);
nor U15335 (N_15335,N_15191,N_15047);
xnor U15336 (N_15336,N_15193,N_15077);
or U15337 (N_15337,N_15087,N_15143);
or U15338 (N_15338,N_15071,N_15019);
nor U15339 (N_15339,N_15230,N_15199);
nor U15340 (N_15340,N_15194,N_15219);
or U15341 (N_15341,N_15105,N_15212);
nand U15342 (N_15342,N_15043,N_15248);
nand U15343 (N_15343,N_15243,N_15166);
xor U15344 (N_15344,N_15195,N_15035);
and U15345 (N_15345,N_15245,N_15006);
nand U15346 (N_15346,N_15135,N_15056);
xnor U15347 (N_15347,N_15224,N_15125);
nand U15348 (N_15348,N_15188,N_15138);
or U15349 (N_15349,N_15240,N_15066);
nor U15350 (N_15350,N_15014,N_15196);
xor U15351 (N_15351,N_15050,N_15048);
xor U15352 (N_15352,N_15238,N_15202);
xor U15353 (N_15353,N_15045,N_15133);
or U15354 (N_15354,N_15137,N_15229);
or U15355 (N_15355,N_15097,N_15239);
or U15356 (N_15356,N_15206,N_15018);
nand U15357 (N_15357,N_15015,N_15246);
nand U15358 (N_15358,N_15033,N_15128);
xor U15359 (N_15359,N_15115,N_15214);
nand U15360 (N_15360,N_15161,N_15118);
and U15361 (N_15361,N_15064,N_15215);
nor U15362 (N_15362,N_15052,N_15074);
nor U15363 (N_15363,N_15088,N_15079);
or U15364 (N_15364,N_15022,N_15149);
nor U15365 (N_15365,N_15009,N_15119);
nand U15366 (N_15366,N_15004,N_15160);
and U15367 (N_15367,N_15134,N_15174);
or U15368 (N_15368,N_15172,N_15146);
or U15369 (N_15369,N_15003,N_15183);
nor U15370 (N_15370,N_15165,N_15070);
xnor U15371 (N_15371,N_15129,N_15198);
or U15372 (N_15372,N_15090,N_15040);
and U15373 (N_15373,N_15111,N_15098);
xnor U15374 (N_15374,N_15179,N_15031);
or U15375 (N_15375,N_15084,N_15000);
nor U15376 (N_15376,N_15022,N_15061);
xor U15377 (N_15377,N_15197,N_15100);
xor U15378 (N_15378,N_15183,N_15047);
nor U15379 (N_15379,N_15200,N_15096);
nand U15380 (N_15380,N_15001,N_15053);
and U15381 (N_15381,N_15103,N_15131);
or U15382 (N_15382,N_15198,N_15245);
or U15383 (N_15383,N_15129,N_15083);
nand U15384 (N_15384,N_15076,N_15178);
nor U15385 (N_15385,N_15071,N_15133);
and U15386 (N_15386,N_15206,N_15061);
nor U15387 (N_15387,N_15173,N_15025);
nor U15388 (N_15388,N_15157,N_15010);
and U15389 (N_15389,N_15022,N_15082);
or U15390 (N_15390,N_15226,N_15170);
and U15391 (N_15391,N_15149,N_15231);
nor U15392 (N_15392,N_15193,N_15114);
nor U15393 (N_15393,N_15166,N_15144);
and U15394 (N_15394,N_15186,N_15231);
or U15395 (N_15395,N_15077,N_15053);
or U15396 (N_15396,N_15030,N_15248);
and U15397 (N_15397,N_15174,N_15142);
xnor U15398 (N_15398,N_15011,N_15018);
nand U15399 (N_15399,N_15041,N_15152);
xor U15400 (N_15400,N_15077,N_15061);
nand U15401 (N_15401,N_15153,N_15053);
xor U15402 (N_15402,N_15113,N_15027);
nand U15403 (N_15403,N_15206,N_15022);
nand U15404 (N_15404,N_15070,N_15143);
xnor U15405 (N_15405,N_15024,N_15176);
nand U15406 (N_15406,N_15024,N_15035);
nor U15407 (N_15407,N_15019,N_15151);
xor U15408 (N_15408,N_15214,N_15116);
nor U15409 (N_15409,N_15073,N_15006);
nor U15410 (N_15410,N_15162,N_15104);
and U15411 (N_15411,N_15007,N_15096);
nand U15412 (N_15412,N_15178,N_15198);
nor U15413 (N_15413,N_15006,N_15207);
nor U15414 (N_15414,N_15085,N_15077);
nand U15415 (N_15415,N_15141,N_15109);
and U15416 (N_15416,N_15041,N_15172);
xnor U15417 (N_15417,N_15104,N_15208);
nand U15418 (N_15418,N_15030,N_15121);
nor U15419 (N_15419,N_15215,N_15084);
nor U15420 (N_15420,N_15020,N_15246);
or U15421 (N_15421,N_15090,N_15175);
nand U15422 (N_15422,N_15189,N_15042);
or U15423 (N_15423,N_15072,N_15240);
nand U15424 (N_15424,N_15140,N_15088);
or U15425 (N_15425,N_15140,N_15221);
nor U15426 (N_15426,N_15036,N_15111);
xnor U15427 (N_15427,N_15160,N_15041);
nor U15428 (N_15428,N_15081,N_15215);
and U15429 (N_15429,N_15086,N_15153);
and U15430 (N_15430,N_15245,N_15099);
nor U15431 (N_15431,N_15012,N_15122);
xor U15432 (N_15432,N_15116,N_15217);
or U15433 (N_15433,N_15227,N_15209);
or U15434 (N_15434,N_15002,N_15007);
and U15435 (N_15435,N_15021,N_15049);
and U15436 (N_15436,N_15052,N_15045);
nor U15437 (N_15437,N_15084,N_15092);
nand U15438 (N_15438,N_15218,N_15192);
nand U15439 (N_15439,N_15154,N_15063);
xnor U15440 (N_15440,N_15108,N_15057);
or U15441 (N_15441,N_15240,N_15095);
nor U15442 (N_15442,N_15207,N_15129);
nor U15443 (N_15443,N_15201,N_15233);
xor U15444 (N_15444,N_15111,N_15051);
or U15445 (N_15445,N_15110,N_15115);
xnor U15446 (N_15446,N_15044,N_15009);
nand U15447 (N_15447,N_15043,N_15080);
and U15448 (N_15448,N_15080,N_15022);
or U15449 (N_15449,N_15245,N_15113);
nor U15450 (N_15450,N_15123,N_15020);
and U15451 (N_15451,N_15030,N_15219);
nand U15452 (N_15452,N_15013,N_15174);
nand U15453 (N_15453,N_15108,N_15113);
and U15454 (N_15454,N_15217,N_15119);
nand U15455 (N_15455,N_15100,N_15136);
nor U15456 (N_15456,N_15191,N_15204);
and U15457 (N_15457,N_15177,N_15081);
xnor U15458 (N_15458,N_15201,N_15194);
or U15459 (N_15459,N_15051,N_15054);
and U15460 (N_15460,N_15096,N_15177);
and U15461 (N_15461,N_15006,N_15080);
nor U15462 (N_15462,N_15243,N_15163);
nand U15463 (N_15463,N_15145,N_15069);
and U15464 (N_15464,N_15220,N_15076);
or U15465 (N_15465,N_15077,N_15133);
or U15466 (N_15466,N_15048,N_15210);
nand U15467 (N_15467,N_15008,N_15242);
and U15468 (N_15468,N_15091,N_15216);
xnor U15469 (N_15469,N_15172,N_15170);
nor U15470 (N_15470,N_15217,N_15083);
or U15471 (N_15471,N_15017,N_15245);
xor U15472 (N_15472,N_15234,N_15240);
nor U15473 (N_15473,N_15142,N_15019);
and U15474 (N_15474,N_15137,N_15086);
or U15475 (N_15475,N_15249,N_15047);
nor U15476 (N_15476,N_15083,N_15088);
nor U15477 (N_15477,N_15213,N_15041);
and U15478 (N_15478,N_15058,N_15156);
and U15479 (N_15479,N_15120,N_15233);
or U15480 (N_15480,N_15123,N_15136);
nor U15481 (N_15481,N_15080,N_15153);
nand U15482 (N_15482,N_15102,N_15071);
nor U15483 (N_15483,N_15222,N_15078);
xnor U15484 (N_15484,N_15160,N_15239);
or U15485 (N_15485,N_15171,N_15144);
nand U15486 (N_15486,N_15121,N_15215);
nand U15487 (N_15487,N_15096,N_15197);
xor U15488 (N_15488,N_15223,N_15129);
or U15489 (N_15489,N_15230,N_15163);
nor U15490 (N_15490,N_15057,N_15087);
xor U15491 (N_15491,N_15115,N_15188);
nand U15492 (N_15492,N_15218,N_15025);
and U15493 (N_15493,N_15008,N_15148);
or U15494 (N_15494,N_15156,N_15096);
nor U15495 (N_15495,N_15035,N_15132);
xor U15496 (N_15496,N_15036,N_15002);
xor U15497 (N_15497,N_15084,N_15099);
or U15498 (N_15498,N_15053,N_15113);
xor U15499 (N_15499,N_15148,N_15069);
nor U15500 (N_15500,N_15377,N_15297);
or U15501 (N_15501,N_15424,N_15455);
and U15502 (N_15502,N_15443,N_15320);
nor U15503 (N_15503,N_15368,N_15394);
and U15504 (N_15504,N_15416,N_15338);
nand U15505 (N_15505,N_15286,N_15303);
xnor U15506 (N_15506,N_15420,N_15433);
xor U15507 (N_15507,N_15415,N_15289);
xor U15508 (N_15508,N_15288,N_15285);
xnor U15509 (N_15509,N_15466,N_15492);
and U15510 (N_15510,N_15306,N_15442);
nand U15511 (N_15511,N_15490,N_15463);
nand U15512 (N_15512,N_15349,N_15421);
xor U15513 (N_15513,N_15400,N_15282);
xnor U15514 (N_15514,N_15329,N_15346);
nor U15515 (N_15515,N_15301,N_15339);
xnor U15516 (N_15516,N_15360,N_15348);
nand U15517 (N_15517,N_15292,N_15486);
or U15518 (N_15518,N_15497,N_15384);
nor U15519 (N_15519,N_15444,N_15454);
and U15520 (N_15520,N_15399,N_15371);
nand U15521 (N_15521,N_15276,N_15491);
and U15522 (N_15522,N_15388,N_15480);
nand U15523 (N_15523,N_15322,N_15387);
nor U15524 (N_15524,N_15418,N_15493);
nand U15525 (N_15525,N_15447,N_15417);
and U15526 (N_15526,N_15390,N_15494);
nor U15527 (N_15527,N_15355,N_15314);
and U15528 (N_15528,N_15337,N_15482);
xor U15529 (N_15529,N_15254,N_15471);
nand U15530 (N_15530,N_15311,N_15495);
xnor U15531 (N_15531,N_15336,N_15462);
nor U15532 (N_15532,N_15344,N_15259);
or U15533 (N_15533,N_15460,N_15313);
xor U15534 (N_15534,N_15253,N_15470);
nor U15535 (N_15535,N_15307,N_15275);
or U15536 (N_15536,N_15333,N_15278);
nand U15537 (N_15537,N_15427,N_15317);
xnor U15538 (N_15538,N_15391,N_15332);
nand U15539 (N_15539,N_15294,N_15284);
nor U15540 (N_15540,N_15477,N_15252);
or U15541 (N_15541,N_15459,N_15476);
xnor U15542 (N_15542,N_15258,N_15413);
nor U15543 (N_15543,N_15488,N_15315);
or U15544 (N_15544,N_15410,N_15283);
nor U15545 (N_15545,N_15481,N_15381);
nand U15546 (N_15546,N_15395,N_15370);
xor U15547 (N_15547,N_15251,N_15450);
xor U15548 (N_15548,N_15255,N_15266);
xnor U15549 (N_15549,N_15318,N_15375);
and U15550 (N_15550,N_15457,N_15334);
nor U15551 (N_15551,N_15468,N_15365);
nor U15552 (N_15552,N_15354,N_15484);
xor U15553 (N_15553,N_15403,N_15352);
xnor U15554 (N_15554,N_15472,N_15369);
nand U15555 (N_15555,N_15386,N_15270);
or U15556 (N_15556,N_15341,N_15478);
nor U15557 (N_15557,N_15498,N_15487);
xor U15558 (N_15558,N_15308,N_15330);
and U15559 (N_15559,N_15483,N_15357);
xnor U15560 (N_15560,N_15411,N_15452);
nand U15561 (N_15561,N_15437,N_15319);
or U15562 (N_15562,N_15309,N_15279);
and U15563 (N_15563,N_15304,N_15268);
or U15564 (N_15564,N_15456,N_15479);
and U15565 (N_15565,N_15287,N_15373);
or U15566 (N_15566,N_15428,N_15412);
or U15567 (N_15567,N_15299,N_15280);
xnor U15568 (N_15568,N_15445,N_15439);
and U15569 (N_15569,N_15359,N_15324);
and U15570 (N_15570,N_15271,N_15353);
nand U15571 (N_15571,N_15300,N_15298);
nor U15572 (N_15572,N_15465,N_15408);
and U15573 (N_15573,N_15293,N_15406);
nand U15574 (N_15574,N_15310,N_15265);
nand U15575 (N_15575,N_15385,N_15389);
and U15576 (N_15576,N_15434,N_15342);
or U15577 (N_15577,N_15264,N_15383);
nand U15578 (N_15578,N_15414,N_15347);
xnor U15579 (N_15579,N_15404,N_15327);
xnor U15580 (N_15580,N_15393,N_15453);
nand U15581 (N_15581,N_15407,N_15379);
nor U15582 (N_15582,N_15267,N_15296);
nand U15583 (N_15583,N_15475,N_15363);
xor U15584 (N_15584,N_15358,N_15473);
or U15585 (N_15585,N_15323,N_15260);
or U15586 (N_15586,N_15446,N_15273);
xor U15587 (N_15587,N_15438,N_15392);
nor U15588 (N_15588,N_15325,N_15351);
or U15589 (N_15589,N_15419,N_15489);
nor U15590 (N_15590,N_15440,N_15356);
xor U15591 (N_15591,N_15382,N_15425);
nor U15592 (N_15592,N_15361,N_15262);
and U15593 (N_15593,N_15272,N_15461);
and U15594 (N_15594,N_15485,N_15441);
or U15595 (N_15595,N_15367,N_15467);
xor U15596 (N_15596,N_15269,N_15448);
and U15597 (N_15597,N_15432,N_15295);
nand U15598 (N_15598,N_15374,N_15364);
and U15599 (N_15599,N_15340,N_15256);
xnor U15600 (N_15600,N_15312,N_15261);
nor U15601 (N_15601,N_15499,N_15328);
nor U15602 (N_15602,N_15401,N_15496);
or U15603 (N_15603,N_15376,N_15305);
and U15604 (N_15604,N_15343,N_15263);
or U15605 (N_15605,N_15316,N_15449);
xor U15606 (N_15606,N_15431,N_15451);
or U15607 (N_15607,N_15435,N_15396);
nor U15608 (N_15608,N_15291,N_15430);
xor U15609 (N_15609,N_15350,N_15372);
xnor U15610 (N_15610,N_15345,N_15326);
or U15611 (N_15611,N_15464,N_15380);
nand U15612 (N_15612,N_15405,N_15422);
or U15613 (N_15613,N_15426,N_15429);
nand U15614 (N_15614,N_15366,N_15423);
xnor U15615 (N_15615,N_15281,N_15362);
or U15616 (N_15616,N_15257,N_15274);
nand U15617 (N_15617,N_15397,N_15290);
nand U15618 (N_15618,N_15335,N_15321);
nor U15619 (N_15619,N_15378,N_15436);
and U15620 (N_15620,N_15277,N_15402);
nand U15621 (N_15621,N_15474,N_15469);
nor U15622 (N_15622,N_15331,N_15458);
or U15623 (N_15623,N_15409,N_15398);
or U15624 (N_15624,N_15302,N_15250);
or U15625 (N_15625,N_15337,N_15428);
or U15626 (N_15626,N_15286,N_15370);
and U15627 (N_15627,N_15364,N_15400);
xnor U15628 (N_15628,N_15378,N_15300);
nor U15629 (N_15629,N_15333,N_15343);
and U15630 (N_15630,N_15372,N_15445);
or U15631 (N_15631,N_15401,N_15493);
or U15632 (N_15632,N_15423,N_15387);
and U15633 (N_15633,N_15302,N_15366);
and U15634 (N_15634,N_15469,N_15417);
and U15635 (N_15635,N_15420,N_15253);
xnor U15636 (N_15636,N_15279,N_15271);
nor U15637 (N_15637,N_15405,N_15319);
xor U15638 (N_15638,N_15428,N_15370);
and U15639 (N_15639,N_15395,N_15353);
nor U15640 (N_15640,N_15295,N_15474);
and U15641 (N_15641,N_15330,N_15372);
nand U15642 (N_15642,N_15437,N_15379);
or U15643 (N_15643,N_15375,N_15365);
or U15644 (N_15644,N_15385,N_15272);
and U15645 (N_15645,N_15416,N_15415);
and U15646 (N_15646,N_15296,N_15390);
and U15647 (N_15647,N_15315,N_15259);
xnor U15648 (N_15648,N_15303,N_15486);
nand U15649 (N_15649,N_15377,N_15286);
and U15650 (N_15650,N_15458,N_15385);
or U15651 (N_15651,N_15302,N_15318);
nand U15652 (N_15652,N_15302,N_15473);
xor U15653 (N_15653,N_15470,N_15488);
and U15654 (N_15654,N_15444,N_15292);
nand U15655 (N_15655,N_15384,N_15446);
and U15656 (N_15656,N_15464,N_15431);
and U15657 (N_15657,N_15428,N_15252);
xnor U15658 (N_15658,N_15358,N_15465);
nor U15659 (N_15659,N_15429,N_15288);
xnor U15660 (N_15660,N_15321,N_15491);
or U15661 (N_15661,N_15363,N_15369);
and U15662 (N_15662,N_15345,N_15429);
and U15663 (N_15663,N_15415,N_15381);
xor U15664 (N_15664,N_15422,N_15350);
nand U15665 (N_15665,N_15466,N_15499);
or U15666 (N_15666,N_15252,N_15276);
and U15667 (N_15667,N_15472,N_15351);
xnor U15668 (N_15668,N_15409,N_15483);
or U15669 (N_15669,N_15399,N_15495);
nand U15670 (N_15670,N_15273,N_15345);
or U15671 (N_15671,N_15252,N_15338);
nand U15672 (N_15672,N_15331,N_15318);
nand U15673 (N_15673,N_15451,N_15280);
and U15674 (N_15674,N_15469,N_15491);
or U15675 (N_15675,N_15393,N_15495);
nor U15676 (N_15676,N_15334,N_15286);
nor U15677 (N_15677,N_15367,N_15364);
and U15678 (N_15678,N_15272,N_15416);
nand U15679 (N_15679,N_15366,N_15489);
xor U15680 (N_15680,N_15446,N_15478);
nand U15681 (N_15681,N_15419,N_15266);
nor U15682 (N_15682,N_15387,N_15372);
nand U15683 (N_15683,N_15259,N_15441);
and U15684 (N_15684,N_15431,N_15428);
and U15685 (N_15685,N_15479,N_15275);
or U15686 (N_15686,N_15312,N_15419);
nor U15687 (N_15687,N_15294,N_15254);
and U15688 (N_15688,N_15262,N_15381);
nor U15689 (N_15689,N_15258,N_15261);
nor U15690 (N_15690,N_15364,N_15451);
or U15691 (N_15691,N_15482,N_15464);
nor U15692 (N_15692,N_15346,N_15477);
and U15693 (N_15693,N_15263,N_15331);
and U15694 (N_15694,N_15471,N_15357);
xor U15695 (N_15695,N_15258,N_15252);
xor U15696 (N_15696,N_15305,N_15476);
or U15697 (N_15697,N_15297,N_15404);
xnor U15698 (N_15698,N_15382,N_15469);
nand U15699 (N_15699,N_15285,N_15364);
xor U15700 (N_15700,N_15476,N_15351);
xor U15701 (N_15701,N_15434,N_15423);
and U15702 (N_15702,N_15462,N_15385);
and U15703 (N_15703,N_15425,N_15350);
nand U15704 (N_15704,N_15474,N_15457);
or U15705 (N_15705,N_15477,N_15259);
nand U15706 (N_15706,N_15276,N_15292);
and U15707 (N_15707,N_15395,N_15303);
nand U15708 (N_15708,N_15414,N_15312);
nand U15709 (N_15709,N_15409,N_15495);
or U15710 (N_15710,N_15314,N_15324);
nand U15711 (N_15711,N_15488,N_15416);
nor U15712 (N_15712,N_15261,N_15406);
nand U15713 (N_15713,N_15303,N_15406);
xnor U15714 (N_15714,N_15456,N_15468);
or U15715 (N_15715,N_15311,N_15498);
xor U15716 (N_15716,N_15255,N_15394);
nand U15717 (N_15717,N_15251,N_15424);
nor U15718 (N_15718,N_15280,N_15330);
xnor U15719 (N_15719,N_15402,N_15467);
and U15720 (N_15720,N_15374,N_15337);
nor U15721 (N_15721,N_15421,N_15405);
or U15722 (N_15722,N_15293,N_15330);
nand U15723 (N_15723,N_15438,N_15477);
nand U15724 (N_15724,N_15484,N_15442);
and U15725 (N_15725,N_15464,N_15426);
nor U15726 (N_15726,N_15283,N_15384);
or U15727 (N_15727,N_15404,N_15257);
or U15728 (N_15728,N_15300,N_15376);
and U15729 (N_15729,N_15317,N_15324);
xor U15730 (N_15730,N_15319,N_15446);
nor U15731 (N_15731,N_15304,N_15496);
xor U15732 (N_15732,N_15436,N_15486);
nor U15733 (N_15733,N_15486,N_15480);
and U15734 (N_15734,N_15477,N_15400);
or U15735 (N_15735,N_15338,N_15486);
and U15736 (N_15736,N_15322,N_15290);
and U15737 (N_15737,N_15305,N_15491);
xnor U15738 (N_15738,N_15292,N_15469);
nor U15739 (N_15739,N_15340,N_15351);
and U15740 (N_15740,N_15493,N_15412);
and U15741 (N_15741,N_15421,N_15493);
nand U15742 (N_15742,N_15393,N_15251);
nor U15743 (N_15743,N_15489,N_15257);
xor U15744 (N_15744,N_15471,N_15386);
nand U15745 (N_15745,N_15389,N_15317);
nand U15746 (N_15746,N_15487,N_15316);
nand U15747 (N_15747,N_15436,N_15406);
and U15748 (N_15748,N_15268,N_15464);
xor U15749 (N_15749,N_15315,N_15375);
or U15750 (N_15750,N_15722,N_15589);
or U15751 (N_15751,N_15731,N_15527);
or U15752 (N_15752,N_15654,N_15582);
nand U15753 (N_15753,N_15694,N_15512);
xnor U15754 (N_15754,N_15528,N_15635);
xnor U15755 (N_15755,N_15604,N_15547);
or U15756 (N_15756,N_15724,N_15537);
and U15757 (N_15757,N_15614,N_15513);
nor U15758 (N_15758,N_15585,N_15663);
or U15759 (N_15759,N_15649,N_15518);
nor U15760 (N_15760,N_15689,N_15639);
and U15761 (N_15761,N_15552,N_15695);
xor U15762 (N_15762,N_15590,N_15599);
or U15763 (N_15763,N_15625,N_15579);
or U15764 (N_15764,N_15530,N_15693);
and U15765 (N_15765,N_15703,N_15706);
nand U15766 (N_15766,N_15610,N_15557);
nor U15767 (N_15767,N_15745,N_15688);
nand U15768 (N_15768,N_15609,N_15619);
nor U15769 (N_15769,N_15562,N_15503);
xnor U15770 (N_15770,N_15515,N_15587);
nand U15771 (N_15771,N_15742,N_15514);
nand U15772 (N_15772,N_15636,N_15718);
and U15773 (N_15773,N_15671,N_15578);
and U15774 (N_15774,N_15738,N_15683);
nor U15775 (N_15775,N_15696,N_15642);
nand U15776 (N_15776,N_15553,N_15598);
xnor U15777 (N_15777,N_15542,N_15573);
or U15778 (N_15778,N_15640,N_15629);
nand U15779 (N_15779,N_15645,N_15680);
or U15780 (N_15780,N_15620,N_15556);
nand U15781 (N_15781,N_15707,N_15611);
xnor U15782 (N_15782,N_15712,N_15653);
nor U15783 (N_15783,N_15621,N_15540);
nand U15784 (N_15784,N_15737,N_15705);
or U15785 (N_15785,N_15743,N_15710);
xnor U15786 (N_15786,N_15728,N_15586);
xnor U15787 (N_15787,N_15520,N_15617);
and U15788 (N_15788,N_15658,N_15595);
nand U15789 (N_15789,N_15721,N_15686);
xor U15790 (N_15790,N_15637,N_15567);
and U15791 (N_15791,N_15575,N_15633);
nor U15792 (N_15792,N_15708,N_15736);
and U15793 (N_15793,N_15646,N_15559);
and U15794 (N_15794,N_15525,N_15650);
nand U15795 (N_15795,N_15676,N_15529);
nor U15796 (N_15796,N_15729,N_15667);
xor U15797 (N_15797,N_15543,N_15510);
nand U15798 (N_15798,N_15730,N_15522);
xnor U15799 (N_15799,N_15555,N_15716);
or U15800 (N_15800,N_15574,N_15698);
or U15801 (N_15801,N_15507,N_15584);
nor U15802 (N_15802,N_15500,N_15602);
or U15803 (N_15803,N_15717,N_15662);
xnor U15804 (N_15804,N_15533,N_15612);
nand U15805 (N_15805,N_15536,N_15534);
xor U15806 (N_15806,N_15613,N_15535);
nor U15807 (N_15807,N_15664,N_15506);
or U15808 (N_15808,N_15577,N_15593);
nor U15809 (N_15809,N_15732,N_15538);
or U15810 (N_15810,N_15624,N_15687);
and U15811 (N_15811,N_15704,N_15700);
nand U15812 (N_15812,N_15501,N_15748);
xor U15813 (N_15813,N_15626,N_15541);
xnor U15814 (N_15814,N_15521,N_15691);
and U15815 (N_15815,N_15692,N_15511);
nand U15816 (N_15816,N_15734,N_15623);
xnor U15817 (N_15817,N_15618,N_15516);
and U15818 (N_15818,N_15709,N_15630);
nand U15819 (N_15819,N_15678,N_15531);
and U15820 (N_15820,N_15651,N_15546);
nand U15821 (N_15821,N_15634,N_15726);
nor U15822 (N_15822,N_15713,N_15727);
and U15823 (N_15823,N_15509,N_15682);
or U15824 (N_15824,N_15545,N_15505);
and U15825 (N_15825,N_15560,N_15670);
xor U15826 (N_15826,N_15632,N_15597);
or U15827 (N_15827,N_15631,N_15656);
nor U15828 (N_15828,N_15564,N_15502);
nor U15829 (N_15829,N_15569,N_15684);
or U15830 (N_15830,N_15615,N_15583);
nand U15831 (N_15831,N_15673,N_15544);
and U15832 (N_15832,N_15566,N_15746);
nor U15833 (N_15833,N_15532,N_15568);
and U15834 (N_15834,N_15668,N_15550);
nor U15835 (N_15835,N_15596,N_15715);
and U15836 (N_15836,N_15719,N_15661);
or U15837 (N_15837,N_15608,N_15600);
and U15838 (N_15838,N_15524,N_15660);
xnor U15839 (N_15839,N_15740,N_15591);
nor U15840 (N_15840,N_15723,N_15666);
or U15841 (N_15841,N_15733,N_15665);
xor U15842 (N_15842,N_15677,N_15647);
xnor U15843 (N_15843,N_15601,N_15565);
or U15844 (N_15844,N_15669,N_15551);
or U15845 (N_15845,N_15741,N_15672);
or U15846 (N_15846,N_15549,N_15607);
xor U15847 (N_15847,N_15580,N_15643);
and U15848 (N_15848,N_15571,N_15606);
xor U15849 (N_15849,N_15526,N_15652);
or U15850 (N_15850,N_15563,N_15657);
nand U15851 (N_15851,N_15554,N_15561);
and U15852 (N_15852,N_15655,N_15628);
or U15853 (N_15853,N_15627,N_15616);
nor U15854 (N_15854,N_15605,N_15659);
or U15855 (N_15855,N_15735,N_15581);
or U15856 (N_15856,N_15539,N_15588);
xor U15857 (N_15857,N_15685,N_15648);
xnor U15858 (N_15858,N_15747,N_15570);
xnor U15859 (N_15859,N_15558,N_15504);
nand U15860 (N_15860,N_15720,N_15576);
and U15861 (N_15861,N_15702,N_15711);
nor U15862 (N_15862,N_15519,N_15622);
nor U15863 (N_15863,N_15638,N_15701);
or U15864 (N_15864,N_15517,N_15679);
xor U15865 (N_15865,N_15744,N_15681);
nand U15866 (N_15866,N_15594,N_15690);
xnor U15867 (N_15867,N_15603,N_15548);
nor U15868 (N_15868,N_15572,N_15523);
and U15869 (N_15869,N_15674,N_15641);
and U15870 (N_15870,N_15592,N_15644);
or U15871 (N_15871,N_15714,N_15739);
nor U15872 (N_15872,N_15749,N_15675);
nand U15873 (N_15873,N_15697,N_15725);
xor U15874 (N_15874,N_15699,N_15508);
nor U15875 (N_15875,N_15538,N_15530);
and U15876 (N_15876,N_15627,N_15605);
nand U15877 (N_15877,N_15568,N_15600);
nor U15878 (N_15878,N_15592,N_15503);
or U15879 (N_15879,N_15714,N_15556);
nor U15880 (N_15880,N_15635,N_15537);
and U15881 (N_15881,N_15552,N_15698);
and U15882 (N_15882,N_15647,N_15565);
nand U15883 (N_15883,N_15593,N_15651);
and U15884 (N_15884,N_15527,N_15733);
nand U15885 (N_15885,N_15594,N_15660);
or U15886 (N_15886,N_15659,N_15719);
or U15887 (N_15887,N_15618,N_15504);
nor U15888 (N_15888,N_15655,N_15580);
nor U15889 (N_15889,N_15741,N_15620);
or U15890 (N_15890,N_15684,N_15584);
xnor U15891 (N_15891,N_15728,N_15627);
nand U15892 (N_15892,N_15662,N_15517);
and U15893 (N_15893,N_15710,N_15688);
nor U15894 (N_15894,N_15736,N_15521);
xnor U15895 (N_15895,N_15747,N_15668);
and U15896 (N_15896,N_15663,N_15588);
xnor U15897 (N_15897,N_15562,N_15717);
nand U15898 (N_15898,N_15565,N_15733);
or U15899 (N_15899,N_15623,N_15708);
nand U15900 (N_15900,N_15651,N_15739);
and U15901 (N_15901,N_15574,N_15688);
nand U15902 (N_15902,N_15548,N_15684);
or U15903 (N_15903,N_15602,N_15599);
nand U15904 (N_15904,N_15667,N_15609);
or U15905 (N_15905,N_15527,N_15742);
xnor U15906 (N_15906,N_15718,N_15578);
nor U15907 (N_15907,N_15698,N_15675);
and U15908 (N_15908,N_15518,N_15720);
xor U15909 (N_15909,N_15735,N_15603);
xnor U15910 (N_15910,N_15640,N_15636);
nand U15911 (N_15911,N_15730,N_15563);
or U15912 (N_15912,N_15540,N_15642);
xor U15913 (N_15913,N_15701,N_15634);
nor U15914 (N_15914,N_15711,N_15699);
xor U15915 (N_15915,N_15671,N_15544);
and U15916 (N_15916,N_15556,N_15712);
and U15917 (N_15917,N_15635,N_15705);
xnor U15918 (N_15918,N_15566,N_15584);
nand U15919 (N_15919,N_15672,N_15564);
and U15920 (N_15920,N_15593,N_15638);
xor U15921 (N_15921,N_15687,N_15703);
nor U15922 (N_15922,N_15712,N_15747);
and U15923 (N_15923,N_15542,N_15525);
xor U15924 (N_15924,N_15520,N_15593);
nand U15925 (N_15925,N_15636,N_15650);
and U15926 (N_15926,N_15509,N_15542);
and U15927 (N_15927,N_15639,N_15601);
nor U15928 (N_15928,N_15630,N_15555);
or U15929 (N_15929,N_15626,N_15616);
or U15930 (N_15930,N_15637,N_15546);
nor U15931 (N_15931,N_15635,N_15669);
xnor U15932 (N_15932,N_15710,N_15606);
and U15933 (N_15933,N_15637,N_15718);
and U15934 (N_15934,N_15680,N_15506);
nor U15935 (N_15935,N_15533,N_15583);
nor U15936 (N_15936,N_15571,N_15729);
nand U15937 (N_15937,N_15616,N_15663);
or U15938 (N_15938,N_15655,N_15687);
or U15939 (N_15939,N_15608,N_15689);
and U15940 (N_15940,N_15697,N_15500);
nand U15941 (N_15941,N_15595,N_15532);
and U15942 (N_15942,N_15728,N_15666);
nor U15943 (N_15943,N_15701,N_15686);
and U15944 (N_15944,N_15713,N_15664);
nand U15945 (N_15945,N_15651,N_15635);
nand U15946 (N_15946,N_15663,N_15577);
or U15947 (N_15947,N_15642,N_15720);
nor U15948 (N_15948,N_15502,N_15665);
nor U15949 (N_15949,N_15690,N_15532);
nand U15950 (N_15950,N_15523,N_15633);
or U15951 (N_15951,N_15711,N_15674);
or U15952 (N_15952,N_15534,N_15682);
and U15953 (N_15953,N_15570,N_15739);
and U15954 (N_15954,N_15553,N_15536);
or U15955 (N_15955,N_15534,N_15607);
nand U15956 (N_15956,N_15730,N_15515);
nor U15957 (N_15957,N_15679,N_15584);
and U15958 (N_15958,N_15562,N_15687);
nor U15959 (N_15959,N_15502,N_15546);
nor U15960 (N_15960,N_15533,N_15509);
or U15961 (N_15961,N_15577,N_15561);
and U15962 (N_15962,N_15534,N_15586);
xor U15963 (N_15963,N_15642,N_15505);
and U15964 (N_15964,N_15523,N_15629);
or U15965 (N_15965,N_15585,N_15504);
nor U15966 (N_15966,N_15587,N_15567);
nand U15967 (N_15967,N_15551,N_15714);
xor U15968 (N_15968,N_15540,N_15512);
nor U15969 (N_15969,N_15563,N_15642);
nor U15970 (N_15970,N_15628,N_15642);
xnor U15971 (N_15971,N_15598,N_15708);
and U15972 (N_15972,N_15632,N_15508);
xnor U15973 (N_15973,N_15512,N_15501);
and U15974 (N_15974,N_15555,N_15556);
or U15975 (N_15975,N_15547,N_15577);
and U15976 (N_15976,N_15658,N_15664);
and U15977 (N_15977,N_15661,N_15687);
nand U15978 (N_15978,N_15533,N_15646);
and U15979 (N_15979,N_15724,N_15602);
nor U15980 (N_15980,N_15657,N_15524);
nand U15981 (N_15981,N_15661,N_15578);
nor U15982 (N_15982,N_15669,N_15503);
and U15983 (N_15983,N_15722,N_15650);
nor U15984 (N_15984,N_15625,N_15593);
xor U15985 (N_15985,N_15501,N_15665);
or U15986 (N_15986,N_15585,N_15575);
nand U15987 (N_15987,N_15672,N_15718);
nand U15988 (N_15988,N_15591,N_15646);
or U15989 (N_15989,N_15630,N_15701);
nand U15990 (N_15990,N_15561,N_15725);
nand U15991 (N_15991,N_15598,N_15677);
nor U15992 (N_15992,N_15549,N_15590);
xnor U15993 (N_15993,N_15605,N_15721);
or U15994 (N_15994,N_15606,N_15629);
xnor U15995 (N_15995,N_15625,N_15587);
and U15996 (N_15996,N_15588,N_15535);
nor U15997 (N_15997,N_15558,N_15548);
xnor U15998 (N_15998,N_15725,N_15596);
and U15999 (N_15999,N_15629,N_15512);
nand U16000 (N_16000,N_15880,N_15909);
nand U16001 (N_16001,N_15923,N_15910);
nand U16002 (N_16002,N_15788,N_15834);
and U16003 (N_16003,N_15874,N_15878);
nand U16004 (N_16004,N_15875,N_15825);
nand U16005 (N_16005,N_15873,N_15978);
or U16006 (N_16006,N_15828,N_15848);
xor U16007 (N_16007,N_15912,N_15781);
nor U16008 (N_16008,N_15915,N_15937);
xor U16009 (N_16009,N_15870,N_15974);
xor U16010 (N_16010,N_15907,N_15888);
nand U16011 (N_16011,N_15751,N_15760);
nand U16012 (N_16012,N_15903,N_15997);
nor U16013 (N_16013,N_15976,N_15829);
or U16014 (N_16014,N_15864,N_15756);
and U16015 (N_16015,N_15835,N_15911);
and U16016 (N_16016,N_15750,N_15922);
nor U16017 (N_16017,N_15883,N_15995);
and U16018 (N_16018,N_15948,N_15863);
or U16019 (N_16019,N_15953,N_15851);
nand U16020 (N_16020,N_15803,N_15979);
and U16021 (N_16021,N_15782,N_15905);
and U16022 (N_16022,N_15849,N_15811);
or U16023 (N_16023,N_15975,N_15898);
and U16024 (N_16024,N_15936,N_15934);
nand U16025 (N_16025,N_15799,N_15792);
nor U16026 (N_16026,N_15805,N_15806);
nand U16027 (N_16027,N_15964,N_15776);
nor U16028 (N_16028,N_15941,N_15988);
nand U16029 (N_16029,N_15869,N_15839);
xnor U16030 (N_16030,N_15761,N_15819);
nor U16031 (N_16031,N_15946,N_15897);
nor U16032 (N_16032,N_15758,N_15753);
xnor U16033 (N_16033,N_15774,N_15815);
and U16034 (N_16034,N_15824,N_15957);
nand U16035 (N_16035,N_15752,N_15924);
nand U16036 (N_16036,N_15812,N_15862);
nand U16037 (N_16037,N_15963,N_15969);
and U16038 (N_16038,N_15780,N_15841);
xor U16039 (N_16039,N_15847,N_15939);
and U16040 (N_16040,N_15944,N_15858);
xor U16041 (N_16041,N_15808,N_15857);
nand U16042 (N_16042,N_15986,N_15861);
xor U16043 (N_16043,N_15790,N_15893);
and U16044 (N_16044,N_15859,N_15767);
nor U16045 (N_16045,N_15884,N_15970);
or U16046 (N_16046,N_15795,N_15867);
nand U16047 (N_16047,N_15956,N_15899);
or U16048 (N_16048,N_15930,N_15991);
nor U16049 (N_16049,N_15967,N_15990);
and U16050 (N_16050,N_15913,N_15791);
xnor U16051 (N_16051,N_15932,N_15826);
xor U16052 (N_16052,N_15968,N_15830);
or U16053 (N_16053,N_15935,N_15852);
and U16054 (N_16054,N_15793,N_15856);
xor U16055 (N_16055,N_15892,N_15854);
and U16056 (N_16056,N_15928,N_15777);
and U16057 (N_16057,N_15794,N_15985);
nor U16058 (N_16058,N_15817,N_15813);
nor U16059 (N_16059,N_15973,N_15980);
nor U16060 (N_16060,N_15994,N_15796);
nand U16061 (N_16061,N_15823,N_15821);
or U16062 (N_16062,N_15797,N_15904);
or U16063 (N_16063,N_15989,N_15925);
xor U16064 (N_16064,N_15787,N_15801);
or U16065 (N_16065,N_15771,N_15755);
xnor U16066 (N_16066,N_15949,N_15872);
xor U16067 (N_16067,N_15929,N_15802);
xnor U16068 (N_16068,N_15977,N_15942);
and U16069 (N_16069,N_15814,N_15959);
xor U16070 (N_16070,N_15764,N_15759);
nor U16071 (N_16071,N_15918,N_15882);
and U16072 (N_16072,N_15783,N_15837);
or U16073 (N_16073,N_15868,N_15916);
and U16074 (N_16074,N_15810,N_15938);
nor U16075 (N_16075,N_15855,N_15769);
xnor U16076 (N_16076,N_15807,N_15853);
nand U16077 (N_16077,N_15955,N_15785);
nor U16078 (N_16078,N_15876,N_15984);
nand U16079 (N_16079,N_15784,N_15779);
and U16080 (N_16080,N_15754,N_15840);
nand U16081 (N_16081,N_15838,N_15998);
nor U16082 (N_16082,N_15800,N_15900);
xor U16083 (N_16083,N_15827,N_15762);
nand U16084 (N_16084,N_15845,N_15917);
and U16085 (N_16085,N_15886,N_15770);
xnor U16086 (N_16086,N_15971,N_15877);
and U16087 (N_16087,N_15972,N_15940);
nand U16088 (N_16088,N_15999,N_15947);
xor U16089 (N_16089,N_15765,N_15775);
nor U16090 (N_16090,N_15921,N_15996);
or U16091 (N_16091,N_15901,N_15960);
or U16092 (N_16092,N_15871,N_15890);
xnor U16093 (N_16093,N_15983,N_15843);
xnor U16094 (N_16094,N_15832,N_15958);
xnor U16095 (N_16095,N_15836,N_15773);
or U16096 (N_16096,N_15914,N_15902);
nor U16097 (N_16097,N_15927,N_15951);
xor U16098 (N_16098,N_15860,N_15831);
xor U16099 (N_16099,N_15961,N_15931);
and U16100 (N_16100,N_15763,N_15757);
and U16101 (N_16101,N_15865,N_15798);
nor U16102 (N_16102,N_15950,N_15866);
nor U16103 (N_16103,N_15850,N_15786);
nand U16104 (N_16104,N_15818,N_15822);
nand U16105 (N_16105,N_15966,N_15993);
xnor U16106 (N_16106,N_15809,N_15842);
nor U16107 (N_16107,N_15926,N_15804);
or U16108 (N_16108,N_15987,N_15820);
nand U16109 (N_16109,N_15896,N_15943);
and U16110 (N_16110,N_15881,N_15945);
or U16111 (N_16111,N_15920,N_15992);
and U16112 (N_16112,N_15908,N_15965);
nand U16113 (N_16113,N_15919,N_15766);
xor U16114 (N_16114,N_15887,N_15962);
xor U16115 (N_16115,N_15981,N_15894);
and U16116 (N_16116,N_15889,N_15952);
nor U16117 (N_16117,N_15906,N_15879);
nand U16118 (N_16118,N_15768,N_15772);
nand U16119 (N_16119,N_15833,N_15982);
nor U16120 (N_16120,N_15885,N_15933);
and U16121 (N_16121,N_15816,N_15895);
xnor U16122 (N_16122,N_15778,N_15844);
xor U16123 (N_16123,N_15846,N_15891);
or U16124 (N_16124,N_15954,N_15789);
and U16125 (N_16125,N_15923,N_15897);
nor U16126 (N_16126,N_15753,N_15914);
or U16127 (N_16127,N_15835,N_15943);
nor U16128 (N_16128,N_15925,N_15759);
nor U16129 (N_16129,N_15850,N_15757);
xor U16130 (N_16130,N_15999,N_15942);
and U16131 (N_16131,N_15959,N_15812);
or U16132 (N_16132,N_15939,N_15998);
nand U16133 (N_16133,N_15817,N_15873);
nand U16134 (N_16134,N_15758,N_15763);
nand U16135 (N_16135,N_15812,N_15820);
nand U16136 (N_16136,N_15800,N_15920);
nor U16137 (N_16137,N_15873,N_15761);
nand U16138 (N_16138,N_15978,N_15874);
and U16139 (N_16139,N_15834,N_15854);
nand U16140 (N_16140,N_15984,N_15859);
nand U16141 (N_16141,N_15855,N_15875);
nor U16142 (N_16142,N_15888,N_15945);
or U16143 (N_16143,N_15816,N_15792);
xor U16144 (N_16144,N_15854,N_15858);
nor U16145 (N_16145,N_15760,N_15887);
or U16146 (N_16146,N_15888,N_15857);
nor U16147 (N_16147,N_15888,N_15791);
xor U16148 (N_16148,N_15977,N_15757);
nand U16149 (N_16149,N_15774,N_15752);
nor U16150 (N_16150,N_15788,N_15874);
nor U16151 (N_16151,N_15950,N_15924);
and U16152 (N_16152,N_15967,N_15842);
or U16153 (N_16153,N_15950,N_15974);
or U16154 (N_16154,N_15864,N_15763);
or U16155 (N_16155,N_15946,N_15799);
or U16156 (N_16156,N_15834,N_15990);
and U16157 (N_16157,N_15798,N_15873);
xnor U16158 (N_16158,N_15885,N_15957);
or U16159 (N_16159,N_15906,N_15978);
xnor U16160 (N_16160,N_15899,N_15759);
nand U16161 (N_16161,N_15758,N_15793);
xor U16162 (N_16162,N_15754,N_15941);
and U16163 (N_16163,N_15961,N_15786);
and U16164 (N_16164,N_15901,N_15850);
and U16165 (N_16165,N_15941,N_15822);
and U16166 (N_16166,N_15791,N_15895);
and U16167 (N_16167,N_15847,N_15894);
nand U16168 (N_16168,N_15806,N_15775);
xnor U16169 (N_16169,N_15993,N_15777);
nand U16170 (N_16170,N_15886,N_15945);
nand U16171 (N_16171,N_15928,N_15981);
xor U16172 (N_16172,N_15896,N_15833);
nor U16173 (N_16173,N_15915,N_15953);
xor U16174 (N_16174,N_15817,N_15838);
and U16175 (N_16175,N_15906,N_15775);
or U16176 (N_16176,N_15912,N_15940);
nor U16177 (N_16177,N_15978,N_15907);
and U16178 (N_16178,N_15939,N_15853);
nor U16179 (N_16179,N_15871,N_15984);
nor U16180 (N_16180,N_15867,N_15785);
or U16181 (N_16181,N_15991,N_15885);
or U16182 (N_16182,N_15798,N_15852);
xnor U16183 (N_16183,N_15949,N_15757);
xnor U16184 (N_16184,N_15987,N_15908);
nand U16185 (N_16185,N_15821,N_15897);
nand U16186 (N_16186,N_15879,N_15851);
nor U16187 (N_16187,N_15981,N_15857);
or U16188 (N_16188,N_15784,N_15939);
xnor U16189 (N_16189,N_15778,N_15907);
or U16190 (N_16190,N_15983,N_15990);
xnor U16191 (N_16191,N_15832,N_15831);
xnor U16192 (N_16192,N_15986,N_15844);
or U16193 (N_16193,N_15864,N_15907);
nand U16194 (N_16194,N_15768,N_15978);
nor U16195 (N_16195,N_15937,N_15769);
and U16196 (N_16196,N_15920,N_15778);
xnor U16197 (N_16197,N_15786,N_15809);
nor U16198 (N_16198,N_15975,N_15885);
or U16199 (N_16199,N_15935,N_15916);
nand U16200 (N_16200,N_15770,N_15981);
nand U16201 (N_16201,N_15957,N_15773);
nor U16202 (N_16202,N_15927,N_15990);
nand U16203 (N_16203,N_15832,N_15826);
xnor U16204 (N_16204,N_15982,N_15821);
or U16205 (N_16205,N_15979,N_15766);
xnor U16206 (N_16206,N_15804,N_15953);
or U16207 (N_16207,N_15794,N_15932);
or U16208 (N_16208,N_15794,N_15891);
nor U16209 (N_16209,N_15777,N_15779);
nor U16210 (N_16210,N_15948,N_15919);
and U16211 (N_16211,N_15827,N_15826);
and U16212 (N_16212,N_15864,N_15929);
nor U16213 (N_16213,N_15787,N_15926);
xor U16214 (N_16214,N_15931,N_15912);
xor U16215 (N_16215,N_15904,N_15968);
or U16216 (N_16216,N_15857,N_15778);
or U16217 (N_16217,N_15988,N_15806);
nor U16218 (N_16218,N_15878,N_15785);
or U16219 (N_16219,N_15810,N_15818);
nand U16220 (N_16220,N_15825,N_15813);
and U16221 (N_16221,N_15902,N_15835);
nand U16222 (N_16222,N_15846,N_15755);
and U16223 (N_16223,N_15974,N_15827);
or U16224 (N_16224,N_15770,N_15764);
nand U16225 (N_16225,N_15953,N_15972);
or U16226 (N_16226,N_15856,N_15917);
or U16227 (N_16227,N_15907,N_15895);
or U16228 (N_16228,N_15926,N_15957);
or U16229 (N_16229,N_15901,N_15788);
or U16230 (N_16230,N_15939,N_15967);
nor U16231 (N_16231,N_15787,N_15902);
or U16232 (N_16232,N_15816,N_15929);
or U16233 (N_16233,N_15752,N_15867);
and U16234 (N_16234,N_15777,N_15896);
nor U16235 (N_16235,N_15857,N_15982);
nand U16236 (N_16236,N_15836,N_15829);
nor U16237 (N_16237,N_15835,N_15975);
xor U16238 (N_16238,N_15833,N_15752);
nor U16239 (N_16239,N_15835,N_15891);
nor U16240 (N_16240,N_15832,N_15808);
or U16241 (N_16241,N_15855,N_15983);
or U16242 (N_16242,N_15967,N_15980);
and U16243 (N_16243,N_15770,N_15906);
nor U16244 (N_16244,N_15811,N_15776);
xnor U16245 (N_16245,N_15991,N_15918);
nor U16246 (N_16246,N_15847,N_15775);
xor U16247 (N_16247,N_15827,N_15979);
xor U16248 (N_16248,N_15827,N_15878);
and U16249 (N_16249,N_15769,N_15872);
nor U16250 (N_16250,N_16133,N_16230);
or U16251 (N_16251,N_16228,N_16086);
and U16252 (N_16252,N_16156,N_16095);
nand U16253 (N_16253,N_16082,N_16234);
or U16254 (N_16254,N_16080,N_16209);
and U16255 (N_16255,N_16180,N_16088);
and U16256 (N_16256,N_16140,N_16241);
nor U16257 (N_16257,N_16046,N_16168);
nor U16258 (N_16258,N_16019,N_16031);
xnor U16259 (N_16259,N_16004,N_16008);
nand U16260 (N_16260,N_16183,N_16128);
nand U16261 (N_16261,N_16021,N_16174);
or U16262 (N_16262,N_16016,N_16189);
xor U16263 (N_16263,N_16101,N_16130);
xor U16264 (N_16264,N_16076,N_16055);
and U16265 (N_16265,N_16247,N_16167);
nand U16266 (N_16266,N_16237,N_16112);
or U16267 (N_16267,N_16041,N_16062);
nand U16268 (N_16268,N_16065,N_16106);
xnor U16269 (N_16269,N_16018,N_16212);
nor U16270 (N_16270,N_16192,N_16064);
xnor U16271 (N_16271,N_16181,N_16075);
nor U16272 (N_16272,N_16150,N_16207);
and U16273 (N_16273,N_16052,N_16114);
and U16274 (N_16274,N_16022,N_16147);
and U16275 (N_16275,N_16170,N_16023);
and U16276 (N_16276,N_16048,N_16227);
or U16277 (N_16277,N_16006,N_16161);
xor U16278 (N_16278,N_16120,N_16193);
nand U16279 (N_16279,N_16217,N_16104);
nor U16280 (N_16280,N_16175,N_16215);
nand U16281 (N_16281,N_16225,N_16173);
xnor U16282 (N_16282,N_16159,N_16162);
or U16283 (N_16283,N_16202,N_16091);
and U16284 (N_16284,N_16049,N_16115);
xor U16285 (N_16285,N_16110,N_16142);
or U16286 (N_16286,N_16063,N_16097);
or U16287 (N_16287,N_16210,N_16148);
xor U16288 (N_16288,N_16200,N_16094);
nor U16289 (N_16289,N_16187,N_16153);
or U16290 (N_16290,N_16007,N_16099);
xnor U16291 (N_16291,N_16155,N_16236);
xnor U16292 (N_16292,N_16047,N_16003);
nor U16293 (N_16293,N_16229,N_16078);
xor U16294 (N_16294,N_16176,N_16085);
and U16295 (N_16295,N_16030,N_16033);
nor U16296 (N_16296,N_16157,N_16073);
xor U16297 (N_16297,N_16043,N_16034);
and U16298 (N_16298,N_16098,N_16137);
nand U16299 (N_16299,N_16131,N_16151);
nor U16300 (N_16300,N_16190,N_16163);
and U16301 (N_16301,N_16077,N_16188);
nor U16302 (N_16302,N_16223,N_16239);
or U16303 (N_16303,N_16214,N_16182);
and U16304 (N_16304,N_16244,N_16070);
nor U16305 (N_16305,N_16017,N_16154);
xnor U16306 (N_16306,N_16011,N_16152);
xor U16307 (N_16307,N_16179,N_16132);
and U16308 (N_16308,N_16012,N_16037);
or U16309 (N_16309,N_16221,N_16029);
xnor U16310 (N_16310,N_16222,N_16040);
xor U16311 (N_16311,N_16145,N_16013);
and U16312 (N_16312,N_16197,N_16143);
or U16313 (N_16313,N_16172,N_16015);
and U16314 (N_16314,N_16010,N_16194);
nor U16315 (N_16315,N_16204,N_16044);
nand U16316 (N_16316,N_16146,N_16224);
or U16317 (N_16317,N_16090,N_16233);
and U16318 (N_16318,N_16054,N_16032);
nor U16319 (N_16319,N_16035,N_16125);
and U16320 (N_16320,N_16108,N_16220);
nor U16321 (N_16321,N_16165,N_16127);
or U16322 (N_16322,N_16045,N_16124);
or U16323 (N_16323,N_16083,N_16169);
nand U16324 (N_16324,N_16240,N_16050);
nor U16325 (N_16325,N_16235,N_16134);
and U16326 (N_16326,N_16116,N_16103);
and U16327 (N_16327,N_16005,N_16122);
nand U16328 (N_16328,N_16129,N_16026);
and U16329 (N_16329,N_16100,N_16199);
or U16330 (N_16330,N_16109,N_16211);
xnor U16331 (N_16331,N_16001,N_16071);
xor U16332 (N_16332,N_16249,N_16246);
or U16333 (N_16333,N_16042,N_16139);
nor U16334 (N_16334,N_16178,N_16198);
or U16335 (N_16335,N_16102,N_16231);
xor U16336 (N_16336,N_16057,N_16081);
nor U16337 (N_16337,N_16123,N_16160);
and U16338 (N_16338,N_16196,N_16009);
and U16339 (N_16339,N_16206,N_16141);
nand U16340 (N_16340,N_16093,N_16068);
nand U16341 (N_16341,N_16158,N_16144);
nand U16342 (N_16342,N_16092,N_16089);
and U16343 (N_16343,N_16038,N_16226);
nand U16344 (N_16344,N_16164,N_16096);
and U16345 (N_16345,N_16014,N_16051);
nand U16346 (N_16346,N_16171,N_16205);
or U16347 (N_16347,N_16105,N_16216);
or U16348 (N_16348,N_16248,N_16061);
xnor U16349 (N_16349,N_16053,N_16079);
nand U16350 (N_16350,N_16219,N_16185);
or U16351 (N_16351,N_16195,N_16232);
xor U16352 (N_16352,N_16119,N_16191);
nor U16353 (N_16353,N_16136,N_16074);
nor U16354 (N_16354,N_16060,N_16177);
nor U16355 (N_16355,N_16208,N_16027);
or U16356 (N_16356,N_16126,N_16121);
xor U16357 (N_16357,N_16201,N_16111);
and U16358 (N_16358,N_16036,N_16072);
or U16359 (N_16359,N_16118,N_16058);
and U16360 (N_16360,N_16242,N_16213);
or U16361 (N_16361,N_16166,N_16084);
or U16362 (N_16362,N_16039,N_16243);
nor U16363 (N_16363,N_16067,N_16028);
nor U16364 (N_16364,N_16069,N_16087);
and U16365 (N_16365,N_16113,N_16024);
and U16366 (N_16366,N_16056,N_16135);
and U16367 (N_16367,N_16186,N_16000);
and U16368 (N_16368,N_16066,N_16025);
nand U16369 (N_16369,N_16149,N_16218);
or U16370 (N_16370,N_16138,N_16117);
nand U16371 (N_16371,N_16184,N_16002);
and U16372 (N_16372,N_16059,N_16020);
nor U16373 (N_16373,N_16107,N_16203);
xor U16374 (N_16374,N_16245,N_16238);
nand U16375 (N_16375,N_16221,N_16165);
xnor U16376 (N_16376,N_16154,N_16108);
nor U16377 (N_16377,N_16130,N_16038);
nand U16378 (N_16378,N_16210,N_16035);
xor U16379 (N_16379,N_16014,N_16015);
or U16380 (N_16380,N_16176,N_16012);
nor U16381 (N_16381,N_16093,N_16063);
xor U16382 (N_16382,N_16206,N_16216);
xnor U16383 (N_16383,N_16070,N_16126);
and U16384 (N_16384,N_16099,N_16179);
and U16385 (N_16385,N_16226,N_16026);
nand U16386 (N_16386,N_16062,N_16129);
xor U16387 (N_16387,N_16003,N_16107);
nand U16388 (N_16388,N_16060,N_16082);
nor U16389 (N_16389,N_16089,N_16040);
or U16390 (N_16390,N_16094,N_16021);
and U16391 (N_16391,N_16083,N_16017);
nor U16392 (N_16392,N_16011,N_16089);
xor U16393 (N_16393,N_16173,N_16027);
xnor U16394 (N_16394,N_16047,N_16087);
xor U16395 (N_16395,N_16002,N_16159);
and U16396 (N_16396,N_16111,N_16232);
nand U16397 (N_16397,N_16227,N_16091);
and U16398 (N_16398,N_16102,N_16066);
xor U16399 (N_16399,N_16106,N_16030);
nor U16400 (N_16400,N_16194,N_16110);
and U16401 (N_16401,N_16014,N_16074);
nand U16402 (N_16402,N_16084,N_16168);
or U16403 (N_16403,N_16093,N_16010);
nand U16404 (N_16404,N_16062,N_16142);
xor U16405 (N_16405,N_16225,N_16157);
xnor U16406 (N_16406,N_16193,N_16035);
nor U16407 (N_16407,N_16173,N_16224);
nand U16408 (N_16408,N_16229,N_16168);
or U16409 (N_16409,N_16190,N_16080);
nor U16410 (N_16410,N_16239,N_16129);
or U16411 (N_16411,N_16055,N_16001);
xnor U16412 (N_16412,N_16007,N_16202);
nor U16413 (N_16413,N_16152,N_16060);
nand U16414 (N_16414,N_16055,N_16212);
or U16415 (N_16415,N_16120,N_16051);
nor U16416 (N_16416,N_16132,N_16047);
xnor U16417 (N_16417,N_16086,N_16233);
xor U16418 (N_16418,N_16050,N_16221);
nor U16419 (N_16419,N_16223,N_16126);
or U16420 (N_16420,N_16077,N_16110);
or U16421 (N_16421,N_16111,N_16118);
and U16422 (N_16422,N_16044,N_16011);
or U16423 (N_16423,N_16058,N_16208);
xnor U16424 (N_16424,N_16098,N_16051);
or U16425 (N_16425,N_16230,N_16035);
nand U16426 (N_16426,N_16099,N_16063);
and U16427 (N_16427,N_16149,N_16029);
nand U16428 (N_16428,N_16026,N_16091);
and U16429 (N_16429,N_16171,N_16075);
nand U16430 (N_16430,N_16088,N_16225);
and U16431 (N_16431,N_16010,N_16185);
and U16432 (N_16432,N_16118,N_16232);
or U16433 (N_16433,N_16094,N_16107);
xnor U16434 (N_16434,N_16038,N_16119);
and U16435 (N_16435,N_16080,N_16018);
nor U16436 (N_16436,N_16121,N_16123);
xnor U16437 (N_16437,N_16072,N_16103);
or U16438 (N_16438,N_16048,N_16122);
or U16439 (N_16439,N_16010,N_16175);
xor U16440 (N_16440,N_16153,N_16031);
xor U16441 (N_16441,N_16210,N_16106);
nand U16442 (N_16442,N_16140,N_16234);
nand U16443 (N_16443,N_16112,N_16216);
nand U16444 (N_16444,N_16161,N_16205);
and U16445 (N_16445,N_16032,N_16226);
nand U16446 (N_16446,N_16096,N_16098);
and U16447 (N_16447,N_16196,N_16002);
xor U16448 (N_16448,N_16194,N_16052);
nor U16449 (N_16449,N_16238,N_16171);
xnor U16450 (N_16450,N_16060,N_16043);
xnor U16451 (N_16451,N_16139,N_16201);
and U16452 (N_16452,N_16213,N_16161);
nor U16453 (N_16453,N_16225,N_16037);
xor U16454 (N_16454,N_16046,N_16188);
and U16455 (N_16455,N_16078,N_16082);
and U16456 (N_16456,N_16183,N_16228);
xor U16457 (N_16457,N_16183,N_16155);
nand U16458 (N_16458,N_16031,N_16160);
or U16459 (N_16459,N_16095,N_16161);
or U16460 (N_16460,N_16029,N_16062);
and U16461 (N_16461,N_16056,N_16036);
or U16462 (N_16462,N_16228,N_16189);
and U16463 (N_16463,N_16088,N_16178);
nand U16464 (N_16464,N_16158,N_16037);
or U16465 (N_16465,N_16223,N_16066);
and U16466 (N_16466,N_16076,N_16037);
or U16467 (N_16467,N_16166,N_16177);
nor U16468 (N_16468,N_16136,N_16168);
nand U16469 (N_16469,N_16178,N_16122);
or U16470 (N_16470,N_16104,N_16097);
nor U16471 (N_16471,N_16044,N_16024);
or U16472 (N_16472,N_16014,N_16064);
and U16473 (N_16473,N_16153,N_16122);
xor U16474 (N_16474,N_16058,N_16205);
and U16475 (N_16475,N_16228,N_16216);
nor U16476 (N_16476,N_16059,N_16014);
nor U16477 (N_16477,N_16083,N_16036);
xor U16478 (N_16478,N_16071,N_16233);
nand U16479 (N_16479,N_16013,N_16108);
and U16480 (N_16480,N_16114,N_16177);
nand U16481 (N_16481,N_16238,N_16205);
xnor U16482 (N_16482,N_16239,N_16073);
xnor U16483 (N_16483,N_16007,N_16080);
and U16484 (N_16484,N_16054,N_16215);
and U16485 (N_16485,N_16176,N_16088);
xor U16486 (N_16486,N_16088,N_16222);
xor U16487 (N_16487,N_16099,N_16011);
and U16488 (N_16488,N_16046,N_16078);
nand U16489 (N_16489,N_16095,N_16107);
and U16490 (N_16490,N_16115,N_16081);
and U16491 (N_16491,N_16066,N_16117);
or U16492 (N_16492,N_16224,N_16119);
nand U16493 (N_16493,N_16119,N_16172);
xnor U16494 (N_16494,N_16035,N_16178);
nor U16495 (N_16495,N_16202,N_16205);
nor U16496 (N_16496,N_16115,N_16052);
or U16497 (N_16497,N_16077,N_16098);
and U16498 (N_16498,N_16010,N_16229);
nand U16499 (N_16499,N_16082,N_16147);
nand U16500 (N_16500,N_16481,N_16342);
and U16501 (N_16501,N_16487,N_16309);
and U16502 (N_16502,N_16498,N_16379);
xnor U16503 (N_16503,N_16336,N_16307);
nand U16504 (N_16504,N_16256,N_16293);
xnor U16505 (N_16505,N_16434,N_16362);
nor U16506 (N_16506,N_16350,N_16308);
nor U16507 (N_16507,N_16426,N_16359);
xnor U16508 (N_16508,N_16430,N_16402);
nand U16509 (N_16509,N_16278,N_16329);
nand U16510 (N_16510,N_16253,N_16288);
xnor U16511 (N_16511,N_16279,N_16399);
and U16512 (N_16512,N_16429,N_16346);
and U16513 (N_16513,N_16281,N_16393);
and U16514 (N_16514,N_16305,N_16444);
nand U16515 (N_16515,N_16284,N_16250);
nand U16516 (N_16516,N_16265,N_16427);
nor U16517 (N_16517,N_16365,N_16277);
and U16518 (N_16518,N_16264,N_16479);
and U16519 (N_16519,N_16302,N_16450);
nand U16520 (N_16520,N_16344,N_16400);
and U16521 (N_16521,N_16283,N_16392);
and U16522 (N_16522,N_16340,N_16316);
nor U16523 (N_16523,N_16396,N_16339);
xor U16524 (N_16524,N_16436,N_16404);
and U16525 (N_16525,N_16272,N_16303);
xor U16526 (N_16526,N_16424,N_16422);
and U16527 (N_16527,N_16294,N_16482);
or U16528 (N_16528,N_16258,N_16297);
and U16529 (N_16529,N_16291,N_16317);
or U16530 (N_16530,N_16347,N_16273);
xor U16531 (N_16531,N_16492,N_16374);
nor U16532 (N_16532,N_16383,N_16420);
xor U16533 (N_16533,N_16386,N_16413);
xnor U16534 (N_16534,N_16301,N_16416);
or U16535 (N_16535,N_16442,N_16299);
or U16536 (N_16536,N_16384,N_16300);
nor U16537 (N_16537,N_16370,N_16364);
or U16538 (N_16538,N_16381,N_16472);
and U16539 (N_16539,N_16356,N_16345);
xnor U16540 (N_16540,N_16490,N_16457);
nor U16541 (N_16541,N_16321,N_16326);
nor U16542 (N_16542,N_16469,N_16263);
xor U16543 (N_16543,N_16330,N_16282);
nand U16544 (N_16544,N_16323,N_16441);
or U16545 (N_16545,N_16463,N_16285);
or U16546 (N_16546,N_16437,N_16335);
nand U16547 (N_16547,N_16403,N_16325);
nor U16548 (N_16548,N_16451,N_16377);
xor U16549 (N_16549,N_16439,N_16331);
nand U16550 (N_16550,N_16435,N_16408);
and U16551 (N_16551,N_16320,N_16310);
nor U16552 (N_16552,N_16462,N_16324);
nand U16553 (N_16553,N_16360,N_16373);
xor U16554 (N_16554,N_16447,N_16296);
and U16555 (N_16555,N_16304,N_16410);
xor U16556 (N_16556,N_16460,N_16419);
or U16557 (N_16557,N_16328,N_16270);
nand U16558 (N_16558,N_16261,N_16476);
nand U16559 (N_16559,N_16448,N_16488);
xnor U16560 (N_16560,N_16438,N_16269);
nand U16561 (N_16561,N_16337,N_16355);
xor U16562 (N_16562,N_16414,N_16327);
nor U16563 (N_16563,N_16489,N_16260);
and U16564 (N_16564,N_16313,N_16391);
and U16565 (N_16565,N_16333,N_16431);
nand U16566 (N_16566,N_16405,N_16372);
nor U16567 (N_16567,N_16385,N_16389);
nor U16568 (N_16568,N_16470,N_16499);
and U16569 (N_16569,N_16415,N_16406);
or U16570 (N_16570,N_16494,N_16466);
and U16571 (N_16571,N_16371,N_16390);
xor U16572 (N_16572,N_16478,N_16252);
nor U16573 (N_16573,N_16351,N_16456);
xnor U16574 (N_16574,N_16358,N_16380);
xnor U16575 (N_16575,N_16375,N_16443);
and U16576 (N_16576,N_16352,N_16266);
nand U16577 (N_16577,N_16480,N_16401);
and U16578 (N_16578,N_16486,N_16425);
nor U16579 (N_16579,N_16421,N_16338);
nor U16580 (N_16580,N_16306,N_16395);
and U16581 (N_16581,N_16254,N_16312);
xnor U16582 (N_16582,N_16423,N_16311);
xor U16583 (N_16583,N_16394,N_16290);
and U16584 (N_16584,N_16268,N_16295);
xnor U16585 (N_16585,N_16286,N_16409);
or U16586 (N_16586,N_16289,N_16428);
nand U16587 (N_16587,N_16348,N_16315);
and U16588 (N_16588,N_16349,N_16475);
xor U16589 (N_16589,N_16334,N_16274);
and U16590 (N_16590,N_16411,N_16267);
xnor U16591 (N_16591,N_16262,N_16407);
nand U16592 (N_16592,N_16388,N_16397);
nor U16593 (N_16593,N_16433,N_16343);
nand U16594 (N_16594,N_16341,N_16257);
xor U16595 (N_16595,N_16467,N_16412);
and U16596 (N_16596,N_16471,N_16477);
xnor U16597 (N_16597,N_16473,N_16496);
xor U16598 (N_16598,N_16276,N_16318);
or U16599 (N_16599,N_16366,N_16271);
or U16600 (N_16600,N_16275,N_16298);
or U16601 (N_16601,N_16465,N_16495);
xnor U16602 (N_16602,N_16418,N_16332);
xor U16603 (N_16603,N_16376,N_16361);
nor U16604 (N_16604,N_16417,N_16251);
and U16605 (N_16605,N_16453,N_16353);
or U16606 (N_16606,N_16483,N_16432);
nand U16607 (N_16607,N_16452,N_16369);
or U16608 (N_16608,N_16398,N_16485);
nand U16609 (N_16609,N_16292,N_16449);
nand U16610 (N_16610,N_16445,N_16491);
or U16611 (N_16611,N_16255,N_16259);
nor U16612 (N_16612,N_16357,N_16319);
nor U16613 (N_16613,N_16314,N_16354);
and U16614 (N_16614,N_16368,N_16387);
nand U16615 (N_16615,N_16363,N_16459);
nand U16616 (N_16616,N_16322,N_16280);
nor U16617 (N_16617,N_16382,N_16484);
nand U16618 (N_16618,N_16287,N_16468);
nand U16619 (N_16619,N_16367,N_16464);
or U16620 (N_16620,N_16497,N_16446);
xor U16621 (N_16621,N_16493,N_16454);
and U16622 (N_16622,N_16474,N_16461);
and U16623 (N_16623,N_16455,N_16458);
nand U16624 (N_16624,N_16440,N_16378);
or U16625 (N_16625,N_16438,N_16468);
xor U16626 (N_16626,N_16347,N_16336);
nand U16627 (N_16627,N_16278,N_16289);
nand U16628 (N_16628,N_16263,N_16319);
nand U16629 (N_16629,N_16490,N_16317);
nor U16630 (N_16630,N_16435,N_16301);
xnor U16631 (N_16631,N_16490,N_16314);
and U16632 (N_16632,N_16478,N_16343);
or U16633 (N_16633,N_16474,N_16396);
or U16634 (N_16634,N_16306,N_16477);
nand U16635 (N_16635,N_16388,N_16292);
nor U16636 (N_16636,N_16316,N_16489);
nor U16637 (N_16637,N_16459,N_16488);
or U16638 (N_16638,N_16457,N_16431);
nand U16639 (N_16639,N_16299,N_16389);
nand U16640 (N_16640,N_16386,N_16398);
and U16641 (N_16641,N_16352,N_16392);
xnor U16642 (N_16642,N_16407,N_16372);
or U16643 (N_16643,N_16379,N_16319);
xor U16644 (N_16644,N_16344,N_16266);
and U16645 (N_16645,N_16274,N_16470);
or U16646 (N_16646,N_16313,N_16280);
nor U16647 (N_16647,N_16499,N_16452);
or U16648 (N_16648,N_16498,N_16416);
nand U16649 (N_16649,N_16345,N_16297);
xor U16650 (N_16650,N_16339,N_16378);
or U16651 (N_16651,N_16411,N_16362);
or U16652 (N_16652,N_16403,N_16421);
nor U16653 (N_16653,N_16251,N_16487);
nor U16654 (N_16654,N_16323,N_16273);
nand U16655 (N_16655,N_16418,N_16307);
nor U16656 (N_16656,N_16473,N_16343);
and U16657 (N_16657,N_16280,N_16357);
and U16658 (N_16658,N_16267,N_16372);
nor U16659 (N_16659,N_16347,N_16457);
or U16660 (N_16660,N_16386,N_16397);
xnor U16661 (N_16661,N_16456,N_16497);
and U16662 (N_16662,N_16252,N_16338);
nand U16663 (N_16663,N_16288,N_16306);
nand U16664 (N_16664,N_16349,N_16369);
nor U16665 (N_16665,N_16384,N_16453);
and U16666 (N_16666,N_16367,N_16374);
nand U16667 (N_16667,N_16293,N_16366);
nand U16668 (N_16668,N_16449,N_16329);
nor U16669 (N_16669,N_16390,N_16380);
or U16670 (N_16670,N_16360,N_16370);
and U16671 (N_16671,N_16303,N_16472);
nor U16672 (N_16672,N_16356,N_16486);
or U16673 (N_16673,N_16397,N_16361);
and U16674 (N_16674,N_16442,N_16413);
nand U16675 (N_16675,N_16331,N_16302);
and U16676 (N_16676,N_16329,N_16383);
nor U16677 (N_16677,N_16432,N_16448);
nand U16678 (N_16678,N_16498,N_16380);
nand U16679 (N_16679,N_16449,N_16389);
xor U16680 (N_16680,N_16373,N_16451);
nor U16681 (N_16681,N_16369,N_16475);
nor U16682 (N_16682,N_16447,N_16292);
nand U16683 (N_16683,N_16359,N_16483);
nand U16684 (N_16684,N_16289,N_16380);
nor U16685 (N_16685,N_16477,N_16446);
or U16686 (N_16686,N_16317,N_16415);
xnor U16687 (N_16687,N_16418,N_16344);
or U16688 (N_16688,N_16370,N_16297);
and U16689 (N_16689,N_16493,N_16270);
or U16690 (N_16690,N_16499,N_16296);
or U16691 (N_16691,N_16318,N_16473);
or U16692 (N_16692,N_16322,N_16467);
xnor U16693 (N_16693,N_16261,N_16433);
nand U16694 (N_16694,N_16454,N_16396);
nand U16695 (N_16695,N_16425,N_16257);
nand U16696 (N_16696,N_16279,N_16322);
or U16697 (N_16697,N_16259,N_16454);
nand U16698 (N_16698,N_16292,N_16252);
xnor U16699 (N_16699,N_16356,N_16283);
or U16700 (N_16700,N_16265,N_16355);
or U16701 (N_16701,N_16325,N_16471);
and U16702 (N_16702,N_16399,N_16418);
nand U16703 (N_16703,N_16481,N_16474);
or U16704 (N_16704,N_16316,N_16404);
nor U16705 (N_16705,N_16345,N_16254);
nor U16706 (N_16706,N_16444,N_16401);
nor U16707 (N_16707,N_16395,N_16381);
nor U16708 (N_16708,N_16409,N_16287);
or U16709 (N_16709,N_16401,N_16405);
nor U16710 (N_16710,N_16415,N_16297);
nor U16711 (N_16711,N_16435,N_16429);
and U16712 (N_16712,N_16308,N_16488);
and U16713 (N_16713,N_16256,N_16276);
nand U16714 (N_16714,N_16270,N_16403);
nand U16715 (N_16715,N_16486,N_16456);
nor U16716 (N_16716,N_16261,N_16305);
and U16717 (N_16717,N_16444,N_16351);
nand U16718 (N_16718,N_16263,N_16434);
xnor U16719 (N_16719,N_16303,N_16487);
nor U16720 (N_16720,N_16387,N_16336);
or U16721 (N_16721,N_16498,N_16424);
nand U16722 (N_16722,N_16459,N_16475);
xnor U16723 (N_16723,N_16291,N_16268);
and U16724 (N_16724,N_16393,N_16443);
or U16725 (N_16725,N_16407,N_16384);
nor U16726 (N_16726,N_16478,N_16294);
and U16727 (N_16727,N_16495,N_16337);
or U16728 (N_16728,N_16295,N_16463);
and U16729 (N_16729,N_16420,N_16251);
and U16730 (N_16730,N_16336,N_16373);
or U16731 (N_16731,N_16365,N_16467);
and U16732 (N_16732,N_16264,N_16273);
nand U16733 (N_16733,N_16293,N_16395);
and U16734 (N_16734,N_16283,N_16273);
nand U16735 (N_16735,N_16345,N_16479);
nand U16736 (N_16736,N_16452,N_16486);
nand U16737 (N_16737,N_16386,N_16305);
or U16738 (N_16738,N_16443,N_16413);
or U16739 (N_16739,N_16397,N_16297);
or U16740 (N_16740,N_16429,N_16326);
nor U16741 (N_16741,N_16454,N_16271);
nand U16742 (N_16742,N_16456,N_16343);
nor U16743 (N_16743,N_16499,N_16439);
or U16744 (N_16744,N_16393,N_16364);
and U16745 (N_16745,N_16424,N_16257);
nor U16746 (N_16746,N_16447,N_16314);
xor U16747 (N_16747,N_16327,N_16297);
and U16748 (N_16748,N_16371,N_16374);
and U16749 (N_16749,N_16316,N_16301);
or U16750 (N_16750,N_16687,N_16733);
or U16751 (N_16751,N_16545,N_16503);
xnor U16752 (N_16752,N_16728,N_16620);
xnor U16753 (N_16753,N_16670,N_16624);
nor U16754 (N_16754,N_16515,N_16698);
and U16755 (N_16755,N_16519,N_16608);
or U16756 (N_16756,N_16638,N_16743);
xnor U16757 (N_16757,N_16626,N_16534);
or U16758 (N_16758,N_16532,N_16573);
or U16759 (N_16759,N_16558,N_16658);
nand U16760 (N_16760,N_16619,N_16560);
and U16761 (N_16761,N_16568,N_16566);
nor U16762 (N_16762,N_16600,N_16644);
nor U16763 (N_16763,N_16712,N_16749);
and U16764 (N_16764,N_16565,N_16648);
xnor U16765 (N_16765,N_16502,N_16668);
and U16766 (N_16766,N_16738,N_16747);
and U16767 (N_16767,N_16744,N_16617);
nand U16768 (N_16768,N_16739,N_16705);
and U16769 (N_16769,N_16537,N_16625);
nor U16770 (N_16770,N_16690,N_16682);
and U16771 (N_16771,N_16587,N_16673);
nor U16772 (N_16772,N_16621,N_16539);
and U16773 (N_16773,N_16671,N_16601);
or U16774 (N_16774,N_16632,N_16631);
or U16775 (N_16775,N_16618,N_16692);
nor U16776 (N_16776,N_16736,N_16581);
nand U16777 (N_16777,N_16527,N_16630);
or U16778 (N_16778,N_16717,N_16583);
xnor U16779 (N_16779,N_16521,N_16641);
or U16780 (N_16780,N_16605,N_16589);
xnor U16781 (N_16781,N_16740,N_16535);
or U16782 (N_16782,N_16741,N_16613);
xor U16783 (N_16783,N_16616,N_16688);
xnor U16784 (N_16784,N_16681,N_16652);
nand U16785 (N_16785,N_16557,N_16533);
or U16786 (N_16786,N_16546,N_16659);
and U16787 (N_16787,N_16639,N_16707);
xor U16788 (N_16788,N_16647,N_16636);
and U16789 (N_16789,N_16724,N_16593);
xor U16790 (N_16790,N_16645,N_16501);
and U16791 (N_16791,N_16525,N_16598);
and U16792 (N_16792,N_16646,N_16553);
and U16793 (N_16793,N_16595,N_16722);
nor U16794 (N_16794,N_16518,N_16703);
nand U16795 (N_16795,N_16552,N_16567);
xor U16796 (N_16796,N_16540,N_16513);
nand U16797 (N_16797,N_16662,N_16665);
or U16798 (N_16798,N_16708,N_16505);
or U16799 (N_16799,N_16653,N_16654);
nor U16800 (N_16800,N_16623,N_16561);
or U16801 (N_16801,N_16602,N_16522);
nand U16802 (N_16802,N_16675,N_16548);
and U16803 (N_16803,N_16742,N_16651);
nor U16804 (N_16804,N_16701,N_16711);
or U16805 (N_16805,N_16536,N_16649);
and U16806 (N_16806,N_16607,N_16661);
and U16807 (N_16807,N_16529,N_16516);
nor U16808 (N_16808,N_16735,N_16563);
or U16809 (N_16809,N_16695,N_16547);
nand U16810 (N_16810,N_16564,N_16572);
and U16811 (N_16811,N_16730,N_16680);
or U16812 (N_16812,N_16660,N_16666);
nand U16813 (N_16813,N_16603,N_16655);
and U16814 (N_16814,N_16562,N_16554);
xnor U16815 (N_16815,N_16584,N_16732);
or U16816 (N_16816,N_16596,N_16628);
or U16817 (N_16817,N_16578,N_16556);
nor U16818 (N_16818,N_16576,N_16574);
and U16819 (N_16819,N_16615,N_16569);
xor U16820 (N_16820,N_16676,N_16721);
or U16821 (N_16821,N_16650,N_16543);
nand U16822 (N_16822,N_16686,N_16716);
nand U16823 (N_16823,N_16571,N_16580);
or U16824 (N_16824,N_16577,N_16590);
and U16825 (N_16825,N_16635,N_16511);
xor U16826 (N_16826,N_16517,N_16640);
xor U16827 (N_16827,N_16642,N_16585);
nor U16828 (N_16828,N_16592,N_16672);
and U16829 (N_16829,N_16702,N_16542);
or U16830 (N_16830,N_16684,N_16657);
and U16831 (N_16831,N_16700,N_16586);
xor U16832 (N_16832,N_16669,N_16531);
and U16833 (N_16833,N_16549,N_16704);
nor U16834 (N_16834,N_16677,N_16709);
xnor U16835 (N_16835,N_16510,N_16663);
nor U16836 (N_16836,N_16610,N_16622);
and U16837 (N_16837,N_16696,N_16746);
xnor U16838 (N_16838,N_16559,N_16725);
and U16839 (N_16839,N_16570,N_16674);
and U16840 (N_16840,N_16678,N_16727);
and U16841 (N_16841,N_16582,N_16504);
xor U16842 (N_16842,N_16734,N_16530);
and U16843 (N_16843,N_16575,N_16611);
nor U16844 (N_16844,N_16667,N_16656);
or U16845 (N_16845,N_16633,N_16689);
nor U16846 (N_16846,N_16514,N_16591);
and U16847 (N_16847,N_16500,N_16588);
xor U16848 (N_16848,N_16637,N_16731);
or U16849 (N_16849,N_16664,N_16526);
nand U16850 (N_16850,N_16685,N_16550);
nand U16851 (N_16851,N_16551,N_16634);
nand U16852 (N_16852,N_16629,N_16520);
nor U16853 (N_16853,N_16579,N_16544);
xnor U16854 (N_16854,N_16729,N_16599);
xnor U16855 (N_16855,N_16714,N_16726);
nor U16856 (N_16856,N_16523,N_16541);
nand U16857 (N_16857,N_16509,N_16507);
nor U16858 (N_16858,N_16612,N_16528);
xnor U16859 (N_16859,N_16597,N_16723);
nand U16860 (N_16860,N_16614,N_16718);
and U16861 (N_16861,N_16713,N_16643);
nor U16862 (N_16862,N_16606,N_16555);
xnor U16863 (N_16863,N_16697,N_16609);
nand U16864 (N_16864,N_16699,N_16627);
nor U16865 (N_16865,N_16679,N_16710);
nor U16866 (N_16866,N_16524,N_16694);
xor U16867 (N_16867,N_16719,N_16594);
nor U16868 (N_16868,N_16512,N_16508);
or U16869 (N_16869,N_16691,N_16604);
or U16870 (N_16870,N_16693,N_16538);
and U16871 (N_16871,N_16745,N_16748);
nor U16872 (N_16872,N_16683,N_16715);
nor U16873 (N_16873,N_16706,N_16737);
or U16874 (N_16874,N_16720,N_16506);
and U16875 (N_16875,N_16597,N_16632);
nand U16876 (N_16876,N_16707,N_16732);
nand U16877 (N_16877,N_16528,N_16565);
or U16878 (N_16878,N_16559,N_16564);
or U16879 (N_16879,N_16544,N_16687);
nand U16880 (N_16880,N_16688,N_16745);
and U16881 (N_16881,N_16594,N_16554);
or U16882 (N_16882,N_16738,N_16543);
or U16883 (N_16883,N_16553,N_16504);
nand U16884 (N_16884,N_16573,N_16571);
xnor U16885 (N_16885,N_16740,N_16729);
nor U16886 (N_16886,N_16519,N_16626);
xor U16887 (N_16887,N_16587,N_16573);
and U16888 (N_16888,N_16526,N_16740);
nand U16889 (N_16889,N_16626,N_16613);
nor U16890 (N_16890,N_16546,N_16647);
nor U16891 (N_16891,N_16515,N_16659);
xnor U16892 (N_16892,N_16597,N_16546);
nand U16893 (N_16893,N_16565,N_16607);
xor U16894 (N_16894,N_16636,N_16514);
and U16895 (N_16895,N_16527,N_16621);
xor U16896 (N_16896,N_16595,N_16574);
or U16897 (N_16897,N_16519,N_16607);
xor U16898 (N_16898,N_16502,N_16609);
nor U16899 (N_16899,N_16746,N_16526);
xor U16900 (N_16900,N_16626,N_16728);
nand U16901 (N_16901,N_16611,N_16580);
or U16902 (N_16902,N_16505,N_16650);
nor U16903 (N_16903,N_16666,N_16704);
nor U16904 (N_16904,N_16561,N_16546);
nand U16905 (N_16905,N_16520,N_16610);
nand U16906 (N_16906,N_16711,N_16607);
nor U16907 (N_16907,N_16661,N_16635);
or U16908 (N_16908,N_16684,N_16506);
and U16909 (N_16909,N_16554,N_16545);
or U16910 (N_16910,N_16704,N_16679);
or U16911 (N_16911,N_16681,N_16742);
or U16912 (N_16912,N_16514,N_16639);
nor U16913 (N_16913,N_16737,N_16732);
xor U16914 (N_16914,N_16632,N_16650);
xnor U16915 (N_16915,N_16712,N_16711);
and U16916 (N_16916,N_16597,N_16611);
and U16917 (N_16917,N_16569,N_16733);
nor U16918 (N_16918,N_16623,N_16638);
or U16919 (N_16919,N_16586,N_16553);
nor U16920 (N_16920,N_16725,N_16570);
nor U16921 (N_16921,N_16568,N_16595);
or U16922 (N_16922,N_16520,N_16579);
xor U16923 (N_16923,N_16576,N_16734);
and U16924 (N_16924,N_16687,N_16703);
and U16925 (N_16925,N_16565,N_16697);
nand U16926 (N_16926,N_16591,N_16655);
nand U16927 (N_16927,N_16701,N_16649);
nor U16928 (N_16928,N_16663,N_16604);
nand U16929 (N_16929,N_16589,N_16541);
nor U16930 (N_16930,N_16545,N_16603);
nand U16931 (N_16931,N_16531,N_16710);
or U16932 (N_16932,N_16663,N_16601);
or U16933 (N_16933,N_16661,N_16634);
xor U16934 (N_16934,N_16557,N_16502);
xor U16935 (N_16935,N_16602,N_16521);
nor U16936 (N_16936,N_16643,N_16545);
nor U16937 (N_16937,N_16545,N_16505);
nand U16938 (N_16938,N_16587,N_16541);
xnor U16939 (N_16939,N_16661,N_16588);
or U16940 (N_16940,N_16616,N_16519);
nand U16941 (N_16941,N_16581,N_16727);
and U16942 (N_16942,N_16670,N_16729);
xnor U16943 (N_16943,N_16737,N_16504);
xnor U16944 (N_16944,N_16528,N_16695);
and U16945 (N_16945,N_16629,N_16528);
nand U16946 (N_16946,N_16543,N_16649);
and U16947 (N_16947,N_16522,N_16745);
xnor U16948 (N_16948,N_16649,N_16707);
xor U16949 (N_16949,N_16674,N_16732);
nand U16950 (N_16950,N_16734,N_16545);
xnor U16951 (N_16951,N_16721,N_16575);
nor U16952 (N_16952,N_16687,N_16630);
nor U16953 (N_16953,N_16512,N_16672);
nor U16954 (N_16954,N_16726,N_16529);
nor U16955 (N_16955,N_16708,N_16733);
xnor U16956 (N_16956,N_16737,N_16593);
nand U16957 (N_16957,N_16648,N_16635);
and U16958 (N_16958,N_16535,N_16633);
xor U16959 (N_16959,N_16635,N_16729);
xor U16960 (N_16960,N_16631,N_16607);
nand U16961 (N_16961,N_16645,N_16529);
nand U16962 (N_16962,N_16573,N_16594);
nand U16963 (N_16963,N_16699,N_16581);
or U16964 (N_16964,N_16651,N_16716);
nand U16965 (N_16965,N_16690,N_16559);
nor U16966 (N_16966,N_16511,N_16657);
xor U16967 (N_16967,N_16632,N_16688);
nand U16968 (N_16968,N_16562,N_16548);
or U16969 (N_16969,N_16618,N_16749);
and U16970 (N_16970,N_16525,N_16658);
or U16971 (N_16971,N_16685,N_16507);
nand U16972 (N_16972,N_16634,N_16719);
and U16973 (N_16973,N_16538,N_16551);
nand U16974 (N_16974,N_16621,N_16584);
xor U16975 (N_16975,N_16564,N_16551);
nor U16976 (N_16976,N_16579,N_16657);
nor U16977 (N_16977,N_16661,N_16563);
or U16978 (N_16978,N_16599,N_16649);
nand U16979 (N_16979,N_16601,N_16578);
xor U16980 (N_16980,N_16632,N_16729);
and U16981 (N_16981,N_16635,N_16639);
and U16982 (N_16982,N_16661,N_16745);
or U16983 (N_16983,N_16591,N_16745);
or U16984 (N_16984,N_16739,N_16731);
or U16985 (N_16985,N_16600,N_16555);
xor U16986 (N_16986,N_16617,N_16628);
or U16987 (N_16987,N_16606,N_16607);
and U16988 (N_16988,N_16712,N_16602);
and U16989 (N_16989,N_16514,N_16700);
nor U16990 (N_16990,N_16574,N_16725);
nand U16991 (N_16991,N_16623,N_16654);
nor U16992 (N_16992,N_16688,N_16716);
or U16993 (N_16993,N_16636,N_16722);
nand U16994 (N_16994,N_16539,N_16538);
nor U16995 (N_16995,N_16742,N_16558);
nor U16996 (N_16996,N_16724,N_16609);
xnor U16997 (N_16997,N_16728,N_16665);
or U16998 (N_16998,N_16688,N_16736);
or U16999 (N_16999,N_16531,N_16641);
nand U17000 (N_17000,N_16855,N_16788);
or U17001 (N_17001,N_16885,N_16955);
and U17002 (N_17002,N_16781,N_16802);
and U17003 (N_17003,N_16764,N_16875);
or U17004 (N_17004,N_16895,N_16849);
or U17005 (N_17005,N_16840,N_16925);
or U17006 (N_17006,N_16751,N_16820);
xnor U17007 (N_17007,N_16923,N_16886);
or U17008 (N_17008,N_16898,N_16932);
nor U17009 (N_17009,N_16954,N_16993);
nor U17010 (N_17010,N_16783,N_16911);
xnor U17011 (N_17011,N_16900,N_16877);
nor U17012 (N_17012,N_16887,N_16874);
or U17013 (N_17013,N_16947,N_16981);
or U17014 (N_17014,N_16978,N_16817);
and U17015 (N_17015,N_16903,N_16798);
nor U17016 (N_17016,N_16857,N_16796);
nor U17017 (N_17017,N_16964,N_16893);
nor U17018 (N_17018,N_16823,N_16844);
and U17019 (N_17019,N_16858,N_16945);
and U17020 (N_17020,N_16938,N_16969);
nand U17021 (N_17021,N_16987,N_16977);
and U17022 (N_17022,N_16755,N_16944);
nor U17023 (N_17023,N_16940,N_16810);
and U17024 (N_17024,N_16864,N_16910);
nor U17025 (N_17025,N_16759,N_16998);
nor U17026 (N_17026,N_16851,N_16958);
nand U17027 (N_17027,N_16989,N_16841);
or U17028 (N_17028,N_16881,N_16884);
or U17029 (N_17029,N_16790,N_16965);
and U17030 (N_17030,N_16752,N_16776);
and U17031 (N_17031,N_16917,N_16768);
or U17032 (N_17032,N_16913,N_16986);
nor U17033 (N_17033,N_16761,N_16856);
and U17034 (N_17034,N_16896,N_16935);
xor U17035 (N_17035,N_16951,N_16952);
or U17036 (N_17036,N_16953,N_16890);
nand U17037 (N_17037,N_16804,N_16828);
xor U17038 (N_17038,N_16985,N_16765);
or U17039 (N_17039,N_16907,N_16774);
or U17040 (N_17040,N_16914,N_16860);
and U17041 (N_17041,N_16793,N_16769);
or U17042 (N_17042,N_16919,N_16878);
nor U17043 (N_17043,N_16797,N_16865);
nor U17044 (N_17044,N_16807,N_16901);
nor U17045 (N_17045,N_16967,N_16848);
nand U17046 (N_17046,N_16800,N_16867);
xor U17047 (N_17047,N_16791,N_16921);
xor U17048 (N_17048,N_16818,N_16786);
xor U17049 (N_17049,N_16760,N_16920);
xor U17050 (N_17050,N_16813,N_16970);
xor U17051 (N_17051,N_16942,N_16972);
xnor U17052 (N_17052,N_16974,N_16843);
and U17053 (N_17053,N_16780,N_16888);
nand U17054 (N_17054,N_16824,N_16766);
or U17055 (N_17055,N_16853,N_16763);
xnor U17056 (N_17056,N_16908,N_16968);
xor U17057 (N_17057,N_16767,N_16931);
nor U17058 (N_17058,N_16883,N_16984);
nor U17059 (N_17059,N_16775,N_16909);
and U17060 (N_17060,N_16982,N_16927);
xnor U17061 (N_17061,N_16937,N_16936);
nor U17062 (N_17062,N_16816,N_16959);
or U17063 (N_17063,N_16957,N_16836);
xor U17064 (N_17064,N_16859,N_16868);
or U17065 (N_17065,N_16812,N_16756);
xor U17066 (N_17066,N_16929,N_16811);
or U17067 (N_17067,N_16999,N_16994);
nand U17068 (N_17068,N_16789,N_16930);
nor U17069 (N_17069,N_16837,N_16905);
nand U17070 (N_17070,N_16990,N_16916);
nor U17071 (N_17071,N_16971,N_16762);
nor U17072 (N_17072,N_16808,N_16803);
nor U17073 (N_17073,N_16961,N_16809);
nor U17074 (N_17074,N_16821,N_16946);
or U17075 (N_17075,N_16778,N_16826);
or U17076 (N_17076,N_16934,N_16805);
and U17077 (N_17077,N_16871,N_16842);
nand U17078 (N_17078,N_16845,N_16799);
or U17079 (N_17079,N_16996,N_16960);
xor U17080 (N_17080,N_16854,N_16831);
nand U17081 (N_17081,N_16819,N_16777);
xor U17082 (N_17082,N_16897,N_16825);
and U17083 (N_17083,N_16794,N_16861);
or U17084 (N_17084,N_16879,N_16889);
nand U17085 (N_17085,N_16850,N_16912);
nor U17086 (N_17086,N_16991,N_16770);
xor U17087 (N_17087,N_16852,N_16975);
nor U17088 (N_17088,N_16976,N_16997);
and U17089 (N_17089,N_16948,N_16894);
nor U17090 (N_17090,N_16785,N_16966);
nand U17091 (N_17091,N_16830,N_16795);
nand U17092 (N_17092,N_16787,N_16847);
or U17093 (N_17093,N_16979,N_16902);
xnor U17094 (N_17094,N_16792,N_16995);
nor U17095 (N_17095,N_16772,N_16815);
or U17096 (N_17096,N_16782,N_16872);
or U17097 (N_17097,N_16906,N_16835);
nor U17098 (N_17098,N_16801,N_16892);
and U17099 (N_17099,N_16939,N_16827);
and U17100 (N_17100,N_16773,N_16928);
or U17101 (N_17101,N_16882,N_16834);
xor U17102 (N_17102,N_16754,N_16838);
nand U17103 (N_17103,N_16870,N_16784);
xor U17104 (N_17104,N_16822,N_16839);
nor U17105 (N_17105,N_16933,N_16926);
and U17106 (N_17106,N_16750,N_16973);
nor U17107 (N_17107,N_16757,N_16846);
nand U17108 (N_17108,N_16873,N_16771);
xnor U17109 (N_17109,N_16899,N_16814);
nor U17110 (N_17110,N_16988,N_16943);
nor U17111 (N_17111,N_16779,N_16922);
and U17112 (N_17112,N_16918,N_16862);
and U17113 (N_17113,N_16962,N_16832);
xnor U17114 (N_17114,N_16950,N_16880);
or U17115 (N_17115,N_16863,N_16876);
and U17116 (N_17116,N_16866,N_16963);
nor U17117 (N_17117,N_16753,N_16949);
xnor U17118 (N_17118,N_16869,N_16758);
xnor U17119 (N_17119,N_16992,N_16983);
or U17120 (N_17120,N_16891,N_16980);
or U17121 (N_17121,N_16806,N_16829);
or U17122 (N_17122,N_16833,N_16904);
xor U17123 (N_17123,N_16956,N_16915);
nand U17124 (N_17124,N_16941,N_16924);
nor U17125 (N_17125,N_16755,N_16991);
nor U17126 (N_17126,N_16917,N_16836);
and U17127 (N_17127,N_16818,N_16856);
and U17128 (N_17128,N_16843,N_16766);
nor U17129 (N_17129,N_16864,N_16962);
or U17130 (N_17130,N_16919,N_16957);
and U17131 (N_17131,N_16798,N_16931);
or U17132 (N_17132,N_16888,N_16945);
nand U17133 (N_17133,N_16786,N_16935);
or U17134 (N_17134,N_16962,N_16876);
and U17135 (N_17135,N_16801,N_16799);
xnor U17136 (N_17136,N_16942,N_16770);
nand U17137 (N_17137,N_16823,N_16857);
nand U17138 (N_17138,N_16864,N_16819);
nor U17139 (N_17139,N_16755,N_16879);
nand U17140 (N_17140,N_16846,N_16956);
or U17141 (N_17141,N_16876,N_16981);
or U17142 (N_17142,N_16786,N_16767);
and U17143 (N_17143,N_16964,N_16909);
and U17144 (N_17144,N_16854,N_16906);
or U17145 (N_17145,N_16925,N_16954);
and U17146 (N_17146,N_16978,N_16859);
nor U17147 (N_17147,N_16909,N_16951);
nand U17148 (N_17148,N_16987,N_16789);
nand U17149 (N_17149,N_16865,N_16778);
and U17150 (N_17150,N_16874,N_16780);
xnor U17151 (N_17151,N_16957,N_16913);
xnor U17152 (N_17152,N_16922,N_16926);
xnor U17153 (N_17153,N_16963,N_16940);
or U17154 (N_17154,N_16939,N_16885);
nor U17155 (N_17155,N_16819,N_16982);
and U17156 (N_17156,N_16866,N_16854);
xnor U17157 (N_17157,N_16859,N_16812);
xnor U17158 (N_17158,N_16780,N_16929);
or U17159 (N_17159,N_16843,N_16958);
nor U17160 (N_17160,N_16984,N_16772);
nor U17161 (N_17161,N_16946,N_16778);
nand U17162 (N_17162,N_16833,N_16936);
and U17163 (N_17163,N_16802,N_16896);
xor U17164 (N_17164,N_16775,N_16853);
nand U17165 (N_17165,N_16937,N_16865);
and U17166 (N_17166,N_16914,N_16894);
or U17167 (N_17167,N_16826,N_16844);
or U17168 (N_17168,N_16810,N_16804);
and U17169 (N_17169,N_16931,N_16927);
nand U17170 (N_17170,N_16781,N_16965);
or U17171 (N_17171,N_16828,N_16820);
nor U17172 (N_17172,N_16947,N_16940);
and U17173 (N_17173,N_16951,N_16957);
or U17174 (N_17174,N_16888,N_16764);
and U17175 (N_17175,N_16947,N_16930);
nor U17176 (N_17176,N_16834,N_16950);
nor U17177 (N_17177,N_16754,N_16971);
or U17178 (N_17178,N_16851,N_16815);
or U17179 (N_17179,N_16884,N_16826);
or U17180 (N_17180,N_16825,N_16885);
xor U17181 (N_17181,N_16912,N_16849);
nor U17182 (N_17182,N_16969,N_16947);
and U17183 (N_17183,N_16764,N_16826);
nor U17184 (N_17184,N_16866,N_16936);
or U17185 (N_17185,N_16923,N_16881);
xnor U17186 (N_17186,N_16916,N_16807);
xnor U17187 (N_17187,N_16964,N_16886);
xor U17188 (N_17188,N_16960,N_16834);
or U17189 (N_17189,N_16767,N_16818);
or U17190 (N_17190,N_16929,N_16779);
xor U17191 (N_17191,N_16848,N_16873);
and U17192 (N_17192,N_16854,N_16926);
xor U17193 (N_17193,N_16875,N_16780);
or U17194 (N_17194,N_16964,N_16953);
xnor U17195 (N_17195,N_16887,N_16948);
nor U17196 (N_17196,N_16832,N_16890);
nand U17197 (N_17197,N_16920,N_16753);
or U17198 (N_17198,N_16993,N_16776);
xnor U17199 (N_17199,N_16844,N_16983);
or U17200 (N_17200,N_16961,N_16953);
nand U17201 (N_17201,N_16791,N_16859);
and U17202 (N_17202,N_16952,N_16873);
and U17203 (N_17203,N_16917,N_16756);
nand U17204 (N_17204,N_16798,N_16924);
xor U17205 (N_17205,N_16756,N_16870);
or U17206 (N_17206,N_16872,N_16973);
or U17207 (N_17207,N_16913,N_16962);
nor U17208 (N_17208,N_16877,N_16929);
or U17209 (N_17209,N_16875,N_16866);
nand U17210 (N_17210,N_16832,N_16888);
or U17211 (N_17211,N_16808,N_16770);
nand U17212 (N_17212,N_16828,N_16846);
nor U17213 (N_17213,N_16788,N_16828);
or U17214 (N_17214,N_16906,N_16977);
nor U17215 (N_17215,N_16767,N_16925);
and U17216 (N_17216,N_16897,N_16818);
or U17217 (N_17217,N_16801,N_16776);
or U17218 (N_17218,N_16835,N_16816);
xor U17219 (N_17219,N_16968,N_16834);
xor U17220 (N_17220,N_16761,N_16767);
xnor U17221 (N_17221,N_16860,N_16751);
or U17222 (N_17222,N_16985,N_16786);
and U17223 (N_17223,N_16792,N_16881);
nand U17224 (N_17224,N_16825,N_16866);
nor U17225 (N_17225,N_16904,N_16959);
nand U17226 (N_17226,N_16912,N_16914);
xnor U17227 (N_17227,N_16835,N_16864);
or U17228 (N_17228,N_16945,N_16943);
and U17229 (N_17229,N_16923,N_16761);
xnor U17230 (N_17230,N_16867,N_16751);
nand U17231 (N_17231,N_16989,N_16811);
xor U17232 (N_17232,N_16958,N_16820);
nand U17233 (N_17233,N_16914,N_16774);
xnor U17234 (N_17234,N_16937,N_16804);
and U17235 (N_17235,N_16893,N_16828);
nor U17236 (N_17236,N_16875,N_16863);
nor U17237 (N_17237,N_16957,N_16984);
nand U17238 (N_17238,N_16750,N_16919);
and U17239 (N_17239,N_16827,N_16811);
xnor U17240 (N_17240,N_16874,N_16836);
nor U17241 (N_17241,N_16930,N_16824);
or U17242 (N_17242,N_16902,N_16941);
or U17243 (N_17243,N_16801,N_16835);
or U17244 (N_17244,N_16929,N_16810);
or U17245 (N_17245,N_16869,N_16974);
and U17246 (N_17246,N_16862,N_16867);
and U17247 (N_17247,N_16809,N_16816);
nor U17248 (N_17248,N_16774,N_16953);
xnor U17249 (N_17249,N_16907,N_16871);
or U17250 (N_17250,N_17027,N_17102);
xnor U17251 (N_17251,N_17196,N_17159);
or U17252 (N_17252,N_17187,N_17123);
and U17253 (N_17253,N_17144,N_17107);
and U17254 (N_17254,N_17248,N_17229);
and U17255 (N_17255,N_17199,N_17191);
nor U17256 (N_17256,N_17099,N_17177);
or U17257 (N_17257,N_17044,N_17008);
and U17258 (N_17258,N_17217,N_17151);
nor U17259 (N_17259,N_17090,N_17215);
or U17260 (N_17260,N_17019,N_17233);
and U17261 (N_17261,N_17238,N_17064);
nand U17262 (N_17262,N_17202,N_17087);
nand U17263 (N_17263,N_17015,N_17097);
xnor U17264 (N_17264,N_17188,N_17034);
nor U17265 (N_17265,N_17111,N_17103);
nand U17266 (N_17266,N_17013,N_17166);
and U17267 (N_17267,N_17112,N_17216);
or U17268 (N_17268,N_17074,N_17073);
or U17269 (N_17269,N_17220,N_17095);
and U17270 (N_17270,N_17232,N_17084);
nor U17271 (N_17271,N_17228,N_17040);
and U17272 (N_17272,N_17176,N_17056);
and U17273 (N_17273,N_17194,N_17240);
and U17274 (N_17274,N_17125,N_17162);
and U17275 (N_17275,N_17136,N_17208);
and U17276 (N_17276,N_17165,N_17158);
and U17277 (N_17277,N_17006,N_17038);
nand U17278 (N_17278,N_17052,N_17204);
nor U17279 (N_17279,N_17245,N_17189);
xnor U17280 (N_17280,N_17219,N_17031);
nor U17281 (N_17281,N_17209,N_17161);
and U17282 (N_17282,N_17007,N_17010);
nor U17283 (N_17283,N_17163,N_17047);
nand U17284 (N_17284,N_17184,N_17033);
xor U17285 (N_17285,N_17004,N_17234);
or U17286 (N_17286,N_17000,N_17201);
nand U17287 (N_17287,N_17172,N_17156);
nor U17288 (N_17288,N_17226,N_17003);
or U17289 (N_17289,N_17032,N_17167);
nor U17290 (N_17290,N_17021,N_17115);
and U17291 (N_17291,N_17246,N_17028);
xnor U17292 (N_17292,N_17025,N_17221);
xnor U17293 (N_17293,N_17049,N_17181);
and U17294 (N_17294,N_17133,N_17236);
and U17295 (N_17295,N_17001,N_17243);
nor U17296 (N_17296,N_17080,N_17134);
or U17297 (N_17297,N_17071,N_17148);
nor U17298 (N_17298,N_17182,N_17160);
and U17299 (N_17299,N_17145,N_17141);
or U17300 (N_17300,N_17164,N_17016);
xnor U17301 (N_17301,N_17244,N_17197);
and U17302 (N_17302,N_17149,N_17089);
or U17303 (N_17303,N_17092,N_17241);
or U17304 (N_17304,N_17193,N_17169);
or U17305 (N_17305,N_17178,N_17043);
nand U17306 (N_17306,N_17078,N_17121);
xnor U17307 (N_17307,N_17114,N_17122);
and U17308 (N_17308,N_17146,N_17230);
nand U17309 (N_17309,N_17018,N_17173);
nor U17310 (N_17310,N_17155,N_17058);
nand U17311 (N_17311,N_17214,N_17060);
or U17312 (N_17312,N_17048,N_17113);
xnor U17313 (N_17313,N_17053,N_17152);
and U17314 (N_17314,N_17185,N_17091);
nand U17315 (N_17315,N_17179,N_17037);
or U17316 (N_17316,N_17190,N_17035);
nand U17317 (N_17317,N_17222,N_17100);
or U17318 (N_17318,N_17067,N_17126);
nand U17319 (N_17319,N_17235,N_17105);
nor U17320 (N_17320,N_17098,N_17192);
xnor U17321 (N_17321,N_17137,N_17130);
or U17322 (N_17322,N_17046,N_17171);
nor U17323 (N_17323,N_17022,N_17094);
nand U17324 (N_17324,N_17083,N_17120);
or U17325 (N_17325,N_17104,N_17030);
xor U17326 (N_17326,N_17142,N_17011);
or U17327 (N_17327,N_17174,N_17157);
nand U17328 (N_17328,N_17088,N_17128);
xnor U17329 (N_17329,N_17070,N_17050);
or U17330 (N_17330,N_17205,N_17012);
nand U17331 (N_17331,N_17153,N_17138);
and U17332 (N_17332,N_17247,N_17079);
nor U17333 (N_17333,N_17020,N_17101);
and U17334 (N_17334,N_17055,N_17132);
and U17335 (N_17335,N_17124,N_17227);
nor U17336 (N_17336,N_17062,N_17042);
or U17337 (N_17337,N_17206,N_17203);
nor U17338 (N_17338,N_17076,N_17116);
or U17339 (N_17339,N_17127,N_17106);
or U17340 (N_17340,N_17065,N_17024);
nor U17341 (N_17341,N_17096,N_17063);
xnor U17342 (N_17342,N_17211,N_17143);
nand U17343 (N_17343,N_17068,N_17005);
nand U17344 (N_17344,N_17045,N_17118);
xor U17345 (N_17345,N_17198,N_17117);
xnor U17346 (N_17346,N_17023,N_17051);
nand U17347 (N_17347,N_17210,N_17186);
and U17348 (N_17348,N_17059,N_17017);
xnor U17349 (N_17349,N_17054,N_17135);
or U17350 (N_17350,N_17093,N_17057);
and U17351 (N_17351,N_17140,N_17223);
xnor U17352 (N_17352,N_17170,N_17077);
or U17353 (N_17353,N_17200,N_17009);
nor U17354 (N_17354,N_17175,N_17036);
xor U17355 (N_17355,N_17237,N_17213);
or U17356 (N_17356,N_17150,N_17131);
nor U17357 (N_17357,N_17129,N_17041);
xor U17358 (N_17358,N_17075,N_17225);
nor U17359 (N_17359,N_17239,N_17242);
or U17360 (N_17360,N_17139,N_17147);
nor U17361 (N_17361,N_17207,N_17224);
nor U17362 (N_17362,N_17081,N_17168);
and U17363 (N_17363,N_17183,N_17072);
xnor U17364 (N_17364,N_17249,N_17002);
xnor U17365 (N_17365,N_17109,N_17014);
and U17366 (N_17366,N_17119,N_17069);
and U17367 (N_17367,N_17108,N_17154);
nand U17368 (N_17368,N_17195,N_17082);
and U17369 (N_17369,N_17085,N_17180);
or U17370 (N_17370,N_17110,N_17231);
xor U17371 (N_17371,N_17026,N_17061);
xnor U17372 (N_17372,N_17218,N_17029);
xnor U17373 (N_17373,N_17066,N_17212);
or U17374 (N_17374,N_17086,N_17039);
nand U17375 (N_17375,N_17147,N_17197);
nand U17376 (N_17376,N_17031,N_17008);
xnor U17377 (N_17377,N_17233,N_17118);
nor U17378 (N_17378,N_17043,N_17187);
or U17379 (N_17379,N_17204,N_17215);
xnor U17380 (N_17380,N_17009,N_17233);
or U17381 (N_17381,N_17205,N_17211);
xnor U17382 (N_17382,N_17243,N_17248);
nor U17383 (N_17383,N_17196,N_17060);
or U17384 (N_17384,N_17005,N_17200);
nor U17385 (N_17385,N_17178,N_17247);
xor U17386 (N_17386,N_17111,N_17146);
or U17387 (N_17387,N_17080,N_17077);
nand U17388 (N_17388,N_17147,N_17155);
xor U17389 (N_17389,N_17097,N_17209);
or U17390 (N_17390,N_17046,N_17066);
nor U17391 (N_17391,N_17045,N_17188);
and U17392 (N_17392,N_17198,N_17134);
nor U17393 (N_17393,N_17026,N_17162);
and U17394 (N_17394,N_17225,N_17243);
or U17395 (N_17395,N_17128,N_17147);
nand U17396 (N_17396,N_17183,N_17009);
nand U17397 (N_17397,N_17120,N_17012);
and U17398 (N_17398,N_17159,N_17111);
or U17399 (N_17399,N_17110,N_17043);
nand U17400 (N_17400,N_17186,N_17167);
xor U17401 (N_17401,N_17171,N_17202);
nor U17402 (N_17402,N_17008,N_17078);
and U17403 (N_17403,N_17185,N_17217);
nor U17404 (N_17404,N_17062,N_17181);
nand U17405 (N_17405,N_17008,N_17134);
nor U17406 (N_17406,N_17242,N_17207);
and U17407 (N_17407,N_17221,N_17248);
xor U17408 (N_17408,N_17032,N_17120);
or U17409 (N_17409,N_17082,N_17023);
xor U17410 (N_17410,N_17062,N_17000);
xnor U17411 (N_17411,N_17021,N_17050);
nor U17412 (N_17412,N_17027,N_17207);
xnor U17413 (N_17413,N_17027,N_17045);
xnor U17414 (N_17414,N_17221,N_17066);
or U17415 (N_17415,N_17092,N_17102);
nor U17416 (N_17416,N_17169,N_17156);
nor U17417 (N_17417,N_17189,N_17168);
and U17418 (N_17418,N_17019,N_17216);
or U17419 (N_17419,N_17203,N_17059);
xor U17420 (N_17420,N_17228,N_17201);
xnor U17421 (N_17421,N_17155,N_17218);
and U17422 (N_17422,N_17000,N_17050);
nand U17423 (N_17423,N_17060,N_17013);
xnor U17424 (N_17424,N_17110,N_17199);
and U17425 (N_17425,N_17091,N_17094);
nand U17426 (N_17426,N_17024,N_17229);
and U17427 (N_17427,N_17116,N_17043);
nor U17428 (N_17428,N_17018,N_17010);
nand U17429 (N_17429,N_17241,N_17081);
or U17430 (N_17430,N_17184,N_17228);
xnor U17431 (N_17431,N_17050,N_17188);
nor U17432 (N_17432,N_17206,N_17172);
nand U17433 (N_17433,N_17058,N_17216);
and U17434 (N_17434,N_17198,N_17212);
nand U17435 (N_17435,N_17058,N_17000);
nand U17436 (N_17436,N_17154,N_17163);
xor U17437 (N_17437,N_17005,N_17244);
nor U17438 (N_17438,N_17176,N_17230);
nand U17439 (N_17439,N_17174,N_17064);
nor U17440 (N_17440,N_17225,N_17052);
or U17441 (N_17441,N_17200,N_17024);
nor U17442 (N_17442,N_17032,N_17070);
xnor U17443 (N_17443,N_17242,N_17127);
xnor U17444 (N_17444,N_17171,N_17198);
xnor U17445 (N_17445,N_17170,N_17141);
nor U17446 (N_17446,N_17094,N_17240);
nand U17447 (N_17447,N_17224,N_17070);
or U17448 (N_17448,N_17154,N_17078);
and U17449 (N_17449,N_17101,N_17127);
xor U17450 (N_17450,N_17172,N_17100);
xor U17451 (N_17451,N_17195,N_17149);
nor U17452 (N_17452,N_17004,N_17057);
or U17453 (N_17453,N_17021,N_17062);
or U17454 (N_17454,N_17016,N_17052);
and U17455 (N_17455,N_17173,N_17132);
nand U17456 (N_17456,N_17087,N_17135);
xnor U17457 (N_17457,N_17152,N_17229);
xnor U17458 (N_17458,N_17109,N_17049);
or U17459 (N_17459,N_17102,N_17107);
nand U17460 (N_17460,N_17007,N_17060);
xnor U17461 (N_17461,N_17148,N_17202);
and U17462 (N_17462,N_17172,N_17144);
xnor U17463 (N_17463,N_17207,N_17190);
xnor U17464 (N_17464,N_17059,N_17122);
nor U17465 (N_17465,N_17155,N_17214);
nand U17466 (N_17466,N_17190,N_17126);
nor U17467 (N_17467,N_17164,N_17224);
or U17468 (N_17468,N_17116,N_17121);
nor U17469 (N_17469,N_17176,N_17192);
xnor U17470 (N_17470,N_17142,N_17031);
nor U17471 (N_17471,N_17036,N_17112);
nand U17472 (N_17472,N_17203,N_17041);
or U17473 (N_17473,N_17183,N_17106);
or U17474 (N_17474,N_17165,N_17129);
nand U17475 (N_17475,N_17206,N_17040);
nand U17476 (N_17476,N_17227,N_17207);
nor U17477 (N_17477,N_17147,N_17134);
xor U17478 (N_17478,N_17201,N_17049);
xnor U17479 (N_17479,N_17040,N_17014);
xor U17480 (N_17480,N_17170,N_17169);
or U17481 (N_17481,N_17221,N_17108);
xnor U17482 (N_17482,N_17159,N_17070);
xor U17483 (N_17483,N_17086,N_17138);
or U17484 (N_17484,N_17129,N_17169);
nand U17485 (N_17485,N_17104,N_17087);
xor U17486 (N_17486,N_17212,N_17023);
nor U17487 (N_17487,N_17049,N_17107);
nand U17488 (N_17488,N_17220,N_17038);
or U17489 (N_17489,N_17105,N_17109);
or U17490 (N_17490,N_17150,N_17233);
nand U17491 (N_17491,N_17117,N_17161);
xnor U17492 (N_17492,N_17094,N_17104);
nor U17493 (N_17493,N_17168,N_17041);
xor U17494 (N_17494,N_17126,N_17087);
or U17495 (N_17495,N_17088,N_17105);
and U17496 (N_17496,N_17212,N_17089);
xor U17497 (N_17497,N_17084,N_17197);
nand U17498 (N_17498,N_17030,N_17115);
nor U17499 (N_17499,N_17185,N_17162);
and U17500 (N_17500,N_17290,N_17432);
and U17501 (N_17501,N_17262,N_17411);
xnor U17502 (N_17502,N_17369,N_17483);
and U17503 (N_17503,N_17257,N_17407);
and U17504 (N_17504,N_17429,N_17459);
and U17505 (N_17505,N_17345,N_17324);
nand U17506 (N_17506,N_17452,N_17457);
or U17507 (N_17507,N_17421,N_17269);
nor U17508 (N_17508,N_17492,N_17319);
or U17509 (N_17509,N_17335,N_17433);
nand U17510 (N_17510,N_17389,N_17448);
xor U17511 (N_17511,N_17293,N_17490);
or U17512 (N_17512,N_17347,N_17382);
and U17513 (N_17513,N_17456,N_17408);
xor U17514 (N_17514,N_17349,N_17258);
and U17515 (N_17515,N_17314,N_17463);
xor U17516 (N_17516,N_17405,N_17413);
nand U17517 (N_17517,N_17326,N_17286);
nor U17518 (N_17518,N_17487,N_17274);
nor U17519 (N_17519,N_17458,N_17395);
nor U17520 (N_17520,N_17361,N_17295);
xnor U17521 (N_17521,N_17303,N_17316);
nand U17522 (N_17522,N_17415,N_17283);
nor U17523 (N_17523,N_17343,N_17477);
and U17524 (N_17524,N_17467,N_17321);
xor U17525 (N_17525,N_17253,N_17461);
and U17526 (N_17526,N_17323,N_17251);
or U17527 (N_17527,N_17380,N_17439);
and U17528 (N_17528,N_17393,N_17489);
nand U17529 (N_17529,N_17400,N_17406);
nor U17530 (N_17530,N_17471,N_17265);
nor U17531 (N_17531,N_17270,N_17329);
or U17532 (N_17532,N_17437,N_17375);
nand U17533 (N_17533,N_17310,N_17351);
or U17534 (N_17534,N_17276,N_17252);
and U17535 (N_17535,N_17261,N_17430);
xnor U17536 (N_17536,N_17311,N_17266);
nand U17537 (N_17537,N_17312,N_17288);
or U17538 (N_17538,N_17379,N_17313);
and U17539 (N_17539,N_17453,N_17280);
nand U17540 (N_17540,N_17436,N_17256);
or U17541 (N_17541,N_17462,N_17255);
nor U17542 (N_17542,N_17447,N_17367);
nor U17543 (N_17543,N_17275,N_17428);
nand U17544 (N_17544,N_17254,N_17404);
and U17545 (N_17545,N_17300,N_17344);
nor U17546 (N_17546,N_17386,N_17480);
nor U17547 (N_17547,N_17473,N_17403);
xor U17548 (N_17548,N_17496,N_17353);
and U17549 (N_17549,N_17469,N_17260);
nor U17550 (N_17550,N_17373,N_17348);
and U17551 (N_17551,N_17376,N_17357);
xor U17552 (N_17552,N_17285,N_17449);
nor U17553 (N_17553,N_17416,N_17297);
nand U17554 (N_17554,N_17412,N_17294);
and U17555 (N_17555,N_17339,N_17468);
xnor U17556 (N_17556,N_17390,N_17277);
and U17557 (N_17557,N_17414,N_17498);
nor U17558 (N_17558,N_17338,N_17341);
and U17559 (N_17559,N_17332,N_17292);
xnor U17560 (N_17560,N_17360,N_17401);
nand U17561 (N_17561,N_17259,N_17278);
or U17562 (N_17562,N_17371,N_17250);
and U17563 (N_17563,N_17454,N_17442);
nor U17564 (N_17564,N_17464,N_17444);
or U17565 (N_17565,N_17315,N_17427);
nand U17566 (N_17566,N_17272,N_17486);
and U17567 (N_17567,N_17465,N_17419);
nand U17568 (N_17568,N_17359,N_17391);
xnor U17569 (N_17569,N_17482,N_17488);
and U17570 (N_17570,N_17481,N_17284);
nor U17571 (N_17571,N_17291,N_17306);
xnor U17572 (N_17572,N_17499,N_17476);
xnor U17573 (N_17573,N_17474,N_17495);
and U17574 (N_17574,N_17381,N_17478);
or U17575 (N_17575,N_17320,N_17308);
and U17576 (N_17576,N_17472,N_17460);
nand U17577 (N_17577,N_17438,N_17370);
nand U17578 (N_17578,N_17440,N_17346);
nand U17579 (N_17579,N_17368,N_17263);
nand U17580 (N_17580,N_17451,N_17420);
nand U17581 (N_17581,N_17383,N_17397);
or U17582 (N_17582,N_17470,N_17441);
and U17583 (N_17583,N_17322,N_17296);
and U17584 (N_17584,N_17385,N_17450);
and U17585 (N_17585,N_17378,N_17434);
and U17586 (N_17586,N_17366,N_17334);
xor U17587 (N_17587,N_17302,N_17299);
nor U17588 (N_17588,N_17350,N_17273);
nand U17589 (N_17589,N_17336,N_17364);
nand U17590 (N_17590,N_17325,N_17374);
xnor U17591 (N_17591,N_17363,N_17497);
nor U17592 (N_17592,N_17392,N_17445);
nor U17593 (N_17593,N_17491,N_17267);
and U17594 (N_17594,N_17402,N_17475);
or U17595 (N_17595,N_17356,N_17396);
nor U17596 (N_17596,N_17493,N_17384);
nor U17597 (N_17597,N_17282,N_17425);
or U17598 (N_17598,N_17443,N_17305);
and U17599 (N_17599,N_17355,N_17365);
or U17600 (N_17600,N_17318,N_17354);
and U17601 (N_17601,N_17387,N_17388);
and U17602 (N_17602,N_17317,N_17394);
xnor U17603 (N_17603,N_17281,N_17309);
xor U17604 (N_17604,N_17328,N_17304);
nand U17605 (N_17605,N_17307,N_17337);
or U17606 (N_17606,N_17327,N_17398);
nor U17607 (N_17607,N_17435,N_17431);
nand U17608 (N_17608,N_17377,N_17494);
xor U17609 (N_17609,N_17340,N_17418);
and U17610 (N_17610,N_17484,N_17298);
xor U17611 (N_17611,N_17333,N_17422);
xor U17612 (N_17612,N_17342,N_17268);
nor U17613 (N_17613,N_17446,N_17466);
xnor U17614 (N_17614,N_17485,N_17301);
or U17615 (N_17615,N_17289,N_17330);
nand U17616 (N_17616,N_17271,N_17423);
xnor U17617 (N_17617,N_17424,N_17426);
and U17618 (N_17618,N_17455,N_17372);
nand U17619 (N_17619,N_17358,N_17362);
nand U17620 (N_17620,N_17352,N_17264);
nand U17621 (N_17621,N_17399,N_17279);
nor U17622 (N_17622,N_17417,N_17331);
and U17623 (N_17623,N_17410,N_17479);
xnor U17624 (N_17624,N_17287,N_17409);
nor U17625 (N_17625,N_17362,N_17495);
nor U17626 (N_17626,N_17391,N_17332);
nand U17627 (N_17627,N_17440,N_17464);
nor U17628 (N_17628,N_17391,N_17470);
or U17629 (N_17629,N_17457,N_17470);
or U17630 (N_17630,N_17430,N_17333);
and U17631 (N_17631,N_17448,N_17459);
xnor U17632 (N_17632,N_17282,N_17452);
nor U17633 (N_17633,N_17479,N_17435);
nor U17634 (N_17634,N_17336,N_17368);
or U17635 (N_17635,N_17444,N_17411);
nor U17636 (N_17636,N_17401,N_17421);
xnor U17637 (N_17637,N_17326,N_17342);
and U17638 (N_17638,N_17392,N_17394);
or U17639 (N_17639,N_17449,N_17335);
xnor U17640 (N_17640,N_17340,N_17389);
and U17641 (N_17641,N_17492,N_17305);
nand U17642 (N_17642,N_17259,N_17424);
or U17643 (N_17643,N_17340,N_17343);
and U17644 (N_17644,N_17478,N_17324);
and U17645 (N_17645,N_17452,N_17267);
nor U17646 (N_17646,N_17282,N_17434);
xor U17647 (N_17647,N_17370,N_17338);
xnor U17648 (N_17648,N_17449,N_17460);
and U17649 (N_17649,N_17262,N_17285);
nor U17650 (N_17650,N_17294,N_17320);
or U17651 (N_17651,N_17454,N_17487);
and U17652 (N_17652,N_17387,N_17348);
and U17653 (N_17653,N_17296,N_17295);
nand U17654 (N_17654,N_17306,N_17267);
xor U17655 (N_17655,N_17351,N_17334);
and U17656 (N_17656,N_17413,N_17437);
nor U17657 (N_17657,N_17306,N_17444);
or U17658 (N_17658,N_17306,N_17473);
xor U17659 (N_17659,N_17277,N_17496);
or U17660 (N_17660,N_17441,N_17264);
nand U17661 (N_17661,N_17424,N_17317);
or U17662 (N_17662,N_17381,N_17473);
nand U17663 (N_17663,N_17323,N_17333);
nor U17664 (N_17664,N_17424,N_17326);
nor U17665 (N_17665,N_17394,N_17292);
nor U17666 (N_17666,N_17485,N_17491);
nand U17667 (N_17667,N_17408,N_17272);
xor U17668 (N_17668,N_17485,N_17252);
and U17669 (N_17669,N_17277,N_17484);
or U17670 (N_17670,N_17385,N_17374);
nor U17671 (N_17671,N_17341,N_17442);
and U17672 (N_17672,N_17405,N_17356);
and U17673 (N_17673,N_17380,N_17267);
nor U17674 (N_17674,N_17382,N_17360);
nor U17675 (N_17675,N_17333,N_17479);
xnor U17676 (N_17676,N_17385,N_17272);
xnor U17677 (N_17677,N_17263,N_17387);
nand U17678 (N_17678,N_17305,N_17379);
nor U17679 (N_17679,N_17355,N_17349);
and U17680 (N_17680,N_17323,N_17492);
and U17681 (N_17681,N_17422,N_17335);
nor U17682 (N_17682,N_17391,N_17285);
nand U17683 (N_17683,N_17378,N_17427);
and U17684 (N_17684,N_17268,N_17332);
nand U17685 (N_17685,N_17430,N_17470);
and U17686 (N_17686,N_17459,N_17471);
xnor U17687 (N_17687,N_17354,N_17405);
or U17688 (N_17688,N_17459,N_17300);
xor U17689 (N_17689,N_17365,N_17490);
xnor U17690 (N_17690,N_17269,N_17365);
nor U17691 (N_17691,N_17492,N_17449);
xnor U17692 (N_17692,N_17346,N_17457);
xnor U17693 (N_17693,N_17300,N_17263);
xor U17694 (N_17694,N_17452,N_17360);
and U17695 (N_17695,N_17324,N_17465);
and U17696 (N_17696,N_17365,N_17398);
and U17697 (N_17697,N_17388,N_17375);
nand U17698 (N_17698,N_17376,N_17322);
and U17699 (N_17699,N_17470,N_17397);
xnor U17700 (N_17700,N_17268,N_17482);
nand U17701 (N_17701,N_17398,N_17453);
or U17702 (N_17702,N_17283,N_17282);
or U17703 (N_17703,N_17351,N_17460);
or U17704 (N_17704,N_17483,N_17385);
nand U17705 (N_17705,N_17314,N_17468);
and U17706 (N_17706,N_17394,N_17393);
or U17707 (N_17707,N_17410,N_17420);
nand U17708 (N_17708,N_17310,N_17259);
or U17709 (N_17709,N_17314,N_17333);
xor U17710 (N_17710,N_17333,N_17296);
or U17711 (N_17711,N_17251,N_17334);
xor U17712 (N_17712,N_17381,N_17385);
or U17713 (N_17713,N_17445,N_17331);
and U17714 (N_17714,N_17464,N_17330);
nand U17715 (N_17715,N_17384,N_17318);
xor U17716 (N_17716,N_17397,N_17497);
and U17717 (N_17717,N_17493,N_17400);
xnor U17718 (N_17718,N_17428,N_17255);
xnor U17719 (N_17719,N_17267,N_17354);
or U17720 (N_17720,N_17403,N_17426);
nor U17721 (N_17721,N_17278,N_17481);
and U17722 (N_17722,N_17314,N_17286);
xor U17723 (N_17723,N_17496,N_17359);
xor U17724 (N_17724,N_17482,N_17351);
nand U17725 (N_17725,N_17439,N_17390);
nor U17726 (N_17726,N_17499,N_17355);
nand U17727 (N_17727,N_17421,N_17469);
nand U17728 (N_17728,N_17291,N_17444);
xnor U17729 (N_17729,N_17259,N_17298);
nor U17730 (N_17730,N_17462,N_17253);
or U17731 (N_17731,N_17347,N_17258);
or U17732 (N_17732,N_17388,N_17477);
and U17733 (N_17733,N_17450,N_17267);
xor U17734 (N_17734,N_17298,N_17275);
nor U17735 (N_17735,N_17354,N_17307);
or U17736 (N_17736,N_17357,N_17432);
nand U17737 (N_17737,N_17332,N_17314);
nor U17738 (N_17738,N_17322,N_17483);
nand U17739 (N_17739,N_17397,N_17439);
and U17740 (N_17740,N_17289,N_17451);
nand U17741 (N_17741,N_17410,N_17320);
or U17742 (N_17742,N_17261,N_17313);
or U17743 (N_17743,N_17349,N_17262);
or U17744 (N_17744,N_17483,N_17261);
and U17745 (N_17745,N_17326,N_17482);
nor U17746 (N_17746,N_17466,N_17350);
nor U17747 (N_17747,N_17303,N_17343);
or U17748 (N_17748,N_17451,N_17262);
and U17749 (N_17749,N_17332,N_17446);
nor U17750 (N_17750,N_17743,N_17538);
xor U17751 (N_17751,N_17584,N_17547);
nor U17752 (N_17752,N_17651,N_17719);
nand U17753 (N_17753,N_17625,N_17532);
and U17754 (N_17754,N_17586,N_17745);
or U17755 (N_17755,N_17548,N_17685);
nor U17756 (N_17756,N_17506,N_17623);
xor U17757 (N_17757,N_17659,N_17711);
xnor U17758 (N_17758,N_17555,N_17663);
nand U17759 (N_17759,N_17724,N_17701);
xnor U17760 (N_17760,N_17527,N_17560);
or U17761 (N_17761,N_17733,N_17604);
xor U17762 (N_17762,N_17723,N_17702);
or U17763 (N_17763,N_17686,N_17741);
and U17764 (N_17764,N_17660,N_17666);
and U17765 (N_17765,N_17540,N_17704);
and U17766 (N_17766,N_17605,N_17742);
nand U17767 (N_17767,N_17646,N_17630);
xor U17768 (N_17768,N_17622,N_17603);
and U17769 (N_17769,N_17717,N_17706);
xnor U17770 (N_17770,N_17677,N_17594);
and U17771 (N_17771,N_17599,N_17728);
nor U17772 (N_17772,N_17620,N_17730);
nand U17773 (N_17773,N_17601,N_17597);
nand U17774 (N_17774,N_17649,N_17636);
nand U17775 (N_17775,N_17600,N_17580);
nor U17776 (N_17776,N_17746,N_17674);
xor U17777 (N_17777,N_17669,N_17641);
nand U17778 (N_17778,N_17579,N_17612);
nor U17779 (N_17779,N_17713,N_17558);
and U17780 (N_17780,N_17526,N_17645);
or U17781 (N_17781,N_17740,N_17553);
nor U17782 (N_17782,N_17696,N_17567);
xnor U17783 (N_17783,N_17593,N_17566);
nor U17784 (N_17784,N_17682,N_17517);
xor U17785 (N_17785,N_17528,N_17609);
and U17786 (N_17786,N_17697,N_17661);
xnor U17787 (N_17787,N_17722,N_17716);
nor U17788 (N_17788,N_17672,N_17511);
nor U17789 (N_17789,N_17546,N_17652);
nand U17790 (N_17790,N_17520,N_17680);
nand U17791 (N_17791,N_17590,N_17735);
or U17792 (N_17792,N_17631,N_17638);
and U17793 (N_17793,N_17705,N_17541);
xnor U17794 (N_17794,N_17642,N_17549);
xor U17795 (N_17795,N_17545,N_17725);
nor U17796 (N_17796,N_17658,N_17667);
xnor U17797 (N_17797,N_17739,N_17662);
nand U17798 (N_17798,N_17691,N_17633);
and U17799 (N_17799,N_17731,N_17512);
and U17800 (N_17800,N_17562,N_17681);
nor U17801 (N_17801,N_17703,N_17515);
nand U17802 (N_17802,N_17665,N_17618);
nor U17803 (N_17803,N_17679,N_17554);
nor U17804 (N_17804,N_17587,N_17644);
or U17805 (N_17805,N_17726,N_17727);
nand U17806 (N_17806,N_17570,N_17577);
and U17807 (N_17807,N_17699,N_17718);
xor U17808 (N_17808,N_17664,N_17502);
nand U17809 (N_17809,N_17606,N_17748);
or U17810 (N_17810,N_17683,N_17708);
and U17811 (N_17811,N_17583,N_17559);
xor U17812 (N_17812,N_17694,N_17585);
nor U17813 (N_17813,N_17564,N_17617);
nand U17814 (N_17814,N_17614,N_17531);
and U17815 (N_17815,N_17533,N_17589);
nand U17816 (N_17816,N_17714,N_17670);
and U17817 (N_17817,N_17552,N_17653);
nand U17818 (N_17818,N_17539,N_17550);
xnor U17819 (N_17819,N_17556,N_17536);
or U17820 (N_17820,N_17687,N_17615);
xor U17821 (N_17821,N_17624,N_17616);
or U17822 (N_17822,N_17632,N_17721);
nand U17823 (N_17823,N_17734,N_17707);
xor U17824 (N_17824,N_17571,N_17688);
nand U17825 (N_17825,N_17598,N_17525);
nand U17826 (N_17826,N_17693,N_17690);
xnor U17827 (N_17827,N_17607,N_17563);
xor U17828 (N_17828,N_17516,N_17640);
and U17829 (N_17829,N_17578,N_17700);
xor U17830 (N_17830,N_17534,N_17749);
and U17831 (N_17831,N_17504,N_17709);
nor U17832 (N_17832,N_17529,N_17509);
nand U17833 (N_17833,N_17592,N_17648);
xor U17834 (N_17834,N_17543,N_17572);
and U17835 (N_17835,N_17710,N_17507);
nand U17836 (N_17836,N_17637,N_17573);
nand U17837 (N_17837,N_17581,N_17591);
nor U17838 (N_17838,N_17565,N_17519);
nor U17839 (N_17839,N_17574,N_17576);
nand U17840 (N_17840,N_17675,N_17602);
and U17841 (N_17841,N_17508,N_17684);
nor U17842 (N_17842,N_17582,N_17628);
and U17843 (N_17843,N_17561,N_17732);
nor U17844 (N_17844,N_17535,N_17657);
xnor U17845 (N_17845,N_17650,N_17627);
xnor U17846 (N_17846,N_17501,N_17613);
xnor U17847 (N_17847,N_17569,N_17629);
or U17848 (N_17848,N_17720,N_17595);
nand U17849 (N_17849,N_17671,N_17514);
or U17850 (N_17850,N_17518,N_17524);
or U17851 (N_17851,N_17712,N_17626);
or U17852 (N_17852,N_17634,N_17737);
nand U17853 (N_17853,N_17715,N_17611);
nand U17854 (N_17854,N_17510,N_17744);
and U17855 (N_17855,N_17736,N_17656);
and U17856 (N_17856,N_17542,N_17557);
nand U17857 (N_17857,N_17676,N_17692);
nand U17858 (N_17858,N_17503,N_17695);
xor U17859 (N_17859,N_17568,N_17505);
or U17860 (N_17860,N_17647,N_17521);
nand U17861 (N_17861,N_17654,N_17530);
nand U17862 (N_17862,N_17621,N_17523);
xor U17863 (N_17863,N_17619,N_17678);
nor U17864 (N_17864,N_17738,N_17689);
or U17865 (N_17865,N_17610,N_17639);
xor U17866 (N_17866,N_17729,N_17668);
nor U17867 (N_17867,N_17522,N_17537);
and U17868 (N_17868,N_17588,N_17655);
xor U17869 (N_17869,N_17643,N_17513);
nand U17870 (N_17870,N_17500,N_17673);
xnor U17871 (N_17871,N_17596,N_17544);
and U17872 (N_17872,N_17747,N_17608);
and U17873 (N_17873,N_17635,N_17698);
or U17874 (N_17874,N_17551,N_17575);
nor U17875 (N_17875,N_17609,N_17624);
and U17876 (N_17876,N_17505,N_17726);
xor U17877 (N_17877,N_17523,N_17700);
and U17878 (N_17878,N_17687,N_17717);
nor U17879 (N_17879,N_17626,N_17695);
nand U17880 (N_17880,N_17702,N_17593);
or U17881 (N_17881,N_17678,N_17613);
and U17882 (N_17882,N_17704,N_17710);
and U17883 (N_17883,N_17611,N_17528);
nand U17884 (N_17884,N_17652,N_17574);
nand U17885 (N_17885,N_17543,N_17696);
and U17886 (N_17886,N_17593,N_17518);
nand U17887 (N_17887,N_17627,N_17601);
and U17888 (N_17888,N_17653,N_17642);
nand U17889 (N_17889,N_17535,N_17599);
xor U17890 (N_17890,N_17690,N_17530);
xor U17891 (N_17891,N_17588,N_17594);
nor U17892 (N_17892,N_17545,N_17542);
nor U17893 (N_17893,N_17726,N_17554);
xnor U17894 (N_17894,N_17662,N_17688);
nor U17895 (N_17895,N_17638,N_17651);
xnor U17896 (N_17896,N_17578,N_17692);
or U17897 (N_17897,N_17566,N_17731);
nand U17898 (N_17898,N_17580,N_17503);
nand U17899 (N_17899,N_17512,N_17667);
nand U17900 (N_17900,N_17502,N_17622);
nand U17901 (N_17901,N_17670,N_17747);
nor U17902 (N_17902,N_17653,N_17596);
nand U17903 (N_17903,N_17677,N_17667);
or U17904 (N_17904,N_17731,N_17730);
nand U17905 (N_17905,N_17692,N_17517);
nand U17906 (N_17906,N_17546,N_17627);
nor U17907 (N_17907,N_17650,N_17633);
and U17908 (N_17908,N_17598,N_17740);
xor U17909 (N_17909,N_17511,N_17592);
nand U17910 (N_17910,N_17543,N_17518);
nor U17911 (N_17911,N_17545,N_17625);
nand U17912 (N_17912,N_17567,N_17662);
and U17913 (N_17913,N_17544,N_17636);
nand U17914 (N_17914,N_17538,N_17534);
or U17915 (N_17915,N_17741,N_17557);
nor U17916 (N_17916,N_17589,N_17619);
xor U17917 (N_17917,N_17594,N_17671);
xor U17918 (N_17918,N_17583,N_17664);
or U17919 (N_17919,N_17528,N_17516);
and U17920 (N_17920,N_17706,N_17672);
nor U17921 (N_17921,N_17506,N_17707);
and U17922 (N_17922,N_17555,N_17679);
nand U17923 (N_17923,N_17586,N_17723);
or U17924 (N_17924,N_17652,N_17672);
nand U17925 (N_17925,N_17662,N_17566);
nand U17926 (N_17926,N_17748,N_17515);
and U17927 (N_17927,N_17547,N_17594);
and U17928 (N_17928,N_17636,N_17613);
xnor U17929 (N_17929,N_17709,N_17621);
nor U17930 (N_17930,N_17524,N_17680);
nor U17931 (N_17931,N_17516,N_17707);
and U17932 (N_17932,N_17735,N_17728);
and U17933 (N_17933,N_17613,N_17553);
nor U17934 (N_17934,N_17515,N_17650);
xnor U17935 (N_17935,N_17615,N_17612);
nand U17936 (N_17936,N_17600,N_17513);
nand U17937 (N_17937,N_17525,N_17587);
nor U17938 (N_17938,N_17650,N_17537);
and U17939 (N_17939,N_17648,N_17657);
nor U17940 (N_17940,N_17734,N_17693);
and U17941 (N_17941,N_17656,N_17569);
or U17942 (N_17942,N_17531,N_17526);
nand U17943 (N_17943,N_17621,N_17596);
xor U17944 (N_17944,N_17722,N_17637);
nor U17945 (N_17945,N_17676,N_17701);
xor U17946 (N_17946,N_17604,N_17744);
nand U17947 (N_17947,N_17688,N_17501);
xor U17948 (N_17948,N_17546,N_17539);
nand U17949 (N_17949,N_17567,N_17611);
nor U17950 (N_17950,N_17734,N_17538);
or U17951 (N_17951,N_17603,N_17687);
or U17952 (N_17952,N_17576,N_17666);
or U17953 (N_17953,N_17513,N_17610);
xnor U17954 (N_17954,N_17680,N_17725);
xor U17955 (N_17955,N_17558,N_17740);
nor U17956 (N_17956,N_17746,N_17683);
xor U17957 (N_17957,N_17600,N_17680);
nor U17958 (N_17958,N_17695,N_17600);
or U17959 (N_17959,N_17707,N_17624);
xor U17960 (N_17960,N_17699,N_17666);
nor U17961 (N_17961,N_17637,N_17543);
and U17962 (N_17962,N_17698,N_17506);
nand U17963 (N_17963,N_17579,N_17560);
and U17964 (N_17964,N_17697,N_17618);
nor U17965 (N_17965,N_17675,N_17679);
nor U17966 (N_17966,N_17737,N_17673);
xnor U17967 (N_17967,N_17690,N_17617);
nor U17968 (N_17968,N_17612,N_17628);
nor U17969 (N_17969,N_17678,N_17531);
nand U17970 (N_17970,N_17502,N_17562);
and U17971 (N_17971,N_17733,N_17728);
or U17972 (N_17972,N_17646,N_17741);
and U17973 (N_17973,N_17611,N_17719);
nand U17974 (N_17974,N_17675,N_17537);
nor U17975 (N_17975,N_17615,N_17679);
and U17976 (N_17976,N_17632,N_17581);
xnor U17977 (N_17977,N_17534,N_17630);
xor U17978 (N_17978,N_17520,N_17589);
nor U17979 (N_17979,N_17651,N_17542);
and U17980 (N_17980,N_17749,N_17503);
nand U17981 (N_17981,N_17641,N_17569);
xnor U17982 (N_17982,N_17516,N_17501);
nand U17983 (N_17983,N_17535,N_17624);
and U17984 (N_17984,N_17627,N_17726);
xnor U17985 (N_17985,N_17746,N_17542);
nand U17986 (N_17986,N_17683,N_17543);
nand U17987 (N_17987,N_17607,N_17595);
nand U17988 (N_17988,N_17579,N_17573);
xnor U17989 (N_17989,N_17572,N_17599);
xnor U17990 (N_17990,N_17516,N_17614);
or U17991 (N_17991,N_17680,N_17503);
nand U17992 (N_17992,N_17580,N_17746);
nor U17993 (N_17993,N_17581,N_17534);
nand U17994 (N_17994,N_17675,N_17628);
nand U17995 (N_17995,N_17690,N_17710);
and U17996 (N_17996,N_17638,N_17600);
or U17997 (N_17997,N_17530,N_17737);
xor U17998 (N_17998,N_17742,N_17636);
or U17999 (N_17999,N_17686,N_17629);
nor U18000 (N_18000,N_17955,N_17839);
xnor U18001 (N_18001,N_17935,N_17929);
and U18002 (N_18002,N_17848,N_17964);
and U18003 (N_18003,N_17825,N_17814);
nand U18004 (N_18004,N_17798,N_17902);
or U18005 (N_18005,N_17898,N_17841);
and U18006 (N_18006,N_17918,N_17916);
and U18007 (N_18007,N_17943,N_17768);
or U18008 (N_18008,N_17996,N_17756);
xnor U18009 (N_18009,N_17881,N_17767);
xnor U18010 (N_18010,N_17805,N_17844);
and U18011 (N_18011,N_17921,N_17928);
and U18012 (N_18012,N_17857,N_17930);
xnor U18013 (N_18013,N_17905,N_17887);
nand U18014 (N_18014,N_17873,N_17884);
xor U18015 (N_18015,N_17937,N_17801);
nand U18016 (N_18016,N_17947,N_17961);
nor U18017 (N_18017,N_17770,N_17863);
and U18018 (N_18018,N_17903,N_17799);
nor U18019 (N_18019,N_17836,N_17892);
and U18020 (N_18020,N_17972,N_17757);
or U18021 (N_18021,N_17861,N_17885);
and U18022 (N_18022,N_17752,N_17904);
or U18023 (N_18023,N_17753,N_17993);
nand U18024 (N_18024,N_17758,N_17889);
and U18025 (N_18025,N_17842,N_17851);
xnor U18026 (N_18026,N_17870,N_17965);
or U18027 (N_18027,N_17948,N_17899);
nor U18028 (N_18028,N_17975,N_17837);
xor U18029 (N_18029,N_17969,N_17938);
xnor U18030 (N_18030,N_17872,N_17761);
or U18031 (N_18031,N_17776,N_17963);
xnor U18032 (N_18032,N_17786,N_17764);
and U18033 (N_18033,N_17787,N_17858);
xor U18034 (N_18034,N_17990,N_17946);
xor U18035 (N_18035,N_17894,N_17852);
nand U18036 (N_18036,N_17981,N_17920);
and U18037 (N_18037,N_17924,N_17931);
xor U18038 (N_18038,N_17925,N_17869);
nand U18039 (N_18039,N_17833,N_17973);
xor U18040 (N_18040,N_17914,N_17783);
or U18041 (N_18041,N_17883,N_17769);
or U18042 (N_18042,N_17960,N_17818);
xor U18043 (N_18043,N_17777,N_17877);
and U18044 (N_18044,N_17835,N_17806);
nor U18045 (N_18045,N_17775,N_17967);
or U18046 (N_18046,N_17803,N_17911);
nor U18047 (N_18047,N_17901,N_17941);
xor U18048 (N_18048,N_17763,N_17840);
and U18049 (N_18049,N_17890,N_17774);
nand U18050 (N_18050,N_17979,N_17838);
nor U18051 (N_18051,N_17864,N_17826);
and U18052 (N_18052,N_17797,N_17988);
xor U18053 (N_18053,N_17765,N_17847);
nor U18054 (N_18054,N_17942,N_17790);
nand U18055 (N_18055,N_17810,N_17895);
and U18056 (N_18056,N_17880,N_17891);
xor U18057 (N_18057,N_17945,N_17773);
xnor U18058 (N_18058,N_17912,N_17854);
and U18059 (N_18059,N_17772,N_17794);
and U18060 (N_18060,N_17927,N_17951);
nand U18061 (N_18061,N_17860,N_17866);
xnor U18062 (N_18062,N_17940,N_17750);
xor U18063 (N_18063,N_17865,N_17817);
and U18064 (N_18064,N_17781,N_17762);
nand U18065 (N_18065,N_17816,N_17754);
nand U18066 (N_18066,N_17824,N_17791);
xor U18067 (N_18067,N_17952,N_17856);
and U18068 (N_18068,N_17954,N_17959);
or U18069 (N_18069,N_17813,N_17867);
xor U18070 (N_18070,N_17811,N_17808);
nand U18071 (N_18071,N_17915,N_17828);
nand U18072 (N_18072,N_17874,N_17888);
xor U18073 (N_18073,N_17751,N_17909);
and U18074 (N_18074,N_17886,N_17819);
nor U18075 (N_18075,N_17986,N_17917);
nand U18076 (N_18076,N_17843,N_17980);
xnor U18077 (N_18077,N_17815,N_17800);
xor U18078 (N_18078,N_17875,N_17983);
and U18079 (N_18079,N_17859,N_17862);
nor U18080 (N_18080,N_17976,N_17778);
nor U18081 (N_18081,N_17760,N_17907);
nand U18082 (N_18082,N_17995,N_17792);
nor U18083 (N_18083,N_17987,N_17936);
or U18084 (N_18084,N_17893,N_17900);
nor U18085 (N_18085,N_17850,N_17823);
or U18086 (N_18086,N_17793,N_17958);
nand U18087 (N_18087,N_17923,N_17978);
nand U18088 (N_18088,N_17785,N_17849);
and U18089 (N_18089,N_17932,N_17796);
or U18090 (N_18090,N_17804,N_17998);
xor U18091 (N_18091,N_17896,N_17919);
and U18092 (N_18092,N_17782,N_17974);
and U18093 (N_18093,N_17910,N_17977);
and U18094 (N_18094,N_17789,N_17784);
nand U18095 (N_18095,N_17812,N_17984);
nand U18096 (N_18096,N_17966,N_17871);
nor U18097 (N_18097,N_17962,N_17985);
xnor U18098 (N_18098,N_17829,N_17795);
or U18099 (N_18099,N_17939,N_17876);
xnor U18100 (N_18100,N_17831,N_17970);
xnor U18101 (N_18101,N_17832,N_17771);
nand U18102 (N_18102,N_17822,N_17950);
xnor U18103 (N_18103,N_17934,N_17991);
and U18104 (N_18104,N_17997,N_17830);
nand U18105 (N_18105,N_17882,N_17992);
nand U18106 (N_18106,N_17913,N_17944);
or U18107 (N_18107,N_17999,N_17827);
or U18108 (N_18108,N_17834,N_17759);
nor U18109 (N_18109,N_17846,N_17855);
nor U18110 (N_18110,N_17788,N_17908);
xor U18111 (N_18111,N_17971,N_17821);
nand U18112 (N_18112,N_17897,N_17802);
and U18113 (N_18113,N_17779,N_17820);
nor U18114 (N_18114,N_17982,N_17989);
or U18115 (N_18115,N_17755,N_17949);
nor U18116 (N_18116,N_17807,N_17853);
nor U18117 (N_18117,N_17922,N_17879);
xor U18118 (N_18118,N_17953,N_17780);
or U18119 (N_18119,N_17933,N_17845);
and U18120 (N_18120,N_17926,N_17957);
nand U18121 (N_18121,N_17956,N_17766);
or U18122 (N_18122,N_17809,N_17868);
nor U18123 (N_18123,N_17878,N_17994);
and U18124 (N_18124,N_17968,N_17906);
nor U18125 (N_18125,N_17885,N_17977);
or U18126 (N_18126,N_17998,N_17951);
or U18127 (N_18127,N_17824,N_17828);
and U18128 (N_18128,N_17990,N_17897);
and U18129 (N_18129,N_17875,N_17985);
or U18130 (N_18130,N_17960,N_17951);
xor U18131 (N_18131,N_17871,N_17878);
xor U18132 (N_18132,N_17964,N_17821);
nand U18133 (N_18133,N_17772,N_17951);
or U18134 (N_18134,N_17795,N_17836);
nand U18135 (N_18135,N_17771,N_17755);
nor U18136 (N_18136,N_17853,N_17931);
or U18137 (N_18137,N_17765,N_17974);
nor U18138 (N_18138,N_17854,N_17920);
xor U18139 (N_18139,N_17974,N_17764);
and U18140 (N_18140,N_17942,N_17923);
nor U18141 (N_18141,N_17811,N_17776);
or U18142 (N_18142,N_17918,N_17846);
nor U18143 (N_18143,N_17842,N_17808);
or U18144 (N_18144,N_17807,N_17841);
or U18145 (N_18145,N_17945,N_17990);
nand U18146 (N_18146,N_17895,N_17764);
nor U18147 (N_18147,N_17795,N_17924);
and U18148 (N_18148,N_17880,N_17824);
nand U18149 (N_18149,N_17821,N_17937);
xor U18150 (N_18150,N_17753,N_17964);
nand U18151 (N_18151,N_17822,N_17977);
nand U18152 (N_18152,N_17794,N_17807);
and U18153 (N_18153,N_17868,N_17893);
or U18154 (N_18154,N_17878,N_17923);
xnor U18155 (N_18155,N_17792,N_17779);
or U18156 (N_18156,N_17934,N_17965);
and U18157 (N_18157,N_17936,N_17898);
xnor U18158 (N_18158,N_17957,N_17946);
or U18159 (N_18159,N_17885,N_17958);
or U18160 (N_18160,N_17978,N_17938);
nor U18161 (N_18161,N_17953,N_17815);
nand U18162 (N_18162,N_17813,N_17864);
and U18163 (N_18163,N_17936,N_17780);
nand U18164 (N_18164,N_17988,N_17777);
nor U18165 (N_18165,N_17816,N_17945);
and U18166 (N_18166,N_17800,N_17998);
or U18167 (N_18167,N_17963,N_17910);
nor U18168 (N_18168,N_17946,N_17998);
and U18169 (N_18169,N_17864,N_17940);
nor U18170 (N_18170,N_17822,N_17908);
nor U18171 (N_18171,N_17962,N_17855);
nor U18172 (N_18172,N_17884,N_17971);
nand U18173 (N_18173,N_17866,N_17922);
and U18174 (N_18174,N_17852,N_17984);
nand U18175 (N_18175,N_17898,N_17991);
or U18176 (N_18176,N_17883,N_17972);
nor U18177 (N_18177,N_17833,N_17971);
and U18178 (N_18178,N_17883,N_17807);
xnor U18179 (N_18179,N_17909,N_17919);
nor U18180 (N_18180,N_17980,N_17938);
and U18181 (N_18181,N_17777,N_17805);
xor U18182 (N_18182,N_17977,N_17965);
nand U18183 (N_18183,N_17790,N_17766);
xor U18184 (N_18184,N_17906,N_17837);
nor U18185 (N_18185,N_17955,N_17996);
nand U18186 (N_18186,N_17970,N_17833);
and U18187 (N_18187,N_17969,N_17935);
or U18188 (N_18188,N_17821,N_17768);
and U18189 (N_18189,N_17943,N_17859);
nand U18190 (N_18190,N_17929,N_17989);
nor U18191 (N_18191,N_17773,N_17856);
or U18192 (N_18192,N_17942,N_17780);
and U18193 (N_18193,N_17832,N_17886);
nor U18194 (N_18194,N_17900,N_17906);
or U18195 (N_18195,N_17988,N_17782);
or U18196 (N_18196,N_17811,N_17861);
or U18197 (N_18197,N_17958,N_17859);
xnor U18198 (N_18198,N_17861,N_17993);
nor U18199 (N_18199,N_17935,N_17759);
or U18200 (N_18200,N_17926,N_17962);
nand U18201 (N_18201,N_17877,N_17832);
nor U18202 (N_18202,N_17750,N_17853);
nand U18203 (N_18203,N_17952,N_17886);
nor U18204 (N_18204,N_17843,N_17767);
nand U18205 (N_18205,N_17826,N_17989);
nor U18206 (N_18206,N_17810,N_17912);
or U18207 (N_18207,N_17956,N_17855);
and U18208 (N_18208,N_17909,N_17797);
and U18209 (N_18209,N_17769,N_17753);
xor U18210 (N_18210,N_17814,N_17834);
nor U18211 (N_18211,N_17995,N_17938);
nor U18212 (N_18212,N_17838,N_17758);
nand U18213 (N_18213,N_17890,N_17814);
or U18214 (N_18214,N_17982,N_17873);
and U18215 (N_18215,N_17969,N_17763);
nor U18216 (N_18216,N_17817,N_17919);
xnor U18217 (N_18217,N_17994,N_17899);
or U18218 (N_18218,N_17835,N_17938);
or U18219 (N_18219,N_17774,N_17871);
xor U18220 (N_18220,N_17833,N_17923);
and U18221 (N_18221,N_17863,N_17887);
xnor U18222 (N_18222,N_17870,N_17950);
nor U18223 (N_18223,N_17869,N_17842);
nor U18224 (N_18224,N_17932,N_17989);
nor U18225 (N_18225,N_17855,N_17889);
xnor U18226 (N_18226,N_17789,N_17838);
nand U18227 (N_18227,N_17821,N_17878);
and U18228 (N_18228,N_17922,N_17932);
nand U18229 (N_18229,N_17752,N_17864);
nor U18230 (N_18230,N_17773,N_17783);
nand U18231 (N_18231,N_17797,N_17921);
or U18232 (N_18232,N_17782,N_17836);
xnor U18233 (N_18233,N_17751,N_17888);
nand U18234 (N_18234,N_17940,N_17947);
xnor U18235 (N_18235,N_17966,N_17944);
and U18236 (N_18236,N_17962,N_17889);
xor U18237 (N_18237,N_17789,N_17943);
and U18238 (N_18238,N_17956,N_17808);
nand U18239 (N_18239,N_17801,N_17945);
nor U18240 (N_18240,N_17898,N_17974);
or U18241 (N_18241,N_17755,N_17822);
nand U18242 (N_18242,N_17754,N_17766);
nand U18243 (N_18243,N_17989,N_17888);
nor U18244 (N_18244,N_17974,N_17902);
nor U18245 (N_18245,N_17785,N_17951);
and U18246 (N_18246,N_17931,N_17769);
nand U18247 (N_18247,N_17955,N_17779);
nand U18248 (N_18248,N_17795,N_17886);
nand U18249 (N_18249,N_17981,N_17864);
nand U18250 (N_18250,N_18210,N_18027);
or U18251 (N_18251,N_18214,N_18238);
xnor U18252 (N_18252,N_18201,N_18002);
nor U18253 (N_18253,N_18096,N_18036);
or U18254 (N_18254,N_18092,N_18045);
and U18255 (N_18255,N_18160,N_18145);
nand U18256 (N_18256,N_18159,N_18018);
nand U18257 (N_18257,N_18161,N_18222);
nand U18258 (N_18258,N_18121,N_18011);
nand U18259 (N_18259,N_18231,N_18078);
nor U18260 (N_18260,N_18111,N_18125);
or U18261 (N_18261,N_18043,N_18024);
or U18262 (N_18262,N_18044,N_18213);
or U18263 (N_18263,N_18193,N_18206);
nand U18264 (N_18264,N_18170,N_18131);
xor U18265 (N_18265,N_18156,N_18042);
and U18266 (N_18266,N_18243,N_18164);
nor U18267 (N_18267,N_18003,N_18079);
or U18268 (N_18268,N_18012,N_18211);
xnor U18269 (N_18269,N_18028,N_18008);
nor U18270 (N_18270,N_18120,N_18014);
nand U18271 (N_18271,N_18127,N_18144);
nor U18272 (N_18272,N_18181,N_18200);
nand U18273 (N_18273,N_18004,N_18103);
and U18274 (N_18274,N_18182,N_18130);
xnor U18275 (N_18275,N_18038,N_18034);
nor U18276 (N_18276,N_18188,N_18098);
xor U18277 (N_18277,N_18245,N_18082);
and U18278 (N_18278,N_18172,N_18063);
nand U18279 (N_18279,N_18219,N_18007);
and U18280 (N_18280,N_18239,N_18178);
nand U18281 (N_18281,N_18023,N_18029);
nand U18282 (N_18282,N_18077,N_18021);
nor U18283 (N_18283,N_18039,N_18241);
and U18284 (N_18284,N_18185,N_18197);
nor U18285 (N_18285,N_18019,N_18115);
nand U18286 (N_18286,N_18208,N_18060);
nand U18287 (N_18287,N_18132,N_18179);
and U18288 (N_18288,N_18158,N_18207);
nand U18289 (N_18289,N_18061,N_18083);
xnor U18290 (N_18290,N_18069,N_18101);
xnor U18291 (N_18291,N_18032,N_18064);
nor U18292 (N_18292,N_18009,N_18123);
or U18293 (N_18293,N_18220,N_18124);
and U18294 (N_18294,N_18076,N_18129);
or U18295 (N_18295,N_18177,N_18048);
and U18296 (N_18296,N_18141,N_18062);
nand U18297 (N_18297,N_18015,N_18110);
and U18298 (N_18298,N_18106,N_18091);
xor U18299 (N_18299,N_18112,N_18246);
nand U18300 (N_18300,N_18215,N_18237);
xnor U18301 (N_18301,N_18035,N_18081);
or U18302 (N_18302,N_18074,N_18031);
or U18303 (N_18303,N_18051,N_18068);
and U18304 (N_18304,N_18094,N_18232);
xor U18305 (N_18305,N_18190,N_18025);
nor U18306 (N_18306,N_18148,N_18065);
xor U18307 (N_18307,N_18105,N_18244);
xor U18308 (N_18308,N_18166,N_18040);
xor U18309 (N_18309,N_18191,N_18187);
and U18310 (N_18310,N_18057,N_18234);
xnor U18311 (N_18311,N_18154,N_18117);
xnor U18312 (N_18312,N_18113,N_18216);
nor U18313 (N_18313,N_18198,N_18122);
or U18314 (N_18314,N_18173,N_18095);
xnor U18315 (N_18315,N_18137,N_18058);
or U18316 (N_18316,N_18202,N_18087);
or U18317 (N_18317,N_18041,N_18054);
xnor U18318 (N_18318,N_18189,N_18152);
nor U18319 (N_18319,N_18184,N_18176);
and U18320 (N_18320,N_18134,N_18247);
xor U18321 (N_18321,N_18142,N_18047);
or U18322 (N_18322,N_18194,N_18180);
xor U18323 (N_18323,N_18192,N_18128);
nand U18324 (N_18324,N_18133,N_18050);
xor U18325 (N_18325,N_18056,N_18093);
and U18326 (N_18326,N_18229,N_18138);
xor U18327 (N_18327,N_18033,N_18140);
xor U18328 (N_18328,N_18135,N_18233);
nand U18329 (N_18329,N_18175,N_18006);
nand U18330 (N_18330,N_18227,N_18049);
or U18331 (N_18331,N_18118,N_18030);
nor U18332 (N_18332,N_18150,N_18174);
xnor U18333 (N_18333,N_18212,N_18114);
or U18334 (N_18334,N_18055,N_18209);
nand U18335 (N_18335,N_18085,N_18109);
xor U18336 (N_18336,N_18223,N_18090);
and U18337 (N_18337,N_18053,N_18016);
nand U18338 (N_18338,N_18204,N_18037);
nor U18339 (N_18339,N_18168,N_18199);
xor U18340 (N_18340,N_18010,N_18071);
or U18341 (N_18341,N_18236,N_18153);
nand U18342 (N_18342,N_18067,N_18242);
nor U18343 (N_18343,N_18205,N_18162);
nand U18344 (N_18344,N_18059,N_18167);
and U18345 (N_18345,N_18235,N_18102);
nor U18346 (N_18346,N_18107,N_18046);
or U18347 (N_18347,N_18119,N_18013);
xnor U18348 (N_18348,N_18217,N_18230);
nand U18349 (N_18349,N_18005,N_18052);
nand U18350 (N_18350,N_18249,N_18163);
and U18351 (N_18351,N_18099,N_18072);
or U18352 (N_18352,N_18139,N_18017);
and U18353 (N_18353,N_18165,N_18196);
nor U18354 (N_18354,N_18066,N_18000);
and U18355 (N_18355,N_18171,N_18100);
nor U18356 (N_18356,N_18224,N_18225);
nor U18357 (N_18357,N_18183,N_18143);
nor U18358 (N_18358,N_18240,N_18151);
and U18359 (N_18359,N_18089,N_18203);
nand U18360 (N_18360,N_18147,N_18146);
and U18361 (N_18361,N_18080,N_18186);
xor U18362 (N_18362,N_18226,N_18086);
or U18363 (N_18363,N_18084,N_18221);
nor U18364 (N_18364,N_18248,N_18075);
nor U18365 (N_18365,N_18195,N_18155);
and U18366 (N_18366,N_18020,N_18136);
xnor U18367 (N_18367,N_18088,N_18026);
and U18368 (N_18368,N_18001,N_18116);
xnor U18369 (N_18369,N_18108,N_18104);
nand U18370 (N_18370,N_18097,N_18073);
nor U18371 (N_18371,N_18169,N_18070);
or U18372 (N_18372,N_18218,N_18022);
nor U18373 (N_18373,N_18228,N_18157);
xnor U18374 (N_18374,N_18149,N_18126);
nor U18375 (N_18375,N_18231,N_18101);
nand U18376 (N_18376,N_18133,N_18224);
xor U18377 (N_18377,N_18131,N_18083);
and U18378 (N_18378,N_18051,N_18209);
or U18379 (N_18379,N_18050,N_18173);
xnor U18380 (N_18380,N_18206,N_18068);
nand U18381 (N_18381,N_18189,N_18240);
or U18382 (N_18382,N_18167,N_18011);
and U18383 (N_18383,N_18105,N_18234);
xor U18384 (N_18384,N_18214,N_18109);
and U18385 (N_18385,N_18157,N_18185);
and U18386 (N_18386,N_18227,N_18123);
nor U18387 (N_18387,N_18226,N_18090);
xnor U18388 (N_18388,N_18219,N_18172);
xor U18389 (N_18389,N_18050,N_18104);
nand U18390 (N_18390,N_18143,N_18120);
or U18391 (N_18391,N_18210,N_18216);
and U18392 (N_18392,N_18046,N_18037);
nand U18393 (N_18393,N_18190,N_18140);
xor U18394 (N_18394,N_18114,N_18139);
or U18395 (N_18395,N_18228,N_18206);
xor U18396 (N_18396,N_18246,N_18152);
xor U18397 (N_18397,N_18136,N_18222);
xor U18398 (N_18398,N_18212,N_18218);
xnor U18399 (N_18399,N_18179,N_18110);
nor U18400 (N_18400,N_18099,N_18100);
nand U18401 (N_18401,N_18094,N_18036);
or U18402 (N_18402,N_18185,N_18183);
nor U18403 (N_18403,N_18077,N_18076);
and U18404 (N_18404,N_18233,N_18152);
nor U18405 (N_18405,N_18176,N_18246);
nand U18406 (N_18406,N_18100,N_18025);
or U18407 (N_18407,N_18017,N_18169);
nand U18408 (N_18408,N_18075,N_18072);
nor U18409 (N_18409,N_18198,N_18088);
nand U18410 (N_18410,N_18176,N_18210);
or U18411 (N_18411,N_18125,N_18004);
nor U18412 (N_18412,N_18244,N_18232);
or U18413 (N_18413,N_18141,N_18093);
and U18414 (N_18414,N_18201,N_18031);
or U18415 (N_18415,N_18091,N_18183);
or U18416 (N_18416,N_18194,N_18133);
nand U18417 (N_18417,N_18116,N_18114);
xnor U18418 (N_18418,N_18059,N_18142);
nand U18419 (N_18419,N_18107,N_18237);
nor U18420 (N_18420,N_18223,N_18180);
xnor U18421 (N_18421,N_18018,N_18012);
or U18422 (N_18422,N_18137,N_18063);
or U18423 (N_18423,N_18051,N_18109);
nand U18424 (N_18424,N_18011,N_18104);
and U18425 (N_18425,N_18198,N_18018);
xor U18426 (N_18426,N_18138,N_18166);
xnor U18427 (N_18427,N_18208,N_18017);
or U18428 (N_18428,N_18174,N_18112);
nor U18429 (N_18429,N_18096,N_18174);
nor U18430 (N_18430,N_18024,N_18037);
or U18431 (N_18431,N_18070,N_18152);
xor U18432 (N_18432,N_18228,N_18040);
nand U18433 (N_18433,N_18065,N_18203);
xor U18434 (N_18434,N_18231,N_18128);
nand U18435 (N_18435,N_18103,N_18199);
or U18436 (N_18436,N_18145,N_18120);
and U18437 (N_18437,N_18199,N_18121);
or U18438 (N_18438,N_18129,N_18019);
nor U18439 (N_18439,N_18054,N_18117);
nand U18440 (N_18440,N_18230,N_18189);
or U18441 (N_18441,N_18198,N_18195);
and U18442 (N_18442,N_18174,N_18179);
xor U18443 (N_18443,N_18208,N_18099);
and U18444 (N_18444,N_18192,N_18181);
nand U18445 (N_18445,N_18112,N_18182);
nor U18446 (N_18446,N_18058,N_18235);
or U18447 (N_18447,N_18010,N_18189);
and U18448 (N_18448,N_18113,N_18062);
nor U18449 (N_18449,N_18024,N_18218);
nand U18450 (N_18450,N_18099,N_18076);
or U18451 (N_18451,N_18180,N_18216);
or U18452 (N_18452,N_18090,N_18064);
nor U18453 (N_18453,N_18204,N_18014);
and U18454 (N_18454,N_18121,N_18158);
nor U18455 (N_18455,N_18117,N_18206);
xnor U18456 (N_18456,N_18053,N_18004);
or U18457 (N_18457,N_18003,N_18001);
or U18458 (N_18458,N_18143,N_18210);
nor U18459 (N_18459,N_18111,N_18094);
xor U18460 (N_18460,N_18024,N_18208);
nand U18461 (N_18461,N_18026,N_18046);
xnor U18462 (N_18462,N_18169,N_18042);
and U18463 (N_18463,N_18078,N_18216);
and U18464 (N_18464,N_18165,N_18119);
nor U18465 (N_18465,N_18140,N_18218);
and U18466 (N_18466,N_18147,N_18136);
or U18467 (N_18467,N_18018,N_18037);
xor U18468 (N_18468,N_18141,N_18232);
and U18469 (N_18469,N_18111,N_18057);
nand U18470 (N_18470,N_18044,N_18131);
nor U18471 (N_18471,N_18143,N_18140);
nand U18472 (N_18472,N_18012,N_18140);
or U18473 (N_18473,N_18207,N_18230);
nor U18474 (N_18474,N_18065,N_18031);
and U18475 (N_18475,N_18215,N_18186);
nand U18476 (N_18476,N_18145,N_18014);
xor U18477 (N_18477,N_18116,N_18063);
or U18478 (N_18478,N_18042,N_18000);
nor U18479 (N_18479,N_18072,N_18125);
or U18480 (N_18480,N_18221,N_18037);
nand U18481 (N_18481,N_18053,N_18148);
xor U18482 (N_18482,N_18166,N_18175);
nor U18483 (N_18483,N_18002,N_18235);
or U18484 (N_18484,N_18189,N_18044);
xor U18485 (N_18485,N_18061,N_18020);
and U18486 (N_18486,N_18035,N_18244);
xnor U18487 (N_18487,N_18149,N_18146);
nand U18488 (N_18488,N_18163,N_18162);
or U18489 (N_18489,N_18153,N_18097);
or U18490 (N_18490,N_18103,N_18015);
and U18491 (N_18491,N_18025,N_18088);
xnor U18492 (N_18492,N_18191,N_18245);
xnor U18493 (N_18493,N_18120,N_18241);
nor U18494 (N_18494,N_18165,N_18033);
nand U18495 (N_18495,N_18196,N_18175);
and U18496 (N_18496,N_18047,N_18183);
or U18497 (N_18497,N_18209,N_18241);
nor U18498 (N_18498,N_18047,N_18158);
xor U18499 (N_18499,N_18237,N_18243);
or U18500 (N_18500,N_18320,N_18368);
and U18501 (N_18501,N_18359,N_18350);
nor U18502 (N_18502,N_18307,N_18460);
nand U18503 (N_18503,N_18291,N_18436);
and U18504 (N_18504,N_18362,N_18272);
nand U18505 (N_18505,N_18377,N_18322);
nor U18506 (N_18506,N_18256,N_18407);
or U18507 (N_18507,N_18454,N_18496);
nand U18508 (N_18508,N_18458,N_18329);
and U18509 (N_18509,N_18472,N_18452);
nor U18510 (N_18510,N_18487,N_18393);
nor U18511 (N_18511,N_18367,N_18493);
or U18512 (N_18512,N_18342,N_18301);
xor U18513 (N_18513,N_18439,N_18463);
xor U18514 (N_18514,N_18478,N_18444);
xor U18515 (N_18515,N_18471,N_18315);
and U18516 (N_18516,N_18293,N_18282);
nor U18517 (N_18517,N_18442,N_18451);
nand U18518 (N_18518,N_18449,N_18354);
xnor U18519 (N_18519,N_18473,N_18404);
or U18520 (N_18520,N_18264,N_18382);
nand U18521 (N_18521,N_18428,N_18250);
or U18522 (N_18522,N_18369,N_18411);
nand U18523 (N_18523,N_18396,N_18319);
nor U18524 (N_18524,N_18426,N_18335);
or U18525 (N_18525,N_18317,N_18314);
and U18526 (N_18526,N_18459,N_18356);
xor U18527 (N_18527,N_18286,N_18448);
or U18528 (N_18528,N_18376,N_18366);
nor U18529 (N_18529,N_18347,N_18297);
nor U18530 (N_18530,N_18267,N_18495);
xor U18531 (N_18531,N_18419,N_18498);
nor U18532 (N_18532,N_18284,N_18421);
or U18533 (N_18533,N_18300,N_18289);
nor U18534 (N_18534,N_18384,N_18371);
xnor U18535 (N_18535,N_18405,N_18295);
or U18536 (N_18536,N_18497,N_18290);
nand U18537 (N_18537,N_18397,N_18346);
or U18538 (N_18538,N_18466,N_18309);
nor U18539 (N_18539,N_18398,N_18408);
or U18540 (N_18540,N_18488,N_18402);
nand U18541 (N_18541,N_18390,N_18255);
and U18542 (N_18542,N_18490,N_18324);
or U18543 (N_18543,N_18383,N_18365);
xor U18544 (N_18544,N_18283,N_18476);
or U18545 (N_18545,N_18406,N_18330);
nand U18546 (N_18546,N_18430,N_18386);
and U18547 (N_18547,N_18344,N_18341);
and U18548 (N_18548,N_18394,N_18468);
nor U18549 (N_18549,N_18378,N_18310);
and U18550 (N_18550,N_18279,N_18361);
nor U18551 (N_18551,N_18296,N_18374);
or U18552 (N_18552,N_18491,N_18380);
nand U18553 (N_18553,N_18266,N_18364);
nor U18554 (N_18554,N_18326,N_18425);
nand U18555 (N_18555,N_18259,N_18446);
or U18556 (N_18556,N_18433,N_18464);
or U18557 (N_18557,N_18265,N_18440);
or U18558 (N_18558,N_18303,N_18323);
or U18559 (N_18559,N_18429,N_18260);
and U18560 (N_18560,N_18263,N_18370);
and U18561 (N_18561,N_18340,N_18399);
xnor U18562 (N_18562,N_18270,N_18328);
and U18563 (N_18563,N_18373,N_18308);
nand U18564 (N_18564,N_18338,N_18312);
nand U18565 (N_18565,N_18434,N_18273);
nor U18566 (N_18566,N_18486,N_18331);
xnor U18567 (N_18567,N_18353,N_18349);
nor U18568 (N_18568,N_18432,N_18418);
nand U18569 (N_18569,N_18274,N_18336);
or U18570 (N_18570,N_18483,N_18254);
and U18571 (N_18571,N_18325,N_18489);
nor U18572 (N_18572,N_18455,N_18343);
or U18573 (N_18573,N_18400,N_18431);
nand U18574 (N_18574,N_18494,N_18392);
nor U18575 (N_18575,N_18253,N_18316);
xnor U18576 (N_18576,N_18420,N_18414);
or U18577 (N_18577,N_18480,N_18287);
and U18578 (N_18578,N_18281,N_18437);
nand U18579 (N_18579,N_18339,N_18299);
nor U18580 (N_18580,N_18288,N_18352);
nand U18581 (N_18581,N_18395,N_18276);
xnor U18582 (N_18582,N_18348,N_18492);
or U18583 (N_18583,N_18381,N_18337);
and U18584 (N_18584,N_18461,N_18484);
nor U18585 (N_18585,N_18363,N_18262);
and U18586 (N_18586,N_18391,N_18305);
or U18587 (N_18587,N_18403,N_18424);
nor U18588 (N_18588,N_18292,N_18360);
nor U18589 (N_18589,N_18306,N_18417);
xor U18590 (N_18590,N_18499,N_18457);
and U18591 (N_18591,N_18422,N_18278);
or U18592 (N_18592,N_18304,N_18470);
nor U18593 (N_18593,N_18401,N_18412);
nor U18594 (N_18594,N_18447,N_18477);
nand U18595 (N_18595,N_18427,N_18327);
nand U18596 (N_18596,N_18481,N_18318);
nor U18597 (N_18597,N_18257,N_18271);
xnor U18598 (N_18598,N_18443,N_18413);
and U18599 (N_18599,N_18475,N_18467);
and U18600 (N_18600,N_18258,N_18357);
or U18601 (N_18601,N_18333,N_18294);
nor U18602 (N_18602,N_18251,N_18261);
xnor U18603 (N_18603,N_18332,N_18416);
nor U18604 (N_18604,N_18479,N_18275);
or U18605 (N_18605,N_18423,N_18269);
nor U18606 (N_18606,N_18438,N_18379);
xor U18607 (N_18607,N_18388,N_18358);
and U18608 (N_18608,N_18387,N_18313);
xor U18609 (N_18609,N_18474,N_18465);
and U18610 (N_18610,N_18385,N_18462);
or U18611 (N_18611,N_18334,N_18456);
nand U18612 (N_18612,N_18445,N_18469);
or U18613 (N_18613,N_18252,N_18453);
nand U18614 (N_18614,N_18302,N_18355);
nand U18615 (N_18615,N_18321,N_18482);
xnor U18616 (N_18616,N_18389,N_18435);
or U18617 (N_18617,N_18375,N_18298);
or U18618 (N_18618,N_18268,N_18311);
xnor U18619 (N_18619,N_18345,N_18485);
nand U18620 (N_18620,N_18409,N_18372);
nand U18621 (N_18621,N_18415,N_18285);
and U18622 (N_18622,N_18351,N_18441);
or U18623 (N_18623,N_18410,N_18450);
nor U18624 (N_18624,N_18277,N_18280);
and U18625 (N_18625,N_18361,N_18331);
and U18626 (N_18626,N_18472,N_18475);
nor U18627 (N_18627,N_18446,N_18460);
or U18628 (N_18628,N_18281,N_18372);
or U18629 (N_18629,N_18479,N_18420);
nand U18630 (N_18630,N_18399,N_18404);
and U18631 (N_18631,N_18274,N_18409);
or U18632 (N_18632,N_18334,N_18388);
and U18633 (N_18633,N_18321,N_18369);
or U18634 (N_18634,N_18311,N_18310);
and U18635 (N_18635,N_18348,N_18265);
and U18636 (N_18636,N_18271,N_18387);
and U18637 (N_18637,N_18444,N_18434);
xnor U18638 (N_18638,N_18329,N_18304);
nor U18639 (N_18639,N_18280,N_18292);
xnor U18640 (N_18640,N_18291,N_18491);
or U18641 (N_18641,N_18298,N_18285);
and U18642 (N_18642,N_18271,N_18265);
and U18643 (N_18643,N_18363,N_18441);
nor U18644 (N_18644,N_18307,N_18356);
or U18645 (N_18645,N_18493,N_18418);
or U18646 (N_18646,N_18299,N_18334);
nor U18647 (N_18647,N_18478,N_18380);
or U18648 (N_18648,N_18383,N_18310);
xnor U18649 (N_18649,N_18469,N_18341);
and U18650 (N_18650,N_18396,N_18485);
and U18651 (N_18651,N_18372,N_18480);
and U18652 (N_18652,N_18277,N_18377);
nor U18653 (N_18653,N_18368,N_18317);
xor U18654 (N_18654,N_18251,N_18389);
or U18655 (N_18655,N_18388,N_18294);
xor U18656 (N_18656,N_18484,N_18455);
xor U18657 (N_18657,N_18356,N_18276);
and U18658 (N_18658,N_18292,N_18474);
and U18659 (N_18659,N_18365,N_18403);
nor U18660 (N_18660,N_18260,N_18345);
nor U18661 (N_18661,N_18483,N_18371);
nand U18662 (N_18662,N_18319,N_18291);
and U18663 (N_18663,N_18456,N_18439);
and U18664 (N_18664,N_18440,N_18292);
nand U18665 (N_18665,N_18493,N_18314);
nand U18666 (N_18666,N_18403,N_18269);
nor U18667 (N_18667,N_18476,N_18417);
nand U18668 (N_18668,N_18355,N_18326);
or U18669 (N_18669,N_18397,N_18443);
xor U18670 (N_18670,N_18379,N_18416);
nand U18671 (N_18671,N_18318,N_18427);
or U18672 (N_18672,N_18346,N_18351);
xnor U18673 (N_18673,N_18285,N_18412);
and U18674 (N_18674,N_18287,N_18297);
nand U18675 (N_18675,N_18393,N_18453);
nor U18676 (N_18676,N_18319,N_18268);
nand U18677 (N_18677,N_18279,N_18434);
and U18678 (N_18678,N_18252,N_18480);
and U18679 (N_18679,N_18332,N_18393);
nand U18680 (N_18680,N_18350,N_18268);
nand U18681 (N_18681,N_18397,N_18309);
or U18682 (N_18682,N_18275,N_18343);
nand U18683 (N_18683,N_18295,N_18279);
or U18684 (N_18684,N_18358,N_18431);
nand U18685 (N_18685,N_18443,N_18261);
xor U18686 (N_18686,N_18416,N_18283);
or U18687 (N_18687,N_18387,N_18320);
xor U18688 (N_18688,N_18298,N_18449);
and U18689 (N_18689,N_18410,N_18379);
nand U18690 (N_18690,N_18322,N_18305);
nor U18691 (N_18691,N_18471,N_18267);
nor U18692 (N_18692,N_18421,N_18345);
and U18693 (N_18693,N_18274,N_18468);
nand U18694 (N_18694,N_18413,N_18292);
nor U18695 (N_18695,N_18486,N_18435);
nand U18696 (N_18696,N_18340,N_18496);
nand U18697 (N_18697,N_18440,N_18359);
or U18698 (N_18698,N_18464,N_18413);
or U18699 (N_18699,N_18344,N_18438);
xnor U18700 (N_18700,N_18303,N_18319);
and U18701 (N_18701,N_18259,N_18380);
nand U18702 (N_18702,N_18457,N_18429);
and U18703 (N_18703,N_18419,N_18389);
nor U18704 (N_18704,N_18445,N_18456);
nor U18705 (N_18705,N_18337,N_18439);
nor U18706 (N_18706,N_18265,N_18443);
xnor U18707 (N_18707,N_18277,N_18426);
and U18708 (N_18708,N_18437,N_18279);
nor U18709 (N_18709,N_18474,N_18464);
xor U18710 (N_18710,N_18449,N_18337);
and U18711 (N_18711,N_18370,N_18435);
and U18712 (N_18712,N_18393,N_18495);
xnor U18713 (N_18713,N_18251,N_18439);
nand U18714 (N_18714,N_18485,N_18480);
nand U18715 (N_18715,N_18333,N_18455);
nor U18716 (N_18716,N_18274,N_18395);
nor U18717 (N_18717,N_18281,N_18260);
xor U18718 (N_18718,N_18466,N_18300);
nand U18719 (N_18719,N_18340,N_18360);
or U18720 (N_18720,N_18415,N_18352);
xor U18721 (N_18721,N_18494,N_18481);
nor U18722 (N_18722,N_18321,N_18415);
xor U18723 (N_18723,N_18366,N_18291);
nor U18724 (N_18724,N_18496,N_18278);
or U18725 (N_18725,N_18291,N_18363);
nor U18726 (N_18726,N_18352,N_18316);
or U18727 (N_18727,N_18405,N_18277);
xnor U18728 (N_18728,N_18339,N_18361);
nand U18729 (N_18729,N_18433,N_18340);
xor U18730 (N_18730,N_18450,N_18250);
nor U18731 (N_18731,N_18390,N_18416);
nor U18732 (N_18732,N_18412,N_18478);
xnor U18733 (N_18733,N_18253,N_18290);
xnor U18734 (N_18734,N_18253,N_18366);
nand U18735 (N_18735,N_18300,N_18354);
nor U18736 (N_18736,N_18422,N_18481);
xnor U18737 (N_18737,N_18284,N_18276);
or U18738 (N_18738,N_18435,N_18446);
nand U18739 (N_18739,N_18280,N_18261);
nand U18740 (N_18740,N_18497,N_18484);
nor U18741 (N_18741,N_18465,N_18351);
and U18742 (N_18742,N_18450,N_18303);
nor U18743 (N_18743,N_18354,N_18433);
nor U18744 (N_18744,N_18449,N_18261);
nand U18745 (N_18745,N_18441,N_18471);
nor U18746 (N_18746,N_18326,N_18336);
nor U18747 (N_18747,N_18496,N_18346);
nand U18748 (N_18748,N_18314,N_18444);
xnor U18749 (N_18749,N_18401,N_18414);
or U18750 (N_18750,N_18745,N_18675);
or U18751 (N_18751,N_18652,N_18696);
or U18752 (N_18752,N_18623,N_18731);
and U18753 (N_18753,N_18723,N_18685);
nor U18754 (N_18754,N_18639,N_18581);
nand U18755 (N_18755,N_18563,N_18559);
xnor U18756 (N_18756,N_18735,N_18688);
or U18757 (N_18757,N_18718,N_18746);
and U18758 (N_18758,N_18749,N_18504);
nor U18759 (N_18759,N_18615,N_18592);
and U18760 (N_18760,N_18620,N_18614);
nor U18761 (N_18761,N_18714,N_18515);
xnor U18762 (N_18762,N_18534,N_18636);
nand U18763 (N_18763,N_18656,N_18740);
nand U18764 (N_18764,N_18719,N_18514);
or U18765 (N_18765,N_18520,N_18642);
or U18766 (N_18766,N_18533,N_18694);
xor U18767 (N_18767,N_18609,N_18687);
and U18768 (N_18768,N_18727,N_18622);
and U18769 (N_18769,N_18627,N_18630);
or U18770 (N_18770,N_18500,N_18683);
xor U18771 (N_18771,N_18513,N_18522);
and U18772 (N_18772,N_18698,N_18655);
xnor U18773 (N_18773,N_18547,N_18743);
xor U18774 (N_18774,N_18552,N_18624);
or U18775 (N_18775,N_18695,N_18692);
xor U18776 (N_18776,N_18607,N_18539);
or U18777 (N_18777,N_18701,N_18549);
or U18778 (N_18778,N_18631,N_18645);
xnor U18779 (N_18779,N_18664,N_18716);
nor U18780 (N_18780,N_18703,N_18670);
nand U18781 (N_18781,N_18728,N_18597);
xor U18782 (N_18782,N_18528,N_18646);
or U18783 (N_18783,N_18674,N_18565);
nand U18784 (N_18784,N_18548,N_18598);
xnor U18785 (N_18785,N_18576,N_18594);
xor U18786 (N_18786,N_18734,N_18681);
xor U18787 (N_18787,N_18566,N_18577);
nor U18788 (N_18788,N_18574,N_18625);
and U18789 (N_18789,N_18556,N_18721);
and U18790 (N_18790,N_18562,N_18715);
nor U18791 (N_18791,N_18545,N_18658);
and U18792 (N_18792,N_18712,N_18693);
nand U18793 (N_18793,N_18617,N_18725);
nor U18794 (N_18794,N_18544,N_18519);
nand U18795 (N_18795,N_18629,N_18575);
and U18796 (N_18796,N_18557,N_18732);
xor U18797 (N_18797,N_18573,N_18593);
xor U18798 (N_18798,N_18708,N_18635);
nor U18799 (N_18799,N_18516,N_18682);
and U18800 (N_18800,N_18705,N_18676);
and U18801 (N_18801,N_18568,N_18741);
nor U18802 (N_18802,N_18700,N_18521);
nand U18803 (N_18803,N_18569,N_18707);
and U18804 (N_18804,N_18668,N_18553);
and U18805 (N_18805,N_18748,N_18579);
nor U18806 (N_18806,N_18659,N_18643);
and U18807 (N_18807,N_18724,N_18512);
nand U18808 (N_18808,N_18738,N_18508);
nor U18809 (N_18809,N_18634,N_18628);
nor U18810 (N_18810,N_18564,N_18689);
and U18811 (N_18811,N_18611,N_18591);
nand U18812 (N_18812,N_18684,N_18587);
nor U18813 (N_18813,N_18527,N_18578);
xor U18814 (N_18814,N_18717,N_18726);
and U18815 (N_18815,N_18526,N_18601);
nor U18816 (N_18816,N_18546,N_18518);
xnor U18817 (N_18817,N_18501,N_18671);
or U18818 (N_18818,N_18686,N_18509);
and U18819 (N_18819,N_18604,N_18637);
nor U18820 (N_18820,N_18644,N_18602);
nor U18821 (N_18821,N_18742,N_18507);
or U18822 (N_18822,N_18543,N_18502);
nor U18823 (N_18823,N_18649,N_18610);
or U18824 (N_18824,N_18603,N_18517);
xnor U18825 (N_18825,N_18572,N_18679);
xor U18826 (N_18826,N_18720,N_18555);
xnor U18827 (N_18827,N_18669,N_18541);
nor U18828 (N_18828,N_18632,N_18678);
xnor U18829 (N_18829,N_18744,N_18747);
xor U18830 (N_18830,N_18595,N_18551);
nand U18831 (N_18831,N_18641,N_18626);
nor U18832 (N_18832,N_18503,N_18638);
nand U18833 (N_18833,N_18648,N_18677);
and U18834 (N_18834,N_18554,N_18506);
nand U18835 (N_18835,N_18699,N_18640);
nor U18836 (N_18836,N_18713,N_18691);
or U18837 (N_18837,N_18733,N_18662);
nor U18838 (N_18838,N_18612,N_18653);
nor U18839 (N_18839,N_18529,N_18661);
nor U18840 (N_18840,N_18524,N_18580);
and U18841 (N_18841,N_18511,N_18672);
or U18842 (N_18842,N_18600,N_18540);
and U18843 (N_18843,N_18505,N_18616);
nor U18844 (N_18844,N_18730,N_18673);
xnor U18845 (N_18845,N_18571,N_18702);
or U18846 (N_18846,N_18599,N_18567);
or U18847 (N_18847,N_18704,N_18589);
nor U18848 (N_18848,N_18537,N_18710);
and U18849 (N_18849,N_18583,N_18584);
xnor U18850 (N_18850,N_18690,N_18558);
xnor U18851 (N_18851,N_18586,N_18621);
nand U18852 (N_18852,N_18585,N_18596);
xor U18853 (N_18853,N_18510,N_18542);
or U18854 (N_18854,N_18561,N_18666);
and U18855 (N_18855,N_18608,N_18737);
nand U18856 (N_18856,N_18657,N_18619);
nand U18857 (N_18857,N_18536,N_18538);
xnor U18858 (N_18858,N_18660,N_18582);
or U18859 (N_18859,N_18618,N_18665);
nor U18860 (N_18860,N_18667,N_18680);
xor U18861 (N_18861,N_18651,N_18532);
or U18862 (N_18862,N_18722,N_18706);
nor U18863 (N_18863,N_18570,N_18729);
and U18864 (N_18864,N_18654,N_18736);
nor U18865 (N_18865,N_18605,N_18739);
nand U18866 (N_18866,N_18590,N_18633);
and U18867 (N_18867,N_18613,N_18606);
nand U18868 (N_18868,N_18535,N_18531);
nor U18869 (N_18869,N_18647,N_18709);
nand U18870 (N_18870,N_18530,N_18525);
nor U18871 (N_18871,N_18697,N_18560);
xor U18872 (N_18872,N_18550,N_18650);
nor U18873 (N_18873,N_18523,N_18663);
and U18874 (N_18874,N_18588,N_18711);
or U18875 (N_18875,N_18587,N_18731);
nand U18876 (N_18876,N_18671,N_18722);
nand U18877 (N_18877,N_18714,N_18565);
xor U18878 (N_18878,N_18714,N_18588);
nor U18879 (N_18879,N_18622,N_18722);
nor U18880 (N_18880,N_18671,N_18658);
nor U18881 (N_18881,N_18670,N_18673);
nor U18882 (N_18882,N_18548,N_18717);
nand U18883 (N_18883,N_18508,N_18611);
nand U18884 (N_18884,N_18568,N_18599);
nor U18885 (N_18885,N_18707,N_18530);
xor U18886 (N_18886,N_18575,N_18581);
nor U18887 (N_18887,N_18678,N_18509);
nand U18888 (N_18888,N_18722,N_18698);
nand U18889 (N_18889,N_18743,N_18580);
or U18890 (N_18890,N_18691,N_18503);
nand U18891 (N_18891,N_18500,N_18509);
and U18892 (N_18892,N_18591,N_18555);
or U18893 (N_18893,N_18561,N_18627);
and U18894 (N_18894,N_18591,N_18725);
xor U18895 (N_18895,N_18585,N_18516);
and U18896 (N_18896,N_18506,N_18717);
xor U18897 (N_18897,N_18641,N_18625);
xor U18898 (N_18898,N_18640,N_18636);
nor U18899 (N_18899,N_18613,N_18533);
nor U18900 (N_18900,N_18521,N_18649);
nor U18901 (N_18901,N_18614,N_18749);
nand U18902 (N_18902,N_18529,N_18710);
and U18903 (N_18903,N_18599,N_18681);
xor U18904 (N_18904,N_18629,N_18569);
nor U18905 (N_18905,N_18582,N_18713);
nand U18906 (N_18906,N_18516,N_18676);
nand U18907 (N_18907,N_18517,N_18656);
or U18908 (N_18908,N_18599,N_18749);
nand U18909 (N_18909,N_18737,N_18561);
xor U18910 (N_18910,N_18528,N_18575);
xor U18911 (N_18911,N_18703,N_18702);
xnor U18912 (N_18912,N_18589,N_18547);
nand U18913 (N_18913,N_18618,N_18507);
and U18914 (N_18914,N_18521,N_18639);
and U18915 (N_18915,N_18717,N_18534);
and U18916 (N_18916,N_18662,N_18515);
xnor U18917 (N_18917,N_18534,N_18723);
or U18918 (N_18918,N_18678,N_18670);
nor U18919 (N_18919,N_18544,N_18717);
or U18920 (N_18920,N_18651,N_18740);
and U18921 (N_18921,N_18619,N_18533);
xnor U18922 (N_18922,N_18525,N_18697);
xor U18923 (N_18923,N_18633,N_18688);
xor U18924 (N_18924,N_18685,N_18586);
or U18925 (N_18925,N_18640,N_18620);
nand U18926 (N_18926,N_18618,N_18605);
and U18927 (N_18927,N_18638,N_18656);
nor U18928 (N_18928,N_18648,N_18511);
nor U18929 (N_18929,N_18500,N_18604);
xnor U18930 (N_18930,N_18722,N_18720);
nand U18931 (N_18931,N_18654,N_18553);
nand U18932 (N_18932,N_18515,N_18703);
or U18933 (N_18933,N_18693,N_18741);
nor U18934 (N_18934,N_18591,N_18582);
and U18935 (N_18935,N_18548,N_18609);
or U18936 (N_18936,N_18510,N_18512);
and U18937 (N_18937,N_18618,N_18564);
or U18938 (N_18938,N_18507,N_18692);
nor U18939 (N_18939,N_18580,N_18677);
nand U18940 (N_18940,N_18729,N_18540);
or U18941 (N_18941,N_18601,N_18696);
nor U18942 (N_18942,N_18503,N_18621);
nand U18943 (N_18943,N_18737,N_18676);
nor U18944 (N_18944,N_18616,N_18684);
nand U18945 (N_18945,N_18609,N_18601);
nor U18946 (N_18946,N_18568,N_18708);
nand U18947 (N_18947,N_18730,N_18662);
xor U18948 (N_18948,N_18677,N_18657);
nand U18949 (N_18949,N_18591,N_18576);
xor U18950 (N_18950,N_18652,N_18732);
or U18951 (N_18951,N_18665,N_18578);
or U18952 (N_18952,N_18633,N_18671);
and U18953 (N_18953,N_18690,N_18579);
xor U18954 (N_18954,N_18691,N_18699);
nor U18955 (N_18955,N_18633,N_18617);
or U18956 (N_18956,N_18617,N_18644);
or U18957 (N_18957,N_18606,N_18669);
xor U18958 (N_18958,N_18621,N_18538);
xor U18959 (N_18959,N_18527,N_18507);
or U18960 (N_18960,N_18514,N_18659);
or U18961 (N_18961,N_18516,N_18746);
nor U18962 (N_18962,N_18747,N_18522);
nand U18963 (N_18963,N_18602,N_18696);
xnor U18964 (N_18964,N_18504,N_18577);
and U18965 (N_18965,N_18607,N_18529);
nand U18966 (N_18966,N_18690,N_18708);
xor U18967 (N_18967,N_18587,N_18694);
and U18968 (N_18968,N_18567,N_18655);
nor U18969 (N_18969,N_18557,N_18527);
and U18970 (N_18970,N_18574,N_18520);
and U18971 (N_18971,N_18651,N_18666);
nand U18972 (N_18972,N_18747,N_18707);
nor U18973 (N_18973,N_18662,N_18724);
and U18974 (N_18974,N_18525,N_18667);
and U18975 (N_18975,N_18555,N_18610);
and U18976 (N_18976,N_18683,N_18574);
nor U18977 (N_18977,N_18579,N_18672);
nor U18978 (N_18978,N_18573,N_18609);
nand U18979 (N_18979,N_18743,N_18530);
xor U18980 (N_18980,N_18627,N_18512);
or U18981 (N_18981,N_18508,N_18549);
and U18982 (N_18982,N_18705,N_18729);
nor U18983 (N_18983,N_18544,N_18709);
or U18984 (N_18984,N_18699,N_18718);
or U18985 (N_18985,N_18736,N_18728);
or U18986 (N_18986,N_18515,N_18562);
nor U18987 (N_18987,N_18538,N_18737);
and U18988 (N_18988,N_18552,N_18600);
nand U18989 (N_18989,N_18683,N_18525);
or U18990 (N_18990,N_18621,N_18679);
xnor U18991 (N_18991,N_18736,N_18743);
nor U18992 (N_18992,N_18588,N_18506);
nor U18993 (N_18993,N_18608,N_18514);
xnor U18994 (N_18994,N_18591,N_18521);
nand U18995 (N_18995,N_18655,N_18597);
or U18996 (N_18996,N_18524,N_18724);
xor U18997 (N_18997,N_18744,N_18736);
and U18998 (N_18998,N_18648,N_18643);
nor U18999 (N_18999,N_18513,N_18748);
and U19000 (N_19000,N_18948,N_18818);
nor U19001 (N_19001,N_18898,N_18793);
or U19002 (N_19002,N_18972,N_18815);
and U19003 (N_19003,N_18849,N_18755);
or U19004 (N_19004,N_18937,N_18891);
nand U19005 (N_19005,N_18901,N_18969);
nor U19006 (N_19006,N_18753,N_18855);
and U19007 (N_19007,N_18922,N_18857);
nor U19008 (N_19008,N_18760,N_18772);
nor U19009 (N_19009,N_18991,N_18863);
or U19010 (N_19010,N_18955,N_18795);
and U19011 (N_19011,N_18750,N_18784);
nand U19012 (N_19012,N_18756,N_18830);
nand U19013 (N_19013,N_18771,N_18912);
and U19014 (N_19014,N_18986,N_18757);
and U19015 (N_19015,N_18866,N_18943);
and U19016 (N_19016,N_18927,N_18981);
and U19017 (N_19017,N_18964,N_18929);
and U19018 (N_19018,N_18900,N_18785);
xor U19019 (N_19019,N_18957,N_18836);
or U19020 (N_19020,N_18769,N_18832);
nand U19021 (N_19021,N_18761,N_18819);
or U19022 (N_19022,N_18966,N_18938);
or U19023 (N_19023,N_18861,N_18848);
nand U19024 (N_19024,N_18873,N_18934);
nand U19025 (N_19025,N_18919,N_18959);
and U19026 (N_19026,N_18965,N_18877);
nor U19027 (N_19027,N_18961,N_18988);
or U19028 (N_19028,N_18839,N_18928);
xor U19029 (N_19029,N_18899,N_18828);
or U19030 (N_19030,N_18767,N_18978);
and U19031 (N_19031,N_18781,N_18896);
nand U19032 (N_19032,N_18773,N_18997);
and U19033 (N_19033,N_18926,N_18947);
nor U19034 (N_19034,N_18810,N_18834);
nand U19035 (N_19035,N_18801,N_18881);
xnor U19036 (N_19036,N_18942,N_18870);
and U19037 (N_19037,N_18921,N_18915);
xnor U19038 (N_19038,N_18875,N_18782);
xor U19039 (N_19039,N_18847,N_18882);
nand U19040 (N_19040,N_18953,N_18951);
and U19041 (N_19041,N_18952,N_18800);
or U19042 (N_19042,N_18917,N_18960);
nor U19043 (N_19043,N_18802,N_18995);
or U19044 (N_19044,N_18876,N_18764);
or U19045 (N_19045,N_18843,N_18987);
xor U19046 (N_19046,N_18977,N_18844);
nand U19047 (N_19047,N_18813,N_18907);
or U19048 (N_19048,N_18910,N_18887);
nor U19049 (N_19049,N_18918,N_18833);
and U19050 (N_19050,N_18804,N_18860);
nand U19051 (N_19051,N_18923,N_18759);
nor U19052 (N_19052,N_18975,N_18998);
xor U19053 (N_19053,N_18854,N_18940);
xnor U19054 (N_19054,N_18913,N_18869);
xnor U19055 (N_19055,N_18858,N_18989);
or U19056 (N_19056,N_18846,N_18797);
and U19057 (N_19057,N_18814,N_18768);
nand U19058 (N_19058,N_18851,N_18897);
and U19059 (N_19059,N_18984,N_18778);
nand U19060 (N_19060,N_18889,N_18976);
xnor U19061 (N_19061,N_18871,N_18852);
and U19062 (N_19062,N_18968,N_18980);
and U19063 (N_19063,N_18974,N_18758);
nor U19064 (N_19064,N_18932,N_18754);
or U19065 (N_19065,N_18763,N_18821);
and U19066 (N_19066,N_18812,N_18809);
or U19067 (N_19067,N_18967,N_18983);
or U19068 (N_19068,N_18874,N_18762);
xnor U19069 (N_19069,N_18894,N_18825);
xor U19070 (N_19070,N_18794,N_18816);
and U19071 (N_19071,N_18783,N_18950);
nor U19072 (N_19072,N_18982,N_18779);
and U19073 (N_19073,N_18787,N_18751);
xor U19074 (N_19074,N_18841,N_18837);
nor U19075 (N_19075,N_18970,N_18798);
xnor U19076 (N_19076,N_18880,N_18935);
and U19077 (N_19077,N_18890,N_18805);
nor U19078 (N_19078,N_18776,N_18808);
nor U19079 (N_19079,N_18840,N_18822);
or U19080 (N_19080,N_18817,N_18905);
and U19081 (N_19081,N_18920,N_18823);
nor U19082 (N_19082,N_18831,N_18916);
nand U19083 (N_19083,N_18909,N_18949);
xnor U19084 (N_19084,N_18936,N_18944);
or U19085 (N_19085,N_18946,N_18850);
and U19086 (N_19086,N_18799,N_18956);
nand U19087 (N_19087,N_18992,N_18806);
or U19088 (N_19088,N_18883,N_18811);
or U19089 (N_19089,N_18902,N_18914);
nand U19090 (N_19090,N_18867,N_18954);
nor U19091 (N_19091,N_18990,N_18985);
and U19092 (N_19092,N_18971,N_18765);
nor U19093 (N_19093,N_18827,N_18796);
and U19094 (N_19094,N_18973,N_18993);
and U19095 (N_19095,N_18963,N_18777);
or U19096 (N_19096,N_18864,N_18885);
and U19097 (N_19097,N_18842,N_18826);
and U19098 (N_19098,N_18792,N_18791);
xor U19099 (N_19099,N_18945,N_18979);
nand U19100 (N_19100,N_18886,N_18911);
nand U19101 (N_19101,N_18930,N_18962);
or U19102 (N_19102,N_18994,N_18924);
nand U19103 (N_19103,N_18892,N_18752);
xor U19104 (N_19104,N_18788,N_18933);
and U19105 (N_19105,N_18824,N_18939);
and U19106 (N_19106,N_18775,N_18879);
xnor U19107 (N_19107,N_18878,N_18770);
xnor U19108 (N_19108,N_18862,N_18853);
xor U19109 (N_19109,N_18895,N_18845);
or U19110 (N_19110,N_18835,N_18856);
xnor U19111 (N_19111,N_18868,N_18931);
or U19112 (N_19112,N_18893,N_18925);
nor U19113 (N_19113,N_18838,N_18872);
nand U19114 (N_19114,N_18884,N_18766);
xor U19115 (N_19115,N_18786,N_18790);
or U19116 (N_19116,N_18903,N_18865);
and U19117 (N_19117,N_18774,N_18958);
and U19118 (N_19118,N_18803,N_18999);
or U19119 (N_19119,N_18941,N_18859);
nor U19120 (N_19120,N_18904,N_18807);
xnor U19121 (N_19121,N_18888,N_18908);
nand U19122 (N_19122,N_18820,N_18780);
and U19123 (N_19123,N_18906,N_18996);
nand U19124 (N_19124,N_18789,N_18829);
or U19125 (N_19125,N_18881,N_18838);
xnor U19126 (N_19126,N_18826,N_18809);
nand U19127 (N_19127,N_18896,N_18798);
xor U19128 (N_19128,N_18751,N_18924);
nand U19129 (N_19129,N_18933,N_18782);
nor U19130 (N_19130,N_18832,N_18810);
xor U19131 (N_19131,N_18925,N_18899);
nor U19132 (N_19132,N_18877,N_18904);
or U19133 (N_19133,N_18826,N_18967);
nand U19134 (N_19134,N_18955,N_18811);
nand U19135 (N_19135,N_18951,N_18821);
and U19136 (N_19136,N_18803,N_18847);
and U19137 (N_19137,N_18904,N_18947);
xor U19138 (N_19138,N_18752,N_18976);
xnor U19139 (N_19139,N_18861,N_18826);
and U19140 (N_19140,N_18955,N_18933);
or U19141 (N_19141,N_18805,N_18995);
or U19142 (N_19142,N_18800,N_18818);
or U19143 (N_19143,N_18916,N_18941);
nand U19144 (N_19144,N_18756,N_18914);
nand U19145 (N_19145,N_18931,N_18774);
nand U19146 (N_19146,N_18760,N_18901);
or U19147 (N_19147,N_18794,N_18869);
nand U19148 (N_19148,N_18804,N_18785);
xnor U19149 (N_19149,N_18865,N_18979);
or U19150 (N_19150,N_18986,N_18950);
or U19151 (N_19151,N_18762,N_18884);
or U19152 (N_19152,N_18805,N_18942);
and U19153 (N_19153,N_18758,N_18871);
nor U19154 (N_19154,N_18812,N_18882);
xnor U19155 (N_19155,N_18753,N_18850);
xnor U19156 (N_19156,N_18792,N_18829);
nor U19157 (N_19157,N_18840,N_18993);
nor U19158 (N_19158,N_18925,N_18954);
and U19159 (N_19159,N_18845,N_18986);
or U19160 (N_19160,N_18822,N_18849);
nand U19161 (N_19161,N_18878,N_18918);
nor U19162 (N_19162,N_18794,N_18776);
nor U19163 (N_19163,N_18978,N_18818);
nand U19164 (N_19164,N_18808,N_18793);
nor U19165 (N_19165,N_18871,N_18895);
and U19166 (N_19166,N_18920,N_18998);
xnor U19167 (N_19167,N_18791,N_18869);
nor U19168 (N_19168,N_18794,N_18918);
xor U19169 (N_19169,N_18904,N_18980);
xnor U19170 (N_19170,N_18790,N_18881);
and U19171 (N_19171,N_18947,N_18851);
xnor U19172 (N_19172,N_18918,N_18954);
or U19173 (N_19173,N_18759,N_18971);
nor U19174 (N_19174,N_18870,N_18754);
or U19175 (N_19175,N_18891,N_18975);
xnor U19176 (N_19176,N_18826,N_18785);
or U19177 (N_19177,N_18883,N_18826);
or U19178 (N_19178,N_18950,N_18888);
xnor U19179 (N_19179,N_18939,N_18797);
nand U19180 (N_19180,N_18896,N_18851);
nand U19181 (N_19181,N_18975,N_18838);
nor U19182 (N_19182,N_18868,N_18893);
nor U19183 (N_19183,N_18993,N_18864);
nor U19184 (N_19184,N_18983,N_18951);
nand U19185 (N_19185,N_18978,N_18807);
and U19186 (N_19186,N_18879,N_18973);
or U19187 (N_19187,N_18901,N_18953);
and U19188 (N_19188,N_18764,N_18998);
and U19189 (N_19189,N_18802,N_18751);
or U19190 (N_19190,N_18874,N_18939);
nor U19191 (N_19191,N_18955,N_18842);
xor U19192 (N_19192,N_18929,N_18943);
nand U19193 (N_19193,N_18999,N_18794);
xnor U19194 (N_19194,N_18822,N_18781);
nor U19195 (N_19195,N_18943,N_18905);
and U19196 (N_19196,N_18961,N_18838);
xnor U19197 (N_19197,N_18969,N_18876);
and U19198 (N_19198,N_18841,N_18923);
nand U19199 (N_19199,N_18912,N_18834);
nor U19200 (N_19200,N_18980,N_18770);
xnor U19201 (N_19201,N_18761,N_18944);
xor U19202 (N_19202,N_18992,N_18765);
nand U19203 (N_19203,N_18988,N_18791);
nand U19204 (N_19204,N_18853,N_18947);
or U19205 (N_19205,N_18878,N_18787);
xor U19206 (N_19206,N_18803,N_18758);
nand U19207 (N_19207,N_18844,N_18976);
or U19208 (N_19208,N_18992,N_18860);
and U19209 (N_19209,N_18998,N_18958);
nand U19210 (N_19210,N_18800,N_18756);
or U19211 (N_19211,N_18959,N_18891);
nand U19212 (N_19212,N_18919,N_18859);
nor U19213 (N_19213,N_18891,N_18953);
and U19214 (N_19214,N_18917,N_18972);
xor U19215 (N_19215,N_18979,N_18760);
xnor U19216 (N_19216,N_18771,N_18876);
nor U19217 (N_19217,N_18849,N_18766);
xor U19218 (N_19218,N_18774,N_18853);
or U19219 (N_19219,N_18872,N_18963);
nand U19220 (N_19220,N_18975,N_18886);
or U19221 (N_19221,N_18950,N_18901);
or U19222 (N_19222,N_18812,N_18919);
xor U19223 (N_19223,N_18778,N_18844);
xnor U19224 (N_19224,N_18862,N_18959);
and U19225 (N_19225,N_18926,N_18863);
nand U19226 (N_19226,N_18972,N_18998);
xor U19227 (N_19227,N_18792,N_18772);
nand U19228 (N_19228,N_18793,N_18995);
and U19229 (N_19229,N_18972,N_18896);
and U19230 (N_19230,N_18804,N_18877);
nor U19231 (N_19231,N_18887,N_18840);
nor U19232 (N_19232,N_18781,N_18972);
nor U19233 (N_19233,N_18815,N_18984);
and U19234 (N_19234,N_18794,N_18808);
nor U19235 (N_19235,N_18829,N_18942);
or U19236 (N_19236,N_18767,N_18845);
or U19237 (N_19237,N_18889,N_18807);
nor U19238 (N_19238,N_18887,N_18777);
xnor U19239 (N_19239,N_18831,N_18909);
nand U19240 (N_19240,N_18945,N_18917);
or U19241 (N_19241,N_18893,N_18963);
nand U19242 (N_19242,N_18882,N_18921);
nand U19243 (N_19243,N_18804,N_18836);
nor U19244 (N_19244,N_18797,N_18935);
or U19245 (N_19245,N_18821,N_18907);
and U19246 (N_19246,N_18826,N_18977);
nor U19247 (N_19247,N_18855,N_18839);
nand U19248 (N_19248,N_18769,N_18835);
nand U19249 (N_19249,N_18880,N_18806);
nor U19250 (N_19250,N_19075,N_19071);
nor U19251 (N_19251,N_19118,N_19058);
and U19252 (N_19252,N_19201,N_19054);
nand U19253 (N_19253,N_19027,N_19206);
xor U19254 (N_19254,N_19034,N_19060);
xor U19255 (N_19255,N_19164,N_19174);
nand U19256 (N_19256,N_19142,N_19045);
nor U19257 (N_19257,N_19148,N_19193);
xor U19258 (N_19258,N_19109,N_19159);
and U19259 (N_19259,N_19093,N_19098);
nand U19260 (N_19260,N_19237,N_19173);
and U19261 (N_19261,N_19223,N_19001);
or U19262 (N_19262,N_19009,N_19056);
or U19263 (N_19263,N_19111,N_19022);
or U19264 (N_19264,N_19171,N_19097);
nor U19265 (N_19265,N_19188,N_19089);
and U19266 (N_19266,N_19131,N_19051);
and U19267 (N_19267,N_19184,N_19062);
xnor U19268 (N_19268,N_19127,N_19140);
xor U19269 (N_19269,N_19208,N_19006);
nand U19270 (N_19270,N_19231,N_19108);
or U19271 (N_19271,N_19130,N_19096);
nand U19272 (N_19272,N_19014,N_19176);
and U19273 (N_19273,N_19037,N_19010);
nor U19274 (N_19274,N_19065,N_19139);
or U19275 (N_19275,N_19163,N_19038);
nand U19276 (N_19276,N_19030,N_19177);
and U19277 (N_19277,N_19221,N_19090);
and U19278 (N_19278,N_19248,N_19064);
and U19279 (N_19279,N_19079,N_19040);
and U19280 (N_19280,N_19123,N_19226);
nor U19281 (N_19281,N_19028,N_19198);
and U19282 (N_19282,N_19165,N_19175);
and U19283 (N_19283,N_19245,N_19247);
and U19284 (N_19284,N_19191,N_19172);
nand U19285 (N_19285,N_19134,N_19241);
or U19286 (N_19286,N_19166,N_19209);
or U19287 (N_19287,N_19026,N_19161);
nand U19288 (N_19288,N_19004,N_19049);
and U19289 (N_19289,N_19200,N_19136);
and U19290 (N_19290,N_19092,N_19194);
xnor U19291 (N_19291,N_19249,N_19196);
or U19292 (N_19292,N_19230,N_19013);
xnor U19293 (N_19293,N_19126,N_19146);
nand U19294 (N_19294,N_19207,N_19224);
nand U19295 (N_19295,N_19239,N_19063);
and U19296 (N_19296,N_19103,N_19059);
nand U19297 (N_19297,N_19082,N_19170);
xor U19298 (N_19298,N_19057,N_19039);
nand U19299 (N_19299,N_19212,N_19106);
or U19300 (N_19300,N_19035,N_19116);
nand U19301 (N_19301,N_19222,N_19102);
and U19302 (N_19302,N_19011,N_19135);
nor U19303 (N_19303,N_19023,N_19189);
nand U19304 (N_19304,N_19144,N_19086);
nor U19305 (N_19305,N_19029,N_19042);
xnor U19306 (N_19306,N_19167,N_19100);
or U19307 (N_19307,N_19156,N_19180);
xnor U19308 (N_19308,N_19073,N_19047);
and U19309 (N_19309,N_19185,N_19072);
nand U19310 (N_19310,N_19203,N_19181);
nor U19311 (N_19311,N_19149,N_19205);
or U19312 (N_19312,N_19032,N_19012);
and U19313 (N_19313,N_19067,N_19115);
xnor U19314 (N_19314,N_19019,N_19085);
and U19315 (N_19315,N_19202,N_19046);
nand U19316 (N_19316,N_19187,N_19124);
or U19317 (N_19317,N_19133,N_19055);
nand U19318 (N_19318,N_19007,N_19053);
nor U19319 (N_19319,N_19077,N_19017);
and U19320 (N_19320,N_19024,N_19122);
xnor U19321 (N_19321,N_19036,N_19217);
or U19322 (N_19322,N_19129,N_19190);
nand U19323 (N_19323,N_19061,N_19094);
xnor U19324 (N_19324,N_19016,N_19052);
nor U19325 (N_19325,N_19150,N_19138);
nor U19326 (N_19326,N_19033,N_19158);
or U19327 (N_19327,N_19025,N_19227);
nor U19328 (N_19328,N_19199,N_19168);
nand U19329 (N_19329,N_19084,N_19160);
or U19330 (N_19330,N_19216,N_19220);
xnor U19331 (N_19331,N_19232,N_19229);
nand U19332 (N_19332,N_19195,N_19143);
and U19333 (N_19333,N_19120,N_19151);
or U19334 (N_19334,N_19169,N_19066);
and U19335 (N_19335,N_19113,N_19182);
nor U19336 (N_19336,N_19048,N_19000);
nor U19337 (N_19337,N_19128,N_19099);
xnor U19338 (N_19338,N_19178,N_19020);
xnor U19339 (N_19339,N_19088,N_19008);
or U19340 (N_19340,N_19179,N_19132);
or U19341 (N_19341,N_19147,N_19080);
or U19342 (N_19342,N_19243,N_19117);
xor U19343 (N_19343,N_19070,N_19210);
nor U19344 (N_19344,N_19242,N_19018);
nand U19345 (N_19345,N_19246,N_19145);
or U19346 (N_19346,N_19068,N_19153);
or U19347 (N_19347,N_19238,N_19104);
and U19348 (N_19348,N_19081,N_19069);
nor U19349 (N_19349,N_19183,N_19107);
nand U19350 (N_19350,N_19215,N_19015);
and U19351 (N_19351,N_19044,N_19121);
nand U19352 (N_19352,N_19244,N_19112);
xor U19353 (N_19353,N_19095,N_19141);
nor U19354 (N_19354,N_19125,N_19091);
nor U19355 (N_19355,N_19234,N_19105);
xor U19356 (N_19356,N_19211,N_19114);
nand U19357 (N_19357,N_19228,N_19154);
nor U19358 (N_19358,N_19157,N_19087);
xnor U19359 (N_19359,N_19235,N_19119);
nand U19360 (N_19360,N_19197,N_19225);
xor U19361 (N_19361,N_19083,N_19204);
or U19362 (N_19362,N_19155,N_19137);
and U19363 (N_19363,N_19213,N_19002);
and U19364 (N_19364,N_19162,N_19076);
xor U19365 (N_19365,N_19214,N_19031);
or U19366 (N_19366,N_19240,N_19074);
xnor U19367 (N_19367,N_19041,N_19050);
nand U19368 (N_19368,N_19152,N_19003);
nor U19369 (N_19369,N_19101,N_19110);
nand U19370 (N_19370,N_19218,N_19005);
nor U19371 (N_19371,N_19021,N_19192);
and U19372 (N_19372,N_19043,N_19219);
xor U19373 (N_19373,N_19186,N_19078);
xnor U19374 (N_19374,N_19233,N_19236);
nor U19375 (N_19375,N_19060,N_19084);
or U19376 (N_19376,N_19150,N_19092);
or U19377 (N_19377,N_19155,N_19069);
nor U19378 (N_19378,N_19145,N_19087);
nor U19379 (N_19379,N_19013,N_19243);
or U19380 (N_19380,N_19063,N_19092);
or U19381 (N_19381,N_19032,N_19050);
xor U19382 (N_19382,N_19078,N_19194);
xor U19383 (N_19383,N_19222,N_19214);
or U19384 (N_19384,N_19083,N_19087);
xnor U19385 (N_19385,N_19045,N_19169);
nand U19386 (N_19386,N_19193,N_19141);
xnor U19387 (N_19387,N_19248,N_19227);
xnor U19388 (N_19388,N_19007,N_19113);
nor U19389 (N_19389,N_19118,N_19114);
xor U19390 (N_19390,N_19176,N_19161);
nor U19391 (N_19391,N_19077,N_19079);
and U19392 (N_19392,N_19067,N_19037);
nand U19393 (N_19393,N_19156,N_19197);
xor U19394 (N_19394,N_19195,N_19222);
nor U19395 (N_19395,N_19042,N_19027);
or U19396 (N_19396,N_19185,N_19097);
nor U19397 (N_19397,N_19111,N_19165);
nand U19398 (N_19398,N_19062,N_19019);
xnor U19399 (N_19399,N_19022,N_19076);
xor U19400 (N_19400,N_19014,N_19109);
or U19401 (N_19401,N_19180,N_19048);
and U19402 (N_19402,N_19087,N_19194);
or U19403 (N_19403,N_19101,N_19237);
xor U19404 (N_19404,N_19115,N_19216);
nor U19405 (N_19405,N_19025,N_19110);
or U19406 (N_19406,N_19083,N_19217);
xor U19407 (N_19407,N_19118,N_19199);
or U19408 (N_19408,N_19190,N_19148);
xnor U19409 (N_19409,N_19099,N_19149);
xnor U19410 (N_19410,N_19189,N_19206);
or U19411 (N_19411,N_19237,N_19091);
nand U19412 (N_19412,N_19096,N_19038);
nand U19413 (N_19413,N_19207,N_19082);
xor U19414 (N_19414,N_19226,N_19146);
nor U19415 (N_19415,N_19130,N_19055);
xnor U19416 (N_19416,N_19146,N_19113);
or U19417 (N_19417,N_19093,N_19068);
or U19418 (N_19418,N_19003,N_19040);
nor U19419 (N_19419,N_19194,N_19064);
nand U19420 (N_19420,N_19167,N_19183);
or U19421 (N_19421,N_19221,N_19072);
nor U19422 (N_19422,N_19055,N_19127);
nand U19423 (N_19423,N_19169,N_19209);
and U19424 (N_19424,N_19133,N_19201);
xnor U19425 (N_19425,N_19146,N_19078);
or U19426 (N_19426,N_19007,N_19116);
nand U19427 (N_19427,N_19076,N_19175);
xnor U19428 (N_19428,N_19147,N_19093);
or U19429 (N_19429,N_19234,N_19047);
or U19430 (N_19430,N_19238,N_19010);
nand U19431 (N_19431,N_19090,N_19115);
and U19432 (N_19432,N_19218,N_19091);
nor U19433 (N_19433,N_19081,N_19040);
and U19434 (N_19434,N_19019,N_19068);
xnor U19435 (N_19435,N_19199,N_19131);
nor U19436 (N_19436,N_19138,N_19029);
nand U19437 (N_19437,N_19028,N_19102);
and U19438 (N_19438,N_19175,N_19213);
xnor U19439 (N_19439,N_19155,N_19082);
and U19440 (N_19440,N_19038,N_19102);
nand U19441 (N_19441,N_19056,N_19006);
or U19442 (N_19442,N_19098,N_19050);
nor U19443 (N_19443,N_19121,N_19107);
xnor U19444 (N_19444,N_19005,N_19139);
nor U19445 (N_19445,N_19043,N_19004);
nor U19446 (N_19446,N_19039,N_19134);
and U19447 (N_19447,N_19192,N_19075);
xnor U19448 (N_19448,N_19121,N_19096);
or U19449 (N_19449,N_19183,N_19095);
and U19450 (N_19450,N_19131,N_19087);
nor U19451 (N_19451,N_19113,N_19143);
or U19452 (N_19452,N_19222,N_19154);
and U19453 (N_19453,N_19247,N_19175);
or U19454 (N_19454,N_19066,N_19144);
xnor U19455 (N_19455,N_19078,N_19133);
nand U19456 (N_19456,N_19011,N_19067);
nand U19457 (N_19457,N_19103,N_19120);
nand U19458 (N_19458,N_19182,N_19189);
and U19459 (N_19459,N_19032,N_19092);
and U19460 (N_19460,N_19083,N_19054);
nor U19461 (N_19461,N_19221,N_19211);
or U19462 (N_19462,N_19068,N_19077);
or U19463 (N_19463,N_19130,N_19192);
and U19464 (N_19464,N_19001,N_19144);
nor U19465 (N_19465,N_19234,N_19166);
nor U19466 (N_19466,N_19217,N_19219);
xnor U19467 (N_19467,N_19006,N_19247);
nand U19468 (N_19468,N_19082,N_19037);
and U19469 (N_19469,N_19232,N_19188);
xnor U19470 (N_19470,N_19100,N_19195);
and U19471 (N_19471,N_19069,N_19132);
nand U19472 (N_19472,N_19232,N_19040);
xor U19473 (N_19473,N_19002,N_19056);
nand U19474 (N_19474,N_19137,N_19147);
or U19475 (N_19475,N_19035,N_19217);
nand U19476 (N_19476,N_19167,N_19044);
nand U19477 (N_19477,N_19134,N_19026);
and U19478 (N_19478,N_19062,N_19172);
xor U19479 (N_19479,N_19049,N_19042);
or U19480 (N_19480,N_19157,N_19200);
xnor U19481 (N_19481,N_19099,N_19058);
or U19482 (N_19482,N_19116,N_19166);
nor U19483 (N_19483,N_19073,N_19058);
nand U19484 (N_19484,N_19199,N_19027);
and U19485 (N_19485,N_19048,N_19018);
or U19486 (N_19486,N_19039,N_19012);
or U19487 (N_19487,N_19063,N_19166);
xnor U19488 (N_19488,N_19138,N_19153);
nor U19489 (N_19489,N_19196,N_19146);
xnor U19490 (N_19490,N_19210,N_19240);
nor U19491 (N_19491,N_19236,N_19159);
nor U19492 (N_19492,N_19035,N_19208);
xnor U19493 (N_19493,N_19192,N_19099);
or U19494 (N_19494,N_19097,N_19245);
nor U19495 (N_19495,N_19182,N_19107);
or U19496 (N_19496,N_19139,N_19104);
nor U19497 (N_19497,N_19196,N_19051);
xnor U19498 (N_19498,N_19000,N_19163);
or U19499 (N_19499,N_19182,N_19160);
xnor U19500 (N_19500,N_19408,N_19290);
nor U19501 (N_19501,N_19334,N_19265);
and U19502 (N_19502,N_19365,N_19450);
or U19503 (N_19503,N_19379,N_19484);
or U19504 (N_19504,N_19264,N_19456);
or U19505 (N_19505,N_19444,N_19493);
nand U19506 (N_19506,N_19439,N_19445);
nor U19507 (N_19507,N_19321,N_19345);
and U19508 (N_19508,N_19342,N_19405);
nand U19509 (N_19509,N_19354,N_19318);
and U19510 (N_19510,N_19384,N_19259);
nand U19511 (N_19511,N_19457,N_19327);
and U19512 (N_19512,N_19383,N_19355);
nor U19513 (N_19513,N_19440,N_19417);
or U19514 (N_19514,N_19428,N_19364);
or U19515 (N_19515,N_19304,N_19394);
and U19516 (N_19516,N_19302,N_19407);
nor U19517 (N_19517,N_19443,N_19399);
or U19518 (N_19518,N_19294,N_19476);
nand U19519 (N_19519,N_19330,N_19402);
and U19520 (N_19520,N_19336,N_19386);
and U19521 (N_19521,N_19404,N_19472);
and U19522 (N_19522,N_19299,N_19397);
nand U19523 (N_19523,N_19328,N_19455);
xnor U19524 (N_19524,N_19357,N_19351);
nand U19525 (N_19525,N_19269,N_19296);
and U19526 (N_19526,N_19250,N_19260);
nor U19527 (N_19527,N_19311,N_19284);
and U19528 (N_19528,N_19436,N_19487);
xnor U19529 (N_19529,N_19434,N_19385);
nor U19530 (N_19530,N_19344,N_19275);
nand U19531 (N_19531,N_19374,N_19261);
or U19532 (N_19532,N_19368,N_19341);
nand U19533 (N_19533,N_19310,N_19409);
nand U19534 (N_19534,N_19497,N_19286);
xor U19535 (N_19535,N_19317,N_19361);
xnor U19536 (N_19536,N_19297,N_19346);
nor U19537 (N_19537,N_19420,N_19413);
or U19538 (N_19538,N_19438,N_19414);
nand U19539 (N_19539,N_19427,N_19422);
xnor U19540 (N_19540,N_19398,N_19347);
xor U19541 (N_19541,N_19274,N_19461);
nand U19542 (N_19542,N_19271,N_19277);
xor U19543 (N_19543,N_19415,N_19481);
nand U19544 (N_19544,N_19370,N_19367);
or U19545 (N_19545,N_19449,N_19483);
xor U19546 (N_19546,N_19293,N_19267);
nand U19547 (N_19547,N_19359,N_19442);
and U19548 (N_19548,N_19431,N_19257);
or U19549 (N_19549,N_19363,N_19320);
nand U19550 (N_19550,N_19362,N_19464);
nor U19551 (N_19551,N_19391,N_19378);
nor U19552 (N_19552,N_19496,N_19376);
or U19553 (N_19553,N_19447,N_19392);
xor U19554 (N_19554,N_19406,N_19278);
xnor U19555 (N_19555,N_19465,N_19446);
nor U19556 (N_19556,N_19255,N_19441);
xnor U19557 (N_19557,N_19498,N_19463);
nand U19558 (N_19558,N_19470,N_19393);
nor U19559 (N_19559,N_19412,N_19479);
nor U19560 (N_19560,N_19469,N_19279);
nand U19561 (N_19561,N_19306,N_19390);
and U19562 (N_19562,N_19256,N_19358);
and U19563 (N_19563,N_19421,N_19262);
or U19564 (N_19564,N_19432,N_19331);
nor U19565 (N_19565,N_19466,N_19338);
xnor U19566 (N_19566,N_19282,N_19325);
xor U19567 (N_19567,N_19473,N_19478);
or U19568 (N_19568,N_19480,N_19486);
or U19569 (N_19569,N_19426,N_19488);
xor U19570 (N_19570,N_19288,N_19356);
xor U19571 (N_19571,N_19353,N_19252);
nor U19572 (N_19572,N_19389,N_19263);
nand U19573 (N_19573,N_19396,N_19322);
nand U19574 (N_19574,N_19454,N_19403);
nor U19575 (N_19575,N_19430,N_19462);
nor U19576 (N_19576,N_19291,N_19416);
nor U19577 (N_19577,N_19329,N_19301);
nand U19578 (N_19578,N_19253,N_19380);
and U19579 (N_19579,N_19268,N_19352);
xnor U19580 (N_19580,N_19468,N_19401);
or U19581 (N_19581,N_19369,N_19307);
nor U19582 (N_19582,N_19276,N_19495);
nor U19583 (N_19583,N_19411,N_19343);
xor U19584 (N_19584,N_19305,N_19283);
xor U19585 (N_19585,N_19339,N_19400);
and U19586 (N_19586,N_19308,N_19323);
xor U19587 (N_19587,N_19435,N_19313);
xor U19588 (N_19588,N_19335,N_19437);
nand U19589 (N_19589,N_19451,N_19314);
nor U19590 (N_19590,N_19485,N_19272);
or U19591 (N_19591,N_19387,N_19377);
xnor U19592 (N_19592,N_19492,N_19375);
or U19593 (N_19593,N_19348,N_19489);
xor U19594 (N_19594,N_19303,N_19423);
or U19595 (N_19595,N_19295,N_19366);
and U19596 (N_19596,N_19425,N_19281);
xor U19597 (N_19597,N_19273,N_19251);
nor U19598 (N_19598,N_19324,N_19337);
xnor U19599 (N_19599,N_19373,N_19258);
or U19600 (N_19600,N_19319,N_19381);
nand U19601 (N_19601,N_19452,N_19289);
xor U19602 (N_19602,N_19309,N_19475);
or U19603 (N_19603,N_19482,N_19418);
nor U19604 (N_19604,N_19471,N_19448);
and U19605 (N_19605,N_19292,N_19395);
and U19606 (N_19606,N_19349,N_19494);
xnor U19607 (N_19607,N_19315,N_19340);
nor U19608 (N_19608,N_19388,N_19499);
nand U19609 (N_19609,N_19467,N_19490);
xnor U19610 (N_19610,N_19419,N_19326);
nand U19611 (N_19611,N_19266,N_19410);
xnor U19612 (N_19612,N_19371,N_19491);
and U19613 (N_19613,N_19360,N_19458);
xor U19614 (N_19614,N_19298,N_19270);
or U19615 (N_19615,N_19382,N_19372);
nand U19616 (N_19616,N_19316,N_19254);
or U19617 (N_19617,N_19459,N_19429);
or U19618 (N_19618,N_19287,N_19424);
xnor U19619 (N_19619,N_19285,N_19477);
and U19620 (N_19620,N_19280,N_19453);
nor U19621 (N_19621,N_19474,N_19350);
or U19622 (N_19622,N_19332,N_19460);
or U19623 (N_19623,N_19312,N_19333);
nand U19624 (N_19624,N_19300,N_19433);
xnor U19625 (N_19625,N_19462,N_19372);
nand U19626 (N_19626,N_19352,N_19360);
and U19627 (N_19627,N_19455,N_19321);
and U19628 (N_19628,N_19310,N_19313);
nand U19629 (N_19629,N_19497,N_19418);
xnor U19630 (N_19630,N_19318,N_19477);
nand U19631 (N_19631,N_19262,N_19414);
nor U19632 (N_19632,N_19342,N_19489);
xnor U19633 (N_19633,N_19436,N_19401);
and U19634 (N_19634,N_19300,N_19362);
nor U19635 (N_19635,N_19368,N_19275);
and U19636 (N_19636,N_19370,N_19383);
or U19637 (N_19637,N_19470,N_19423);
nand U19638 (N_19638,N_19282,N_19483);
xor U19639 (N_19639,N_19407,N_19290);
and U19640 (N_19640,N_19316,N_19294);
and U19641 (N_19641,N_19296,N_19361);
xor U19642 (N_19642,N_19300,N_19429);
or U19643 (N_19643,N_19476,N_19343);
and U19644 (N_19644,N_19354,N_19465);
or U19645 (N_19645,N_19337,N_19262);
nand U19646 (N_19646,N_19296,N_19252);
and U19647 (N_19647,N_19336,N_19371);
nor U19648 (N_19648,N_19430,N_19444);
or U19649 (N_19649,N_19292,N_19484);
or U19650 (N_19650,N_19405,N_19287);
and U19651 (N_19651,N_19393,N_19479);
or U19652 (N_19652,N_19341,N_19378);
nand U19653 (N_19653,N_19447,N_19473);
xnor U19654 (N_19654,N_19391,N_19332);
and U19655 (N_19655,N_19315,N_19299);
nand U19656 (N_19656,N_19412,N_19252);
xnor U19657 (N_19657,N_19319,N_19375);
nand U19658 (N_19658,N_19322,N_19467);
xor U19659 (N_19659,N_19487,N_19279);
xnor U19660 (N_19660,N_19278,N_19315);
nor U19661 (N_19661,N_19318,N_19268);
xor U19662 (N_19662,N_19488,N_19350);
nor U19663 (N_19663,N_19399,N_19431);
xnor U19664 (N_19664,N_19477,N_19406);
or U19665 (N_19665,N_19271,N_19283);
nand U19666 (N_19666,N_19344,N_19380);
or U19667 (N_19667,N_19331,N_19384);
nor U19668 (N_19668,N_19289,N_19443);
or U19669 (N_19669,N_19428,N_19288);
or U19670 (N_19670,N_19472,N_19303);
or U19671 (N_19671,N_19441,N_19304);
xor U19672 (N_19672,N_19253,N_19322);
or U19673 (N_19673,N_19263,N_19362);
xnor U19674 (N_19674,N_19398,N_19297);
xor U19675 (N_19675,N_19358,N_19312);
and U19676 (N_19676,N_19279,N_19433);
nor U19677 (N_19677,N_19265,N_19485);
and U19678 (N_19678,N_19474,N_19313);
nor U19679 (N_19679,N_19364,N_19444);
xor U19680 (N_19680,N_19466,N_19485);
nand U19681 (N_19681,N_19284,N_19344);
nor U19682 (N_19682,N_19481,N_19263);
or U19683 (N_19683,N_19368,N_19430);
xnor U19684 (N_19684,N_19367,N_19356);
nor U19685 (N_19685,N_19498,N_19299);
xor U19686 (N_19686,N_19388,N_19471);
nor U19687 (N_19687,N_19375,N_19436);
nand U19688 (N_19688,N_19398,N_19456);
xor U19689 (N_19689,N_19279,N_19461);
nor U19690 (N_19690,N_19499,N_19369);
nand U19691 (N_19691,N_19417,N_19253);
or U19692 (N_19692,N_19310,N_19402);
nor U19693 (N_19693,N_19441,N_19298);
nor U19694 (N_19694,N_19451,N_19482);
nand U19695 (N_19695,N_19298,N_19274);
nand U19696 (N_19696,N_19473,N_19448);
nor U19697 (N_19697,N_19401,N_19346);
and U19698 (N_19698,N_19445,N_19360);
nand U19699 (N_19699,N_19268,N_19266);
xnor U19700 (N_19700,N_19405,N_19279);
nor U19701 (N_19701,N_19403,N_19467);
or U19702 (N_19702,N_19406,N_19326);
and U19703 (N_19703,N_19450,N_19474);
xnor U19704 (N_19704,N_19422,N_19328);
nor U19705 (N_19705,N_19400,N_19432);
nor U19706 (N_19706,N_19446,N_19267);
xnor U19707 (N_19707,N_19320,N_19420);
or U19708 (N_19708,N_19402,N_19342);
nand U19709 (N_19709,N_19445,N_19260);
or U19710 (N_19710,N_19310,N_19343);
nor U19711 (N_19711,N_19319,N_19348);
or U19712 (N_19712,N_19267,N_19380);
xor U19713 (N_19713,N_19381,N_19499);
and U19714 (N_19714,N_19428,N_19472);
nor U19715 (N_19715,N_19429,N_19302);
or U19716 (N_19716,N_19255,N_19298);
xnor U19717 (N_19717,N_19256,N_19448);
nand U19718 (N_19718,N_19388,N_19418);
xor U19719 (N_19719,N_19393,N_19357);
xnor U19720 (N_19720,N_19466,N_19266);
and U19721 (N_19721,N_19425,N_19277);
nand U19722 (N_19722,N_19429,N_19497);
or U19723 (N_19723,N_19438,N_19418);
nor U19724 (N_19724,N_19294,N_19498);
xnor U19725 (N_19725,N_19273,N_19415);
or U19726 (N_19726,N_19314,N_19265);
or U19727 (N_19727,N_19422,N_19338);
nand U19728 (N_19728,N_19292,N_19266);
or U19729 (N_19729,N_19312,N_19394);
xor U19730 (N_19730,N_19319,N_19302);
and U19731 (N_19731,N_19325,N_19481);
or U19732 (N_19732,N_19395,N_19428);
xnor U19733 (N_19733,N_19384,N_19340);
or U19734 (N_19734,N_19317,N_19427);
xnor U19735 (N_19735,N_19447,N_19390);
or U19736 (N_19736,N_19252,N_19323);
and U19737 (N_19737,N_19461,N_19401);
xnor U19738 (N_19738,N_19277,N_19360);
and U19739 (N_19739,N_19452,N_19459);
xor U19740 (N_19740,N_19476,N_19344);
and U19741 (N_19741,N_19421,N_19393);
and U19742 (N_19742,N_19390,N_19364);
and U19743 (N_19743,N_19283,N_19298);
or U19744 (N_19744,N_19429,N_19252);
nand U19745 (N_19745,N_19334,N_19350);
nor U19746 (N_19746,N_19252,N_19371);
or U19747 (N_19747,N_19337,N_19490);
nor U19748 (N_19748,N_19272,N_19326);
and U19749 (N_19749,N_19374,N_19434);
nor U19750 (N_19750,N_19591,N_19725);
nand U19751 (N_19751,N_19695,N_19631);
nand U19752 (N_19752,N_19506,N_19696);
nand U19753 (N_19753,N_19686,N_19613);
or U19754 (N_19754,N_19539,N_19688);
xor U19755 (N_19755,N_19660,N_19608);
xnor U19756 (N_19756,N_19709,N_19707);
and U19757 (N_19757,N_19656,N_19558);
xor U19758 (N_19758,N_19627,N_19690);
nor U19759 (N_19759,N_19685,N_19502);
xnor U19760 (N_19760,N_19535,N_19645);
xnor U19761 (N_19761,N_19635,N_19720);
nand U19762 (N_19762,N_19700,N_19677);
and U19763 (N_19763,N_19593,N_19714);
nand U19764 (N_19764,N_19657,N_19702);
and U19765 (N_19765,N_19723,N_19745);
nor U19766 (N_19766,N_19743,N_19708);
nand U19767 (N_19767,N_19546,N_19553);
nor U19768 (N_19768,N_19733,N_19736);
nor U19769 (N_19769,N_19640,N_19730);
xnor U19770 (N_19770,N_19572,N_19687);
xor U19771 (N_19771,N_19523,N_19655);
xnor U19772 (N_19772,N_19620,N_19567);
nor U19773 (N_19773,N_19564,N_19654);
nand U19774 (N_19774,N_19525,N_19632);
nor U19775 (N_19775,N_19548,N_19671);
or U19776 (N_19776,N_19512,N_19735);
nand U19777 (N_19777,N_19536,N_19526);
nand U19778 (N_19778,N_19500,N_19592);
or U19779 (N_19779,N_19747,N_19665);
xnor U19780 (N_19780,N_19565,N_19749);
nand U19781 (N_19781,N_19594,N_19722);
or U19782 (N_19782,N_19547,N_19522);
and U19783 (N_19783,N_19584,N_19568);
xnor U19784 (N_19784,N_19617,N_19544);
nand U19785 (N_19785,N_19555,N_19721);
nor U19786 (N_19786,N_19596,N_19606);
nor U19787 (N_19787,N_19663,N_19744);
nand U19788 (N_19788,N_19728,N_19740);
and U19789 (N_19789,N_19543,N_19549);
or U19790 (N_19790,N_19586,N_19646);
or U19791 (N_19791,N_19521,N_19604);
nor U19792 (N_19792,N_19731,N_19524);
nand U19793 (N_19793,N_19724,N_19541);
nand U19794 (N_19794,N_19533,N_19699);
and U19795 (N_19795,N_19621,N_19674);
and U19796 (N_19796,N_19559,N_19662);
xor U19797 (N_19797,N_19692,N_19636);
xor U19798 (N_19798,N_19659,N_19563);
or U19799 (N_19799,N_19551,N_19597);
xor U19800 (N_19800,N_19711,N_19668);
or U19801 (N_19801,N_19732,N_19644);
or U19802 (N_19802,N_19667,N_19738);
and U19803 (N_19803,N_19746,N_19530);
nand U19804 (N_19804,N_19516,N_19611);
nor U19805 (N_19805,N_19737,N_19628);
and U19806 (N_19806,N_19580,N_19748);
xor U19807 (N_19807,N_19630,N_19557);
xnor U19808 (N_19808,N_19566,N_19508);
and U19809 (N_19809,N_19504,N_19562);
xor U19810 (N_19810,N_19518,N_19639);
nor U19811 (N_19811,N_19583,N_19710);
and U19812 (N_19812,N_19715,N_19704);
nor U19813 (N_19813,N_19588,N_19673);
and U19814 (N_19814,N_19560,N_19573);
nand U19815 (N_19815,N_19581,N_19609);
nand U19816 (N_19816,N_19734,N_19509);
or U19817 (N_19817,N_19589,N_19625);
or U19818 (N_19818,N_19698,N_19545);
xnor U19819 (N_19819,N_19712,N_19612);
and U19820 (N_19820,N_19716,N_19706);
nand U19821 (N_19821,N_19614,N_19653);
or U19822 (N_19822,N_19742,N_19629);
and U19823 (N_19823,N_19529,N_19624);
nor U19824 (N_19824,N_19561,N_19507);
nand U19825 (N_19825,N_19683,N_19651);
and U19826 (N_19826,N_19729,N_19664);
or U19827 (N_19827,N_19610,N_19600);
or U19828 (N_19828,N_19542,N_19576);
nor U19829 (N_19829,N_19701,N_19517);
nor U19830 (N_19830,N_19575,N_19638);
xnor U19831 (N_19831,N_19574,N_19510);
nor U19832 (N_19832,N_19626,N_19669);
nand U19833 (N_19833,N_19577,N_19672);
and U19834 (N_19834,N_19684,N_19511);
and U19835 (N_19835,N_19676,N_19605);
xnor U19836 (N_19836,N_19534,N_19717);
nor U19837 (N_19837,N_19554,N_19719);
xor U19838 (N_19838,N_19595,N_19598);
or U19839 (N_19839,N_19615,N_19505);
nand U19840 (N_19840,N_19515,N_19649);
xnor U19841 (N_19841,N_19528,N_19680);
and U19842 (N_19842,N_19599,N_19643);
and U19843 (N_19843,N_19666,N_19650);
nand U19844 (N_19844,N_19520,N_19691);
nand U19845 (N_19845,N_19634,N_19607);
and U19846 (N_19846,N_19718,N_19622);
nand U19847 (N_19847,N_19503,N_19532);
xor U19848 (N_19848,N_19726,N_19585);
xor U19849 (N_19849,N_19582,N_19675);
and U19850 (N_19850,N_19519,N_19647);
nand U19851 (N_19851,N_19616,N_19623);
nand U19852 (N_19852,N_19578,N_19697);
nand U19853 (N_19853,N_19679,N_19703);
nor U19854 (N_19854,N_19556,N_19538);
nand U19855 (N_19855,N_19540,N_19641);
nor U19856 (N_19856,N_19571,N_19642);
and U19857 (N_19857,N_19661,N_19601);
xnor U19858 (N_19858,N_19579,N_19570);
nor U19859 (N_19859,N_19527,N_19514);
and U19860 (N_19860,N_19658,N_19741);
and U19861 (N_19861,N_19587,N_19689);
or U19862 (N_19862,N_19569,N_19682);
or U19863 (N_19863,N_19693,N_19633);
or U19864 (N_19864,N_19531,N_19652);
and U19865 (N_19865,N_19681,N_19739);
nand U19866 (N_19866,N_19727,N_19619);
xnor U19867 (N_19867,N_19705,N_19637);
xnor U19868 (N_19868,N_19670,N_19694);
or U19869 (N_19869,N_19603,N_19552);
nand U19870 (N_19870,N_19602,N_19550);
and U19871 (N_19871,N_19501,N_19618);
and U19872 (N_19872,N_19513,N_19590);
nor U19873 (N_19873,N_19678,N_19713);
nor U19874 (N_19874,N_19537,N_19648);
nor U19875 (N_19875,N_19553,N_19709);
nand U19876 (N_19876,N_19725,N_19593);
nand U19877 (N_19877,N_19640,N_19541);
and U19878 (N_19878,N_19527,N_19692);
nor U19879 (N_19879,N_19507,N_19698);
xnor U19880 (N_19880,N_19540,N_19587);
nand U19881 (N_19881,N_19581,N_19691);
or U19882 (N_19882,N_19542,N_19525);
and U19883 (N_19883,N_19579,N_19629);
xnor U19884 (N_19884,N_19587,N_19521);
nand U19885 (N_19885,N_19522,N_19508);
or U19886 (N_19886,N_19594,N_19728);
and U19887 (N_19887,N_19678,N_19544);
xor U19888 (N_19888,N_19720,N_19563);
nand U19889 (N_19889,N_19525,N_19725);
and U19890 (N_19890,N_19738,N_19740);
nand U19891 (N_19891,N_19512,N_19600);
and U19892 (N_19892,N_19545,N_19623);
or U19893 (N_19893,N_19717,N_19571);
nand U19894 (N_19894,N_19506,N_19593);
or U19895 (N_19895,N_19564,N_19615);
nand U19896 (N_19896,N_19564,N_19734);
xnor U19897 (N_19897,N_19587,N_19596);
nor U19898 (N_19898,N_19724,N_19741);
and U19899 (N_19899,N_19558,N_19746);
or U19900 (N_19900,N_19702,N_19504);
or U19901 (N_19901,N_19586,N_19730);
nor U19902 (N_19902,N_19667,N_19602);
xnor U19903 (N_19903,N_19683,N_19537);
nand U19904 (N_19904,N_19590,N_19514);
and U19905 (N_19905,N_19743,N_19535);
nand U19906 (N_19906,N_19626,N_19651);
or U19907 (N_19907,N_19649,N_19607);
xor U19908 (N_19908,N_19503,N_19655);
and U19909 (N_19909,N_19690,N_19632);
and U19910 (N_19910,N_19664,N_19632);
nand U19911 (N_19911,N_19522,N_19576);
xnor U19912 (N_19912,N_19532,N_19727);
nor U19913 (N_19913,N_19609,N_19655);
or U19914 (N_19914,N_19608,N_19526);
or U19915 (N_19915,N_19745,N_19692);
nor U19916 (N_19916,N_19738,N_19605);
and U19917 (N_19917,N_19665,N_19645);
xnor U19918 (N_19918,N_19704,N_19613);
or U19919 (N_19919,N_19733,N_19638);
nor U19920 (N_19920,N_19578,N_19549);
nand U19921 (N_19921,N_19724,N_19733);
nand U19922 (N_19922,N_19542,N_19684);
nand U19923 (N_19923,N_19523,N_19685);
and U19924 (N_19924,N_19596,N_19649);
nand U19925 (N_19925,N_19669,N_19618);
or U19926 (N_19926,N_19571,N_19728);
xor U19927 (N_19927,N_19684,N_19640);
or U19928 (N_19928,N_19696,N_19732);
and U19929 (N_19929,N_19584,N_19508);
nor U19930 (N_19930,N_19610,N_19556);
xor U19931 (N_19931,N_19582,N_19655);
xor U19932 (N_19932,N_19700,N_19549);
nand U19933 (N_19933,N_19610,N_19637);
and U19934 (N_19934,N_19716,N_19554);
and U19935 (N_19935,N_19737,N_19746);
nand U19936 (N_19936,N_19675,N_19524);
xnor U19937 (N_19937,N_19717,N_19597);
and U19938 (N_19938,N_19683,N_19507);
nand U19939 (N_19939,N_19666,N_19536);
xor U19940 (N_19940,N_19694,N_19652);
nand U19941 (N_19941,N_19599,N_19606);
and U19942 (N_19942,N_19679,N_19733);
or U19943 (N_19943,N_19585,N_19744);
and U19944 (N_19944,N_19677,N_19627);
and U19945 (N_19945,N_19654,N_19676);
and U19946 (N_19946,N_19501,N_19730);
or U19947 (N_19947,N_19657,N_19527);
nor U19948 (N_19948,N_19568,N_19605);
and U19949 (N_19949,N_19603,N_19533);
and U19950 (N_19950,N_19676,N_19556);
nor U19951 (N_19951,N_19643,N_19627);
xnor U19952 (N_19952,N_19709,N_19737);
and U19953 (N_19953,N_19554,N_19683);
nand U19954 (N_19954,N_19586,N_19561);
and U19955 (N_19955,N_19630,N_19681);
xnor U19956 (N_19956,N_19666,N_19623);
or U19957 (N_19957,N_19569,N_19675);
nor U19958 (N_19958,N_19690,N_19540);
xor U19959 (N_19959,N_19619,N_19721);
or U19960 (N_19960,N_19580,N_19521);
xnor U19961 (N_19961,N_19737,N_19710);
xnor U19962 (N_19962,N_19640,N_19522);
nor U19963 (N_19963,N_19634,N_19729);
nor U19964 (N_19964,N_19524,N_19554);
xor U19965 (N_19965,N_19587,N_19537);
xnor U19966 (N_19966,N_19608,N_19720);
nand U19967 (N_19967,N_19617,N_19540);
or U19968 (N_19968,N_19561,N_19532);
nand U19969 (N_19969,N_19660,N_19634);
or U19970 (N_19970,N_19722,N_19542);
and U19971 (N_19971,N_19678,N_19559);
and U19972 (N_19972,N_19607,N_19699);
nor U19973 (N_19973,N_19523,N_19659);
nand U19974 (N_19974,N_19593,N_19612);
xnor U19975 (N_19975,N_19639,N_19644);
nor U19976 (N_19976,N_19583,N_19505);
nand U19977 (N_19977,N_19580,N_19578);
and U19978 (N_19978,N_19741,N_19655);
xnor U19979 (N_19979,N_19642,N_19508);
xnor U19980 (N_19980,N_19663,N_19725);
nor U19981 (N_19981,N_19591,N_19645);
xor U19982 (N_19982,N_19565,N_19600);
and U19983 (N_19983,N_19740,N_19575);
nand U19984 (N_19984,N_19618,N_19680);
and U19985 (N_19985,N_19561,N_19706);
xor U19986 (N_19986,N_19683,N_19519);
nand U19987 (N_19987,N_19696,N_19671);
and U19988 (N_19988,N_19745,N_19733);
xor U19989 (N_19989,N_19730,N_19736);
nand U19990 (N_19990,N_19705,N_19549);
and U19991 (N_19991,N_19630,N_19607);
nand U19992 (N_19992,N_19589,N_19515);
or U19993 (N_19993,N_19573,N_19743);
xnor U19994 (N_19994,N_19615,N_19572);
xor U19995 (N_19995,N_19619,N_19674);
xnor U19996 (N_19996,N_19593,N_19695);
nand U19997 (N_19997,N_19640,N_19693);
and U19998 (N_19998,N_19511,N_19553);
xor U19999 (N_19999,N_19596,N_19617);
and U20000 (N_20000,N_19961,N_19787);
nor U20001 (N_20001,N_19758,N_19969);
and U20002 (N_20002,N_19899,N_19893);
nor U20003 (N_20003,N_19793,N_19892);
nor U20004 (N_20004,N_19950,N_19777);
xnor U20005 (N_20005,N_19873,N_19866);
xnor U20006 (N_20006,N_19874,N_19806);
nor U20007 (N_20007,N_19759,N_19953);
and U20008 (N_20008,N_19816,N_19859);
nand U20009 (N_20009,N_19924,N_19905);
nand U20010 (N_20010,N_19811,N_19978);
nand U20011 (N_20011,N_19938,N_19926);
and U20012 (N_20012,N_19987,N_19890);
or U20013 (N_20013,N_19923,N_19869);
xor U20014 (N_20014,N_19982,N_19846);
nand U20015 (N_20015,N_19775,N_19943);
nand U20016 (N_20016,N_19805,N_19959);
nor U20017 (N_20017,N_19891,N_19855);
or U20018 (N_20018,N_19827,N_19940);
or U20019 (N_20019,N_19954,N_19886);
nand U20020 (N_20020,N_19754,N_19861);
or U20021 (N_20021,N_19776,N_19825);
or U20022 (N_20022,N_19856,N_19962);
nor U20023 (N_20023,N_19770,N_19809);
nor U20024 (N_20024,N_19966,N_19843);
nor U20025 (N_20025,N_19997,N_19860);
xor U20026 (N_20026,N_19983,N_19965);
or U20027 (N_20027,N_19884,N_19837);
and U20028 (N_20028,N_19850,N_19753);
or U20029 (N_20029,N_19974,N_19995);
and U20030 (N_20030,N_19931,N_19824);
and U20031 (N_20031,N_19799,N_19922);
and U20032 (N_20032,N_19885,N_19844);
nor U20033 (N_20033,N_19852,N_19839);
and U20034 (N_20034,N_19956,N_19761);
and U20035 (N_20035,N_19882,N_19985);
and U20036 (N_20036,N_19848,N_19797);
or U20037 (N_20037,N_19796,N_19771);
nand U20038 (N_20038,N_19750,N_19911);
nor U20039 (N_20039,N_19802,N_19894);
and U20040 (N_20040,N_19916,N_19834);
and U20041 (N_20041,N_19845,N_19981);
and U20042 (N_20042,N_19773,N_19900);
nand U20043 (N_20043,N_19889,N_19989);
xor U20044 (N_20044,N_19986,N_19783);
xor U20045 (N_20045,N_19851,N_19919);
xor U20046 (N_20046,N_19990,N_19871);
nand U20047 (N_20047,N_19790,N_19947);
or U20048 (N_20048,N_19785,N_19842);
xnor U20049 (N_20049,N_19883,N_19779);
nand U20050 (N_20050,N_19898,N_19774);
nor U20051 (N_20051,N_19766,N_19801);
or U20052 (N_20052,N_19955,N_19870);
nand U20053 (N_20053,N_19991,N_19765);
nor U20054 (N_20054,N_19833,N_19863);
nor U20055 (N_20055,N_19904,N_19936);
xor U20056 (N_20056,N_19928,N_19907);
xnor U20057 (N_20057,N_19935,N_19920);
nand U20058 (N_20058,N_19820,N_19791);
and U20059 (N_20059,N_19930,N_19914);
nor U20060 (N_20060,N_19878,N_19912);
nor U20061 (N_20061,N_19823,N_19772);
xor U20062 (N_20062,N_19967,N_19901);
or U20063 (N_20063,N_19932,N_19862);
xor U20064 (N_20064,N_19810,N_19757);
nor U20065 (N_20065,N_19946,N_19888);
xor U20066 (N_20066,N_19917,N_19815);
nand U20067 (N_20067,N_19993,N_19996);
or U20068 (N_20068,N_19988,N_19768);
or U20069 (N_20069,N_19849,N_19877);
nand U20070 (N_20070,N_19933,N_19755);
or U20071 (N_20071,N_19944,N_19854);
nand U20072 (N_20072,N_19879,N_19822);
or U20073 (N_20073,N_19857,N_19868);
nor U20074 (N_20074,N_19840,N_19975);
and U20075 (N_20075,N_19934,N_19853);
or U20076 (N_20076,N_19949,N_19830);
and U20077 (N_20077,N_19832,N_19941);
and U20078 (N_20078,N_19972,N_19829);
nand U20079 (N_20079,N_19915,N_19864);
xor U20080 (N_20080,N_19963,N_19751);
xnor U20081 (N_20081,N_19992,N_19756);
xnor U20082 (N_20082,N_19813,N_19788);
xor U20083 (N_20083,N_19887,N_19752);
and U20084 (N_20084,N_19817,N_19786);
nor U20085 (N_20085,N_19925,N_19767);
xor U20086 (N_20086,N_19808,N_19875);
or U20087 (N_20087,N_19906,N_19826);
xnor U20088 (N_20088,N_19828,N_19812);
nor U20089 (N_20089,N_19764,N_19831);
and U20090 (N_20090,N_19769,N_19798);
nor U20091 (N_20091,N_19979,N_19867);
or U20092 (N_20092,N_19804,N_19937);
and U20093 (N_20093,N_19794,N_19881);
and U20094 (N_20094,N_19803,N_19903);
and U20095 (N_20095,N_19897,N_19964);
or U20096 (N_20096,N_19939,N_19781);
nand U20097 (N_20097,N_19970,N_19872);
and U20098 (N_20098,N_19945,N_19865);
and U20099 (N_20099,N_19980,N_19763);
and U20100 (N_20100,N_19960,N_19902);
or U20101 (N_20101,N_19895,N_19818);
or U20102 (N_20102,N_19896,N_19835);
xor U20103 (N_20103,N_19958,N_19921);
or U20104 (N_20104,N_19957,N_19836);
or U20105 (N_20105,N_19847,N_19984);
or U20106 (N_20106,N_19821,N_19951);
and U20107 (N_20107,N_19784,N_19942);
nor U20108 (N_20108,N_19841,N_19819);
nand U20109 (N_20109,N_19782,N_19807);
nor U20110 (N_20110,N_19973,N_19908);
nand U20111 (N_20111,N_19795,N_19971);
xor U20112 (N_20112,N_19913,N_19999);
or U20113 (N_20113,N_19760,N_19910);
and U20114 (N_20114,N_19780,N_19792);
nor U20115 (N_20115,N_19814,N_19998);
and U20116 (N_20116,N_19927,N_19838);
or U20117 (N_20117,N_19948,N_19929);
or U20118 (N_20118,N_19800,N_19994);
nor U20119 (N_20119,N_19762,N_19880);
nand U20120 (N_20120,N_19976,N_19952);
nor U20121 (N_20121,N_19778,N_19968);
or U20122 (N_20122,N_19789,N_19858);
nand U20123 (N_20123,N_19876,N_19977);
nor U20124 (N_20124,N_19918,N_19909);
xnor U20125 (N_20125,N_19940,N_19861);
or U20126 (N_20126,N_19759,N_19773);
nor U20127 (N_20127,N_19977,N_19983);
and U20128 (N_20128,N_19785,N_19790);
or U20129 (N_20129,N_19912,N_19837);
or U20130 (N_20130,N_19858,N_19758);
nor U20131 (N_20131,N_19902,N_19892);
nand U20132 (N_20132,N_19928,N_19894);
nand U20133 (N_20133,N_19896,N_19894);
nor U20134 (N_20134,N_19966,N_19897);
nand U20135 (N_20135,N_19776,N_19949);
nand U20136 (N_20136,N_19960,N_19986);
nor U20137 (N_20137,N_19846,N_19995);
nor U20138 (N_20138,N_19957,N_19785);
nor U20139 (N_20139,N_19851,N_19825);
xnor U20140 (N_20140,N_19995,N_19890);
nor U20141 (N_20141,N_19753,N_19770);
xor U20142 (N_20142,N_19992,N_19782);
or U20143 (N_20143,N_19966,N_19765);
xor U20144 (N_20144,N_19785,N_19951);
and U20145 (N_20145,N_19915,N_19876);
nor U20146 (N_20146,N_19885,N_19910);
nand U20147 (N_20147,N_19756,N_19836);
nor U20148 (N_20148,N_19974,N_19961);
and U20149 (N_20149,N_19852,N_19980);
and U20150 (N_20150,N_19883,N_19868);
or U20151 (N_20151,N_19839,N_19844);
xnor U20152 (N_20152,N_19775,N_19902);
xor U20153 (N_20153,N_19922,N_19910);
xnor U20154 (N_20154,N_19875,N_19861);
nand U20155 (N_20155,N_19816,N_19771);
and U20156 (N_20156,N_19979,N_19998);
and U20157 (N_20157,N_19945,N_19922);
and U20158 (N_20158,N_19816,N_19909);
xnor U20159 (N_20159,N_19823,N_19963);
nor U20160 (N_20160,N_19753,N_19799);
nand U20161 (N_20161,N_19941,N_19820);
and U20162 (N_20162,N_19928,N_19839);
and U20163 (N_20163,N_19887,N_19906);
and U20164 (N_20164,N_19821,N_19874);
and U20165 (N_20165,N_19783,N_19836);
nor U20166 (N_20166,N_19911,N_19822);
nand U20167 (N_20167,N_19835,N_19942);
nor U20168 (N_20168,N_19829,N_19848);
nor U20169 (N_20169,N_19852,N_19979);
or U20170 (N_20170,N_19994,N_19848);
nand U20171 (N_20171,N_19946,N_19758);
xor U20172 (N_20172,N_19794,N_19852);
and U20173 (N_20173,N_19805,N_19835);
and U20174 (N_20174,N_19790,N_19853);
and U20175 (N_20175,N_19791,N_19750);
or U20176 (N_20176,N_19895,N_19957);
xor U20177 (N_20177,N_19969,N_19860);
xor U20178 (N_20178,N_19759,N_19819);
and U20179 (N_20179,N_19778,N_19922);
nor U20180 (N_20180,N_19839,N_19869);
nand U20181 (N_20181,N_19930,N_19954);
nor U20182 (N_20182,N_19808,N_19777);
xor U20183 (N_20183,N_19979,N_19847);
nor U20184 (N_20184,N_19817,N_19909);
or U20185 (N_20185,N_19964,N_19925);
nor U20186 (N_20186,N_19828,N_19894);
and U20187 (N_20187,N_19942,N_19787);
nand U20188 (N_20188,N_19765,N_19796);
nor U20189 (N_20189,N_19843,N_19814);
nor U20190 (N_20190,N_19935,N_19790);
nor U20191 (N_20191,N_19811,N_19790);
and U20192 (N_20192,N_19875,N_19786);
xor U20193 (N_20193,N_19783,N_19951);
nor U20194 (N_20194,N_19824,N_19755);
or U20195 (N_20195,N_19896,N_19759);
nor U20196 (N_20196,N_19877,N_19969);
nor U20197 (N_20197,N_19992,N_19996);
nor U20198 (N_20198,N_19770,N_19908);
nand U20199 (N_20199,N_19920,N_19859);
xor U20200 (N_20200,N_19968,N_19823);
nand U20201 (N_20201,N_19844,N_19830);
nand U20202 (N_20202,N_19797,N_19922);
xor U20203 (N_20203,N_19847,N_19907);
and U20204 (N_20204,N_19968,N_19806);
or U20205 (N_20205,N_19838,N_19947);
xnor U20206 (N_20206,N_19993,N_19972);
and U20207 (N_20207,N_19831,N_19880);
xnor U20208 (N_20208,N_19806,N_19833);
nor U20209 (N_20209,N_19981,N_19836);
nor U20210 (N_20210,N_19796,N_19873);
or U20211 (N_20211,N_19989,N_19807);
xor U20212 (N_20212,N_19968,N_19936);
or U20213 (N_20213,N_19808,N_19800);
xnor U20214 (N_20214,N_19781,N_19989);
nor U20215 (N_20215,N_19962,N_19754);
nand U20216 (N_20216,N_19817,N_19863);
nand U20217 (N_20217,N_19981,N_19937);
xnor U20218 (N_20218,N_19998,N_19809);
nand U20219 (N_20219,N_19876,N_19855);
nor U20220 (N_20220,N_19872,N_19918);
or U20221 (N_20221,N_19952,N_19953);
or U20222 (N_20222,N_19779,N_19946);
nand U20223 (N_20223,N_19921,N_19813);
nand U20224 (N_20224,N_19942,N_19884);
or U20225 (N_20225,N_19937,N_19987);
nand U20226 (N_20226,N_19804,N_19926);
and U20227 (N_20227,N_19925,N_19756);
nand U20228 (N_20228,N_19856,N_19932);
xnor U20229 (N_20229,N_19848,N_19995);
or U20230 (N_20230,N_19800,N_19998);
xnor U20231 (N_20231,N_19833,N_19795);
xnor U20232 (N_20232,N_19951,N_19830);
and U20233 (N_20233,N_19958,N_19891);
or U20234 (N_20234,N_19821,N_19816);
and U20235 (N_20235,N_19845,N_19998);
xnor U20236 (N_20236,N_19787,N_19769);
nor U20237 (N_20237,N_19822,N_19903);
nand U20238 (N_20238,N_19958,N_19789);
nor U20239 (N_20239,N_19816,N_19765);
or U20240 (N_20240,N_19859,N_19793);
nand U20241 (N_20241,N_19976,N_19944);
nor U20242 (N_20242,N_19751,N_19960);
nand U20243 (N_20243,N_19845,N_19771);
or U20244 (N_20244,N_19926,N_19845);
xnor U20245 (N_20245,N_19969,N_19996);
nand U20246 (N_20246,N_19880,N_19997);
nor U20247 (N_20247,N_19874,N_19927);
or U20248 (N_20248,N_19759,N_19944);
nor U20249 (N_20249,N_19765,N_19775);
xor U20250 (N_20250,N_20194,N_20076);
and U20251 (N_20251,N_20001,N_20026);
or U20252 (N_20252,N_20225,N_20229);
nand U20253 (N_20253,N_20034,N_20049);
nor U20254 (N_20254,N_20226,N_20006);
xnor U20255 (N_20255,N_20198,N_20205);
nand U20256 (N_20256,N_20074,N_20000);
nand U20257 (N_20257,N_20172,N_20022);
nand U20258 (N_20258,N_20035,N_20090);
nor U20259 (N_20259,N_20152,N_20030);
and U20260 (N_20260,N_20106,N_20143);
nor U20261 (N_20261,N_20244,N_20188);
nand U20262 (N_20262,N_20222,N_20095);
and U20263 (N_20263,N_20096,N_20159);
and U20264 (N_20264,N_20230,N_20206);
nand U20265 (N_20265,N_20080,N_20204);
and U20266 (N_20266,N_20011,N_20081);
nor U20267 (N_20267,N_20154,N_20068);
nand U20268 (N_20268,N_20043,N_20217);
nor U20269 (N_20269,N_20157,N_20147);
nand U20270 (N_20270,N_20187,N_20200);
nor U20271 (N_20271,N_20211,N_20097);
and U20272 (N_20272,N_20041,N_20228);
xor U20273 (N_20273,N_20137,N_20042);
or U20274 (N_20274,N_20027,N_20105);
and U20275 (N_20275,N_20162,N_20248);
nor U20276 (N_20276,N_20117,N_20184);
nand U20277 (N_20277,N_20048,N_20242);
xor U20278 (N_20278,N_20039,N_20218);
and U20279 (N_20279,N_20123,N_20046);
xnor U20280 (N_20280,N_20122,N_20167);
xnor U20281 (N_20281,N_20209,N_20085);
and U20282 (N_20282,N_20234,N_20063);
xnor U20283 (N_20283,N_20249,N_20127);
nand U20284 (N_20284,N_20082,N_20164);
and U20285 (N_20285,N_20240,N_20091);
and U20286 (N_20286,N_20212,N_20107);
nor U20287 (N_20287,N_20037,N_20195);
and U20288 (N_20288,N_20020,N_20138);
xnor U20289 (N_20289,N_20136,N_20017);
xnor U20290 (N_20290,N_20088,N_20216);
nand U20291 (N_20291,N_20060,N_20170);
nor U20292 (N_20292,N_20126,N_20062);
nor U20293 (N_20293,N_20141,N_20231);
or U20294 (N_20294,N_20031,N_20176);
and U20295 (N_20295,N_20189,N_20196);
nand U20296 (N_20296,N_20233,N_20246);
xnor U20297 (N_20297,N_20185,N_20044);
nand U20298 (N_20298,N_20086,N_20078);
and U20299 (N_20299,N_20066,N_20111);
and U20300 (N_20300,N_20092,N_20148);
or U20301 (N_20301,N_20207,N_20243);
and U20302 (N_20302,N_20210,N_20003);
or U20303 (N_20303,N_20239,N_20101);
nand U20304 (N_20304,N_20221,N_20102);
nand U20305 (N_20305,N_20114,N_20150);
nand U20306 (N_20306,N_20015,N_20193);
nor U20307 (N_20307,N_20131,N_20174);
nand U20308 (N_20308,N_20168,N_20202);
nand U20309 (N_20309,N_20009,N_20007);
xnor U20310 (N_20310,N_20171,N_20112);
nand U20311 (N_20311,N_20104,N_20247);
and U20312 (N_20312,N_20100,N_20077);
and U20313 (N_20313,N_20245,N_20156);
nor U20314 (N_20314,N_20047,N_20093);
or U20315 (N_20315,N_20010,N_20014);
nand U20316 (N_20316,N_20002,N_20232);
and U20317 (N_20317,N_20110,N_20181);
or U20318 (N_20318,N_20197,N_20169);
or U20319 (N_20319,N_20103,N_20113);
nor U20320 (N_20320,N_20235,N_20199);
nor U20321 (N_20321,N_20072,N_20178);
and U20322 (N_20322,N_20055,N_20144);
and U20323 (N_20323,N_20213,N_20099);
or U20324 (N_20324,N_20050,N_20087);
xnor U20325 (N_20325,N_20177,N_20132);
and U20326 (N_20326,N_20089,N_20019);
nand U20327 (N_20327,N_20203,N_20237);
nand U20328 (N_20328,N_20033,N_20018);
and U20329 (N_20329,N_20115,N_20130);
or U20330 (N_20330,N_20149,N_20139);
nand U20331 (N_20331,N_20182,N_20094);
nand U20332 (N_20332,N_20160,N_20153);
xnor U20333 (N_20333,N_20201,N_20215);
and U20334 (N_20334,N_20016,N_20128);
or U20335 (N_20335,N_20029,N_20125);
xor U20336 (N_20336,N_20109,N_20052);
nand U20337 (N_20337,N_20163,N_20053);
xor U20338 (N_20338,N_20040,N_20175);
or U20339 (N_20339,N_20173,N_20038);
and U20340 (N_20340,N_20238,N_20056);
nand U20341 (N_20341,N_20071,N_20057);
or U20342 (N_20342,N_20223,N_20116);
xnor U20343 (N_20343,N_20023,N_20183);
nor U20344 (N_20344,N_20108,N_20191);
xor U20345 (N_20345,N_20224,N_20166);
or U20346 (N_20346,N_20145,N_20059);
and U20347 (N_20347,N_20075,N_20151);
and U20348 (N_20348,N_20008,N_20058);
and U20349 (N_20349,N_20241,N_20012);
and U20350 (N_20350,N_20236,N_20051);
or U20351 (N_20351,N_20054,N_20155);
and U20352 (N_20352,N_20120,N_20079);
and U20353 (N_20353,N_20158,N_20045);
xnor U20354 (N_20354,N_20124,N_20161);
nor U20355 (N_20355,N_20013,N_20118);
and U20356 (N_20356,N_20121,N_20024);
xor U20357 (N_20357,N_20069,N_20192);
or U20358 (N_20358,N_20180,N_20219);
nand U20359 (N_20359,N_20140,N_20186);
nor U20360 (N_20360,N_20165,N_20032);
or U20361 (N_20361,N_20064,N_20208);
or U20362 (N_20362,N_20025,N_20227);
nor U20363 (N_20363,N_20146,N_20004);
nand U20364 (N_20364,N_20119,N_20005);
xnor U20365 (N_20365,N_20028,N_20129);
xor U20366 (N_20366,N_20021,N_20083);
nand U20367 (N_20367,N_20036,N_20179);
xnor U20368 (N_20368,N_20084,N_20134);
xor U20369 (N_20369,N_20061,N_20220);
or U20370 (N_20370,N_20133,N_20067);
xor U20371 (N_20371,N_20065,N_20214);
and U20372 (N_20372,N_20070,N_20098);
or U20373 (N_20373,N_20073,N_20142);
xnor U20374 (N_20374,N_20135,N_20190);
and U20375 (N_20375,N_20011,N_20223);
xnor U20376 (N_20376,N_20161,N_20148);
or U20377 (N_20377,N_20196,N_20234);
or U20378 (N_20378,N_20233,N_20146);
or U20379 (N_20379,N_20190,N_20009);
nor U20380 (N_20380,N_20116,N_20213);
nand U20381 (N_20381,N_20182,N_20018);
nor U20382 (N_20382,N_20215,N_20004);
nand U20383 (N_20383,N_20183,N_20207);
or U20384 (N_20384,N_20091,N_20157);
nand U20385 (N_20385,N_20187,N_20060);
or U20386 (N_20386,N_20220,N_20094);
nor U20387 (N_20387,N_20135,N_20164);
and U20388 (N_20388,N_20197,N_20074);
and U20389 (N_20389,N_20021,N_20056);
nor U20390 (N_20390,N_20072,N_20198);
and U20391 (N_20391,N_20209,N_20100);
and U20392 (N_20392,N_20136,N_20219);
and U20393 (N_20393,N_20244,N_20182);
nor U20394 (N_20394,N_20121,N_20031);
and U20395 (N_20395,N_20152,N_20011);
or U20396 (N_20396,N_20213,N_20093);
or U20397 (N_20397,N_20041,N_20118);
and U20398 (N_20398,N_20145,N_20199);
and U20399 (N_20399,N_20197,N_20045);
xnor U20400 (N_20400,N_20161,N_20232);
nor U20401 (N_20401,N_20105,N_20018);
nand U20402 (N_20402,N_20135,N_20170);
nand U20403 (N_20403,N_20166,N_20108);
xnor U20404 (N_20404,N_20090,N_20060);
nand U20405 (N_20405,N_20000,N_20024);
nand U20406 (N_20406,N_20105,N_20035);
nand U20407 (N_20407,N_20207,N_20091);
xnor U20408 (N_20408,N_20072,N_20107);
nor U20409 (N_20409,N_20006,N_20092);
and U20410 (N_20410,N_20095,N_20218);
and U20411 (N_20411,N_20153,N_20106);
and U20412 (N_20412,N_20211,N_20138);
nor U20413 (N_20413,N_20076,N_20117);
nand U20414 (N_20414,N_20236,N_20152);
nand U20415 (N_20415,N_20070,N_20242);
or U20416 (N_20416,N_20096,N_20111);
nand U20417 (N_20417,N_20237,N_20011);
or U20418 (N_20418,N_20102,N_20132);
nand U20419 (N_20419,N_20199,N_20116);
xnor U20420 (N_20420,N_20197,N_20065);
or U20421 (N_20421,N_20216,N_20137);
or U20422 (N_20422,N_20209,N_20169);
nor U20423 (N_20423,N_20090,N_20087);
nor U20424 (N_20424,N_20242,N_20116);
nor U20425 (N_20425,N_20034,N_20100);
nor U20426 (N_20426,N_20095,N_20076);
nor U20427 (N_20427,N_20244,N_20075);
xnor U20428 (N_20428,N_20157,N_20179);
xor U20429 (N_20429,N_20015,N_20187);
nor U20430 (N_20430,N_20077,N_20048);
xor U20431 (N_20431,N_20104,N_20082);
xnor U20432 (N_20432,N_20109,N_20054);
or U20433 (N_20433,N_20226,N_20183);
and U20434 (N_20434,N_20118,N_20024);
or U20435 (N_20435,N_20208,N_20222);
and U20436 (N_20436,N_20186,N_20183);
or U20437 (N_20437,N_20186,N_20181);
nand U20438 (N_20438,N_20099,N_20190);
nor U20439 (N_20439,N_20218,N_20172);
and U20440 (N_20440,N_20192,N_20207);
or U20441 (N_20441,N_20232,N_20206);
nand U20442 (N_20442,N_20146,N_20071);
nand U20443 (N_20443,N_20137,N_20228);
and U20444 (N_20444,N_20039,N_20227);
nand U20445 (N_20445,N_20070,N_20136);
nor U20446 (N_20446,N_20001,N_20139);
nor U20447 (N_20447,N_20172,N_20149);
and U20448 (N_20448,N_20136,N_20059);
and U20449 (N_20449,N_20214,N_20213);
nor U20450 (N_20450,N_20140,N_20238);
nor U20451 (N_20451,N_20195,N_20152);
or U20452 (N_20452,N_20093,N_20078);
and U20453 (N_20453,N_20186,N_20056);
nand U20454 (N_20454,N_20181,N_20108);
xnor U20455 (N_20455,N_20168,N_20142);
nand U20456 (N_20456,N_20149,N_20201);
nand U20457 (N_20457,N_20059,N_20206);
xnor U20458 (N_20458,N_20102,N_20133);
nand U20459 (N_20459,N_20217,N_20227);
nor U20460 (N_20460,N_20145,N_20082);
or U20461 (N_20461,N_20104,N_20088);
and U20462 (N_20462,N_20090,N_20174);
or U20463 (N_20463,N_20194,N_20175);
nor U20464 (N_20464,N_20243,N_20187);
and U20465 (N_20465,N_20007,N_20248);
and U20466 (N_20466,N_20176,N_20170);
nor U20467 (N_20467,N_20076,N_20201);
or U20468 (N_20468,N_20050,N_20043);
or U20469 (N_20469,N_20112,N_20188);
xor U20470 (N_20470,N_20008,N_20236);
xnor U20471 (N_20471,N_20014,N_20186);
xnor U20472 (N_20472,N_20245,N_20107);
or U20473 (N_20473,N_20126,N_20201);
or U20474 (N_20474,N_20014,N_20192);
or U20475 (N_20475,N_20151,N_20088);
or U20476 (N_20476,N_20102,N_20087);
nor U20477 (N_20477,N_20113,N_20166);
and U20478 (N_20478,N_20021,N_20038);
xor U20479 (N_20479,N_20015,N_20151);
nor U20480 (N_20480,N_20209,N_20113);
xor U20481 (N_20481,N_20240,N_20199);
nor U20482 (N_20482,N_20239,N_20169);
nand U20483 (N_20483,N_20164,N_20210);
xor U20484 (N_20484,N_20066,N_20070);
and U20485 (N_20485,N_20246,N_20097);
xor U20486 (N_20486,N_20134,N_20129);
and U20487 (N_20487,N_20007,N_20111);
nor U20488 (N_20488,N_20033,N_20102);
nor U20489 (N_20489,N_20175,N_20057);
nor U20490 (N_20490,N_20243,N_20181);
or U20491 (N_20491,N_20184,N_20205);
xor U20492 (N_20492,N_20129,N_20191);
nand U20493 (N_20493,N_20062,N_20166);
or U20494 (N_20494,N_20148,N_20001);
nand U20495 (N_20495,N_20045,N_20021);
and U20496 (N_20496,N_20127,N_20074);
xor U20497 (N_20497,N_20230,N_20123);
nand U20498 (N_20498,N_20097,N_20126);
nor U20499 (N_20499,N_20059,N_20119);
or U20500 (N_20500,N_20262,N_20358);
xor U20501 (N_20501,N_20296,N_20275);
xor U20502 (N_20502,N_20485,N_20497);
or U20503 (N_20503,N_20289,N_20364);
xnor U20504 (N_20504,N_20436,N_20339);
nor U20505 (N_20505,N_20373,N_20430);
nand U20506 (N_20506,N_20429,N_20444);
and U20507 (N_20507,N_20383,N_20439);
nand U20508 (N_20508,N_20405,N_20381);
nor U20509 (N_20509,N_20366,N_20449);
nor U20510 (N_20510,N_20377,N_20338);
nor U20511 (N_20511,N_20269,N_20354);
nand U20512 (N_20512,N_20412,N_20406);
and U20513 (N_20513,N_20433,N_20431);
xnor U20514 (N_20514,N_20445,N_20257);
nand U20515 (N_20515,N_20499,N_20476);
or U20516 (N_20516,N_20276,N_20318);
nand U20517 (N_20517,N_20477,N_20341);
or U20518 (N_20518,N_20435,N_20492);
xor U20519 (N_20519,N_20349,N_20409);
xor U20520 (N_20520,N_20376,N_20374);
or U20521 (N_20521,N_20407,N_20311);
and U20522 (N_20522,N_20400,N_20454);
nand U20523 (N_20523,N_20333,N_20369);
xnor U20524 (N_20524,N_20288,N_20388);
nor U20525 (N_20525,N_20284,N_20325);
nand U20526 (N_20526,N_20292,N_20302);
or U20527 (N_20527,N_20352,N_20357);
nand U20528 (N_20528,N_20294,N_20490);
and U20529 (N_20529,N_20448,N_20372);
xnor U20530 (N_20530,N_20415,N_20368);
xnor U20531 (N_20531,N_20460,N_20346);
nand U20532 (N_20532,N_20273,N_20469);
or U20533 (N_20533,N_20321,N_20272);
nor U20534 (N_20534,N_20422,N_20270);
xnor U20535 (N_20535,N_20336,N_20319);
and U20536 (N_20536,N_20278,N_20393);
or U20537 (N_20537,N_20252,N_20471);
nor U20538 (N_20538,N_20256,N_20451);
or U20539 (N_20539,N_20378,N_20255);
and U20540 (N_20540,N_20335,N_20259);
nand U20541 (N_20541,N_20323,N_20283);
or U20542 (N_20542,N_20466,N_20457);
or U20543 (N_20543,N_20455,N_20394);
xnor U20544 (N_20544,N_20390,N_20313);
xor U20545 (N_20545,N_20450,N_20332);
and U20546 (N_20546,N_20356,N_20309);
or U20547 (N_20547,N_20481,N_20307);
xnor U20548 (N_20548,N_20297,N_20316);
nor U20549 (N_20549,N_20367,N_20385);
or U20550 (N_20550,N_20462,N_20387);
and U20551 (N_20551,N_20280,N_20446);
nor U20552 (N_20552,N_20310,N_20464);
nor U20553 (N_20553,N_20375,N_20285);
or U20554 (N_20554,N_20482,N_20343);
and U20555 (N_20555,N_20402,N_20328);
nand U20556 (N_20556,N_20331,N_20326);
or U20557 (N_20557,N_20324,N_20350);
nor U20558 (N_20558,N_20303,N_20437);
or U20559 (N_20559,N_20342,N_20487);
nand U20560 (N_20560,N_20353,N_20362);
or U20561 (N_20561,N_20291,N_20371);
or U20562 (N_20562,N_20399,N_20317);
or U20563 (N_20563,N_20484,N_20271);
nand U20564 (N_20564,N_20461,N_20473);
nor U20565 (N_20565,N_20401,N_20327);
and U20566 (N_20566,N_20410,N_20403);
or U20567 (N_20567,N_20480,N_20470);
and U20568 (N_20568,N_20467,N_20298);
or U20569 (N_20569,N_20475,N_20465);
nor U20570 (N_20570,N_20413,N_20299);
nand U20571 (N_20571,N_20428,N_20261);
and U20572 (N_20572,N_20293,N_20258);
nor U20573 (N_20573,N_20396,N_20404);
nand U20574 (N_20574,N_20295,N_20389);
nand U20575 (N_20575,N_20495,N_20419);
xnor U20576 (N_20576,N_20264,N_20488);
nor U20577 (N_20577,N_20370,N_20434);
nor U20578 (N_20578,N_20282,N_20498);
xor U20579 (N_20579,N_20260,N_20384);
xor U20580 (N_20580,N_20496,N_20427);
xnor U20581 (N_20581,N_20398,N_20305);
and U20582 (N_20582,N_20315,N_20330);
nand U20583 (N_20583,N_20474,N_20363);
and U20584 (N_20584,N_20306,N_20438);
or U20585 (N_20585,N_20421,N_20416);
or U20586 (N_20586,N_20486,N_20453);
nor U20587 (N_20587,N_20301,N_20253);
or U20588 (N_20588,N_20365,N_20340);
or U20589 (N_20589,N_20494,N_20263);
or U20590 (N_20590,N_20268,N_20489);
nor U20591 (N_20591,N_20254,N_20382);
and U20592 (N_20592,N_20347,N_20432);
and U20593 (N_20593,N_20267,N_20287);
nor U20594 (N_20594,N_20392,N_20379);
or U20595 (N_20595,N_20265,N_20440);
xnor U20596 (N_20596,N_20290,N_20277);
and U20597 (N_20597,N_20337,N_20493);
and U20598 (N_20598,N_20459,N_20345);
and U20599 (N_20599,N_20463,N_20443);
or U20600 (N_20600,N_20414,N_20478);
or U20601 (N_20601,N_20314,N_20423);
or U20602 (N_20602,N_20420,N_20408);
and U20603 (N_20603,N_20411,N_20344);
nand U20604 (N_20604,N_20322,N_20397);
xnor U20605 (N_20605,N_20380,N_20458);
xnor U20606 (N_20606,N_20266,N_20251);
nor U20607 (N_20607,N_20351,N_20360);
and U20608 (N_20608,N_20424,N_20417);
nor U20609 (N_20609,N_20359,N_20447);
nand U20610 (N_20610,N_20418,N_20472);
nor U20611 (N_20611,N_20274,N_20361);
nor U20612 (N_20612,N_20468,N_20355);
or U20613 (N_20613,N_20483,N_20386);
and U20614 (N_20614,N_20391,N_20491);
nand U20615 (N_20615,N_20320,N_20286);
nor U20616 (N_20616,N_20304,N_20452);
nand U20617 (N_20617,N_20250,N_20300);
and U20618 (N_20618,N_20348,N_20456);
nand U20619 (N_20619,N_20308,N_20479);
xnor U20620 (N_20620,N_20329,N_20441);
and U20621 (N_20621,N_20425,N_20426);
and U20622 (N_20622,N_20312,N_20279);
and U20623 (N_20623,N_20395,N_20334);
nor U20624 (N_20624,N_20281,N_20442);
xnor U20625 (N_20625,N_20431,N_20392);
nor U20626 (N_20626,N_20448,N_20421);
xnor U20627 (N_20627,N_20311,N_20422);
nand U20628 (N_20628,N_20485,N_20259);
or U20629 (N_20629,N_20325,N_20254);
nand U20630 (N_20630,N_20389,N_20468);
or U20631 (N_20631,N_20358,N_20309);
or U20632 (N_20632,N_20335,N_20458);
or U20633 (N_20633,N_20336,N_20390);
nand U20634 (N_20634,N_20256,N_20336);
xor U20635 (N_20635,N_20470,N_20273);
or U20636 (N_20636,N_20436,N_20293);
xnor U20637 (N_20637,N_20253,N_20252);
nand U20638 (N_20638,N_20447,N_20298);
xor U20639 (N_20639,N_20288,N_20359);
nor U20640 (N_20640,N_20385,N_20404);
and U20641 (N_20641,N_20254,N_20465);
nor U20642 (N_20642,N_20406,N_20255);
xor U20643 (N_20643,N_20262,N_20494);
nor U20644 (N_20644,N_20345,N_20282);
nor U20645 (N_20645,N_20366,N_20487);
or U20646 (N_20646,N_20326,N_20265);
or U20647 (N_20647,N_20336,N_20466);
and U20648 (N_20648,N_20327,N_20307);
or U20649 (N_20649,N_20429,N_20451);
nand U20650 (N_20650,N_20400,N_20294);
or U20651 (N_20651,N_20486,N_20419);
and U20652 (N_20652,N_20458,N_20324);
or U20653 (N_20653,N_20386,N_20369);
or U20654 (N_20654,N_20363,N_20272);
nor U20655 (N_20655,N_20324,N_20255);
or U20656 (N_20656,N_20382,N_20371);
nand U20657 (N_20657,N_20446,N_20309);
xor U20658 (N_20658,N_20470,N_20406);
and U20659 (N_20659,N_20356,N_20437);
xor U20660 (N_20660,N_20294,N_20283);
or U20661 (N_20661,N_20359,N_20327);
nand U20662 (N_20662,N_20309,N_20496);
xor U20663 (N_20663,N_20410,N_20407);
and U20664 (N_20664,N_20415,N_20393);
xor U20665 (N_20665,N_20317,N_20287);
and U20666 (N_20666,N_20430,N_20441);
xnor U20667 (N_20667,N_20356,N_20381);
and U20668 (N_20668,N_20377,N_20494);
nor U20669 (N_20669,N_20286,N_20252);
xnor U20670 (N_20670,N_20348,N_20388);
nor U20671 (N_20671,N_20327,N_20347);
and U20672 (N_20672,N_20486,N_20476);
and U20673 (N_20673,N_20499,N_20406);
or U20674 (N_20674,N_20478,N_20371);
nor U20675 (N_20675,N_20400,N_20314);
xnor U20676 (N_20676,N_20443,N_20491);
nand U20677 (N_20677,N_20383,N_20479);
and U20678 (N_20678,N_20295,N_20481);
and U20679 (N_20679,N_20278,N_20299);
xnor U20680 (N_20680,N_20336,N_20352);
xnor U20681 (N_20681,N_20349,N_20406);
and U20682 (N_20682,N_20308,N_20397);
xnor U20683 (N_20683,N_20408,N_20320);
nand U20684 (N_20684,N_20371,N_20304);
nand U20685 (N_20685,N_20371,N_20457);
nand U20686 (N_20686,N_20405,N_20459);
xor U20687 (N_20687,N_20328,N_20280);
nor U20688 (N_20688,N_20432,N_20428);
nor U20689 (N_20689,N_20417,N_20415);
and U20690 (N_20690,N_20408,N_20288);
or U20691 (N_20691,N_20278,N_20345);
nand U20692 (N_20692,N_20466,N_20317);
and U20693 (N_20693,N_20373,N_20344);
or U20694 (N_20694,N_20355,N_20410);
nor U20695 (N_20695,N_20319,N_20346);
xnor U20696 (N_20696,N_20441,N_20270);
nor U20697 (N_20697,N_20467,N_20485);
and U20698 (N_20698,N_20485,N_20311);
nor U20699 (N_20699,N_20383,N_20258);
nand U20700 (N_20700,N_20376,N_20388);
or U20701 (N_20701,N_20326,N_20302);
and U20702 (N_20702,N_20331,N_20334);
xor U20703 (N_20703,N_20467,N_20330);
or U20704 (N_20704,N_20281,N_20318);
xnor U20705 (N_20705,N_20458,N_20486);
nand U20706 (N_20706,N_20425,N_20483);
or U20707 (N_20707,N_20416,N_20374);
nor U20708 (N_20708,N_20358,N_20491);
nand U20709 (N_20709,N_20392,N_20269);
and U20710 (N_20710,N_20298,N_20377);
or U20711 (N_20711,N_20435,N_20406);
nor U20712 (N_20712,N_20431,N_20263);
nor U20713 (N_20713,N_20453,N_20441);
and U20714 (N_20714,N_20395,N_20419);
xnor U20715 (N_20715,N_20319,N_20445);
nor U20716 (N_20716,N_20483,N_20448);
nor U20717 (N_20717,N_20490,N_20259);
and U20718 (N_20718,N_20253,N_20281);
or U20719 (N_20719,N_20364,N_20474);
nor U20720 (N_20720,N_20416,N_20267);
nand U20721 (N_20721,N_20381,N_20280);
nor U20722 (N_20722,N_20372,N_20304);
or U20723 (N_20723,N_20266,N_20331);
and U20724 (N_20724,N_20477,N_20332);
nand U20725 (N_20725,N_20312,N_20419);
nor U20726 (N_20726,N_20262,N_20317);
nor U20727 (N_20727,N_20256,N_20285);
nor U20728 (N_20728,N_20342,N_20453);
nor U20729 (N_20729,N_20487,N_20369);
nand U20730 (N_20730,N_20358,N_20316);
nor U20731 (N_20731,N_20401,N_20486);
and U20732 (N_20732,N_20269,N_20479);
xor U20733 (N_20733,N_20455,N_20341);
or U20734 (N_20734,N_20426,N_20454);
xor U20735 (N_20735,N_20406,N_20308);
nand U20736 (N_20736,N_20351,N_20405);
and U20737 (N_20737,N_20455,N_20471);
or U20738 (N_20738,N_20317,N_20438);
nand U20739 (N_20739,N_20402,N_20292);
or U20740 (N_20740,N_20288,N_20382);
and U20741 (N_20741,N_20265,N_20269);
or U20742 (N_20742,N_20405,N_20370);
xnor U20743 (N_20743,N_20321,N_20367);
or U20744 (N_20744,N_20315,N_20450);
nand U20745 (N_20745,N_20324,N_20455);
xnor U20746 (N_20746,N_20261,N_20454);
or U20747 (N_20747,N_20300,N_20356);
and U20748 (N_20748,N_20462,N_20469);
nand U20749 (N_20749,N_20497,N_20309);
nand U20750 (N_20750,N_20625,N_20651);
or U20751 (N_20751,N_20736,N_20618);
xnor U20752 (N_20752,N_20731,N_20504);
xnor U20753 (N_20753,N_20602,N_20746);
or U20754 (N_20754,N_20717,N_20701);
or U20755 (N_20755,N_20588,N_20559);
nor U20756 (N_20756,N_20562,N_20571);
or U20757 (N_20757,N_20688,N_20531);
and U20758 (N_20758,N_20724,N_20520);
or U20759 (N_20759,N_20560,N_20727);
or U20760 (N_20760,N_20681,N_20598);
nand U20761 (N_20761,N_20711,N_20595);
xnor U20762 (N_20762,N_20726,N_20600);
xnor U20763 (N_20763,N_20697,N_20555);
xor U20764 (N_20764,N_20526,N_20699);
xor U20765 (N_20765,N_20572,N_20645);
or U20766 (N_20766,N_20592,N_20657);
nor U20767 (N_20767,N_20505,N_20536);
nor U20768 (N_20768,N_20742,N_20668);
nand U20769 (N_20769,N_20741,N_20515);
nor U20770 (N_20770,N_20629,N_20690);
nand U20771 (N_20771,N_20709,N_20604);
or U20772 (N_20772,N_20579,N_20548);
or U20773 (N_20773,N_20619,N_20590);
xor U20774 (N_20774,N_20606,N_20691);
or U20775 (N_20775,N_20587,N_20671);
nor U20776 (N_20776,N_20540,N_20740);
and U20777 (N_20777,N_20612,N_20518);
xnor U20778 (N_20778,N_20738,N_20553);
nand U20779 (N_20779,N_20630,N_20650);
nor U20780 (N_20780,N_20733,N_20719);
nand U20781 (N_20781,N_20569,N_20644);
nor U20782 (N_20782,N_20667,N_20693);
or U20783 (N_20783,N_20643,N_20543);
nand U20784 (N_20784,N_20609,N_20591);
nor U20785 (N_20785,N_20581,N_20685);
nand U20786 (N_20786,N_20516,N_20537);
xor U20787 (N_20787,N_20639,N_20689);
xor U20788 (N_20788,N_20652,N_20649);
or U20789 (N_20789,N_20694,N_20509);
nor U20790 (N_20790,N_20605,N_20570);
or U20791 (N_20791,N_20554,N_20622);
nor U20792 (N_20792,N_20730,N_20669);
and U20793 (N_20793,N_20599,N_20656);
xor U20794 (N_20794,N_20675,N_20616);
nand U20795 (N_20795,N_20544,N_20692);
xor U20796 (N_20796,N_20682,N_20721);
and U20797 (N_20797,N_20603,N_20673);
nand U20798 (N_20798,N_20610,N_20703);
nor U20799 (N_20799,N_20678,N_20556);
nand U20800 (N_20800,N_20653,N_20666);
or U20801 (N_20801,N_20723,N_20614);
and U20802 (N_20802,N_20702,N_20617);
nor U20803 (N_20803,N_20745,N_20715);
nor U20804 (N_20804,N_20646,N_20734);
nand U20805 (N_20805,N_20743,N_20535);
nand U20806 (N_20806,N_20687,N_20718);
and U20807 (N_20807,N_20528,N_20534);
and U20808 (N_20808,N_20672,N_20561);
nor U20809 (N_20809,N_20541,N_20568);
nor U20810 (N_20810,N_20708,N_20503);
or U20811 (N_20811,N_20748,N_20589);
xor U20812 (N_20812,N_20552,N_20529);
or U20813 (N_20813,N_20729,N_20508);
xnor U20814 (N_20814,N_20707,N_20628);
nor U20815 (N_20815,N_20580,N_20514);
or U20816 (N_20816,N_20686,N_20547);
xnor U20817 (N_20817,N_20532,N_20513);
nor U20818 (N_20818,N_20608,N_20512);
nand U20819 (N_20819,N_20684,N_20549);
nand U20820 (N_20820,N_20594,N_20665);
or U20821 (N_20821,N_20533,N_20521);
and U20822 (N_20822,N_20631,N_20573);
or U20823 (N_20823,N_20615,N_20519);
nor U20824 (N_20824,N_20582,N_20525);
nand U20825 (N_20825,N_20524,N_20507);
nand U20826 (N_20826,N_20744,N_20621);
xor U20827 (N_20827,N_20725,N_20680);
nor U20828 (N_20828,N_20706,N_20500);
nor U20829 (N_20829,N_20597,N_20627);
nand U20830 (N_20830,N_20674,N_20527);
or U20831 (N_20831,N_20659,N_20633);
nand U20832 (N_20832,N_20623,N_20670);
and U20833 (N_20833,N_20558,N_20596);
and U20834 (N_20834,N_20655,N_20735);
nand U20835 (N_20835,N_20704,N_20698);
or U20836 (N_20836,N_20705,N_20530);
xor U20837 (N_20837,N_20576,N_20636);
and U20838 (N_20838,N_20574,N_20632);
nand U20839 (N_20839,N_20637,N_20586);
xnor U20840 (N_20840,N_20564,N_20722);
xnor U20841 (N_20841,N_20737,N_20695);
xor U20842 (N_20842,N_20663,N_20749);
and U20843 (N_20843,N_20660,N_20700);
xnor U20844 (N_20844,N_20662,N_20714);
and U20845 (N_20845,N_20506,N_20567);
nand U20846 (N_20846,N_20634,N_20739);
nor U20847 (N_20847,N_20575,N_20563);
nor U20848 (N_20848,N_20550,N_20511);
or U20849 (N_20849,N_20565,N_20523);
xnor U20850 (N_20850,N_20710,N_20578);
nand U20851 (N_20851,N_20638,N_20676);
or U20852 (N_20852,N_20557,N_20654);
nand U20853 (N_20853,N_20641,N_20640);
nand U20854 (N_20854,N_20611,N_20664);
or U20855 (N_20855,N_20585,N_20747);
xnor U20856 (N_20856,N_20517,N_20677);
xnor U20857 (N_20857,N_20607,N_20583);
and U20858 (N_20858,N_20716,N_20679);
nor U20859 (N_20859,N_20642,N_20593);
nor U20860 (N_20860,N_20683,N_20613);
nor U20861 (N_20861,N_20712,N_20728);
and U20862 (N_20862,N_20577,N_20648);
xor U20863 (N_20863,N_20696,N_20658);
nand U20864 (N_20864,N_20635,N_20601);
and U20865 (N_20865,N_20501,N_20732);
or U20866 (N_20866,N_20502,N_20626);
or U20867 (N_20867,N_20720,N_20624);
xor U20868 (N_20868,N_20647,N_20522);
xor U20869 (N_20869,N_20545,N_20510);
nor U20870 (N_20870,N_20620,N_20551);
and U20871 (N_20871,N_20584,N_20661);
nand U20872 (N_20872,N_20546,N_20713);
or U20873 (N_20873,N_20538,N_20539);
and U20874 (N_20874,N_20542,N_20566);
nor U20875 (N_20875,N_20614,N_20619);
or U20876 (N_20876,N_20549,N_20526);
xor U20877 (N_20877,N_20534,N_20637);
nand U20878 (N_20878,N_20585,N_20690);
nor U20879 (N_20879,N_20544,N_20615);
nand U20880 (N_20880,N_20558,N_20614);
or U20881 (N_20881,N_20595,N_20548);
xnor U20882 (N_20882,N_20552,N_20691);
nor U20883 (N_20883,N_20535,N_20733);
xnor U20884 (N_20884,N_20521,N_20543);
nand U20885 (N_20885,N_20741,N_20744);
nand U20886 (N_20886,N_20584,N_20540);
xor U20887 (N_20887,N_20589,N_20636);
nor U20888 (N_20888,N_20711,N_20693);
xnor U20889 (N_20889,N_20698,N_20563);
nor U20890 (N_20890,N_20566,N_20630);
nor U20891 (N_20891,N_20555,N_20554);
xor U20892 (N_20892,N_20567,N_20627);
or U20893 (N_20893,N_20746,N_20568);
nor U20894 (N_20894,N_20615,N_20709);
xnor U20895 (N_20895,N_20560,N_20631);
xnor U20896 (N_20896,N_20609,N_20541);
nor U20897 (N_20897,N_20672,N_20682);
and U20898 (N_20898,N_20592,N_20555);
and U20899 (N_20899,N_20631,N_20734);
nand U20900 (N_20900,N_20693,N_20707);
nor U20901 (N_20901,N_20663,N_20743);
nor U20902 (N_20902,N_20686,N_20587);
xor U20903 (N_20903,N_20630,N_20551);
nand U20904 (N_20904,N_20629,N_20528);
nand U20905 (N_20905,N_20547,N_20650);
nor U20906 (N_20906,N_20507,N_20702);
xnor U20907 (N_20907,N_20582,N_20528);
and U20908 (N_20908,N_20550,N_20687);
nor U20909 (N_20909,N_20528,N_20702);
nand U20910 (N_20910,N_20536,N_20538);
nor U20911 (N_20911,N_20709,N_20623);
nand U20912 (N_20912,N_20533,N_20586);
xor U20913 (N_20913,N_20533,N_20743);
nor U20914 (N_20914,N_20700,N_20637);
nor U20915 (N_20915,N_20507,N_20579);
xor U20916 (N_20916,N_20544,N_20583);
xor U20917 (N_20917,N_20613,N_20700);
nor U20918 (N_20918,N_20624,N_20600);
and U20919 (N_20919,N_20741,N_20684);
and U20920 (N_20920,N_20540,N_20524);
or U20921 (N_20921,N_20604,N_20692);
nand U20922 (N_20922,N_20659,N_20541);
or U20923 (N_20923,N_20527,N_20723);
nor U20924 (N_20924,N_20682,N_20674);
xor U20925 (N_20925,N_20603,N_20713);
nand U20926 (N_20926,N_20638,N_20669);
xnor U20927 (N_20927,N_20728,N_20599);
or U20928 (N_20928,N_20703,N_20587);
xor U20929 (N_20929,N_20609,N_20535);
nor U20930 (N_20930,N_20552,N_20515);
nand U20931 (N_20931,N_20679,N_20516);
xor U20932 (N_20932,N_20661,N_20729);
nor U20933 (N_20933,N_20700,N_20738);
xnor U20934 (N_20934,N_20595,N_20586);
xnor U20935 (N_20935,N_20509,N_20636);
nand U20936 (N_20936,N_20690,N_20616);
nand U20937 (N_20937,N_20735,N_20638);
nor U20938 (N_20938,N_20739,N_20645);
xnor U20939 (N_20939,N_20587,N_20540);
nor U20940 (N_20940,N_20568,N_20649);
and U20941 (N_20941,N_20701,N_20620);
xnor U20942 (N_20942,N_20530,N_20569);
and U20943 (N_20943,N_20657,N_20640);
nor U20944 (N_20944,N_20574,N_20702);
nand U20945 (N_20945,N_20539,N_20547);
or U20946 (N_20946,N_20657,N_20607);
nand U20947 (N_20947,N_20617,N_20682);
nor U20948 (N_20948,N_20604,N_20592);
nor U20949 (N_20949,N_20615,N_20677);
xnor U20950 (N_20950,N_20574,N_20718);
or U20951 (N_20951,N_20738,N_20617);
nor U20952 (N_20952,N_20715,N_20674);
and U20953 (N_20953,N_20506,N_20606);
nand U20954 (N_20954,N_20564,N_20538);
and U20955 (N_20955,N_20606,N_20717);
xnor U20956 (N_20956,N_20644,N_20694);
nand U20957 (N_20957,N_20654,N_20680);
nor U20958 (N_20958,N_20533,N_20558);
xor U20959 (N_20959,N_20544,N_20678);
nand U20960 (N_20960,N_20661,N_20510);
xor U20961 (N_20961,N_20627,N_20608);
xor U20962 (N_20962,N_20593,N_20726);
nor U20963 (N_20963,N_20741,N_20606);
or U20964 (N_20964,N_20653,N_20692);
or U20965 (N_20965,N_20651,N_20730);
nor U20966 (N_20966,N_20622,N_20638);
nor U20967 (N_20967,N_20672,N_20522);
xnor U20968 (N_20968,N_20542,N_20550);
nand U20969 (N_20969,N_20630,N_20660);
nor U20970 (N_20970,N_20737,N_20677);
nor U20971 (N_20971,N_20654,N_20590);
and U20972 (N_20972,N_20695,N_20688);
nor U20973 (N_20973,N_20596,N_20574);
nor U20974 (N_20974,N_20554,N_20634);
xnor U20975 (N_20975,N_20645,N_20578);
and U20976 (N_20976,N_20572,N_20541);
xnor U20977 (N_20977,N_20714,N_20520);
and U20978 (N_20978,N_20645,N_20664);
or U20979 (N_20979,N_20736,N_20665);
nor U20980 (N_20980,N_20682,N_20568);
nand U20981 (N_20981,N_20534,N_20567);
and U20982 (N_20982,N_20722,N_20738);
nor U20983 (N_20983,N_20618,N_20653);
xnor U20984 (N_20984,N_20723,N_20508);
or U20985 (N_20985,N_20567,N_20652);
xor U20986 (N_20986,N_20684,N_20552);
xnor U20987 (N_20987,N_20648,N_20646);
nor U20988 (N_20988,N_20646,N_20601);
xor U20989 (N_20989,N_20561,N_20620);
and U20990 (N_20990,N_20699,N_20585);
nor U20991 (N_20991,N_20519,N_20671);
xor U20992 (N_20992,N_20594,N_20510);
or U20993 (N_20993,N_20640,N_20701);
nand U20994 (N_20994,N_20695,N_20570);
xnor U20995 (N_20995,N_20554,N_20553);
nand U20996 (N_20996,N_20688,N_20537);
or U20997 (N_20997,N_20543,N_20696);
nor U20998 (N_20998,N_20737,N_20664);
or U20999 (N_20999,N_20549,N_20523);
xor U21000 (N_21000,N_20946,N_20994);
nand U21001 (N_21001,N_20862,N_20770);
xnor U21002 (N_21002,N_20964,N_20773);
or U21003 (N_21003,N_20819,N_20801);
and U21004 (N_21004,N_20932,N_20929);
xnor U21005 (N_21005,N_20910,N_20784);
nand U21006 (N_21006,N_20754,N_20891);
nand U21007 (N_21007,N_20860,N_20868);
xnor U21008 (N_21008,N_20813,N_20757);
or U21009 (N_21009,N_20959,N_20824);
and U21010 (N_21010,N_20919,N_20768);
and U21011 (N_21011,N_20978,N_20841);
and U21012 (N_21012,N_20962,N_20853);
or U21013 (N_21013,N_20986,N_20942);
xor U21014 (N_21014,N_20980,N_20923);
nor U21015 (N_21015,N_20976,N_20990);
nand U21016 (N_21016,N_20882,N_20949);
or U21017 (N_21017,N_20921,N_20933);
xnor U21018 (N_21018,N_20763,N_20952);
or U21019 (N_21019,N_20844,N_20792);
nor U21020 (N_21020,N_20890,N_20900);
or U21021 (N_21021,N_20960,N_20966);
and U21022 (N_21022,N_20835,N_20920);
nand U21023 (N_21023,N_20846,N_20941);
xor U21024 (N_21024,N_20951,N_20859);
and U21025 (N_21025,N_20796,N_20826);
xnor U21026 (N_21026,N_20797,N_20774);
and U21027 (N_21027,N_20988,N_20809);
xnor U21028 (N_21028,N_20857,N_20888);
nor U21029 (N_21029,N_20911,N_20790);
nor U21030 (N_21030,N_20788,N_20908);
nor U21031 (N_21031,N_20789,N_20756);
nor U21032 (N_21032,N_20970,N_20979);
xnor U21033 (N_21033,N_20850,N_20897);
xnor U21034 (N_21034,N_20800,N_20798);
nand U21035 (N_21035,N_20927,N_20963);
or U21036 (N_21036,N_20861,N_20836);
nor U21037 (N_21037,N_20937,N_20840);
xor U21038 (N_21038,N_20977,N_20777);
nor U21039 (N_21039,N_20917,N_20981);
and U21040 (N_21040,N_20764,N_20879);
nand U21041 (N_21041,N_20945,N_20944);
or U21042 (N_21042,N_20805,N_20761);
nand U21043 (N_21043,N_20810,N_20828);
and U21044 (N_21044,N_20998,N_20856);
xor U21045 (N_21045,N_20765,N_20975);
or U21046 (N_21046,N_20995,N_20875);
or U21047 (N_21047,N_20876,N_20881);
nor U21048 (N_21048,N_20851,N_20845);
nand U21049 (N_21049,N_20827,N_20779);
xnor U21050 (N_21050,N_20926,N_20829);
nand U21051 (N_21051,N_20934,N_20930);
nor U21052 (N_21052,N_20795,N_20902);
or U21053 (N_21053,N_20913,N_20928);
xor U21054 (N_21054,N_20794,N_20968);
nor U21055 (N_21055,N_20948,N_20993);
nor U21056 (N_21056,N_20954,N_20907);
nor U21057 (N_21057,N_20989,N_20936);
nor U21058 (N_21058,N_20894,N_20984);
and U21059 (N_21059,N_20940,N_20867);
xor U21060 (N_21060,N_20807,N_20895);
or U21061 (N_21061,N_20755,N_20969);
or U21062 (N_21062,N_20950,N_20778);
xor U21063 (N_21063,N_20837,N_20781);
nand U21064 (N_21064,N_20814,N_20839);
nand U21065 (N_21065,N_20838,N_20922);
nor U21066 (N_21066,N_20785,N_20865);
nand U21067 (N_21067,N_20766,N_20991);
xor U21068 (N_21068,N_20831,N_20904);
nand U21069 (N_21069,N_20909,N_20752);
nand U21070 (N_21070,N_20855,N_20912);
nand U21071 (N_21071,N_20870,N_20915);
xor U21072 (N_21072,N_20762,N_20997);
and U21073 (N_21073,N_20808,N_20822);
and U21074 (N_21074,N_20769,N_20958);
or U21075 (N_21075,N_20873,N_20974);
nand U21076 (N_21076,N_20914,N_20820);
xor U21077 (N_21077,N_20804,N_20871);
nand U21078 (N_21078,N_20925,N_20877);
xnor U21079 (N_21079,N_20869,N_20996);
and U21080 (N_21080,N_20815,N_20898);
xor U21081 (N_21081,N_20823,N_20965);
nor U21082 (N_21082,N_20818,N_20812);
nand U21083 (N_21083,N_20906,N_20834);
or U21084 (N_21084,N_20772,N_20816);
or U21085 (N_21085,N_20759,N_20866);
and U21086 (N_21086,N_20874,N_20767);
or U21087 (N_21087,N_20848,N_20987);
nor U21088 (N_21088,N_20905,N_20939);
nor U21089 (N_21089,N_20901,N_20825);
or U21090 (N_21090,N_20854,N_20982);
nand U21091 (N_21091,N_20776,N_20889);
nand U21092 (N_21092,N_20892,N_20842);
nand U21093 (N_21093,N_20878,N_20863);
xor U21094 (N_21094,N_20791,N_20751);
nand U21095 (N_21095,N_20953,N_20832);
or U21096 (N_21096,N_20771,N_20864);
and U21097 (N_21097,N_20880,N_20985);
or U21098 (N_21098,N_20817,N_20786);
xnor U21099 (N_21099,N_20799,N_20811);
nand U21100 (N_21100,N_20775,N_20852);
xor U21101 (N_21101,N_20955,N_20780);
xor U21102 (N_21102,N_20787,N_20957);
and U21103 (N_21103,N_20821,N_20803);
and U21104 (N_21104,N_20903,N_20849);
and U21105 (N_21105,N_20971,N_20961);
and U21106 (N_21106,N_20899,N_20847);
or U21107 (N_21107,N_20806,N_20843);
or U21108 (N_21108,N_20887,N_20872);
or U21109 (N_21109,N_20830,N_20802);
nand U21110 (N_21110,N_20967,N_20924);
nor U21111 (N_21111,N_20999,N_20883);
nor U21112 (N_21112,N_20938,N_20858);
nor U21113 (N_21113,N_20758,N_20893);
or U21114 (N_21114,N_20884,N_20833);
nand U21115 (N_21115,N_20886,N_20956);
xor U21116 (N_21116,N_20931,N_20782);
nor U21117 (N_21117,N_20916,N_20935);
and U21118 (N_21118,N_20943,N_20793);
nand U21119 (N_21119,N_20972,N_20973);
and U21120 (N_21120,N_20760,N_20750);
or U21121 (N_21121,N_20896,N_20753);
and U21122 (N_21122,N_20992,N_20783);
nor U21123 (N_21123,N_20918,N_20947);
and U21124 (N_21124,N_20885,N_20983);
or U21125 (N_21125,N_20766,N_20883);
or U21126 (N_21126,N_20786,N_20753);
and U21127 (N_21127,N_20795,N_20830);
or U21128 (N_21128,N_20891,N_20854);
nor U21129 (N_21129,N_20929,N_20759);
nor U21130 (N_21130,N_20960,N_20838);
nand U21131 (N_21131,N_20979,N_20807);
or U21132 (N_21132,N_20828,N_20758);
or U21133 (N_21133,N_20895,N_20767);
xnor U21134 (N_21134,N_20880,N_20909);
or U21135 (N_21135,N_20780,N_20864);
nor U21136 (N_21136,N_20921,N_20826);
xor U21137 (N_21137,N_20974,N_20827);
or U21138 (N_21138,N_20847,N_20944);
nand U21139 (N_21139,N_20949,N_20796);
nand U21140 (N_21140,N_20915,N_20882);
and U21141 (N_21141,N_20901,N_20992);
and U21142 (N_21142,N_20751,N_20854);
or U21143 (N_21143,N_20987,N_20909);
xor U21144 (N_21144,N_20764,N_20952);
nor U21145 (N_21145,N_20758,N_20876);
xnor U21146 (N_21146,N_20811,N_20786);
nor U21147 (N_21147,N_20931,N_20819);
nand U21148 (N_21148,N_20834,N_20795);
and U21149 (N_21149,N_20971,N_20893);
nor U21150 (N_21150,N_20883,N_20876);
nor U21151 (N_21151,N_20913,N_20934);
nand U21152 (N_21152,N_20928,N_20866);
xnor U21153 (N_21153,N_20844,N_20957);
or U21154 (N_21154,N_20879,N_20854);
and U21155 (N_21155,N_20881,N_20781);
nand U21156 (N_21156,N_20921,N_20889);
nand U21157 (N_21157,N_20844,N_20959);
nor U21158 (N_21158,N_20943,N_20921);
xor U21159 (N_21159,N_20907,N_20919);
and U21160 (N_21160,N_20864,N_20797);
or U21161 (N_21161,N_20922,N_20823);
and U21162 (N_21162,N_20845,N_20966);
nand U21163 (N_21163,N_20779,N_20757);
nand U21164 (N_21164,N_20756,N_20942);
xnor U21165 (N_21165,N_20860,N_20854);
or U21166 (N_21166,N_20934,N_20905);
xnor U21167 (N_21167,N_20976,N_20776);
nand U21168 (N_21168,N_20996,N_20978);
or U21169 (N_21169,N_20832,N_20808);
xnor U21170 (N_21170,N_20945,N_20992);
or U21171 (N_21171,N_20775,N_20862);
and U21172 (N_21172,N_20854,N_20881);
xnor U21173 (N_21173,N_20829,N_20850);
nor U21174 (N_21174,N_20945,N_20972);
xor U21175 (N_21175,N_20997,N_20892);
xnor U21176 (N_21176,N_20890,N_20764);
or U21177 (N_21177,N_20767,N_20890);
xor U21178 (N_21178,N_20927,N_20851);
and U21179 (N_21179,N_20778,N_20881);
nor U21180 (N_21180,N_20859,N_20920);
nor U21181 (N_21181,N_20834,N_20769);
xor U21182 (N_21182,N_20877,N_20779);
xor U21183 (N_21183,N_20765,N_20894);
xor U21184 (N_21184,N_20992,N_20761);
or U21185 (N_21185,N_20824,N_20773);
xnor U21186 (N_21186,N_20922,N_20869);
or U21187 (N_21187,N_20821,N_20779);
and U21188 (N_21188,N_20880,N_20791);
xnor U21189 (N_21189,N_20965,N_20855);
and U21190 (N_21190,N_20799,N_20915);
and U21191 (N_21191,N_20909,N_20805);
nand U21192 (N_21192,N_20757,N_20973);
nand U21193 (N_21193,N_20781,N_20767);
or U21194 (N_21194,N_20766,N_20947);
xnor U21195 (N_21195,N_20997,N_20901);
nor U21196 (N_21196,N_20795,N_20858);
and U21197 (N_21197,N_20786,N_20777);
or U21198 (N_21198,N_20833,N_20913);
xnor U21199 (N_21199,N_20971,N_20954);
xnor U21200 (N_21200,N_20803,N_20770);
nor U21201 (N_21201,N_20972,N_20904);
nor U21202 (N_21202,N_20982,N_20768);
or U21203 (N_21203,N_20943,N_20930);
nand U21204 (N_21204,N_20859,N_20901);
or U21205 (N_21205,N_20870,N_20818);
nor U21206 (N_21206,N_20906,N_20774);
xnor U21207 (N_21207,N_20895,N_20814);
nor U21208 (N_21208,N_20877,N_20798);
nand U21209 (N_21209,N_20915,N_20969);
xor U21210 (N_21210,N_20852,N_20964);
nor U21211 (N_21211,N_20795,N_20891);
nor U21212 (N_21212,N_20928,N_20750);
or U21213 (N_21213,N_20891,N_20889);
or U21214 (N_21214,N_20763,N_20991);
and U21215 (N_21215,N_20963,N_20972);
xnor U21216 (N_21216,N_20945,N_20816);
nor U21217 (N_21217,N_20961,N_20778);
and U21218 (N_21218,N_20820,N_20992);
and U21219 (N_21219,N_20919,N_20826);
xnor U21220 (N_21220,N_20816,N_20979);
or U21221 (N_21221,N_20876,N_20906);
and U21222 (N_21222,N_20849,N_20914);
and U21223 (N_21223,N_20818,N_20825);
nor U21224 (N_21224,N_20857,N_20991);
and U21225 (N_21225,N_20773,N_20779);
or U21226 (N_21226,N_20911,N_20908);
nor U21227 (N_21227,N_20763,N_20822);
or U21228 (N_21228,N_20952,N_20932);
or U21229 (N_21229,N_20832,N_20964);
or U21230 (N_21230,N_20777,N_20825);
and U21231 (N_21231,N_20781,N_20834);
nand U21232 (N_21232,N_20949,N_20759);
xor U21233 (N_21233,N_20794,N_20857);
nor U21234 (N_21234,N_20921,N_20759);
or U21235 (N_21235,N_20809,N_20973);
nand U21236 (N_21236,N_20919,N_20873);
or U21237 (N_21237,N_20750,N_20888);
or U21238 (N_21238,N_20769,N_20818);
and U21239 (N_21239,N_20816,N_20821);
and U21240 (N_21240,N_20921,N_20872);
xor U21241 (N_21241,N_20809,N_20822);
nand U21242 (N_21242,N_20806,N_20781);
nand U21243 (N_21243,N_20945,N_20890);
or U21244 (N_21244,N_20850,N_20903);
or U21245 (N_21245,N_20953,N_20987);
xnor U21246 (N_21246,N_20781,N_20754);
nor U21247 (N_21247,N_20945,N_20796);
and U21248 (N_21248,N_20979,N_20856);
xnor U21249 (N_21249,N_20902,N_20951);
and U21250 (N_21250,N_21087,N_21112);
and U21251 (N_21251,N_21211,N_21127);
and U21252 (N_21252,N_21222,N_21081);
nor U21253 (N_21253,N_21073,N_21241);
or U21254 (N_21254,N_21044,N_21062);
xor U21255 (N_21255,N_21102,N_21111);
xor U21256 (N_21256,N_21025,N_21061);
xnor U21257 (N_21257,N_21089,N_21224);
and U21258 (N_21258,N_21085,N_21210);
or U21259 (N_21259,N_21139,N_21043);
nor U21260 (N_21260,N_21167,N_21131);
or U21261 (N_21261,N_21200,N_21124);
nand U21262 (N_21262,N_21153,N_21152);
xnor U21263 (N_21263,N_21171,N_21020);
nor U21264 (N_21264,N_21180,N_21094);
nor U21265 (N_21265,N_21203,N_21132);
xor U21266 (N_21266,N_21235,N_21060);
and U21267 (N_21267,N_21077,N_21202);
xnor U21268 (N_21268,N_21105,N_21100);
xnor U21269 (N_21269,N_21023,N_21158);
or U21270 (N_21270,N_21176,N_21246);
and U21271 (N_21271,N_21238,N_21206);
nand U21272 (N_21272,N_21101,N_21187);
nand U21273 (N_21273,N_21198,N_21122);
and U21274 (N_21274,N_21134,N_21244);
or U21275 (N_21275,N_21226,N_21192);
nand U21276 (N_21276,N_21026,N_21018);
xnor U21277 (N_21277,N_21097,N_21181);
xor U21278 (N_21278,N_21215,N_21107);
nand U21279 (N_21279,N_21109,N_21248);
or U21280 (N_21280,N_21118,N_21195);
xnor U21281 (N_21281,N_21228,N_21136);
nand U21282 (N_21282,N_21027,N_21146);
xor U21283 (N_21283,N_21239,N_21116);
nor U21284 (N_21284,N_21040,N_21220);
xor U21285 (N_21285,N_21185,N_21186);
xnor U21286 (N_21286,N_21042,N_21227);
and U21287 (N_21287,N_21028,N_21247);
nor U21288 (N_21288,N_21141,N_21047);
and U21289 (N_21289,N_21166,N_21050);
nor U21290 (N_21290,N_21155,N_21205);
xor U21291 (N_21291,N_21173,N_21039);
and U21292 (N_21292,N_21191,N_21005);
nor U21293 (N_21293,N_21083,N_21189);
and U21294 (N_21294,N_21175,N_21138);
xnor U21295 (N_21295,N_21163,N_21148);
nor U21296 (N_21296,N_21168,N_21196);
or U21297 (N_21297,N_21236,N_21204);
or U21298 (N_21298,N_21119,N_21017);
nor U21299 (N_21299,N_21177,N_21135);
or U21300 (N_21300,N_21151,N_21022);
or U21301 (N_21301,N_21213,N_21065);
nor U21302 (N_21302,N_21103,N_21066);
nand U21303 (N_21303,N_21037,N_21174);
nand U21304 (N_21304,N_21019,N_21048);
or U21305 (N_21305,N_21142,N_21030);
and U21306 (N_21306,N_21096,N_21003);
nor U21307 (N_21307,N_21183,N_21034);
xor U21308 (N_21308,N_21046,N_21133);
and U21309 (N_21309,N_21216,N_21120);
or U21310 (N_21310,N_21117,N_21006);
nand U21311 (N_21311,N_21115,N_21075);
and U21312 (N_21312,N_21172,N_21218);
or U21313 (N_21313,N_21114,N_21147);
and U21314 (N_21314,N_21193,N_21179);
xor U21315 (N_21315,N_21063,N_21113);
and U21316 (N_21316,N_21240,N_21029);
and U21317 (N_21317,N_21064,N_21086);
and U21318 (N_21318,N_21217,N_21032);
nand U21319 (N_21319,N_21225,N_21232);
nand U21320 (N_21320,N_21011,N_21001);
xor U21321 (N_21321,N_21194,N_21130);
xnor U21322 (N_21322,N_21093,N_21229);
or U21323 (N_21323,N_21150,N_21201);
xnor U21324 (N_21324,N_21098,N_21121);
xnor U21325 (N_21325,N_21002,N_21071);
or U21326 (N_21326,N_21178,N_21092);
xnor U21327 (N_21327,N_21184,N_21234);
or U21328 (N_21328,N_21084,N_21008);
and U21329 (N_21329,N_21014,N_21049);
nor U21330 (N_21330,N_21095,N_21214);
nor U21331 (N_21331,N_21154,N_21208);
or U21332 (N_21332,N_21242,N_21016);
or U21333 (N_21333,N_21012,N_21143);
nor U21334 (N_21334,N_21038,N_21056);
and U21335 (N_21335,N_21041,N_21129);
nand U21336 (N_21336,N_21212,N_21207);
xor U21337 (N_21337,N_21233,N_21074);
xor U21338 (N_21338,N_21000,N_21007);
and U21339 (N_21339,N_21165,N_21024);
xnor U21340 (N_21340,N_21058,N_21080);
or U21341 (N_21341,N_21072,N_21188);
nor U21342 (N_21342,N_21209,N_21068);
nor U21343 (N_21343,N_21004,N_21013);
xor U21344 (N_21344,N_21045,N_21144);
nand U21345 (N_21345,N_21149,N_21125);
nand U21346 (N_21346,N_21159,N_21057);
nand U21347 (N_21347,N_21099,N_21082);
or U21348 (N_21348,N_21035,N_21108);
xor U21349 (N_21349,N_21182,N_21104);
xor U21350 (N_21350,N_21052,N_21164);
nor U21351 (N_21351,N_21090,N_21128);
or U21352 (N_21352,N_21157,N_21126);
nand U21353 (N_21353,N_21243,N_21033);
nor U21354 (N_21354,N_21055,N_21162);
xor U21355 (N_21355,N_21123,N_21145);
and U21356 (N_21356,N_21169,N_21223);
and U21357 (N_21357,N_21088,N_21076);
xor U21358 (N_21358,N_21110,N_21078);
xnor U21359 (N_21359,N_21010,N_21051);
xnor U21360 (N_21360,N_21031,N_21221);
and U21361 (N_21361,N_21036,N_21161);
or U21362 (N_21362,N_21160,N_21069);
nor U21363 (N_21363,N_21219,N_21079);
nand U21364 (N_21364,N_21059,N_21237);
or U21365 (N_21365,N_21156,N_21199);
nor U21366 (N_21366,N_21190,N_21231);
or U21367 (N_21367,N_21091,N_21106);
and U21368 (N_21368,N_21137,N_21009);
and U21369 (N_21369,N_21140,N_21054);
or U21370 (N_21370,N_21021,N_21053);
nand U21371 (N_21371,N_21230,N_21249);
and U21372 (N_21372,N_21245,N_21197);
xnor U21373 (N_21373,N_21067,N_21015);
nor U21374 (N_21374,N_21070,N_21170);
and U21375 (N_21375,N_21074,N_21208);
nor U21376 (N_21376,N_21000,N_21142);
and U21377 (N_21377,N_21176,N_21221);
or U21378 (N_21378,N_21143,N_21173);
and U21379 (N_21379,N_21243,N_21045);
nor U21380 (N_21380,N_21094,N_21159);
or U21381 (N_21381,N_21050,N_21078);
xnor U21382 (N_21382,N_21157,N_21034);
nand U21383 (N_21383,N_21202,N_21028);
nor U21384 (N_21384,N_21057,N_21247);
nor U21385 (N_21385,N_21042,N_21153);
nor U21386 (N_21386,N_21186,N_21239);
xor U21387 (N_21387,N_21210,N_21046);
nor U21388 (N_21388,N_21087,N_21214);
nand U21389 (N_21389,N_21052,N_21071);
nor U21390 (N_21390,N_21041,N_21193);
nor U21391 (N_21391,N_21033,N_21143);
and U21392 (N_21392,N_21154,N_21132);
and U21393 (N_21393,N_21225,N_21209);
and U21394 (N_21394,N_21187,N_21128);
and U21395 (N_21395,N_21033,N_21026);
nand U21396 (N_21396,N_21234,N_21066);
nand U21397 (N_21397,N_21072,N_21081);
nand U21398 (N_21398,N_21244,N_21060);
nand U21399 (N_21399,N_21121,N_21199);
and U21400 (N_21400,N_21083,N_21009);
nor U21401 (N_21401,N_21032,N_21243);
xnor U21402 (N_21402,N_21147,N_21203);
or U21403 (N_21403,N_21203,N_21034);
or U21404 (N_21404,N_21212,N_21151);
xnor U21405 (N_21405,N_21135,N_21228);
and U21406 (N_21406,N_21222,N_21111);
and U21407 (N_21407,N_21006,N_21029);
or U21408 (N_21408,N_21102,N_21216);
or U21409 (N_21409,N_21044,N_21115);
or U21410 (N_21410,N_21012,N_21105);
nor U21411 (N_21411,N_21142,N_21111);
or U21412 (N_21412,N_21163,N_21044);
or U21413 (N_21413,N_21231,N_21018);
and U21414 (N_21414,N_21119,N_21113);
or U21415 (N_21415,N_21107,N_21037);
and U21416 (N_21416,N_21004,N_21067);
or U21417 (N_21417,N_21239,N_21229);
xnor U21418 (N_21418,N_21137,N_21247);
or U21419 (N_21419,N_21014,N_21080);
xnor U21420 (N_21420,N_21249,N_21141);
xnor U21421 (N_21421,N_21240,N_21245);
nand U21422 (N_21422,N_21180,N_21131);
or U21423 (N_21423,N_21143,N_21036);
nand U21424 (N_21424,N_21140,N_21209);
and U21425 (N_21425,N_21129,N_21246);
nand U21426 (N_21426,N_21018,N_21073);
or U21427 (N_21427,N_21036,N_21187);
or U21428 (N_21428,N_21003,N_21110);
or U21429 (N_21429,N_21108,N_21218);
and U21430 (N_21430,N_21036,N_21120);
xnor U21431 (N_21431,N_21216,N_21206);
or U21432 (N_21432,N_21116,N_21060);
or U21433 (N_21433,N_21098,N_21087);
nor U21434 (N_21434,N_21196,N_21217);
nor U21435 (N_21435,N_21057,N_21018);
xnor U21436 (N_21436,N_21235,N_21206);
nor U21437 (N_21437,N_21062,N_21027);
or U21438 (N_21438,N_21233,N_21172);
or U21439 (N_21439,N_21224,N_21140);
or U21440 (N_21440,N_21161,N_21043);
and U21441 (N_21441,N_21196,N_21210);
nor U21442 (N_21442,N_21072,N_21076);
and U21443 (N_21443,N_21090,N_21116);
or U21444 (N_21444,N_21138,N_21235);
nor U21445 (N_21445,N_21180,N_21228);
or U21446 (N_21446,N_21136,N_21035);
nor U21447 (N_21447,N_21197,N_21209);
xor U21448 (N_21448,N_21000,N_21192);
xnor U21449 (N_21449,N_21056,N_21054);
nor U21450 (N_21450,N_21016,N_21123);
nand U21451 (N_21451,N_21093,N_21035);
nand U21452 (N_21452,N_21226,N_21116);
nand U21453 (N_21453,N_21089,N_21225);
or U21454 (N_21454,N_21009,N_21140);
nand U21455 (N_21455,N_21166,N_21098);
and U21456 (N_21456,N_21172,N_21043);
xnor U21457 (N_21457,N_21127,N_21015);
nor U21458 (N_21458,N_21052,N_21147);
nand U21459 (N_21459,N_21236,N_21177);
nor U21460 (N_21460,N_21119,N_21100);
nand U21461 (N_21461,N_21160,N_21124);
nand U21462 (N_21462,N_21188,N_21231);
nand U21463 (N_21463,N_21220,N_21004);
nor U21464 (N_21464,N_21080,N_21248);
and U21465 (N_21465,N_21200,N_21204);
nand U21466 (N_21466,N_21106,N_21161);
nor U21467 (N_21467,N_21199,N_21041);
xor U21468 (N_21468,N_21076,N_21030);
nand U21469 (N_21469,N_21037,N_21211);
nor U21470 (N_21470,N_21046,N_21016);
and U21471 (N_21471,N_21096,N_21066);
nor U21472 (N_21472,N_21026,N_21230);
nand U21473 (N_21473,N_21005,N_21131);
nor U21474 (N_21474,N_21133,N_21028);
nor U21475 (N_21475,N_21119,N_21210);
nand U21476 (N_21476,N_21080,N_21046);
or U21477 (N_21477,N_21237,N_21207);
xnor U21478 (N_21478,N_21037,N_21198);
or U21479 (N_21479,N_21001,N_21076);
or U21480 (N_21480,N_21033,N_21040);
and U21481 (N_21481,N_21027,N_21171);
and U21482 (N_21482,N_21085,N_21231);
and U21483 (N_21483,N_21059,N_21129);
nor U21484 (N_21484,N_21027,N_21213);
and U21485 (N_21485,N_21002,N_21069);
xor U21486 (N_21486,N_21073,N_21245);
nand U21487 (N_21487,N_21127,N_21042);
nor U21488 (N_21488,N_21071,N_21145);
and U21489 (N_21489,N_21056,N_21076);
nor U21490 (N_21490,N_21145,N_21221);
or U21491 (N_21491,N_21225,N_21038);
nor U21492 (N_21492,N_21173,N_21223);
nor U21493 (N_21493,N_21111,N_21104);
xor U21494 (N_21494,N_21078,N_21179);
nor U21495 (N_21495,N_21113,N_21057);
nand U21496 (N_21496,N_21031,N_21175);
or U21497 (N_21497,N_21183,N_21102);
nor U21498 (N_21498,N_21090,N_21200);
and U21499 (N_21499,N_21072,N_21053);
xnor U21500 (N_21500,N_21499,N_21336);
nand U21501 (N_21501,N_21391,N_21470);
nor U21502 (N_21502,N_21332,N_21421);
nand U21503 (N_21503,N_21330,N_21275);
or U21504 (N_21504,N_21286,N_21351);
nor U21505 (N_21505,N_21278,N_21405);
xor U21506 (N_21506,N_21316,N_21369);
nor U21507 (N_21507,N_21443,N_21265);
and U21508 (N_21508,N_21495,N_21374);
and U21509 (N_21509,N_21429,N_21488);
nor U21510 (N_21510,N_21462,N_21385);
and U21511 (N_21511,N_21306,N_21367);
or U21512 (N_21512,N_21277,N_21494);
nand U21513 (N_21513,N_21445,N_21427);
or U21514 (N_21514,N_21423,N_21304);
or U21515 (N_21515,N_21381,N_21363);
xnor U21516 (N_21516,N_21435,N_21296);
and U21517 (N_21517,N_21279,N_21409);
xnor U21518 (N_21518,N_21475,N_21344);
and U21519 (N_21519,N_21281,N_21384);
or U21520 (N_21520,N_21284,N_21267);
or U21521 (N_21521,N_21403,N_21297);
or U21522 (N_21522,N_21302,N_21266);
and U21523 (N_21523,N_21342,N_21340);
xnor U21524 (N_21524,N_21473,N_21371);
nand U21525 (N_21525,N_21451,N_21274);
and U21526 (N_21526,N_21411,N_21383);
nor U21527 (N_21527,N_21493,N_21379);
nand U21528 (N_21528,N_21437,N_21280);
nand U21529 (N_21529,N_21386,N_21317);
or U21530 (N_21530,N_21335,N_21366);
or U21531 (N_21531,N_21460,N_21326);
nor U21532 (N_21532,N_21394,N_21431);
or U21533 (N_21533,N_21322,N_21350);
nand U21534 (N_21534,N_21287,N_21273);
or U21535 (N_21535,N_21430,N_21308);
xnor U21536 (N_21536,N_21324,N_21331);
nand U21537 (N_21537,N_21321,N_21390);
nor U21538 (N_21538,N_21492,N_21415);
or U21539 (N_21539,N_21256,N_21270);
nand U21540 (N_21540,N_21455,N_21418);
or U21541 (N_21541,N_21291,N_21404);
nand U21542 (N_21542,N_21444,N_21360);
nor U21543 (N_21543,N_21259,N_21318);
and U21544 (N_21544,N_21257,N_21373);
nor U21545 (N_21545,N_21387,N_21454);
nor U21546 (N_21546,N_21380,N_21433);
or U21547 (N_21547,N_21252,N_21376);
nor U21548 (N_21548,N_21496,N_21292);
or U21549 (N_21549,N_21327,N_21453);
nand U21550 (N_21550,N_21276,N_21424);
or U21551 (N_21551,N_21377,N_21410);
xnor U21552 (N_21552,N_21343,N_21489);
or U21553 (N_21553,N_21354,N_21357);
nand U21554 (N_21554,N_21348,N_21481);
nor U21555 (N_21555,N_21483,N_21255);
nor U21556 (N_21556,N_21485,N_21397);
nand U21557 (N_21557,N_21476,N_21484);
or U21558 (N_21558,N_21300,N_21395);
nor U21559 (N_21559,N_21414,N_21457);
nand U21560 (N_21560,N_21293,N_21434);
nand U21561 (N_21561,N_21378,N_21258);
nand U21562 (N_21562,N_21355,N_21389);
xor U21563 (N_21563,N_21420,N_21312);
nor U21564 (N_21564,N_21400,N_21295);
and U21565 (N_21565,N_21347,N_21364);
and U21566 (N_21566,N_21487,N_21337);
nand U21567 (N_21567,N_21474,N_21345);
and U21568 (N_21568,N_21469,N_21449);
and U21569 (N_21569,N_21283,N_21479);
and U21570 (N_21570,N_21311,N_21352);
and U21571 (N_21571,N_21422,N_21334);
or U21572 (N_21572,N_21353,N_21325);
and U21573 (N_21573,N_21490,N_21254);
xnor U21574 (N_21574,N_21251,N_21468);
or U21575 (N_21575,N_21426,N_21438);
xor U21576 (N_21576,N_21250,N_21467);
or U21577 (N_21577,N_21263,N_21464);
nor U21578 (N_21578,N_21253,N_21362);
xnor U21579 (N_21579,N_21271,N_21328);
xnor U21580 (N_21580,N_21382,N_21465);
or U21581 (N_21581,N_21341,N_21461);
nor U21582 (N_21582,N_21262,N_21448);
nor U21583 (N_21583,N_21272,N_21365);
nor U21584 (N_21584,N_21425,N_21375);
or U21585 (N_21585,N_21333,N_21440);
nand U21586 (N_21586,N_21401,N_21356);
nand U21587 (N_21587,N_21412,N_21269);
nor U21588 (N_21588,N_21456,N_21294);
nor U21589 (N_21589,N_21298,N_21338);
nor U21590 (N_21590,N_21486,N_21303);
xor U21591 (N_21591,N_21310,N_21349);
or U21592 (N_21592,N_21413,N_21313);
nor U21593 (N_21593,N_21299,N_21406);
nor U21594 (N_21594,N_21416,N_21441);
nand U21595 (N_21595,N_21288,N_21320);
and U21596 (N_21596,N_21361,N_21472);
or U21597 (N_21597,N_21466,N_21393);
and U21598 (N_21598,N_21260,N_21319);
nor U21599 (N_21599,N_21264,N_21459);
nor U21600 (N_21600,N_21396,N_21268);
or U21601 (N_21601,N_21478,N_21419);
or U21602 (N_21602,N_21372,N_21282);
or U21603 (N_21603,N_21399,N_21482);
and U21604 (N_21604,N_21498,N_21471);
or U21605 (N_21605,N_21398,N_21439);
nand U21606 (N_21606,N_21309,N_21301);
and U21607 (N_21607,N_21285,N_21370);
or U21608 (N_21608,N_21491,N_21323);
and U21609 (N_21609,N_21480,N_21392);
xor U21610 (N_21610,N_21359,N_21289);
and U21611 (N_21611,N_21315,N_21368);
nor U21612 (N_21612,N_21329,N_21497);
nor U21613 (N_21613,N_21446,N_21314);
xnor U21614 (N_21614,N_21450,N_21436);
nor U21615 (N_21615,N_21447,N_21305);
nor U21616 (N_21616,N_21408,N_21417);
xor U21617 (N_21617,N_21346,N_21442);
nor U21618 (N_21618,N_21358,N_21477);
nor U21619 (N_21619,N_21407,N_21458);
xor U21620 (N_21620,N_21307,N_21428);
nor U21621 (N_21621,N_21402,N_21339);
nor U21622 (N_21622,N_21290,N_21388);
or U21623 (N_21623,N_21463,N_21432);
nand U21624 (N_21624,N_21261,N_21452);
xnor U21625 (N_21625,N_21342,N_21469);
or U21626 (N_21626,N_21312,N_21340);
xor U21627 (N_21627,N_21495,N_21296);
nand U21628 (N_21628,N_21444,N_21413);
nor U21629 (N_21629,N_21295,N_21371);
and U21630 (N_21630,N_21302,N_21345);
and U21631 (N_21631,N_21414,N_21493);
xnor U21632 (N_21632,N_21334,N_21284);
or U21633 (N_21633,N_21455,N_21260);
xor U21634 (N_21634,N_21439,N_21386);
and U21635 (N_21635,N_21471,N_21419);
nand U21636 (N_21636,N_21280,N_21450);
nand U21637 (N_21637,N_21347,N_21303);
or U21638 (N_21638,N_21369,N_21481);
xnor U21639 (N_21639,N_21477,N_21467);
nand U21640 (N_21640,N_21334,N_21380);
and U21641 (N_21641,N_21254,N_21323);
nand U21642 (N_21642,N_21284,N_21499);
nor U21643 (N_21643,N_21344,N_21284);
nor U21644 (N_21644,N_21356,N_21284);
nand U21645 (N_21645,N_21398,N_21253);
and U21646 (N_21646,N_21336,N_21436);
nor U21647 (N_21647,N_21488,N_21333);
xor U21648 (N_21648,N_21479,N_21391);
or U21649 (N_21649,N_21311,N_21340);
and U21650 (N_21650,N_21443,N_21362);
and U21651 (N_21651,N_21325,N_21264);
and U21652 (N_21652,N_21327,N_21458);
or U21653 (N_21653,N_21497,N_21451);
nand U21654 (N_21654,N_21466,N_21406);
nand U21655 (N_21655,N_21461,N_21286);
nand U21656 (N_21656,N_21425,N_21263);
xor U21657 (N_21657,N_21429,N_21265);
and U21658 (N_21658,N_21495,N_21452);
nand U21659 (N_21659,N_21268,N_21403);
nand U21660 (N_21660,N_21411,N_21434);
or U21661 (N_21661,N_21414,N_21367);
and U21662 (N_21662,N_21263,N_21273);
xor U21663 (N_21663,N_21477,N_21421);
xnor U21664 (N_21664,N_21287,N_21473);
xnor U21665 (N_21665,N_21405,N_21403);
xor U21666 (N_21666,N_21413,N_21457);
or U21667 (N_21667,N_21326,N_21253);
and U21668 (N_21668,N_21309,N_21332);
xnor U21669 (N_21669,N_21455,N_21289);
xor U21670 (N_21670,N_21417,N_21411);
nor U21671 (N_21671,N_21465,N_21445);
nand U21672 (N_21672,N_21334,N_21337);
nand U21673 (N_21673,N_21490,N_21425);
nand U21674 (N_21674,N_21265,N_21284);
nand U21675 (N_21675,N_21449,N_21280);
nor U21676 (N_21676,N_21435,N_21404);
nand U21677 (N_21677,N_21422,N_21336);
nor U21678 (N_21678,N_21326,N_21425);
or U21679 (N_21679,N_21427,N_21410);
or U21680 (N_21680,N_21417,N_21462);
xor U21681 (N_21681,N_21315,N_21256);
nand U21682 (N_21682,N_21272,N_21446);
or U21683 (N_21683,N_21421,N_21268);
and U21684 (N_21684,N_21413,N_21280);
and U21685 (N_21685,N_21423,N_21303);
xor U21686 (N_21686,N_21400,N_21364);
nor U21687 (N_21687,N_21361,N_21271);
nor U21688 (N_21688,N_21493,N_21325);
or U21689 (N_21689,N_21295,N_21362);
and U21690 (N_21690,N_21438,N_21429);
or U21691 (N_21691,N_21406,N_21373);
xor U21692 (N_21692,N_21454,N_21463);
or U21693 (N_21693,N_21405,N_21336);
nor U21694 (N_21694,N_21313,N_21296);
nand U21695 (N_21695,N_21256,N_21371);
and U21696 (N_21696,N_21347,N_21471);
xor U21697 (N_21697,N_21434,N_21355);
and U21698 (N_21698,N_21336,N_21311);
nand U21699 (N_21699,N_21428,N_21399);
nand U21700 (N_21700,N_21315,N_21348);
nand U21701 (N_21701,N_21300,N_21408);
and U21702 (N_21702,N_21427,N_21253);
nor U21703 (N_21703,N_21432,N_21487);
and U21704 (N_21704,N_21462,N_21427);
and U21705 (N_21705,N_21432,N_21255);
xor U21706 (N_21706,N_21428,N_21256);
and U21707 (N_21707,N_21352,N_21458);
and U21708 (N_21708,N_21428,N_21450);
nand U21709 (N_21709,N_21433,N_21266);
or U21710 (N_21710,N_21252,N_21425);
or U21711 (N_21711,N_21405,N_21372);
or U21712 (N_21712,N_21302,N_21470);
nand U21713 (N_21713,N_21265,N_21313);
xnor U21714 (N_21714,N_21427,N_21457);
nor U21715 (N_21715,N_21313,N_21366);
xnor U21716 (N_21716,N_21419,N_21442);
nor U21717 (N_21717,N_21441,N_21254);
nor U21718 (N_21718,N_21421,N_21469);
or U21719 (N_21719,N_21291,N_21321);
nand U21720 (N_21720,N_21394,N_21266);
or U21721 (N_21721,N_21406,N_21326);
and U21722 (N_21722,N_21366,N_21343);
and U21723 (N_21723,N_21412,N_21302);
or U21724 (N_21724,N_21252,N_21321);
xor U21725 (N_21725,N_21420,N_21495);
xor U21726 (N_21726,N_21378,N_21470);
nor U21727 (N_21727,N_21293,N_21336);
xor U21728 (N_21728,N_21261,N_21313);
xor U21729 (N_21729,N_21382,N_21352);
and U21730 (N_21730,N_21455,N_21474);
nor U21731 (N_21731,N_21387,N_21467);
and U21732 (N_21732,N_21298,N_21388);
nor U21733 (N_21733,N_21322,N_21430);
nand U21734 (N_21734,N_21251,N_21403);
xor U21735 (N_21735,N_21384,N_21259);
and U21736 (N_21736,N_21304,N_21390);
nor U21737 (N_21737,N_21480,N_21260);
or U21738 (N_21738,N_21333,N_21280);
nand U21739 (N_21739,N_21347,N_21279);
nor U21740 (N_21740,N_21390,N_21292);
nand U21741 (N_21741,N_21449,N_21300);
nor U21742 (N_21742,N_21370,N_21473);
or U21743 (N_21743,N_21291,N_21392);
xnor U21744 (N_21744,N_21410,N_21296);
and U21745 (N_21745,N_21408,N_21428);
nand U21746 (N_21746,N_21407,N_21474);
or U21747 (N_21747,N_21454,N_21378);
and U21748 (N_21748,N_21316,N_21288);
xor U21749 (N_21749,N_21282,N_21489);
and U21750 (N_21750,N_21657,N_21707);
and U21751 (N_21751,N_21741,N_21747);
or U21752 (N_21752,N_21608,N_21711);
nor U21753 (N_21753,N_21739,N_21651);
nand U21754 (N_21754,N_21700,N_21592);
nor U21755 (N_21755,N_21639,N_21577);
xor U21756 (N_21756,N_21602,N_21599);
and U21757 (N_21757,N_21656,N_21712);
and U21758 (N_21758,N_21718,N_21648);
xnor U21759 (N_21759,N_21525,N_21562);
nand U21760 (N_21760,N_21686,N_21553);
or U21761 (N_21761,N_21542,N_21566);
or U21762 (N_21762,N_21728,N_21568);
or U21763 (N_21763,N_21575,N_21505);
nand U21764 (N_21764,N_21719,N_21581);
and U21765 (N_21765,N_21646,N_21604);
or U21766 (N_21766,N_21501,N_21723);
or U21767 (N_21767,N_21538,N_21622);
xor U21768 (N_21768,N_21563,N_21669);
nor U21769 (N_21769,N_21742,N_21716);
or U21770 (N_21770,N_21559,N_21614);
nor U21771 (N_21771,N_21515,N_21605);
or U21772 (N_21772,N_21603,N_21724);
nand U21773 (N_21773,N_21694,N_21612);
nand U21774 (N_21774,N_21520,N_21607);
and U21775 (N_21775,N_21737,N_21643);
or U21776 (N_21776,N_21615,N_21660);
or U21777 (N_21777,N_21541,N_21588);
nand U21778 (N_21778,N_21658,N_21600);
nand U21779 (N_21779,N_21654,N_21572);
and U21780 (N_21780,N_21632,N_21531);
nor U21781 (N_21781,N_21672,N_21726);
or U21782 (N_21782,N_21578,N_21703);
and U21783 (N_21783,N_21667,N_21624);
and U21784 (N_21784,N_21552,N_21674);
nor U21785 (N_21785,N_21571,N_21540);
or U21786 (N_21786,N_21611,N_21635);
xor U21787 (N_21787,N_21693,N_21625);
and U21788 (N_21788,N_21734,N_21670);
and U21789 (N_21789,N_21616,N_21731);
xnor U21790 (N_21790,N_21629,N_21543);
nor U21791 (N_21791,N_21699,N_21527);
or U21792 (N_21792,N_21579,N_21630);
nand U21793 (N_21793,N_21606,N_21587);
nor U21794 (N_21794,N_21627,N_21685);
xnor U21795 (N_21795,N_21659,N_21744);
nand U21796 (N_21796,N_21601,N_21597);
nand U21797 (N_21797,N_21545,N_21702);
and U21798 (N_21798,N_21569,N_21655);
nor U21799 (N_21799,N_21596,N_21555);
xnor U21800 (N_21800,N_21508,N_21560);
or U21801 (N_21801,N_21585,N_21595);
or U21802 (N_21802,N_21690,N_21749);
or U21803 (N_21803,N_21500,N_21536);
and U21804 (N_21804,N_21636,N_21677);
xor U21805 (N_21805,N_21637,N_21547);
xor U21806 (N_21806,N_21633,N_21745);
nand U21807 (N_21807,N_21705,N_21692);
and U21808 (N_21808,N_21729,N_21590);
nand U21809 (N_21809,N_21518,N_21556);
or U21810 (N_21810,N_21710,N_21638);
and U21811 (N_21811,N_21521,N_21610);
or U21812 (N_21812,N_21671,N_21583);
and U21813 (N_21813,N_21539,N_21619);
nor U21814 (N_21814,N_21589,N_21652);
nand U21815 (N_21815,N_21725,N_21668);
nor U21816 (N_21816,N_21598,N_21551);
nor U21817 (N_21817,N_21529,N_21537);
and U21818 (N_21818,N_21512,N_21550);
and U21819 (N_21819,N_21573,N_21675);
nor U21820 (N_21820,N_21628,N_21682);
nor U21821 (N_21821,N_21663,N_21748);
xnor U21822 (N_21822,N_21733,N_21673);
nor U21823 (N_21823,N_21696,N_21664);
xor U21824 (N_21824,N_21634,N_21691);
nor U21825 (N_21825,N_21684,N_21662);
xnor U21826 (N_21826,N_21558,N_21620);
and U21827 (N_21827,N_21535,N_21511);
xnor U21828 (N_21828,N_21546,N_21576);
or U21829 (N_21829,N_21516,N_21704);
and U21830 (N_21830,N_21514,N_21644);
nor U21831 (N_21831,N_21513,N_21736);
and U21832 (N_21832,N_21641,N_21567);
xor U21833 (N_21833,N_21532,N_21591);
nand U21834 (N_21834,N_21502,N_21526);
and U21835 (N_21835,N_21594,N_21561);
nor U21836 (N_21836,N_21683,N_21649);
or U21837 (N_21837,N_21510,N_21701);
and U21838 (N_21838,N_21695,N_21676);
xnor U21839 (N_21839,N_21661,N_21680);
nand U21840 (N_21840,N_21743,N_21609);
or U21841 (N_21841,N_21689,N_21507);
or U21842 (N_21842,N_21582,N_21557);
and U21843 (N_21843,N_21697,N_21640);
nor U21844 (N_21844,N_21530,N_21717);
and U21845 (N_21845,N_21580,N_21746);
and U21846 (N_21846,N_21714,N_21544);
xnor U21847 (N_21847,N_21618,N_21735);
xnor U21848 (N_21848,N_21523,N_21650);
xnor U21849 (N_21849,N_21653,N_21548);
nor U21850 (N_21850,N_21715,N_21738);
xor U21851 (N_21851,N_21574,N_21666);
nand U21852 (N_21852,N_21631,N_21713);
nand U21853 (N_21853,N_21570,N_21681);
xor U21854 (N_21854,N_21554,N_21730);
nand U21855 (N_21855,N_21534,N_21688);
nand U21856 (N_21856,N_21509,N_21506);
nor U21857 (N_21857,N_21549,N_21564);
and U21858 (N_21858,N_21621,N_21647);
or U21859 (N_21859,N_21533,N_21586);
xnor U21860 (N_21860,N_21623,N_21687);
xnor U21861 (N_21861,N_21565,N_21722);
and U21862 (N_21862,N_21706,N_21740);
nor U21863 (N_21863,N_21617,N_21698);
nor U21864 (N_21864,N_21524,N_21626);
or U21865 (N_21865,N_21503,N_21665);
nor U21866 (N_21866,N_21584,N_21519);
or U21867 (N_21867,N_21720,N_21708);
nor U21868 (N_21868,N_21678,N_21517);
nor U21869 (N_21869,N_21645,N_21642);
nand U21870 (N_21870,N_21727,N_21732);
xor U21871 (N_21871,N_21528,N_21613);
nand U21872 (N_21872,N_21504,N_21679);
and U21873 (N_21873,N_21709,N_21593);
nor U21874 (N_21874,N_21721,N_21522);
and U21875 (N_21875,N_21718,N_21541);
or U21876 (N_21876,N_21631,N_21603);
xnor U21877 (N_21877,N_21580,N_21597);
or U21878 (N_21878,N_21566,N_21614);
or U21879 (N_21879,N_21515,N_21576);
nand U21880 (N_21880,N_21538,N_21690);
or U21881 (N_21881,N_21547,N_21726);
or U21882 (N_21882,N_21642,N_21585);
nor U21883 (N_21883,N_21695,N_21598);
and U21884 (N_21884,N_21656,N_21737);
nand U21885 (N_21885,N_21708,N_21600);
nand U21886 (N_21886,N_21644,N_21743);
or U21887 (N_21887,N_21638,N_21640);
xnor U21888 (N_21888,N_21593,N_21744);
or U21889 (N_21889,N_21532,N_21590);
nand U21890 (N_21890,N_21557,N_21680);
xor U21891 (N_21891,N_21702,N_21716);
nor U21892 (N_21892,N_21606,N_21554);
nand U21893 (N_21893,N_21645,N_21501);
or U21894 (N_21894,N_21729,N_21608);
nand U21895 (N_21895,N_21701,N_21573);
nor U21896 (N_21896,N_21632,N_21525);
or U21897 (N_21897,N_21628,N_21687);
and U21898 (N_21898,N_21596,N_21691);
nor U21899 (N_21899,N_21500,N_21686);
nand U21900 (N_21900,N_21638,N_21613);
nand U21901 (N_21901,N_21631,N_21539);
nor U21902 (N_21902,N_21530,N_21670);
or U21903 (N_21903,N_21634,N_21670);
nor U21904 (N_21904,N_21710,N_21709);
xnor U21905 (N_21905,N_21725,N_21629);
nor U21906 (N_21906,N_21681,N_21642);
nand U21907 (N_21907,N_21643,N_21729);
xor U21908 (N_21908,N_21640,N_21739);
and U21909 (N_21909,N_21647,N_21508);
or U21910 (N_21910,N_21679,N_21686);
nand U21911 (N_21911,N_21598,N_21514);
and U21912 (N_21912,N_21610,N_21546);
nand U21913 (N_21913,N_21581,N_21532);
and U21914 (N_21914,N_21641,N_21543);
xnor U21915 (N_21915,N_21593,N_21705);
xnor U21916 (N_21916,N_21524,N_21519);
or U21917 (N_21917,N_21736,N_21518);
or U21918 (N_21918,N_21656,N_21609);
and U21919 (N_21919,N_21699,N_21655);
nand U21920 (N_21920,N_21694,N_21610);
nor U21921 (N_21921,N_21663,N_21585);
nor U21922 (N_21922,N_21675,N_21510);
and U21923 (N_21923,N_21624,N_21662);
xor U21924 (N_21924,N_21502,N_21671);
nand U21925 (N_21925,N_21631,N_21530);
xor U21926 (N_21926,N_21636,N_21501);
xor U21927 (N_21927,N_21508,N_21637);
or U21928 (N_21928,N_21579,N_21509);
xnor U21929 (N_21929,N_21524,N_21610);
and U21930 (N_21930,N_21554,N_21551);
nand U21931 (N_21931,N_21658,N_21696);
or U21932 (N_21932,N_21556,N_21572);
xnor U21933 (N_21933,N_21522,N_21516);
nor U21934 (N_21934,N_21566,N_21606);
or U21935 (N_21935,N_21593,N_21528);
nand U21936 (N_21936,N_21743,N_21642);
and U21937 (N_21937,N_21602,N_21690);
and U21938 (N_21938,N_21646,N_21747);
or U21939 (N_21939,N_21746,N_21688);
and U21940 (N_21940,N_21623,N_21616);
nand U21941 (N_21941,N_21626,N_21591);
or U21942 (N_21942,N_21584,N_21676);
or U21943 (N_21943,N_21612,N_21531);
nand U21944 (N_21944,N_21709,N_21517);
or U21945 (N_21945,N_21706,N_21707);
xnor U21946 (N_21946,N_21503,N_21613);
or U21947 (N_21947,N_21737,N_21715);
nand U21948 (N_21948,N_21629,N_21685);
xor U21949 (N_21949,N_21652,N_21702);
xor U21950 (N_21950,N_21612,N_21688);
nand U21951 (N_21951,N_21580,N_21639);
or U21952 (N_21952,N_21654,N_21729);
nor U21953 (N_21953,N_21537,N_21592);
nor U21954 (N_21954,N_21673,N_21682);
or U21955 (N_21955,N_21717,N_21542);
nor U21956 (N_21956,N_21668,N_21596);
nand U21957 (N_21957,N_21619,N_21536);
nand U21958 (N_21958,N_21551,N_21737);
xnor U21959 (N_21959,N_21723,N_21643);
nand U21960 (N_21960,N_21528,N_21686);
nand U21961 (N_21961,N_21639,N_21640);
nand U21962 (N_21962,N_21511,N_21553);
xor U21963 (N_21963,N_21647,N_21711);
or U21964 (N_21964,N_21556,N_21655);
and U21965 (N_21965,N_21525,N_21546);
and U21966 (N_21966,N_21734,N_21563);
and U21967 (N_21967,N_21539,N_21607);
xor U21968 (N_21968,N_21595,N_21649);
and U21969 (N_21969,N_21519,N_21710);
nor U21970 (N_21970,N_21513,N_21504);
xnor U21971 (N_21971,N_21672,N_21606);
and U21972 (N_21972,N_21542,N_21524);
and U21973 (N_21973,N_21504,N_21534);
xor U21974 (N_21974,N_21585,N_21587);
xor U21975 (N_21975,N_21697,N_21522);
or U21976 (N_21976,N_21556,N_21594);
and U21977 (N_21977,N_21557,N_21656);
xor U21978 (N_21978,N_21552,N_21581);
or U21979 (N_21979,N_21694,N_21507);
xnor U21980 (N_21980,N_21735,N_21659);
or U21981 (N_21981,N_21564,N_21706);
or U21982 (N_21982,N_21574,N_21587);
nor U21983 (N_21983,N_21737,N_21511);
and U21984 (N_21984,N_21575,N_21536);
nor U21985 (N_21985,N_21653,N_21606);
or U21986 (N_21986,N_21601,N_21589);
or U21987 (N_21987,N_21615,N_21592);
or U21988 (N_21988,N_21724,N_21516);
or U21989 (N_21989,N_21643,N_21649);
nor U21990 (N_21990,N_21633,N_21643);
xnor U21991 (N_21991,N_21596,N_21677);
and U21992 (N_21992,N_21711,N_21526);
nor U21993 (N_21993,N_21681,N_21685);
nor U21994 (N_21994,N_21611,N_21745);
nand U21995 (N_21995,N_21598,N_21518);
or U21996 (N_21996,N_21648,N_21733);
xor U21997 (N_21997,N_21573,N_21687);
and U21998 (N_21998,N_21603,N_21686);
or U21999 (N_21999,N_21604,N_21678);
nand U22000 (N_22000,N_21763,N_21869);
and U22001 (N_22001,N_21851,N_21778);
and U22002 (N_22002,N_21895,N_21911);
nor U22003 (N_22003,N_21910,N_21948);
and U22004 (N_22004,N_21986,N_21962);
nand U22005 (N_22005,N_21881,N_21825);
nor U22006 (N_22006,N_21921,N_21788);
and U22007 (N_22007,N_21859,N_21956);
xnor U22008 (N_22008,N_21958,N_21949);
nand U22009 (N_22009,N_21840,N_21953);
nor U22010 (N_22010,N_21929,N_21753);
and U22011 (N_22011,N_21812,N_21944);
nor U22012 (N_22012,N_21837,N_21978);
or U22013 (N_22013,N_21992,N_21764);
and U22014 (N_22014,N_21931,N_21789);
and U22015 (N_22015,N_21920,N_21977);
nand U22016 (N_22016,N_21793,N_21782);
or U22017 (N_22017,N_21967,N_21896);
nand U22018 (N_22018,N_21892,N_21796);
nand U22019 (N_22019,N_21885,N_21824);
and U22020 (N_22020,N_21987,N_21762);
or U22021 (N_22021,N_21932,N_21976);
xor U22022 (N_22022,N_21807,N_21844);
xnor U22023 (N_22023,N_21783,N_21871);
nand U22024 (N_22024,N_21898,N_21854);
xnor U22025 (N_22025,N_21902,N_21882);
and U22026 (N_22026,N_21817,N_21918);
nand U22027 (N_22027,N_21959,N_21755);
and U22028 (N_22028,N_21880,N_21803);
and U22029 (N_22029,N_21974,N_21985);
nand U22030 (N_22030,N_21815,N_21914);
and U22031 (N_22031,N_21969,N_21973);
nor U22032 (N_22032,N_21846,N_21894);
or U22033 (N_22033,N_21877,N_21960);
nand U22034 (N_22034,N_21954,N_21774);
nor U22035 (N_22035,N_21759,N_21820);
or U22036 (N_22036,N_21994,N_21757);
nand U22037 (N_22037,N_21988,N_21845);
nor U22038 (N_22038,N_21831,N_21769);
or U22039 (N_22039,N_21756,N_21795);
nor U22040 (N_22040,N_21772,N_21883);
xor U22041 (N_22041,N_21773,N_21775);
and U22042 (N_22042,N_21804,N_21760);
or U22043 (N_22043,N_21916,N_21945);
xor U22044 (N_22044,N_21938,N_21968);
or U22045 (N_22045,N_21850,N_21990);
nand U22046 (N_22046,N_21867,N_21903);
nand U22047 (N_22047,N_21779,N_21981);
nand U22048 (N_22048,N_21873,N_21843);
nand U22049 (N_22049,N_21842,N_21876);
or U22050 (N_22050,N_21865,N_21800);
nand U22051 (N_22051,N_21951,N_21848);
xnor U22052 (N_22052,N_21947,N_21889);
nand U22053 (N_22053,N_21887,N_21982);
nand U22054 (N_22054,N_21868,N_21808);
nor U22055 (N_22055,N_21856,N_21901);
nand U22056 (N_22056,N_21835,N_21776);
and U22057 (N_22057,N_21847,N_21765);
or U22058 (N_22058,N_21770,N_21863);
nor U22059 (N_22059,N_21907,N_21830);
and U22060 (N_22060,N_21946,N_21975);
nand U22061 (N_22061,N_21899,N_21879);
xor U22062 (N_22062,N_21943,N_21838);
or U22063 (N_22063,N_21936,N_21833);
nand U22064 (N_22064,N_21852,N_21829);
nand U22065 (N_22065,N_21821,N_21926);
and U22066 (N_22066,N_21905,N_21754);
nand U22067 (N_22067,N_21792,N_21997);
nand U22068 (N_22068,N_21878,N_21802);
nor U22069 (N_22069,N_21891,N_21853);
nand U22070 (N_22070,N_21798,N_21771);
xor U22071 (N_22071,N_21874,N_21836);
and U22072 (N_22072,N_21940,N_21816);
or U22073 (N_22073,N_21781,N_21766);
nand U22074 (N_22074,N_21928,N_21989);
xor U22075 (N_22075,N_21827,N_21806);
xnor U22076 (N_22076,N_21758,N_21991);
nand U22077 (N_22077,N_21979,N_21915);
or U22078 (N_22078,N_21998,N_21791);
nor U22079 (N_22079,N_21797,N_21858);
and U22080 (N_22080,N_21906,N_21884);
nor U22081 (N_22081,N_21750,N_21950);
nor U22082 (N_22082,N_21924,N_21866);
or U22083 (N_22083,N_21923,N_21900);
and U22084 (N_22084,N_21875,N_21805);
nand U22085 (N_22085,N_21857,N_21955);
nand U22086 (N_22086,N_21813,N_21855);
nand U22087 (N_22087,N_21768,N_21849);
and U22088 (N_22088,N_21909,N_21925);
nor U22089 (N_22089,N_21939,N_21993);
or U22090 (N_22090,N_21966,N_21886);
nor U22091 (N_22091,N_21786,N_21908);
xor U22092 (N_22092,N_21935,N_21818);
nand U22093 (N_22093,N_21961,N_21922);
nand U22094 (N_22094,N_21934,N_21784);
nor U22095 (N_22095,N_21777,N_21927);
xor U22096 (N_22096,N_21794,N_21823);
or U22097 (N_22097,N_21761,N_21767);
nand U22098 (N_22098,N_21860,N_21893);
nand U22099 (N_22099,N_21828,N_21930);
or U22100 (N_22100,N_21822,N_21919);
nand U22101 (N_22101,N_21984,N_21752);
nor U22102 (N_22102,N_21864,N_21913);
or U22103 (N_22103,N_21861,N_21963);
nor U22104 (N_22104,N_21888,N_21952);
nor U22105 (N_22105,N_21751,N_21970);
nand U22106 (N_22106,N_21799,N_21780);
nand U22107 (N_22107,N_21942,N_21999);
nor U22108 (N_22108,N_21964,N_21832);
xnor U22109 (N_22109,N_21995,N_21790);
and U22110 (N_22110,N_21870,N_21965);
nand U22111 (N_22111,N_21912,N_21814);
or U22112 (N_22112,N_21841,N_21983);
and U22113 (N_22113,N_21897,N_21980);
nor U22114 (N_22114,N_21834,N_21996);
nor U22115 (N_22115,N_21839,N_21957);
nand U22116 (N_22116,N_21862,N_21872);
and U22117 (N_22117,N_21787,N_21809);
nor U22118 (N_22118,N_21941,N_21811);
or U22119 (N_22119,N_21972,N_21819);
and U22120 (N_22120,N_21937,N_21917);
or U22121 (N_22121,N_21810,N_21890);
xnor U22122 (N_22122,N_21801,N_21826);
nor U22123 (N_22123,N_21933,N_21904);
nand U22124 (N_22124,N_21785,N_21971);
nor U22125 (N_22125,N_21826,N_21872);
and U22126 (N_22126,N_21951,N_21907);
nor U22127 (N_22127,N_21891,N_21782);
nand U22128 (N_22128,N_21761,N_21791);
nor U22129 (N_22129,N_21902,N_21827);
or U22130 (N_22130,N_21993,N_21969);
nand U22131 (N_22131,N_21797,N_21946);
or U22132 (N_22132,N_21877,N_21861);
or U22133 (N_22133,N_21792,N_21943);
nand U22134 (N_22134,N_21864,N_21927);
or U22135 (N_22135,N_21927,N_21800);
or U22136 (N_22136,N_21790,N_21778);
nand U22137 (N_22137,N_21915,N_21868);
nor U22138 (N_22138,N_21755,N_21811);
and U22139 (N_22139,N_21981,N_21947);
nor U22140 (N_22140,N_21807,N_21753);
and U22141 (N_22141,N_21875,N_21856);
nand U22142 (N_22142,N_21864,N_21807);
nor U22143 (N_22143,N_21947,N_21877);
and U22144 (N_22144,N_21827,N_21936);
nor U22145 (N_22145,N_21942,N_21969);
nor U22146 (N_22146,N_21858,N_21764);
xor U22147 (N_22147,N_21750,N_21887);
or U22148 (N_22148,N_21866,N_21907);
nand U22149 (N_22149,N_21852,N_21969);
xor U22150 (N_22150,N_21830,N_21996);
nand U22151 (N_22151,N_21839,N_21809);
nor U22152 (N_22152,N_21854,N_21988);
and U22153 (N_22153,N_21962,N_21814);
nand U22154 (N_22154,N_21947,N_21790);
nor U22155 (N_22155,N_21772,N_21845);
or U22156 (N_22156,N_21802,N_21848);
nor U22157 (N_22157,N_21936,N_21760);
nand U22158 (N_22158,N_21800,N_21991);
xor U22159 (N_22159,N_21904,N_21966);
or U22160 (N_22160,N_21969,N_21832);
nand U22161 (N_22161,N_21852,N_21779);
or U22162 (N_22162,N_21785,N_21837);
xor U22163 (N_22163,N_21861,N_21802);
or U22164 (N_22164,N_21872,N_21775);
xor U22165 (N_22165,N_21970,N_21875);
and U22166 (N_22166,N_21926,N_21819);
xnor U22167 (N_22167,N_21789,N_21861);
nand U22168 (N_22168,N_21941,N_21979);
nor U22169 (N_22169,N_21849,N_21964);
nor U22170 (N_22170,N_21906,N_21820);
or U22171 (N_22171,N_21797,N_21864);
or U22172 (N_22172,N_21965,N_21944);
nand U22173 (N_22173,N_21992,N_21875);
or U22174 (N_22174,N_21912,N_21956);
or U22175 (N_22175,N_21775,N_21893);
or U22176 (N_22176,N_21765,N_21947);
nor U22177 (N_22177,N_21918,N_21775);
nand U22178 (N_22178,N_21986,N_21840);
nand U22179 (N_22179,N_21891,N_21761);
xnor U22180 (N_22180,N_21995,N_21917);
xor U22181 (N_22181,N_21950,N_21805);
xnor U22182 (N_22182,N_21865,N_21952);
xor U22183 (N_22183,N_21960,N_21939);
or U22184 (N_22184,N_21802,N_21787);
xnor U22185 (N_22185,N_21876,N_21863);
nand U22186 (N_22186,N_21938,N_21778);
xor U22187 (N_22187,N_21940,N_21920);
nor U22188 (N_22188,N_21978,N_21876);
nand U22189 (N_22189,N_21907,N_21998);
and U22190 (N_22190,N_21773,N_21812);
nand U22191 (N_22191,N_21838,N_21882);
or U22192 (N_22192,N_21991,N_21774);
xor U22193 (N_22193,N_21963,N_21810);
or U22194 (N_22194,N_21811,N_21766);
or U22195 (N_22195,N_21894,N_21886);
nor U22196 (N_22196,N_21939,N_21874);
nand U22197 (N_22197,N_21962,N_21906);
or U22198 (N_22198,N_21909,N_21877);
and U22199 (N_22199,N_21805,N_21976);
nor U22200 (N_22200,N_21786,N_21938);
xnor U22201 (N_22201,N_21883,N_21787);
nand U22202 (N_22202,N_21832,N_21916);
nor U22203 (N_22203,N_21820,N_21776);
and U22204 (N_22204,N_21840,N_21981);
nand U22205 (N_22205,N_21972,N_21909);
nand U22206 (N_22206,N_21815,N_21873);
nor U22207 (N_22207,N_21949,N_21966);
xor U22208 (N_22208,N_21765,N_21992);
and U22209 (N_22209,N_21866,N_21925);
and U22210 (N_22210,N_21755,N_21890);
and U22211 (N_22211,N_21777,N_21889);
nand U22212 (N_22212,N_21936,N_21985);
xor U22213 (N_22213,N_21815,N_21927);
xor U22214 (N_22214,N_21919,N_21760);
or U22215 (N_22215,N_21855,N_21840);
or U22216 (N_22216,N_21798,N_21866);
xnor U22217 (N_22217,N_21962,N_21931);
nand U22218 (N_22218,N_21893,N_21902);
nand U22219 (N_22219,N_21972,N_21776);
or U22220 (N_22220,N_21972,N_21880);
and U22221 (N_22221,N_21869,N_21981);
nor U22222 (N_22222,N_21851,N_21971);
or U22223 (N_22223,N_21914,N_21840);
xor U22224 (N_22224,N_21954,N_21940);
or U22225 (N_22225,N_21877,N_21840);
nor U22226 (N_22226,N_21790,N_21866);
nor U22227 (N_22227,N_21998,N_21989);
nor U22228 (N_22228,N_21945,N_21806);
nand U22229 (N_22229,N_21807,N_21955);
xor U22230 (N_22230,N_21751,N_21779);
nor U22231 (N_22231,N_21787,N_21936);
or U22232 (N_22232,N_21813,N_21807);
and U22233 (N_22233,N_21839,N_21949);
xor U22234 (N_22234,N_21796,N_21787);
and U22235 (N_22235,N_21773,N_21924);
nor U22236 (N_22236,N_21947,N_21847);
and U22237 (N_22237,N_21814,N_21792);
nor U22238 (N_22238,N_21817,N_21932);
or U22239 (N_22239,N_21779,N_21963);
nand U22240 (N_22240,N_21830,N_21942);
and U22241 (N_22241,N_21965,N_21925);
and U22242 (N_22242,N_21854,N_21857);
and U22243 (N_22243,N_21832,N_21792);
xor U22244 (N_22244,N_21895,N_21865);
nor U22245 (N_22245,N_21915,N_21763);
and U22246 (N_22246,N_21754,N_21837);
or U22247 (N_22247,N_21763,N_21925);
nand U22248 (N_22248,N_21858,N_21788);
xnor U22249 (N_22249,N_21997,N_21968);
nor U22250 (N_22250,N_22222,N_22129);
nand U22251 (N_22251,N_22115,N_22176);
and U22252 (N_22252,N_22242,N_22118);
or U22253 (N_22253,N_22223,N_22019);
and U22254 (N_22254,N_22010,N_22091);
nor U22255 (N_22255,N_22026,N_22138);
nor U22256 (N_22256,N_22191,N_22024);
nand U22257 (N_22257,N_22113,N_22128);
xor U22258 (N_22258,N_22066,N_22043);
or U22259 (N_22259,N_22062,N_22081);
or U22260 (N_22260,N_22084,N_22224);
nand U22261 (N_22261,N_22053,N_22049);
nor U22262 (N_22262,N_22007,N_22188);
and U22263 (N_22263,N_22092,N_22199);
xnor U22264 (N_22264,N_22204,N_22239);
nor U22265 (N_22265,N_22123,N_22104);
xnor U22266 (N_22266,N_22107,N_22217);
nor U22267 (N_22267,N_22187,N_22087);
nand U22268 (N_22268,N_22042,N_22126);
or U22269 (N_22269,N_22121,N_22082);
nor U22270 (N_22270,N_22073,N_22040);
xnor U22271 (N_22271,N_22150,N_22172);
and U22272 (N_22272,N_22000,N_22016);
or U22273 (N_22273,N_22094,N_22100);
nand U22274 (N_22274,N_22200,N_22205);
xnor U22275 (N_22275,N_22163,N_22028);
nor U22276 (N_22276,N_22075,N_22157);
nand U22277 (N_22277,N_22167,N_22122);
and U22278 (N_22278,N_22106,N_22111);
and U22279 (N_22279,N_22011,N_22041);
and U22280 (N_22280,N_22018,N_22056);
nor U22281 (N_22281,N_22114,N_22022);
nand U22282 (N_22282,N_22141,N_22186);
or U22283 (N_22283,N_22211,N_22076);
or U22284 (N_22284,N_22185,N_22183);
and U22285 (N_22285,N_22130,N_22153);
nor U22286 (N_22286,N_22021,N_22063);
nor U22287 (N_22287,N_22203,N_22144);
xnor U22288 (N_22288,N_22055,N_22212);
and U22289 (N_22289,N_22101,N_22072);
and U22290 (N_22290,N_22168,N_22093);
nor U22291 (N_22291,N_22248,N_22231);
nand U22292 (N_22292,N_22109,N_22232);
nand U22293 (N_22293,N_22182,N_22083);
or U22294 (N_22294,N_22177,N_22152);
or U22295 (N_22295,N_22134,N_22173);
xor U22296 (N_22296,N_22050,N_22038);
and U22297 (N_22297,N_22181,N_22192);
nor U22298 (N_22298,N_22164,N_22034);
or U22299 (N_22299,N_22120,N_22090);
and U22300 (N_22300,N_22061,N_22238);
nor U22301 (N_22301,N_22003,N_22029);
and U22302 (N_22302,N_22229,N_22135);
or U22303 (N_22303,N_22088,N_22015);
nor U22304 (N_22304,N_22046,N_22098);
or U22305 (N_22305,N_22190,N_22033);
and U22306 (N_22306,N_22160,N_22099);
and U22307 (N_22307,N_22161,N_22154);
and U22308 (N_22308,N_22193,N_22180);
nor U22309 (N_22309,N_22236,N_22143);
and U22310 (N_22310,N_22149,N_22105);
or U22311 (N_22311,N_22095,N_22045);
and U22312 (N_22312,N_22097,N_22071);
or U22313 (N_22313,N_22039,N_22174);
nor U22314 (N_22314,N_22060,N_22155);
nor U22315 (N_22315,N_22175,N_22233);
nand U22316 (N_22316,N_22027,N_22245);
nor U22317 (N_22317,N_22179,N_22080);
nor U22318 (N_22318,N_22035,N_22156);
xnor U22319 (N_22319,N_22009,N_22057);
or U22320 (N_22320,N_22201,N_22218);
xor U22321 (N_22321,N_22228,N_22131);
and U22322 (N_22322,N_22103,N_22146);
nor U22323 (N_22323,N_22208,N_22032);
nor U22324 (N_22324,N_22124,N_22147);
or U22325 (N_22325,N_22221,N_22012);
or U22326 (N_22326,N_22006,N_22165);
xor U22327 (N_22327,N_22184,N_22102);
nand U22328 (N_22328,N_22044,N_22202);
and U22329 (N_22329,N_22210,N_22078);
xor U22330 (N_22330,N_22225,N_22158);
nand U22331 (N_22331,N_22030,N_22085);
nor U22332 (N_22332,N_22089,N_22142);
nand U22333 (N_22333,N_22117,N_22133);
nand U22334 (N_22334,N_22137,N_22214);
and U22335 (N_22335,N_22001,N_22054);
or U22336 (N_22336,N_22206,N_22079);
nand U22337 (N_22337,N_22059,N_22148);
and U22338 (N_22338,N_22220,N_22178);
and U22339 (N_22339,N_22025,N_22096);
xor U22340 (N_22340,N_22132,N_22215);
nand U22341 (N_22341,N_22159,N_22207);
and U22342 (N_22342,N_22145,N_22197);
or U22343 (N_22343,N_22068,N_22031);
nand U22344 (N_22344,N_22125,N_22070);
or U22345 (N_22345,N_22244,N_22008);
and U22346 (N_22346,N_22086,N_22213);
xnor U22347 (N_22347,N_22112,N_22127);
nor U22348 (N_22348,N_22247,N_22198);
nor U22349 (N_22349,N_22219,N_22047);
or U22350 (N_22350,N_22065,N_22194);
nor U22351 (N_22351,N_22226,N_22002);
nor U22352 (N_22352,N_22013,N_22249);
xor U22353 (N_22353,N_22108,N_22067);
nor U22354 (N_22354,N_22209,N_22037);
nand U22355 (N_22355,N_22237,N_22074);
nor U22356 (N_22356,N_22036,N_22048);
nor U22357 (N_22357,N_22064,N_22235);
nor U22358 (N_22358,N_22169,N_22151);
xor U22359 (N_22359,N_22014,N_22241);
nor U22360 (N_22360,N_22196,N_22230);
xnor U22361 (N_22361,N_22020,N_22166);
or U22362 (N_22362,N_22240,N_22116);
and U22363 (N_22363,N_22246,N_22139);
nand U22364 (N_22364,N_22017,N_22077);
nor U22365 (N_22365,N_22170,N_22069);
or U22366 (N_22366,N_22216,N_22140);
xnor U22367 (N_22367,N_22119,N_22005);
xor U22368 (N_22368,N_22171,N_22195);
xnor U22369 (N_22369,N_22227,N_22189);
nor U22370 (N_22370,N_22004,N_22058);
nor U22371 (N_22371,N_22052,N_22136);
and U22372 (N_22372,N_22051,N_22243);
nand U22373 (N_22373,N_22110,N_22023);
xnor U22374 (N_22374,N_22234,N_22162);
and U22375 (N_22375,N_22125,N_22077);
and U22376 (N_22376,N_22020,N_22192);
or U22377 (N_22377,N_22067,N_22163);
and U22378 (N_22378,N_22081,N_22102);
nor U22379 (N_22379,N_22193,N_22102);
and U22380 (N_22380,N_22212,N_22148);
xnor U22381 (N_22381,N_22077,N_22142);
xnor U22382 (N_22382,N_22136,N_22218);
nand U22383 (N_22383,N_22091,N_22195);
nor U22384 (N_22384,N_22149,N_22137);
and U22385 (N_22385,N_22130,N_22077);
or U22386 (N_22386,N_22200,N_22029);
xor U22387 (N_22387,N_22072,N_22051);
nor U22388 (N_22388,N_22177,N_22033);
and U22389 (N_22389,N_22090,N_22067);
and U22390 (N_22390,N_22011,N_22079);
and U22391 (N_22391,N_22154,N_22105);
nor U22392 (N_22392,N_22047,N_22078);
and U22393 (N_22393,N_22072,N_22112);
or U22394 (N_22394,N_22012,N_22007);
nand U22395 (N_22395,N_22221,N_22199);
xor U22396 (N_22396,N_22091,N_22004);
and U22397 (N_22397,N_22192,N_22082);
nor U22398 (N_22398,N_22024,N_22047);
nor U22399 (N_22399,N_22164,N_22114);
and U22400 (N_22400,N_22072,N_22194);
nand U22401 (N_22401,N_22243,N_22211);
nor U22402 (N_22402,N_22172,N_22033);
nor U22403 (N_22403,N_22206,N_22143);
xor U22404 (N_22404,N_22021,N_22054);
or U22405 (N_22405,N_22003,N_22061);
and U22406 (N_22406,N_22198,N_22170);
or U22407 (N_22407,N_22144,N_22182);
xor U22408 (N_22408,N_22139,N_22239);
nor U22409 (N_22409,N_22138,N_22089);
xnor U22410 (N_22410,N_22211,N_22058);
nor U22411 (N_22411,N_22167,N_22001);
xor U22412 (N_22412,N_22142,N_22084);
nor U22413 (N_22413,N_22083,N_22150);
xor U22414 (N_22414,N_22035,N_22021);
or U22415 (N_22415,N_22085,N_22040);
or U22416 (N_22416,N_22112,N_22126);
nor U22417 (N_22417,N_22176,N_22083);
nand U22418 (N_22418,N_22083,N_22126);
nand U22419 (N_22419,N_22147,N_22183);
and U22420 (N_22420,N_22205,N_22120);
nor U22421 (N_22421,N_22118,N_22086);
or U22422 (N_22422,N_22220,N_22246);
nor U22423 (N_22423,N_22218,N_22102);
and U22424 (N_22424,N_22150,N_22062);
nor U22425 (N_22425,N_22053,N_22062);
xnor U22426 (N_22426,N_22115,N_22032);
nand U22427 (N_22427,N_22053,N_22006);
nor U22428 (N_22428,N_22161,N_22159);
xnor U22429 (N_22429,N_22013,N_22199);
xor U22430 (N_22430,N_22140,N_22161);
nand U22431 (N_22431,N_22049,N_22226);
xnor U22432 (N_22432,N_22138,N_22220);
xnor U22433 (N_22433,N_22050,N_22219);
nor U22434 (N_22434,N_22115,N_22046);
nand U22435 (N_22435,N_22062,N_22112);
or U22436 (N_22436,N_22110,N_22133);
nor U22437 (N_22437,N_22146,N_22162);
or U22438 (N_22438,N_22121,N_22049);
nand U22439 (N_22439,N_22200,N_22001);
nor U22440 (N_22440,N_22167,N_22152);
xnor U22441 (N_22441,N_22046,N_22205);
nand U22442 (N_22442,N_22058,N_22060);
xor U22443 (N_22443,N_22239,N_22181);
or U22444 (N_22444,N_22191,N_22171);
or U22445 (N_22445,N_22110,N_22206);
and U22446 (N_22446,N_22093,N_22090);
xor U22447 (N_22447,N_22060,N_22182);
xnor U22448 (N_22448,N_22003,N_22051);
nor U22449 (N_22449,N_22144,N_22133);
and U22450 (N_22450,N_22162,N_22222);
nor U22451 (N_22451,N_22186,N_22123);
nor U22452 (N_22452,N_22095,N_22249);
xor U22453 (N_22453,N_22154,N_22026);
xor U22454 (N_22454,N_22076,N_22183);
or U22455 (N_22455,N_22076,N_22160);
xor U22456 (N_22456,N_22115,N_22098);
or U22457 (N_22457,N_22054,N_22058);
nand U22458 (N_22458,N_22170,N_22226);
nor U22459 (N_22459,N_22031,N_22108);
and U22460 (N_22460,N_22245,N_22117);
xnor U22461 (N_22461,N_22243,N_22169);
or U22462 (N_22462,N_22215,N_22124);
nand U22463 (N_22463,N_22108,N_22010);
xnor U22464 (N_22464,N_22103,N_22142);
xnor U22465 (N_22465,N_22087,N_22247);
xor U22466 (N_22466,N_22043,N_22065);
xnor U22467 (N_22467,N_22116,N_22073);
or U22468 (N_22468,N_22086,N_22237);
nor U22469 (N_22469,N_22045,N_22083);
xor U22470 (N_22470,N_22080,N_22201);
and U22471 (N_22471,N_22004,N_22040);
or U22472 (N_22472,N_22151,N_22073);
or U22473 (N_22473,N_22103,N_22169);
and U22474 (N_22474,N_22210,N_22110);
or U22475 (N_22475,N_22028,N_22210);
xnor U22476 (N_22476,N_22039,N_22092);
nor U22477 (N_22477,N_22209,N_22146);
and U22478 (N_22478,N_22211,N_22157);
and U22479 (N_22479,N_22081,N_22040);
nand U22480 (N_22480,N_22057,N_22200);
or U22481 (N_22481,N_22060,N_22090);
nand U22482 (N_22482,N_22020,N_22139);
nor U22483 (N_22483,N_22136,N_22190);
nand U22484 (N_22484,N_22071,N_22009);
nor U22485 (N_22485,N_22153,N_22058);
and U22486 (N_22486,N_22191,N_22078);
or U22487 (N_22487,N_22165,N_22052);
or U22488 (N_22488,N_22134,N_22079);
nand U22489 (N_22489,N_22000,N_22033);
nand U22490 (N_22490,N_22079,N_22164);
nand U22491 (N_22491,N_22052,N_22074);
and U22492 (N_22492,N_22101,N_22025);
nand U22493 (N_22493,N_22196,N_22029);
or U22494 (N_22494,N_22095,N_22246);
nor U22495 (N_22495,N_22016,N_22083);
nand U22496 (N_22496,N_22248,N_22072);
xor U22497 (N_22497,N_22245,N_22153);
xor U22498 (N_22498,N_22213,N_22021);
or U22499 (N_22499,N_22136,N_22087);
nand U22500 (N_22500,N_22327,N_22292);
xor U22501 (N_22501,N_22486,N_22331);
nand U22502 (N_22502,N_22280,N_22323);
nor U22503 (N_22503,N_22342,N_22430);
and U22504 (N_22504,N_22329,N_22371);
nand U22505 (N_22505,N_22419,N_22318);
nand U22506 (N_22506,N_22469,N_22309);
nor U22507 (N_22507,N_22254,N_22338);
nor U22508 (N_22508,N_22296,N_22375);
or U22509 (N_22509,N_22363,N_22355);
xor U22510 (N_22510,N_22438,N_22386);
nand U22511 (N_22511,N_22420,N_22380);
or U22512 (N_22512,N_22449,N_22457);
nor U22513 (N_22513,N_22391,N_22266);
nor U22514 (N_22514,N_22427,N_22320);
xor U22515 (N_22515,N_22263,N_22284);
or U22516 (N_22516,N_22300,N_22312);
and U22517 (N_22517,N_22436,N_22479);
or U22518 (N_22518,N_22405,N_22255);
nand U22519 (N_22519,N_22305,N_22361);
nor U22520 (N_22520,N_22389,N_22297);
xor U22521 (N_22521,N_22426,N_22416);
nand U22522 (N_22522,N_22450,N_22448);
and U22523 (N_22523,N_22294,N_22475);
and U22524 (N_22524,N_22392,N_22325);
nand U22525 (N_22525,N_22442,N_22362);
xnor U22526 (N_22526,N_22378,N_22489);
xnor U22527 (N_22527,N_22395,N_22262);
and U22528 (N_22528,N_22374,N_22494);
nor U22529 (N_22529,N_22330,N_22418);
nor U22530 (N_22530,N_22287,N_22252);
and U22531 (N_22531,N_22307,N_22270);
or U22532 (N_22532,N_22335,N_22346);
xnor U22533 (N_22533,N_22465,N_22369);
xor U22534 (N_22534,N_22359,N_22310);
nor U22535 (N_22535,N_22495,N_22417);
nor U22536 (N_22536,N_22488,N_22352);
or U22537 (N_22537,N_22313,N_22453);
xor U22538 (N_22538,N_22261,N_22439);
nand U22539 (N_22539,N_22347,N_22385);
nand U22540 (N_22540,N_22289,N_22492);
or U22541 (N_22541,N_22259,N_22275);
xnor U22542 (N_22542,N_22291,N_22383);
xor U22543 (N_22543,N_22343,N_22372);
nand U22544 (N_22544,N_22433,N_22308);
nor U22545 (N_22545,N_22303,N_22403);
xor U22546 (N_22546,N_22390,N_22274);
nor U22547 (N_22547,N_22299,N_22444);
nor U22548 (N_22548,N_22264,N_22301);
or U22549 (N_22549,N_22487,N_22401);
nand U22550 (N_22550,N_22445,N_22468);
nand U22551 (N_22551,N_22463,N_22435);
nor U22552 (N_22552,N_22476,N_22277);
and U22553 (N_22553,N_22467,N_22348);
xor U22554 (N_22554,N_22499,N_22339);
and U22555 (N_22555,N_22459,N_22269);
or U22556 (N_22556,N_22394,N_22317);
and U22557 (N_22557,N_22422,N_22452);
nor U22558 (N_22558,N_22461,N_22334);
nor U22559 (N_22559,N_22484,N_22421);
or U22560 (N_22560,N_22413,N_22258);
or U22561 (N_22561,N_22491,N_22324);
xor U22562 (N_22562,N_22472,N_22271);
nor U22563 (N_22563,N_22454,N_22431);
or U22564 (N_22564,N_22481,N_22437);
nor U22565 (N_22565,N_22493,N_22290);
nand U22566 (N_22566,N_22283,N_22336);
and U22567 (N_22567,N_22498,N_22408);
and U22568 (N_22568,N_22256,N_22356);
nor U22569 (N_22569,N_22311,N_22281);
xnor U22570 (N_22570,N_22434,N_22279);
or U22571 (N_22571,N_22314,N_22466);
nand U22572 (N_22572,N_22441,N_22407);
and U22573 (N_22573,N_22251,N_22388);
xnor U22574 (N_22574,N_22377,N_22354);
xor U22575 (N_22575,N_22474,N_22477);
nand U22576 (N_22576,N_22397,N_22304);
or U22577 (N_22577,N_22253,N_22332);
nand U22578 (N_22578,N_22285,N_22273);
nor U22579 (N_22579,N_22473,N_22267);
and U22580 (N_22580,N_22447,N_22382);
nand U22581 (N_22581,N_22351,N_22482);
nand U22582 (N_22582,N_22257,N_22370);
xnor U22583 (N_22583,N_22478,N_22268);
nand U22584 (N_22584,N_22393,N_22399);
and U22585 (N_22585,N_22402,N_22298);
and U22586 (N_22586,N_22398,N_22497);
and U22587 (N_22587,N_22432,N_22440);
xnor U22588 (N_22588,N_22470,N_22429);
and U22589 (N_22589,N_22455,N_22373);
xnor U22590 (N_22590,N_22490,N_22344);
xor U22591 (N_22591,N_22295,N_22368);
xor U22592 (N_22592,N_22349,N_22316);
and U22593 (N_22593,N_22387,N_22328);
nand U22594 (N_22594,N_22272,N_22278);
nand U22595 (N_22595,N_22451,N_22341);
nor U22596 (N_22596,N_22333,N_22428);
and U22597 (N_22597,N_22443,N_22282);
nor U22598 (N_22598,N_22384,N_22423);
or U22599 (N_22599,N_22326,N_22412);
or U22600 (N_22600,N_22496,N_22471);
or U22601 (N_22601,N_22315,N_22462);
xor U22602 (N_22602,N_22424,N_22456);
nand U22603 (N_22603,N_22276,N_22250);
or U22604 (N_22604,N_22485,N_22286);
nand U22605 (N_22605,N_22265,N_22350);
xnor U22606 (N_22606,N_22414,N_22410);
nor U22607 (N_22607,N_22381,N_22458);
and U22608 (N_22608,N_22464,N_22404);
nand U22609 (N_22609,N_22340,N_22288);
nor U22610 (N_22610,N_22406,N_22400);
xor U22611 (N_22611,N_22376,N_22260);
or U22612 (N_22612,N_22337,N_22409);
and U22613 (N_22613,N_22358,N_22302);
nor U22614 (N_22614,N_22415,N_22366);
or U22615 (N_22615,N_22367,N_22345);
xor U22616 (N_22616,N_22365,N_22446);
nor U22617 (N_22617,N_22425,N_22360);
or U22618 (N_22618,N_22480,N_22293);
or U22619 (N_22619,N_22460,N_22364);
and U22620 (N_22620,N_22411,N_22322);
xnor U22621 (N_22621,N_22353,N_22319);
nand U22622 (N_22622,N_22396,N_22306);
xor U22623 (N_22623,N_22357,N_22321);
and U22624 (N_22624,N_22379,N_22483);
xnor U22625 (N_22625,N_22270,N_22492);
nand U22626 (N_22626,N_22455,N_22402);
xor U22627 (N_22627,N_22331,N_22307);
or U22628 (N_22628,N_22270,N_22437);
xor U22629 (N_22629,N_22293,N_22452);
nand U22630 (N_22630,N_22410,N_22437);
xor U22631 (N_22631,N_22336,N_22263);
or U22632 (N_22632,N_22353,N_22451);
nor U22633 (N_22633,N_22308,N_22391);
nand U22634 (N_22634,N_22337,N_22467);
and U22635 (N_22635,N_22497,N_22409);
nand U22636 (N_22636,N_22419,N_22250);
xnor U22637 (N_22637,N_22336,N_22359);
or U22638 (N_22638,N_22341,N_22291);
xnor U22639 (N_22639,N_22381,N_22439);
nand U22640 (N_22640,N_22280,N_22460);
or U22641 (N_22641,N_22485,N_22429);
and U22642 (N_22642,N_22464,N_22458);
nand U22643 (N_22643,N_22391,N_22392);
or U22644 (N_22644,N_22270,N_22279);
xnor U22645 (N_22645,N_22386,N_22467);
and U22646 (N_22646,N_22412,N_22463);
xnor U22647 (N_22647,N_22347,N_22466);
or U22648 (N_22648,N_22449,N_22317);
xnor U22649 (N_22649,N_22385,N_22267);
xnor U22650 (N_22650,N_22443,N_22295);
nor U22651 (N_22651,N_22316,N_22313);
nand U22652 (N_22652,N_22267,N_22453);
xnor U22653 (N_22653,N_22267,N_22374);
nand U22654 (N_22654,N_22277,N_22478);
nand U22655 (N_22655,N_22285,N_22325);
or U22656 (N_22656,N_22350,N_22428);
or U22657 (N_22657,N_22369,N_22462);
or U22658 (N_22658,N_22253,N_22475);
nand U22659 (N_22659,N_22251,N_22286);
nor U22660 (N_22660,N_22313,N_22296);
nand U22661 (N_22661,N_22351,N_22359);
and U22662 (N_22662,N_22389,N_22426);
xor U22663 (N_22663,N_22446,N_22459);
and U22664 (N_22664,N_22305,N_22323);
xor U22665 (N_22665,N_22422,N_22474);
or U22666 (N_22666,N_22324,N_22471);
xnor U22667 (N_22667,N_22368,N_22442);
or U22668 (N_22668,N_22296,N_22331);
nor U22669 (N_22669,N_22489,N_22286);
nor U22670 (N_22670,N_22292,N_22316);
nand U22671 (N_22671,N_22393,N_22407);
xnor U22672 (N_22672,N_22401,N_22362);
and U22673 (N_22673,N_22443,N_22396);
or U22674 (N_22674,N_22335,N_22453);
xor U22675 (N_22675,N_22376,N_22369);
nor U22676 (N_22676,N_22342,N_22421);
xnor U22677 (N_22677,N_22348,N_22331);
nand U22678 (N_22678,N_22401,N_22445);
and U22679 (N_22679,N_22489,N_22443);
and U22680 (N_22680,N_22392,N_22253);
nand U22681 (N_22681,N_22369,N_22391);
xor U22682 (N_22682,N_22482,N_22444);
or U22683 (N_22683,N_22351,N_22373);
or U22684 (N_22684,N_22289,N_22470);
and U22685 (N_22685,N_22365,N_22281);
nor U22686 (N_22686,N_22327,N_22458);
and U22687 (N_22687,N_22464,N_22332);
nor U22688 (N_22688,N_22363,N_22375);
nand U22689 (N_22689,N_22472,N_22343);
or U22690 (N_22690,N_22494,N_22496);
nand U22691 (N_22691,N_22450,N_22451);
and U22692 (N_22692,N_22283,N_22482);
nand U22693 (N_22693,N_22289,N_22400);
or U22694 (N_22694,N_22374,N_22263);
nor U22695 (N_22695,N_22383,N_22381);
xnor U22696 (N_22696,N_22480,N_22325);
nor U22697 (N_22697,N_22260,N_22277);
xor U22698 (N_22698,N_22413,N_22309);
nor U22699 (N_22699,N_22488,N_22379);
nand U22700 (N_22700,N_22365,N_22427);
nand U22701 (N_22701,N_22495,N_22265);
xor U22702 (N_22702,N_22477,N_22348);
xor U22703 (N_22703,N_22271,N_22278);
nor U22704 (N_22704,N_22383,N_22445);
nand U22705 (N_22705,N_22281,N_22320);
nand U22706 (N_22706,N_22298,N_22379);
and U22707 (N_22707,N_22251,N_22403);
xnor U22708 (N_22708,N_22296,N_22432);
nor U22709 (N_22709,N_22491,N_22360);
nand U22710 (N_22710,N_22389,N_22484);
xor U22711 (N_22711,N_22417,N_22422);
or U22712 (N_22712,N_22315,N_22454);
nand U22713 (N_22713,N_22459,N_22413);
nor U22714 (N_22714,N_22347,N_22370);
and U22715 (N_22715,N_22392,N_22254);
nand U22716 (N_22716,N_22307,N_22265);
and U22717 (N_22717,N_22289,N_22323);
or U22718 (N_22718,N_22390,N_22361);
and U22719 (N_22719,N_22489,N_22453);
nand U22720 (N_22720,N_22258,N_22344);
nor U22721 (N_22721,N_22415,N_22265);
xor U22722 (N_22722,N_22383,N_22281);
nor U22723 (N_22723,N_22436,N_22390);
or U22724 (N_22724,N_22277,N_22493);
xor U22725 (N_22725,N_22362,N_22393);
or U22726 (N_22726,N_22343,N_22393);
or U22727 (N_22727,N_22365,N_22445);
xnor U22728 (N_22728,N_22290,N_22328);
and U22729 (N_22729,N_22454,N_22316);
nor U22730 (N_22730,N_22276,N_22440);
or U22731 (N_22731,N_22266,N_22375);
xor U22732 (N_22732,N_22294,N_22429);
nand U22733 (N_22733,N_22391,N_22259);
nand U22734 (N_22734,N_22339,N_22413);
xor U22735 (N_22735,N_22463,N_22409);
or U22736 (N_22736,N_22311,N_22258);
or U22737 (N_22737,N_22270,N_22335);
and U22738 (N_22738,N_22463,N_22414);
and U22739 (N_22739,N_22385,N_22406);
nand U22740 (N_22740,N_22496,N_22493);
nor U22741 (N_22741,N_22394,N_22496);
or U22742 (N_22742,N_22291,N_22274);
nand U22743 (N_22743,N_22403,N_22441);
xor U22744 (N_22744,N_22392,N_22333);
and U22745 (N_22745,N_22355,N_22479);
nor U22746 (N_22746,N_22364,N_22314);
nand U22747 (N_22747,N_22364,N_22287);
nand U22748 (N_22748,N_22335,N_22482);
xor U22749 (N_22749,N_22423,N_22339);
or U22750 (N_22750,N_22647,N_22507);
nor U22751 (N_22751,N_22712,N_22695);
nor U22752 (N_22752,N_22685,N_22736);
xnor U22753 (N_22753,N_22508,N_22699);
and U22754 (N_22754,N_22510,N_22636);
nand U22755 (N_22755,N_22526,N_22564);
nor U22756 (N_22756,N_22539,N_22735);
xor U22757 (N_22757,N_22714,N_22541);
nor U22758 (N_22758,N_22590,N_22502);
nor U22759 (N_22759,N_22648,N_22689);
or U22760 (N_22760,N_22536,N_22542);
nand U22761 (N_22761,N_22683,N_22646);
xor U22762 (N_22762,N_22743,N_22623);
nand U22763 (N_22763,N_22557,N_22571);
or U22764 (N_22764,N_22687,N_22522);
nor U22765 (N_22765,N_22578,N_22651);
xnor U22766 (N_22766,N_22744,N_22739);
nor U22767 (N_22767,N_22628,N_22654);
and U22768 (N_22768,N_22707,N_22708);
nor U22769 (N_22769,N_22731,N_22580);
or U22770 (N_22770,N_22677,N_22527);
or U22771 (N_22771,N_22514,N_22547);
xnor U22772 (N_22772,N_22504,N_22546);
and U22773 (N_22773,N_22729,N_22706);
nor U22774 (N_22774,N_22548,N_22663);
nor U22775 (N_22775,N_22671,N_22723);
nand U22776 (N_22776,N_22741,N_22724);
nand U22777 (N_22777,N_22650,N_22516);
nand U22778 (N_22778,N_22703,N_22675);
xnor U22779 (N_22779,N_22748,N_22612);
or U22780 (N_22780,N_22622,N_22566);
xnor U22781 (N_22781,N_22607,N_22725);
or U22782 (N_22782,N_22589,N_22558);
and U22783 (N_22783,N_22596,N_22694);
xor U22784 (N_22784,N_22637,N_22627);
and U22785 (N_22785,N_22704,N_22626);
or U22786 (N_22786,N_22710,N_22652);
nand U22787 (N_22787,N_22599,N_22574);
or U22788 (N_22788,N_22512,N_22718);
and U22789 (N_22789,N_22586,N_22561);
xnor U22790 (N_22790,N_22594,N_22719);
or U22791 (N_22791,N_22713,N_22524);
xor U22792 (N_22792,N_22641,N_22538);
nor U22793 (N_22793,N_22584,N_22597);
nand U22794 (N_22794,N_22501,N_22696);
and U22795 (N_22795,N_22598,N_22544);
or U22796 (N_22796,N_22575,N_22552);
or U22797 (N_22797,N_22616,N_22554);
or U22798 (N_22798,N_22738,N_22611);
xnor U22799 (N_22799,N_22519,N_22635);
or U22800 (N_22800,N_22667,N_22701);
nor U22801 (N_22801,N_22656,N_22533);
xnor U22802 (N_22802,N_22692,N_22661);
and U22803 (N_22803,N_22669,N_22601);
xnor U22804 (N_22804,N_22520,N_22509);
nand U22805 (N_22805,N_22543,N_22732);
or U22806 (N_22806,N_22749,N_22591);
nor U22807 (N_22807,N_22624,N_22528);
and U22808 (N_22808,N_22585,N_22549);
nor U22809 (N_22809,N_22716,N_22730);
or U22810 (N_22810,N_22700,N_22556);
nand U22811 (N_22811,N_22605,N_22600);
xnor U22812 (N_22812,N_22746,N_22702);
xor U22813 (N_22813,N_22532,N_22506);
and U22814 (N_22814,N_22657,N_22518);
nand U22815 (N_22815,N_22614,N_22666);
and U22816 (N_22816,N_22634,N_22503);
nor U22817 (N_22817,N_22745,N_22662);
nor U22818 (N_22818,N_22540,N_22631);
and U22819 (N_22819,N_22682,N_22582);
xor U22820 (N_22820,N_22620,N_22587);
xor U22821 (N_22821,N_22545,N_22728);
xnor U22822 (N_22822,N_22581,N_22705);
xor U22823 (N_22823,N_22595,N_22569);
or U22824 (N_22824,N_22638,N_22680);
nand U22825 (N_22825,N_22643,N_22619);
xnor U22826 (N_22826,N_22555,N_22727);
or U22827 (N_22827,N_22747,N_22523);
nand U22828 (N_22828,N_22511,N_22668);
and U22829 (N_22829,N_22686,N_22500);
and U22830 (N_22830,N_22665,N_22640);
and U22831 (N_22831,N_22726,N_22579);
nor U22832 (N_22832,N_22563,N_22525);
nand U22833 (N_22833,N_22577,N_22602);
xnor U22834 (N_22834,N_22551,N_22664);
and U22835 (N_22835,N_22603,N_22537);
and U22836 (N_22836,N_22698,N_22606);
or U22837 (N_22837,N_22573,N_22717);
xor U22838 (N_22838,N_22676,N_22608);
nor U22839 (N_22839,N_22560,N_22632);
and U22840 (N_22840,N_22562,N_22733);
nor U22841 (N_22841,N_22588,N_22642);
and U22842 (N_22842,N_22618,N_22658);
nand U22843 (N_22843,N_22550,N_22672);
nand U22844 (N_22844,N_22720,N_22565);
or U22845 (N_22845,N_22655,N_22576);
or U22846 (N_22846,N_22709,N_22678);
nor U22847 (N_22847,N_22583,N_22531);
xnor U22848 (N_22848,N_22572,N_22553);
xor U22849 (N_22849,N_22670,N_22567);
and U22850 (N_22850,N_22535,N_22721);
nor U22851 (N_22851,N_22534,N_22633);
and U22852 (N_22852,N_22688,N_22734);
and U22853 (N_22853,N_22715,N_22711);
or U22854 (N_22854,N_22593,N_22659);
and U22855 (N_22855,N_22610,N_22570);
xnor U22856 (N_22856,N_22697,N_22517);
or U22857 (N_22857,N_22604,N_22737);
xnor U22858 (N_22858,N_22621,N_22568);
and U22859 (N_22859,N_22530,N_22521);
and U22860 (N_22860,N_22691,N_22592);
nor U22861 (N_22861,N_22684,N_22681);
nor U22862 (N_22862,N_22660,N_22690);
or U22863 (N_22863,N_22679,N_22505);
or U22864 (N_22864,N_22630,N_22515);
nand U22865 (N_22865,N_22629,N_22740);
or U22866 (N_22866,N_22529,N_22613);
nand U22867 (N_22867,N_22615,N_22649);
and U22868 (N_22868,N_22625,N_22673);
or U22869 (N_22869,N_22639,N_22644);
or U22870 (N_22870,N_22693,N_22559);
and U22871 (N_22871,N_22674,N_22609);
or U22872 (N_22872,N_22722,N_22742);
nand U22873 (N_22873,N_22513,N_22653);
and U22874 (N_22874,N_22617,N_22645);
nor U22875 (N_22875,N_22558,N_22557);
nand U22876 (N_22876,N_22578,N_22733);
or U22877 (N_22877,N_22660,N_22686);
nor U22878 (N_22878,N_22555,N_22521);
or U22879 (N_22879,N_22564,N_22599);
and U22880 (N_22880,N_22648,N_22577);
and U22881 (N_22881,N_22585,N_22623);
or U22882 (N_22882,N_22609,N_22720);
or U22883 (N_22883,N_22634,N_22605);
xnor U22884 (N_22884,N_22613,N_22693);
nor U22885 (N_22885,N_22726,N_22669);
or U22886 (N_22886,N_22717,N_22617);
xor U22887 (N_22887,N_22730,N_22661);
nand U22888 (N_22888,N_22606,N_22509);
nor U22889 (N_22889,N_22725,N_22545);
xor U22890 (N_22890,N_22575,N_22502);
nand U22891 (N_22891,N_22585,N_22560);
nand U22892 (N_22892,N_22638,N_22729);
xor U22893 (N_22893,N_22652,N_22596);
xnor U22894 (N_22894,N_22549,N_22555);
nor U22895 (N_22895,N_22690,N_22685);
nor U22896 (N_22896,N_22553,N_22703);
or U22897 (N_22897,N_22523,N_22535);
or U22898 (N_22898,N_22540,N_22502);
or U22899 (N_22899,N_22537,N_22650);
nand U22900 (N_22900,N_22602,N_22576);
xnor U22901 (N_22901,N_22669,N_22629);
nor U22902 (N_22902,N_22548,N_22734);
xnor U22903 (N_22903,N_22743,N_22600);
and U22904 (N_22904,N_22702,N_22542);
xor U22905 (N_22905,N_22536,N_22730);
or U22906 (N_22906,N_22557,N_22740);
and U22907 (N_22907,N_22742,N_22636);
or U22908 (N_22908,N_22648,N_22711);
xor U22909 (N_22909,N_22554,N_22567);
xnor U22910 (N_22910,N_22716,N_22611);
and U22911 (N_22911,N_22548,N_22673);
nor U22912 (N_22912,N_22638,N_22616);
and U22913 (N_22913,N_22548,N_22633);
and U22914 (N_22914,N_22506,N_22592);
or U22915 (N_22915,N_22719,N_22727);
and U22916 (N_22916,N_22575,N_22613);
or U22917 (N_22917,N_22602,N_22533);
and U22918 (N_22918,N_22537,N_22647);
and U22919 (N_22919,N_22735,N_22690);
xnor U22920 (N_22920,N_22536,N_22532);
nand U22921 (N_22921,N_22504,N_22535);
nand U22922 (N_22922,N_22681,N_22650);
nand U22923 (N_22923,N_22535,N_22690);
nor U22924 (N_22924,N_22613,N_22609);
xor U22925 (N_22925,N_22559,N_22708);
nor U22926 (N_22926,N_22583,N_22742);
nor U22927 (N_22927,N_22703,N_22546);
and U22928 (N_22928,N_22554,N_22687);
and U22929 (N_22929,N_22602,N_22643);
nand U22930 (N_22930,N_22636,N_22605);
nor U22931 (N_22931,N_22574,N_22582);
or U22932 (N_22932,N_22662,N_22715);
or U22933 (N_22933,N_22740,N_22516);
nor U22934 (N_22934,N_22738,N_22684);
and U22935 (N_22935,N_22625,N_22569);
xor U22936 (N_22936,N_22724,N_22674);
nand U22937 (N_22937,N_22581,N_22725);
xor U22938 (N_22938,N_22719,N_22691);
or U22939 (N_22939,N_22578,N_22530);
or U22940 (N_22940,N_22639,N_22706);
or U22941 (N_22941,N_22562,N_22686);
or U22942 (N_22942,N_22684,N_22578);
nor U22943 (N_22943,N_22622,N_22636);
nor U22944 (N_22944,N_22623,N_22544);
nor U22945 (N_22945,N_22725,N_22518);
nor U22946 (N_22946,N_22550,N_22515);
nor U22947 (N_22947,N_22570,N_22528);
nor U22948 (N_22948,N_22593,N_22648);
and U22949 (N_22949,N_22604,N_22721);
and U22950 (N_22950,N_22524,N_22632);
nand U22951 (N_22951,N_22577,N_22671);
or U22952 (N_22952,N_22719,N_22577);
or U22953 (N_22953,N_22666,N_22649);
nor U22954 (N_22954,N_22700,N_22742);
nand U22955 (N_22955,N_22681,N_22718);
nor U22956 (N_22956,N_22567,N_22585);
xor U22957 (N_22957,N_22602,N_22556);
xnor U22958 (N_22958,N_22705,N_22508);
or U22959 (N_22959,N_22625,N_22616);
and U22960 (N_22960,N_22513,N_22684);
xor U22961 (N_22961,N_22626,N_22612);
nor U22962 (N_22962,N_22604,N_22689);
nor U22963 (N_22963,N_22719,N_22718);
or U22964 (N_22964,N_22531,N_22521);
nor U22965 (N_22965,N_22534,N_22697);
and U22966 (N_22966,N_22672,N_22671);
xor U22967 (N_22967,N_22532,N_22745);
xor U22968 (N_22968,N_22699,N_22536);
xor U22969 (N_22969,N_22735,N_22588);
or U22970 (N_22970,N_22528,N_22640);
nand U22971 (N_22971,N_22704,N_22617);
or U22972 (N_22972,N_22729,N_22687);
nand U22973 (N_22973,N_22707,N_22683);
or U22974 (N_22974,N_22509,N_22540);
and U22975 (N_22975,N_22708,N_22744);
nand U22976 (N_22976,N_22721,N_22638);
xor U22977 (N_22977,N_22546,N_22631);
and U22978 (N_22978,N_22576,N_22732);
xnor U22979 (N_22979,N_22725,N_22601);
or U22980 (N_22980,N_22670,N_22628);
nor U22981 (N_22981,N_22741,N_22701);
or U22982 (N_22982,N_22745,N_22623);
nor U22983 (N_22983,N_22590,N_22535);
nor U22984 (N_22984,N_22692,N_22577);
nand U22985 (N_22985,N_22558,N_22565);
nand U22986 (N_22986,N_22576,N_22605);
or U22987 (N_22987,N_22574,N_22596);
and U22988 (N_22988,N_22719,N_22536);
nand U22989 (N_22989,N_22606,N_22637);
nor U22990 (N_22990,N_22512,N_22687);
and U22991 (N_22991,N_22562,N_22583);
xnor U22992 (N_22992,N_22517,N_22552);
or U22993 (N_22993,N_22741,N_22653);
and U22994 (N_22994,N_22513,N_22739);
and U22995 (N_22995,N_22749,N_22504);
nor U22996 (N_22996,N_22727,N_22583);
xnor U22997 (N_22997,N_22682,N_22729);
nand U22998 (N_22998,N_22612,N_22515);
xor U22999 (N_22999,N_22725,N_22719);
nand U23000 (N_23000,N_22857,N_22981);
nand U23001 (N_23001,N_22910,N_22845);
nor U23002 (N_23002,N_22827,N_22868);
nand U23003 (N_23003,N_22894,N_22799);
or U23004 (N_23004,N_22779,N_22817);
and U23005 (N_23005,N_22835,N_22923);
nand U23006 (N_23006,N_22931,N_22965);
xnor U23007 (N_23007,N_22980,N_22874);
xnor U23008 (N_23008,N_22829,N_22977);
and U23009 (N_23009,N_22888,N_22998);
xnor U23010 (N_23010,N_22880,N_22922);
nand U23011 (N_23011,N_22819,N_22760);
and U23012 (N_23012,N_22918,N_22841);
and U23013 (N_23013,N_22935,N_22772);
and U23014 (N_23014,N_22899,N_22833);
and U23015 (N_23015,N_22852,N_22952);
nor U23016 (N_23016,N_22974,N_22797);
or U23017 (N_23017,N_22863,N_22756);
or U23018 (N_23018,N_22893,N_22768);
nor U23019 (N_23019,N_22896,N_22940);
and U23020 (N_23020,N_22867,N_22966);
xor U23021 (N_23021,N_22808,N_22987);
nand U23022 (N_23022,N_22961,N_22785);
xnor U23023 (N_23023,N_22956,N_22959);
nand U23024 (N_23024,N_22790,N_22786);
xnor U23025 (N_23025,N_22881,N_22984);
nand U23026 (N_23026,N_22944,N_22828);
and U23027 (N_23027,N_22955,N_22812);
xnor U23028 (N_23028,N_22842,N_22866);
and U23029 (N_23029,N_22905,N_22869);
nor U23030 (N_23030,N_22810,N_22891);
xor U23031 (N_23031,N_22846,N_22793);
or U23032 (N_23032,N_22764,N_22825);
nor U23033 (N_23033,N_22858,N_22982);
nand U23034 (N_23034,N_22872,N_22826);
or U23035 (N_23035,N_22989,N_22757);
and U23036 (N_23036,N_22775,N_22850);
and U23037 (N_23037,N_22912,N_22851);
and U23038 (N_23038,N_22898,N_22946);
and U23039 (N_23039,N_22798,N_22876);
nor U23040 (N_23040,N_22773,N_22892);
or U23041 (N_23041,N_22902,N_22770);
nor U23042 (N_23042,N_22767,N_22886);
or U23043 (N_23043,N_22934,N_22838);
nand U23044 (N_23044,N_22873,N_22854);
xnor U23045 (N_23045,N_22967,N_22803);
nand U23046 (N_23046,N_22992,N_22921);
nor U23047 (N_23047,N_22818,N_22945);
or U23048 (N_23048,N_22849,N_22929);
xor U23049 (N_23049,N_22788,N_22871);
nor U23050 (N_23050,N_22901,N_22976);
and U23051 (N_23051,N_22914,N_22909);
nand U23052 (N_23052,N_22837,N_22795);
nand U23053 (N_23053,N_22957,N_22784);
and U23054 (N_23054,N_22993,N_22811);
nand U23055 (N_23055,N_22939,N_22942);
xor U23056 (N_23056,N_22995,N_22947);
or U23057 (N_23057,N_22840,N_22755);
and U23058 (N_23058,N_22792,N_22776);
nor U23059 (N_23059,N_22823,N_22853);
nor U23060 (N_23060,N_22975,N_22904);
nor U23061 (N_23061,N_22794,N_22862);
nor U23062 (N_23062,N_22927,N_22883);
or U23063 (N_23063,N_22752,N_22978);
nand U23064 (N_23064,N_22807,N_22937);
or U23065 (N_23065,N_22796,N_22990);
and U23066 (N_23066,N_22844,N_22916);
nor U23067 (N_23067,N_22915,N_22753);
and U23068 (N_23068,N_22890,N_22814);
or U23069 (N_23069,N_22781,N_22815);
nor U23070 (N_23070,N_22761,N_22831);
nor U23071 (N_23071,N_22991,N_22865);
xor U23072 (N_23072,N_22970,N_22908);
or U23073 (N_23073,N_22996,N_22791);
and U23074 (N_23074,N_22839,N_22830);
nand U23075 (N_23075,N_22800,N_22948);
xnor U23076 (N_23076,N_22924,N_22994);
nor U23077 (N_23077,N_22895,N_22843);
nand U23078 (N_23078,N_22877,N_22780);
and U23079 (N_23079,N_22906,N_22802);
nand U23080 (N_23080,N_22885,N_22986);
and U23081 (N_23081,N_22787,N_22925);
nand U23082 (N_23082,N_22953,N_22928);
and U23083 (N_23083,N_22856,N_22907);
nor U23084 (N_23084,N_22884,N_22809);
or U23085 (N_23085,N_22765,N_22801);
nor U23086 (N_23086,N_22848,N_22778);
nor U23087 (N_23087,N_22950,N_22962);
xnor U23088 (N_23088,N_22887,N_22821);
nor U23089 (N_23089,N_22930,N_22762);
nand U23090 (N_23090,N_22932,N_22971);
xor U23091 (N_23091,N_22882,N_22820);
xnor U23092 (N_23092,N_22861,N_22926);
or U23093 (N_23093,N_22750,N_22911);
and U23094 (N_23094,N_22783,N_22759);
and U23095 (N_23095,N_22999,N_22960);
nand U23096 (N_23096,N_22954,N_22903);
nand U23097 (N_23097,N_22813,N_22972);
and U23098 (N_23098,N_22943,N_22963);
and U23099 (N_23099,N_22754,N_22836);
or U23100 (N_23100,N_22941,N_22864);
nand U23101 (N_23101,N_22988,N_22964);
or U23102 (N_23102,N_22920,N_22889);
or U23103 (N_23103,N_22860,N_22859);
nand U23104 (N_23104,N_22805,N_22938);
or U23105 (N_23105,N_22968,N_22997);
nand U23106 (N_23106,N_22913,N_22816);
nor U23107 (N_23107,N_22951,N_22777);
xor U23108 (N_23108,N_22834,N_22985);
xnor U23109 (N_23109,N_22804,N_22822);
and U23110 (N_23110,N_22758,N_22969);
xor U23111 (N_23111,N_22832,N_22771);
xor U23112 (N_23112,N_22789,N_22919);
and U23113 (N_23113,N_22870,N_22983);
xor U23114 (N_23114,N_22751,N_22900);
nor U23115 (N_23115,N_22763,N_22958);
nor U23116 (N_23116,N_22782,N_22769);
and U23117 (N_23117,N_22847,N_22824);
and U23118 (N_23118,N_22774,N_22875);
nor U23119 (N_23119,N_22973,N_22766);
nor U23120 (N_23120,N_22933,N_22936);
nand U23121 (N_23121,N_22879,N_22979);
xnor U23122 (N_23122,N_22949,N_22878);
nand U23123 (N_23123,N_22806,N_22897);
or U23124 (N_23124,N_22855,N_22917);
xor U23125 (N_23125,N_22895,N_22975);
and U23126 (N_23126,N_22819,N_22774);
and U23127 (N_23127,N_22969,N_22899);
and U23128 (N_23128,N_22935,N_22825);
xor U23129 (N_23129,N_22996,N_22955);
xor U23130 (N_23130,N_22850,N_22970);
xor U23131 (N_23131,N_22922,N_22933);
and U23132 (N_23132,N_22856,N_22923);
and U23133 (N_23133,N_22764,N_22879);
and U23134 (N_23134,N_22889,N_22891);
xnor U23135 (N_23135,N_22759,N_22861);
or U23136 (N_23136,N_22923,N_22846);
nor U23137 (N_23137,N_22835,N_22891);
or U23138 (N_23138,N_22784,N_22811);
nor U23139 (N_23139,N_22956,N_22802);
or U23140 (N_23140,N_22993,N_22836);
or U23141 (N_23141,N_22837,N_22811);
and U23142 (N_23142,N_22920,N_22827);
nand U23143 (N_23143,N_22935,N_22858);
or U23144 (N_23144,N_22990,N_22913);
and U23145 (N_23145,N_22892,N_22937);
and U23146 (N_23146,N_22821,N_22990);
nor U23147 (N_23147,N_22868,N_22885);
and U23148 (N_23148,N_22848,N_22893);
xor U23149 (N_23149,N_22910,N_22755);
nor U23150 (N_23150,N_22951,N_22926);
and U23151 (N_23151,N_22934,N_22979);
nand U23152 (N_23152,N_22861,N_22862);
xor U23153 (N_23153,N_22939,N_22843);
and U23154 (N_23154,N_22789,N_22892);
or U23155 (N_23155,N_22989,N_22971);
xor U23156 (N_23156,N_22773,N_22966);
xnor U23157 (N_23157,N_22877,N_22764);
and U23158 (N_23158,N_22811,N_22761);
nand U23159 (N_23159,N_22753,N_22958);
and U23160 (N_23160,N_22967,N_22902);
nor U23161 (N_23161,N_22804,N_22865);
and U23162 (N_23162,N_22904,N_22850);
and U23163 (N_23163,N_22779,N_22953);
nand U23164 (N_23164,N_22813,N_22791);
nor U23165 (N_23165,N_22768,N_22930);
nor U23166 (N_23166,N_22788,N_22957);
and U23167 (N_23167,N_22808,N_22819);
and U23168 (N_23168,N_22939,N_22930);
nor U23169 (N_23169,N_22957,N_22914);
or U23170 (N_23170,N_22770,N_22766);
xnor U23171 (N_23171,N_22974,N_22993);
nor U23172 (N_23172,N_22847,N_22803);
or U23173 (N_23173,N_22950,N_22816);
or U23174 (N_23174,N_22845,N_22900);
or U23175 (N_23175,N_22948,N_22885);
nor U23176 (N_23176,N_22861,N_22990);
xnor U23177 (N_23177,N_22932,N_22774);
and U23178 (N_23178,N_22835,N_22907);
xnor U23179 (N_23179,N_22797,N_22898);
and U23180 (N_23180,N_22803,N_22931);
or U23181 (N_23181,N_22901,N_22767);
nand U23182 (N_23182,N_22799,N_22814);
nor U23183 (N_23183,N_22894,N_22834);
or U23184 (N_23184,N_22780,N_22762);
or U23185 (N_23185,N_22998,N_22986);
nand U23186 (N_23186,N_22752,N_22804);
or U23187 (N_23187,N_22817,N_22801);
and U23188 (N_23188,N_22806,N_22778);
nand U23189 (N_23189,N_22946,N_22844);
nor U23190 (N_23190,N_22827,N_22922);
nand U23191 (N_23191,N_22970,N_22861);
xnor U23192 (N_23192,N_22903,N_22816);
nand U23193 (N_23193,N_22836,N_22892);
nor U23194 (N_23194,N_22935,N_22784);
nand U23195 (N_23195,N_22926,N_22833);
or U23196 (N_23196,N_22962,N_22795);
nand U23197 (N_23197,N_22904,N_22996);
or U23198 (N_23198,N_22944,N_22910);
nand U23199 (N_23199,N_22820,N_22847);
nand U23200 (N_23200,N_22756,N_22930);
xor U23201 (N_23201,N_22942,N_22840);
and U23202 (N_23202,N_22962,N_22948);
and U23203 (N_23203,N_22873,N_22988);
or U23204 (N_23204,N_22970,N_22886);
and U23205 (N_23205,N_22906,N_22929);
nand U23206 (N_23206,N_22909,N_22913);
and U23207 (N_23207,N_22959,N_22952);
nand U23208 (N_23208,N_22920,N_22938);
nor U23209 (N_23209,N_22894,N_22853);
nand U23210 (N_23210,N_22811,N_22907);
and U23211 (N_23211,N_22925,N_22786);
and U23212 (N_23212,N_22896,N_22880);
and U23213 (N_23213,N_22921,N_22806);
nand U23214 (N_23214,N_22883,N_22778);
and U23215 (N_23215,N_22974,N_22763);
nor U23216 (N_23216,N_22880,N_22838);
nor U23217 (N_23217,N_22828,N_22756);
nand U23218 (N_23218,N_22990,N_22846);
nand U23219 (N_23219,N_22772,N_22756);
nor U23220 (N_23220,N_22914,N_22803);
nand U23221 (N_23221,N_22965,N_22809);
nor U23222 (N_23222,N_22909,N_22776);
nor U23223 (N_23223,N_22943,N_22864);
xor U23224 (N_23224,N_22815,N_22795);
and U23225 (N_23225,N_22795,N_22980);
and U23226 (N_23226,N_22770,N_22881);
nand U23227 (N_23227,N_22974,N_22753);
nand U23228 (N_23228,N_22965,N_22941);
or U23229 (N_23229,N_22861,N_22873);
nand U23230 (N_23230,N_22909,N_22781);
xor U23231 (N_23231,N_22946,N_22835);
nor U23232 (N_23232,N_22893,N_22978);
xnor U23233 (N_23233,N_22762,N_22878);
xor U23234 (N_23234,N_22955,N_22882);
nand U23235 (N_23235,N_22862,N_22970);
and U23236 (N_23236,N_22892,N_22998);
and U23237 (N_23237,N_22903,N_22797);
nand U23238 (N_23238,N_22807,N_22997);
or U23239 (N_23239,N_22959,N_22829);
nand U23240 (N_23240,N_22929,N_22770);
nor U23241 (N_23241,N_22966,N_22762);
nor U23242 (N_23242,N_22943,N_22892);
nor U23243 (N_23243,N_22961,N_22945);
and U23244 (N_23244,N_22916,N_22756);
xor U23245 (N_23245,N_22826,N_22991);
nor U23246 (N_23246,N_22783,N_22996);
nor U23247 (N_23247,N_22827,N_22986);
nor U23248 (N_23248,N_22783,N_22754);
nand U23249 (N_23249,N_22783,N_22806);
nand U23250 (N_23250,N_23021,N_23183);
or U23251 (N_23251,N_23200,N_23005);
xnor U23252 (N_23252,N_23020,N_23161);
and U23253 (N_23253,N_23007,N_23099);
nand U23254 (N_23254,N_23228,N_23106);
or U23255 (N_23255,N_23185,N_23057);
nor U23256 (N_23256,N_23157,N_23216);
and U23257 (N_23257,N_23165,N_23048);
and U23258 (N_23258,N_23065,N_23122);
and U23259 (N_23259,N_23178,N_23140);
or U23260 (N_23260,N_23231,N_23088);
nand U23261 (N_23261,N_23008,N_23215);
nor U23262 (N_23262,N_23126,N_23025);
or U23263 (N_23263,N_23062,N_23100);
and U23264 (N_23264,N_23222,N_23085);
nand U23265 (N_23265,N_23040,N_23138);
and U23266 (N_23266,N_23019,N_23198);
xnor U23267 (N_23267,N_23219,N_23091);
xor U23268 (N_23268,N_23024,N_23217);
nor U23269 (N_23269,N_23131,N_23236);
or U23270 (N_23270,N_23006,N_23243);
nor U23271 (N_23271,N_23066,N_23064);
nor U23272 (N_23272,N_23061,N_23029);
nand U23273 (N_23273,N_23030,N_23001);
nor U23274 (N_23274,N_23150,N_23156);
nand U23275 (N_23275,N_23022,N_23071);
nand U23276 (N_23276,N_23074,N_23238);
nor U23277 (N_23277,N_23118,N_23063);
or U23278 (N_23278,N_23086,N_23214);
and U23279 (N_23279,N_23162,N_23110);
nand U23280 (N_23280,N_23059,N_23234);
and U23281 (N_23281,N_23158,N_23143);
nor U23282 (N_23282,N_23245,N_23130);
and U23283 (N_23283,N_23211,N_23123);
and U23284 (N_23284,N_23016,N_23056);
or U23285 (N_23285,N_23155,N_23010);
nor U23286 (N_23286,N_23046,N_23232);
or U23287 (N_23287,N_23032,N_23179);
nor U23288 (N_23288,N_23166,N_23244);
nand U23289 (N_23289,N_23141,N_23055);
xor U23290 (N_23290,N_23120,N_23213);
nand U23291 (N_23291,N_23180,N_23047);
nor U23292 (N_23292,N_23146,N_23090);
or U23293 (N_23293,N_23013,N_23102);
or U23294 (N_23294,N_23172,N_23104);
xor U23295 (N_23295,N_23109,N_23044);
xnor U23296 (N_23296,N_23240,N_23014);
and U23297 (N_23297,N_23193,N_23164);
nor U23298 (N_23298,N_23176,N_23073);
nor U23299 (N_23299,N_23194,N_23116);
xnor U23300 (N_23300,N_23145,N_23149);
nor U23301 (N_23301,N_23197,N_23127);
nor U23302 (N_23302,N_23224,N_23171);
or U23303 (N_23303,N_23049,N_23015);
nand U23304 (N_23304,N_23092,N_23079);
nand U23305 (N_23305,N_23169,N_23002);
nor U23306 (N_23306,N_23201,N_23163);
or U23307 (N_23307,N_23195,N_23009);
and U23308 (N_23308,N_23137,N_23208);
nand U23309 (N_23309,N_23050,N_23142);
nor U23310 (N_23310,N_23026,N_23045);
nand U23311 (N_23311,N_23115,N_23038);
and U23312 (N_23312,N_23136,N_23139);
nand U23313 (N_23313,N_23230,N_23188);
nor U23314 (N_23314,N_23018,N_23000);
nand U23315 (N_23315,N_23089,N_23082);
nor U23316 (N_23316,N_23237,N_23075);
and U23317 (N_23317,N_23170,N_23233);
nor U23318 (N_23318,N_23067,N_23028);
or U23319 (N_23319,N_23248,N_23107);
xnor U23320 (N_23320,N_23031,N_23069);
xor U23321 (N_23321,N_23241,N_23043);
nor U23322 (N_23322,N_23209,N_23175);
nor U23323 (N_23323,N_23182,N_23152);
nor U23324 (N_23324,N_23084,N_23058);
xor U23325 (N_23325,N_23148,N_23221);
or U23326 (N_23326,N_23192,N_23205);
nand U23327 (N_23327,N_23135,N_23226);
or U23328 (N_23328,N_23220,N_23206);
nor U23329 (N_23329,N_23174,N_23167);
or U23330 (N_23330,N_23225,N_23027);
and U23331 (N_23331,N_23042,N_23052);
or U23332 (N_23332,N_23097,N_23189);
or U23333 (N_23333,N_23103,N_23117);
or U23334 (N_23334,N_23060,N_23054);
xnor U23335 (N_23335,N_23078,N_23105);
nor U23336 (N_23336,N_23087,N_23053);
or U23337 (N_23337,N_23023,N_23114);
nand U23338 (N_23338,N_23111,N_23246);
nor U23339 (N_23339,N_23003,N_23101);
or U23340 (N_23340,N_23108,N_23177);
xnor U23341 (N_23341,N_23129,N_23168);
xor U23342 (N_23342,N_23153,N_23017);
nand U23343 (N_23343,N_23147,N_23098);
and U23344 (N_23344,N_23113,N_23077);
nor U23345 (N_23345,N_23159,N_23112);
nand U23346 (N_23346,N_23184,N_23199);
or U23347 (N_23347,N_23207,N_23235);
and U23348 (N_23348,N_23190,N_23051);
and U23349 (N_23349,N_23096,N_23154);
nor U23350 (N_23350,N_23218,N_23173);
nor U23351 (N_23351,N_23076,N_23041);
xnor U23352 (N_23352,N_23144,N_23212);
nor U23353 (N_23353,N_23033,N_23204);
or U23354 (N_23354,N_23004,N_23132);
and U23355 (N_23355,N_23068,N_23247);
nand U23356 (N_23356,N_23011,N_23070);
nand U23357 (N_23357,N_23012,N_23034);
xnor U23358 (N_23358,N_23202,N_23036);
and U23359 (N_23359,N_23242,N_23191);
nor U23360 (N_23360,N_23124,N_23083);
xor U23361 (N_23361,N_23121,N_23187);
or U23362 (N_23362,N_23196,N_23072);
and U23363 (N_23363,N_23125,N_23203);
or U23364 (N_23364,N_23080,N_23095);
xnor U23365 (N_23365,N_23128,N_23239);
and U23366 (N_23366,N_23181,N_23134);
nand U23367 (N_23367,N_23160,N_23227);
nand U23368 (N_23368,N_23229,N_23081);
nand U23369 (N_23369,N_23186,N_23119);
or U23370 (N_23370,N_23210,N_23151);
or U23371 (N_23371,N_23094,N_23037);
nor U23372 (N_23372,N_23039,N_23093);
or U23373 (N_23373,N_23035,N_23223);
nand U23374 (N_23374,N_23133,N_23249);
and U23375 (N_23375,N_23193,N_23212);
nor U23376 (N_23376,N_23040,N_23151);
xnor U23377 (N_23377,N_23052,N_23201);
nor U23378 (N_23378,N_23020,N_23241);
nand U23379 (N_23379,N_23102,N_23232);
nand U23380 (N_23380,N_23189,N_23192);
xnor U23381 (N_23381,N_23099,N_23134);
or U23382 (N_23382,N_23015,N_23162);
or U23383 (N_23383,N_23238,N_23225);
or U23384 (N_23384,N_23083,N_23187);
nand U23385 (N_23385,N_23241,N_23110);
nor U23386 (N_23386,N_23087,N_23031);
xor U23387 (N_23387,N_23164,N_23206);
nand U23388 (N_23388,N_23200,N_23031);
nand U23389 (N_23389,N_23212,N_23072);
nor U23390 (N_23390,N_23064,N_23210);
xor U23391 (N_23391,N_23084,N_23033);
nand U23392 (N_23392,N_23028,N_23074);
or U23393 (N_23393,N_23216,N_23150);
xnor U23394 (N_23394,N_23056,N_23130);
nand U23395 (N_23395,N_23061,N_23083);
nor U23396 (N_23396,N_23047,N_23196);
nor U23397 (N_23397,N_23140,N_23021);
or U23398 (N_23398,N_23242,N_23202);
nor U23399 (N_23399,N_23080,N_23190);
xor U23400 (N_23400,N_23136,N_23011);
nor U23401 (N_23401,N_23057,N_23084);
and U23402 (N_23402,N_23116,N_23068);
xor U23403 (N_23403,N_23129,N_23011);
and U23404 (N_23404,N_23185,N_23092);
or U23405 (N_23405,N_23068,N_23165);
xor U23406 (N_23406,N_23051,N_23035);
nor U23407 (N_23407,N_23004,N_23114);
or U23408 (N_23408,N_23150,N_23242);
and U23409 (N_23409,N_23211,N_23000);
and U23410 (N_23410,N_23223,N_23008);
nor U23411 (N_23411,N_23005,N_23087);
or U23412 (N_23412,N_23114,N_23210);
nor U23413 (N_23413,N_23048,N_23009);
or U23414 (N_23414,N_23046,N_23078);
xor U23415 (N_23415,N_23099,N_23123);
or U23416 (N_23416,N_23077,N_23136);
nand U23417 (N_23417,N_23161,N_23195);
xnor U23418 (N_23418,N_23120,N_23128);
nor U23419 (N_23419,N_23127,N_23200);
or U23420 (N_23420,N_23140,N_23036);
and U23421 (N_23421,N_23212,N_23017);
nor U23422 (N_23422,N_23038,N_23023);
or U23423 (N_23423,N_23034,N_23014);
nand U23424 (N_23424,N_23232,N_23245);
and U23425 (N_23425,N_23206,N_23014);
nand U23426 (N_23426,N_23080,N_23082);
or U23427 (N_23427,N_23100,N_23208);
and U23428 (N_23428,N_23191,N_23124);
or U23429 (N_23429,N_23158,N_23084);
xnor U23430 (N_23430,N_23209,N_23085);
and U23431 (N_23431,N_23077,N_23187);
or U23432 (N_23432,N_23151,N_23052);
and U23433 (N_23433,N_23149,N_23100);
xor U23434 (N_23434,N_23195,N_23231);
and U23435 (N_23435,N_23209,N_23048);
xor U23436 (N_23436,N_23197,N_23184);
and U23437 (N_23437,N_23195,N_23211);
nor U23438 (N_23438,N_23241,N_23222);
and U23439 (N_23439,N_23220,N_23121);
xnor U23440 (N_23440,N_23249,N_23002);
nor U23441 (N_23441,N_23134,N_23170);
and U23442 (N_23442,N_23128,N_23135);
and U23443 (N_23443,N_23232,N_23189);
and U23444 (N_23444,N_23078,N_23175);
nand U23445 (N_23445,N_23195,N_23018);
xor U23446 (N_23446,N_23069,N_23133);
or U23447 (N_23447,N_23133,N_23216);
or U23448 (N_23448,N_23211,N_23101);
nor U23449 (N_23449,N_23235,N_23118);
xor U23450 (N_23450,N_23186,N_23042);
nor U23451 (N_23451,N_23041,N_23078);
or U23452 (N_23452,N_23087,N_23235);
and U23453 (N_23453,N_23105,N_23149);
or U23454 (N_23454,N_23015,N_23011);
and U23455 (N_23455,N_23199,N_23169);
nor U23456 (N_23456,N_23112,N_23059);
or U23457 (N_23457,N_23116,N_23167);
and U23458 (N_23458,N_23125,N_23170);
xnor U23459 (N_23459,N_23135,N_23167);
xnor U23460 (N_23460,N_23144,N_23151);
and U23461 (N_23461,N_23017,N_23180);
and U23462 (N_23462,N_23078,N_23025);
or U23463 (N_23463,N_23166,N_23239);
and U23464 (N_23464,N_23098,N_23141);
and U23465 (N_23465,N_23185,N_23248);
or U23466 (N_23466,N_23218,N_23196);
xnor U23467 (N_23467,N_23100,N_23127);
xnor U23468 (N_23468,N_23199,N_23242);
nand U23469 (N_23469,N_23204,N_23092);
nand U23470 (N_23470,N_23203,N_23006);
or U23471 (N_23471,N_23174,N_23155);
and U23472 (N_23472,N_23033,N_23174);
nor U23473 (N_23473,N_23080,N_23108);
nor U23474 (N_23474,N_23173,N_23127);
nand U23475 (N_23475,N_23163,N_23017);
or U23476 (N_23476,N_23149,N_23079);
or U23477 (N_23477,N_23092,N_23158);
nor U23478 (N_23478,N_23132,N_23178);
nand U23479 (N_23479,N_23084,N_23002);
nor U23480 (N_23480,N_23219,N_23089);
nor U23481 (N_23481,N_23188,N_23100);
nand U23482 (N_23482,N_23012,N_23201);
nand U23483 (N_23483,N_23025,N_23190);
nor U23484 (N_23484,N_23155,N_23014);
nor U23485 (N_23485,N_23249,N_23211);
and U23486 (N_23486,N_23170,N_23085);
nand U23487 (N_23487,N_23076,N_23194);
or U23488 (N_23488,N_23094,N_23197);
or U23489 (N_23489,N_23194,N_23171);
and U23490 (N_23490,N_23046,N_23049);
nand U23491 (N_23491,N_23131,N_23015);
nand U23492 (N_23492,N_23106,N_23117);
and U23493 (N_23493,N_23189,N_23218);
nor U23494 (N_23494,N_23143,N_23208);
xor U23495 (N_23495,N_23164,N_23081);
and U23496 (N_23496,N_23179,N_23162);
xor U23497 (N_23497,N_23185,N_23155);
and U23498 (N_23498,N_23240,N_23133);
nand U23499 (N_23499,N_23015,N_23199);
nor U23500 (N_23500,N_23420,N_23367);
xnor U23501 (N_23501,N_23415,N_23302);
and U23502 (N_23502,N_23257,N_23478);
xor U23503 (N_23503,N_23431,N_23459);
or U23504 (N_23504,N_23316,N_23439);
nor U23505 (N_23505,N_23380,N_23476);
nor U23506 (N_23506,N_23301,N_23406);
nor U23507 (N_23507,N_23388,N_23340);
nor U23508 (N_23508,N_23352,N_23409);
and U23509 (N_23509,N_23314,N_23335);
and U23510 (N_23510,N_23371,N_23346);
or U23511 (N_23511,N_23399,N_23275);
nand U23512 (N_23512,N_23258,N_23325);
xnor U23513 (N_23513,N_23261,N_23324);
xor U23514 (N_23514,N_23473,N_23370);
and U23515 (N_23515,N_23477,N_23393);
or U23516 (N_23516,N_23444,N_23437);
or U23517 (N_23517,N_23338,N_23482);
and U23518 (N_23518,N_23354,N_23432);
or U23519 (N_23519,N_23445,N_23383);
or U23520 (N_23520,N_23462,N_23284);
nand U23521 (N_23521,N_23457,N_23305);
and U23522 (N_23522,N_23429,N_23253);
xor U23523 (N_23523,N_23372,N_23312);
or U23524 (N_23524,N_23475,N_23488);
xnor U23525 (N_23525,N_23298,N_23272);
nand U23526 (N_23526,N_23260,N_23493);
nor U23527 (N_23527,N_23452,N_23414);
or U23528 (N_23528,N_23355,N_23397);
and U23529 (N_23529,N_23296,N_23471);
nor U23530 (N_23530,N_23436,N_23299);
nor U23531 (N_23531,N_23274,N_23480);
xnor U23532 (N_23532,N_23322,N_23288);
nor U23533 (N_23533,N_23489,N_23492);
and U23534 (N_23534,N_23313,N_23448);
nand U23535 (N_23535,N_23470,N_23417);
and U23536 (N_23536,N_23333,N_23485);
xnor U23537 (N_23537,N_23418,N_23486);
nor U23538 (N_23538,N_23347,N_23433);
nand U23539 (N_23539,N_23369,N_23252);
nor U23540 (N_23540,N_23395,N_23401);
or U23541 (N_23541,N_23277,N_23293);
or U23542 (N_23542,N_23330,N_23434);
and U23543 (N_23543,N_23491,N_23270);
nor U23544 (N_23544,N_23430,N_23343);
and U23545 (N_23545,N_23311,N_23297);
nor U23546 (N_23546,N_23469,N_23494);
xnor U23547 (N_23547,N_23273,N_23416);
xnor U23548 (N_23548,N_23443,N_23267);
nor U23549 (N_23549,N_23402,N_23255);
nand U23550 (N_23550,N_23378,N_23421);
nor U23551 (N_23551,N_23425,N_23283);
xor U23552 (N_23552,N_23295,N_23349);
nor U23553 (N_23553,N_23392,N_23329);
xor U23554 (N_23554,N_23321,N_23428);
and U23555 (N_23555,N_23403,N_23407);
nor U23556 (N_23556,N_23308,N_23481);
or U23557 (N_23557,N_23483,N_23440);
xnor U23558 (N_23558,N_23353,N_23282);
or U23559 (N_23559,N_23398,N_23341);
or U23560 (N_23560,N_23490,N_23337);
xnor U23561 (N_23561,N_23310,N_23344);
nand U23562 (N_23562,N_23342,N_23495);
and U23563 (N_23563,N_23400,N_23360);
and U23564 (N_23564,N_23262,N_23307);
and U23565 (N_23565,N_23379,N_23405);
and U23566 (N_23566,N_23435,N_23366);
or U23567 (N_23567,N_23410,N_23396);
nand U23568 (N_23568,N_23384,N_23479);
nor U23569 (N_23569,N_23423,N_23368);
xnor U23570 (N_23570,N_23474,N_23467);
nor U23571 (N_23571,N_23361,N_23408);
xor U23572 (N_23572,N_23332,N_23362);
or U23573 (N_23573,N_23458,N_23454);
nor U23574 (N_23574,N_23281,N_23461);
or U23575 (N_23575,N_23315,N_23455);
nand U23576 (N_23576,N_23287,N_23442);
or U23577 (N_23577,N_23456,N_23358);
and U23578 (N_23578,N_23351,N_23345);
and U23579 (N_23579,N_23386,N_23357);
nand U23580 (N_23580,N_23375,N_23292);
and U23581 (N_23581,N_23278,N_23254);
xnor U23582 (N_23582,N_23496,N_23286);
nand U23583 (N_23583,N_23365,N_23450);
nor U23584 (N_23584,N_23256,N_23291);
and U23585 (N_23585,N_23497,N_23449);
nor U23586 (N_23586,N_23300,N_23447);
nand U23587 (N_23587,N_23466,N_23359);
nand U23588 (N_23588,N_23382,N_23327);
nand U23589 (N_23589,N_23276,N_23373);
nand U23590 (N_23590,N_23279,N_23460);
and U23591 (N_23591,N_23499,N_23320);
xnor U23592 (N_23592,N_23377,N_23427);
nor U23593 (N_23593,N_23289,N_23438);
nand U23594 (N_23594,N_23389,N_23463);
and U23595 (N_23595,N_23381,N_23309);
and U23596 (N_23596,N_23348,N_23451);
and U23597 (N_23597,N_23374,N_23364);
or U23598 (N_23598,N_23326,N_23391);
and U23599 (N_23599,N_23334,N_23350);
or U23600 (N_23600,N_23468,N_23411);
xnor U23601 (N_23601,N_23304,N_23356);
or U23602 (N_23602,N_23394,N_23317);
nand U23603 (N_23603,N_23303,N_23318);
or U23604 (N_23604,N_23285,N_23422);
xor U23605 (N_23605,N_23426,N_23336);
and U23606 (N_23606,N_23265,N_23419);
nand U23607 (N_23607,N_23453,N_23250);
or U23608 (N_23608,N_23363,N_23387);
nor U23609 (N_23609,N_23465,N_23264);
or U23610 (N_23610,N_23328,N_23263);
and U23611 (N_23611,N_23271,N_23331);
or U23612 (N_23612,N_23266,N_23424);
nand U23613 (N_23613,N_23269,N_23251);
nor U23614 (N_23614,N_23385,N_23376);
and U23615 (N_23615,N_23498,N_23472);
nor U23616 (N_23616,N_23294,N_23446);
xor U23617 (N_23617,N_23290,N_23268);
nand U23618 (N_23618,N_23319,N_23390);
nor U23619 (N_23619,N_23259,N_23280);
nand U23620 (N_23620,N_23306,N_23339);
xnor U23621 (N_23621,N_23412,N_23441);
or U23622 (N_23622,N_23413,N_23487);
xor U23623 (N_23623,N_23323,N_23484);
or U23624 (N_23624,N_23464,N_23404);
xnor U23625 (N_23625,N_23499,N_23348);
and U23626 (N_23626,N_23324,N_23457);
nor U23627 (N_23627,N_23387,N_23329);
nor U23628 (N_23628,N_23316,N_23253);
xor U23629 (N_23629,N_23358,N_23293);
nor U23630 (N_23630,N_23451,N_23491);
and U23631 (N_23631,N_23372,N_23253);
xor U23632 (N_23632,N_23415,N_23286);
xnor U23633 (N_23633,N_23265,N_23460);
xnor U23634 (N_23634,N_23437,N_23441);
nor U23635 (N_23635,N_23499,N_23428);
nand U23636 (N_23636,N_23423,N_23416);
nand U23637 (N_23637,N_23477,N_23294);
xnor U23638 (N_23638,N_23445,N_23448);
and U23639 (N_23639,N_23422,N_23367);
xor U23640 (N_23640,N_23342,N_23483);
or U23641 (N_23641,N_23450,N_23472);
xnor U23642 (N_23642,N_23359,N_23430);
or U23643 (N_23643,N_23290,N_23265);
or U23644 (N_23644,N_23401,N_23425);
nand U23645 (N_23645,N_23344,N_23251);
and U23646 (N_23646,N_23300,N_23277);
and U23647 (N_23647,N_23437,N_23364);
nand U23648 (N_23648,N_23283,N_23284);
nand U23649 (N_23649,N_23397,N_23496);
or U23650 (N_23650,N_23397,N_23448);
or U23651 (N_23651,N_23404,N_23281);
nand U23652 (N_23652,N_23477,N_23428);
or U23653 (N_23653,N_23397,N_23263);
xnor U23654 (N_23654,N_23482,N_23472);
or U23655 (N_23655,N_23360,N_23334);
and U23656 (N_23656,N_23365,N_23281);
xor U23657 (N_23657,N_23279,N_23375);
nor U23658 (N_23658,N_23425,N_23297);
xnor U23659 (N_23659,N_23487,N_23499);
nor U23660 (N_23660,N_23299,N_23284);
nor U23661 (N_23661,N_23416,N_23283);
and U23662 (N_23662,N_23374,N_23336);
nor U23663 (N_23663,N_23280,N_23494);
nand U23664 (N_23664,N_23478,N_23270);
xnor U23665 (N_23665,N_23277,N_23472);
xnor U23666 (N_23666,N_23296,N_23386);
xnor U23667 (N_23667,N_23412,N_23337);
and U23668 (N_23668,N_23455,N_23372);
nor U23669 (N_23669,N_23494,N_23327);
nand U23670 (N_23670,N_23423,N_23251);
and U23671 (N_23671,N_23370,N_23294);
nor U23672 (N_23672,N_23254,N_23308);
xor U23673 (N_23673,N_23374,N_23263);
nand U23674 (N_23674,N_23482,N_23381);
and U23675 (N_23675,N_23477,N_23258);
nor U23676 (N_23676,N_23464,N_23319);
and U23677 (N_23677,N_23282,N_23388);
nor U23678 (N_23678,N_23473,N_23351);
or U23679 (N_23679,N_23387,N_23337);
or U23680 (N_23680,N_23259,N_23348);
nor U23681 (N_23681,N_23280,N_23440);
or U23682 (N_23682,N_23432,N_23454);
nand U23683 (N_23683,N_23396,N_23458);
or U23684 (N_23684,N_23353,N_23259);
nor U23685 (N_23685,N_23433,N_23458);
or U23686 (N_23686,N_23404,N_23482);
or U23687 (N_23687,N_23344,N_23413);
nand U23688 (N_23688,N_23270,N_23285);
xor U23689 (N_23689,N_23468,N_23405);
and U23690 (N_23690,N_23498,N_23365);
nor U23691 (N_23691,N_23330,N_23341);
or U23692 (N_23692,N_23292,N_23401);
xor U23693 (N_23693,N_23325,N_23344);
nand U23694 (N_23694,N_23479,N_23336);
and U23695 (N_23695,N_23436,N_23347);
and U23696 (N_23696,N_23275,N_23408);
nand U23697 (N_23697,N_23469,N_23295);
nor U23698 (N_23698,N_23454,N_23256);
or U23699 (N_23699,N_23382,N_23416);
and U23700 (N_23700,N_23398,N_23417);
nor U23701 (N_23701,N_23451,N_23276);
xor U23702 (N_23702,N_23332,N_23369);
or U23703 (N_23703,N_23322,N_23302);
xnor U23704 (N_23704,N_23445,N_23389);
and U23705 (N_23705,N_23411,N_23420);
nor U23706 (N_23706,N_23403,N_23386);
xnor U23707 (N_23707,N_23306,N_23493);
nand U23708 (N_23708,N_23389,N_23353);
nor U23709 (N_23709,N_23388,N_23318);
or U23710 (N_23710,N_23408,N_23382);
nor U23711 (N_23711,N_23376,N_23485);
nor U23712 (N_23712,N_23422,N_23308);
xor U23713 (N_23713,N_23441,N_23429);
or U23714 (N_23714,N_23464,N_23435);
or U23715 (N_23715,N_23317,N_23444);
nor U23716 (N_23716,N_23409,N_23405);
and U23717 (N_23717,N_23410,N_23312);
and U23718 (N_23718,N_23333,N_23479);
or U23719 (N_23719,N_23263,N_23470);
and U23720 (N_23720,N_23285,N_23293);
and U23721 (N_23721,N_23263,N_23293);
nor U23722 (N_23722,N_23291,N_23408);
nor U23723 (N_23723,N_23423,N_23347);
xnor U23724 (N_23724,N_23413,N_23277);
nand U23725 (N_23725,N_23375,N_23364);
nor U23726 (N_23726,N_23387,N_23290);
xnor U23727 (N_23727,N_23414,N_23315);
or U23728 (N_23728,N_23427,N_23433);
or U23729 (N_23729,N_23370,N_23458);
xnor U23730 (N_23730,N_23278,N_23280);
xor U23731 (N_23731,N_23295,N_23487);
and U23732 (N_23732,N_23483,N_23320);
nor U23733 (N_23733,N_23305,N_23310);
nand U23734 (N_23734,N_23377,N_23477);
nor U23735 (N_23735,N_23343,N_23276);
and U23736 (N_23736,N_23353,N_23260);
nor U23737 (N_23737,N_23461,N_23472);
xor U23738 (N_23738,N_23250,N_23297);
nor U23739 (N_23739,N_23304,N_23293);
xnor U23740 (N_23740,N_23430,N_23379);
or U23741 (N_23741,N_23337,N_23390);
nand U23742 (N_23742,N_23450,N_23421);
nor U23743 (N_23743,N_23481,N_23290);
nor U23744 (N_23744,N_23410,N_23481);
or U23745 (N_23745,N_23433,N_23290);
nor U23746 (N_23746,N_23333,N_23425);
and U23747 (N_23747,N_23358,N_23329);
xor U23748 (N_23748,N_23253,N_23454);
nor U23749 (N_23749,N_23334,N_23389);
or U23750 (N_23750,N_23709,N_23573);
or U23751 (N_23751,N_23540,N_23735);
nor U23752 (N_23752,N_23680,N_23628);
nand U23753 (N_23753,N_23620,N_23506);
nor U23754 (N_23754,N_23626,N_23704);
and U23755 (N_23755,N_23731,N_23632);
nor U23756 (N_23756,N_23706,N_23523);
and U23757 (N_23757,N_23671,N_23600);
nor U23758 (N_23758,N_23705,N_23719);
xnor U23759 (N_23759,N_23589,N_23641);
or U23760 (N_23760,N_23592,N_23558);
nand U23761 (N_23761,N_23668,N_23739);
nor U23762 (N_23762,N_23733,N_23539);
nand U23763 (N_23763,N_23595,N_23529);
and U23764 (N_23764,N_23681,N_23684);
nor U23765 (N_23765,N_23574,N_23610);
xor U23766 (N_23766,N_23513,N_23655);
and U23767 (N_23767,N_23563,N_23745);
xnor U23768 (N_23768,N_23673,N_23640);
or U23769 (N_23769,N_23687,N_23561);
nor U23770 (N_23770,N_23581,N_23517);
nor U23771 (N_23771,N_23515,N_23617);
or U23772 (N_23772,N_23519,N_23518);
and U23773 (N_23773,N_23549,N_23612);
or U23774 (N_23774,N_23691,N_23500);
and U23775 (N_23775,N_23649,N_23590);
and U23776 (N_23776,N_23526,N_23746);
nand U23777 (N_23777,N_23550,N_23598);
xnor U23778 (N_23778,N_23588,N_23631);
xnor U23779 (N_23779,N_23737,N_23670);
and U23780 (N_23780,N_23696,N_23586);
nor U23781 (N_23781,N_23578,N_23742);
xnor U23782 (N_23782,N_23699,N_23514);
nor U23783 (N_23783,N_23591,N_23710);
nor U23784 (N_23784,N_23690,N_23676);
nand U23785 (N_23785,N_23535,N_23703);
xnor U23786 (N_23786,N_23524,N_23736);
xnor U23787 (N_23787,N_23516,N_23633);
xnor U23788 (N_23788,N_23510,N_23530);
or U23789 (N_23789,N_23553,N_23654);
nor U23790 (N_23790,N_23532,N_23570);
nand U23791 (N_23791,N_23741,N_23575);
or U23792 (N_23792,N_23643,N_23554);
nand U23793 (N_23793,N_23701,N_23718);
nor U23794 (N_23794,N_23541,N_23698);
and U23795 (N_23795,N_23527,N_23738);
and U23796 (N_23796,N_23501,N_23659);
or U23797 (N_23797,N_23700,N_23577);
and U23798 (N_23798,N_23548,N_23616);
xnor U23799 (N_23799,N_23707,N_23638);
xor U23800 (N_23800,N_23688,N_23503);
xor U23801 (N_23801,N_23666,N_23693);
or U23802 (N_23802,N_23722,N_23723);
xnor U23803 (N_23803,N_23508,N_23507);
or U23804 (N_23804,N_23725,N_23682);
xor U23805 (N_23805,N_23715,N_23579);
or U23806 (N_23806,N_23646,N_23656);
or U23807 (N_23807,N_23650,N_23545);
nand U23808 (N_23808,N_23502,N_23653);
and U23809 (N_23809,N_23686,N_23505);
or U23810 (N_23810,N_23747,N_23582);
xor U23811 (N_23811,N_23694,N_23645);
xor U23812 (N_23812,N_23615,N_23702);
and U23813 (N_23813,N_23717,N_23726);
nand U23814 (N_23814,N_23663,N_23629);
nand U23815 (N_23815,N_23713,N_23636);
xor U23816 (N_23816,N_23651,N_23544);
nand U23817 (N_23817,N_23624,N_23748);
and U23818 (N_23818,N_23622,N_23662);
xnor U23819 (N_23819,N_23607,N_23660);
xnor U23820 (N_23820,N_23634,N_23627);
and U23821 (N_23821,N_23674,N_23608);
nor U23822 (N_23822,N_23734,N_23743);
or U23823 (N_23823,N_23714,N_23728);
or U23824 (N_23824,N_23534,N_23552);
or U23825 (N_23825,N_23613,N_23611);
or U23826 (N_23826,N_23614,N_23585);
xnor U23827 (N_23827,N_23677,N_23587);
and U23828 (N_23828,N_23664,N_23565);
or U23829 (N_23829,N_23580,N_23732);
nor U23830 (N_23830,N_23559,N_23672);
or U23831 (N_23831,N_23716,N_23556);
or U23832 (N_23832,N_23547,N_23504);
nand U23833 (N_23833,N_23551,N_23536);
and U23834 (N_23834,N_23560,N_23749);
and U23835 (N_23835,N_23692,N_23685);
and U23836 (N_23836,N_23568,N_23623);
xor U23837 (N_23837,N_23721,N_23618);
xor U23838 (N_23838,N_23531,N_23630);
xnor U23839 (N_23839,N_23678,N_23555);
and U23840 (N_23840,N_23720,N_23724);
or U23841 (N_23841,N_23683,N_23730);
nor U23842 (N_23842,N_23571,N_23695);
nand U23843 (N_23843,N_23652,N_23667);
nand U23844 (N_23844,N_23657,N_23528);
nand U23845 (N_23845,N_23557,N_23594);
xnor U23846 (N_23846,N_23708,N_23661);
nor U23847 (N_23847,N_23546,N_23542);
xor U23848 (N_23848,N_23729,N_23711);
and U23849 (N_23849,N_23744,N_23522);
xnor U23850 (N_23850,N_23543,N_23603);
nand U23851 (N_23851,N_23605,N_23679);
nor U23852 (N_23852,N_23509,N_23583);
and U23853 (N_23853,N_23647,N_23689);
nand U23854 (N_23854,N_23533,N_23697);
xor U23855 (N_23855,N_23644,N_23538);
and U23856 (N_23856,N_23566,N_23621);
xor U23857 (N_23857,N_23512,N_23511);
nand U23858 (N_23858,N_23597,N_23625);
nand U23859 (N_23859,N_23601,N_23576);
nor U23860 (N_23860,N_23648,N_23599);
and U23861 (N_23861,N_23619,N_23604);
nand U23862 (N_23862,N_23637,N_23596);
nor U23863 (N_23863,N_23606,N_23569);
nand U23864 (N_23864,N_23521,N_23669);
or U23865 (N_23865,N_23639,N_23572);
nor U23866 (N_23866,N_23642,N_23537);
or U23867 (N_23867,N_23520,N_23635);
or U23868 (N_23868,N_23602,N_23584);
nor U23869 (N_23869,N_23727,N_23665);
or U23870 (N_23870,N_23609,N_23593);
or U23871 (N_23871,N_23564,N_23658);
nand U23872 (N_23872,N_23740,N_23567);
or U23873 (N_23873,N_23525,N_23712);
nor U23874 (N_23874,N_23562,N_23675);
nor U23875 (N_23875,N_23699,N_23554);
and U23876 (N_23876,N_23621,N_23510);
and U23877 (N_23877,N_23727,N_23688);
xnor U23878 (N_23878,N_23721,N_23682);
and U23879 (N_23879,N_23564,N_23737);
nand U23880 (N_23880,N_23700,N_23551);
or U23881 (N_23881,N_23570,N_23665);
nand U23882 (N_23882,N_23563,N_23744);
nor U23883 (N_23883,N_23521,N_23703);
and U23884 (N_23884,N_23588,N_23700);
xnor U23885 (N_23885,N_23613,N_23742);
nor U23886 (N_23886,N_23624,N_23562);
nand U23887 (N_23887,N_23721,N_23670);
xnor U23888 (N_23888,N_23596,N_23528);
and U23889 (N_23889,N_23622,N_23523);
nor U23890 (N_23890,N_23682,N_23500);
nor U23891 (N_23891,N_23657,N_23561);
xor U23892 (N_23892,N_23500,N_23617);
and U23893 (N_23893,N_23642,N_23736);
nor U23894 (N_23894,N_23619,N_23571);
and U23895 (N_23895,N_23720,N_23625);
or U23896 (N_23896,N_23718,N_23537);
xnor U23897 (N_23897,N_23699,N_23574);
nor U23898 (N_23898,N_23530,N_23583);
nor U23899 (N_23899,N_23661,N_23523);
nand U23900 (N_23900,N_23621,N_23705);
or U23901 (N_23901,N_23642,N_23687);
or U23902 (N_23902,N_23504,N_23681);
and U23903 (N_23903,N_23578,N_23696);
or U23904 (N_23904,N_23743,N_23594);
nand U23905 (N_23905,N_23685,N_23538);
nor U23906 (N_23906,N_23681,N_23622);
and U23907 (N_23907,N_23637,N_23723);
nand U23908 (N_23908,N_23628,N_23558);
and U23909 (N_23909,N_23661,N_23684);
or U23910 (N_23910,N_23644,N_23588);
xnor U23911 (N_23911,N_23586,N_23530);
nand U23912 (N_23912,N_23542,N_23744);
nor U23913 (N_23913,N_23656,N_23634);
nor U23914 (N_23914,N_23697,N_23625);
and U23915 (N_23915,N_23687,N_23570);
nor U23916 (N_23916,N_23676,N_23677);
or U23917 (N_23917,N_23529,N_23574);
nor U23918 (N_23918,N_23671,N_23633);
xor U23919 (N_23919,N_23629,N_23626);
and U23920 (N_23920,N_23591,N_23638);
or U23921 (N_23921,N_23601,N_23698);
nor U23922 (N_23922,N_23564,N_23688);
and U23923 (N_23923,N_23509,N_23663);
xnor U23924 (N_23924,N_23695,N_23747);
nor U23925 (N_23925,N_23659,N_23671);
nor U23926 (N_23926,N_23733,N_23713);
nor U23927 (N_23927,N_23641,N_23616);
or U23928 (N_23928,N_23711,N_23635);
or U23929 (N_23929,N_23541,N_23649);
xnor U23930 (N_23930,N_23673,N_23566);
nand U23931 (N_23931,N_23652,N_23712);
nand U23932 (N_23932,N_23701,N_23681);
nor U23933 (N_23933,N_23642,N_23578);
and U23934 (N_23934,N_23698,N_23645);
nand U23935 (N_23935,N_23690,N_23581);
nand U23936 (N_23936,N_23554,N_23508);
xor U23937 (N_23937,N_23528,N_23521);
nand U23938 (N_23938,N_23670,N_23636);
nand U23939 (N_23939,N_23737,N_23524);
or U23940 (N_23940,N_23651,N_23503);
xor U23941 (N_23941,N_23597,N_23686);
and U23942 (N_23942,N_23573,N_23530);
xor U23943 (N_23943,N_23741,N_23724);
nor U23944 (N_23944,N_23594,N_23698);
and U23945 (N_23945,N_23585,N_23700);
or U23946 (N_23946,N_23713,N_23704);
xor U23947 (N_23947,N_23709,N_23546);
nand U23948 (N_23948,N_23584,N_23632);
nor U23949 (N_23949,N_23738,N_23559);
nor U23950 (N_23950,N_23558,N_23749);
nor U23951 (N_23951,N_23622,N_23542);
nand U23952 (N_23952,N_23636,N_23691);
nor U23953 (N_23953,N_23590,N_23506);
or U23954 (N_23954,N_23721,N_23637);
xor U23955 (N_23955,N_23558,N_23694);
xor U23956 (N_23956,N_23508,N_23696);
and U23957 (N_23957,N_23600,N_23636);
xor U23958 (N_23958,N_23636,N_23512);
nor U23959 (N_23959,N_23598,N_23529);
xor U23960 (N_23960,N_23654,N_23604);
or U23961 (N_23961,N_23594,N_23573);
nand U23962 (N_23962,N_23661,N_23560);
nor U23963 (N_23963,N_23604,N_23516);
nor U23964 (N_23964,N_23645,N_23656);
or U23965 (N_23965,N_23685,N_23671);
and U23966 (N_23966,N_23566,N_23554);
nand U23967 (N_23967,N_23547,N_23693);
or U23968 (N_23968,N_23740,N_23539);
nor U23969 (N_23969,N_23542,N_23506);
xor U23970 (N_23970,N_23710,N_23717);
or U23971 (N_23971,N_23721,N_23591);
or U23972 (N_23972,N_23740,N_23735);
and U23973 (N_23973,N_23533,N_23739);
xnor U23974 (N_23974,N_23686,N_23711);
nor U23975 (N_23975,N_23696,N_23617);
nand U23976 (N_23976,N_23710,N_23663);
nor U23977 (N_23977,N_23569,N_23673);
and U23978 (N_23978,N_23587,N_23700);
xor U23979 (N_23979,N_23556,N_23650);
nand U23980 (N_23980,N_23538,N_23731);
nand U23981 (N_23981,N_23721,N_23559);
nor U23982 (N_23982,N_23736,N_23738);
nand U23983 (N_23983,N_23548,N_23742);
or U23984 (N_23984,N_23730,N_23681);
nand U23985 (N_23985,N_23632,N_23505);
xor U23986 (N_23986,N_23620,N_23641);
nand U23987 (N_23987,N_23577,N_23623);
or U23988 (N_23988,N_23534,N_23717);
xnor U23989 (N_23989,N_23518,N_23510);
or U23990 (N_23990,N_23574,N_23506);
and U23991 (N_23991,N_23685,N_23748);
or U23992 (N_23992,N_23666,N_23687);
and U23993 (N_23993,N_23544,N_23729);
xnor U23994 (N_23994,N_23507,N_23558);
nor U23995 (N_23995,N_23511,N_23667);
or U23996 (N_23996,N_23641,N_23728);
nor U23997 (N_23997,N_23679,N_23745);
and U23998 (N_23998,N_23650,N_23712);
or U23999 (N_23999,N_23721,N_23517);
xor U24000 (N_24000,N_23947,N_23924);
and U24001 (N_24001,N_23772,N_23964);
and U24002 (N_24002,N_23974,N_23796);
and U24003 (N_24003,N_23936,N_23976);
and U24004 (N_24004,N_23833,N_23789);
nand U24005 (N_24005,N_23793,N_23786);
and U24006 (N_24006,N_23930,N_23882);
nand U24007 (N_24007,N_23889,N_23783);
nand U24008 (N_24008,N_23944,N_23809);
nor U24009 (N_24009,N_23760,N_23826);
or U24010 (N_24010,N_23819,N_23825);
nand U24011 (N_24011,N_23913,N_23777);
nand U24012 (N_24012,N_23822,N_23850);
and U24013 (N_24013,N_23957,N_23784);
or U24014 (N_24014,N_23869,N_23755);
nor U24015 (N_24015,N_23762,N_23846);
nor U24016 (N_24016,N_23842,N_23958);
xnor U24017 (N_24017,N_23855,N_23968);
nand U24018 (N_24018,N_23778,N_23960);
nand U24019 (N_24019,N_23851,N_23770);
nand U24020 (N_24020,N_23798,N_23890);
xor U24021 (N_24021,N_23971,N_23990);
xnor U24022 (N_24022,N_23844,N_23907);
or U24023 (N_24023,N_23986,N_23830);
xnor U24024 (N_24024,N_23916,N_23909);
xor U24025 (N_24025,N_23982,N_23969);
and U24026 (N_24026,N_23859,N_23802);
xor U24027 (N_24027,N_23921,N_23884);
nand U24028 (N_24028,N_23813,N_23901);
and U24029 (N_24029,N_23781,N_23761);
nand U24030 (N_24030,N_23827,N_23775);
xnor U24031 (N_24031,N_23945,N_23911);
nor U24032 (N_24032,N_23992,N_23979);
or U24033 (N_24033,N_23956,N_23984);
nor U24034 (N_24034,N_23896,N_23991);
xor U24035 (N_24035,N_23865,N_23828);
xor U24036 (N_24036,N_23817,N_23995);
xor U24037 (N_24037,N_23792,N_23765);
xor U24038 (N_24038,N_23906,N_23811);
xnor U24039 (N_24039,N_23900,N_23878);
and U24040 (N_24040,N_23949,N_23997);
nand U24041 (N_24041,N_23815,N_23973);
nand U24042 (N_24042,N_23863,N_23885);
and U24043 (N_24043,N_23816,N_23894);
and U24044 (N_24044,N_23933,N_23773);
nand U24045 (N_24045,N_23860,N_23920);
or U24046 (N_24046,N_23763,N_23790);
and U24047 (N_24047,N_23751,N_23866);
nor U24048 (N_24048,N_23998,N_23797);
or U24049 (N_24049,N_23824,N_23862);
and U24050 (N_24050,N_23961,N_23795);
and U24051 (N_24051,N_23852,N_23895);
nand U24052 (N_24052,N_23867,N_23829);
nand U24053 (N_24053,N_23953,N_23768);
xnor U24054 (N_24054,N_23854,N_23805);
or U24055 (N_24055,N_23937,N_23899);
or U24056 (N_24056,N_23931,N_23800);
or U24057 (N_24057,N_23856,N_23983);
or U24058 (N_24058,N_23774,N_23905);
and U24059 (N_24059,N_23837,N_23951);
nand U24060 (N_24060,N_23987,N_23922);
xor U24061 (N_24061,N_23950,N_23831);
or U24062 (N_24062,N_23888,N_23902);
nand U24063 (N_24063,N_23893,N_23794);
nor U24064 (N_24064,N_23874,N_23972);
and U24065 (N_24065,N_23988,N_23750);
nand U24066 (N_24066,N_23757,N_23870);
nand U24067 (N_24067,N_23771,N_23927);
nor U24068 (N_24068,N_23941,N_23847);
nand U24069 (N_24069,N_23868,N_23977);
or U24070 (N_24070,N_23806,N_23864);
xor U24071 (N_24071,N_23914,N_23871);
nand U24072 (N_24072,N_23999,N_23919);
xor U24073 (N_24073,N_23801,N_23845);
nor U24074 (N_24074,N_23980,N_23952);
and U24075 (N_24075,N_23994,N_23766);
xnor U24076 (N_24076,N_23932,N_23873);
or U24077 (N_24077,N_23915,N_23752);
nor U24078 (N_24078,N_23823,N_23756);
xnor U24079 (N_24079,N_23883,N_23904);
nor U24080 (N_24080,N_23876,N_23776);
nand U24081 (N_24081,N_23887,N_23807);
xor U24082 (N_24082,N_23935,N_23955);
nor U24083 (N_24083,N_23892,N_23965);
nor U24084 (N_24084,N_23840,N_23926);
xnor U24085 (N_24085,N_23903,N_23767);
nand U24086 (N_24086,N_23942,N_23910);
or U24087 (N_24087,N_23934,N_23948);
and U24088 (N_24088,N_23804,N_23978);
and U24089 (N_24089,N_23908,N_23753);
or U24090 (N_24090,N_23966,N_23970);
and U24091 (N_24091,N_23923,N_23897);
or U24092 (N_24092,N_23848,N_23779);
or U24093 (N_24093,N_23985,N_23791);
or U24094 (N_24094,N_23917,N_23843);
xnor U24095 (N_24095,N_23981,N_23853);
or U24096 (N_24096,N_23818,N_23993);
and U24097 (N_24097,N_23954,N_23886);
nand U24098 (N_24098,N_23785,N_23989);
nand U24099 (N_24099,N_23839,N_23759);
xor U24100 (N_24100,N_23912,N_23879);
or U24101 (N_24101,N_23803,N_23808);
nor U24102 (N_24102,N_23925,N_23754);
or U24103 (N_24103,N_23857,N_23861);
nor U24104 (N_24104,N_23872,N_23769);
nor U24105 (N_24105,N_23943,N_23836);
and U24106 (N_24106,N_23963,N_23929);
xnor U24107 (N_24107,N_23996,N_23849);
xnor U24108 (N_24108,N_23810,N_23940);
nand U24109 (N_24109,N_23780,N_23799);
and U24110 (N_24110,N_23814,N_23881);
or U24111 (N_24111,N_23832,N_23939);
nor U24112 (N_24112,N_23788,N_23918);
and U24113 (N_24113,N_23938,N_23834);
nand U24114 (N_24114,N_23975,N_23898);
nand U24115 (N_24115,N_23959,N_23821);
nor U24116 (N_24116,N_23838,N_23891);
nor U24117 (N_24117,N_23758,N_23764);
or U24118 (N_24118,N_23787,N_23835);
or U24119 (N_24119,N_23820,N_23880);
nand U24120 (N_24120,N_23782,N_23946);
nand U24121 (N_24121,N_23928,N_23858);
nand U24122 (N_24122,N_23877,N_23812);
xnor U24123 (N_24123,N_23841,N_23875);
nand U24124 (N_24124,N_23967,N_23962);
and U24125 (N_24125,N_23999,N_23766);
xor U24126 (N_24126,N_23765,N_23979);
and U24127 (N_24127,N_23830,N_23883);
or U24128 (N_24128,N_23838,N_23813);
nand U24129 (N_24129,N_23752,N_23918);
or U24130 (N_24130,N_23923,N_23763);
nor U24131 (N_24131,N_23899,N_23985);
xor U24132 (N_24132,N_23853,N_23795);
nand U24133 (N_24133,N_23981,N_23882);
nand U24134 (N_24134,N_23925,N_23848);
nand U24135 (N_24135,N_23846,N_23965);
xor U24136 (N_24136,N_23985,N_23754);
or U24137 (N_24137,N_23974,N_23797);
xor U24138 (N_24138,N_23988,N_23946);
nor U24139 (N_24139,N_23838,N_23879);
or U24140 (N_24140,N_23750,N_23897);
and U24141 (N_24141,N_23912,N_23759);
nor U24142 (N_24142,N_23806,N_23931);
or U24143 (N_24143,N_23831,N_23879);
or U24144 (N_24144,N_23982,N_23994);
and U24145 (N_24145,N_23882,N_23860);
nor U24146 (N_24146,N_23868,N_23982);
xor U24147 (N_24147,N_23856,N_23792);
or U24148 (N_24148,N_23904,N_23874);
or U24149 (N_24149,N_23876,N_23902);
nor U24150 (N_24150,N_23820,N_23983);
nor U24151 (N_24151,N_23940,N_23839);
nand U24152 (N_24152,N_23765,N_23755);
xor U24153 (N_24153,N_23974,N_23898);
xor U24154 (N_24154,N_23770,N_23771);
nand U24155 (N_24155,N_23859,N_23964);
and U24156 (N_24156,N_23992,N_23785);
xnor U24157 (N_24157,N_23922,N_23982);
and U24158 (N_24158,N_23872,N_23856);
and U24159 (N_24159,N_23834,N_23832);
xor U24160 (N_24160,N_23856,N_23841);
xnor U24161 (N_24161,N_23806,N_23779);
nor U24162 (N_24162,N_23924,N_23888);
and U24163 (N_24163,N_23768,N_23823);
xnor U24164 (N_24164,N_23773,N_23846);
or U24165 (N_24165,N_23948,N_23971);
or U24166 (N_24166,N_23790,N_23921);
xnor U24167 (N_24167,N_23756,N_23983);
nor U24168 (N_24168,N_23753,N_23808);
nor U24169 (N_24169,N_23948,N_23897);
nand U24170 (N_24170,N_23857,N_23845);
nand U24171 (N_24171,N_23806,N_23814);
or U24172 (N_24172,N_23898,N_23938);
and U24173 (N_24173,N_23886,N_23916);
nand U24174 (N_24174,N_23963,N_23968);
and U24175 (N_24175,N_23830,N_23884);
and U24176 (N_24176,N_23955,N_23773);
or U24177 (N_24177,N_23793,N_23859);
and U24178 (N_24178,N_23992,N_23900);
nand U24179 (N_24179,N_23979,N_23895);
xnor U24180 (N_24180,N_23959,N_23998);
or U24181 (N_24181,N_23855,N_23954);
nand U24182 (N_24182,N_23921,N_23775);
or U24183 (N_24183,N_23796,N_23809);
nand U24184 (N_24184,N_23951,N_23906);
and U24185 (N_24185,N_23938,N_23809);
nand U24186 (N_24186,N_23887,N_23995);
and U24187 (N_24187,N_23977,N_23878);
and U24188 (N_24188,N_23769,N_23802);
xor U24189 (N_24189,N_23786,N_23800);
and U24190 (N_24190,N_23872,N_23768);
or U24191 (N_24191,N_23879,N_23871);
nor U24192 (N_24192,N_23900,N_23861);
and U24193 (N_24193,N_23953,N_23887);
and U24194 (N_24194,N_23933,N_23869);
or U24195 (N_24195,N_23991,N_23887);
nor U24196 (N_24196,N_23989,N_23828);
and U24197 (N_24197,N_23820,N_23989);
and U24198 (N_24198,N_23857,N_23997);
xnor U24199 (N_24199,N_23870,N_23806);
and U24200 (N_24200,N_23769,N_23853);
and U24201 (N_24201,N_23929,N_23826);
nand U24202 (N_24202,N_23796,N_23752);
and U24203 (N_24203,N_23930,N_23927);
xnor U24204 (N_24204,N_23990,N_23891);
xnor U24205 (N_24205,N_23979,N_23990);
and U24206 (N_24206,N_23957,N_23939);
and U24207 (N_24207,N_23784,N_23897);
xor U24208 (N_24208,N_23868,N_23785);
nor U24209 (N_24209,N_23814,N_23750);
nand U24210 (N_24210,N_23758,N_23937);
nand U24211 (N_24211,N_23925,N_23808);
nand U24212 (N_24212,N_23845,N_23914);
and U24213 (N_24213,N_23969,N_23779);
or U24214 (N_24214,N_23993,N_23932);
nand U24215 (N_24215,N_23771,N_23932);
or U24216 (N_24216,N_23898,N_23754);
nor U24217 (N_24217,N_23930,N_23801);
xor U24218 (N_24218,N_23887,N_23852);
nor U24219 (N_24219,N_23844,N_23989);
nand U24220 (N_24220,N_23984,N_23780);
and U24221 (N_24221,N_23897,N_23961);
nand U24222 (N_24222,N_23930,N_23964);
nand U24223 (N_24223,N_23963,N_23822);
nand U24224 (N_24224,N_23805,N_23996);
xnor U24225 (N_24225,N_23834,N_23833);
nor U24226 (N_24226,N_23862,N_23877);
and U24227 (N_24227,N_23951,N_23942);
or U24228 (N_24228,N_23766,N_23988);
nand U24229 (N_24229,N_23954,N_23989);
and U24230 (N_24230,N_23864,N_23786);
and U24231 (N_24231,N_23970,N_23905);
and U24232 (N_24232,N_23900,N_23894);
or U24233 (N_24233,N_23918,N_23770);
nor U24234 (N_24234,N_23773,N_23839);
nand U24235 (N_24235,N_23774,N_23766);
and U24236 (N_24236,N_23859,N_23871);
nor U24237 (N_24237,N_23947,N_23996);
or U24238 (N_24238,N_23973,N_23971);
or U24239 (N_24239,N_23976,N_23938);
and U24240 (N_24240,N_23856,N_23879);
or U24241 (N_24241,N_23978,N_23955);
nor U24242 (N_24242,N_23837,N_23919);
and U24243 (N_24243,N_23944,N_23948);
nor U24244 (N_24244,N_23826,N_23906);
or U24245 (N_24245,N_23757,N_23888);
xnor U24246 (N_24246,N_23853,N_23846);
nor U24247 (N_24247,N_23914,N_23911);
xnor U24248 (N_24248,N_23823,N_23884);
nand U24249 (N_24249,N_23881,N_23866);
and U24250 (N_24250,N_24055,N_24149);
and U24251 (N_24251,N_24027,N_24021);
and U24252 (N_24252,N_24126,N_24164);
xnor U24253 (N_24253,N_24185,N_24045);
or U24254 (N_24254,N_24060,N_24096);
or U24255 (N_24255,N_24051,N_24201);
or U24256 (N_24256,N_24176,N_24030);
and U24257 (N_24257,N_24139,N_24024);
nor U24258 (N_24258,N_24241,N_24142);
nor U24259 (N_24259,N_24206,N_24076);
xor U24260 (N_24260,N_24050,N_24087);
xnor U24261 (N_24261,N_24239,N_24015);
nor U24262 (N_24262,N_24049,N_24160);
and U24263 (N_24263,N_24235,N_24177);
nor U24264 (N_24264,N_24012,N_24029);
or U24265 (N_24265,N_24213,N_24210);
and U24266 (N_24266,N_24218,N_24208);
and U24267 (N_24267,N_24072,N_24028);
nand U24268 (N_24268,N_24156,N_24234);
and U24269 (N_24269,N_24220,N_24165);
nor U24270 (N_24270,N_24007,N_24247);
nand U24271 (N_24271,N_24046,N_24033);
nor U24272 (N_24272,N_24248,N_24170);
xor U24273 (N_24273,N_24143,N_24097);
nand U24274 (N_24274,N_24168,N_24152);
and U24275 (N_24275,N_24074,N_24070);
nor U24276 (N_24276,N_24205,N_24184);
or U24277 (N_24277,N_24061,N_24082);
nor U24278 (N_24278,N_24124,N_24047);
xnor U24279 (N_24279,N_24132,N_24243);
nor U24280 (N_24280,N_24141,N_24219);
nand U24281 (N_24281,N_24066,N_24058);
xnor U24282 (N_24282,N_24180,N_24067);
xnor U24283 (N_24283,N_24145,N_24036);
xnor U24284 (N_24284,N_24018,N_24221);
and U24285 (N_24285,N_24212,N_24071);
or U24286 (N_24286,N_24113,N_24104);
nor U24287 (N_24287,N_24122,N_24068);
nand U24288 (N_24288,N_24056,N_24001);
nand U24289 (N_24289,N_24038,N_24016);
xnor U24290 (N_24290,N_24137,N_24034);
nand U24291 (N_24291,N_24227,N_24059);
nand U24292 (N_24292,N_24150,N_24065);
or U24293 (N_24293,N_24192,N_24217);
and U24294 (N_24294,N_24228,N_24188);
xor U24295 (N_24295,N_24080,N_24053);
nand U24296 (N_24296,N_24092,N_24231);
and U24297 (N_24297,N_24014,N_24040);
or U24298 (N_24298,N_24244,N_24002);
nor U24299 (N_24299,N_24005,N_24200);
nor U24300 (N_24300,N_24008,N_24009);
nor U24301 (N_24301,N_24109,N_24181);
xor U24302 (N_24302,N_24240,N_24166);
nor U24303 (N_24303,N_24173,N_24161);
nor U24304 (N_24304,N_24107,N_24086);
nand U24305 (N_24305,N_24245,N_24020);
xor U24306 (N_24306,N_24062,N_24064);
xnor U24307 (N_24307,N_24136,N_24182);
and U24308 (N_24308,N_24138,N_24171);
nand U24309 (N_24309,N_24083,N_24195);
or U24310 (N_24310,N_24183,N_24130);
nand U24311 (N_24311,N_24098,N_24088);
nand U24312 (N_24312,N_24127,N_24131);
nand U24313 (N_24313,N_24154,N_24000);
nand U24314 (N_24314,N_24054,N_24091);
and U24315 (N_24315,N_24148,N_24134);
nor U24316 (N_24316,N_24155,N_24224);
and U24317 (N_24317,N_24174,N_24204);
and U24318 (N_24318,N_24095,N_24202);
or U24319 (N_24319,N_24114,N_24099);
or U24320 (N_24320,N_24193,N_24031);
nand U24321 (N_24321,N_24026,N_24004);
nor U24322 (N_24322,N_24094,N_24222);
and U24323 (N_24323,N_24118,N_24246);
xor U24324 (N_24324,N_24108,N_24189);
nor U24325 (N_24325,N_24112,N_24159);
xor U24326 (N_24326,N_24163,N_24116);
nor U24327 (N_24327,N_24078,N_24199);
or U24328 (N_24328,N_24135,N_24090);
nor U24329 (N_24329,N_24207,N_24057);
and U24330 (N_24330,N_24025,N_24223);
nand U24331 (N_24331,N_24215,N_24129);
and U24332 (N_24332,N_24191,N_24117);
or U24333 (N_24333,N_24011,N_24186);
nor U24334 (N_24334,N_24119,N_24037);
nand U24335 (N_24335,N_24102,N_24178);
xnor U24336 (N_24336,N_24225,N_24172);
nor U24337 (N_24337,N_24237,N_24035);
or U24338 (N_24338,N_24209,N_24106);
and U24339 (N_24339,N_24190,N_24187);
or U24340 (N_24340,N_24133,N_24100);
xor U24341 (N_24341,N_24075,N_24003);
nand U24342 (N_24342,N_24214,N_24048);
nor U24343 (N_24343,N_24128,N_24196);
and U24344 (N_24344,N_24044,N_24052);
xnor U24345 (N_24345,N_24194,N_24063);
and U24346 (N_24346,N_24238,N_24022);
nor U24347 (N_24347,N_24023,N_24085);
nand U24348 (N_24348,N_24013,N_24144);
and U24349 (N_24349,N_24169,N_24110);
xnor U24350 (N_24350,N_24198,N_24147);
or U24351 (N_24351,N_24242,N_24069);
and U24352 (N_24352,N_24249,N_24121);
and U24353 (N_24353,N_24236,N_24089);
or U24354 (N_24354,N_24032,N_24115);
nor U24355 (N_24355,N_24230,N_24146);
and U24356 (N_24356,N_24081,N_24093);
nor U24357 (N_24357,N_24216,N_24006);
and U24358 (N_24358,N_24010,N_24203);
and U24359 (N_24359,N_24151,N_24120);
nor U24360 (N_24360,N_24105,N_24197);
or U24361 (N_24361,N_24140,N_24157);
xnor U24362 (N_24362,N_24211,N_24229);
nand U24363 (N_24363,N_24162,N_24232);
nor U24364 (N_24364,N_24084,N_24158);
or U24365 (N_24365,N_24017,N_24077);
or U24366 (N_24366,N_24101,N_24167);
or U24367 (N_24367,N_24043,N_24233);
or U24368 (N_24368,N_24153,N_24079);
nand U24369 (N_24369,N_24175,N_24039);
and U24370 (N_24370,N_24019,N_24042);
or U24371 (N_24371,N_24123,N_24041);
nor U24372 (N_24372,N_24111,N_24073);
and U24373 (N_24373,N_24179,N_24226);
xnor U24374 (N_24374,N_24103,N_24125);
xnor U24375 (N_24375,N_24120,N_24152);
and U24376 (N_24376,N_24060,N_24205);
nor U24377 (N_24377,N_24092,N_24083);
or U24378 (N_24378,N_24090,N_24106);
nor U24379 (N_24379,N_24127,N_24228);
nand U24380 (N_24380,N_24207,N_24217);
or U24381 (N_24381,N_24047,N_24154);
xnor U24382 (N_24382,N_24125,N_24212);
or U24383 (N_24383,N_24245,N_24040);
and U24384 (N_24384,N_24222,N_24091);
nand U24385 (N_24385,N_24218,N_24077);
or U24386 (N_24386,N_24042,N_24222);
or U24387 (N_24387,N_24166,N_24070);
nand U24388 (N_24388,N_24246,N_24093);
nor U24389 (N_24389,N_24243,N_24065);
nand U24390 (N_24390,N_24001,N_24245);
xnor U24391 (N_24391,N_24124,N_24204);
nor U24392 (N_24392,N_24012,N_24228);
nor U24393 (N_24393,N_24241,N_24189);
nor U24394 (N_24394,N_24043,N_24020);
or U24395 (N_24395,N_24237,N_24143);
nor U24396 (N_24396,N_24048,N_24241);
nand U24397 (N_24397,N_24031,N_24026);
nand U24398 (N_24398,N_24083,N_24003);
nand U24399 (N_24399,N_24139,N_24245);
nand U24400 (N_24400,N_24217,N_24110);
and U24401 (N_24401,N_24120,N_24169);
or U24402 (N_24402,N_24052,N_24149);
or U24403 (N_24403,N_24032,N_24096);
and U24404 (N_24404,N_24116,N_24139);
xnor U24405 (N_24405,N_24151,N_24148);
and U24406 (N_24406,N_24138,N_24011);
nand U24407 (N_24407,N_24075,N_24004);
and U24408 (N_24408,N_24096,N_24049);
or U24409 (N_24409,N_24154,N_24126);
or U24410 (N_24410,N_24142,N_24205);
or U24411 (N_24411,N_24158,N_24170);
or U24412 (N_24412,N_24153,N_24031);
xor U24413 (N_24413,N_24218,N_24034);
or U24414 (N_24414,N_24091,N_24167);
nor U24415 (N_24415,N_24096,N_24076);
nand U24416 (N_24416,N_24083,N_24156);
or U24417 (N_24417,N_24109,N_24160);
or U24418 (N_24418,N_24122,N_24196);
or U24419 (N_24419,N_24000,N_24004);
xor U24420 (N_24420,N_24207,N_24186);
xnor U24421 (N_24421,N_24093,N_24201);
nand U24422 (N_24422,N_24055,N_24137);
or U24423 (N_24423,N_24061,N_24211);
and U24424 (N_24424,N_24175,N_24074);
nand U24425 (N_24425,N_24139,N_24119);
nor U24426 (N_24426,N_24219,N_24111);
nor U24427 (N_24427,N_24118,N_24134);
nor U24428 (N_24428,N_24146,N_24164);
nor U24429 (N_24429,N_24071,N_24185);
or U24430 (N_24430,N_24118,N_24122);
and U24431 (N_24431,N_24065,N_24163);
and U24432 (N_24432,N_24239,N_24228);
nand U24433 (N_24433,N_24139,N_24198);
and U24434 (N_24434,N_24086,N_24119);
or U24435 (N_24435,N_24139,N_24200);
xnor U24436 (N_24436,N_24159,N_24071);
nand U24437 (N_24437,N_24111,N_24023);
or U24438 (N_24438,N_24197,N_24217);
xor U24439 (N_24439,N_24097,N_24206);
nand U24440 (N_24440,N_24000,N_24060);
nand U24441 (N_24441,N_24135,N_24056);
or U24442 (N_24442,N_24179,N_24028);
and U24443 (N_24443,N_24015,N_24221);
xor U24444 (N_24444,N_24056,N_24185);
nand U24445 (N_24445,N_24011,N_24192);
xnor U24446 (N_24446,N_24049,N_24231);
xor U24447 (N_24447,N_24236,N_24245);
xor U24448 (N_24448,N_24131,N_24011);
nand U24449 (N_24449,N_24073,N_24205);
xnor U24450 (N_24450,N_24172,N_24201);
or U24451 (N_24451,N_24014,N_24000);
nand U24452 (N_24452,N_24065,N_24204);
nand U24453 (N_24453,N_24168,N_24240);
and U24454 (N_24454,N_24172,N_24128);
and U24455 (N_24455,N_24131,N_24021);
nand U24456 (N_24456,N_24025,N_24242);
and U24457 (N_24457,N_24035,N_24197);
nor U24458 (N_24458,N_24112,N_24111);
and U24459 (N_24459,N_24238,N_24019);
nand U24460 (N_24460,N_24191,N_24216);
nor U24461 (N_24461,N_24044,N_24036);
or U24462 (N_24462,N_24068,N_24179);
xor U24463 (N_24463,N_24245,N_24232);
or U24464 (N_24464,N_24156,N_24072);
nor U24465 (N_24465,N_24033,N_24100);
nand U24466 (N_24466,N_24141,N_24100);
and U24467 (N_24467,N_24224,N_24202);
or U24468 (N_24468,N_24160,N_24186);
nor U24469 (N_24469,N_24152,N_24022);
nor U24470 (N_24470,N_24205,N_24041);
nor U24471 (N_24471,N_24017,N_24023);
xor U24472 (N_24472,N_24087,N_24145);
nor U24473 (N_24473,N_24176,N_24014);
xor U24474 (N_24474,N_24081,N_24013);
and U24475 (N_24475,N_24162,N_24212);
xor U24476 (N_24476,N_24167,N_24243);
nand U24477 (N_24477,N_24210,N_24249);
nor U24478 (N_24478,N_24035,N_24056);
xor U24479 (N_24479,N_24102,N_24222);
and U24480 (N_24480,N_24174,N_24161);
and U24481 (N_24481,N_24133,N_24170);
nand U24482 (N_24482,N_24214,N_24010);
xnor U24483 (N_24483,N_24127,N_24115);
nor U24484 (N_24484,N_24202,N_24226);
xnor U24485 (N_24485,N_24115,N_24121);
and U24486 (N_24486,N_24021,N_24112);
nor U24487 (N_24487,N_24212,N_24088);
or U24488 (N_24488,N_24016,N_24197);
and U24489 (N_24489,N_24082,N_24170);
nor U24490 (N_24490,N_24050,N_24070);
nor U24491 (N_24491,N_24000,N_24151);
or U24492 (N_24492,N_24214,N_24153);
xor U24493 (N_24493,N_24085,N_24044);
or U24494 (N_24494,N_24138,N_24001);
xnor U24495 (N_24495,N_24053,N_24115);
and U24496 (N_24496,N_24249,N_24240);
nand U24497 (N_24497,N_24106,N_24166);
and U24498 (N_24498,N_24006,N_24198);
nand U24499 (N_24499,N_24116,N_24083);
nor U24500 (N_24500,N_24320,N_24397);
nand U24501 (N_24501,N_24414,N_24260);
or U24502 (N_24502,N_24360,N_24310);
and U24503 (N_24503,N_24454,N_24257);
and U24504 (N_24504,N_24271,N_24351);
or U24505 (N_24505,N_24490,N_24424);
or U24506 (N_24506,N_24412,N_24350);
nor U24507 (N_24507,N_24492,N_24438);
nand U24508 (N_24508,N_24436,N_24488);
and U24509 (N_24509,N_24285,N_24406);
nand U24510 (N_24510,N_24461,N_24371);
nand U24511 (N_24511,N_24275,N_24370);
xnor U24512 (N_24512,N_24264,N_24347);
and U24513 (N_24513,N_24384,N_24443);
or U24514 (N_24514,N_24317,N_24319);
and U24515 (N_24515,N_24330,N_24445);
xnor U24516 (N_24516,N_24250,N_24314);
nor U24517 (N_24517,N_24372,N_24368);
nand U24518 (N_24518,N_24463,N_24324);
or U24519 (N_24519,N_24427,N_24491);
xor U24520 (N_24520,N_24263,N_24392);
or U24521 (N_24521,N_24423,N_24383);
nand U24522 (N_24522,N_24439,N_24378);
and U24523 (N_24523,N_24356,N_24440);
xor U24524 (N_24524,N_24312,N_24309);
and U24525 (N_24525,N_24286,N_24410);
or U24526 (N_24526,N_24321,N_24366);
or U24527 (N_24527,N_24281,N_24333);
and U24528 (N_24528,N_24477,N_24459);
nor U24529 (N_24529,N_24484,N_24299);
xor U24530 (N_24530,N_24395,N_24270);
and U24531 (N_24531,N_24290,N_24465);
and U24532 (N_24532,N_24448,N_24399);
and U24533 (N_24533,N_24442,N_24404);
nor U24534 (N_24534,N_24352,N_24482);
or U24535 (N_24535,N_24498,N_24437);
nor U24536 (N_24536,N_24287,N_24307);
xor U24537 (N_24537,N_24369,N_24365);
nand U24538 (N_24538,N_24481,N_24435);
xnor U24539 (N_24539,N_24431,N_24421);
and U24540 (N_24540,N_24425,N_24466);
xor U24541 (N_24541,N_24272,N_24306);
nor U24542 (N_24542,N_24411,N_24475);
nor U24543 (N_24543,N_24456,N_24326);
nor U24544 (N_24544,N_24362,N_24273);
nor U24545 (N_24545,N_24485,N_24432);
or U24546 (N_24546,N_24495,N_24297);
nor U24547 (N_24547,N_24305,N_24296);
xor U24548 (N_24548,N_24478,N_24429);
and U24549 (N_24549,N_24345,N_24358);
nor U24550 (N_24550,N_24403,N_24308);
or U24551 (N_24551,N_24487,N_24269);
nand U24552 (N_24552,N_24434,N_24256);
nor U24553 (N_24553,N_24254,N_24420);
nand U24554 (N_24554,N_24262,N_24449);
or U24555 (N_24555,N_24496,N_24280);
xor U24556 (N_24556,N_24494,N_24340);
nor U24557 (N_24557,N_24289,N_24328);
nor U24558 (N_24558,N_24258,N_24470);
or U24559 (N_24559,N_24323,N_24376);
or U24560 (N_24560,N_24381,N_24278);
xor U24561 (N_24561,N_24288,N_24332);
xnor U24562 (N_24562,N_24268,N_24348);
nand U24563 (N_24563,N_24302,N_24407);
or U24564 (N_24564,N_24355,N_24468);
nand U24565 (N_24565,N_24359,N_24329);
and U24566 (N_24566,N_24253,N_24393);
nor U24567 (N_24567,N_24325,N_24460);
or U24568 (N_24568,N_24451,N_24398);
xor U24569 (N_24569,N_24417,N_24419);
nand U24570 (N_24570,N_24444,N_24473);
nor U24571 (N_24571,N_24334,N_24400);
or U24572 (N_24572,N_24251,N_24318);
xor U24573 (N_24573,N_24388,N_24474);
nand U24574 (N_24574,N_24430,N_24316);
nor U24575 (N_24575,N_24338,N_24480);
xnor U24576 (N_24576,N_24416,N_24402);
nor U24577 (N_24577,N_24337,N_24277);
or U24578 (N_24578,N_24386,N_24300);
nand U24579 (N_24579,N_24266,N_24315);
nor U24580 (N_24580,N_24301,N_24489);
xnor U24581 (N_24581,N_24426,N_24422);
nand U24582 (N_24582,N_24298,N_24344);
or U24583 (N_24583,N_24303,N_24469);
or U24584 (N_24584,N_24394,N_24295);
nor U24585 (N_24585,N_24457,N_24343);
xnor U24586 (N_24586,N_24331,N_24339);
and U24587 (N_24587,N_24364,N_24354);
nor U24588 (N_24588,N_24472,N_24396);
nor U24589 (N_24589,N_24336,N_24294);
nor U24590 (N_24590,N_24390,N_24479);
nand U24591 (N_24591,N_24433,N_24346);
and U24592 (N_24592,N_24274,N_24313);
or U24593 (N_24593,N_24265,N_24453);
or U24594 (N_24594,N_24405,N_24375);
nand U24595 (N_24595,N_24379,N_24493);
nor U24596 (N_24596,N_24455,N_24483);
nand U24597 (N_24597,N_24418,N_24342);
or U24598 (N_24598,N_24322,N_24497);
and U24599 (N_24599,N_24335,N_24367);
nor U24600 (N_24600,N_24374,N_24450);
nand U24601 (N_24601,N_24284,N_24380);
nand U24602 (N_24602,N_24471,N_24349);
or U24603 (N_24603,N_24255,N_24408);
nand U24604 (N_24604,N_24283,N_24292);
or U24605 (N_24605,N_24259,N_24357);
nor U24606 (N_24606,N_24293,N_24389);
nand U24607 (N_24607,N_24464,N_24387);
xor U24608 (N_24608,N_24462,N_24291);
nor U24609 (N_24609,N_24252,N_24363);
and U24610 (N_24610,N_24327,N_24447);
or U24611 (N_24611,N_24353,N_24361);
and U24612 (N_24612,N_24452,N_24377);
or U24613 (N_24613,N_24428,N_24415);
nor U24614 (N_24614,N_24304,N_24476);
xor U24615 (N_24615,N_24279,N_24341);
or U24616 (N_24616,N_24373,N_24276);
nor U24617 (N_24617,N_24413,N_24267);
nor U24618 (N_24618,N_24382,N_24499);
or U24619 (N_24619,N_24391,N_24401);
nor U24620 (N_24620,N_24385,N_24486);
and U24621 (N_24621,N_24409,N_24311);
or U24622 (N_24622,N_24282,N_24446);
nand U24623 (N_24623,N_24441,N_24467);
and U24624 (N_24624,N_24261,N_24458);
nor U24625 (N_24625,N_24303,N_24431);
nand U24626 (N_24626,N_24432,N_24479);
nor U24627 (N_24627,N_24401,N_24424);
nand U24628 (N_24628,N_24497,N_24423);
or U24629 (N_24629,N_24358,N_24269);
nand U24630 (N_24630,N_24279,N_24250);
nand U24631 (N_24631,N_24255,N_24275);
nand U24632 (N_24632,N_24398,N_24294);
xnor U24633 (N_24633,N_24404,N_24405);
nand U24634 (N_24634,N_24336,N_24399);
xor U24635 (N_24635,N_24361,N_24316);
nor U24636 (N_24636,N_24416,N_24385);
or U24637 (N_24637,N_24270,N_24399);
or U24638 (N_24638,N_24490,N_24369);
or U24639 (N_24639,N_24389,N_24350);
nor U24640 (N_24640,N_24339,N_24361);
or U24641 (N_24641,N_24274,N_24391);
xor U24642 (N_24642,N_24396,N_24491);
nand U24643 (N_24643,N_24389,N_24304);
or U24644 (N_24644,N_24324,N_24473);
nand U24645 (N_24645,N_24459,N_24294);
nand U24646 (N_24646,N_24284,N_24444);
xor U24647 (N_24647,N_24496,N_24369);
xnor U24648 (N_24648,N_24407,N_24403);
nand U24649 (N_24649,N_24378,N_24323);
nor U24650 (N_24650,N_24425,N_24412);
nor U24651 (N_24651,N_24484,N_24457);
nor U24652 (N_24652,N_24367,N_24344);
nand U24653 (N_24653,N_24302,N_24369);
xnor U24654 (N_24654,N_24357,N_24403);
nand U24655 (N_24655,N_24483,N_24472);
or U24656 (N_24656,N_24311,N_24380);
nand U24657 (N_24657,N_24311,N_24357);
and U24658 (N_24658,N_24410,N_24401);
nor U24659 (N_24659,N_24361,N_24449);
xor U24660 (N_24660,N_24471,N_24493);
and U24661 (N_24661,N_24448,N_24394);
nor U24662 (N_24662,N_24354,N_24482);
xor U24663 (N_24663,N_24457,N_24472);
nand U24664 (N_24664,N_24374,N_24424);
xor U24665 (N_24665,N_24278,N_24423);
nand U24666 (N_24666,N_24360,N_24458);
and U24667 (N_24667,N_24377,N_24463);
or U24668 (N_24668,N_24424,N_24451);
or U24669 (N_24669,N_24453,N_24469);
or U24670 (N_24670,N_24285,N_24398);
nor U24671 (N_24671,N_24426,N_24399);
and U24672 (N_24672,N_24272,N_24369);
nand U24673 (N_24673,N_24280,N_24404);
or U24674 (N_24674,N_24488,N_24287);
nand U24675 (N_24675,N_24321,N_24396);
xor U24676 (N_24676,N_24402,N_24437);
nand U24677 (N_24677,N_24440,N_24381);
nand U24678 (N_24678,N_24383,N_24314);
nor U24679 (N_24679,N_24360,N_24402);
nor U24680 (N_24680,N_24320,N_24485);
xor U24681 (N_24681,N_24385,N_24254);
nand U24682 (N_24682,N_24453,N_24263);
or U24683 (N_24683,N_24266,N_24400);
and U24684 (N_24684,N_24272,N_24417);
or U24685 (N_24685,N_24276,N_24492);
nand U24686 (N_24686,N_24337,N_24369);
nand U24687 (N_24687,N_24457,N_24482);
nor U24688 (N_24688,N_24296,N_24326);
or U24689 (N_24689,N_24257,N_24281);
xor U24690 (N_24690,N_24407,N_24315);
xor U24691 (N_24691,N_24460,N_24290);
xor U24692 (N_24692,N_24288,N_24283);
xor U24693 (N_24693,N_24319,N_24483);
nand U24694 (N_24694,N_24434,N_24496);
nor U24695 (N_24695,N_24304,N_24429);
and U24696 (N_24696,N_24272,N_24478);
nor U24697 (N_24697,N_24479,N_24254);
and U24698 (N_24698,N_24496,N_24324);
xor U24699 (N_24699,N_24467,N_24369);
or U24700 (N_24700,N_24481,N_24262);
xor U24701 (N_24701,N_24329,N_24455);
xor U24702 (N_24702,N_24372,N_24497);
nand U24703 (N_24703,N_24394,N_24319);
nor U24704 (N_24704,N_24258,N_24317);
nand U24705 (N_24705,N_24391,N_24366);
or U24706 (N_24706,N_24276,N_24439);
nor U24707 (N_24707,N_24379,N_24477);
or U24708 (N_24708,N_24438,N_24406);
nand U24709 (N_24709,N_24253,N_24447);
or U24710 (N_24710,N_24304,N_24448);
xnor U24711 (N_24711,N_24463,N_24308);
nand U24712 (N_24712,N_24300,N_24344);
nor U24713 (N_24713,N_24362,N_24418);
nand U24714 (N_24714,N_24367,N_24283);
xnor U24715 (N_24715,N_24436,N_24393);
or U24716 (N_24716,N_24310,N_24354);
xnor U24717 (N_24717,N_24441,N_24283);
nor U24718 (N_24718,N_24325,N_24461);
nor U24719 (N_24719,N_24476,N_24300);
or U24720 (N_24720,N_24383,N_24421);
nand U24721 (N_24721,N_24381,N_24288);
and U24722 (N_24722,N_24376,N_24281);
nand U24723 (N_24723,N_24262,N_24474);
or U24724 (N_24724,N_24256,N_24338);
or U24725 (N_24725,N_24275,N_24351);
nor U24726 (N_24726,N_24398,N_24390);
or U24727 (N_24727,N_24394,N_24476);
nand U24728 (N_24728,N_24269,N_24310);
nand U24729 (N_24729,N_24334,N_24346);
nand U24730 (N_24730,N_24399,N_24381);
xor U24731 (N_24731,N_24345,N_24301);
or U24732 (N_24732,N_24388,N_24429);
or U24733 (N_24733,N_24318,N_24393);
nor U24734 (N_24734,N_24403,N_24477);
nor U24735 (N_24735,N_24458,N_24369);
xor U24736 (N_24736,N_24358,N_24417);
and U24737 (N_24737,N_24375,N_24250);
xor U24738 (N_24738,N_24346,N_24491);
or U24739 (N_24739,N_24260,N_24408);
and U24740 (N_24740,N_24420,N_24366);
nand U24741 (N_24741,N_24269,N_24413);
nand U24742 (N_24742,N_24351,N_24374);
or U24743 (N_24743,N_24273,N_24347);
xor U24744 (N_24744,N_24477,N_24352);
nor U24745 (N_24745,N_24251,N_24433);
nor U24746 (N_24746,N_24330,N_24471);
or U24747 (N_24747,N_24267,N_24258);
nor U24748 (N_24748,N_24260,N_24441);
xnor U24749 (N_24749,N_24471,N_24426);
nand U24750 (N_24750,N_24680,N_24513);
or U24751 (N_24751,N_24661,N_24718);
nor U24752 (N_24752,N_24635,N_24583);
or U24753 (N_24753,N_24567,N_24674);
nand U24754 (N_24754,N_24686,N_24707);
xnor U24755 (N_24755,N_24730,N_24521);
xnor U24756 (N_24756,N_24526,N_24738);
xnor U24757 (N_24757,N_24664,N_24594);
xnor U24758 (N_24758,N_24740,N_24511);
nor U24759 (N_24759,N_24610,N_24589);
xnor U24760 (N_24760,N_24532,N_24667);
nor U24761 (N_24761,N_24590,N_24616);
or U24762 (N_24762,N_24705,N_24697);
xnor U24763 (N_24763,N_24563,N_24681);
or U24764 (N_24764,N_24595,N_24617);
or U24765 (N_24765,N_24582,N_24679);
nor U24766 (N_24766,N_24712,N_24646);
and U24767 (N_24767,N_24519,N_24500);
nor U24768 (N_24768,N_24554,N_24572);
nand U24769 (N_24769,N_24578,N_24742);
and U24770 (N_24770,N_24503,N_24613);
and U24771 (N_24771,N_24621,N_24630);
nand U24772 (N_24772,N_24651,N_24638);
nand U24773 (N_24773,N_24642,N_24668);
nor U24774 (N_24774,N_24660,N_24748);
nor U24775 (N_24775,N_24569,N_24605);
nor U24776 (N_24776,N_24531,N_24555);
nor U24777 (N_24777,N_24598,N_24645);
or U24778 (N_24778,N_24706,N_24538);
and U24779 (N_24779,N_24641,N_24637);
nor U24780 (N_24780,N_24746,N_24544);
xnor U24781 (N_24781,N_24525,N_24696);
and U24782 (N_24782,N_24647,N_24708);
nor U24783 (N_24783,N_24650,N_24643);
and U24784 (N_24784,N_24741,N_24684);
xor U24785 (N_24785,N_24655,N_24510);
or U24786 (N_24786,N_24716,N_24722);
nand U24787 (N_24787,N_24723,N_24656);
xor U24788 (N_24788,N_24600,N_24714);
nand U24789 (N_24789,N_24733,N_24715);
xnor U24790 (N_24790,N_24677,N_24729);
nand U24791 (N_24791,N_24559,N_24632);
xnor U24792 (N_24792,N_24506,N_24556);
or U24793 (N_24793,N_24739,N_24703);
and U24794 (N_24794,N_24626,N_24634);
nand U24795 (N_24795,N_24720,N_24585);
and U24796 (N_24796,N_24501,N_24725);
and U24797 (N_24797,N_24537,N_24601);
nor U24798 (N_24798,N_24719,N_24573);
nand U24799 (N_24799,N_24628,N_24694);
and U24800 (N_24800,N_24542,N_24522);
xor U24801 (N_24801,N_24553,N_24608);
and U24802 (N_24802,N_24709,N_24691);
nor U24803 (N_24803,N_24736,N_24614);
and U24804 (N_24804,N_24700,N_24695);
xor U24805 (N_24805,N_24744,N_24631);
xnor U24806 (N_24806,N_24561,N_24579);
or U24807 (N_24807,N_24574,N_24524);
nand U24808 (N_24808,N_24689,N_24508);
and U24809 (N_24809,N_24625,N_24570);
nand U24810 (N_24810,N_24704,N_24682);
xnor U24811 (N_24811,N_24548,N_24654);
nor U24812 (N_24812,N_24669,N_24512);
or U24813 (N_24813,N_24504,N_24665);
xor U24814 (N_24814,N_24575,N_24732);
nor U24815 (N_24815,N_24698,N_24530);
xor U24816 (N_24816,N_24534,N_24620);
nor U24817 (N_24817,N_24676,N_24586);
nor U24818 (N_24818,N_24612,N_24653);
nor U24819 (N_24819,N_24721,N_24566);
nor U24820 (N_24820,N_24547,N_24516);
xnor U24821 (N_24821,N_24685,N_24591);
nor U24822 (N_24822,N_24536,N_24564);
nand U24823 (N_24823,N_24520,N_24603);
nor U24824 (N_24824,N_24673,N_24692);
and U24825 (N_24825,N_24747,N_24727);
xor U24826 (N_24826,N_24699,N_24640);
and U24827 (N_24827,N_24558,N_24675);
nand U24828 (N_24828,N_24662,N_24701);
nand U24829 (N_24829,N_24596,N_24545);
or U24830 (N_24830,N_24517,N_24629);
nand U24831 (N_24831,N_24728,N_24606);
nor U24832 (N_24832,N_24502,N_24568);
and U24833 (N_24833,N_24562,N_24514);
or U24834 (N_24834,N_24607,N_24602);
nand U24835 (N_24835,N_24518,N_24731);
xnor U24836 (N_24836,N_24659,N_24505);
and U24837 (N_24837,N_24549,N_24584);
nand U24838 (N_24838,N_24541,N_24551);
nand U24839 (N_24839,N_24533,N_24648);
nand U24840 (N_24840,N_24576,N_24749);
nor U24841 (N_24841,N_24611,N_24627);
nor U24842 (N_24842,N_24507,N_24652);
or U24843 (N_24843,N_24609,N_24672);
nand U24844 (N_24844,N_24633,N_24529);
nand U24845 (N_24845,N_24670,N_24539);
nor U24846 (N_24846,N_24509,N_24565);
xor U24847 (N_24847,N_24587,N_24683);
or U24848 (N_24848,N_24717,N_24571);
nand U24849 (N_24849,N_24619,N_24639);
xor U24850 (N_24850,N_24688,N_24552);
xnor U24851 (N_24851,N_24693,N_24711);
nor U24852 (N_24852,N_24702,N_24624);
nor U24853 (N_24853,N_24649,N_24540);
nor U24854 (N_24854,N_24557,N_24726);
nand U24855 (N_24855,N_24527,N_24724);
nor U24856 (N_24856,N_24710,N_24644);
and U24857 (N_24857,N_24618,N_24604);
or U24858 (N_24858,N_24599,N_24523);
and U24859 (N_24859,N_24658,N_24622);
xor U24860 (N_24860,N_24615,N_24593);
nand U24861 (N_24861,N_24690,N_24687);
nor U24862 (N_24862,N_24543,N_24623);
nor U24863 (N_24863,N_24592,N_24528);
or U24864 (N_24864,N_24745,N_24743);
nor U24865 (N_24865,N_24588,N_24577);
nor U24866 (N_24866,N_24515,N_24597);
and U24867 (N_24867,N_24657,N_24581);
and U24868 (N_24868,N_24678,N_24737);
nand U24869 (N_24869,N_24580,N_24713);
and U24870 (N_24870,N_24734,N_24546);
nor U24871 (N_24871,N_24735,N_24663);
nand U24872 (N_24872,N_24636,N_24666);
nor U24873 (N_24873,N_24671,N_24535);
or U24874 (N_24874,N_24560,N_24550);
and U24875 (N_24875,N_24656,N_24585);
xor U24876 (N_24876,N_24516,N_24633);
and U24877 (N_24877,N_24654,N_24746);
nor U24878 (N_24878,N_24673,N_24737);
and U24879 (N_24879,N_24701,N_24720);
and U24880 (N_24880,N_24527,N_24583);
xnor U24881 (N_24881,N_24545,N_24724);
nand U24882 (N_24882,N_24726,N_24749);
xnor U24883 (N_24883,N_24639,N_24594);
or U24884 (N_24884,N_24649,N_24546);
nor U24885 (N_24885,N_24650,N_24515);
or U24886 (N_24886,N_24508,N_24723);
nor U24887 (N_24887,N_24718,N_24731);
xor U24888 (N_24888,N_24696,N_24545);
nand U24889 (N_24889,N_24561,N_24727);
or U24890 (N_24890,N_24510,N_24526);
nand U24891 (N_24891,N_24732,N_24613);
xnor U24892 (N_24892,N_24657,N_24736);
nor U24893 (N_24893,N_24722,N_24665);
xnor U24894 (N_24894,N_24592,N_24632);
or U24895 (N_24895,N_24562,N_24529);
or U24896 (N_24896,N_24643,N_24518);
xnor U24897 (N_24897,N_24723,N_24633);
and U24898 (N_24898,N_24510,N_24728);
xor U24899 (N_24899,N_24575,N_24725);
xnor U24900 (N_24900,N_24747,N_24577);
xnor U24901 (N_24901,N_24655,N_24654);
and U24902 (N_24902,N_24531,N_24505);
xnor U24903 (N_24903,N_24650,N_24664);
and U24904 (N_24904,N_24702,N_24732);
nand U24905 (N_24905,N_24722,N_24654);
and U24906 (N_24906,N_24523,N_24605);
nand U24907 (N_24907,N_24712,N_24593);
or U24908 (N_24908,N_24558,N_24684);
and U24909 (N_24909,N_24620,N_24537);
nand U24910 (N_24910,N_24538,N_24516);
nor U24911 (N_24911,N_24566,N_24694);
or U24912 (N_24912,N_24528,N_24559);
nand U24913 (N_24913,N_24674,N_24740);
xnor U24914 (N_24914,N_24730,N_24563);
nor U24915 (N_24915,N_24611,N_24725);
or U24916 (N_24916,N_24503,N_24725);
xor U24917 (N_24917,N_24562,N_24617);
nand U24918 (N_24918,N_24536,N_24684);
xnor U24919 (N_24919,N_24656,N_24523);
and U24920 (N_24920,N_24705,N_24669);
and U24921 (N_24921,N_24679,N_24724);
nand U24922 (N_24922,N_24640,N_24548);
nor U24923 (N_24923,N_24506,N_24722);
nand U24924 (N_24924,N_24590,N_24648);
nand U24925 (N_24925,N_24524,N_24590);
nand U24926 (N_24926,N_24591,N_24592);
nor U24927 (N_24927,N_24629,N_24686);
nand U24928 (N_24928,N_24731,N_24584);
nand U24929 (N_24929,N_24616,N_24651);
and U24930 (N_24930,N_24666,N_24670);
nand U24931 (N_24931,N_24634,N_24625);
nor U24932 (N_24932,N_24591,N_24634);
nor U24933 (N_24933,N_24643,N_24723);
and U24934 (N_24934,N_24719,N_24743);
nor U24935 (N_24935,N_24522,N_24562);
and U24936 (N_24936,N_24600,N_24585);
and U24937 (N_24937,N_24579,N_24557);
xor U24938 (N_24938,N_24695,N_24574);
nand U24939 (N_24939,N_24746,N_24712);
nor U24940 (N_24940,N_24696,N_24543);
or U24941 (N_24941,N_24614,N_24677);
or U24942 (N_24942,N_24735,N_24501);
or U24943 (N_24943,N_24727,N_24549);
and U24944 (N_24944,N_24504,N_24742);
nand U24945 (N_24945,N_24713,N_24575);
xnor U24946 (N_24946,N_24671,N_24533);
nand U24947 (N_24947,N_24638,N_24728);
xnor U24948 (N_24948,N_24573,N_24726);
xor U24949 (N_24949,N_24650,N_24595);
xnor U24950 (N_24950,N_24616,N_24547);
or U24951 (N_24951,N_24610,N_24715);
nor U24952 (N_24952,N_24514,N_24703);
xor U24953 (N_24953,N_24520,N_24591);
nor U24954 (N_24954,N_24636,N_24630);
xnor U24955 (N_24955,N_24708,N_24619);
nand U24956 (N_24956,N_24546,N_24718);
or U24957 (N_24957,N_24532,N_24588);
or U24958 (N_24958,N_24615,N_24643);
xor U24959 (N_24959,N_24717,N_24582);
nand U24960 (N_24960,N_24679,N_24601);
nor U24961 (N_24961,N_24683,N_24620);
or U24962 (N_24962,N_24603,N_24541);
nand U24963 (N_24963,N_24665,N_24530);
and U24964 (N_24964,N_24633,N_24514);
and U24965 (N_24965,N_24596,N_24582);
xnor U24966 (N_24966,N_24746,N_24720);
nand U24967 (N_24967,N_24721,N_24589);
and U24968 (N_24968,N_24729,N_24633);
or U24969 (N_24969,N_24546,N_24612);
or U24970 (N_24970,N_24717,N_24657);
xor U24971 (N_24971,N_24584,N_24738);
or U24972 (N_24972,N_24675,N_24598);
and U24973 (N_24973,N_24563,N_24651);
or U24974 (N_24974,N_24681,N_24705);
or U24975 (N_24975,N_24536,N_24682);
nand U24976 (N_24976,N_24729,N_24583);
nand U24977 (N_24977,N_24687,N_24570);
nor U24978 (N_24978,N_24540,N_24697);
xor U24979 (N_24979,N_24727,N_24595);
and U24980 (N_24980,N_24651,N_24746);
nand U24981 (N_24981,N_24703,N_24501);
nor U24982 (N_24982,N_24687,N_24746);
nor U24983 (N_24983,N_24524,N_24515);
or U24984 (N_24984,N_24640,N_24623);
and U24985 (N_24985,N_24732,N_24664);
nand U24986 (N_24986,N_24679,N_24583);
xnor U24987 (N_24987,N_24667,N_24572);
nor U24988 (N_24988,N_24655,N_24516);
xnor U24989 (N_24989,N_24702,N_24585);
and U24990 (N_24990,N_24651,N_24594);
xor U24991 (N_24991,N_24547,N_24602);
nor U24992 (N_24992,N_24674,N_24586);
nand U24993 (N_24993,N_24675,N_24714);
and U24994 (N_24994,N_24500,N_24736);
or U24995 (N_24995,N_24627,N_24624);
and U24996 (N_24996,N_24731,N_24507);
or U24997 (N_24997,N_24658,N_24578);
and U24998 (N_24998,N_24623,N_24510);
or U24999 (N_24999,N_24535,N_24693);
and U25000 (N_25000,N_24821,N_24871);
xor U25001 (N_25001,N_24964,N_24895);
nor U25002 (N_25002,N_24826,N_24990);
and U25003 (N_25003,N_24856,N_24979);
nor U25004 (N_25004,N_24845,N_24893);
xnor U25005 (N_25005,N_24973,N_24811);
xor U25006 (N_25006,N_24862,N_24864);
or U25007 (N_25007,N_24995,N_24839);
and U25008 (N_25008,N_24897,N_24974);
or U25009 (N_25009,N_24789,N_24752);
or U25010 (N_25010,N_24955,N_24779);
nor U25011 (N_25011,N_24967,N_24928);
nand U25012 (N_25012,N_24970,N_24798);
nand U25013 (N_25013,N_24874,N_24932);
or U25014 (N_25014,N_24926,N_24805);
nand U25015 (N_25015,N_24940,N_24914);
nor U25016 (N_25016,N_24983,N_24911);
nand U25017 (N_25017,N_24832,N_24971);
or U25018 (N_25018,N_24807,N_24818);
and U25019 (N_25019,N_24880,N_24925);
xnor U25020 (N_25020,N_24896,N_24778);
nand U25021 (N_25021,N_24793,N_24799);
nand U25022 (N_25022,N_24959,N_24987);
nor U25023 (N_25023,N_24849,N_24867);
nor U25024 (N_25024,N_24958,N_24943);
nor U25025 (N_25025,N_24755,N_24878);
nor U25026 (N_25026,N_24782,N_24840);
or U25027 (N_25027,N_24763,N_24823);
or U25028 (N_25028,N_24868,N_24774);
and U25029 (N_25029,N_24873,N_24976);
or U25030 (N_25030,N_24942,N_24927);
xor U25031 (N_25031,N_24820,N_24800);
nand U25032 (N_25032,N_24848,N_24772);
nand U25033 (N_25033,N_24788,N_24853);
and U25034 (N_25034,N_24946,N_24756);
or U25035 (N_25035,N_24757,N_24859);
xnor U25036 (N_25036,N_24750,N_24773);
nor U25037 (N_25037,N_24751,N_24830);
or U25038 (N_25038,N_24934,N_24919);
and U25039 (N_25039,N_24888,N_24760);
xor U25040 (N_25040,N_24828,N_24953);
nand U25041 (N_25041,N_24858,N_24909);
xor U25042 (N_25042,N_24803,N_24775);
and U25043 (N_25043,N_24816,N_24819);
nand U25044 (N_25044,N_24835,N_24978);
or U25045 (N_25045,N_24836,N_24908);
nor U25046 (N_25046,N_24781,N_24777);
nor U25047 (N_25047,N_24851,N_24977);
and U25048 (N_25048,N_24872,N_24804);
nand U25049 (N_25049,N_24857,N_24981);
or U25050 (N_25050,N_24843,N_24956);
or U25051 (N_25051,N_24808,N_24762);
and U25052 (N_25052,N_24822,N_24949);
xor U25053 (N_25053,N_24861,N_24850);
or U25054 (N_25054,N_24935,N_24838);
and U25055 (N_25055,N_24992,N_24863);
nand U25056 (N_25056,N_24910,N_24892);
xor U25057 (N_25057,N_24969,N_24837);
nand U25058 (N_25058,N_24931,N_24792);
and U25059 (N_25059,N_24802,N_24882);
nor U25060 (N_25060,N_24814,N_24783);
or U25061 (N_25061,N_24945,N_24817);
and U25062 (N_25062,N_24986,N_24997);
nand U25063 (N_25063,N_24759,N_24860);
nand U25064 (N_25064,N_24769,N_24916);
xnor U25065 (N_25065,N_24869,N_24930);
nor U25066 (N_25066,N_24846,N_24922);
nand U25067 (N_25067,N_24771,N_24877);
and U25068 (N_25068,N_24827,N_24797);
nand U25069 (N_25069,N_24966,N_24766);
nor U25070 (N_25070,N_24950,N_24963);
and U25071 (N_25071,N_24954,N_24770);
and U25072 (N_25072,N_24883,N_24948);
or U25073 (N_25073,N_24847,N_24993);
or U25074 (N_25074,N_24902,N_24806);
nor U25075 (N_25075,N_24885,N_24938);
or U25076 (N_25076,N_24984,N_24785);
or U25077 (N_25077,N_24894,N_24913);
xor U25078 (N_25078,N_24903,N_24982);
or U25079 (N_25079,N_24812,N_24960);
nor U25080 (N_25080,N_24929,N_24917);
nand U25081 (N_25081,N_24944,N_24939);
or U25082 (N_25082,N_24923,N_24865);
or U25083 (N_25083,N_24852,N_24936);
or U25084 (N_25084,N_24933,N_24780);
or U25085 (N_25085,N_24975,N_24831);
nand U25086 (N_25086,N_24899,N_24957);
xor U25087 (N_25087,N_24898,N_24810);
or U25088 (N_25088,N_24972,N_24854);
nor U25089 (N_25089,N_24906,N_24794);
and U25090 (N_25090,N_24924,N_24891);
or U25091 (N_25091,N_24786,N_24824);
xnor U25092 (N_25092,N_24920,N_24904);
nor U25093 (N_25093,N_24825,N_24952);
and U25094 (N_25094,N_24765,N_24889);
or U25095 (N_25095,N_24855,N_24844);
xnor U25096 (N_25096,N_24753,N_24881);
and U25097 (N_25097,N_24767,N_24886);
nand U25098 (N_25098,N_24833,N_24890);
nor U25099 (N_25099,N_24876,N_24790);
and U25100 (N_25100,N_24829,N_24784);
nor U25101 (N_25101,N_24998,N_24761);
and U25102 (N_25102,N_24965,N_24879);
xnor U25103 (N_25103,N_24980,N_24884);
xnor U25104 (N_25104,N_24776,N_24866);
xnor U25105 (N_25105,N_24764,N_24842);
nor U25106 (N_25106,N_24921,N_24999);
and U25107 (N_25107,N_24915,N_24795);
nor U25108 (N_25108,N_24937,N_24901);
nand U25109 (N_25109,N_24947,N_24815);
and U25110 (N_25110,N_24809,N_24887);
nor U25111 (N_25111,N_24905,N_24968);
xor U25112 (N_25112,N_24841,N_24801);
or U25113 (N_25113,N_24961,N_24941);
or U25114 (N_25114,N_24988,N_24951);
nor U25115 (N_25115,N_24989,N_24791);
nand U25116 (N_25116,N_24813,N_24796);
or U25117 (N_25117,N_24787,N_24994);
and U25118 (N_25118,N_24834,N_24991);
and U25119 (N_25119,N_24907,N_24985);
nand U25120 (N_25120,N_24996,N_24912);
xor U25121 (N_25121,N_24962,N_24900);
nand U25122 (N_25122,N_24875,N_24918);
or U25123 (N_25123,N_24754,N_24758);
nand U25124 (N_25124,N_24768,N_24870);
and U25125 (N_25125,N_24966,N_24894);
nand U25126 (N_25126,N_24808,N_24927);
nor U25127 (N_25127,N_24948,N_24804);
and U25128 (N_25128,N_24840,N_24844);
or U25129 (N_25129,N_24865,N_24879);
nand U25130 (N_25130,N_24799,N_24920);
or U25131 (N_25131,N_24780,N_24961);
or U25132 (N_25132,N_24822,N_24868);
or U25133 (N_25133,N_24802,N_24878);
and U25134 (N_25134,N_24986,N_24930);
or U25135 (N_25135,N_24902,N_24880);
nand U25136 (N_25136,N_24921,N_24953);
nor U25137 (N_25137,N_24935,N_24753);
nand U25138 (N_25138,N_24903,N_24930);
nand U25139 (N_25139,N_24863,N_24774);
nand U25140 (N_25140,N_24931,N_24767);
xnor U25141 (N_25141,N_24898,N_24991);
xnor U25142 (N_25142,N_24860,N_24979);
xnor U25143 (N_25143,N_24936,N_24974);
xnor U25144 (N_25144,N_24867,N_24785);
or U25145 (N_25145,N_24919,N_24875);
xnor U25146 (N_25146,N_24965,N_24795);
or U25147 (N_25147,N_24987,N_24992);
xnor U25148 (N_25148,N_24842,N_24893);
or U25149 (N_25149,N_24802,N_24801);
or U25150 (N_25150,N_24981,N_24889);
nand U25151 (N_25151,N_24905,N_24806);
or U25152 (N_25152,N_24992,N_24919);
and U25153 (N_25153,N_24920,N_24780);
or U25154 (N_25154,N_24915,N_24919);
nor U25155 (N_25155,N_24953,N_24779);
xnor U25156 (N_25156,N_24807,N_24816);
and U25157 (N_25157,N_24761,N_24943);
nand U25158 (N_25158,N_24866,N_24843);
nand U25159 (N_25159,N_24753,N_24988);
nand U25160 (N_25160,N_24891,N_24810);
or U25161 (N_25161,N_24834,N_24875);
nor U25162 (N_25162,N_24923,N_24902);
or U25163 (N_25163,N_24984,N_24838);
nand U25164 (N_25164,N_24765,N_24949);
xor U25165 (N_25165,N_24953,N_24897);
and U25166 (N_25166,N_24959,N_24817);
nor U25167 (N_25167,N_24869,N_24981);
nor U25168 (N_25168,N_24804,N_24869);
nor U25169 (N_25169,N_24859,N_24908);
and U25170 (N_25170,N_24955,N_24899);
nor U25171 (N_25171,N_24951,N_24795);
xor U25172 (N_25172,N_24961,N_24765);
and U25173 (N_25173,N_24971,N_24809);
nor U25174 (N_25174,N_24879,N_24863);
nand U25175 (N_25175,N_24810,N_24856);
nor U25176 (N_25176,N_24882,N_24765);
and U25177 (N_25177,N_24857,N_24843);
or U25178 (N_25178,N_24867,N_24874);
nor U25179 (N_25179,N_24946,N_24815);
xor U25180 (N_25180,N_24761,N_24804);
nand U25181 (N_25181,N_24780,N_24791);
nand U25182 (N_25182,N_24997,N_24929);
nor U25183 (N_25183,N_24918,N_24887);
xnor U25184 (N_25184,N_24877,N_24861);
or U25185 (N_25185,N_24922,N_24825);
xor U25186 (N_25186,N_24887,N_24986);
xnor U25187 (N_25187,N_24826,N_24790);
and U25188 (N_25188,N_24977,N_24792);
or U25189 (N_25189,N_24776,N_24845);
nand U25190 (N_25190,N_24957,N_24965);
and U25191 (N_25191,N_24974,N_24904);
xnor U25192 (N_25192,N_24915,N_24889);
nand U25193 (N_25193,N_24996,N_24864);
and U25194 (N_25194,N_24960,N_24884);
or U25195 (N_25195,N_24890,N_24773);
nand U25196 (N_25196,N_24816,N_24815);
xnor U25197 (N_25197,N_24763,N_24751);
xnor U25198 (N_25198,N_24823,N_24856);
xor U25199 (N_25199,N_24970,N_24923);
nor U25200 (N_25200,N_24792,N_24810);
or U25201 (N_25201,N_24762,N_24861);
and U25202 (N_25202,N_24818,N_24761);
xnor U25203 (N_25203,N_24787,N_24856);
and U25204 (N_25204,N_24828,N_24760);
nor U25205 (N_25205,N_24962,N_24976);
or U25206 (N_25206,N_24855,N_24824);
xor U25207 (N_25207,N_24935,N_24949);
nand U25208 (N_25208,N_24917,N_24964);
xnor U25209 (N_25209,N_24751,N_24753);
nand U25210 (N_25210,N_24833,N_24962);
xor U25211 (N_25211,N_24954,N_24788);
nor U25212 (N_25212,N_24933,N_24981);
xor U25213 (N_25213,N_24938,N_24960);
nand U25214 (N_25214,N_24893,N_24983);
or U25215 (N_25215,N_24755,N_24955);
nor U25216 (N_25216,N_24783,N_24954);
nand U25217 (N_25217,N_24958,N_24920);
or U25218 (N_25218,N_24971,N_24896);
xor U25219 (N_25219,N_24973,N_24952);
and U25220 (N_25220,N_24844,N_24766);
or U25221 (N_25221,N_24796,N_24937);
xor U25222 (N_25222,N_24930,N_24896);
nor U25223 (N_25223,N_24919,N_24899);
xor U25224 (N_25224,N_24877,N_24823);
nor U25225 (N_25225,N_24936,N_24862);
nor U25226 (N_25226,N_24789,N_24804);
nand U25227 (N_25227,N_24895,N_24994);
xor U25228 (N_25228,N_24967,N_24942);
and U25229 (N_25229,N_24825,N_24767);
xnor U25230 (N_25230,N_24778,N_24843);
xor U25231 (N_25231,N_24942,N_24798);
nor U25232 (N_25232,N_24901,N_24917);
and U25233 (N_25233,N_24981,N_24943);
nor U25234 (N_25234,N_24868,N_24920);
nand U25235 (N_25235,N_24998,N_24800);
nand U25236 (N_25236,N_24819,N_24917);
or U25237 (N_25237,N_24995,N_24797);
or U25238 (N_25238,N_24845,N_24848);
nor U25239 (N_25239,N_24908,N_24973);
or U25240 (N_25240,N_24771,N_24910);
and U25241 (N_25241,N_24889,N_24898);
xor U25242 (N_25242,N_24761,N_24893);
xnor U25243 (N_25243,N_24899,N_24799);
xor U25244 (N_25244,N_24763,N_24993);
nor U25245 (N_25245,N_24887,N_24770);
xor U25246 (N_25246,N_24951,N_24913);
nand U25247 (N_25247,N_24980,N_24894);
nand U25248 (N_25248,N_24857,N_24996);
and U25249 (N_25249,N_24896,N_24910);
xnor U25250 (N_25250,N_25057,N_25146);
nor U25251 (N_25251,N_25204,N_25189);
xor U25252 (N_25252,N_25173,N_25177);
nor U25253 (N_25253,N_25107,N_25078);
or U25254 (N_25254,N_25128,N_25133);
or U25255 (N_25255,N_25009,N_25161);
nand U25256 (N_25256,N_25164,N_25096);
nand U25257 (N_25257,N_25007,N_25059);
nand U25258 (N_25258,N_25222,N_25139);
nor U25259 (N_25259,N_25051,N_25241);
nand U25260 (N_25260,N_25150,N_25236);
and U25261 (N_25261,N_25027,N_25171);
nor U25262 (N_25262,N_25235,N_25145);
and U25263 (N_25263,N_25246,N_25207);
nor U25264 (N_25264,N_25187,N_25157);
xnor U25265 (N_25265,N_25101,N_25125);
nor U25266 (N_25266,N_25024,N_25152);
nor U25267 (N_25267,N_25242,N_25072);
nor U25268 (N_25268,N_25182,N_25217);
or U25269 (N_25269,N_25114,N_25028);
nand U25270 (N_25270,N_25109,N_25071);
xnor U25271 (N_25271,N_25010,N_25126);
nor U25272 (N_25272,N_25120,N_25215);
or U25273 (N_25273,N_25084,N_25111);
nor U25274 (N_25274,N_25122,N_25248);
or U25275 (N_25275,N_25046,N_25158);
nand U25276 (N_25276,N_25023,N_25208);
nor U25277 (N_25277,N_25240,N_25226);
nor U25278 (N_25278,N_25165,N_25121);
nand U25279 (N_25279,N_25004,N_25201);
and U25280 (N_25280,N_25013,N_25117);
or U25281 (N_25281,N_25003,N_25202);
or U25282 (N_25282,N_25079,N_25091);
or U25283 (N_25283,N_25154,N_25233);
nor U25284 (N_25284,N_25025,N_25063);
nor U25285 (N_25285,N_25210,N_25098);
and U25286 (N_25286,N_25016,N_25088);
xnor U25287 (N_25287,N_25223,N_25232);
or U25288 (N_25288,N_25090,N_25034);
nor U25289 (N_25289,N_25245,N_25019);
nor U25290 (N_25290,N_25001,N_25155);
or U25291 (N_25291,N_25018,N_25080);
nor U25292 (N_25292,N_25069,N_25216);
or U25293 (N_25293,N_25219,N_25149);
xnor U25294 (N_25294,N_25190,N_25032);
or U25295 (N_25295,N_25144,N_25082);
and U25296 (N_25296,N_25138,N_25188);
and U25297 (N_25297,N_25002,N_25026);
xor U25298 (N_25298,N_25230,N_25218);
and U25299 (N_25299,N_25148,N_25200);
nor U25300 (N_25300,N_25085,N_25163);
or U25301 (N_25301,N_25053,N_25108);
nor U25302 (N_25302,N_25067,N_25213);
and U25303 (N_25303,N_25102,N_25172);
or U25304 (N_25304,N_25045,N_25074);
or U25305 (N_25305,N_25168,N_25129);
nand U25306 (N_25306,N_25214,N_25176);
and U25307 (N_25307,N_25017,N_25075);
nand U25308 (N_25308,N_25127,N_25021);
and U25309 (N_25309,N_25175,N_25183);
nor U25310 (N_25310,N_25156,N_25185);
xnor U25311 (N_25311,N_25064,N_25077);
nor U25312 (N_25312,N_25060,N_25008);
nor U25313 (N_25313,N_25151,N_25056);
xnor U25314 (N_25314,N_25020,N_25143);
nor U25315 (N_25315,N_25170,N_25211);
xor U25316 (N_25316,N_25100,N_25159);
xor U25317 (N_25317,N_25011,N_25012);
or U25318 (N_25318,N_25179,N_25162);
and U25319 (N_25319,N_25052,N_25036);
nand U25320 (N_25320,N_25030,N_25061);
nor U25321 (N_25321,N_25099,N_25224);
and U25322 (N_25322,N_25244,N_25000);
nor U25323 (N_25323,N_25199,N_25054);
nand U25324 (N_25324,N_25086,N_25195);
xnor U25325 (N_25325,N_25206,N_25174);
xor U25326 (N_25326,N_25227,N_25035);
nor U25327 (N_25327,N_25105,N_25137);
nand U25328 (N_25328,N_25033,N_25073);
nor U25329 (N_25329,N_25039,N_25153);
xor U25330 (N_25330,N_25049,N_25197);
nor U25331 (N_25331,N_25065,N_25167);
and U25332 (N_25332,N_25238,N_25134);
nand U25333 (N_25333,N_25043,N_25089);
and U25334 (N_25334,N_25135,N_25247);
nor U25335 (N_25335,N_25076,N_25212);
nand U25336 (N_25336,N_25234,N_25180);
or U25337 (N_25337,N_25198,N_25106);
nor U25338 (N_25338,N_25022,N_25066);
nor U25339 (N_25339,N_25047,N_25070);
nor U25340 (N_25340,N_25239,N_25040);
nand U25341 (N_25341,N_25140,N_25147);
or U25342 (N_25342,N_25087,N_25115);
nand U25343 (N_25343,N_25042,N_25194);
or U25344 (N_25344,N_25130,N_25103);
nand U25345 (N_25345,N_25029,N_25123);
or U25346 (N_25346,N_25092,N_25237);
nor U25347 (N_25347,N_25094,N_25229);
and U25348 (N_25348,N_25005,N_25184);
or U25349 (N_25349,N_25132,N_25015);
or U25350 (N_25350,N_25249,N_25178);
xnor U25351 (N_25351,N_25044,N_25231);
or U25352 (N_25352,N_25062,N_25209);
xnor U25353 (N_25353,N_25136,N_25118);
or U25354 (N_25354,N_25031,N_25131);
xnor U25355 (N_25355,N_25097,N_25083);
xnor U25356 (N_25356,N_25014,N_25095);
and U25357 (N_25357,N_25058,N_25110);
nand U25358 (N_25358,N_25191,N_25196);
and U25359 (N_25359,N_25166,N_25124);
nand U25360 (N_25360,N_25055,N_25142);
or U25361 (N_25361,N_25228,N_25193);
xnor U25362 (N_25362,N_25116,N_25041);
nand U25363 (N_25363,N_25038,N_25243);
or U25364 (N_25364,N_25081,N_25037);
xor U25365 (N_25365,N_25169,N_25141);
nor U25366 (N_25366,N_25050,N_25203);
nor U25367 (N_25367,N_25093,N_25068);
or U25368 (N_25368,N_25221,N_25220);
xor U25369 (N_25369,N_25225,N_25113);
nor U25370 (N_25370,N_25112,N_25192);
or U25371 (N_25371,N_25119,N_25104);
or U25372 (N_25372,N_25205,N_25160);
nand U25373 (N_25373,N_25048,N_25006);
and U25374 (N_25374,N_25186,N_25181);
xor U25375 (N_25375,N_25071,N_25248);
or U25376 (N_25376,N_25202,N_25133);
nor U25377 (N_25377,N_25242,N_25011);
nand U25378 (N_25378,N_25215,N_25114);
and U25379 (N_25379,N_25069,N_25140);
nand U25380 (N_25380,N_25073,N_25091);
xor U25381 (N_25381,N_25064,N_25089);
nor U25382 (N_25382,N_25121,N_25111);
nand U25383 (N_25383,N_25237,N_25141);
or U25384 (N_25384,N_25045,N_25141);
or U25385 (N_25385,N_25175,N_25160);
xnor U25386 (N_25386,N_25135,N_25073);
or U25387 (N_25387,N_25028,N_25086);
or U25388 (N_25388,N_25102,N_25162);
nor U25389 (N_25389,N_25074,N_25208);
and U25390 (N_25390,N_25035,N_25210);
and U25391 (N_25391,N_25124,N_25207);
nor U25392 (N_25392,N_25114,N_25057);
and U25393 (N_25393,N_25165,N_25033);
or U25394 (N_25394,N_25094,N_25062);
xor U25395 (N_25395,N_25105,N_25178);
nand U25396 (N_25396,N_25234,N_25203);
or U25397 (N_25397,N_25115,N_25057);
nand U25398 (N_25398,N_25027,N_25202);
and U25399 (N_25399,N_25088,N_25202);
xnor U25400 (N_25400,N_25012,N_25244);
xnor U25401 (N_25401,N_25244,N_25225);
nand U25402 (N_25402,N_25224,N_25112);
nor U25403 (N_25403,N_25088,N_25177);
xnor U25404 (N_25404,N_25121,N_25025);
xor U25405 (N_25405,N_25101,N_25017);
nand U25406 (N_25406,N_25042,N_25050);
nor U25407 (N_25407,N_25235,N_25080);
nand U25408 (N_25408,N_25228,N_25004);
and U25409 (N_25409,N_25063,N_25109);
and U25410 (N_25410,N_25133,N_25225);
nor U25411 (N_25411,N_25073,N_25216);
xor U25412 (N_25412,N_25199,N_25187);
and U25413 (N_25413,N_25078,N_25212);
nand U25414 (N_25414,N_25029,N_25100);
nand U25415 (N_25415,N_25083,N_25248);
xnor U25416 (N_25416,N_25241,N_25064);
and U25417 (N_25417,N_25248,N_25060);
nor U25418 (N_25418,N_25121,N_25234);
and U25419 (N_25419,N_25242,N_25082);
xnor U25420 (N_25420,N_25228,N_25147);
nor U25421 (N_25421,N_25136,N_25032);
or U25422 (N_25422,N_25192,N_25096);
or U25423 (N_25423,N_25118,N_25180);
xor U25424 (N_25424,N_25126,N_25072);
nor U25425 (N_25425,N_25202,N_25012);
nand U25426 (N_25426,N_25131,N_25054);
nor U25427 (N_25427,N_25063,N_25022);
nor U25428 (N_25428,N_25080,N_25147);
or U25429 (N_25429,N_25112,N_25078);
nor U25430 (N_25430,N_25019,N_25142);
nor U25431 (N_25431,N_25026,N_25217);
xor U25432 (N_25432,N_25225,N_25085);
nor U25433 (N_25433,N_25128,N_25032);
and U25434 (N_25434,N_25037,N_25202);
nor U25435 (N_25435,N_25023,N_25016);
nor U25436 (N_25436,N_25132,N_25190);
nor U25437 (N_25437,N_25159,N_25228);
nor U25438 (N_25438,N_25127,N_25113);
and U25439 (N_25439,N_25040,N_25117);
nor U25440 (N_25440,N_25002,N_25203);
nor U25441 (N_25441,N_25004,N_25098);
and U25442 (N_25442,N_25056,N_25177);
nand U25443 (N_25443,N_25137,N_25031);
nor U25444 (N_25444,N_25049,N_25043);
or U25445 (N_25445,N_25102,N_25030);
xor U25446 (N_25446,N_25190,N_25044);
nand U25447 (N_25447,N_25121,N_25182);
and U25448 (N_25448,N_25236,N_25174);
nand U25449 (N_25449,N_25075,N_25214);
xor U25450 (N_25450,N_25125,N_25010);
nor U25451 (N_25451,N_25180,N_25164);
and U25452 (N_25452,N_25049,N_25201);
and U25453 (N_25453,N_25082,N_25157);
nand U25454 (N_25454,N_25223,N_25156);
nor U25455 (N_25455,N_25200,N_25093);
nor U25456 (N_25456,N_25150,N_25144);
nand U25457 (N_25457,N_25090,N_25202);
xnor U25458 (N_25458,N_25054,N_25112);
nor U25459 (N_25459,N_25036,N_25176);
nor U25460 (N_25460,N_25132,N_25129);
nand U25461 (N_25461,N_25010,N_25177);
xnor U25462 (N_25462,N_25160,N_25035);
nor U25463 (N_25463,N_25107,N_25075);
xnor U25464 (N_25464,N_25005,N_25057);
and U25465 (N_25465,N_25122,N_25128);
nor U25466 (N_25466,N_25020,N_25099);
or U25467 (N_25467,N_25081,N_25247);
nor U25468 (N_25468,N_25197,N_25134);
xnor U25469 (N_25469,N_25035,N_25169);
and U25470 (N_25470,N_25100,N_25074);
nor U25471 (N_25471,N_25151,N_25064);
xor U25472 (N_25472,N_25242,N_25042);
nand U25473 (N_25473,N_25208,N_25035);
or U25474 (N_25474,N_25131,N_25142);
or U25475 (N_25475,N_25087,N_25188);
nor U25476 (N_25476,N_25031,N_25165);
nor U25477 (N_25477,N_25095,N_25059);
xnor U25478 (N_25478,N_25030,N_25212);
and U25479 (N_25479,N_25061,N_25141);
and U25480 (N_25480,N_25079,N_25186);
and U25481 (N_25481,N_25118,N_25203);
xnor U25482 (N_25482,N_25167,N_25032);
nor U25483 (N_25483,N_25026,N_25145);
nor U25484 (N_25484,N_25200,N_25018);
or U25485 (N_25485,N_25079,N_25156);
nor U25486 (N_25486,N_25195,N_25194);
nand U25487 (N_25487,N_25031,N_25243);
or U25488 (N_25488,N_25121,N_25051);
nor U25489 (N_25489,N_25110,N_25180);
nand U25490 (N_25490,N_25044,N_25083);
nand U25491 (N_25491,N_25160,N_25235);
nor U25492 (N_25492,N_25226,N_25134);
nor U25493 (N_25493,N_25059,N_25188);
and U25494 (N_25494,N_25157,N_25147);
or U25495 (N_25495,N_25201,N_25110);
nand U25496 (N_25496,N_25102,N_25129);
and U25497 (N_25497,N_25092,N_25178);
nor U25498 (N_25498,N_25053,N_25054);
nor U25499 (N_25499,N_25128,N_25211);
nand U25500 (N_25500,N_25294,N_25469);
and U25501 (N_25501,N_25372,N_25406);
or U25502 (N_25502,N_25475,N_25359);
xnor U25503 (N_25503,N_25340,N_25276);
or U25504 (N_25504,N_25396,N_25362);
or U25505 (N_25505,N_25354,N_25456);
or U25506 (N_25506,N_25379,N_25483);
and U25507 (N_25507,N_25336,N_25348);
xor U25508 (N_25508,N_25452,N_25443);
nor U25509 (N_25509,N_25433,N_25314);
and U25510 (N_25510,N_25446,N_25395);
or U25511 (N_25511,N_25489,N_25338);
nand U25512 (N_25512,N_25450,N_25417);
xor U25513 (N_25513,N_25335,N_25384);
nor U25514 (N_25514,N_25327,N_25284);
nor U25515 (N_25515,N_25312,N_25451);
and U25516 (N_25516,N_25289,N_25437);
or U25517 (N_25517,N_25495,N_25304);
and U25518 (N_25518,N_25321,N_25325);
xnor U25519 (N_25519,N_25411,N_25371);
nor U25520 (N_25520,N_25316,N_25268);
or U25521 (N_25521,N_25346,N_25322);
nor U25522 (N_25522,N_25301,N_25264);
nor U25523 (N_25523,N_25271,N_25458);
xnor U25524 (N_25524,N_25415,N_25375);
nor U25525 (N_25525,N_25465,N_25389);
or U25526 (N_25526,N_25370,N_25470);
xor U25527 (N_25527,N_25329,N_25493);
or U25528 (N_25528,N_25390,N_25453);
or U25529 (N_25529,N_25377,N_25297);
nor U25530 (N_25530,N_25461,N_25420);
and U25531 (N_25531,N_25445,N_25353);
nand U25532 (N_25532,N_25455,N_25488);
xnor U25533 (N_25533,N_25324,N_25449);
or U25534 (N_25534,N_25290,N_25333);
xnor U25535 (N_25535,N_25405,N_25293);
or U25536 (N_25536,N_25430,N_25317);
nand U25537 (N_25537,N_25360,N_25341);
or U25538 (N_25538,N_25376,N_25299);
or U25539 (N_25539,N_25288,N_25291);
xnor U25540 (N_25540,N_25496,N_25349);
or U25541 (N_25541,N_25302,N_25410);
and U25542 (N_25542,N_25497,N_25432);
or U25543 (N_25543,N_25463,N_25356);
and U25544 (N_25544,N_25295,N_25344);
nand U25545 (N_25545,N_25318,N_25482);
or U25546 (N_25546,N_25421,N_25459);
or U25547 (N_25547,N_25454,N_25266);
or U25548 (N_25548,N_25412,N_25478);
xnor U25549 (N_25549,N_25251,N_25498);
xor U25550 (N_25550,N_25391,N_25457);
or U25551 (N_25551,N_25323,N_25388);
nand U25552 (N_25552,N_25307,N_25416);
or U25553 (N_25553,N_25479,N_25466);
or U25554 (N_25554,N_25260,N_25380);
or U25555 (N_25555,N_25343,N_25368);
nand U25556 (N_25556,N_25448,N_25355);
and U25557 (N_25557,N_25259,N_25279);
nand U25558 (N_25558,N_25403,N_25485);
nand U25559 (N_25559,N_25331,N_25392);
and U25560 (N_25560,N_25490,N_25278);
or U25561 (N_25561,N_25369,N_25422);
or U25562 (N_25562,N_25480,N_25434);
or U25563 (N_25563,N_25427,N_25309);
and U25564 (N_25564,N_25281,N_25319);
or U25565 (N_25565,N_25444,N_25352);
nand U25566 (N_25566,N_25270,N_25441);
and U25567 (N_25567,N_25471,N_25409);
and U25568 (N_25568,N_25460,N_25287);
nor U25569 (N_25569,N_25298,N_25313);
and U25570 (N_25570,N_25413,N_25258);
nor U25571 (N_25571,N_25467,N_25252);
nor U25572 (N_25572,N_25358,N_25428);
nand U25573 (N_25573,N_25419,N_25499);
nand U25574 (N_25574,N_25363,N_25387);
or U25575 (N_25575,N_25261,N_25339);
nor U25576 (N_25576,N_25397,N_25404);
xor U25577 (N_25577,N_25275,N_25274);
xor U25578 (N_25578,N_25292,N_25254);
and U25579 (N_25579,N_25486,N_25267);
nor U25580 (N_25580,N_25357,N_25350);
nand U25581 (N_25581,N_25378,N_25367);
nand U25582 (N_25582,N_25386,N_25381);
nor U25583 (N_25583,N_25364,N_25337);
or U25584 (N_25584,N_25347,N_25382);
nor U25585 (N_25585,N_25481,N_25474);
nand U25586 (N_25586,N_25402,N_25425);
and U25587 (N_25587,N_25345,N_25351);
xnor U25588 (N_25588,N_25334,N_25280);
and U25589 (N_25589,N_25286,N_25426);
nor U25590 (N_25590,N_25383,N_25408);
or U25591 (N_25591,N_25414,N_25300);
or U25592 (N_25592,N_25435,N_25436);
and U25593 (N_25593,N_25257,N_25310);
nor U25594 (N_25594,N_25431,N_25255);
nand U25595 (N_25595,N_25262,N_25423);
nand U25596 (N_25596,N_25285,N_25462);
nand U25597 (N_25597,N_25418,N_25365);
or U25598 (N_25598,N_25468,N_25308);
nor U25599 (N_25599,N_25429,N_25473);
xnor U25600 (N_25600,N_25311,N_25494);
nand U25601 (N_25601,N_25447,N_25442);
xor U25602 (N_25602,N_25272,N_25328);
and U25603 (N_25603,N_25283,N_25477);
and U25604 (N_25604,N_25464,N_25424);
nor U25605 (N_25605,N_25373,N_25374);
nand U25606 (N_25606,N_25282,N_25439);
and U25607 (N_25607,N_25401,N_25305);
nor U25608 (N_25608,N_25326,N_25263);
or U25609 (N_25609,N_25393,N_25250);
nor U25610 (N_25610,N_25277,N_25342);
or U25611 (N_25611,N_25487,N_25273);
xnor U25612 (N_25612,N_25492,N_25491);
nor U25613 (N_25613,N_25361,N_25315);
nand U25614 (N_25614,N_25407,N_25400);
and U25615 (N_25615,N_25265,N_25385);
or U25616 (N_25616,N_25366,N_25332);
nor U25617 (N_25617,N_25438,N_25330);
and U25618 (N_25618,N_25472,N_25399);
and U25619 (N_25619,N_25394,N_25306);
or U25620 (N_25620,N_25398,N_25476);
xnor U25621 (N_25621,N_25296,N_25256);
and U25622 (N_25622,N_25303,N_25269);
or U25623 (N_25623,N_25253,N_25440);
nand U25624 (N_25624,N_25320,N_25484);
and U25625 (N_25625,N_25471,N_25278);
xnor U25626 (N_25626,N_25357,N_25472);
xor U25627 (N_25627,N_25484,N_25455);
nand U25628 (N_25628,N_25366,N_25324);
or U25629 (N_25629,N_25397,N_25333);
or U25630 (N_25630,N_25463,N_25451);
and U25631 (N_25631,N_25433,N_25459);
xor U25632 (N_25632,N_25411,N_25424);
nor U25633 (N_25633,N_25299,N_25426);
or U25634 (N_25634,N_25407,N_25460);
nor U25635 (N_25635,N_25343,N_25370);
nand U25636 (N_25636,N_25267,N_25284);
or U25637 (N_25637,N_25317,N_25473);
and U25638 (N_25638,N_25324,N_25271);
or U25639 (N_25639,N_25382,N_25493);
nor U25640 (N_25640,N_25445,N_25264);
xnor U25641 (N_25641,N_25350,N_25457);
and U25642 (N_25642,N_25498,N_25383);
or U25643 (N_25643,N_25299,N_25269);
and U25644 (N_25644,N_25333,N_25302);
and U25645 (N_25645,N_25304,N_25370);
nand U25646 (N_25646,N_25415,N_25385);
or U25647 (N_25647,N_25252,N_25424);
nor U25648 (N_25648,N_25367,N_25452);
nor U25649 (N_25649,N_25424,N_25339);
and U25650 (N_25650,N_25356,N_25471);
xor U25651 (N_25651,N_25467,N_25403);
and U25652 (N_25652,N_25450,N_25299);
or U25653 (N_25653,N_25413,N_25294);
or U25654 (N_25654,N_25305,N_25429);
or U25655 (N_25655,N_25270,N_25357);
or U25656 (N_25656,N_25309,N_25406);
and U25657 (N_25657,N_25438,N_25421);
or U25658 (N_25658,N_25432,N_25266);
nand U25659 (N_25659,N_25380,N_25282);
nor U25660 (N_25660,N_25384,N_25388);
nor U25661 (N_25661,N_25297,N_25386);
and U25662 (N_25662,N_25379,N_25253);
xnor U25663 (N_25663,N_25485,N_25323);
or U25664 (N_25664,N_25326,N_25450);
nor U25665 (N_25665,N_25410,N_25436);
nand U25666 (N_25666,N_25283,N_25262);
and U25667 (N_25667,N_25291,N_25345);
and U25668 (N_25668,N_25314,N_25323);
or U25669 (N_25669,N_25344,N_25322);
xor U25670 (N_25670,N_25357,N_25449);
nor U25671 (N_25671,N_25303,N_25474);
nand U25672 (N_25672,N_25343,N_25287);
nand U25673 (N_25673,N_25417,N_25444);
nor U25674 (N_25674,N_25365,N_25399);
or U25675 (N_25675,N_25440,N_25252);
nand U25676 (N_25676,N_25452,N_25402);
nor U25677 (N_25677,N_25350,N_25342);
nand U25678 (N_25678,N_25253,N_25358);
nor U25679 (N_25679,N_25410,N_25411);
or U25680 (N_25680,N_25262,N_25418);
xor U25681 (N_25681,N_25499,N_25425);
and U25682 (N_25682,N_25305,N_25477);
nor U25683 (N_25683,N_25256,N_25274);
nand U25684 (N_25684,N_25323,N_25316);
xnor U25685 (N_25685,N_25304,N_25316);
or U25686 (N_25686,N_25365,N_25298);
nor U25687 (N_25687,N_25482,N_25349);
nor U25688 (N_25688,N_25447,N_25499);
nor U25689 (N_25689,N_25277,N_25410);
nand U25690 (N_25690,N_25361,N_25456);
nor U25691 (N_25691,N_25333,N_25426);
xnor U25692 (N_25692,N_25449,N_25416);
or U25693 (N_25693,N_25320,N_25494);
nand U25694 (N_25694,N_25494,N_25331);
xnor U25695 (N_25695,N_25406,N_25485);
or U25696 (N_25696,N_25424,N_25297);
or U25697 (N_25697,N_25358,N_25448);
nor U25698 (N_25698,N_25491,N_25459);
xor U25699 (N_25699,N_25364,N_25391);
xnor U25700 (N_25700,N_25308,N_25268);
and U25701 (N_25701,N_25273,N_25410);
and U25702 (N_25702,N_25312,N_25399);
nor U25703 (N_25703,N_25441,N_25297);
nor U25704 (N_25704,N_25454,N_25250);
or U25705 (N_25705,N_25263,N_25281);
xor U25706 (N_25706,N_25325,N_25256);
nand U25707 (N_25707,N_25447,N_25395);
xor U25708 (N_25708,N_25281,N_25265);
or U25709 (N_25709,N_25375,N_25442);
xnor U25710 (N_25710,N_25346,N_25435);
nor U25711 (N_25711,N_25327,N_25307);
and U25712 (N_25712,N_25275,N_25318);
nor U25713 (N_25713,N_25251,N_25311);
or U25714 (N_25714,N_25346,N_25395);
nor U25715 (N_25715,N_25284,N_25352);
or U25716 (N_25716,N_25433,N_25404);
nand U25717 (N_25717,N_25313,N_25441);
xnor U25718 (N_25718,N_25412,N_25291);
xor U25719 (N_25719,N_25312,N_25460);
xnor U25720 (N_25720,N_25422,N_25328);
or U25721 (N_25721,N_25363,N_25464);
and U25722 (N_25722,N_25476,N_25496);
nor U25723 (N_25723,N_25262,N_25472);
nand U25724 (N_25724,N_25441,N_25404);
nand U25725 (N_25725,N_25386,N_25424);
nand U25726 (N_25726,N_25331,N_25321);
or U25727 (N_25727,N_25383,N_25421);
xnor U25728 (N_25728,N_25363,N_25444);
and U25729 (N_25729,N_25264,N_25374);
nand U25730 (N_25730,N_25257,N_25420);
and U25731 (N_25731,N_25309,N_25294);
nand U25732 (N_25732,N_25267,N_25279);
and U25733 (N_25733,N_25336,N_25486);
nand U25734 (N_25734,N_25486,N_25335);
and U25735 (N_25735,N_25291,N_25459);
and U25736 (N_25736,N_25281,N_25361);
nor U25737 (N_25737,N_25341,N_25398);
or U25738 (N_25738,N_25450,N_25436);
nor U25739 (N_25739,N_25410,N_25308);
and U25740 (N_25740,N_25430,N_25432);
nand U25741 (N_25741,N_25457,N_25261);
nand U25742 (N_25742,N_25455,N_25285);
nor U25743 (N_25743,N_25303,N_25329);
nor U25744 (N_25744,N_25366,N_25405);
xor U25745 (N_25745,N_25498,N_25404);
or U25746 (N_25746,N_25293,N_25374);
nor U25747 (N_25747,N_25416,N_25331);
xnor U25748 (N_25748,N_25433,N_25484);
nand U25749 (N_25749,N_25381,N_25338);
nor U25750 (N_25750,N_25741,N_25668);
and U25751 (N_25751,N_25579,N_25658);
nand U25752 (N_25752,N_25719,N_25709);
or U25753 (N_25753,N_25550,N_25647);
xor U25754 (N_25754,N_25586,N_25514);
nand U25755 (N_25755,N_25555,N_25618);
xor U25756 (N_25756,N_25643,N_25602);
nand U25757 (N_25757,N_25612,N_25540);
nand U25758 (N_25758,N_25530,N_25508);
nand U25759 (N_25759,N_25687,N_25721);
or U25760 (N_25760,N_25746,N_25608);
nand U25761 (N_25761,N_25718,N_25609);
or U25762 (N_25762,N_25605,N_25717);
nor U25763 (N_25763,N_25676,N_25636);
xor U25764 (N_25764,N_25626,N_25648);
and U25765 (N_25765,N_25696,N_25597);
or U25766 (N_25766,N_25716,N_25500);
nand U25767 (N_25767,N_25679,N_25673);
nand U25768 (N_25768,N_25567,N_25532);
and U25769 (N_25769,N_25659,N_25544);
or U25770 (N_25770,N_25526,N_25691);
and U25771 (N_25771,N_25733,N_25584);
and U25772 (N_25772,N_25683,N_25685);
xor U25773 (N_25773,N_25649,N_25727);
or U25774 (N_25774,N_25537,N_25601);
xor U25775 (N_25775,N_25698,N_25507);
xor U25776 (N_25776,N_25592,N_25682);
and U25777 (N_25777,N_25724,N_25552);
and U25778 (N_25778,N_25638,N_25703);
nand U25779 (N_25779,N_25599,N_25681);
nor U25780 (N_25780,N_25661,N_25501);
or U25781 (N_25781,N_25695,N_25688);
and U25782 (N_25782,N_25726,N_25651);
nand U25783 (N_25783,N_25670,N_25705);
xnor U25784 (N_25784,N_25669,N_25723);
and U25785 (N_25785,N_25725,N_25512);
xor U25786 (N_25786,N_25556,N_25631);
and U25787 (N_25787,N_25564,N_25606);
or U25788 (N_25788,N_25619,N_25642);
nand U25789 (N_25789,N_25667,N_25672);
and U25790 (N_25790,N_25522,N_25662);
nor U25791 (N_25791,N_25557,N_25577);
nor U25792 (N_25792,N_25694,N_25546);
nor U25793 (N_25793,N_25737,N_25749);
nand U25794 (N_25794,N_25699,N_25735);
or U25795 (N_25795,N_25657,N_25663);
nand U25796 (N_25796,N_25632,N_25607);
and U25797 (N_25797,N_25553,N_25732);
nor U25798 (N_25798,N_25536,N_25736);
nand U25799 (N_25799,N_25713,N_25692);
xor U25800 (N_25800,N_25538,N_25678);
nor U25801 (N_25801,N_25534,N_25562);
nand U25802 (N_25802,N_25574,N_25640);
and U25803 (N_25803,N_25547,N_25585);
nand U25804 (N_25804,N_25671,N_25548);
and U25805 (N_25805,N_25588,N_25656);
nor U25806 (N_25806,N_25639,N_25622);
and U25807 (N_25807,N_25518,N_25533);
nor U25808 (N_25808,N_25589,N_25702);
and U25809 (N_25809,N_25653,N_25519);
and U25810 (N_25810,N_25571,N_25520);
or U25811 (N_25811,N_25621,N_25646);
or U25812 (N_25812,N_25637,N_25568);
or U25813 (N_25813,N_25630,N_25566);
nor U25814 (N_25814,N_25712,N_25624);
and U25815 (N_25815,N_25660,N_25549);
or U25816 (N_25816,N_25742,N_25611);
nor U25817 (N_25817,N_25652,N_25596);
or U25818 (N_25818,N_25710,N_25582);
or U25819 (N_25819,N_25511,N_25715);
and U25820 (N_25820,N_25677,N_25504);
and U25821 (N_25821,N_25542,N_25559);
nand U25822 (N_25822,N_25595,N_25560);
and U25823 (N_25823,N_25744,N_25634);
xor U25824 (N_25824,N_25583,N_25541);
and U25825 (N_25825,N_25615,N_25629);
nor U25826 (N_25826,N_25563,N_25701);
or U25827 (N_25827,N_25515,N_25711);
and U25828 (N_25828,N_25697,N_25700);
or U25829 (N_25829,N_25513,N_25527);
nor U25830 (N_25830,N_25503,N_25573);
nand U25831 (N_25831,N_25516,N_25675);
nor U25832 (N_25832,N_25598,N_25600);
xnor U25833 (N_25833,N_25731,N_25509);
nor U25834 (N_25834,N_25680,N_25635);
and U25835 (N_25835,N_25551,N_25529);
and U25836 (N_25836,N_25617,N_25578);
nand U25837 (N_25837,N_25505,N_25525);
nand U25838 (N_25838,N_25614,N_25706);
xnor U25839 (N_25839,N_25510,N_25561);
or U25840 (N_25840,N_25641,N_25603);
xnor U25841 (N_25841,N_25572,N_25545);
and U25842 (N_25842,N_25693,N_25591);
nor U25843 (N_25843,N_25627,N_25565);
nand U25844 (N_25844,N_25745,N_25575);
nand U25845 (N_25845,N_25517,N_25730);
nor U25846 (N_25846,N_25729,N_25665);
or U25847 (N_25847,N_25708,N_25623);
or U25848 (N_25848,N_25739,N_25690);
nand U25849 (N_25849,N_25610,N_25689);
nor U25850 (N_25850,N_25748,N_25554);
or U25851 (N_25851,N_25613,N_25616);
nand U25852 (N_25852,N_25524,N_25521);
nand U25853 (N_25853,N_25644,N_25707);
or U25854 (N_25854,N_25628,N_25543);
nor U25855 (N_25855,N_25664,N_25593);
nand U25856 (N_25856,N_25720,N_25506);
xnor U25857 (N_25857,N_25523,N_25587);
nand U25858 (N_25858,N_25576,N_25655);
and U25859 (N_25859,N_25633,N_25674);
nand U25860 (N_25860,N_25580,N_25728);
nand U25861 (N_25861,N_25740,N_25738);
nor U25862 (N_25862,N_25539,N_25747);
nor U25863 (N_25863,N_25528,N_25625);
or U25864 (N_25864,N_25650,N_25570);
nand U25865 (N_25865,N_25734,N_25569);
and U25866 (N_25866,N_25535,N_25654);
nand U25867 (N_25867,N_25558,N_25581);
nand U25868 (N_25868,N_25502,N_25590);
or U25869 (N_25869,N_25684,N_25531);
nor U25870 (N_25870,N_25686,N_25604);
and U25871 (N_25871,N_25645,N_25666);
and U25872 (N_25872,N_25743,N_25620);
and U25873 (N_25873,N_25704,N_25722);
xor U25874 (N_25874,N_25594,N_25714);
nand U25875 (N_25875,N_25691,N_25685);
nand U25876 (N_25876,N_25648,N_25585);
or U25877 (N_25877,N_25731,N_25604);
nor U25878 (N_25878,N_25726,N_25624);
nand U25879 (N_25879,N_25632,N_25512);
and U25880 (N_25880,N_25682,N_25560);
or U25881 (N_25881,N_25509,N_25689);
xor U25882 (N_25882,N_25629,N_25597);
nand U25883 (N_25883,N_25594,N_25670);
nor U25884 (N_25884,N_25621,N_25520);
nand U25885 (N_25885,N_25704,N_25572);
xor U25886 (N_25886,N_25694,N_25564);
nand U25887 (N_25887,N_25672,N_25731);
or U25888 (N_25888,N_25596,N_25515);
nand U25889 (N_25889,N_25667,N_25648);
nand U25890 (N_25890,N_25623,N_25571);
nor U25891 (N_25891,N_25742,N_25703);
nor U25892 (N_25892,N_25722,N_25567);
and U25893 (N_25893,N_25726,N_25682);
nor U25894 (N_25894,N_25585,N_25601);
nand U25895 (N_25895,N_25603,N_25686);
nor U25896 (N_25896,N_25704,N_25600);
nand U25897 (N_25897,N_25616,N_25698);
or U25898 (N_25898,N_25584,N_25746);
nor U25899 (N_25899,N_25504,N_25681);
nand U25900 (N_25900,N_25508,N_25607);
nor U25901 (N_25901,N_25651,N_25660);
xor U25902 (N_25902,N_25524,N_25711);
xnor U25903 (N_25903,N_25581,N_25579);
and U25904 (N_25904,N_25728,N_25649);
and U25905 (N_25905,N_25518,N_25521);
or U25906 (N_25906,N_25702,N_25525);
xnor U25907 (N_25907,N_25558,N_25690);
nand U25908 (N_25908,N_25624,N_25655);
nor U25909 (N_25909,N_25711,N_25512);
nor U25910 (N_25910,N_25526,N_25632);
or U25911 (N_25911,N_25613,N_25588);
nor U25912 (N_25912,N_25555,N_25633);
nor U25913 (N_25913,N_25528,N_25541);
xor U25914 (N_25914,N_25671,N_25604);
or U25915 (N_25915,N_25704,N_25592);
or U25916 (N_25916,N_25739,N_25624);
xnor U25917 (N_25917,N_25670,N_25668);
xor U25918 (N_25918,N_25626,N_25593);
nor U25919 (N_25919,N_25723,N_25664);
xor U25920 (N_25920,N_25611,N_25668);
or U25921 (N_25921,N_25550,N_25561);
or U25922 (N_25922,N_25679,N_25735);
nand U25923 (N_25923,N_25622,N_25620);
nand U25924 (N_25924,N_25503,N_25613);
nand U25925 (N_25925,N_25728,N_25628);
or U25926 (N_25926,N_25562,N_25687);
xnor U25927 (N_25927,N_25567,N_25729);
nand U25928 (N_25928,N_25662,N_25548);
xor U25929 (N_25929,N_25612,N_25689);
xnor U25930 (N_25930,N_25713,N_25577);
xor U25931 (N_25931,N_25726,N_25536);
and U25932 (N_25932,N_25558,N_25664);
nand U25933 (N_25933,N_25502,N_25575);
or U25934 (N_25934,N_25616,N_25604);
xnor U25935 (N_25935,N_25517,N_25570);
nand U25936 (N_25936,N_25743,N_25677);
or U25937 (N_25937,N_25694,N_25620);
or U25938 (N_25938,N_25559,N_25705);
nand U25939 (N_25939,N_25620,N_25580);
nand U25940 (N_25940,N_25653,N_25568);
nand U25941 (N_25941,N_25647,N_25554);
nand U25942 (N_25942,N_25540,N_25634);
xor U25943 (N_25943,N_25609,N_25639);
or U25944 (N_25944,N_25528,N_25532);
nor U25945 (N_25945,N_25537,N_25694);
and U25946 (N_25946,N_25665,N_25710);
nor U25947 (N_25947,N_25584,N_25523);
and U25948 (N_25948,N_25745,N_25643);
nor U25949 (N_25949,N_25536,N_25628);
nand U25950 (N_25950,N_25704,N_25675);
xor U25951 (N_25951,N_25652,N_25712);
and U25952 (N_25952,N_25651,N_25696);
and U25953 (N_25953,N_25595,N_25578);
or U25954 (N_25954,N_25538,N_25699);
and U25955 (N_25955,N_25638,N_25652);
or U25956 (N_25956,N_25567,N_25624);
nand U25957 (N_25957,N_25707,N_25648);
and U25958 (N_25958,N_25579,N_25626);
and U25959 (N_25959,N_25602,N_25720);
nand U25960 (N_25960,N_25556,N_25612);
or U25961 (N_25961,N_25743,N_25746);
and U25962 (N_25962,N_25509,N_25606);
nand U25963 (N_25963,N_25514,N_25682);
or U25964 (N_25964,N_25718,N_25744);
nor U25965 (N_25965,N_25516,N_25692);
nor U25966 (N_25966,N_25578,N_25580);
and U25967 (N_25967,N_25563,N_25637);
or U25968 (N_25968,N_25630,N_25606);
nor U25969 (N_25969,N_25600,N_25560);
xnor U25970 (N_25970,N_25692,N_25565);
nand U25971 (N_25971,N_25540,N_25616);
and U25972 (N_25972,N_25524,N_25585);
nand U25973 (N_25973,N_25671,N_25554);
nand U25974 (N_25974,N_25697,N_25662);
nand U25975 (N_25975,N_25710,N_25704);
and U25976 (N_25976,N_25606,N_25679);
or U25977 (N_25977,N_25710,N_25617);
and U25978 (N_25978,N_25544,N_25713);
nor U25979 (N_25979,N_25682,N_25681);
and U25980 (N_25980,N_25618,N_25685);
nor U25981 (N_25981,N_25610,N_25723);
nand U25982 (N_25982,N_25657,N_25514);
or U25983 (N_25983,N_25557,N_25703);
or U25984 (N_25984,N_25740,N_25669);
and U25985 (N_25985,N_25545,N_25676);
xnor U25986 (N_25986,N_25661,N_25524);
nor U25987 (N_25987,N_25707,N_25641);
nor U25988 (N_25988,N_25708,N_25545);
and U25989 (N_25989,N_25681,N_25543);
or U25990 (N_25990,N_25583,N_25652);
nor U25991 (N_25991,N_25735,N_25669);
or U25992 (N_25992,N_25588,N_25514);
or U25993 (N_25993,N_25642,N_25612);
nand U25994 (N_25994,N_25579,N_25594);
or U25995 (N_25995,N_25609,N_25699);
or U25996 (N_25996,N_25565,N_25629);
nor U25997 (N_25997,N_25585,N_25622);
nand U25998 (N_25998,N_25595,N_25502);
nor U25999 (N_25999,N_25549,N_25615);
nand U26000 (N_26000,N_25936,N_25997);
xor U26001 (N_26001,N_25963,N_25855);
or U26002 (N_26002,N_25755,N_25767);
nor U26003 (N_26003,N_25846,N_25921);
nand U26004 (N_26004,N_25954,N_25874);
and U26005 (N_26005,N_25891,N_25901);
nor U26006 (N_26006,N_25838,N_25839);
nand U26007 (N_26007,N_25831,N_25800);
nand U26008 (N_26008,N_25906,N_25923);
or U26009 (N_26009,N_25845,N_25784);
and U26010 (N_26010,N_25961,N_25938);
nor U26011 (N_26011,N_25916,N_25824);
nor U26012 (N_26012,N_25822,N_25994);
nor U26013 (N_26013,N_25774,N_25865);
and U26014 (N_26014,N_25962,N_25934);
nand U26015 (N_26015,N_25917,N_25849);
xor U26016 (N_26016,N_25975,N_25763);
or U26017 (N_26017,N_25984,N_25853);
or U26018 (N_26018,N_25816,N_25796);
nand U26019 (N_26019,N_25752,N_25932);
nand U26020 (N_26020,N_25929,N_25753);
xnor U26021 (N_26021,N_25948,N_25858);
or U26022 (N_26022,N_25843,N_25996);
nor U26023 (N_26023,N_25789,N_25928);
nand U26024 (N_26024,N_25945,N_25804);
nor U26025 (N_26025,N_25818,N_25803);
and U26026 (N_26026,N_25903,N_25918);
xor U26027 (N_26027,N_25777,N_25915);
or U26028 (N_26028,N_25904,N_25905);
and U26029 (N_26029,N_25913,N_25968);
and U26030 (N_26030,N_25872,N_25814);
nor U26031 (N_26031,N_25942,N_25983);
nand U26032 (N_26032,N_25786,N_25992);
xnor U26033 (N_26033,N_25991,N_25788);
nand U26034 (N_26034,N_25958,N_25826);
nor U26035 (N_26035,N_25877,N_25890);
and U26036 (N_26036,N_25761,N_25880);
and U26037 (N_26037,N_25969,N_25768);
nand U26038 (N_26038,N_25980,N_25869);
nand U26039 (N_26039,N_25791,N_25893);
nor U26040 (N_26040,N_25909,N_25985);
nor U26041 (N_26041,N_25848,N_25771);
nand U26042 (N_26042,N_25940,N_25933);
nand U26043 (N_26043,N_25987,N_25993);
xnor U26044 (N_26044,N_25960,N_25896);
and U26045 (N_26045,N_25766,N_25785);
or U26046 (N_26046,N_25972,N_25805);
xor U26047 (N_26047,N_25790,N_25758);
or U26048 (N_26048,N_25876,N_25861);
nand U26049 (N_26049,N_25835,N_25782);
xor U26050 (N_26050,N_25943,N_25819);
xnor U26051 (N_26051,N_25939,N_25823);
nor U26052 (N_26052,N_25878,N_25998);
nand U26053 (N_26053,N_25799,N_25922);
nand U26054 (N_26054,N_25920,N_25829);
and U26055 (N_26055,N_25947,N_25851);
xnor U26056 (N_26056,N_25926,N_25908);
xor U26057 (N_26057,N_25817,N_25875);
or U26058 (N_26058,N_25952,N_25966);
nand U26059 (N_26059,N_25895,N_25836);
xnor U26060 (N_26060,N_25950,N_25854);
nand U26061 (N_26061,N_25937,N_25820);
nor U26062 (N_26062,N_25825,N_25783);
nor U26063 (N_26063,N_25981,N_25859);
nor U26064 (N_26064,N_25870,N_25931);
xnor U26065 (N_26065,N_25828,N_25863);
or U26066 (N_26066,N_25976,N_25852);
nor U26067 (N_26067,N_25965,N_25775);
nor U26068 (N_26068,N_25873,N_25941);
and U26069 (N_26069,N_25956,N_25759);
or U26070 (N_26070,N_25779,N_25889);
nor U26071 (N_26071,N_25770,N_25949);
xnor U26072 (N_26072,N_25812,N_25776);
xnor U26073 (N_26073,N_25794,N_25862);
nand U26074 (N_26074,N_25887,N_25857);
and U26075 (N_26075,N_25850,N_25955);
or U26076 (N_26076,N_25864,N_25807);
or U26077 (N_26077,N_25912,N_25971);
nor U26078 (N_26078,N_25888,N_25750);
nor U26079 (N_26079,N_25856,N_25982);
nand U26080 (N_26080,N_25977,N_25798);
xor U26081 (N_26081,N_25990,N_25795);
and U26082 (N_26082,N_25860,N_25793);
or U26083 (N_26083,N_25765,N_25867);
nand U26084 (N_26084,N_25757,N_25964);
or U26085 (N_26085,N_25897,N_25914);
xor U26086 (N_26086,N_25830,N_25844);
nor U26087 (N_26087,N_25847,N_25959);
nand U26088 (N_26088,N_25886,N_25935);
or U26089 (N_26089,N_25883,N_25810);
nor U26090 (N_26090,N_25986,N_25866);
nand U26091 (N_26091,N_25762,N_25988);
and U26092 (N_26092,N_25871,N_25885);
nor U26093 (N_26093,N_25751,N_25815);
or U26094 (N_26094,N_25780,N_25868);
nand U26095 (N_26095,N_25884,N_25892);
xor U26096 (N_26096,N_25787,N_25910);
and U26097 (N_26097,N_25879,N_25808);
xor U26098 (N_26098,N_25953,N_25999);
or U26099 (N_26099,N_25806,N_25827);
nand U26100 (N_26100,N_25927,N_25773);
nand U26101 (N_26101,N_25973,N_25772);
and U26102 (N_26102,N_25778,N_25967);
and U26103 (N_26103,N_25809,N_25989);
nand U26104 (N_26104,N_25813,N_25769);
nand U26105 (N_26105,N_25833,N_25811);
or U26106 (N_26106,N_25754,N_25925);
nor U26107 (N_26107,N_25894,N_25781);
nand U26108 (N_26108,N_25902,N_25802);
and U26109 (N_26109,N_25837,N_25801);
nor U26110 (N_26110,N_25842,N_25821);
nand U26111 (N_26111,N_25907,N_25957);
and U26112 (N_26112,N_25979,N_25832);
xor U26113 (N_26113,N_25840,N_25995);
nor U26114 (N_26114,N_25951,N_25797);
or U26115 (N_26115,N_25834,N_25930);
nand U26116 (N_26116,N_25899,N_25756);
nand U26117 (N_26117,N_25882,N_25944);
nand U26118 (N_26118,N_25919,N_25911);
xnor U26119 (N_26119,N_25900,N_25764);
nand U26120 (N_26120,N_25970,N_25898);
or U26121 (N_26121,N_25760,N_25924);
nor U26122 (N_26122,N_25978,N_25841);
xnor U26123 (N_26123,N_25881,N_25792);
nand U26124 (N_26124,N_25974,N_25946);
xor U26125 (N_26125,N_25893,N_25795);
and U26126 (N_26126,N_25979,N_25930);
nor U26127 (N_26127,N_25987,N_25875);
or U26128 (N_26128,N_25759,N_25945);
nand U26129 (N_26129,N_25848,N_25876);
xor U26130 (N_26130,N_25848,N_25905);
and U26131 (N_26131,N_25783,N_25797);
or U26132 (N_26132,N_25895,N_25917);
xor U26133 (N_26133,N_25750,N_25762);
nand U26134 (N_26134,N_25833,N_25834);
nor U26135 (N_26135,N_25841,N_25961);
or U26136 (N_26136,N_25881,N_25763);
nor U26137 (N_26137,N_25931,N_25849);
and U26138 (N_26138,N_25930,N_25806);
nand U26139 (N_26139,N_25883,N_25862);
nand U26140 (N_26140,N_25970,N_25791);
or U26141 (N_26141,N_25981,N_25951);
nand U26142 (N_26142,N_25853,N_25999);
or U26143 (N_26143,N_25807,N_25910);
nor U26144 (N_26144,N_25944,N_25811);
and U26145 (N_26145,N_25796,N_25907);
nand U26146 (N_26146,N_25995,N_25915);
or U26147 (N_26147,N_25878,N_25953);
or U26148 (N_26148,N_25793,N_25828);
or U26149 (N_26149,N_25758,N_25901);
nand U26150 (N_26150,N_25758,N_25927);
xor U26151 (N_26151,N_25894,N_25910);
and U26152 (N_26152,N_25781,N_25804);
xnor U26153 (N_26153,N_25778,N_25814);
or U26154 (N_26154,N_25783,N_25753);
nor U26155 (N_26155,N_25782,N_25947);
nand U26156 (N_26156,N_25822,N_25952);
and U26157 (N_26157,N_25937,N_25964);
nand U26158 (N_26158,N_25888,N_25991);
and U26159 (N_26159,N_25903,N_25864);
and U26160 (N_26160,N_25953,N_25875);
nor U26161 (N_26161,N_25831,N_25906);
xor U26162 (N_26162,N_25980,N_25761);
xor U26163 (N_26163,N_25929,N_25885);
xor U26164 (N_26164,N_25990,N_25943);
nor U26165 (N_26165,N_25774,N_25840);
nor U26166 (N_26166,N_25886,N_25779);
nand U26167 (N_26167,N_25824,N_25754);
and U26168 (N_26168,N_25797,N_25819);
or U26169 (N_26169,N_25851,N_25773);
and U26170 (N_26170,N_25857,N_25767);
or U26171 (N_26171,N_25858,N_25918);
or U26172 (N_26172,N_25840,N_25914);
nor U26173 (N_26173,N_25912,N_25791);
xor U26174 (N_26174,N_25999,N_25842);
xor U26175 (N_26175,N_25987,N_25765);
xor U26176 (N_26176,N_25986,N_25993);
nand U26177 (N_26177,N_25807,N_25889);
xnor U26178 (N_26178,N_25900,N_25822);
nor U26179 (N_26179,N_25853,N_25820);
nor U26180 (N_26180,N_25843,N_25948);
xor U26181 (N_26181,N_25787,N_25774);
nand U26182 (N_26182,N_25920,N_25897);
nor U26183 (N_26183,N_25773,N_25784);
and U26184 (N_26184,N_25983,N_25796);
nor U26185 (N_26185,N_25871,N_25889);
nand U26186 (N_26186,N_25855,N_25770);
nor U26187 (N_26187,N_25969,N_25940);
nor U26188 (N_26188,N_25840,N_25815);
nand U26189 (N_26189,N_25918,N_25895);
nand U26190 (N_26190,N_25881,N_25874);
or U26191 (N_26191,N_25779,N_25907);
or U26192 (N_26192,N_25980,N_25931);
or U26193 (N_26193,N_25878,N_25849);
xor U26194 (N_26194,N_25984,N_25937);
or U26195 (N_26195,N_25902,N_25815);
and U26196 (N_26196,N_25914,N_25779);
and U26197 (N_26197,N_25969,N_25990);
nand U26198 (N_26198,N_25801,N_25996);
nor U26199 (N_26199,N_25947,N_25866);
or U26200 (N_26200,N_25805,N_25919);
and U26201 (N_26201,N_25952,N_25944);
or U26202 (N_26202,N_25894,N_25849);
xnor U26203 (N_26203,N_25781,N_25964);
nor U26204 (N_26204,N_25947,N_25985);
nor U26205 (N_26205,N_25918,N_25814);
xnor U26206 (N_26206,N_25924,N_25932);
or U26207 (N_26207,N_25981,N_25833);
and U26208 (N_26208,N_25844,N_25976);
xor U26209 (N_26209,N_25984,N_25796);
and U26210 (N_26210,N_25877,N_25943);
xnor U26211 (N_26211,N_25851,N_25878);
or U26212 (N_26212,N_25849,N_25927);
nor U26213 (N_26213,N_25782,N_25859);
and U26214 (N_26214,N_25936,N_25852);
xor U26215 (N_26215,N_25919,N_25908);
or U26216 (N_26216,N_25818,N_25900);
nand U26217 (N_26217,N_25955,N_25921);
nor U26218 (N_26218,N_25805,N_25774);
nand U26219 (N_26219,N_25843,N_25920);
nor U26220 (N_26220,N_25772,N_25789);
nor U26221 (N_26221,N_25935,N_25814);
xnor U26222 (N_26222,N_25951,N_25769);
nand U26223 (N_26223,N_25887,N_25787);
nor U26224 (N_26224,N_25754,N_25847);
xor U26225 (N_26225,N_25944,N_25878);
or U26226 (N_26226,N_25904,N_25765);
or U26227 (N_26227,N_25909,N_25848);
xor U26228 (N_26228,N_25759,N_25859);
and U26229 (N_26229,N_25968,N_25879);
or U26230 (N_26230,N_25859,N_25832);
xor U26231 (N_26231,N_25838,N_25934);
or U26232 (N_26232,N_25791,N_25760);
xor U26233 (N_26233,N_25933,N_25838);
or U26234 (N_26234,N_25993,N_25983);
nor U26235 (N_26235,N_25834,N_25920);
nor U26236 (N_26236,N_25946,N_25759);
and U26237 (N_26237,N_25790,N_25893);
xor U26238 (N_26238,N_25855,N_25910);
nor U26239 (N_26239,N_25940,N_25798);
or U26240 (N_26240,N_25843,N_25896);
nor U26241 (N_26241,N_25945,N_25756);
and U26242 (N_26242,N_25926,N_25990);
nor U26243 (N_26243,N_25852,N_25895);
and U26244 (N_26244,N_25863,N_25797);
and U26245 (N_26245,N_25951,N_25816);
nor U26246 (N_26246,N_25754,N_25926);
nor U26247 (N_26247,N_25896,N_25950);
xnor U26248 (N_26248,N_25837,N_25952);
or U26249 (N_26249,N_25985,N_25781);
xor U26250 (N_26250,N_26170,N_26040);
xor U26251 (N_26251,N_26147,N_26199);
nand U26252 (N_26252,N_26210,N_26217);
nand U26253 (N_26253,N_26052,N_26214);
nand U26254 (N_26254,N_26127,N_26169);
nor U26255 (N_26255,N_26013,N_26070);
and U26256 (N_26256,N_26102,N_26134);
or U26257 (N_26257,N_26032,N_26002);
nand U26258 (N_26258,N_26171,N_26145);
nand U26259 (N_26259,N_26229,N_26004);
nand U26260 (N_26260,N_26187,N_26164);
or U26261 (N_26261,N_26248,N_26200);
or U26262 (N_26262,N_26131,N_26192);
nor U26263 (N_26263,N_26156,N_26238);
xnor U26264 (N_26264,N_26003,N_26189);
nand U26265 (N_26265,N_26057,N_26188);
nor U26266 (N_26266,N_26218,N_26033);
nand U26267 (N_26267,N_26235,N_26031);
nor U26268 (N_26268,N_26198,N_26072);
nor U26269 (N_26269,N_26159,N_26101);
and U26270 (N_26270,N_26028,N_26104);
or U26271 (N_26271,N_26008,N_26154);
xnor U26272 (N_26272,N_26020,N_26148);
xor U26273 (N_26273,N_26236,N_26026);
and U26274 (N_26274,N_26015,N_26066);
nand U26275 (N_26275,N_26086,N_26146);
or U26276 (N_26276,N_26074,N_26046);
and U26277 (N_26277,N_26185,N_26044);
or U26278 (N_26278,N_26120,N_26021);
and U26279 (N_26279,N_26191,N_26163);
and U26280 (N_26280,N_26166,N_26065);
nand U26281 (N_26281,N_26241,N_26000);
nor U26282 (N_26282,N_26230,N_26081);
xnor U26283 (N_26283,N_26228,N_26119);
nor U26284 (N_26284,N_26221,N_26062);
nand U26285 (N_26285,N_26149,N_26056);
and U26286 (N_26286,N_26224,N_26155);
nand U26287 (N_26287,N_26007,N_26245);
nor U26288 (N_26288,N_26115,N_26121);
nand U26289 (N_26289,N_26076,N_26075);
nand U26290 (N_26290,N_26247,N_26097);
nand U26291 (N_26291,N_26124,N_26093);
and U26292 (N_26292,N_26181,N_26012);
xor U26293 (N_26293,N_26205,N_26014);
and U26294 (N_26294,N_26165,N_26157);
xor U26295 (N_26295,N_26135,N_26116);
and U26296 (N_26296,N_26233,N_26047);
nor U26297 (N_26297,N_26035,N_26091);
nor U26298 (N_26298,N_26058,N_26197);
nor U26299 (N_26299,N_26136,N_26055);
nand U26300 (N_26300,N_26195,N_26194);
xor U26301 (N_26301,N_26051,N_26069);
xnor U26302 (N_26302,N_26025,N_26078);
and U26303 (N_26303,N_26034,N_26050);
xor U26304 (N_26304,N_26161,N_26118);
and U26305 (N_26305,N_26213,N_26193);
and U26306 (N_26306,N_26173,N_26010);
or U26307 (N_26307,N_26080,N_26130);
nand U26308 (N_26308,N_26107,N_26018);
and U26309 (N_26309,N_26137,N_26158);
and U26310 (N_26310,N_26242,N_26222);
and U26311 (N_26311,N_26125,N_26207);
or U26312 (N_26312,N_26095,N_26140);
xor U26313 (N_26313,N_26223,N_26182);
xor U26314 (N_26314,N_26098,N_26001);
xnor U26315 (N_26315,N_26152,N_26184);
xor U26316 (N_26316,N_26243,N_26085);
nor U26317 (N_26317,N_26246,N_26240);
or U26318 (N_26318,N_26216,N_26175);
and U26319 (N_26319,N_26123,N_26082);
or U26320 (N_26320,N_26167,N_26005);
xor U26321 (N_26321,N_26024,N_26160);
nor U26322 (N_26322,N_26249,N_26179);
nor U26323 (N_26323,N_26113,N_26105);
nand U26324 (N_26324,N_26144,N_26022);
or U26325 (N_26325,N_26211,N_26029);
nor U26326 (N_26326,N_26219,N_26079);
and U26327 (N_26327,N_26030,N_26094);
nand U26328 (N_26328,N_26239,N_26183);
nand U26329 (N_26329,N_26049,N_26225);
or U26330 (N_26330,N_26178,N_26206);
xor U26331 (N_26331,N_26162,N_26109);
xor U26332 (N_26332,N_26073,N_26176);
and U26333 (N_26333,N_26133,N_26016);
xnor U26334 (N_26334,N_26111,N_26043);
nand U26335 (N_26335,N_26132,N_26143);
nor U26336 (N_26336,N_26009,N_26168);
nor U26337 (N_26337,N_26174,N_26090);
nand U26338 (N_26338,N_26060,N_26038);
xnor U26339 (N_26339,N_26063,N_26037);
nand U26340 (N_26340,N_26054,N_26017);
xnor U26341 (N_26341,N_26208,N_26201);
xnor U26342 (N_26342,N_26106,N_26108);
nand U26343 (N_26343,N_26226,N_26244);
nor U26344 (N_26344,N_26019,N_26142);
and U26345 (N_26345,N_26128,N_26129);
nor U26346 (N_26346,N_26084,N_26203);
or U26347 (N_26347,N_26077,N_26064);
xnor U26348 (N_26348,N_26138,N_26041);
or U26349 (N_26349,N_26067,N_26153);
and U26350 (N_26350,N_26122,N_26089);
nand U26351 (N_26351,N_26087,N_26204);
nand U26352 (N_26352,N_26103,N_26068);
nor U26353 (N_26353,N_26011,N_26100);
nand U26354 (N_26354,N_26112,N_26150);
nor U26355 (N_26355,N_26039,N_26045);
nor U26356 (N_26356,N_26096,N_26083);
or U26357 (N_26357,N_26006,N_26220);
or U26358 (N_26358,N_26231,N_26186);
nand U26359 (N_26359,N_26036,N_26126);
nor U26360 (N_26360,N_26053,N_26172);
xnor U26361 (N_26361,N_26227,N_26092);
nor U26362 (N_26362,N_26237,N_26042);
nor U26363 (N_26363,N_26048,N_26151);
xnor U26364 (N_26364,N_26023,N_26059);
nand U26365 (N_26365,N_26190,N_26099);
nand U26366 (N_26366,N_26071,N_26027);
or U26367 (N_26367,N_26180,N_26232);
nor U26368 (N_26368,N_26139,N_26117);
or U26369 (N_26369,N_26215,N_26088);
nor U26370 (N_26370,N_26061,N_26212);
nand U26371 (N_26371,N_26196,N_26209);
and U26372 (N_26372,N_26110,N_26114);
and U26373 (N_26373,N_26202,N_26234);
nor U26374 (N_26374,N_26177,N_26141);
nor U26375 (N_26375,N_26032,N_26067);
nand U26376 (N_26376,N_26144,N_26047);
and U26377 (N_26377,N_26090,N_26103);
and U26378 (N_26378,N_26244,N_26025);
and U26379 (N_26379,N_26092,N_26086);
nand U26380 (N_26380,N_26140,N_26185);
or U26381 (N_26381,N_26234,N_26136);
or U26382 (N_26382,N_26182,N_26161);
nor U26383 (N_26383,N_26058,N_26127);
nor U26384 (N_26384,N_26159,N_26172);
and U26385 (N_26385,N_26066,N_26164);
and U26386 (N_26386,N_26044,N_26225);
xor U26387 (N_26387,N_26039,N_26154);
nor U26388 (N_26388,N_26148,N_26146);
nand U26389 (N_26389,N_26052,N_26177);
or U26390 (N_26390,N_26073,N_26239);
nor U26391 (N_26391,N_26136,N_26007);
nand U26392 (N_26392,N_26020,N_26221);
or U26393 (N_26393,N_26192,N_26082);
xnor U26394 (N_26394,N_26235,N_26009);
and U26395 (N_26395,N_26080,N_26150);
or U26396 (N_26396,N_26249,N_26155);
nand U26397 (N_26397,N_26200,N_26112);
or U26398 (N_26398,N_26175,N_26240);
or U26399 (N_26399,N_26239,N_26000);
or U26400 (N_26400,N_26018,N_26015);
and U26401 (N_26401,N_26188,N_26098);
nor U26402 (N_26402,N_26184,N_26025);
xor U26403 (N_26403,N_26117,N_26176);
nor U26404 (N_26404,N_26241,N_26155);
or U26405 (N_26405,N_26091,N_26037);
nand U26406 (N_26406,N_26211,N_26021);
xnor U26407 (N_26407,N_26184,N_26105);
and U26408 (N_26408,N_26087,N_26191);
or U26409 (N_26409,N_26100,N_26146);
xor U26410 (N_26410,N_26064,N_26045);
nand U26411 (N_26411,N_26105,N_26229);
nand U26412 (N_26412,N_26013,N_26201);
xnor U26413 (N_26413,N_26154,N_26092);
nor U26414 (N_26414,N_26045,N_26152);
or U26415 (N_26415,N_26037,N_26217);
xnor U26416 (N_26416,N_26164,N_26050);
nor U26417 (N_26417,N_26210,N_26156);
nor U26418 (N_26418,N_26245,N_26230);
and U26419 (N_26419,N_26034,N_26151);
and U26420 (N_26420,N_26131,N_26030);
xnor U26421 (N_26421,N_26043,N_26081);
nand U26422 (N_26422,N_26218,N_26075);
nand U26423 (N_26423,N_26134,N_26234);
xnor U26424 (N_26424,N_26156,N_26189);
nor U26425 (N_26425,N_26160,N_26169);
or U26426 (N_26426,N_26041,N_26006);
nor U26427 (N_26427,N_26197,N_26236);
xnor U26428 (N_26428,N_26219,N_26109);
and U26429 (N_26429,N_26187,N_26234);
and U26430 (N_26430,N_26164,N_26149);
nor U26431 (N_26431,N_26141,N_26077);
xnor U26432 (N_26432,N_26133,N_26104);
nand U26433 (N_26433,N_26035,N_26144);
or U26434 (N_26434,N_26244,N_26190);
nand U26435 (N_26435,N_26221,N_26018);
or U26436 (N_26436,N_26179,N_26243);
nand U26437 (N_26437,N_26239,N_26039);
and U26438 (N_26438,N_26146,N_26074);
xor U26439 (N_26439,N_26216,N_26077);
nor U26440 (N_26440,N_26069,N_26041);
nor U26441 (N_26441,N_26177,N_26161);
nand U26442 (N_26442,N_26012,N_26066);
nor U26443 (N_26443,N_26204,N_26009);
xnor U26444 (N_26444,N_26104,N_26011);
xor U26445 (N_26445,N_26173,N_26157);
and U26446 (N_26446,N_26000,N_26040);
and U26447 (N_26447,N_26120,N_26076);
nand U26448 (N_26448,N_26182,N_26096);
nand U26449 (N_26449,N_26236,N_26242);
or U26450 (N_26450,N_26030,N_26044);
xnor U26451 (N_26451,N_26118,N_26059);
or U26452 (N_26452,N_26037,N_26054);
xnor U26453 (N_26453,N_26137,N_26134);
xor U26454 (N_26454,N_26213,N_26079);
and U26455 (N_26455,N_26059,N_26140);
xnor U26456 (N_26456,N_26009,N_26148);
xnor U26457 (N_26457,N_26079,N_26086);
or U26458 (N_26458,N_26126,N_26135);
or U26459 (N_26459,N_26163,N_26038);
nor U26460 (N_26460,N_26058,N_26043);
xor U26461 (N_26461,N_26097,N_26121);
nor U26462 (N_26462,N_26193,N_26123);
or U26463 (N_26463,N_26031,N_26217);
nor U26464 (N_26464,N_26111,N_26150);
nor U26465 (N_26465,N_26072,N_26178);
and U26466 (N_26466,N_26237,N_26095);
nand U26467 (N_26467,N_26124,N_26212);
nor U26468 (N_26468,N_26077,N_26106);
nor U26469 (N_26469,N_26173,N_26175);
or U26470 (N_26470,N_26182,N_26045);
nand U26471 (N_26471,N_26186,N_26183);
or U26472 (N_26472,N_26072,N_26067);
and U26473 (N_26473,N_26237,N_26111);
nor U26474 (N_26474,N_26228,N_26010);
nor U26475 (N_26475,N_26189,N_26146);
xnor U26476 (N_26476,N_26077,N_26149);
xor U26477 (N_26477,N_26228,N_26120);
and U26478 (N_26478,N_26102,N_26248);
nand U26479 (N_26479,N_26046,N_26165);
nor U26480 (N_26480,N_26168,N_26046);
and U26481 (N_26481,N_26198,N_26135);
and U26482 (N_26482,N_26233,N_26080);
and U26483 (N_26483,N_26162,N_26032);
xor U26484 (N_26484,N_26023,N_26109);
nor U26485 (N_26485,N_26099,N_26113);
and U26486 (N_26486,N_26212,N_26095);
nor U26487 (N_26487,N_26138,N_26010);
nor U26488 (N_26488,N_26217,N_26062);
xnor U26489 (N_26489,N_26061,N_26115);
nor U26490 (N_26490,N_26090,N_26060);
nor U26491 (N_26491,N_26183,N_26227);
and U26492 (N_26492,N_26005,N_26243);
xor U26493 (N_26493,N_26051,N_26186);
or U26494 (N_26494,N_26199,N_26208);
nor U26495 (N_26495,N_26194,N_26187);
nand U26496 (N_26496,N_26103,N_26146);
nor U26497 (N_26497,N_26003,N_26114);
nand U26498 (N_26498,N_26129,N_26207);
nand U26499 (N_26499,N_26106,N_26140);
nor U26500 (N_26500,N_26352,N_26250);
or U26501 (N_26501,N_26439,N_26410);
and U26502 (N_26502,N_26337,N_26457);
or U26503 (N_26503,N_26325,N_26458);
nor U26504 (N_26504,N_26252,N_26422);
nand U26505 (N_26505,N_26329,N_26398);
nor U26506 (N_26506,N_26386,N_26481);
nor U26507 (N_26507,N_26276,N_26326);
xor U26508 (N_26508,N_26357,N_26469);
or U26509 (N_26509,N_26254,N_26423);
nand U26510 (N_26510,N_26344,N_26478);
nor U26511 (N_26511,N_26402,N_26354);
xnor U26512 (N_26512,N_26408,N_26346);
nand U26513 (N_26513,N_26287,N_26328);
xor U26514 (N_26514,N_26496,N_26345);
xor U26515 (N_26515,N_26373,N_26332);
or U26516 (N_26516,N_26343,N_26451);
or U26517 (N_26517,N_26445,N_26434);
xor U26518 (N_26518,N_26319,N_26286);
or U26519 (N_26519,N_26347,N_26342);
nor U26520 (N_26520,N_26427,N_26259);
and U26521 (N_26521,N_26388,N_26257);
nand U26522 (N_26522,N_26338,N_26455);
xor U26523 (N_26523,N_26487,N_26311);
or U26524 (N_26524,N_26269,N_26376);
or U26525 (N_26525,N_26355,N_26403);
and U26526 (N_26526,N_26281,N_26494);
xor U26527 (N_26527,N_26264,N_26300);
nand U26528 (N_26528,N_26397,N_26277);
nor U26529 (N_26529,N_26375,N_26415);
and U26530 (N_26530,N_26411,N_26335);
nor U26531 (N_26531,N_26413,N_26462);
nand U26532 (N_26532,N_26380,N_26409);
or U26533 (N_26533,N_26449,N_26468);
nor U26534 (N_26534,N_26480,N_26392);
xnor U26535 (N_26535,N_26255,N_26369);
nand U26536 (N_26536,N_26285,N_26336);
and U26537 (N_26537,N_26479,N_26266);
nor U26538 (N_26538,N_26321,N_26459);
or U26539 (N_26539,N_26327,N_26492);
nor U26540 (N_26540,N_26367,N_26293);
xor U26541 (N_26541,N_26384,N_26333);
nor U26542 (N_26542,N_26348,N_26491);
and U26543 (N_26543,N_26283,N_26405);
or U26544 (N_26544,N_26467,N_26256);
nor U26545 (N_26545,N_26289,N_26273);
nand U26546 (N_26546,N_26251,N_26441);
nor U26547 (N_26547,N_26443,N_26368);
nand U26548 (N_26548,N_26301,N_26452);
and U26549 (N_26549,N_26359,N_26331);
nor U26550 (N_26550,N_26280,N_26262);
and U26551 (N_26551,N_26378,N_26450);
xor U26552 (N_26552,N_26270,N_26362);
and U26553 (N_26553,N_26340,N_26486);
xnor U26554 (N_26554,N_26391,N_26282);
xor U26555 (N_26555,N_26475,N_26278);
nand U26556 (N_26556,N_26428,N_26490);
and U26557 (N_26557,N_26306,N_26431);
and U26558 (N_26558,N_26253,N_26417);
or U26559 (N_26559,N_26330,N_26353);
and U26560 (N_26560,N_26498,N_26298);
xor U26561 (N_26561,N_26303,N_26361);
nand U26562 (N_26562,N_26442,N_26387);
and U26563 (N_26563,N_26472,N_26482);
and U26564 (N_26564,N_26260,N_26297);
xnor U26565 (N_26565,N_26320,N_26390);
nand U26566 (N_26566,N_26274,N_26272);
or U26567 (N_26567,N_26485,N_26460);
nand U26568 (N_26568,N_26436,N_26495);
nor U26569 (N_26569,N_26477,N_26341);
and U26570 (N_26570,N_26322,N_26385);
nor U26571 (N_26571,N_26324,N_26315);
and U26572 (N_26572,N_26424,N_26399);
and U26573 (N_26573,N_26493,N_26377);
nor U26574 (N_26574,N_26371,N_26407);
xnor U26575 (N_26575,N_26454,N_26383);
or U26576 (N_26576,N_26379,N_26316);
nor U26577 (N_26577,N_26366,N_26265);
nand U26578 (N_26578,N_26288,N_26483);
nor U26579 (N_26579,N_26295,N_26263);
and U26580 (N_26580,N_26365,N_26464);
and U26581 (N_26581,N_26356,N_26395);
nor U26582 (N_26582,N_26374,N_26444);
and U26583 (N_26583,N_26349,N_26425);
nand U26584 (N_26584,N_26406,N_26430);
xor U26585 (N_26585,N_26393,N_26473);
nand U26586 (N_26586,N_26302,N_26292);
and U26587 (N_26587,N_26418,N_26489);
xor U26588 (N_26588,N_26275,N_26317);
nor U26589 (N_26589,N_26394,N_26279);
or U26590 (N_26590,N_26318,N_26404);
or U26591 (N_26591,N_26463,N_26305);
nor U26592 (N_26592,N_26358,N_26401);
and U26593 (N_26593,N_26261,N_26372);
or U26594 (N_26594,N_26351,N_26304);
and U26595 (N_26595,N_26446,N_26291);
or U26596 (N_26596,N_26440,N_26309);
nand U26597 (N_26597,N_26433,N_26313);
nand U26598 (N_26598,N_26334,N_26381);
or U26599 (N_26599,N_26310,N_26299);
nand U26600 (N_26600,N_26453,N_26471);
nor U26601 (N_26601,N_26426,N_26438);
or U26602 (N_26602,N_26448,N_26465);
and U26603 (N_26603,N_26360,N_26497);
nor U26604 (N_26604,N_26466,N_26284);
xnor U26605 (N_26605,N_26400,N_26421);
nor U26606 (N_26606,N_26470,N_26461);
or U26607 (N_26607,N_26432,N_26420);
nor U26608 (N_26608,N_26416,N_26307);
and U26609 (N_26609,N_26258,N_26267);
and U26610 (N_26610,N_26419,N_26364);
nor U26611 (N_26611,N_26294,N_26429);
or U26612 (N_26612,N_26323,N_26474);
nand U26613 (N_26613,N_26499,N_26339);
nor U26614 (N_26614,N_26350,N_26363);
nand U26615 (N_26615,N_26271,N_26447);
or U26616 (N_26616,N_26312,N_26382);
or U26617 (N_26617,N_26389,N_26308);
nor U26618 (N_26618,N_26268,N_26412);
or U26619 (N_26619,N_26488,N_26476);
and U26620 (N_26620,N_26296,N_26437);
or U26621 (N_26621,N_26314,N_26484);
or U26622 (N_26622,N_26370,N_26414);
xnor U26623 (N_26623,N_26435,N_26456);
nor U26624 (N_26624,N_26290,N_26396);
nor U26625 (N_26625,N_26337,N_26443);
xor U26626 (N_26626,N_26477,N_26282);
nand U26627 (N_26627,N_26482,N_26356);
and U26628 (N_26628,N_26268,N_26338);
and U26629 (N_26629,N_26267,N_26280);
nor U26630 (N_26630,N_26370,N_26452);
and U26631 (N_26631,N_26307,N_26363);
or U26632 (N_26632,N_26331,N_26470);
nand U26633 (N_26633,N_26484,N_26383);
or U26634 (N_26634,N_26472,N_26256);
nand U26635 (N_26635,N_26335,N_26499);
and U26636 (N_26636,N_26452,N_26261);
or U26637 (N_26637,N_26491,N_26416);
or U26638 (N_26638,N_26419,N_26494);
and U26639 (N_26639,N_26382,N_26482);
xnor U26640 (N_26640,N_26419,N_26283);
or U26641 (N_26641,N_26353,N_26415);
nand U26642 (N_26642,N_26251,N_26253);
nor U26643 (N_26643,N_26305,N_26387);
or U26644 (N_26644,N_26476,N_26445);
xor U26645 (N_26645,N_26267,N_26300);
xor U26646 (N_26646,N_26343,N_26287);
and U26647 (N_26647,N_26489,N_26368);
and U26648 (N_26648,N_26277,N_26359);
nand U26649 (N_26649,N_26311,N_26295);
or U26650 (N_26650,N_26263,N_26474);
or U26651 (N_26651,N_26353,N_26297);
and U26652 (N_26652,N_26364,N_26315);
nor U26653 (N_26653,N_26289,N_26357);
and U26654 (N_26654,N_26268,N_26319);
nand U26655 (N_26655,N_26351,N_26359);
and U26656 (N_26656,N_26261,N_26483);
or U26657 (N_26657,N_26489,N_26275);
nand U26658 (N_26658,N_26479,N_26302);
or U26659 (N_26659,N_26424,N_26270);
nor U26660 (N_26660,N_26457,N_26468);
nor U26661 (N_26661,N_26308,N_26368);
and U26662 (N_26662,N_26310,N_26309);
xnor U26663 (N_26663,N_26496,N_26415);
nand U26664 (N_26664,N_26476,N_26439);
nor U26665 (N_26665,N_26366,N_26365);
nor U26666 (N_26666,N_26304,N_26335);
and U26667 (N_26667,N_26338,N_26401);
or U26668 (N_26668,N_26310,N_26368);
nand U26669 (N_26669,N_26335,N_26259);
nor U26670 (N_26670,N_26425,N_26251);
nor U26671 (N_26671,N_26373,N_26325);
or U26672 (N_26672,N_26253,N_26372);
nand U26673 (N_26673,N_26285,N_26360);
nor U26674 (N_26674,N_26291,N_26441);
or U26675 (N_26675,N_26267,N_26380);
or U26676 (N_26676,N_26266,N_26415);
and U26677 (N_26677,N_26416,N_26274);
nand U26678 (N_26678,N_26373,N_26412);
nand U26679 (N_26679,N_26360,N_26450);
nand U26680 (N_26680,N_26255,N_26285);
nor U26681 (N_26681,N_26320,N_26497);
and U26682 (N_26682,N_26300,N_26256);
nor U26683 (N_26683,N_26420,N_26460);
and U26684 (N_26684,N_26452,N_26366);
nor U26685 (N_26685,N_26455,N_26339);
or U26686 (N_26686,N_26485,N_26276);
xnor U26687 (N_26687,N_26430,N_26440);
nand U26688 (N_26688,N_26428,N_26346);
xor U26689 (N_26689,N_26446,N_26375);
or U26690 (N_26690,N_26387,N_26372);
or U26691 (N_26691,N_26332,N_26418);
or U26692 (N_26692,N_26401,N_26259);
xnor U26693 (N_26693,N_26485,N_26439);
and U26694 (N_26694,N_26474,N_26328);
nor U26695 (N_26695,N_26359,N_26325);
and U26696 (N_26696,N_26352,N_26397);
and U26697 (N_26697,N_26356,N_26496);
nand U26698 (N_26698,N_26476,N_26320);
or U26699 (N_26699,N_26336,N_26465);
nor U26700 (N_26700,N_26364,N_26367);
nand U26701 (N_26701,N_26376,N_26293);
or U26702 (N_26702,N_26287,N_26453);
or U26703 (N_26703,N_26320,N_26499);
xnor U26704 (N_26704,N_26462,N_26437);
nand U26705 (N_26705,N_26486,N_26363);
and U26706 (N_26706,N_26405,N_26295);
nand U26707 (N_26707,N_26364,N_26417);
nand U26708 (N_26708,N_26316,N_26265);
and U26709 (N_26709,N_26261,N_26425);
nor U26710 (N_26710,N_26262,N_26347);
nand U26711 (N_26711,N_26330,N_26369);
or U26712 (N_26712,N_26259,N_26374);
nor U26713 (N_26713,N_26472,N_26358);
or U26714 (N_26714,N_26316,N_26287);
xnor U26715 (N_26715,N_26479,N_26405);
xnor U26716 (N_26716,N_26385,N_26456);
or U26717 (N_26717,N_26427,N_26417);
and U26718 (N_26718,N_26479,N_26443);
xnor U26719 (N_26719,N_26279,N_26405);
and U26720 (N_26720,N_26366,N_26266);
nand U26721 (N_26721,N_26347,N_26259);
nor U26722 (N_26722,N_26264,N_26371);
nor U26723 (N_26723,N_26407,N_26391);
and U26724 (N_26724,N_26338,N_26289);
or U26725 (N_26725,N_26465,N_26353);
nand U26726 (N_26726,N_26492,N_26335);
nand U26727 (N_26727,N_26369,N_26343);
nor U26728 (N_26728,N_26365,N_26413);
nand U26729 (N_26729,N_26402,N_26319);
and U26730 (N_26730,N_26432,N_26425);
nor U26731 (N_26731,N_26350,N_26487);
nor U26732 (N_26732,N_26348,N_26444);
or U26733 (N_26733,N_26451,N_26327);
nand U26734 (N_26734,N_26451,N_26365);
nand U26735 (N_26735,N_26417,N_26331);
and U26736 (N_26736,N_26343,N_26381);
nor U26737 (N_26737,N_26444,N_26319);
or U26738 (N_26738,N_26453,N_26301);
nor U26739 (N_26739,N_26296,N_26398);
nor U26740 (N_26740,N_26415,N_26277);
and U26741 (N_26741,N_26324,N_26362);
xor U26742 (N_26742,N_26279,N_26389);
nand U26743 (N_26743,N_26329,N_26386);
xnor U26744 (N_26744,N_26343,N_26358);
nand U26745 (N_26745,N_26324,N_26450);
nand U26746 (N_26746,N_26332,N_26279);
and U26747 (N_26747,N_26287,N_26459);
nor U26748 (N_26748,N_26393,N_26253);
and U26749 (N_26749,N_26428,N_26390);
xnor U26750 (N_26750,N_26525,N_26688);
or U26751 (N_26751,N_26509,N_26616);
nor U26752 (N_26752,N_26531,N_26574);
or U26753 (N_26753,N_26579,N_26638);
and U26754 (N_26754,N_26599,N_26520);
nor U26755 (N_26755,N_26503,N_26584);
and U26756 (N_26756,N_26534,N_26566);
nor U26757 (N_26757,N_26643,N_26550);
or U26758 (N_26758,N_26535,N_26749);
nand U26759 (N_26759,N_26596,N_26645);
xor U26760 (N_26760,N_26721,N_26567);
nor U26761 (N_26761,N_26694,N_26555);
nor U26762 (N_26762,N_26601,N_26640);
nand U26763 (N_26763,N_26637,N_26593);
nand U26764 (N_26764,N_26612,N_26678);
and U26765 (N_26765,N_26676,N_26513);
xnor U26766 (N_26766,N_26674,N_26700);
nand U26767 (N_26767,N_26583,N_26528);
nor U26768 (N_26768,N_26727,N_26732);
or U26769 (N_26769,N_26719,N_26679);
nor U26770 (N_26770,N_26667,N_26614);
or U26771 (N_26771,N_26648,N_26551);
and U26772 (N_26772,N_26634,N_26632);
xor U26773 (N_26773,N_26553,N_26661);
nor U26774 (N_26774,N_26742,N_26507);
nand U26775 (N_26775,N_26672,N_26714);
and U26776 (N_26776,N_26627,N_26538);
and U26777 (N_26777,N_26532,N_26666);
xor U26778 (N_26778,N_26728,N_26615);
or U26779 (N_26779,N_26689,N_26501);
nand U26780 (N_26780,N_26620,N_26745);
and U26781 (N_26781,N_26657,N_26682);
xnor U26782 (N_26782,N_26565,N_26647);
and U26783 (N_26783,N_26518,N_26512);
or U26784 (N_26784,N_26548,N_26624);
nand U26785 (N_26785,N_26547,N_26543);
nand U26786 (N_26786,N_26625,N_26602);
xor U26787 (N_26787,N_26686,N_26580);
nand U26788 (N_26788,N_26698,N_26564);
nor U26789 (N_26789,N_26590,N_26709);
nand U26790 (N_26790,N_26663,N_26511);
or U26791 (N_26791,N_26581,N_26633);
xnor U26792 (N_26792,N_26658,N_26635);
nand U26793 (N_26793,N_26636,N_26746);
xnor U26794 (N_26794,N_26716,N_26597);
nor U26795 (N_26795,N_26556,N_26575);
nor U26796 (N_26796,N_26652,N_26655);
nand U26797 (N_26797,N_26649,N_26675);
nand U26798 (N_26798,N_26573,N_26699);
nor U26799 (N_26799,N_26591,N_26603);
nand U26800 (N_26800,N_26702,N_26552);
and U26801 (N_26801,N_26619,N_26631);
xnor U26802 (N_26802,N_26621,N_26641);
nand U26803 (N_26803,N_26696,N_26653);
nand U26804 (N_26804,N_26585,N_26517);
nand U26805 (N_26805,N_26617,N_26740);
nor U26806 (N_26806,N_26669,N_26651);
xor U26807 (N_26807,N_26595,N_26715);
xor U26808 (N_26808,N_26610,N_26527);
or U26809 (N_26809,N_26729,N_26561);
xnor U26810 (N_26810,N_26592,N_26546);
nand U26811 (N_26811,N_26571,N_26560);
nor U26812 (N_26812,N_26735,N_26731);
nand U26813 (N_26813,N_26730,N_26544);
and U26814 (N_26814,N_26650,N_26611);
nor U26815 (N_26815,N_26613,N_26519);
nor U26816 (N_26816,N_26598,N_26588);
nor U26817 (N_26817,N_26521,N_26733);
or U26818 (N_26818,N_26701,N_26662);
xnor U26819 (N_26819,N_26738,N_26541);
or U26820 (N_26820,N_26673,N_26707);
or U26821 (N_26821,N_26505,N_26744);
and U26822 (N_26822,N_26671,N_26572);
nand U26823 (N_26823,N_26708,N_26515);
nand U26824 (N_26824,N_26712,N_26629);
or U26825 (N_26825,N_26609,N_26722);
xor U26826 (N_26826,N_26526,N_26720);
or U26827 (N_26827,N_26705,N_26623);
or U26828 (N_26828,N_26697,N_26710);
xor U26829 (N_26829,N_26604,N_26736);
nor U26830 (N_26830,N_26539,N_26724);
xnor U26831 (N_26831,N_26586,N_26523);
or U26832 (N_26832,N_26514,N_26656);
or U26833 (N_26833,N_26741,N_26606);
and U26834 (N_26834,N_26516,N_26681);
and U26835 (N_26835,N_26578,N_26589);
and U26836 (N_26836,N_26563,N_26660);
nand U26837 (N_26837,N_26542,N_26693);
and U26838 (N_26838,N_26684,N_26510);
and U26839 (N_26839,N_26734,N_26748);
and U26840 (N_26840,N_26659,N_26726);
nand U26841 (N_26841,N_26506,N_26630);
or U26842 (N_26842,N_26607,N_26706);
nand U26843 (N_26843,N_26618,N_26536);
xnor U26844 (N_26844,N_26677,N_26529);
and U26845 (N_26845,N_26522,N_26554);
or U26846 (N_26846,N_26549,N_26703);
nand U26847 (N_26847,N_26644,N_26664);
nand U26848 (N_26848,N_26695,N_26713);
or U26849 (N_26849,N_26557,N_26743);
nor U26850 (N_26850,N_26723,N_26594);
nor U26851 (N_26851,N_26545,N_26622);
nor U26852 (N_26852,N_26605,N_26747);
or U26853 (N_26853,N_26680,N_26508);
nor U26854 (N_26854,N_26502,N_26717);
xnor U26855 (N_26855,N_26577,N_26558);
nor U26856 (N_26856,N_26587,N_26626);
nand U26857 (N_26857,N_26537,N_26540);
xor U26858 (N_26858,N_26582,N_26600);
nor U26859 (N_26859,N_26725,N_26628);
xnor U26860 (N_26860,N_26568,N_26692);
xnor U26861 (N_26861,N_26530,N_26569);
or U26862 (N_26862,N_26737,N_26687);
nor U26863 (N_26863,N_26665,N_26704);
nor U26864 (N_26864,N_26500,N_26570);
nand U26865 (N_26865,N_26668,N_26711);
nor U26866 (N_26866,N_26646,N_26670);
xor U26867 (N_26867,N_26639,N_26576);
and U26868 (N_26868,N_26690,N_26691);
nand U26869 (N_26869,N_26608,N_26642);
and U26870 (N_26870,N_26562,N_26685);
or U26871 (N_26871,N_26739,N_26533);
xor U26872 (N_26872,N_26559,N_26718);
nand U26873 (N_26873,N_26524,N_26504);
or U26874 (N_26874,N_26654,N_26683);
and U26875 (N_26875,N_26739,N_26710);
nand U26876 (N_26876,N_26528,N_26620);
nor U26877 (N_26877,N_26681,N_26662);
and U26878 (N_26878,N_26615,N_26727);
or U26879 (N_26879,N_26563,N_26686);
xnor U26880 (N_26880,N_26637,N_26687);
or U26881 (N_26881,N_26670,N_26552);
or U26882 (N_26882,N_26521,N_26530);
nand U26883 (N_26883,N_26685,N_26746);
nor U26884 (N_26884,N_26730,N_26749);
nand U26885 (N_26885,N_26680,N_26656);
nor U26886 (N_26886,N_26639,N_26520);
xnor U26887 (N_26887,N_26741,N_26698);
or U26888 (N_26888,N_26689,N_26732);
nand U26889 (N_26889,N_26541,N_26666);
nand U26890 (N_26890,N_26662,N_26749);
or U26891 (N_26891,N_26674,N_26516);
or U26892 (N_26892,N_26582,N_26661);
or U26893 (N_26893,N_26639,N_26535);
or U26894 (N_26894,N_26601,N_26646);
xnor U26895 (N_26895,N_26662,N_26536);
and U26896 (N_26896,N_26578,N_26592);
nand U26897 (N_26897,N_26739,N_26732);
nor U26898 (N_26898,N_26708,N_26646);
nand U26899 (N_26899,N_26608,N_26520);
nor U26900 (N_26900,N_26734,N_26746);
nand U26901 (N_26901,N_26534,N_26641);
nand U26902 (N_26902,N_26741,N_26661);
nor U26903 (N_26903,N_26522,N_26580);
nor U26904 (N_26904,N_26737,N_26727);
and U26905 (N_26905,N_26693,N_26680);
nor U26906 (N_26906,N_26722,N_26733);
nor U26907 (N_26907,N_26713,N_26545);
or U26908 (N_26908,N_26501,N_26552);
nor U26909 (N_26909,N_26650,N_26641);
nand U26910 (N_26910,N_26600,N_26695);
and U26911 (N_26911,N_26552,N_26674);
and U26912 (N_26912,N_26634,N_26714);
xor U26913 (N_26913,N_26516,N_26595);
xnor U26914 (N_26914,N_26612,N_26549);
xor U26915 (N_26915,N_26738,N_26655);
xnor U26916 (N_26916,N_26536,N_26554);
nand U26917 (N_26917,N_26535,N_26587);
and U26918 (N_26918,N_26682,N_26662);
or U26919 (N_26919,N_26715,N_26537);
or U26920 (N_26920,N_26626,N_26640);
and U26921 (N_26921,N_26563,N_26564);
nand U26922 (N_26922,N_26601,N_26506);
or U26923 (N_26923,N_26563,N_26749);
and U26924 (N_26924,N_26502,N_26583);
or U26925 (N_26925,N_26506,N_26504);
xor U26926 (N_26926,N_26665,N_26508);
nor U26927 (N_26927,N_26682,N_26707);
nor U26928 (N_26928,N_26701,N_26568);
or U26929 (N_26929,N_26575,N_26724);
nand U26930 (N_26930,N_26529,N_26691);
and U26931 (N_26931,N_26667,N_26615);
nand U26932 (N_26932,N_26594,N_26602);
or U26933 (N_26933,N_26536,N_26611);
nand U26934 (N_26934,N_26500,N_26644);
or U26935 (N_26935,N_26583,N_26563);
nand U26936 (N_26936,N_26659,N_26699);
xnor U26937 (N_26937,N_26657,N_26508);
nor U26938 (N_26938,N_26506,N_26538);
and U26939 (N_26939,N_26741,N_26616);
or U26940 (N_26940,N_26749,N_26616);
xor U26941 (N_26941,N_26553,N_26646);
xor U26942 (N_26942,N_26686,N_26688);
xor U26943 (N_26943,N_26542,N_26640);
nor U26944 (N_26944,N_26579,N_26609);
and U26945 (N_26945,N_26659,N_26572);
and U26946 (N_26946,N_26713,N_26637);
nor U26947 (N_26947,N_26603,N_26597);
nor U26948 (N_26948,N_26532,N_26582);
or U26949 (N_26949,N_26663,N_26567);
nand U26950 (N_26950,N_26549,N_26743);
or U26951 (N_26951,N_26701,N_26549);
and U26952 (N_26952,N_26664,N_26709);
nand U26953 (N_26953,N_26536,N_26682);
nor U26954 (N_26954,N_26518,N_26698);
xor U26955 (N_26955,N_26615,N_26666);
xnor U26956 (N_26956,N_26717,N_26668);
and U26957 (N_26957,N_26585,N_26574);
xnor U26958 (N_26958,N_26665,N_26516);
nand U26959 (N_26959,N_26747,N_26712);
nand U26960 (N_26960,N_26523,N_26542);
and U26961 (N_26961,N_26718,N_26648);
or U26962 (N_26962,N_26727,N_26703);
nand U26963 (N_26963,N_26734,N_26582);
nand U26964 (N_26964,N_26715,N_26590);
and U26965 (N_26965,N_26659,N_26505);
nor U26966 (N_26966,N_26663,N_26627);
nor U26967 (N_26967,N_26714,N_26588);
or U26968 (N_26968,N_26592,N_26628);
or U26969 (N_26969,N_26682,N_26708);
nand U26970 (N_26970,N_26563,N_26524);
and U26971 (N_26971,N_26671,N_26501);
xnor U26972 (N_26972,N_26587,N_26705);
nor U26973 (N_26973,N_26561,N_26626);
and U26974 (N_26974,N_26543,N_26596);
nand U26975 (N_26975,N_26601,N_26681);
and U26976 (N_26976,N_26556,N_26660);
and U26977 (N_26977,N_26596,N_26623);
xnor U26978 (N_26978,N_26727,N_26531);
or U26979 (N_26979,N_26620,N_26726);
xnor U26980 (N_26980,N_26585,N_26614);
nor U26981 (N_26981,N_26601,N_26724);
nand U26982 (N_26982,N_26656,N_26551);
or U26983 (N_26983,N_26588,N_26684);
nand U26984 (N_26984,N_26661,N_26659);
and U26985 (N_26985,N_26676,N_26503);
nor U26986 (N_26986,N_26666,N_26580);
xor U26987 (N_26987,N_26746,N_26680);
nand U26988 (N_26988,N_26730,N_26560);
nor U26989 (N_26989,N_26595,N_26630);
nand U26990 (N_26990,N_26533,N_26682);
nand U26991 (N_26991,N_26578,N_26726);
and U26992 (N_26992,N_26678,N_26549);
nor U26993 (N_26993,N_26656,N_26501);
xor U26994 (N_26994,N_26560,N_26538);
nand U26995 (N_26995,N_26572,N_26622);
xnor U26996 (N_26996,N_26635,N_26645);
nor U26997 (N_26997,N_26742,N_26500);
or U26998 (N_26998,N_26668,N_26509);
or U26999 (N_26999,N_26675,N_26616);
nor U27000 (N_27000,N_26938,N_26978);
nor U27001 (N_27001,N_26961,N_26966);
nor U27002 (N_27002,N_26770,N_26889);
xor U27003 (N_27003,N_26915,N_26766);
and U27004 (N_27004,N_26886,N_26990);
xor U27005 (N_27005,N_26983,N_26795);
nand U27006 (N_27006,N_26758,N_26905);
xor U27007 (N_27007,N_26787,N_26981);
xnor U27008 (N_27008,N_26871,N_26831);
nand U27009 (N_27009,N_26776,N_26971);
nor U27010 (N_27010,N_26959,N_26874);
or U27011 (N_27011,N_26826,N_26888);
xnor U27012 (N_27012,N_26865,N_26877);
nand U27013 (N_27013,N_26750,N_26809);
xor U27014 (N_27014,N_26980,N_26979);
or U27015 (N_27015,N_26753,N_26757);
nor U27016 (N_27016,N_26964,N_26891);
and U27017 (N_27017,N_26863,N_26868);
or U27018 (N_27018,N_26847,N_26939);
or U27019 (N_27019,N_26823,N_26986);
nor U27020 (N_27020,N_26946,N_26968);
or U27021 (N_27021,N_26756,N_26832);
or U27022 (N_27022,N_26783,N_26898);
nand U27023 (N_27023,N_26948,N_26909);
xor U27024 (N_27024,N_26929,N_26907);
nand U27025 (N_27025,N_26772,N_26952);
or U27026 (N_27026,N_26916,N_26880);
nand U27027 (N_27027,N_26890,N_26763);
nor U27028 (N_27028,N_26984,N_26957);
and U27029 (N_27029,N_26860,N_26912);
xnor U27030 (N_27030,N_26872,N_26881);
or U27031 (N_27031,N_26902,N_26820);
or U27032 (N_27032,N_26967,N_26914);
nor U27033 (N_27033,N_26927,N_26822);
and U27034 (N_27034,N_26791,N_26900);
and U27035 (N_27035,N_26834,N_26810);
xor U27036 (N_27036,N_26958,N_26935);
or U27037 (N_27037,N_26879,N_26835);
nor U27038 (N_27038,N_26816,N_26794);
nand U27039 (N_27039,N_26841,N_26975);
and U27040 (N_27040,N_26882,N_26956);
or U27041 (N_27041,N_26796,N_26904);
nor U27042 (N_27042,N_26910,N_26790);
nand U27043 (N_27043,N_26908,N_26911);
nor U27044 (N_27044,N_26942,N_26953);
nand U27045 (N_27045,N_26943,N_26767);
nand U27046 (N_27046,N_26764,N_26875);
xnor U27047 (N_27047,N_26870,N_26901);
xor U27048 (N_27048,N_26784,N_26846);
nand U27049 (N_27049,N_26988,N_26924);
xor U27050 (N_27050,N_26923,N_26827);
nor U27051 (N_27051,N_26782,N_26936);
and U27052 (N_27052,N_26812,N_26960);
nor U27053 (N_27053,N_26857,N_26862);
nor U27054 (N_27054,N_26906,N_26897);
xnor U27055 (N_27055,N_26970,N_26815);
or U27056 (N_27056,N_26840,N_26768);
xor U27057 (N_27057,N_26876,N_26844);
and U27058 (N_27058,N_26937,N_26785);
nor U27059 (N_27059,N_26925,N_26833);
xnor U27060 (N_27060,N_26775,N_26802);
xnor U27061 (N_27061,N_26899,N_26845);
nand U27062 (N_27062,N_26856,N_26913);
nor U27063 (N_27063,N_26761,N_26934);
and U27064 (N_27064,N_26991,N_26853);
xor U27065 (N_27065,N_26931,N_26792);
nand U27066 (N_27066,N_26836,N_26921);
and U27067 (N_27067,N_26837,N_26955);
or U27068 (N_27068,N_26949,N_26779);
and U27069 (N_27069,N_26851,N_26752);
or U27070 (N_27070,N_26962,N_26864);
xnor U27071 (N_27071,N_26850,N_26765);
nand U27072 (N_27072,N_26996,N_26808);
nor U27073 (N_27073,N_26806,N_26965);
nand U27074 (N_27074,N_26974,N_26829);
nor U27075 (N_27075,N_26869,N_26998);
or U27076 (N_27076,N_26895,N_26769);
or U27077 (N_27077,N_26989,N_26892);
nand U27078 (N_27078,N_26963,N_26760);
nor U27079 (N_27079,N_26818,N_26885);
nor U27080 (N_27080,N_26803,N_26976);
nand U27081 (N_27081,N_26788,N_26941);
or U27082 (N_27082,N_26859,N_26954);
xnor U27083 (N_27083,N_26755,N_26993);
and U27084 (N_27084,N_26814,N_26817);
and U27085 (N_27085,N_26842,N_26821);
nor U27086 (N_27086,N_26995,N_26994);
nor U27087 (N_27087,N_26786,N_26855);
and U27088 (N_27088,N_26797,N_26839);
and U27089 (N_27089,N_26798,N_26819);
nand U27090 (N_27090,N_26903,N_26751);
or U27091 (N_27091,N_26781,N_26997);
or U27092 (N_27092,N_26883,N_26922);
nand U27093 (N_27093,N_26973,N_26950);
and U27094 (N_27094,N_26777,N_26945);
nor U27095 (N_27095,N_26754,N_26800);
nand U27096 (N_27096,N_26807,N_26811);
and U27097 (N_27097,N_26838,N_26799);
nand U27098 (N_27098,N_26867,N_26762);
or U27099 (N_27099,N_26932,N_26789);
xor U27100 (N_27100,N_26759,N_26825);
nand U27101 (N_27101,N_26933,N_26848);
nand U27102 (N_27102,N_26917,N_26992);
nand U27103 (N_27103,N_26985,N_26919);
nor U27104 (N_27104,N_26805,N_26824);
nor U27105 (N_27105,N_26930,N_26926);
nor U27106 (N_27106,N_26884,N_26894);
xor U27107 (N_27107,N_26866,N_26896);
nand U27108 (N_27108,N_26947,N_26813);
or U27109 (N_27109,N_26773,N_26982);
and U27110 (N_27110,N_26969,N_26918);
and U27111 (N_27111,N_26804,N_26944);
or U27112 (N_27112,N_26873,N_26828);
or U27113 (N_27113,N_26887,N_26928);
xnor U27114 (N_27114,N_26852,N_26920);
nand U27115 (N_27115,N_26771,N_26893);
nor U27116 (N_27116,N_26972,N_26780);
or U27117 (N_27117,N_26849,N_26878);
and U27118 (N_27118,N_26774,N_26858);
and U27119 (N_27119,N_26778,N_26793);
xor U27120 (N_27120,N_26987,N_26940);
nand U27121 (N_27121,N_26854,N_26861);
and U27122 (N_27122,N_26843,N_26801);
or U27123 (N_27123,N_26830,N_26977);
nor U27124 (N_27124,N_26951,N_26999);
or U27125 (N_27125,N_26804,N_26823);
nand U27126 (N_27126,N_26833,N_26908);
or U27127 (N_27127,N_26866,N_26806);
or U27128 (N_27128,N_26912,N_26956);
or U27129 (N_27129,N_26965,N_26932);
and U27130 (N_27130,N_26850,N_26794);
nand U27131 (N_27131,N_26847,N_26962);
nand U27132 (N_27132,N_26957,N_26828);
nand U27133 (N_27133,N_26948,N_26778);
nor U27134 (N_27134,N_26837,N_26934);
nor U27135 (N_27135,N_26754,N_26825);
and U27136 (N_27136,N_26939,N_26998);
nor U27137 (N_27137,N_26751,N_26817);
and U27138 (N_27138,N_26823,N_26833);
or U27139 (N_27139,N_26858,N_26924);
xnor U27140 (N_27140,N_26794,N_26752);
and U27141 (N_27141,N_26810,N_26887);
xnor U27142 (N_27142,N_26782,N_26978);
xnor U27143 (N_27143,N_26935,N_26874);
and U27144 (N_27144,N_26957,N_26919);
or U27145 (N_27145,N_26858,N_26837);
or U27146 (N_27146,N_26780,N_26913);
xnor U27147 (N_27147,N_26959,N_26819);
nand U27148 (N_27148,N_26890,N_26898);
and U27149 (N_27149,N_26823,N_26776);
and U27150 (N_27150,N_26810,N_26763);
nor U27151 (N_27151,N_26859,N_26809);
nor U27152 (N_27152,N_26940,N_26883);
nor U27153 (N_27153,N_26817,N_26877);
nand U27154 (N_27154,N_26981,N_26950);
and U27155 (N_27155,N_26799,N_26878);
xor U27156 (N_27156,N_26932,N_26984);
nor U27157 (N_27157,N_26981,N_26836);
or U27158 (N_27158,N_26786,N_26960);
or U27159 (N_27159,N_26979,N_26918);
nor U27160 (N_27160,N_26995,N_26754);
nor U27161 (N_27161,N_26768,N_26934);
xnor U27162 (N_27162,N_26761,N_26836);
nor U27163 (N_27163,N_26945,N_26921);
nor U27164 (N_27164,N_26843,N_26778);
xor U27165 (N_27165,N_26890,N_26812);
xor U27166 (N_27166,N_26857,N_26820);
and U27167 (N_27167,N_26798,N_26974);
nand U27168 (N_27168,N_26955,N_26898);
nand U27169 (N_27169,N_26779,N_26826);
or U27170 (N_27170,N_26826,N_26951);
and U27171 (N_27171,N_26869,N_26858);
and U27172 (N_27172,N_26774,N_26869);
and U27173 (N_27173,N_26846,N_26913);
nor U27174 (N_27174,N_26813,N_26755);
and U27175 (N_27175,N_26994,N_26889);
and U27176 (N_27176,N_26899,N_26987);
and U27177 (N_27177,N_26961,N_26875);
xor U27178 (N_27178,N_26949,N_26905);
xor U27179 (N_27179,N_26833,N_26810);
or U27180 (N_27180,N_26959,N_26902);
and U27181 (N_27181,N_26811,N_26935);
nor U27182 (N_27182,N_26867,N_26860);
nor U27183 (N_27183,N_26887,N_26909);
xnor U27184 (N_27184,N_26939,N_26760);
and U27185 (N_27185,N_26807,N_26758);
xnor U27186 (N_27186,N_26877,N_26957);
or U27187 (N_27187,N_26952,N_26806);
xor U27188 (N_27188,N_26950,N_26847);
and U27189 (N_27189,N_26987,N_26802);
nand U27190 (N_27190,N_26791,N_26969);
or U27191 (N_27191,N_26819,N_26836);
or U27192 (N_27192,N_26908,N_26978);
nor U27193 (N_27193,N_26832,N_26827);
or U27194 (N_27194,N_26750,N_26924);
or U27195 (N_27195,N_26940,N_26763);
or U27196 (N_27196,N_26949,N_26968);
xnor U27197 (N_27197,N_26980,N_26797);
nor U27198 (N_27198,N_26984,N_26951);
nand U27199 (N_27199,N_26839,N_26857);
or U27200 (N_27200,N_26865,N_26987);
nand U27201 (N_27201,N_26760,N_26826);
or U27202 (N_27202,N_26945,N_26861);
xor U27203 (N_27203,N_26789,N_26890);
xor U27204 (N_27204,N_26751,N_26967);
xnor U27205 (N_27205,N_26905,N_26839);
xnor U27206 (N_27206,N_26927,N_26832);
or U27207 (N_27207,N_26921,N_26835);
nand U27208 (N_27208,N_26939,N_26944);
nand U27209 (N_27209,N_26865,N_26845);
nand U27210 (N_27210,N_26774,N_26796);
or U27211 (N_27211,N_26872,N_26769);
nor U27212 (N_27212,N_26970,N_26856);
xor U27213 (N_27213,N_26963,N_26984);
or U27214 (N_27214,N_26790,N_26888);
and U27215 (N_27215,N_26885,N_26911);
and U27216 (N_27216,N_26833,N_26861);
xnor U27217 (N_27217,N_26797,N_26915);
or U27218 (N_27218,N_26795,N_26779);
nand U27219 (N_27219,N_26755,N_26980);
nand U27220 (N_27220,N_26987,N_26850);
and U27221 (N_27221,N_26780,N_26959);
xor U27222 (N_27222,N_26758,N_26868);
nand U27223 (N_27223,N_26780,N_26871);
or U27224 (N_27224,N_26780,N_26944);
nor U27225 (N_27225,N_26894,N_26753);
nor U27226 (N_27226,N_26937,N_26921);
nor U27227 (N_27227,N_26957,N_26895);
nor U27228 (N_27228,N_26810,N_26769);
or U27229 (N_27229,N_26764,N_26882);
nor U27230 (N_27230,N_26998,N_26782);
nand U27231 (N_27231,N_26866,N_26939);
and U27232 (N_27232,N_26791,N_26756);
or U27233 (N_27233,N_26831,N_26761);
xnor U27234 (N_27234,N_26952,N_26878);
and U27235 (N_27235,N_26895,N_26826);
nand U27236 (N_27236,N_26810,N_26789);
nor U27237 (N_27237,N_26949,N_26971);
nor U27238 (N_27238,N_26981,N_26941);
nand U27239 (N_27239,N_26936,N_26851);
nand U27240 (N_27240,N_26877,N_26808);
nor U27241 (N_27241,N_26824,N_26943);
xnor U27242 (N_27242,N_26977,N_26989);
nor U27243 (N_27243,N_26854,N_26942);
xor U27244 (N_27244,N_26834,N_26860);
xnor U27245 (N_27245,N_26987,N_26904);
nor U27246 (N_27246,N_26873,N_26933);
and U27247 (N_27247,N_26950,N_26827);
xnor U27248 (N_27248,N_26797,N_26870);
or U27249 (N_27249,N_26966,N_26918);
nand U27250 (N_27250,N_27089,N_27037);
nand U27251 (N_27251,N_27147,N_27148);
nand U27252 (N_27252,N_27129,N_27202);
or U27253 (N_27253,N_27143,N_27080);
nand U27254 (N_27254,N_27170,N_27241);
nor U27255 (N_27255,N_27152,N_27018);
and U27256 (N_27256,N_27087,N_27090);
nand U27257 (N_27257,N_27001,N_27109);
nand U27258 (N_27258,N_27032,N_27052);
nand U27259 (N_27259,N_27222,N_27011);
and U27260 (N_27260,N_27210,N_27104);
nor U27261 (N_27261,N_27248,N_27226);
nand U27262 (N_27262,N_27231,N_27204);
and U27263 (N_27263,N_27043,N_27211);
xnor U27264 (N_27264,N_27091,N_27000);
nand U27265 (N_27265,N_27099,N_27181);
and U27266 (N_27266,N_27137,N_27036);
nor U27267 (N_27267,N_27081,N_27098);
nor U27268 (N_27268,N_27096,N_27111);
nor U27269 (N_27269,N_27200,N_27128);
nor U27270 (N_27270,N_27031,N_27155);
nor U27271 (N_27271,N_27078,N_27165);
or U27272 (N_27272,N_27179,N_27192);
or U27273 (N_27273,N_27088,N_27042);
nor U27274 (N_27274,N_27049,N_27110);
and U27275 (N_27275,N_27033,N_27140);
nand U27276 (N_27276,N_27132,N_27125);
and U27277 (N_27277,N_27063,N_27071);
xor U27278 (N_27278,N_27227,N_27045);
or U27279 (N_27279,N_27188,N_27027);
or U27280 (N_27280,N_27006,N_27105);
nand U27281 (N_27281,N_27159,N_27067);
nand U27282 (N_27282,N_27162,N_27075);
nand U27283 (N_27283,N_27208,N_27223);
xor U27284 (N_27284,N_27100,N_27025);
nor U27285 (N_27285,N_27236,N_27160);
and U27286 (N_27286,N_27176,N_27156);
nand U27287 (N_27287,N_27002,N_27215);
nand U27288 (N_27288,N_27169,N_27057);
and U27289 (N_27289,N_27038,N_27108);
nand U27290 (N_27290,N_27246,N_27219);
xor U27291 (N_27291,N_27154,N_27149);
or U27292 (N_27292,N_27164,N_27103);
nand U27293 (N_27293,N_27083,N_27177);
xnor U27294 (N_27294,N_27190,N_27051);
nand U27295 (N_27295,N_27191,N_27050);
nand U27296 (N_27296,N_27145,N_27058);
and U27297 (N_27297,N_27123,N_27184);
nor U27298 (N_27298,N_27040,N_27174);
nand U27299 (N_27299,N_27186,N_27163);
and U27300 (N_27300,N_27072,N_27126);
or U27301 (N_27301,N_27234,N_27082);
or U27302 (N_27302,N_27112,N_27247);
xor U27303 (N_27303,N_27185,N_27122);
xnor U27304 (N_27304,N_27013,N_27118);
and U27305 (N_27305,N_27238,N_27066);
or U27306 (N_27306,N_27173,N_27114);
nand U27307 (N_27307,N_27245,N_27073);
nand U27308 (N_27308,N_27124,N_27240);
and U27309 (N_27309,N_27133,N_27218);
or U27310 (N_27310,N_27139,N_27022);
and U27311 (N_27311,N_27019,N_27077);
and U27312 (N_27312,N_27230,N_27054);
nand U27313 (N_27313,N_27196,N_27034);
or U27314 (N_27314,N_27180,N_27168);
nand U27315 (N_27315,N_27024,N_27189);
nand U27316 (N_27316,N_27010,N_27209);
nand U27317 (N_27317,N_27171,N_27007);
nand U27318 (N_27318,N_27138,N_27225);
xor U27319 (N_27319,N_27115,N_27203);
xnor U27320 (N_27320,N_27161,N_27061);
nand U27321 (N_27321,N_27249,N_27144);
xnor U27322 (N_27322,N_27199,N_27084);
xor U27323 (N_27323,N_27150,N_27008);
and U27324 (N_27324,N_27229,N_27107);
nor U27325 (N_27325,N_27020,N_27069);
xor U27326 (N_27326,N_27151,N_27182);
and U27327 (N_27327,N_27106,N_27232);
nand U27328 (N_27328,N_27172,N_27135);
xnor U27329 (N_27329,N_27065,N_27092);
nor U27330 (N_27330,N_27060,N_27217);
xnor U27331 (N_27331,N_27064,N_27039);
or U27332 (N_27332,N_27167,N_27243);
or U27333 (N_27333,N_27016,N_27017);
or U27334 (N_27334,N_27004,N_27014);
nor U27335 (N_27335,N_27093,N_27197);
or U27336 (N_27336,N_27198,N_27193);
and U27337 (N_27337,N_27021,N_27213);
and U27338 (N_27338,N_27003,N_27023);
nand U27339 (N_27339,N_27005,N_27194);
or U27340 (N_27340,N_27086,N_27175);
nor U27341 (N_27341,N_27206,N_27074);
nor U27342 (N_27342,N_27195,N_27207);
nand U27343 (N_27343,N_27166,N_27127);
xnor U27344 (N_27344,N_27076,N_27120);
xor U27345 (N_27345,N_27158,N_27233);
or U27346 (N_27346,N_27079,N_27102);
and U27347 (N_27347,N_27047,N_27244);
xnor U27348 (N_27348,N_27153,N_27068);
or U27349 (N_27349,N_27235,N_27015);
nand U27350 (N_27350,N_27239,N_27030);
nor U27351 (N_27351,N_27131,N_27201);
nor U27352 (N_27352,N_27116,N_27187);
and U27353 (N_27353,N_27035,N_27121);
nor U27354 (N_27354,N_27205,N_27183);
or U27355 (N_27355,N_27070,N_27130);
nand U27356 (N_27356,N_27157,N_27048);
nor U27357 (N_27357,N_27041,N_27134);
or U27358 (N_27358,N_27119,N_27237);
or U27359 (N_27359,N_27228,N_27044);
or U27360 (N_27360,N_27146,N_27221);
and U27361 (N_27361,N_27026,N_27056);
or U27362 (N_27362,N_27094,N_27062);
or U27363 (N_27363,N_27113,N_27053);
nor U27364 (N_27364,N_27142,N_27095);
nand U27365 (N_27365,N_27085,N_27097);
xor U27366 (N_27366,N_27216,N_27055);
and U27367 (N_27367,N_27009,N_27212);
or U27368 (N_27368,N_27220,N_27046);
or U27369 (N_27369,N_27117,N_27224);
and U27370 (N_27370,N_27136,N_27012);
nor U27371 (N_27371,N_27141,N_27028);
nor U27372 (N_27372,N_27029,N_27101);
xor U27373 (N_27373,N_27059,N_27214);
and U27374 (N_27374,N_27178,N_27242);
xor U27375 (N_27375,N_27188,N_27065);
xor U27376 (N_27376,N_27082,N_27180);
nand U27377 (N_27377,N_27178,N_27241);
and U27378 (N_27378,N_27118,N_27151);
or U27379 (N_27379,N_27142,N_27068);
xor U27380 (N_27380,N_27066,N_27032);
nand U27381 (N_27381,N_27207,N_27068);
nand U27382 (N_27382,N_27157,N_27180);
nand U27383 (N_27383,N_27028,N_27134);
xnor U27384 (N_27384,N_27119,N_27245);
or U27385 (N_27385,N_27193,N_27107);
and U27386 (N_27386,N_27019,N_27164);
nor U27387 (N_27387,N_27200,N_27142);
xor U27388 (N_27388,N_27150,N_27016);
and U27389 (N_27389,N_27089,N_27095);
nor U27390 (N_27390,N_27068,N_27245);
xor U27391 (N_27391,N_27065,N_27052);
nor U27392 (N_27392,N_27171,N_27162);
nand U27393 (N_27393,N_27037,N_27238);
xor U27394 (N_27394,N_27094,N_27246);
nand U27395 (N_27395,N_27228,N_27054);
nor U27396 (N_27396,N_27157,N_27000);
and U27397 (N_27397,N_27052,N_27078);
nand U27398 (N_27398,N_27158,N_27084);
nor U27399 (N_27399,N_27084,N_27015);
and U27400 (N_27400,N_27056,N_27097);
or U27401 (N_27401,N_27144,N_27099);
nand U27402 (N_27402,N_27215,N_27210);
and U27403 (N_27403,N_27129,N_27030);
xor U27404 (N_27404,N_27014,N_27176);
or U27405 (N_27405,N_27219,N_27068);
xor U27406 (N_27406,N_27068,N_27152);
nor U27407 (N_27407,N_27010,N_27092);
nor U27408 (N_27408,N_27150,N_27110);
xor U27409 (N_27409,N_27131,N_27030);
nand U27410 (N_27410,N_27028,N_27081);
nor U27411 (N_27411,N_27090,N_27164);
nand U27412 (N_27412,N_27042,N_27031);
and U27413 (N_27413,N_27048,N_27190);
or U27414 (N_27414,N_27101,N_27178);
xnor U27415 (N_27415,N_27176,N_27158);
nor U27416 (N_27416,N_27056,N_27043);
nor U27417 (N_27417,N_27174,N_27025);
xor U27418 (N_27418,N_27077,N_27113);
xor U27419 (N_27419,N_27097,N_27145);
and U27420 (N_27420,N_27179,N_27194);
and U27421 (N_27421,N_27167,N_27068);
nand U27422 (N_27422,N_27106,N_27121);
xor U27423 (N_27423,N_27143,N_27214);
and U27424 (N_27424,N_27079,N_27168);
and U27425 (N_27425,N_27243,N_27046);
nand U27426 (N_27426,N_27157,N_27243);
xnor U27427 (N_27427,N_27228,N_27206);
or U27428 (N_27428,N_27044,N_27018);
nand U27429 (N_27429,N_27167,N_27049);
nor U27430 (N_27430,N_27079,N_27011);
nand U27431 (N_27431,N_27227,N_27144);
or U27432 (N_27432,N_27166,N_27219);
xnor U27433 (N_27433,N_27059,N_27119);
nand U27434 (N_27434,N_27176,N_27146);
or U27435 (N_27435,N_27223,N_27155);
xnor U27436 (N_27436,N_27082,N_27193);
nand U27437 (N_27437,N_27085,N_27060);
xor U27438 (N_27438,N_27229,N_27086);
and U27439 (N_27439,N_27216,N_27207);
or U27440 (N_27440,N_27076,N_27117);
or U27441 (N_27441,N_27059,N_27222);
nand U27442 (N_27442,N_27212,N_27022);
nor U27443 (N_27443,N_27058,N_27190);
xnor U27444 (N_27444,N_27177,N_27118);
xnor U27445 (N_27445,N_27129,N_27159);
nand U27446 (N_27446,N_27060,N_27210);
nor U27447 (N_27447,N_27211,N_27018);
xor U27448 (N_27448,N_27115,N_27134);
nand U27449 (N_27449,N_27122,N_27087);
nor U27450 (N_27450,N_27005,N_27162);
or U27451 (N_27451,N_27240,N_27028);
nor U27452 (N_27452,N_27213,N_27168);
or U27453 (N_27453,N_27086,N_27084);
nand U27454 (N_27454,N_27003,N_27123);
or U27455 (N_27455,N_27091,N_27149);
nand U27456 (N_27456,N_27233,N_27080);
or U27457 (N_27457,N_27156,N_27048);
or U27458 (N_27458,N_27055,N_27169);
nand U27459 (N_27459,N_27057,N_27231);
and U27460 (N_27460,N_27070,N_27101);
xnor U27461 (N_27461,N_27023,N_27249);
nor U27462 (N_27462,N_27244,N_27185);
or U27463 (N_27463,N_27071,N_27114);
and U27464 (N_27464,N_27096,N_27009);
xnor U27465 (N_27465,N_27000,N_27011);
and U27466 (N_27466,N_27202,N_27010);
or U27467 (N_27467,N_27248,N_27015);
or U27468 (N_27468,N_27156,N_27007);
xor U27469 (N_27469,N_27179,N_27121);
xor U27470 (N_27470,N_27035,N_27236);
or U27471 (N_27471,N_27050,N_27031);
xor U27472 (N_27472,N_27080,N_27015);
nand U27473 (N_27473,N_27003,N_27163);
and U27474 (N_27474,N_27096,N_27021);
nor U27475 (N_27475,N_27034,N_27222);
and U27476 (N_27476,N_27094,N_27078);
nand U27477 (N_27477,N_27224,N_27025);
xor U27478 (N_27478,N_27102,N_27080);
nor U27479 (N_27479,N_27115,N_27030);
xnor U27480 (N_27480,N_27211,N_27157);
xnor U27481 (N_27481,N_27233,N_27172);
and U27482 (N_27482,N_27049,N_27093);
xnor U27483 (N_27483,N_27138,N_27153);
nor U27484 (N_27484,N_27243,N_27042);
xor U27485 (N_27485,N_27237,N_27062);
xnor U27486 (N_27486,N_27139,N_27133);
or U27487 (N_27487,N_27231,N_27121);
and U27488 (N_27488,N_27128,N_27193);
or U27489 (N_27489,N_27113,N_27241);
or U27490 (N_27490,N_27151,N_27128);
and U27491 (N_27491,N_27080,N_27189);
nor U27492 (N_27492,N_27081,N_27027);
xnor U27493 (N_27493,N_27077,N_27159);
xnor U27494 (N_27494,N_27032,N_27153);
nor U27495 (N_27495,N_27149,N_27075);
and U27496 (N_27496,N_27038,N_27128);
nand U27497 (N_27497,N_27102,N_27166);
or U27498 (N_27498,N_27203,N_27095);
or U27499 (N_27499,N_27055,N_27033);
and U27500 (N_27500,N_27385,N_27355);
nor U27501 (N_27501,N_27456,N_27361);
xnor U27502 (N_27502,N_27419,N_27283);
xor U27503 (N_27503,N_27449,N_27400);
xor U27504 (N_27504,N_27371,N_27286);
nand U27505 (N_27505,N_27434,N_27433);
nand U27506 (N_27506,N_27308,N_27478);
nor U27507 (N_27507,N_27324,N_27275);
nor U27508 (N_27508,N_27437,N_27289);
nand U27509 (N_27509,N_27299,N_27326);
xor U27510 (N_27510,N_27392,N_27423);
xnor U27511 (N_27511,N_27421,N_27332);
nand U27512 (N_27512,N_27390,N_27397);
xor U27513 (N_27513,N_27328,N_27269);
nor U27514 (N_27514,N_27325,N_27410);
xor U27515 (N_27515,N_27473,N_27462);
nand U27516 (N_27516,N_27300,N_27295);
and U27517 (N_27517,N_27448,N_27458);
or U27518 (N_27518,N_27352,N_27364);
xnor U27519 (N_27519,N_27321,N_27468);
and U27520 (N_27520,N_27431,N_27335);
xnor U27521 (N_27521,N_27271,N_27329);
and U27522 (N_27522,N_27469,N_27402);
nor U27523 (N_27523,N_27334,N_27253);
or U27524 (N_27524,N_27342,N_27406);
xor U27525 (N_27525,N_27305,N_27409);
nor U27526 (N_27526,N_27493,N_27333);
nor U27527 (N_27527,N_27454,N_27327);
and U27528 (N_27528,N_27272,N_27280);
or U27529 (N_27529,N_27441,N_27340);
nand U27530 (N_27530,N_27386,N_27401);
xnor U27531 (N_27531,N_27360,N_27389);
or U27532 (N_27532,N_27293,N_27398);
nand U27533 (N_27533,N_27311,N_27339);
and U27534 (N_27534,N_27396,N_27378);
and U27535 (N_27535,N_27315,N_27276);
nand U27536 (N_27536,N_27277,N_27250);
xnor U27537 (N_27537,N_27351,N_27413);
or U27538 (N_27538,N_27480,N_27257);
xnor U27539 (N_27539,N_27499,N_27363);
nor U27540 (N_27540,N_27347,N_27306);
and U27541 (N_27541,N_27407,N_27452);
nor U27542 (N_27542,N_27376,N_27255);
or U27543 (N_27543,N_27393,N_27297);
xnor U27544 (N_27544,N_27345,N_27470);
nand U27545 (N_27545,N_27415,N_27443);
nor U27546 (N_27546,N_27490,N_27476);
and U27547 (N_27547,N_27284,N_27404);
or U27548 (N_27548,N_27254,N_27318);
or U27549 (N_27549,N_27491,N_27313);
nor U27550 (N_27550,N_27445,N_27348);
nand U27551 (N_27551,N_27258,N_27270);
nand U27552 (N_27552,N_27304,N_27358);
nor U27553 (N_27553,N_27291,N_27472);
or U27554 (N_27554,N_27440,N_27294);
nand U27555 (N_27555,N_27338,N_27412);
and U27556 (N_27556,N_27420,N_27290);
nand U27557 (N_27557,N_27354,N_27450);
xnor U27558 (N_27558,N_27282,N_27482);
or U27559 (N_27559,N_27455,N_27251);
xor U27560 (N_27560,N_27343,N_27486);
xor U27561 (N_27561,N_27461,N_27395);
and U27562 (N_27562,N_27488,N_27307);
nand U27563 (N_27563,N_27375,N_27274);
nand U27564 (N_27564,N_27383,N_27467);
nand U27565 (N_27565,N_27322,N_27356);
and U27566 (N_27566,N_27463,N_27384);
and U27567 (N_27567,N_27439,N_27436);
xor U27568 (N_27568,N_27372,N_27273);
or U27569 (N_27569,N_27496,N_27310);
nand U27570 (N_27570,N_27362,N_27391);
and U27571 (N_27571,N_27466,N_27465);
and U27572 (N_27572,N_27316,N_27483);
and U27573 (N_27573,N_27494,N_27288);
nand U27574 (N_27574,N_27424,N_27459);
nor U27575 (N_27575,N_27414,N_27314);
nand U27576 (N_27576,N_27312,N_27319);
xnor U27577 (N_27577,N_27377,N_27349);
xnor U27578 (N_27578,N_27485,N_27418);
and U27579 (N_27579,N_27408,N_27266);
or U27580 (N_27580,N_27320,N_27498);
or U27581 (N_27581,N_27484,N_27460);
or U27582 (N_27582,N_27474,N_27353);
and U27583 (N_27583,N_27442,N_27481);
and U27584 (N_27584,N_27438,N_27428);
or U27585 (N_27585,N_27479,N_27337);
nor U27586 (N_27586,N_27411,N_27366);
or U27587 (N_27587,N_27487,N_27264);
or U27588 (N_27588,N_27350,N_27367);
or U27589 (N_27589,N_27489,N_27259);
xnor U27590 (N_27590,N_27256,N_27477);
xor U27591 (N_27591,N_27451,N_27471);
nor U27592 (N_27592,N_27382,N_27262);
nor U27593 (N_27593,N_27444,N_27296);
and U27594 (N_27594,N_27399,N_27427);
or U27595 (N_27595,N_27475,N_27403);
nand U27596 (N_27596,N_27330,N_27301);
xnor U27597 (N_27597,N_27446,N_27373);
and U27598 (N_27598,N_27380,N_27394);
nor U27599 (N_27599,N_27359,N_27422);
and U27600 (N_27600,N_27344,N_27292);
nor U27601 (N_27601,N_27425,N_27252);
xor U27602 (N_27602,N_27495,N_27265);
or U27603 (N_27603,N_27369,N_27260);
and U27604 (N_27604,N_27303,N_27374);
or U27605 (N_27605,N_27298,N_27492);
nor U27606 (N_27606,N_27357,N_27268);
nor U27607 (N_27607,N_27336,N_27346);
xnor U27608 (N_27608,N_27464,N_27281);
nor U27609 (N_27609,N_27368,N_27279);
xnor U27610 (N_27610,N_27278,N_27430);
or U27611 (N_27611,N_27453,N_27435);
nand U27612 (N_27612,N_27287,N_27417);
nand U27613 (N_27613,N_27457,N_27309);
nor U27614 (N_27614,N_27416,N_27432);
nor U27615 (N_27615,N_27317,N_27261);
nand U27616 (N_27616,N_27405,N_27379);
xnor U27617 (N_27617,N_27302,N_27370);
nor U27618 (N_27618,N_27365,N_27381);
nand U27619 (N_27619,N_27387,N_27285);
and U27620 (N_27620,N_27263,N_27497);
nand U27621 (N_27621,N_27429,N_27388);
xnor U27622 (N_27622,N_27323,N_27267);
nand U27623 (N_27623,N_27341,N_27447);
xnor U27624 (N_27624,N_27331,N_27426);
nor U27625 (N_27625,N_27491,N_27346);
nand U27626 (N_27626,N_27417,N_27433);
nand U27627 (N_27627,N_27391,N_27289);
or U27628 (N_27628,N_27274,N_27266);
or U27629 (N_27629,N_27300,N_27450);
nand U27630 (N_27630,N_27334,N_27386);
and U27631 (N_27631,N_27306,N_27318);
xnor U27632 (N_27632,N_27345,N_27428);
nand U27633 (N_27633,N_27361,N_27467);
or U27634 (N_27634,N_27496,N_27464);
nor U27635 (N_27635,N_27321,N_27355);
xor U27636 (N_27636,N_27273,N_27427);
nand U27637 (N_27637,N_27389,N_27377);
nand U27638 (N_27638,N_27268,N_27426);
xor U27639 (N_27639,N_27403,N_27269);
xnor U27640 (N_27640,N_27402,N_27292);
nor U27641 (N_27641,N_27343,N_27443);
nand U27642 (N_27642,N_27452,N_27398);
nor U27643 (N_27643,N_27256,N_27276);
nor U27644 (N_27644,N_27394,N_27473);
xor U27645 (N_27645,N_27440,N_27481);
nor U27646 (N_27646,N_27496,N_27329);
xor U27647 (N_27647,N_27366,N_27456);
or U27648 (N_27648,N_27288,N_27318);
xor U27649 (N_27649,N_27450,N_27333);
nand U27650 (N_27650,N_27451,N_27303);
nand U27651 (N_27651,N_27414,N_27292);
xnor U27652 (N_27652,N_27407,N_27314);
nor U27653 (N_27653,N_27472,N_27446);
xnor U27654 (N_27654,N_27314,N_27494);
nand U27655 (N_27655,N_27462,N_27443);
xnor U27656 (N_27656,N_27417,N_27447);
or U27657 (N_27657,N_27329,N_27322);
and U27658 (N_27658,N_27383,N_27492);
and U27659 (N_27659,N_27435,N_27312);
or U27660 (N_27660,N_27305,N_27355);
and U27661 (N_27661,N_27410,N_27304);
or U27662 (N_27662,N_27360,N_27458);
nor U27663 (N_27663,N_27450,N_27430);
nor U27664 (N_27664,N_27298,N_27326);
or U27665 (N_27665,N_27359,N_27477);
xor U27666 (N_27666,N_27495,N_27334);
xor U27667 (N_27667,N_27371,N_27469);
xor U27668 (N_27668,N_27405,N_27479);
xnor U27669 (N_27669,N_27266,N_27364);
nor U27670 (N_27670,N_27251,N_27472);
and U27671 (N_27671,N_27433,N_27366);
nand U27672 (N_27672,N_27417,N_27424);
nand U27673 (N_27673,N_27329,N_27252);
nor U27674 (N_27674,N_27359,N_27309);
xor U27675 (N_27675,N_27282,N_27315);
xnor U27676 (N_27676,N_27407,N_27356);
xnor U27677 (N_27677,N_27436,N_27451);
or U27678 (N_27678,N_27286,N_27258);
nor U27679 (N_27679,N_27292,N_27342);
and U27680 (N_27680,N_27372,N_27354);
and U27681 (N_27681,N_27317,N_27432);
and U27682 (N_27682,N_27274,N_27271);
nand U27683 (N_27683,N_27269,N_27415);
xnor U27684 (N_27684,N_27497,N_27341);
xor U27685 (N_27685,N_27253,N_27333);
nor U27686 (N_27686,N_27493,N_27361);
xnor U27687 (N_27687,N_27331,N_27497);
nor U27688 (N_27688,N_27383,N_27414);
and U27689 (N_27689,N_27339,N_27361);
xor U27690 (N_27690,N_27469,N_27272);
nor U27691 (N_27691,N_27415,N_27484);
nand U27692 (N_27692,N_27335,N_27403);
nor U27693 (N_27693,N_27391,N_27258);
or U27694 (N_27694,N_27296,N_27360);
or U27695 (N_27695,N_27475,N_27351);
or U27696 (N_27696,N_27394,N_27295);
nand U27697 (N_27697,N_27463,N_27415);
or U27698 (N_27698,N_27295,N_27372);
nor U27699 (N_27699,N_27346,N_27310);
nor U27700 (N_27700,N_27396,N_27328);
nor U27701 (N_27701,N_27452,N_27291);
nand U27702 (N_27702,N_27366,N_27498);
nor U27703 (N_27703,N_27499,N_27479);
xnor U27704 (N_27704,N_27328,N_27453);
and U27705 (N_27705,N_27443,N_27440);
xor U27706 (N_27706,N_27281,N_27384);
or U27707 (N_27707,N_27485,N_27390);
nand U27708 (N_27708,N_27386,N_27345);
xor U27709 (N_27709,N_27425,N_27437);
or U27710 (N_27710,N_27483,N_27337);
nor U27711 (N_27711,N_27435,N_27284);
and U27712 (N_27712,N_27284,N_27363);
nand U27713 (N_27713,N_27280,N_27287);
xnor U27714 (N_27714,N_27283,N_27260);
or U27715 (N_27715,N_27259,N_27380);
or U27716 (N_27716,N_27338,N_27339);
nand U27717 (N_27717,N_27301,N_27391);
xor U27718 (N_27718,N_27400,N_27374);
nand U27719 (N_27719,N_27455,N_27487);
nor U27720 (N_27720,N_27300,N_27435);
or U27721 (N_27721,N_27429,N_27330);
nor U27722 (N_27722,N_27458,N_27412);
nand U27723 (N_27723,N_27274,N_27252);
or U27724 (N_27724,N_27332,N_27302);
or U27725 (N_27725,N_27372,N_27471);
nor U27726 (N_27726,N_27320,N_27259);
nand U27727 (N_27727,N_27477,N_27381);
and U27728 (N_27728,N_27350,N_27262);
and U27729 (N_27729,N_27439,N_27323);
xor U27730 (N_27730,N_27368,N_27369);
and U27731 (N_27731,N_27303,N_27320);
and U27732 (N_27732,N_27421,N_27368);
nand U27733 (N_27733,N_27479,N_27278);
nand U27734 (N_27734,N_27461,N_27319);
and U27735 (N_27735,N_27421,N_27319);
nor U27736 (N_27736,N_27334,N_27491);
nand U27737 (N_27737,N_27255,N_27372);
xor U27738 (N_27738,N_27273,N_27295);
or U27739 (N_27739,N_27450,N_27474);
nor U27740 (N_27740,N_27436,N_27307);
xor U27741 (N_27741,N_27390,N_27401);
xnor U27742 (N_27742,N_27341,N_27378);
nor U27743 (N_27743,N_27494,N_27491);
nor U27744 (N_27744,N_27301,N_27325);
and U27745 (N_27745,N_27477,N_27292);
and U27746 (N_27746,N_27465,N_27273);
nor U27747 (N_27747,N_27445,N_27420);
or U27748 (N_27748,N_27360,N_27432);
nor U27749 (N_27749,N_27377,N_27422);
or U27750 (N_27750,N_27561,N_27514);
xnor U27751 (N_27751,N_27716,N_27629);
or U27752 (N_27752,N_27733,N_27671);
and U27753 (N_27753,N_27732,N_27618);
and U27754 (N_27754,N_27515,N_27516);
nor U27755 (N_27755,N_27533,N_27700);
xnor U27756 (N_27756,N_27593,N_27710);
and U27757 (N_27757,N_27506,N_27695);
xor U27758 (N_27758,N_27510,N_27678);
nor U27759 (N_27759,N_27699,N_27508);
nand U27760 (N_27760,N_27702,N_27646);
or U27761 (N_27761,N_27609,N_27685);
nand U27762 (N_27762,N_27590,N_27651);
or U27763 (N_27763,N_27635,N_27610);
and U27764 (N_27764,N_27626,N_27604);
xor U27765 (N_27765,N_27743,N_27689);
nand U27766 (N_27766,N_27624,N_27595);
xnor U27767 (N_27767,N_27535,N_27569);
xnor U27768 (N_27768,N_27532,N_27547);
nor U27769 (N_27769,N_27589,N_27641);
or U27770 (N_27770,N_27501,N_27705);
nor U27771 (N_27771,N_27513,N_27548);
nor U27772 (N_27772,N_27742,N_27544);
or U27773 (N_27773,N_27542,N_27679);
nor U27774 (N_27774,N_27594,N_27658);
or U27775 (N_27775,N_27541,N_27718);
nand U27776 (N_27776,N_27522,N_27579);
or U27777 (N_27777,N_27656,N_27586);
or U27778 (N_27778,N_27562,N_27555);
or U27779 (N_27779,N_27625,N_27676);
nor U27780 (N_27780,N_27713,N_27525);
and U27781 (N_27781,N_27712,N_27729);
xnor U27782 (N_27782,N_27583,N_27709);
xor U27783 (N_27783,N_27740,N_27736);
and U27784 (N_27784,N_27645,N_27636);
nor U27785 (N_27785,N_27719,N_27615);
xor U27786 (N_27786,N_27563,N_27691);
or U27787 (N_27787,N_27576,N_27673);
and U27788 (N_27788,N_27597,N_27505);
or U27789 (N_27789,N_27520,N_27644);
nor U27790 (N_27790,N_27581,N_27662);
xnor U27791 (N_27791,N_27580,N_27613);
nor U27792 (N_27792,N_27741,N_27665);
or U27793 (N_27793,N_27703,N_27731);
nand U27794 (N_27794,N_27694,N_27565);
nand U27795 (N_27795,N_27526,N_27707);
nor U27796 (N_27796,N_27577,N_27518);
or U27797 (N_27797,N_27529,N_27603);
or U27798 (N_27798,N_27749,N_27727);
nand U27799 (N_27799,N_27531,N_27682);
nor U27800 (N_27800,N_27660,N_27500);
and U27801 (N_27801,N_27728,N_27666);
xnor U27802 (N_27802,N_27557,N_27623);
xnor U27803 (N_27803,N_27642,N_27628);
nor U27804 (N_27804,N_27524,N_27551);
or U27805 (N_27805,N_27739,N_27670);
or U27806 (N_27806,N_27746,N_27503);
nor U27807 (N_27807,N_27643,N_27621);
nor U27808 (N_27808,N_27616,N_27509);
and U27809 (N_27809,N_27546,N_27737);
nand U27810 (N_27810,N_27714,N_27744);
nor U27811 (N_27811,N_27654,N_27745);
or U27812 (N_27812,N_27564,N_27725);
or U27813 (N_27813,N_27696,N_27688);
nor U27814 (N_27814,N_27521,N_27686);
or U27815 (N_27815,N_27596,N_27652);
and U27816 (N_27816,N_27647,N_27704);
and U27817 (N_27817,N_27748,N_27669);
or U27818 (N_27818,N_27684,N_27722);
nor U27819 (N_27819,N_27553,N_27552);
xor U27820 (N_27820,N_27587,N_27661);
xor U27821 (N_27821,N_27664,N_27608);
and U27822 (N_27822,N_27734,N_27517);
and U27823 (N_27823,N_27598,N_27692);
and U27824 (N_27824,N_27730,N_27549);
or U27825 (N_27825,N_27599,N_27721);
and U27826 (N_27826,N_27674,N_27659);
xor U27827 (N_27827,N_27578,N_27631);
nor U27828 (N_27828,N_27675,N_27648);
or U27829 (N_27829,N_27637,N_27554);
xor U27830 (N_27830,N_27627,N_27698);
xor U27831 (N_27831,N_27612,N_27680);
and U27832 (N_27832,N_27512,N_27536);
and U27833 (N_27833,N_27558,N_27523);
and U27834 (N_27834,N_27632,N_27572);
xnor U27835 (N_27835,N_27573,N_27735);
nand U27836 (N_27836,N_27630,N_27534);
nand U27837 (N_27837,N_27708,N_27622);
and U27838 (N_27838,N_27527,N_27607);
nor U27839 (N_27839,N_27556,N_27693);
and U27840 (N_27840,N_27575,N_27639);
nor U27841 (N_27841,N_27584,N_27677);
xnor U27842 (N_27842,N_27697,N_27657);
nand U27843 (N_27843,N_27605,N_27570);
xor U27844 (N_27844,N_27653,N_27611);
nand U27845 (N_27845,N_27747,N_27614);
nand U27846 (N_27846,N_27687,N_27540);
nor U27847 (N_27847,N_27530,N_27550);
xnor U27848 (N_27848,N_27667,N_27668);
and U27849 (N_27849,N_27711,N_27568);
xor U27850 (N_27850,N_27726,N_27507);
xnor U27851 (N_27851,N_27619,N_27502);
xnor U27852 (N_27852,N_27592,N_27591);
xor U27853 (N_27853,N_27620,N_27617);
and U27854 (N_27854,N_27640,N_27638);
and U27855 (N_27855,N_27574,N_27566);
or U27856 (N_27856,N_27602,N_27601);
xnor U27857 (N_27857,N_27519,N_27571);
or U27858 (N_27858,N_27738,N_27582);
or U27859 (N_27859,N_27606,N_27655);
and U27860 (N_27860,N_27633,N_27723);
xor U27861 (N_27861,N_27683,N_27634);
or U27862 (N_27862,N_27706,N_27717);
nand U27863 (N_27863,N_27649,N_27539);
xnor U27864 (N_27864,N_27681,N_27504);
or U27865 (N_27865,N_27701,N_27538);
xor U27866 (N_27866,N_27585,N_27724);
or U27867 (N_27867,N_27690,N_27663);
nand U27868 (N_27868,N_27720,N_27567);
nor U27869 (N_27869,N_27672,N_27560);
and U27870 (N_27870,N_27715,N_27543);
or U27871 (N_27871,N_27600,N_27537);
xor U27872 (N_27872,N_27511,N_27650);
nor U27873 (N_27873,N_27545,N_27588);
or U27874 (N_27874,N_27528,N_27559);
nor U27875 (N_27875,N_27585,N_27749);
or U27876 (N_27876,N_27698,N_27633);
and U27877 (N_27877,N_27697,N_27609);
xor U27878 (N_27878,N_27620,N_27676);
xnor U27879 (N_27879,N_27520,N_27659);
xor U27880 (N_27880,N_27565,N_27517);
and U27881 (N_27881,N_27708,N_27648);
nor U27882 (N_27882,N_27705,N_27606);
and U27883 (N_27883,N_27566,N_27545);
and U27884 (N_27884,N_27711,N_27741);
nor U27885 (N_27885,N_27680,N_27640);
xnor U27886 (N_27886,N_27607,N_27654);
nand U27887 (N_27887,N_27664,N_27596);
and U27888 (N_27888,N_27618,N_27709);
nor U27889 (N_27889,N_27600,N_27586);
and U27890 (N_27890,N_27652,N_27737);
nor U27891 (N_27891,N_27703,N_27689);
and U27892 (N_27892,N_27577,N_27631);
or U27893 (N_27893,N_27630,N_27603);
xnor U27894 (N_27894,N_27623,N_27591);
nand U27895 (N_27895,N_27637,N_27619);
nor U27896 (N_27896,N_27735,N_27691);
nor U27897 (N_27897,N_27675,N_27542);
and U27898 (N_27898,N_27713,N_27539);
or U27899 (N_27899,N_27745,N_27719);
xnor U27900 (N_27900,N_27622,N_27597);
xor U27901 (N_27901,N_27549,N_27576);
nand U27902 (N_27902,N_27748,N_27519);
or U27903 (N_27903,N_27544,N_27711);
xnor U27904 (N_27904,N_27618,N_27510);
or U27905 (N_27905,N_27566,N_27704);
nor U27906 (N_27906,N_27523,N_27704);
or U27907 (N_27907,N_27517,N_27707);
nand U27908 (N_27908,N_27716,N_27684);
or U27909 (N_27909,N_27745,N_27678);
nand U27910 (N_27910,N_27665,N_27585);
nor U27911 (N_27911,N_27652,N_27638);
xor U27912 (N_27912,N_27526,N_27704);
or U27913 (N_27913,N_27530,N_27713);
and U27914 (N_27914,N_27651,N_27692);
and U27915 (N_27915,N_27640,N_27553);
or U27916 (N_27916,N_27572,N_27610);
and U27917 (N_27917,N_27531,N_27624);
or U27918 (N_27918,N_27723,N_27711);
or U27919 (N_27919,N_27570,N_27574);
and U27920 (N_27920,N_27748,N_27581);
and U27921 (N_27921,N_27629,N_27678);
nand U27922 (N_27922,N_27530,N_27739);
and U27923 (N_27923,N_27510,N_27550);
or U27924 (N_27924,N_27595,N_27533);
xnor U27925 (N_27925,N_27527,N_27723);
nand U27926 (N_27926,N_27545,N_27647);
nand U27927 (N_27927,N_27637,N_27536);
or U27928 (N_27928,N_27746,N_27549);
xnor U27929 (N_27929,N_27726,N_27642);
and U27930 (N_27930,N_27514,N_27608);
nor U27931 (N_27931,N_27583,N_27582);
nand U27932 (N_27932,N_27683,N_27731);
and U27933 (N_27933,N_27585,N_27712);
and U27934 (N_27934,N_27534,N_27542);
xor U27935 (N_27935,N_27509,N_27703);
nor U27936 (N_27936,N_27602,N_27598);
nor U27937 (N_27937,N_27682,N_27721);
or U27938 (N_27938,N_27702,N_27531);
nand U27939 (N_27939,N_27651,N_27536);
nor U27940 (N_27940,N_27561,N_27553);
nor U27941 (N_27941,N_27742,N_27500);
xnor U27942 (N_27942,N_27607,N_27508);
nor U27943 (N_27943,N_27678,N_27618);
nand U27944 (N_27944,N_27511,N_27516);
xor U27945 (N_27945,N_27502,N_27581);
or U27946 (N_27946,N_27614,N_27687);
and U27947 (N_27947,N_27635,N_27625);
and U27948 (N_27948,N_27552,N_27501);
nand U27949 (N_27949,N_27607,N_27611);
xnor U27950 (N_27950,N_27516,N_27595);
nand U27951 (N_27951,N_27664,N_27723);
nor U27952 (N_27952,N_27624,N_27530);
xnor U27953 (N_27953,N_27515,N_27687);
nor U27954 (N_27954,N_27708,N_27692);
nand U27955 (N_27955,N_27511,N_27740);
xnor U27956 (N_27956,N_27607,N_27681);
nand U27957 (N_27957,N_27572,N_27739);
xor U27958 (N_27958,N_27522,N_27558);
nand U27959 (N_27959,N_27527,N_27594);
and U27960 (N_27960,N_27717,N_27732);
and U27961 (N_27961,N_27561,N_27509);
nor U27962 (N_27962,N_27728,N_27725);
nand U27963 (N_27963,N_27579,N_27578);
xnor U27964 (N_27964,N_27506,N_27532);
nor U27965 (N_27965,N_27685,N_27644);
and U27966 (N_27966,N_27743,N_27562);
or U27967 (N_27967,N_27543,N_27574);
and U27968 (N_27968,N_27689,N_27724);
and U27969 (N_27969,N_27716,N_27682);
nor U27970 (N_27970,N_27744,N_27595);
and U27971 (N_27971,N_27656,N_27715);
nand U27972 (N_27972,N_27626,N_27557);
xnor U27973 (N_27973,N_27581,N_27562);
xnor U27974 (N_27974,N_27730,N_27637);
nand U27975 (N_27975,N_27535,N_27595);
or U27976 (N_27976,N_27615,N_27729);
and U27977 (N_27977,N_27643,N_27569);
xor U27978 (N_27978,N_27664,N_27557);
nand U27979 (N_27979,N_27535,N_27733);
nor U27980 (N_27980,N_27570,N_27637);
or U27981 (N_27981,N_27517,N_27637);
xnor U27982 (N_27982,N_27552,N_27539);
nor U27983 (N_27983,N_27656,N_27558);
nor U27984 (N_27984,N_27644,N_27733);
nor U27985 (N_27985,N_27588,N_27526);
xnor U27986 (N_27986,N_27615,N_27692);
nor U27987 (N_27987,N_27601,N_27561);
and U27988 (N_27988,N_27608,N_27626);
xnor U27989 (N_27989,N_27536,N_27626);
and U27990 (N_27990,N_27622,N_27534);
or U27991 (N_27991,N_27720,N_27513);
nor U27992 (N_27992,N_27520,N_27539);
and U27993 (N_27993,N_27689,N_27512);
and U27994 (N_27994,N_27677,N_27617);
and U27995 (N_27995,N_27625,N_27581);
nor U27996 (N_27996,N_27727,N_27585);
or U27997 (N_27997,N_27548,N_27607);
or U27998 (N_27998,N_27643,N_27722);
or U27999 (N_27999,N_27609,N_27616);
nand U28000 (N_28000,N_27979,N_27978);
or U28001 (N_28001,N_27844,N_27933);
xnor U28002 (N_28002,N_27943,N_27928);
xnor U28003 (N_28003,N_27785,N_27894);
nand U28004 (N_28004,N_27937,N_27836);
and U28005 (N_28005,N_27919,N_27828);
or U28006 (N_28006,N_27835,N_27807);
and U28007 (N_28007,N_27968,N_27855);
nor U28008 (N_28008,N_27955,N_27797);
or U28009 (N_28009,N_27804,N_27848);
xnor U28010 (N_28010,N_27900,N_27983);
nor U28011 (N_28011,N_27877,N_27774);
nand U28012 (N_28012,N_27930,N_27852);
nor U28013 (N_28013,N_27934,N_27795);
nor U28014 (N_28014,N_27791,N_27811);
or U28015 (N_28015,N_27873,N_27778);
and U28016 (N_28016,N_27911,N_27851);
xor U28017 (N_28017,N_27879,N_27862);
xor U28018 (N_28018,N_27856,N_27945);
nor U28019 (N_28019,N_27845,N_27962);
xor U28020 (N_28020,N_27751,N_27808);
and U28021 (N_28021,N_27763,N_27980);
xor U28022 (N_28022,N_27782,N_27938);
nand U28023 (N_28023,N_27770,N_27947);
nor U28024 (N_28024,N_27802,N_27949);
xor U28025 (N_28025,N_27820,N_27936);
or U28026 (N_28026,N_27875,N_27769);
or U28027 (N_28027,N_27914,N_27970);
xnor U28028 (N_28028,N_27896,N_27765);
and U28029 (N_28029,N_27815,N_27893);
xnor U28030 (N_28030,N_27889,N_27939);
or U28031 (N_28031,N_27923,N_27841);
and U28032 (N_28032,N_27837,N_27957);
or U28033 (N_28033,N_27982,N_27948);
and U28034 (N_28034,N_27903,N_27756);
nor U28035 (N_28035,N_27927,N_27798);
nand U28036 (N_28036,N_27908,N_27926);
xor U28037 (N_28037,N_27822,N_27762);
xor U28038 (N_28038,N_27959,N_27790);
xnor U28039 (N_28039,N_27783,N_27816);
xor U28040 (N_28040,N_27986,N_27975);
nor U28041 (N_28041,N_27898,N_27831);
nor U28042 (N_28042,N_27932,N_27915);
and U28043 (N_28043,N_27784,N_27918);
xor U28044 (N_28044,N_27787,N_27752);
and U28045 (N_28045,N_27990,N_27843);
or U28046 (N_28046,N_27840,N_27806);
and U28047 (N_28047,N_27964,N_27832);
xnor U28048 (N_28048,N_27897,N_27818);
or U28049 (N_28049,N_27772,N_27773);
and U28050 (N_28050,N_27868,N_27985);
nand U28051 (N_28051,N_27882,N_27767);
xnor U28052 (N_28052,N_27940,N_27917);
or U28053 (N_28053,N_27942,N_27850);
or U28054 (N_28054,N_27906,N_27809);
and U28055 (N_28055,N_27865,N_27971);
and U28056 (N_28056,N_27965,N_27866);
nand U28057 (N_28057,N_27776,N_27988);
or U28058 (N_28058,N_27824,N_27973);
nand U28059 (N_28059,N_27922,N_27853);
nand U28060 (N_28060,N_27909,N_27929);
xor U28061 (N_28061,N_27895,N_27876);
and U28062 (N_28062,N_27830,N_27952);
or U28063 (N_28063,N_27913,N_27833);
nand U28064 (N_28064,N_27759,N_27810);
xnor U28065 (N_28065,N_27825,N_27887);
nand U28066 (N_28066,N_27786,N_27958);
or U28067 (N_28067,N_27977,N_27801);
and U28068 (N_28068,N_27800,N_27966);
nand U28069 (N_28069,N_27757,N_27967);
and U28070 (N_28070,N_27997,N_27881);
nor U28071 (N_28071,N_27885,N_27951);
xor U28072 (N_28072,N_27781,N_27974);
or U28073 (N_28073,N_27849,N_27863);
and U28074 (N_28074,N_27771,N_27976);
nand U28075 (N_28075,N_27766,N_27874);
nand U28076 (N_28076,N_27750,N_27969);
or U28077 (N_28077,N_27880,N_27871);
and U28078 (N_28078,N_27907,N_27813);
and U28079 (N_28079,N_27861,N_27788);
nor U28080 (N_28080,N_27817,N_27864);
and U28081 (N_28081,N_27854,N_27796);
xor U28082 (N_28082,N_27847,N_27944);
nor U28083 (N_28083,N_27753,N_27870);
nand U28084 (N_28084,N_27912,N_27960);
or U28085 (N_28085,N_27891,N_27827);
nor U28086 (N_28086,N_27996,N_27755);
and U28087 (N_28087,N_27814,N_27991);
nor U28088 (N_28088,N_27920,N_27886);
or U28089 (N_28089,N_27892,N_27777);
xnor U28090 (N_28090,N_27910,N_27994);
nand U28091 (N_28091,N_27883,N_27799);
or U28092 (N_28092,N_27789,N_27987);
nand U28093 (N_28093,N_27992,N_27867);
and U28094 (N_28094,N_27823,N_27950);
xnor U28095 (N_28095,N_27834,N_27935);
and U28096 (N_28096,N_27916,N_27860);
nor U28097 (N_28097,N_27805,N_27754);
xnor U28098 (N_28098,N_27931,N_27995);
xnor U28099 (N_28099,N_27899,N_27956);
nor U28100 (N_28100,N_27998,N_27946);
or U28101 (N_28101,N_27921,N_27963);
xnor U28102 (N_28102,N_27925,N_27826);
xnor U28103 (N_28103,N_27981,N_27768);
xnor U28104 (N_28104,N_27839,N_27792);
xnor U28105 (N_28105,N_27794,N_27954);
xor U28106 (N_28106,N_27842,N_27905);
and U28107 (N_28107,N_27760,N_27872);
xnor U28108 (N_28108,N_27780,N_27884);
xnor U28109 (N_28109,N_27858,N_27793);
xor U28110 (N_28110,N_27924,N_27941);
nand U28111 (N_28111,N_27993,N_27764);
and U28112 (N_28112,N_27999,N_27857);
nand U28113 (N_28113,N_27838,N_27829);
nand U28114 (N_28114,N_27775,N_27859);
or U28115 (N_28115,N_27812,N_27888);
or U28116 (N_28116,N_27761,N_27972);
nand U28117 (N_28117,N_27984,N_27890);
and U28118 (N_28118,N_27989,N_27902);
xnor U28119 (N_28119,N_27869,N_27819);
or U28120 (N_28120,N_27846,N_27878);
xor U28121 (N_28121,N_27803,N_27821);
nand U28122 (N_28122,N_27961,N_27904);
and U28123 (N_28123,N_27779,N_27901);
xor U28124 (N_28124,N_27758,N_27953);
and U28125 (N_28125,N_27760,N_27909);
or U28126 (N_28126,N_27954,N_27911);
or U28127 (N_28127,N_27935,N_27956);
xor U28128 (N_28128,N_27933,N_27940);
xor U28129 (N_28129,N_27789,N_27899);
xor U28130 (N_28130,N_27816,N_27853);
xnor U28131 (N_28131,N_27912,N_27861);
xor U28132 (N_28132,N_27940,N_27969);
nand U28133 (N_28133,N_27837,N_27896);
nand U28134 (N_28134,N_27822,N_27880);
xnor U28135 (N_28135,N_27930,N_27996);
xor U28136 (N_28136,N_27933,N_27904);
or U28137 (N_28137,N_27781,N_27898);
and U28138 (N_28138,N_27973,N_27793);
or U28139 (N_28139,N_27867,N_27976);
or U28140 (N_28140,N_27900,N_27833);
xor U28141 (N_28141,N_27912,N_27940);
nand U28142 (N_28142,N_27910,N_27794);
xor U28143 (N_28143,N_27930,N_27949);
or U28144 (N_28144,N_27840,N_27969);
xnor U28145 (N_28145,N_27948,N_27816);
nor U28146 (N_28146,N_27861,N_27976);
and U28147 (N_28147,N_27912,N_27785);
and U28148 (N_28148,N_27926,N_27779);
xor U28149 (N_28149,N_27979,N_27783);
nand U28150 (N_28150,N_27884,N_27964);
or U28151 (N_28151,N_27960,N_27943);
and U28152 (N_28152,N_27900,N_27921);
xnor U28153 (N_28153,N_27753,N_27992);
or U28154 (N_28154,N_27794,N_27868);
and U28155 (N_28155,N_27796,N_27795);
and U28156 (N_28156,N_27815,N_27898);
nand U28157 (N_28157,N_27969,N_27867);
nor U28158 (N_28158,N_27921,N_27819);
xor U28159 (N_28159,N_27874,N_27862);
nand U28160 (N_28160,N_27875,N_27948);
nand U28161 (N_28161,N_27976,N_27768);
nor U28162 (N_28162,N_27865,N_27885);
and U28163 (N_28163,N_27801,N_27874);
nor U28164 (N_28164,N_27919,N_27765);
or U28165 (N_28165,N_27872,N_27994);
nand U28166 (N_28166,N_27864,N_27993);
nand U28167 (N_28167,N_27862,N_27997);
and U28168 (N_28168,N_27770,N_27761);
nor U28169 (N_28169,N_27792,N_27802);
nor U28170 (N_28170,N_27865,N_27853);
nor U28171 (N_28171,N_27778,N_27869);
or U28172 (N_28172,N_27811,N_27849);
nor U28173 (N_28173,N_27866,N_27873);
nand U28174 (N_28174,N_27972,N_27774);
nor U28175 (N_28175,N_27939,N_27885);
and U28176 (N_28176,N_27888,N_27958);
or U28177 (N_28177,N_27963,N_27929);
nand U28178 (N_28178,N_27895,N_27842);
nor U28179 (N_28179,N_27816,N_27767);
and U28180 (N_28180,N_27794,N_27859);
xnor U28181 (N_28181,N_27988,N_27961);
or U28182 (N_28182,N_27757,N_27756);
xor U28183 (N_28183,N_27854,N_27969);
nand U28184 (N_28184,N_27989,N_27760);
nor U28185 (N_28185,N_27789,N_27914);
nor U28186 (N_28186,N_27832,N_27987);
and U28187 (N_28187,N_27758,N_27773);
nor U28188 (N_28188,N_27864,N_27808);
and U28189 (N_28189,N_27876,N_27832);
or U28190 (N_28190,N_27760,N_27997);
nor U28191 (N_28191,N_27961,N_27759);
nor U28192 (N_28192,N_27822,N_27804);
xor U28193 (N_28193,N_27929,N_27785);
and U28194 (N_28194,N_27971,N_27996);
or U28195 (N_28195,N_27973,N_27873);
xor U28196 (N_28196,N_27854,N_27840);
and U28197 (N_28197,N_27908,N_27967);
nand U28198 (N_28198,N_27757,N_27946);
xnor U28199 (N_28199,N_27864,N_27858);
and U28200 (N_28200,N_27880,N_27891);
nor U28201 (N_28201,N_27759,N_27879);
and U28202 (N_28202,N_27818,N_27845);
and U28203 (N_28203,N_27848,N_27790);
nand U28204 (N_28204,N_27927,N_27994);
nor U28205 (N_28205,N_27936,N_27870);
nand U28206 (N_28206,N_27930,N_27889);
and U28207 (N_28207,N_27818,N_27966);
nand U28208 (N_28208,N_27992,N_27905);
nand U28209 (N_28209,N_27958,N_27761);
or U28210 (N_28210,N_27776,N_27886);
nor U28211 (N_28211,N_27976,N_27850);
and U28212 (N_28212,N_27892,N_27906);
nand U28213 (N_28213,N_27947,N_27964);
and U28214 (N_28214,N_27777,N_27991);
and U28215 (N_28215,N_27812,N_27869);
and U28216 (N_28216,N_27880,N_27878);
and U28217 (N_28217,N_27820,N_27770);
and U28218 (N_28218,N_27861,N_27955);
or U28219 (N_28219,N_27962,N_27937);
nand U28220 (N_28220,N_27815,N_27878);
xnor U28221 (N_28221,N_27865,N_27946);
xnor U28222 (N_28222,N_27775,N_27974);
or U28223 (N_28223,N_27814,N_27817);
nand U28224 (N_28224,N_27863,N_27829);
nand U28225 (N_28225,N_27893,N_27938);
and U28226 (N_28226,N_27830,N_27822);
nand U28227 (N_28227,N_27773,N_27940);
nor U28228 (N_28228,N_27864,N_27981);
xnor U28229 (N_28229,N_27984,N_27877);
and U28230 (N_28230,N_27841,N_27947);
nand U28231 (N_28231,N_27916,N_27791);
nor U28232 (N_28232,N_27964,N_27890);
nor U28233 (N_28233,N_27964,N_27974);
nor U28234 (N_28234,N_27960,N_27897);
nor U28235 (N_28235,N_27826,N_27960);
xnor U28236 (N_28236,N_27833,N_27788);
and U28237 (N_28237,N_27910,N_27820);
xnor U28238 (N_28238,N_27932,N_27980);
or U28239 (N_28239,N_27928,N_27961);
xor U28240 (N_28240,N_27928,N_27892);
xor U28241 (N_28241,N_27759,N_27945);
nor U28242 (N_28242,N_27954,N_27882);
and U28243 (N_28243,N_27894,N_27979);
xnor U28244 (N_28244,N_27794,N_27960);
or U28245 (N_28245,N_27776,N_27752);
or U28246 (N_28246,N_27979,N_27781);
nand U28247 (N_28247,N_27831,N_27756);
xor U28248 (N_28248,N_27917,N_27948);
xor U28249 (N_28249,N_27960,N_27765);
xor U28250 (N_28250,N_28189,N_28158);
xnor U28251 (N_28251,N_28167,N_28246);
xnor U28252 (N_28252,N_28171,N_28088);
nand U28253 (N_28253,N_28185,N_28075);
nand U28254 (N_28254,N_28245,N_28012);
nor U28255 (N_28255,N_28102,N_28145);
and U28256 (N_28256,N_28148,N_28034);
xnor U28257 (N_28257,N_28107,N_28108);
nor U28258 (N_28258,N_28015,N_28045);
and U28259 (N_28259,N_28050,N_28043);
xor U28260 (N_28260,N_28217,N_28164);
nand U28261 (N_28261,N_28198,N_28220);
or U28262 (N_28262,N_28090,N_28060);
xor U28263 (N_28263,N_28177,N_28097);
and U28264 (N_28264,N_28183,N_28115);
or U28265 (N_28265,N_28131,N_28091);
and U28266 (N_28266,N_28149,N_28044);
nor U28267 (N_28267,N_28071,N_28182);
nor U28268 (N_28268,N_28008,N_28187);
nor U28269 (N_28269,N_28074,N_28132);
xor U28270 (N_28270,N_28014,N_28138);
xnor U28271 (N_28271,N_28048,N_28006);
or U28272 (N_28272,N_28221,N_28018);
or U28273 (N_28273,N_28168,N_28092);
nand U28274 (N_28274,N_28111,N_28248);
xnor U28275 (N_28275,N_28101,N_28104);
nor U28276 (N_28276,N_28000,N_28144);
nor U28277 (N_28277,N_28042,N_28002);
xnor U28278 (N_28278,N_28021,N_28166);
or U28279 (N_28279,N_28224,N_28037);
nand U28280 (N_28280,N_28064,N_28094);
xor U28281 (N_28281,N_28159,N_28228);
and U28282 (N_28282,N_28204,N_28249);
or U28283 (N_28283,N_28047,N_28157);
or U28284 (N_28284,N_28233,N_28103);
and U28285 (N_28285,N_28197,N_28054);
nand U28286 (N_28286,N_28143,N_28001);
and U28287 (N_28287,N_28030,N_28160);
nor U28288 (N_28288,N_28087,N_28243);
and U28289 (N_28289,N_28058,N_28128);
nor U28290 (N_28290,N_28239,N_28055);
nand U28291 (N_28291,N_28084,N_28114);
or U28292 (N_28292,N_28009,N_28162);
nor U28293 (N_28293,N_28086,N_28033);
nand U28294 (N_28294,N_28242,N_28146);
nor U28295 (N_28295,N_28121,N_28209);
or U28296 (N_28296,N_28240,N_28192);
xor U28297 (N_28297,N_28175,N_28024);
and U28298 (N_28298,N_28215,N_28218);
nand U28299 (N_28299,N_28142,N_28029);
nand U28300 (N_28300,N_28027,N_28200);
nand U28301 (N_28301,N_28163,N_28036);
nor U28302 (N_28302,N_28190,N_28078);
nand U28303 (N_28303,N_28057,N_28193);
nor U28304 (N_28304,N_28203,N_28093);
or U28305 (N_28305,N_28105,N_28098);
xor U28306 (N_28306,N_28123,N_28174);
and U28307 (N_28307,N_28089,N_28120);
nor U28308 (N_28308,N_28134,N_28213);
xnor U28309 (N_28309,N_28161,N_28095);
nand U28310 (N_28310,N_28053,N_28178);
or U28311 (N_28311,N_28010,N_28194);
nor U28312 (N_28312,N_28096,N_28234);
xnor U28313 (N_28313,N_28100,N_28022);
nand U28314 (N_28314,N_28026,N_28133);
nand U28315 (N_28315,N_28226,N_28152);
and U28316 (N_28316,N_28230,N_28184);
or U28317 (N_28317,N_28020,N_28049);
or U28318 (N_28318,N_28082,N_28025);
or U28319 (N_28319,N_28031,N_28135);
and U28320 (N_28320,N_28176,N_28028);
nand U28321 (N_28321,N_28188,N_28068);
or U28322 (N_28322,N_28196,N_28117);
nor U28323 (N_28323,N_28165,N_28023);
xor U28324 (N_28324,N_28223,N_28040);
xor U28325 (N_28325,N_28214,N_28169);
nand U28326 (N_28326,N_28059,N_28173);
and U28327 (N_28327,N_28195,N_28052);
or U28328 (N_28328,N_28005,N_28099);
nor U28329 (N_28329,N_28129,N_28211);
or U28330 (N_28330,N_28072,N_28191);
xor U28331 (N_28331,N_28127,N_28083);
xor U28332 (N_28332,N_28017,N_28153);
or U28333 (N_28333,N_28210,N_28238);
xnor U28334 (N_28334,N_28062,N_28051);
and U28335 (N_28335,N_28170,N_28179);
nand U28336 (N_28336,N_28130,N_28003);
and U28337 (N_28337,N_28080,N_28122);
nand U28338 (N_28338,N_28113,N_28229);
xor U28339 (N_28339,N_28155,N_28208);
or U28340 (N_28340,N_28181,N_28201);
nor U28341 (N_28341,N_28067,N_28186);
nand U28342 (N_28342,N_28079,N_28244);
nor U28343 (N_28343,N_28066,N_28219);
xor U28344 (N_28344,N_28225,N_28140);
xnor U28345 (N_28345,N_28180,N_28013);
and U28346 (N_28346,N_28202,N_28235);
xnor U28347 (N_28347,N_28126,N_28124);
and U28348 (N_28348,N_28041,N_28231);
or U28349 (N_28349,N_28065,N_28137);
xor U28350 (N_28350,N_28061,N_28038);
xor U28351 (N_28351,N_28116,N_28112);
nor U28352 (N_28352,N_28119,N_28136);
nor U28353 (N_28353,N_28085,N_28222);
xnor U28354 (N_28354,N_28011,N_28063);
nand U28355 (N_28355,N_28156,N_28172);
nand U28356 (N_28356,N_28077,N_28207);
nor U28357 (N_28357,N_28118,N_28150);
or U28358 (N_28358,N_28035,N_28069);
xnor U28359 (N_28359,N_28073,N_28199);
nand U28360 (N_28360,N_28039,N_28004);
or U28361 (N_28361,N_28106,N_28032);
xnor U28362 (N_28362,N_28007,N_28016);
nor U28363 (N_28363,N_28236,N_28019);
nor U28364 (N_28364,N_28046,N_28076);
nor U28365 (N_28365,N_28205,N_28227);
and U28366 (N_28366,N_28241,N_28237);
or U28367 (N_28367,N_28147,N_28154);
nor U28368 (N_28368,N_28216,N_28109);
xor U28369 (N_28369,N_28151,N_28110);
or U28370 (N_28370,N_28141,N_28125);
nand U28371 (N_28371,N_28070,N_28056);
nor U28372 (N_28372,N_28081,N_28247);
xor U28373 (N_28373,N_28139,N_28232);
and U28374 (N_28374,N_28206,N_28212);
xnor U28375 (N_28375,N_28087,N_28076);
xnor U28376 (N_28376,N_28055,N_28141);
nand U28377 (N_28377,N_28081,N_28015);
nand U28378 (N_28378,N_28021,N_28208);
or U28379 (N_28379,N_28181,N_28073);
and U28380 (N_28380,N_28071,N_28243);
and U28381 (N_28381,N_28142,N_28075);
nor U28382 (N_28382,N_28086,N_28002);
or U28383 (N_28383,N_28157,N_28132);
nand U28384 (N_28384,N_28024,N_28205);
xnor U28385 (N_28385,N_28086,N_28056);
and U28386 (N_28386,N_28027,N_28107);
and U28387 (N_28387,N_28024,N_28098);
xnor U28388 (N_28388,N_28033,N_28249);
xor U28389 (N_28389,N_28073,N_28005);
or U28390 (N_28390,N_28032,N_28060);
or U28391 (N_28391,N_28236,N_28235);
nand U28392 (N_28392,N_28018,N_28075);
nand U28393 (N_28393,N_28059,N_28238);
and U28394 (N_28394,N_28146,N_28238);
and U28395 (N_28395,N_28042,N_28119);
and U28396 (N_28396,N_28103,N_28098);
or U28397 (N_28397,N_28060,N_28008);
xnor U28398 (N_28398,N_28103,N_28095);
xnor U28399 (N_28399,N_28110,N_28006);
or U28400 (N_28400,N_28058,N_28238);
nor U28401 (N_28401,N_28159,N_28065);
and U28402 (N_28402,N_28161,N_28040);
and U28403 (N_28403,N_28113,N_28243);
nand U28404 (N_28404,N_28205,N_28101);
or U28405 (N_28405,N_28014,N_28000);
xor U28406 (N_28406,N_28188,N_28109);
nand U28407 (N_28407,N_28244,N_28069);
nor U28408 (N_28408,N_28150,N_28160);
or U28409 (N_28409,N_28093,N_28138);
or U28410 (N_28410,N_28202,N_28227);
and U28411 (N_28411,N_28194,N_28038);
or U28412 (N_28412,N_28120,N_28144);
xnor U28413 (N_28413,N_28050,N_28249);
nand U28414 (N_28414,N_28019,N_28222);
nor U28415 (N_28415,N_28174,N_28234);
and U28416 (N_28416,N_28200,N_28030);
and U28417 (N_28417,N_28112,N_28203);
xnor U28418 (N_28418,N_28024,N_28167);
or U28419 (N_28419,N_28006,N_28143);
or U28420 (N_28420,N_28076,N_28206);
xor U28421 (N_28421,N_28160,N_28209);
nor U28422 (N_28422,N_28100,N_28150);
or U28423 (N_28423,N_28019,N_28113);
nor U28424 (N_28424,N_28012,N_28150);
and U28425 (N_28425,N_28094,N_28012);
and U28426 (N_28426,N_28090,N_28219);
nand U28427 (N_28427,N_28162,N_28098);
and U28428 (N_28428,N_28242,N_28007);
and U28429 (N_28429,N_28089,N_28058);
and U28430 (N_28430,N_28127,N_28244);
or U28431 (N_28431,N_28059,N_28103);
xor U28432 (N_28432,N_28131,N_28129);
xor U28433 (N_28433,N_28227,N_28182);
or U28434 (N_28434,N_28233,N_28041);
xnor U28435 (N_28435,N_28116,N_28025);
and U28436 (N_28436,N_28249,N_28016);
nor U28437 (N_28437,N_28096,N_28187);
xor U28438 (N_28438,N_28061,N_28063);
nor U28439 (N_28439,N_28047,N_28002);
or U28440 (N_28440,N_28099,N_28041);
nor U28441 (N_28441,N_28013,N_28003);
xnor U28442 (N_28442,N_28115,N_28189);
or U28443 (N_28443,N_28046,N_28125);
and U28444 (N_28444,N_28109,N_28241);
or U28445 (N_28445,N_28228,N_28037);
or U28446 (N_28446,N_28221,N_28201);
nor U28447 (N_28447,N_28048,N_28092);
or U28448 (N_28448,N_28027,N_28197);
xor U28449 (N_28449,N_28142,N_28184);
nand U28450 (N_28450,N_28026,N_28055);
nand U28451 (N_28451,N_28135,N_28148);
nand U28452 (N_28452,N_28091,N_28231);
xor U28453 (N_28453,N_28048,N_28152);
nor U28454 (N_28454,N_28017,N_28026);
xnor U28455 (N_28455,N_28143,N_28049);
nor U28456 (N_28456,N_28021,N_28168);
xnor U28457 (N_28457,N_28249,N_28006);
nor U28458 (N_28458,N_28189,N_28135);
xor U28459 (N_28459,N_28028,N_28224);
nor U28460 (N_28460,N_28221,N_28073);
xnor U28461 (N_28461,N_28227,N_28060);
or U28462 (N_28462,N_28101,N_28171);
or U28463 (N_28463,N_28027,N_28239);
nand U28464 (N_28464,N_28232,N_28153);
xor U28465 (N_28465,N_28173,N_28213);
or U28466 (N_28466,N_28128,N_28202);
nand U28467 (N_28467,N_28013,N_28095);
and U28468 (N_28468,N_28015,N_28054);
nor U28469 (N_28469,N_28013,N_28049);
nand U28470 (N_28470,N_28225,N_28121);
or U28471 (N_28471,N_28058,N_28135);
nand U28472 (N_28472,N_28172,N_28162);
nor U28473 (N_28473,N_28122,N_28019);
or U28474 (N_28474,N_28113,N_28178);
nor U28475 (N_28475,N_28212,N_28077);
or U28476 (N_28476,N_28133,N_28246);
nand U28477 (N_28477,N_28097,N_28044);
nand U28478 (N_28478,N_28145,N_28249);
nor U28479 (N_28479,N_28132,N_28165);
and U28480 (N_28480,N_28071,N_28179);
nor U28481 (N_28481,N_28144,N_28165);
nor U28482 (N_28482,N_28245,N_28212);
nor U28483 (N_28483,N_28059,N_28037);
and U28484 (N_28484,N_28214,N_28032);
and U28485 (N_28485,N_28117,N_28060);
nor U28486 (N_28486,N_28179,N_28009);
xor U28487 (N_28487,N_28041,N_28020);
or U28488 (N_28488,N_28053,N_28074);
or U28489 (N_28489,N_28036,N_28153);
and U28490 (N_28490,N_28064,N_28209);
or U28491 (N_28491,N_28122,N_28211);
or U28492 (N_28492,N_28143,N_28229);
or U28493 (N_28493,N_28174,N_28044);
nor U28494 (N_28494,N_28200,N_28214);
and U28495 (N_28495,N_28043,N_28194);
xor U28496 (N_28496,N_28169,N_28184);
and U28497 (N_28497,N_28158,N_28205);
xnor U28498 (N_28498,N_28057,N_28095);
or U28499 (N_28499,N_28034,N_28127);
nor U28500 (N_28500,N_28276,N_28357);
nor U28501 (N_28501,N_28467,N_28438);
xnor U28502 (N_28502,N_28418,N_28407);
and U28503 (N_28503,N_28273,N_28347);
nor U28504 (N_28504,N_28495,N_28258);
nand U28505 (N_28505,N_28296,N_28382);
nand U28506 (N_28506,N_28486,N_28399);
or U28507 (N_28507,N_28391,N_28309);
or U28508 (N_28508,N_28275,N_28494);
nor U28509 (N_28509,N_28255,N_28343);
nand U28510 (N_28510,N_28412,N_28465);
nand U28511 (N_28511,N_28388,N_28351);
nand U28512 (N_28512,N_28381,N_28436);
or U28513 (N_28513,N_28476,N_28342);
nand U28514 (N_28514,N_28284,N_28352);
or U28515 (N_28515,N_28410,N_28350);
and U28516 (N_28516,N_28338,N_28453);
or U28517 (N_28517,N_28462,N_28251);
nor U28518 (N_28518,N_28425,N_28355);
and U28519 (N_28519,N_28283,N_28400);
xnor U28520 (N_28520,N_28334,N_28300);
and U28521 (N_28521,N_28333,N_28403);
xor U28522 (N_28522,N_28493,N_28393);
nor U28523 (N_28523,N_28370,N_28487);
xnor U28524 (N_28524,N_28405,N_28499);
and U28525 (N_28525,N_28329,N_28398);
xnor U28526 (N_28526,N_28371,N_28423);
or U28527 (N_28527,N_28291,N_28435);
and U28528 (N_28528,N_28426,N_28409);
or U28529 (N_28529,N_28253,N_28298);
nand U28530 (N_28530,N_28460,N_28481);
nand U28531 (N_28531,N_28377,N_28361);
nand U28532 (N_28532,N_28379,N_28431);
or U28533 (N_28533,N_28348,N_28312);
or U28534 (N_28534,N_28261,N_28353);
and U28535 (N_28535,N_28301,N_28252);
nor U28536 (N_28536,N_28433,N_28455);
nor U28537 (N_28537,N_28411,N_28443);
nand U28538 (N_28538,N_28360,N_28359);
and U28539 (N_28539,N_28277,N_28290);
xnor U28540 (N_28540,N_28386,N_28406);
xnor U28541 (N_28541,N_28306,N_28268);
or U28542 (N_28542,N_28363,N_28389);
and U28543 (N_28543,N_28264,N_28445);
and U28544 (N_28544,N_28419,N_28485);
or U28545 (N_28545,N_28437,N_28307);
and U28546 (N_28546,N_28451,N_28447);
or U28547 (N_28547,N_28375,N_28368);
or U28548 (N_28548,N_28341,N_28414);
nand U28549 (N_28549,N_28280,N_28470);
nor U28550 (N_28550,N_28285,N_28478);
and U28551 (N_28551,N_28332,N_28325);
or U28552 (N_28552,N_28452,N_28317);
nand U28553 (N_28553,N_28305,N_28318);
nor U28554 (N_28554,N_28430,N_28254);
nor U28555 (N_28555,N_28297,N_28269);
and U28556 (N_28556,N_28482,N_28302);
nand U28557 (N_28557,N_28427,N_28415);
nor U28558 (N_28558,N_28311,N_28266);
nand U28559 (N_28559,N_28295,N_28314);
or U28560 (N_28560,N_28271,N_28424);
and U28561 (N_28561,N_28369,N_28364);
and U28562 (N_28562,N_28315,N_28344);
nor U28563 (N_28563,N_28491,N_28428);
nor U28564 (N_28564,N_28278,N_28473);
nand U28565 (N_28565,N_28260,N_28265);
and U28566 (N_28566,N_28463,N_28413);
nand U28567 (N_28567,N_28469,N_28257);
and U28568 (N_28568,N_28444,N_28440);
nand U28569 (N_28569,N_28328,N_28489);
nor U28570 (N_28570,N_28456,N_28339);
nand U28571 (N_28571,N_28335,N_28294);
and U28572 (N_28572,N_28378,N_28281);
xor U28573 (N_28573,N_28446,N_28262);
xor U28574 (N_28574,N_28390,N_28349);
nand U28575 (N_28575,N_28448,N_28387);
or U28576 (N_28576,N_28282,N_28279);
or U28577 (N_28577,N_28422,N_28374);
xor U28578 (N_28578,N_28497,N_28383);
nand U28579 (N_28579,N_28397,N_28472);
or U28580 (N_28580,N_28292,N_28492);
and U28581 (N_28581,N_28466,N_28490);
and U28582 (N_28582,N_28356,N_28496);
nor U28583 (N_28583,N_28458,N_28330);
and U28584 (N_28584,N_28346,N_28385);
and U28585 (N_28585,N_28464,N_28256);
or U28586 (N_28586,N_28484,N_28286);
nor U28587 (N_28587,N_28471,N_28474);
xor U28588 (N_28588,N_28392,N_28336);
nor U28589 (N_28589,N_28366,N_28322);
or U28590 (N_28590,N_28404,N_28439);
and U28591 (N_28591,N_28373,N_28417);
and U28592 (N_28592,N_28340,N_28308);
or U28593 (N_28593,N_28432,N_28316);
nor U28594 (N_28594,N_28416,N_28274);
nor U28595 (N_28595,N_28358,N_28420);
and U28596 (N_28596,N_28310,N_28326);
nor U28597 (N_28597,N_28401,N_28498);
or U28598 (N_28598,N_28408,N_28289);
nor U28599 (N_28599,N_28331,N_28394);
xnor U28600 (N_28600,N_28396,N_28362);
nor U28601 (N_28601,N_28488,N_28479);
or U28602 (N_28602,N_28457,N_28337);
xnor U28603 (N_28603,N_28468,N_28429);
and U28604 (N_28604,N_28459,N_28477);
xnor U28605 (N_28605,N_28288,N_28259);
xor U28606 (N_28606,N_28345,N_28313);
nor U28607 (N_28607,N_28441,N_28321);
xnor U28608 (N_28608,N_28304,N_28327);
and U28609 (N_28609,N_28287,N_28250);
or U28610 (N_28610,N_28454,N_28323);
or U28611 (N_28611,N_28365,N_28320);
or U28612 (N_28612,N_28376,N_28319);
or U28613 (N_28613,N_28449,N_28263);
or U28614 (N_28614,N_28402,N_28372);
nand U28615 (N_28615,N_28324,N_28434);
nand U28616 (N_28616,N_28272,N_28303);
nand U28617 (N_28617,N_28267,N_28461);
nor U28618 (N_28618,N_28480,N_28354);
and U28619 (N_28619,N_28442,N_28367);
xnor U28620 (N_28620,N_28450,N_28395);
nor U28621 (N_28621,N_28384,N_28270);
nor U28622 (N_28622,N_28483,N_28380);
and U28623 (N_28623,N_28293,N_28299);
nand U28624 (N_28624,N_28475,N_28421);
or U28625 (N_28625,N_28342,N_28427);
nand U28626 (N_28626,N_28375,N_28355);
and U28627 (N_28627,N_28329,N_28348);
nor U28628 (N_28628,N_28278,N_28450);
xor U28629 (N_28629,N_28258,N_28425);
or U28630 (N_28630,N_28342,N_28329);
xnor U28631 (N_28631,N_28391,N_28374);
xor U28632 (N_28632,N_28475,N_28299);
nor U28633 (N_28633,N_28364,N_28370);
nor U28634 (N_28634,N_28482,N_28386);
nand U28635 (N_28635,N_28428,N_28448);
xnor U28636 (N_28636,N_28396,N_28346);
nor U28637 (N_28637,N_28338,N_28390);
or U28638 (N_28638,N_28416,N_28492);
or U28639 (N_28639,N_28254,N_28421);
or U28640 (N_28640,N_28496,N_28426);
and U28641 (N_28641,N_28396,N_28283);
and U28642 (N_28642,N_28271,N_28490);
xnor U28643 (N_28643,N_28437,N_28443);
xnor U28644 (N_28644,N_28361,N_28451);
or U28645 (N_28645,N_28284,N_28429);
nor U28646 (N_28646,N_28442,N_28292);
and U28647 (N_28647,N_28453,N_28251);
nor U28648 (N_28648,N_28463,N_28267);
xor U28649 (N_28649,N_28449,N_28269);
nor U28650 (N_28650,N_28400,N_28268);
nand U28651 (N_28651,N_28422,N_28315);
and U28652 (N_28652,N_28385,N_28347);
nor U28653 (N_28653,N_28320,N_28382);
and U28654 (N_28654,N_28292,N_28467);
nor U28655 (N_28655,N_28289,N_28477);
xor U28656 (N_28656,N_28288,N_28404);
or U28657 (N_28657,N_28330,N_28457);
and U28658 (N_28658,N_28446,N_28407);
xnor U28659 (N_28659,N_28414,N_28275);
and U28660 (N_28660,N_28291,N_28344);
and U28661 (N_28661,N_28462,N_28490);
and U28662 (N_28662,N_28294,N_28324);
nor U28663 (N_28663,N_28348,N_28322);
nor U28664 (N_28664,N_28352,N_28499);
xor U28665 (N_28665,N_28466,N_28260);
xor U28666 (N_28666,N_28490,N_28474);
nand U28667 (N_28667,N_28374,N_28365);
nand U28668 (N_28668,N_28292,N_28269);
or U28669 (N_28669,N_28318,N_28366);
nor U28670 (N_28670,N_28474,N_28328);
xor U28671 (N_28671,N_28360,N_28399);
nor U28672 (N_28672,N_28315,N_28376);
xnor U28673 (N_28673,N_28490,N_28382);
or U28674 (N_28674,N_28435,N_28422);
and U28675 (N_28675,N_28308,N_28331);
or U28676 (N_28676,N_28275,N_28477);
nand U28677 (N_28677,N_28348,N_28433);
and U28678 (N_28678,N_28384,N_28466);
nor U28679 (N_28679,N_28483,N_28309);
or U28680 (N_28680,N_28302,N_28372);
or U28681 (N_28681,N_28465,N_28439);
xnor U28682 (N_28682,N_28321,N_28259);
and U28683 (N_28683,N_28308,N_28443);
nand U28684 (N_28684,N_28399,N_28337);
or U28685 (N_28685,N_28256,N_28318);
nor U28686 (N_28686,N_28362,N_28307);
xor U28687 (N_28687,N_28336,N_28316);
and U28688 (N_28688,N_28450,N_28359);
nor U28689 (N_28689,N_28255,N_28416);
and U28690 (N_28690,N_28418,N_28470);
and U28691 (N_28691,N_28304,N_28379);
or U28692 (N_28692,N_28250,N_28252);
or U28693 (N_28693,N_28294,N_28326);
nor U28694 (N_28694,N_28301,N_28424);
nor U28695 (N_28695,N_28458,N_28445);
and U28696 (N_28696,N_28489,N_28317);
and U28697 (N_28697,N_28489,N_28462);
nand U28698 (N_28698,N_28373,N_28308);
nor U28699 (N_28699,N_28430,N_28299);
xnor U28700 (N_28700,N_28426,N_28349);
and U28701 (N_28701,N_28314,N_28428);
xnor U28702 (N_28702,N_28439,N_28344);
and U28703 (N_28703,N_28401,N_28499);
nor U28704 (N_28704,N_28334,N_28335);
nor U28705 (N_28705,N_28356,N_28486);
xnor U28706 (N_28706,N_28467,N_28278);
and U28707 (N_28707,N_28349,N_28419);
or U28708 (N_28708,N_28436,N_28465);
and U28709 (N_28709,N_28376,N_28493);
or U28710 (N_28710,N_28486,N_28305);
xor U28711 (N_28711,N_28306,N_28256);
xnor U28712 (N_28712,N_28283,N_28402);
xor U28713 (N_28713,N_28361,N_28285);
nor U28714 (N_28714,N_28384,N_28382);
nor U28715 (N_28715,N_28363,N_28334);
nand U28716 (N_28716,N_28389,N_28392);
xor U28717 (N_28717,N_28369,N_28482);
and U28718 (N_28718,N_28270,N_28265);
or U28719 (N_28719,N_28345,N_28343);
or U28720 (N_28720,N_28463,N_28403);
nand U28721 (N_28721,N_28349,N_28443);
xor U28722 (N_28722,N_28335,N_28338);
xnor U28723 (N_28723,N_28393,N_28454);
or U28724 (N_28724,N_28299,N_28372);
or U28725 (N_28725,N_28390,N_28371);
and U28726 (N_28726,N_28350,N_28484);
xor U28727 (N_28727,N_28282,N_28290);
nand U28728 (N_28728,N_28258,N_28276);
and U28729 (N_28729,N_28387,N_28436);
xnor U28730 (N_28730,N_28390,N_28495);
xnor U28731 (N_28731,N_28391,N_28318);
nand U28732 (N_28732,N_28359,N_28487);
or U28733 (N_28733,N_28290,N_28401);
or U28734 (N_28734,N_28358,N_28426);
nor U28735 (N_28735,N_28368,N_28261);
and U28736 (N_28736,N_28482,N_28334);
nand U28737 (N_28737,N_28403,N_28408);
and U28738 (N_28738,N_28264,N_28343);
nand U28739 (N_28739,N_28304,N_28438);
or U28740 (N_28740,N_28478,N_28351);
or U28741 (N_28741,N_28287,N_28316);
or U28742 (N_28742,N_28459,N_28320);
nand U28743 (N_28743,N_28273,N_28481);
nor U28744 (N_28744,N_28280,N_28490);
nor U28745 (N_28745,N_28495,N_28455);
nand U28746 (N_28746,N_28283,N_28379);
nor U28747 (N_28747,N_28338,N_28329);
xnor U28748 (N_28748,N_28395,N_28396);
nand U28749 (N_28749,N_28449,N_28319);
nand U28750 (N_28750,N_28580,N_28560);
and U28751 (N_28751,N_28582,N_28590);
nor U28752 (N_28752,N_28569,N_28734);
xnor U28753 (N_28753,N_28508,N_28566);
nand U28754 (N_28754,N_28662,N_28550);
or U28755 (N_28755,N_28528,N_28543);
xor U28756 (N_28756,N_28748,N_28611);
and U28757 (N_28757,N_28553,N_28724);
nor U28758 (N_28758,N_28591,N_28549);
and U28759 (N_28759,N_28594,N_28521);
or U28760 (N_28760,N_28608,N_28607);
nand U28761 (N_28761,N_28583,N_28720);
or U28762 (N_28762,N_28727,N_28527);
nand U28763 (N_28763,N_28686,N_28600);
or U28764 (N_28764,N_28663,N_28692);
and U28765 (N_28765,N_28532,N_28643);
xor U28766 (N_28766,N_28575,N_28661);
or U28767 (N_28767,N_28559,N_28697);
nor U28768 (N_28768,N_28693,N_28517);
xnor U28769 (N_28769,N_28584,N_28630);
nand U28770 (N_28770,N_28670,N_28647);
nand U28771 (N_28771,N_28555,N_28519);
and U28772 (N_28772,N_28636,N_28565);
nor U28773 (N_28773,N_28721,N_28633);
nor U28774 (N_28774,N_28731,N_28657);
nand U28775 (N_28775,N_28563,N_28551);
nor U28776 (N_28776,N_28533,N_28530);
and U28777 (N_28777,N_28523,N_28579);
and U28778 (N_28778,N_28604,N_28631);
or U28779 (N_28779,N_28511,N_28544);
nor U28780 (N_28780,N_28561,N_28616);
or U28781 (N_28781,N_28703,N_28699);
nor U28782 (N_28782,N_28539,N_28678);
xor U28783 (N_28783,N_28696,N_28688);
nand U28784 (N_28784,N_28638,N_28656);
nand U28785 (N_28785,N_28749,N_28504);
and U28786 (N_28786,N_28619,N_28624);
and U28787 (N_28787,N_28725,N_28618);
nand U28788 (N_28788,N_28667,N_28664);
nand U28789 (N_28789,N_28547,N_28743);
nand U28790 (N_28790,N_28674,N_28609);
and U28791 (N_28791,N_28716,N_28715);
and U28792 (N_28792,N_28573,N_28672);
xor U28793 (N_28793,N_28685,N_28660);
nor U28794 (N_28794,N_28687,N_28601);
nor U28795 (N_28795,N_28546,N_28714);
and U28796 (N_28796,N_28717,N_28700);
and U28797 (N_28797,N_28645,N_28535);
or U28798 (N_28798,N_28708,N_28556);
nor U28799 (N_28799,N_28634,N_28689);
or U28800 (N_28800,N_28669,N_28726);
and U28801 (N_28801,N_28621,N_28640);
nor U28802 (N_28802,N_28562,N_28723);
nor U28803 (N_28803,N_28512,N_28707);
nor U28804 (N_28804,N_28680,N_28529);
and U28805 (N_28805,N_28506,N_28733);
nor U28806 (N_28806,N_28642,N_28612);
and U28807 (N_28807,N_28735,N_28691);
and U28808 (N_28808,N_28541,N_28620);
nand U28809 (N_28809,N_28745,N_28627);
xnor U28810 (N_28810,N_28679,N_28596);
nor U28811 (N_28811,N_28558,N_28729);
and U28812 (N_28812,N_28581,N_28719);
nor U28813 (N_28813,N_28578,N_28500);
nor U28814 (N_28814,N_28671,N_28648);
and U28815 (N_28815,N_28510,N_28652);
and U28816 (N_28816,N_28589,N_28730);
and U28817 (N_28817,N_28653,N_28732);
xnor U28818 (N_28818,N_28538,N_28518);
and U28819 (N_28819,N_28628,N_28586);
and U28820 (N_28820,N_28675,N_28668);
or U28821 (N_28821,N_28552,N_28570);
nand U28822 (N_28822,N_28577,N_28606);
nand U28823 (N_28823,N_28592,N_28629);
and U28824 (N_28824,N_28659,N_28593);
nand U28825 (N_28825,N_28705,N_28650);
xor U28826 (N_28826,N_28644,N_28542);
and U28827 (N_28827,N_28637,N_28507);
nor U28828 (N_28828,N_28654,N_28614);
nor U28829 (N_28829,N_28515,N_28513);
and U28830 (N_28830,N_28603,N_28639);
nand U28831 (N_28831,N_28595,N_28572);
nand U28832 (N_28832,N_28567,N_28677);
nor U28833 (N_28833,N_28557,N_28649);
and U28834 (N_28834,N_28540,N_28509);
and U28835 (N_28835,N_28681,N_28706);
and U28836 (N_28836,N_28599,N_28564);
or U28837 (N_28837,N_28554,N_28673);
or U28838 (N_28838,N_28626,N_28746);
xor U28839 (N_28839,N_28682,N_28520);
nand U28840 (N_28840,N_28587,N_28514);
and U28841 (N_28841,N_28548,N_28739);
and U28842 (N_28842,N_28525,N_28622);
xor U28843 (N_28843,N_28701,N_28576);
nand U28844 (N_28844,N_28741,N_28702);
nand U28845 (N_28845,N_28588,N_28623);
nor U28846 (N_28846,N_28531,N_28625);
xnor U28847 (N_28847,N_28501,N_28505);
xnor U28848 (N_28848,N_28646,N_28712);
nand U28849 (N_28849,N_28574,N_28737);
nand U28850 (N_28850,N_28665,N_28524);
nand U28851 (N_28851,N_28522,N_28615);
and U28852 (N_28852,N_28571,N_28698);
xor U28853 (N_28853,N_28740,N_28728);
or U28854 (N_28854,N_28658,N_28502);
and U28855 (N_28855,N_28602,N_28536);
xor U28856 (N_28856,N_28676,N_28613);
and U28857 (N_28857,N_28516,N_28537);
nand U28858 (N_28858,N_28713,N_28655);
or U28859 (N_28859,N_28704,N_28610);
xor U28860 (N_28860,N_28683,N_28666);
xor U28861 (N_28861,N_28651,N_28503);
nor U28862 (N_28862,N_28710,N_28744);
nand U28863 (N_28863,N_28694,N_28585);
xnor U28864 (N_28864,N_28632,N_28568);
xnor U28865 (N_28865,N_28709,N_28742);
or U28866 (N_28866,N_28598,N_28605);
or U28867 (N_28867,N_28641,N_28718);
xor U28868 (N_28868,N_28597,N_28684);
nor U28869 (N_28869,N_28736,N_28738);
nand U28870 (N_28870,N_28635,N_28617);
nand U28871 (N_28871,N_28545,N_28711);
xor U28872 (N_28872,N_28690,N_28747);
nand U28873 (N_28873,N_28695,N_28534);
or U28874 (N_28874,N_28526,N_28722);
nand U28875 (N_28875,N_28580,N_28554);
or U28876 (N_28876,N_28668,N_28609);
xnor U28877 (N_28877,N_28724,N_28669);
or U28878 (N_28878,N_28665,N_28533);
xor U28879 (N_28879,N_28744,N_28538);
nor U28880 (N_28880,N_28533,N_28595);
nor U28881 (N_28881,N_28609,N_28642);
xor U28882 (N_28882,N_28510,N_28573);
or U28883 (N_28883,N_28541,N_28644);
xnor U28884 (N_28884,N_28681,N_28735);
xor U28885 (N_28885,N_28626,N_28553);
xor U28886 (N_28886,N_28671,N_28511);
nor U28887 (N_28887,N_28546,N_28662);
and U28888 (N_28888,N_28749,N_28664);
nor U28889 (N_28889,N_28628,N_28743);
nor U28890 (N_28890,N_28664,N_28550);
nor U28891 (N_28891,N_28627,N_28656);
or U28892 (N_28892,N_28574,N_28562);
xor U28893 (N_28893,N_28701,N_28516);
nand U28894 (N_28894,N_28727,N_28661);
or U28895 (N_28895,N_28640,N_28524);
nand U28896 (N_28896,N_28736,N_28519);
nor U28897 (N_28897,N_28647,N_28650);
nor U28898 (N_28898,N_28507,N_28537);
nor U28899 (N_28899,N_28713,N_28603);
xor U28900 (N_28900,N_28545,N_28733);
nor U28901 (N_28901,N_28659,N_28506);
nor U28902 (N_28902,N_28712,N_28633);
and U28903 (N_28903,N_28580,N_28677);
nand U28904 (N_28904,N_28684,N_28551);
xor U28905 (N_28905,N_28654,N_28651);
and U28906 (N_28906,N_28732,N_28645);
nand U28907 (N_28907,N_28625,N_28522);
and U28908 (N_28908,N_28538,N_28576);
nor U28909 (N_28909,N_28664,N_28703);
and U28910 (N_28910,N_28666,N_28606);
xor U28911 (N_28911,N_28578,N_28651);
and U28912 (N_28912,N_28733,N_28510);
nor U28913 (N_28913,N_28695,N_28621);
nand U28914 (N_28914,N_28637,N_28725);
xor U28915 (N_28915,N_28576,N_28615);
nand U28916 (N_28916,N_28696,N_28727);
nand U28917 (N_28917,N_28654,N_28685);
nand U28918 (N_28918,N_28581,N_28554);
and U28919 (N_28919,N_28633,N_28657);
nor U28920 (N_28920,N_28651,N_28658);
and U28921 (N_28921,N_28711,N_28675);
nand U28922 (N_28922,N_28515,N_28625);
nor U28923 (N_28923,N_28580,N_28690);
nand U28924 (N_28924,N_28664,N_28610);
and U28925 (N_28925,N_28662,N_28530);
and U28926 (N_28926,N_28715,N_28585);
nor U28927 (N_28927,N_28705,N_28712);
nor U28928 (N_28928,N_28658,N_28606);
and U28929 (N_28929,N_28513,N_28689);
nor U28930 (N_28930,N_28530,N_28607);
nor U28931 (N_28931,N_28644,N_28576);
and U28932 (N_28932,N_28552,N_28662);
nand U28933 (N_28933,N_28540,N_28649);
nand U28934 (N_28934,N_28590,N_28622);
nand U28935 (N_28935,N_28605,N_28723);
nand U28936 (N_28936,N_28556,N_28514);
and U28937 (N_28937,N_28715,N_28534);
nand U28938 (N_28938,N_28576,N_28524);
nand U28939 (N_28939,N_28735,N_28632);
and U28940 (N_28940,N_28663,N_28633);
nor U28941 (N_28941,N_28531,N_28608);
or U28942 (N_28942,N_28619,N_28589);
nor U28943 (N_28943,N_28643,N_28615);
xnor U28944 (N_28944,N_28552,N_28625);
nor U28945 (N_28945,N_28606,N_28583);
nand U28946 (N_28946,N_28704,N_28502);
xnor U28947 (N_28947,N_28559,N_28731);
xnor U28948 (N_28948,N_28678,N_28747);
xnor U28949 (N_28949,N_28636,N_28574);
nor U28950 (N_28950,N_28662,N_28589);
xnor U28951 (N_28951,N_28561,N_28680);
nand U28952 (N_28952,N_28568,N_28583);
xor U28953 (N_28953,N_28566,N_28590);
or U28954 (N_28954,N_28729,N_28646);
nor U28955 (N_28955,N_28542,N_28585);
or U28956 (N_28956,N_28602,N_28678);
or U28957 (N_28957,N_28578,N_28605);
xor U28958 (N_28958,N_28516,N_28599);
nor U28959 (N_28959,N_28740,N_28580);
nor U28960 (N_28960,N_28555,N_28576);
and U28961 (N_28961,N_28528,N_28614);
nand U28962 (N_28962,N_28533,N_28735);
or U28963 (N_28963,N_28715,N_28502);
nand U28964 (N_28964,N_28655,N_28521);
and U28965 (N_28965,N_28546,N_28744);
or U28966 (N_28966,N_28647,N_28522);
or U28967 (N_28967,N_28673,N_28588);
nor U28968 (N_28968,N_28662,N_28725);
nand U28969 (N_28969,N_28538,N_28611);
and U28970 (N_28970,N_28684,N_28733);
nand U28971 (N_28971,N_28633,N_28646);
xor U28972 (N_28972,N_28689,N_28690);
nor U28973 (N_28973,N_28689,N_28608);
nand U28974 (N_28974,N_28573,N_28592);
nor U28975 (N_28975,N_28673,N_28735);
nand U28976 (N_28976,N_28565,N_28687);
or U28977 (N_28977,N_28512,N_28621);
xnor U28978 (N_28978,N_28613,N_28662);
xor U28979 (N_28979,N_28660,N_28538);
xor U28980 (N_28980,N_28740,N_28679);
xor U28981 (N_28981,N_28589,N_28586);
xnor U28982 (N_28982,N_28656,N_28647);
xnor U28983 (N_28983,N_28689,N_28565);
and U28984 (N_28984,N_28501,N_28506);
nand U28985 (N_28985,N_28641,N_28553);
xor U28986 (N_28986,N_28526,N_28749);
and U28987 (N_28987,N_28560,N_28645);
nor U28988 (N_28988,N_28707,N_28748);
xnor U28989 (N_28989,N_28568,N_28738);
or U28990 (N_28990,N_28594,N_28502);
nand U28991 (N_28991,N_28621,N_28562);
nor U28992 (N_28992,N_28586,N_28519);
nand U28993 (N_28993,N_28707,N_28640);
xor U28994 (N_28994,N_28566,N_28559);
nor U28995 (N_28995,N_28727,N_28712);
and U28996 (N_28996,N_28744,N_28571);
and U28997 (N_28997,N_28500,N_28744);
or U28998 (N_28998,N_28704,N_28705);
and U28999 (N_28999,N_28643,N_28698);
xnor U29000 (N_29000,N_28801,N_28988);
xnor U29001 (N_29001,N_28980,N_28794);
xnor U29002 (N_29002,N_28879,N_28918);
and U29003 (N_29003,N_28992,N_28840);
nor U29004 (N_29004,N_28983,N_28771);
or U29005 (N_29005,N_28796,N_28960);
xnor U29006 (N_29006,N_28826,N_28819);
and U29007 (N_29007,N_28889,N_28795);
or U29008 (N_29008,N_28906,N_28791);
and U29009 (N_29009,N_28890,N_28777);
xnor U29010 (N_29010,N_28790,N_28940);
xor U29011 (N_29011,N_28915,N_28903);
nand U29012 (N_29012,N_28836,N_28877);
xor U29013 (N_29013,N_28870,N_28816);
nand U29014 (N_29014,N_28834,N_28900);
nor U29015 (N_29015,N_28961,N_28893);
and U29016 (N_29016,N_28865,N_28752);
or U29017 (N_29017,N_28912,N_28872);
nand U29018 (N_29018,N_28813,N_28979);
nor U29019 (N_29019,N_28999,N_28804);
and U29020 (N_29020,N_28841,N_28892);
xor U29021 (N_29021,N_28937,N_28994);
or U29022 (N_29022,N_28966,N_28754);
nor U29023 (N_29023,N_28965,N_28799);
xnor U29024 (N_29024,N_28783,N_28962);
nor U29025 (N_29025,N_28786,N_28942);
nand U29026 (N_29026,N_28830,N_28956);
and U29027 (N_29027,N_28871,N_28843);
and U29028 (N_29028,N_28936,N_28914);
and U29029 (N_29029,N_28846,N_28907);
or U29030 (N_29030,N_28986,N_28957);
or U29031 (N_29031,N_28993,N_28935);
nor U29032 (N_29032,N_28954,N_28904);
nand U29033 (N_29033,N_28932,N_28793);
xor U29034 (N_29034,N_28823,N_28897);
and U29035 (N_29035,N_28943,N_28989);
or U29036 (N_29036,N_28873,N_28821);
and U29037 (N_29037,N_28827,N_28985);
nor U29038 (N_29038,N_28750,N_28859);
xor U29039 (N_29039,N_28762,N_28856);
nor U29040 (N_29040,N_28929,N_28883);
or U29041 (N_29041,N_28968,N_28921);
or U29042 (N_29042,N_28959,N_28978);
nand U29043 (N_29043,N_28951,N_28916);
nand U29044 (N_29044,N_28781,N_28756);
or U29045 (N_29045,N_28928,N_28922);
or U29046 (N_29046,N_28953,N_28759);
and U29047 (N_29047,N_28829,N_28778);
and U29048 (N_29048,N_28802,N_28996);
xor U29049 (N_29049,N_28852,N_28758);
xor U29050 (N_29050,N_28851,N_28963);
xor U29051 (N_29051,N_28910,N_28886);
nand U29052 (N_29052,N_28981,N_28853);
or U29053 (N_29053,N_28824,N_28876);
xor U29054 (N_29054,N_28933,N_28849);
nor U29055 (N_29055,N_28974,N_28971);
nor U29056 (N_29056,N_28972,N_28848);
xor U29057 (N_29057,N_28908,N_28895);
nand U29058 (N_29058,N_28831,N_28815);
or U29059 (N_29059,N_28995,N_28751);
and U29060 (N_29060,N_28882,N_28768);
nor U29061 (N_29061,N_28760,N_28761);
nand U29062 (N_29062,N_28814,N_28792);
or U29063 (N_29063,N_28925,N_28991);
or U29064 (N_29064,N_28764,N_28812);
nand U29065 (N_29065,N_28898,N_28917);
xor U29066 (N_29066,N_28803,N_28874);
xor U29067 (N_29067,N_28977,N_28780);
or U29068 (N_29068,N_28911,N_28769);
xor U29069 (N_29069,N_28807,N_28975);
nand U29070 (N_29070,N_28930,N_28884);
and U29071 (N_29071,N_28931,N_28800);
nand U29072 (N_29072,N_28952,N_28976);
nand U29073 (N_29073,N_28896,N_28941);
and U29074 (N_29074,N_28818,N_28919);
or U29075 (N_29075,N_28775,N_28880);
and U29076 (N_29076,N_28920,N_28969);
nand U29077 (N_29077,N_28868,N_28878);
or U29078 (N_29078,N_28997,N_28863);
nand U29079 (N_29079,N_28772,N_28939);
and U29080 (N_29080,N_28765,N_28946);
xnor U29081 (N_29081,N_28964,N_28787);
xor U29082 (N_29082,N_28847,N_28855);
nand U29083 (N_29083,N_28885,N_28967);
xor U29084 (N_29084,N_28755,N_28955);
xnor U29085 (N_29085,N_28833,N_28810);
nor U29086 (N_29086,N_28854,N_28987);
or U29087 (N_29087,N_28913,N_28805);
nand U29088 (N_29088,N_28798,N_28782);
nor U29089 (N_29089,N_28909,N_28881);
nor U29090 (N_29090,N_28926,N_28773);
nor U29091 (N_29091,N_28842,N_28806);
xnor U29092 (N_29092,N_28808,N_28763);
and U29093 (N_29093,N_28770,N_28864);
nand U29094 (N_29094,N_28902,N_28838);
nor U29095 (N_29095,N_28861,N_28860);
xnor U29096 (N_29096,N_28757,N_28788);
xnor U29097 (N_29097,N_28809,N_28867);
and U29098 (N_29098,N_28958,N_28845);
nor U29099 (N_29099,N_28837,N_28924);
nand U29100 (N_29100,N_28905,N_28832);
or U29101 (N_29101,N_28984,N_28891);
and U29102 (N_29102,N_28839,N_28875);
nand U29103 (N_29103,N_28779,N_28822);
or U29104 (N_29104,N_28774,N_28857);
xor U29105 (N_29105,N_28899,N_28923);
and U29106 (N_29106,N_28828,N_28817);
nor U29107 (N_29107,N_28767,N_28789);
or U29108 (N_29108,N_28866,N_28970);
and U29109 (N_29109,N_28797,N_28820);
and U29110 (N_29110,N_28753,N_28825);
and U29111 (N_29111,N_28934,N_28998);
nand U29112 (N_29112,N_28850,N_28947);
or U29113 (N_29113,N_28784,N_28949);
nand U29114 (N_29114,N_28766,N_28948);
nor U29115 (N_29115,N_28858,N_28844);
and U29116 (N_29116,N_28869,N_28973);
xnor U29117 (N_29117,N_28945,N_28982);
xor U29118 (N_29118,N_28927,N_28862);
or U29119 (N_29119,N_28776,N_28888);
or U29120 (N_29120,N_28901,N_28894);
and U29121 (N_29121,N_28944,N_28990);
or U29122 (N_29122,N_28785,N_28938);
and U29123 (N_29123,N_28835,N_28887);
or U29124 (N_29124,N_28811,N_28950);
nor U29125 (N_29125,N_28896,N_28955);
nand U29126 (N_29126,N_28945,N_28885);
and U29127 (N_29127,N_28842,N_28816);
or U29128 (N_29128,N_28872,N_28925);
nor U29129 (N_29129,N_28863,N_28776);
or U29130 (N_29130,N_28814,N_28987);
nor U29131 (N_29131,N_28787,N_28932);
nand U29132 (N_29132,N_28913,N_28762);
nand U29133 (N_29133,N_28890,N_28968);
xnor U29134 (N_29134,N_28753,N_28986);
nor U29135 (N_29135,N_28850,N_28866);
or U29136 (N_29136,N_28882,N_28759);
nor U29137 (N_29137,N_28913,N_28998);
nand U29138 (N_29138,N_28797,N_28808);
xor U29139 (N_29139,N_28769,N_28762);
or U29140 (N_29140,N_28886,N_28971);
nand U29141 (N_29141,N_28941,N_28948);
or U29142 (N_29142,N_28951,N_28924);
xnor U29143 (N_29143,N_28964,N_28815);
nand U29144 (N_29144,N_28948,N_28754);
or U29145 (N_29145,N_28898,N_28965);
or U29146 (N_29146,N_28821,N_28938);
nand U29147 (N_29147,N_28778,N_28751);
nor U29148 (N_29148,N_28908,N_28998);
xnor U29149 (N_29149,N_28847,N_28853);
and U29150 (N_29150,N_28782,N_28795);
or U29151 (N_29151,N_28901,N_28921);
nor U29152 (N_29152,N_28881,N_28876);
nor U29153 (N_29153,N_28850,N_28986);
and U29154 (N_29154,N_28827,N_28990);
xnor U29155 (N_29155,N_28760,N_28886);
nor U29156 (N_29156,N_28875,N_28887);
and U29157 (N_29157,N_28912,N_28915);
or U29158 (N_29158,N_28754,N_28889);
nor U29159 (N_29159,N_28904,N_28851);
or U29160 (N_29160,N_28857,N_28896);
nor U29161 (N_29161,N_28926,N_28892);
nor U29162 (N_29162,N_28799,N_28981);
nand U29163 (N_29163,N_28929,N_28987);
or U29164 (N_29164,N_28835,N_28980);
and U29165 (N_29165,N_28792,N_28918);
and U29166 (N_29166,N_28904,N_28878);
nor U29167 (N_29167,N_28920,N_28994);
nor U29168 (N_29168,N_28978,N_28952);
xnor U29169 (N_29169,N_28979,N_28892);
nor U29170 (N_29170,N_28784,N_28787);
and U29171 (N_29171,N_28879,N_28834);
nand U29172 (N_29172,N_28944,N_28889);
or U29173 (N_29173,N_28879,N_28787);
nor U29174 (N_29174,N_28812,N_28943);
nor U29175 (N_29175,N_28787,N_28981);
nor U29176 (N_29176,N_28839,N_28760);
nor U29177 (N_29177,N_28818,N_28937);
xnor U29178 (N_29178,N_28907,N_28958);
nand U29179 (N_29179,N_28981,N_28841);
nor U29180 (N_29180,N_28968,N_28840);
and U29181 (N_29181,N_28969,N_28776);
nand U29182 (N_29182,N_28868,N_28879);
xnor U29183 (N_29183,N_28846,N_28887);
xor U29184 (N_29184,N_28964,N_28897);
or U29185 (N_29185,N_28800,N_28946);
nor U29186 (N_29186,N_28908,N_28802);
xnor U29187 (N_29187,N_28784,N_28894);
xnor U29188 (N_29188,N_28984,N_28785);
nand U29189 (N_29189,N_28771,N_28872);
nor U29190 (N_29190,N_28847,N_28807);
xor U29191 (N_29191,N_28831,N_28861);
or U29192 (N_29192,N_28997,N_28940);
xnor U29193 (N_29193,N_28987,N_28909);
and U29194 (N_29194,N_28890,N_28766);
nor U29195 (N_29195,N_28766,N_28908);
or U29196 (N_29196,N_28898,N_28786);
and U29197 (N_29197,N_28907,N_28772);
nand U29198 (N_29198,N_28962,N_28977);
and U29199 (N_29199,N_28841,N_28752);
nand U29200 (N_29200,N_28980,N_28942);
xor U29201 (N_29201,N_28991,N_28918);
nand U29202 (N_29202,N_28961,N_28806);
xnor U29203 (N_29203,N_28977,N_28928);
nor U29204 (N_29204,N_28915,N_28931);
or U29205 (N_29205,N_28770,N_28865);
or U29206 (N_29206,N_28809,N_28812);
or U29207 (N_29207,N_28853,N_28865);
nand U29208 (N_29208,N_28809,N_28778);
and U29209 (N_29209,N_28948,N_28852);
and U29210 (N_29210,N_28828,N_28879);
nor U29211 (N_29211,N_28839,N_28781);
or U29212 (N_29212,N_28980,N_28905);
nor U29213 (N_29213,N_28866,N_28830);
or U29214 (N_29214,N_28866,N_28877);
nand U29215 (N_29215,N_28783,N_28849);
or U29216 (N_29216,N_28910,N_28817);
nand U29217 (N_29217,N_28909,N_28936);
and U29218 (N_29218,N_28993,N_28845);
xnor U29219 (N_29219,N_28962,N_28875);
and U29220 (N_29220,N_28994,N_28901);
nor U29221 (N_29221,N_28920,N_28908);
or U29222 (N_29222,N_28811,N_28801);
nor U29223 (N_29223,N_28910,N_28777);
or U29224 (N_29224,N_28877,N_28937);
or U29225 (N_29225,N_28806,N_28753);
or U29226 (N_29226,N_28863,N_28798);
xnor U29227 (N_29227,N_28851,N_28886);
nor U29228 (N_29228,N_28788,N_28803);
xor U29229 (N_29229,N_28837,N_28788);
or U29230 (N_29230,N_28951,N_28939);
or U29231 (N_29231,N_28959,N_28907);
nand U29232 (N_29232,N_28962,N_28943);
xnor U29233 (N_29233,N_28812,N_28842);
or U29234 (N_29234,N_28827,N_28955);
nor U29235 (N_29235,N_28953,N_28850);
or U29236 (N_29236,N_28781,N_28977);
nor U29237 (N_29237,N_28883,N_28876);
nand U29238 (N_29238,N_28783,N_28885);
or U29239 (N_29239,N_28800,N_28974);
and U29240 (N_29240,N_28802,N_28978);
nor U29241 (N_29241,N_28762,N_28966);
xor U29242 (N_29242,N_28798,N_28937);
or U29243 (N_29243,N_28839,N_28919);
or U29244 (N_29244,N_28930,N_28855);
and U29245 (N_29245,N_28957,N_28851);
and U29246 (N_29246,N_28968,N_28913);
nand U29247 (N_29247,N_28989,N_28997);
and U29248 (N_29248,N_28937,N_28891);
xor U29249 (N_29249,N_28805,N_28841);
and U29250 (N_29250,N_29185,N_29050);
nand U29251 (N_29251,N_29119,N_29056);
and U29252 (N_29252,N_29061,N_29117);
or U29253 (N_29253,N_29113,N_29041);
or U29254 (N_29254,N_29149,N_29221);
or U29255 (N_29255,N_29093,N_29247);
xor U29256 (N_29256,N_29108,N_29168);
and U29257 (N_29257,N_29230,N_29223);
and U29258 (N_29258,N_29195,N_29210);
nor U29259 (N_29259,N_29123,N_29240);
and U29260 (N_29260,N_29073,N_29064);
xor U29261 (N_29261,N_29146,N_29044);
nor U29262 (N_29262,N_29095,N_29163);
nand U29263 (N_29263,N_29091,N_29155);
nand U29264 (N_29264,N_29085,N_29231);
nor U29265 (N_29265,N_29074,N_29014);
xnor U29266 (N_29266,N_29128,N_29054);
nand U29267 (N_29267,N_29200,N_29121);
xor U29268 (N_29268,N_29238,N_29244);
nor U29269 (N_29269,N_29015,N_29171);
nor U29270 (N_29270,N_29024,N_29191);
and U29271 (N_29271,N_29033,N_29190);
nand U29272 (N_29272,N_29241,N_29233);
nor U29273 (N_29273,N_29122,N_29236);
and U29274 (N_29274,N_29063,N_29109);
xor U29275 (N_29275,N_29013,N_29141);
nor U29276 (N_29276,N_29207,N_29177);
and U29277 (N_29277,N_29107,N_29226);
nand U29278 (N_29278,N_29138,N_29118);
nor U29279 (N_29279,N_29099,N_29018);
and U29280 (N_29280,N_29219,N_29048);
nor U29281 (N_29281,N_29178,N_29071);
and U29282 (N_29282,N_29017,N_29008);
xnor U29283 (N_29283,N_29016,N_29039);
nor U29284 (N_29284,N_29087,N_29145);
xnor U29285 (N_29285,N_29060,N_29235);
or U29286 (N_29286,N_29129,N_29058);
and U29287 (N_29287,N_29005,N_29172);
nand U29288 (N_29288,N_29088,N_29089);
or U29289 (N_29289,N_29237,N_29180);
nand U29290 (N_29290,N_29102,N_29007);
or U29291 (N_29291,N_29218,N_29246);
and U29292 (N_29292,N_29130,N_29051);
and U29293 (N_29293,N_29152,N_29096);
or U29294 (N_29294,N_29011,N_29182);
xor U29295 (N_29295,N_29143,N_29103);
xor U29296 (N_29296,N_29053,N_29194);
nor U29297 (N_29297,N_29181,N_29009);
or U29298 (N_29298,N_29112,N_29169);
or U29299 (N_29299,N_29214,N_29076);
nor U29300 (N_29300,N_29116,N_29010);
and U29301 (N_29301,N_29166,N_29057);
nand U29302 (N_29302,N_29106,N_29232);
xor U29303 (N_29303,N_29147,N_29153);
and U29304 (N_29304,N_29154,N_29249);
xor U29305 (N_29305,N_29126,N_29062);
nand U29306 (N_29306,N_29020,N_29183);
and U29307 (N_29307,N_29234,N_29225);
or U29308 (N_29308,N_29055,N_29125);
xor U29309 (N_29309,N_29227,N_29100);
xor U29310 (N_29310,N_29174,N_29204);
nor U29311 (N_29311,N_29111,N_29159);
or U29312 (N_29312,N_29066,N_29114);
nor U29313 (N_29313,N_29068,N_29000);
and U29314 (N_29314,N_29019,N_29037);
and U29315 (N_29315,N_29124,N_29160);
nand U29316 (N_29316,N_29031,N_29080);
and U29317 (N_29317,N_29150,N_29028);
nand U29318 (N_29318,N_29245,N_29025);
nand U29319 (N_29319,N_29196,N_29156);
or U29320 (N_29320,N_29032,N_29029);
and U29321 (N_29321,N_29094,N_29035);
nand U29322 (N_29322,N_29002,N_29110);
nand U29323 (N_29323,N_29078,N_29042);
or U29324 (N_29324,N_29248,N_29139);
xor U29325 (N_29325,N_29192,N_29133);
nor U29326 (N_29326,N_29215,N_29047);
and U29327 (N_29327,N_29187,N_29206);
nor U29328 (N_29328,N_29092,N_29097);
nand U29329 (N_29329,N_29229,N_29144);
xor U29330 (N_29330,N_29081,N_29217);
nor U29331 (N_29331,N_29189,N_29090);
xnor U29332 (N_29332,N_29083,N_29098);
nor U29333 (N_29333,N_29162,N_29069);
and U29334 (N_29334,N_29043,N_29164);
nor U29335 (N_29335,N_29201,N_29120);
or U29336 (N_29336,N_29030,N_29193);
nor U29337 (N_29337,N_29197,N_29115);
nor U29338 (N_29338,N_29127,N_29132);
nand U29339 (N_29339,N_29184,N_29198);
and U29340 (N_29340,N_29079,N_29101);
and U29341 (N_29341,N_29003,N_29158);
nand U29342 (N_29342,N_29173,N_29026);
and U29343 (N_29343,N_29075,N_29151);
and U29344 (N_29344,N_29176,N_29023);
or U29345 (N_29345,N_29165,N_29243);
xnor U29346 (N_29346,N_29065,N_29170);
and U29347 (N_29347,N_29213,N_29086);
xor U29348 (N_29348,N_29239,N_29208);
nand U29349 (N_29349,N_29228,N_29212);
or U29350 (N_29350,N_29186,N_29188);
or U29351 (N_29351,N_29049,N_29082);
and U29352 (N_29352,N_29211,N_29216);
xor U29353 (N_29353,N_29167,N_29203);
nor U29354 (N_29354,N_29072,N_29021);
nor U29355 (N_29355,N_29220,N_29222);
nand U29356 (N_29356,N_29135,N_29148);
and U29357 (N_29357,N_29209,N_29224);
xnor U29358 (N_29358,N_29004,N_29136);
and U29359 (N_29359,N_29045,N_29052);
nor U29360 (N_29360,N_29140,N_29006);
and U29361 (N_29361,N_29036,N_29104);
xor U29362 (N_29362,N_29067,N_29027);
nor U29363 (N_29363,N_29012,N_29161);
and U29364 (N_29364,N_29157,N_29038);
xnor U29365 (N_29365,N_29242,N_29040);
nor U29366 (N_29366,N_29175,N_29046);
nand U29367 (N_29367,N_29070,N_29179);
xnor U29368 (N_29368,N_29105,N_29084);
or U29369 (N_29369,N_29134,N_29034);
nor U29370 (N_29370,N_29077,N_29131);
and U29371 (N_29371,N_29205,N_29142);
and U29372 (N_29372,N_29059,N_29202);
xnor U29373 (N_29373,N_29001,N_29137);
and U29374 (N_29374,N_29022,N_29199);
nor U29375 (N_29375,N_29122,N_29063);
and U29376 (N_29376,N_29015,N_29195);
xor U29377 (N_29377,N_29225,N_29020);
nand U29378 (N_29378,N_29064,N_29130);
and U29379 (N_29379,N_29098,N_29100);
and U29380 (N_29380,N_29194,N_29168);
xnor U29381 (N_29381,N_29104,N_29081);
or U29382 (N_29382,N_29041,N_29135);
and U29383 (N_29383,N_29160,N_29042);
nor U29384 (N_29384,N_29105,N_29156);
xnor U29385 (N_29385,N_29049,N_29034);
xnor U29386 (N_29386,N_29245,N_29065);
nor U29387 (N_29387,N_29168,N_29059);
nand U29388 (N_29388,N_29072,N_29078);
nor U29389 (N_29389,N_29097,N_29172);
nand U29390 (N_29390,N_29010,N_29110);
nor U29391 (N_29391,N_29008,N_29163);
nand U29392 (N_29392,N_29182,N_29237);
xor U29393 (N_29393,N_29217,N_29014);
or U29394 (N_29394,N_29048,N_29180);
or U29395 (N_29395,N_29166,N_29008);
and U29396 (N_29396,N_29217,N_29136);
and U29397 (N_29397,N_29152,N_29125);
nand U29398 (N_29398,N_29213,N_29236);
xnor U29399 (N_29399,N_29043,N_29209);
nand U29400 (N_29400,N_29094,N_29149);
nand U29401 (N_29401,N_29083,N_29238);
nand U29402 (N_29402,N_29009,N_29223);
and U29403 (N_29403,N_29190,N_29215);
or U29404 (N_29404,N_29179,N_29182);
nand U29405 (N_29405,N_29045,N_29107);
or U29406 (N_29406,N_29204,N_29096);
nor U29407 (N_29407,N_29222,N_29196);
and U29408 (N_29408,N_29179,N_29233);
nand U29409 (N_29409,N_29081,N_29056);
or U29410 (N_29410,N_29103,N_29208);
xnor U29411 (N_29411,N_29154,N_29026);
or U29412 (N_29412,N_29246,N_29057);
nor U29413 (N_29413,N_29088,N_29234);
nor U29414 (N_29414,N_29022,N_29239);
xnor U29415 (N_29415,N_29237,N_29190);
or U29416 (N_29416,N_29082,N_29046);
xnor U29417 (N_29417,N_29115,N_29167);
and U29418 (N_29418,N_29039,N_29079);
or U29419 (N_29419,N_29137,N_29070);
or U29420 (N_29420,N_29065,N_29176);
nand U29421 (N_29421,N_29136,N_29117);
or U29422 (N_29422,N_29073,N_29238);
nor U29423 (N_29423,N_29247,N_29072);
and U29424 (N_29424,N_29200,N_29128);
xor U29425 (N_29425,N_29230,N_29090);
xnor U29426 (N_29426,N_29154,N_29213);
nand U29427 (N_29427,N_29183,N_29147);
nor U29428 (N_29428,N_29097,N_29117);
xnor U29429 (N_29429,N_29172,N_29111);
nand U29430 (N_29430,N_29022,N_29102);
xor U29431 (N_29431,N_29019,N_29002);
nor U29432 (N_29432,N_29023,N_29167);
nand U29433 (N_29433,N_29244,N_29221);
or U29434 (N_29434,N_29246,N_29185);
and U29435 (N_29435,N_29244,N_29186);
xnor U29436 (N_29436,N_29047,N_29032);
xnor U29437 (N_29437,N_29140,N_29131);
and U29438 (N_29438,N_29125,N_29242);
or U29439 (N_29439,N_29093,N_29106);
xnor U29440 (N_29440,N_29029,N_29072);
or U29441 (N_29441,N_29140,N_29018);
nand U29442 (N_29442,N_29094,N_29181);
or U29443 (N_29443,N_29246,N_29244);
or U29444 (N_29444,N_29224,N_29244);
nor U29445 (N_29445,N_29137,N_29158);
nand U29446 (N_29446,N_29059,N_29164);
nor U29447 (N_29447,N_29203,N_29110);
nor U29448 (N_29448,N_29142,N_29164);
xnor U29449 (N_29449,N_29105,N_29058);
xor U29450 (N_29450,N_29060,N_29105);
nand U29451 (N_29451,N_29084,N_29091);
and U29452 (N_29452,N_29036,N_29166);
nor U29453 (N_29453,N_29248,N_29022);
xnor U29454 (N_29454,N_29057,N_29198);
xnor U29455 (N_29455,N_29231,N_29158);
or U29456 (N_29456,N_29127,N_29086);
and U29457 (N_29457,N_29149,N_29238);
or U29458 (N_29458,N_29169,N_29096);
xor U29459 (N_29459,N_29210,N_29006);
and U29460 (N_29460,N_29142,N_29216);
and U29461 (N_29461,N_29184,N_29096);
nand U29462 (N_29462,N_29150,N_29080);
nor U29463 (N_29463,N_29155,N_29129);
and U29464 (N_29464,N_29223,N_29215);
nand U29465 (N_29465,N_29192,N_29082);
or U29466 (N_29466,N_29164,N_29239);
nor U29467 (N_29467,N_29076,N_29227);
nor U29468 (N_29468,N_29189,N_29017);
nor U29469 (N_29469,N_29238,N_29176);
and U29470 (N_29470,N_29232,N_29098);
xor U29471 (N_29471,N_29134,N_29169);
or U29472 (N_29472,N_29223,N_29193);
and U29473 (N_29473,N_29110,N_29031);
and U29474 (N_29474,N_29095,N_29187);
xor U29475 (N_29475,N_29104,N_29185);
or U29476 (N_29476,N_29067,N_29025);
xor U29477 (N_29477,N_29248,N_29118);
and U29478 (N_29478,N_29181,N_29017);
nor U29479 (N_29479,N_29186,N_29143);
nor U29480 (N_29480,N_29154,N_29130);
xor U29481 (N_29481,N_29009,N_29045);
nand U29482 (N_29482,N_29193,N_29005);
and U29483 (N_29483,N_29151,N_29145);
nor U29484 (N_29484,N_29055,N_29241);
xor U29485 (N_29485,N_29080,N_29212);
xor U29486 (N_29486,N_29034,N_29073);
nor U29487 (N_29487,N_29179,N_29096);
xnor U29488 (N_29488,N_29164,N_29127);
or U29489 (N_29489,N_29036,N_29095);
and U29490 (N_29490,N_29058,N_29138);
nand U29491 (N_29491,N_29193,N_29246);
nand U29492 (N_29492,N_29057,N_29237);
xnor U29493 (N_29493,N_29205,N_29099);
nand U29494 (N_29494,N_29029,N_29010);
nand U29495 (N_29495,N_29020,N_29093);
or U29496 (N_29496,N_29159,N_29065);
xnor U29497 (N_29497,N_29097,N_29212);
and U29498 (N_29498,N_29025,N_29044);
and U29499 (N_29499,N_29158,N_29086);
nand U29500 (N_29500,N_29419,N_29355);
and U29501 (N_29501,N_29330,N_29477);
nand U29502 (N_29502,N_29420,N_29277);
or U29503 (N_29503,N_29475,N_29497);
nor U29504 (N_29504,N_29486,N_29309);
and U29505 (N_29505,N_29401,N_29491);
nand U29506 (N_29506,N_29307,N_29364);
nand U29507 (N_29507,N_29451,N_29259);
nand U29508 (N_29508,N_29279,N_29343);
nor U29509 (N_29509,N_29255,N_29337);
xnor U29510 (N_29510,N_29263,N_29435);
nor U29511 (N_29511,N_29415,N_29427);
and U29512 (N_29512,N_29411,N_29288);
and U29513 (N_29513,N_29456,N_29294);
nand U29514 (N_29514,N_29315,N_29320);
xnor U29515 (N_29515,N_29302,N_29390);
nand U29516 (N_29516,N_29371,N_29374);
and U29517 (N_29517,N_29474,N_29322);
nand U29518 (N_29518,N_29421,N_29382);
nand U29519 (N_29519,N_29430,N_29453);
nor U29520 (N_29520,N_29447,N_29373);
nor U29521 (N_29521,N_29352,N_29327);
nand U29522 (N_29522,N_29338,N_29264);
and U29523 (N_29523,N_29490,N_29344);
xnor U29524 (N_29524,N_29367,N_29360);
and U29525 (N_29525,N_29462,N_29299);
and U29526 (N_29526,N_29296,N_29471);
or U29527 (N_29527,N_29339,N_29481);
or U29528 (N_29528,N_29312,N_29458);
xor U29529 (N_29529,N_29250,N_29479);
nor U29530 (N_29530,N_29267,N_29341);
and U29531 (N_29531,N_29356,N_29410);
or U29532 (N_29532,N_29304,N_29325);
nand U29533 (N_29533,N_29256,N_29293);
nor U29534 (N_29534,N_29448,N_29345);
nand U29535 (N_29535,N_29386,N_29489);
or U29536 (N_29536,N_29400,N_29380);
or U29537 (N_29537,N_29464,N_29314);
nand U29538 (N_29538,N_29383,N_29463);
and U29539 (N_29539,N_29340,N_29377);
and U29540 (N_29540,N_29289,N_29283);
and U29541 (N_29541,N_29482,N_29287);
xnor U29542 (N_29542,N_29442,N_29336);
nand U29543 (N_29543,N_29441,N_29426);
nor U29544 (N_29544,N_29365,N_29413);
and U29545 (N_29545,N_29412,N_29466);
and U29546 (N_29546,N_29303,N_29317);
or U29547 (N_29547,N_29284,N_29408);
and U29548 (N_29548,N_29372,N_29483);
and U29549 (N_29549,N_29359,N_29273);
or U29550 (N_29550,N_29271,N_29472);
or U29551 (N_29551,N_29282,N_29258);
and U29552 (N_29552,N_29403,N_29381);
or U29553 (N_29553,N_29478,N_29260);
nand U29554 (N_29554,N_29457,N_29487);
nand U29555 (N_29555,N_29286,N_29459);
xor U29556 (N_29556,N_29261,N_29370);
nand U29557 (N_29557,N_29305,N_29342);
xnor U29558 (N_29558,N_29333,N_29353);
or U29559 (N_29559,N_29358,N_29285);
nor U29560 (N_29560,N_29366,N_29484);
xor U29561 (N_29561,N_29300,N_29349);
nand U29562 (N_29562,N_29266,N_29473);
or U29563 (N_29563,N_29280,N_29298);
nor U29564 (N_29564,N_29375,N_29402);
nand U29565 (N_29565,N_29319,N_29318);
and U29566 (N_29566,N_29297,N_29436);
nand U29567 (N_29567,N_29492,N_29423);
nand U29568 (N_29568,N_29424,N_29440);
xnor U29569 (N_29569,N_29398,N_29399);
nor U29570 (N_29570,N_29392,N_29445);
xnor U29571 (N_29571,N_29384,N_29379);
xnor U29572 (N_29572,N_29272,N_29452);
nor U29573 (N_29573,N_29437,N_29499);
nand U29574 (N_29574,N_29488,N_29389);
or U29575 (N_29575,N_29417,N_29308);
xor U29576 (N_29576,N_29433,N_29316);
or U29577 (N_29577,N_29251,N_29265);
xor U29578 (N_29578,N_29257,N_29311);
or U29579 (N_29579,N_29439,N_29495);
and U29580 (N_29580,N_29268,N_29388);
nor U29581 (N_29581,N_29444,N_29357);
nand U29582 (N_29582,N_29476,N_29429);
or U29583 (N_29583,N_29404,N_29274);
xnor U29584 (N_29584,N_29281,N_29460);
nand U29585 (N_29585,N_29465,N_29480);
or U29586 (N_29586,N_29493,N_29438);
or U29587 (N_29587,N_29295,N_29292);
nor U29588 (N_29588,N_29310,N_29394);
and U29589 (N_29589,N_29498,N_29469);
or U29590 (N_29590,N_29306,N_29414);
nand U29591 (N_29591,N_29328,N_29335);
nand U29592 (N_29592,N_29431,N_29406);
xor U29593 (N_29593,N_29334,N_29378);
nor U29594 (N_29594,N_29253,N_29350);
and U29595 (N_29595,N_29395,N_29409);
nor U29596 (N_29596,N_29324,N_29363);
nand U29597 (N_29597,N_29276,N_29354);
nand U29598 (N_29598,N_29494,N_29275);
xnor U29599 (N_29599,N_29291,N_29290);
nand U29600 (N_29600,N_29301,N_29262);
xor U29601 (N_29601,N_29362,N_29270);
or U29602 (N_29602,N_29351,N_29332);
nand U29603 (N_29603,N_29252,N_29269);
nor U29604 (N_29604,N_29329,N_29361);
xnor U29605 (N_29605,N_29323,N_29455);
and U29606 (N_29606,N_29434,N_29313);
nand U29607 (N_29607,N_29443,N_29331);
and U29608 (N_29608,N_29449,N_29346);
xnor U29609 (N_29609,N_29397,N_29428);
nand U29610 (N_29610,N_29391,N_29278);
nand U29611 (N_29611,N_29461,N_29418);
and U29612 (N_29612,N_29446,N_29468);
xor U29613 (N_29613,N_29369,N_29422);
nor U29614 (N_29614,N_29321,N_29393);
nand U29615 (N_29615,N_29485,N_29467);
nor U29616 (N_29616,N_29376,N_29450);
or U29617 (N_29617,N_29416,N_29387);
or U29618 (N_29618,N_29396,N_29347);
and U29619 (N_29619,N_29432,N_29470);
xnor U29620 (N_29620,N_29326,N_29368);
and U29621 (N_29621,N_29454,N_29425);
and U29622 (N_29622,N_29405,N_29348);
nor U29623 (N_29623,N_29407,N_29385);
nand U29624 (N_29624,N_29496,N_29254);
xor U29625 (N_29625,N_29477,N_29288);
xnor U29626 (N_29626,N_29304,N_29254);
nand U29627 (N_29627,N_29370,N_29373);
or U29628 (N_29628,N_29425,N_29338);
nand U29629 (N_29629,N_29332,N_29423);
nand U29630 (N_29630,N_29374,N_29386);
and U29631 (N_29631,N_29350,N_29469);
nor U29632 (N_29632,N_29426,N_29489);
or U29633 (N_29633,N_29482,N_29499);
nor U29634 (N_29634,N_29464,N_29301);
nand U29635 (N_29635,N_29453,N_29360);
and U29636 (N_29636,N_29458,N_29459);
or U29637 (N_29637,N_29263,N_29367);
nand U29638 (N_29638,N_29396,N_29409);
or U29639 (N_29639,N_29325,N_29443);
or U29640 (N_29640,N_29428,N_29317);
and U29641 (N_29641,N_29369,N_29432);
nand U29642 (N_29642,N_29320,N_29380);
nand U29643 (N_29643,N_29470,N_29324);
nor U29644 (N_29644,N_29352,N_29435);
and U29645 (N_29645,N_29343,N_29271);
xnor U29646 (N_29646,N_29488,N_29452);
nor U29647 (N_29647,N_29390,N_29493);
and U29648 (N_29648,N_29311,N_29338);
nor U29649 (N_29649,N_29410,N_29346);
nor U29650 (N_29650,N_29346,N_29280);
xnor U29651 (N_29651,N_29253,N_29287);
or U29652 (N_29652,N_29401,N_29380);
xor U29653 (N_29653,N_29438,N_29338);
or U29654 (N_29654,N_29439,N_29370);
and U29655 (N_29655,N_29279,N_29440);
or U29656 (N_29656,N_29359,N_29394);
or U29657 (N_29657,N_29363,N_29348);
xor U29658 (N_29658,N_29410,N_29260);
or U29659 (N_29659,N_29345,N_29462);
nor U29660 (N_29660,N_29334,N_29403);
or U29661 (N_29661,N_29437,N_29445);
xor U29662 (N_29662,N_29435,N_29392);
xnor U29663 (N_29663,N_29419,N_29296);
xor U29664 (N_29664,N_29334,N_29444);
nand U29665 (N_29665,N_29345,N_29256);
nand U29666 (N_29666,N_29396,N_29326);
and U29667 (N_29667,N_29365,N_29355);
nand U29668 (N_29668,N_29343,N_29432);
nand U29669 (N_29669,N_29365,N_29264);
and U29670 (N_29670,N_29269,N_29285);
nand U29671 (N_29671,N_29425,N_29491);
and U29672 (N_29672,N_29374,N_29490);
xnor U29673 (N_29673,N_29348,N_29297);
xnor U29674 (N_29674,N_29444,N_29375);
nand U29675 (N_29675,N_29490,N_29363);
nor U29676 (N_29676,N_29335,N_29344);
and U29677 (N_29677,N_29442,N_29315);
xor U29678 (N_29678,N_29387,N_29317);
and U29679 (N_29679,N_29286,N_29423);
nand U29680 (N_29680,N_29368,N_29287);
or U29681 (N_29681,N_29336,N_29401);
nor U29682 (N_29682,N_29481,N_29315);
or U29683 (N_29683,N_29274,N_29336);
nand U29684 (N_29684,N_29348,N_29487);
and U29685 (N_29685,N_29250,N_29405);
nor U29686 (N_29686,N_29328,N_29258);
or U29687 (N_29687,N_29480,N_29367);
nand U29688 (N_29688,N_29252,N_29497);
or U29689 (N_29689,N_29368,N_29332);
xor U29690 (N_29690,N_29347,N_29412);
nand U29691 (N_29691,N_29271,N_29412);
and U29692 (N_29692,N_29419,N_29461);
nand U29693 (N_29693,N_29448,N_29287);
or U29694 (N_29694,N_29262,N_29434);
nand U29695 (N_29695,N_29253,N_29474);
nor U29696 (N_29696,N_29360,N_29254);
and U29697 (N_29697,N_29358,N_29399);
or U29698 (N_29698,N_29384,N_29424);
nor U29699 (N_29699,N_29312,N_29371);
or U29700 (N_29700,N_29272,N_29284);
nor U29701 (N_29701,N_29488,N_29416);
nand U29702 (N_29702,N_29402,N_29495);
and U29703 (N_29703,N_29354,N_29331);
or U29704 (N_29704,N_29283,N_29399);
or U29705 (N_29705,N_29377,N_29394);
and U29706 (N_29706,N_29486,N_29350);
or U29707 (N_29707,N_29289,N_29273);
xor U29708 (N_29708,N_29410,N_29355);
and U29709 (N_29709,N_29377,N_29416);
nor U29710 (N_29710,N_29265,N_29433);
nand U29711 (N_29711,N_29270,N_29431);
nor U29712 (N_29712,N_29285,N_29421);
nand U29713 (N_29713,N_29346,N_29363);
xor U29714 (N_29714,N_29424,N_29429);
or U29715 (N_29715,N_29325,N_29335);
nand U29716 (N_29716,N_29463,N_29467);
xor U29717 (N_29717,N_29441,N_29412);
xnor U29718 (N_29718,N_29304,N_29335);
nor U29719 (N_29719,N_29457,N_29397);
xor U29720 (N_29720,N_29407,N_29452);
and U29721 (N_29721,N_29430,N_29469);
nor U29722 (N_29722,N_29338,N_29381);
or U29723 (N_29723,N_29452,N_29498);
or U29724 (N_29724,N_29437,N_29389);
xor U29725 (N_29725,N_29268,N_29455);
nand U29726 (N_29726,N_29428,N_29480);
or U29727 (N_29727,N_29314,N_29499);
nand U29728 (N_29728,N_29292,N_29466);
xnor U29729 (N_29729,N_29409,N_29346);
xor U29730 (N_29730,N_29279,N_29459);
nor U29731 (N_29731,N_29323,N_29345);
nand U29732 (N_29732,N_29339,N_29455);
and U29733 (N_29733,N_29447,N_29390);
xnor U29734 (N_29734,N_29448,N_29296);
xor U29735 (N_29735,N_29324,N_29490);
xor U29736 (N_29736,N_29441,N_29480);
nand U29737 (N_29737,N_29335,N_29389);
nor U29738 (N_29738,N_29316,N_29325);
or U29739 (N_29739,N_29292,N_29339);
nor U29740 (N_29740,N_29338,N_29409);
and U29741 (N_29741,N_29401,N_29369);
or U29742 (N_29742,N_29306,N_29394);
xnor U29743 (N_29743,N_29326,N_29259);
nor U29744 (N_29744,N_29448,N_29259);
xnor U29745 (N_29745,N_29320,N_29265);
nand U29746 (N_29746,N_29274,N_29288);
nand U29747 (N_29747,N_29344,N_29275);
and U29748 (N_29748,N_29306,N_29449);
nand U29749 (N_29749,N_29278,N_29267);
and U29750 (N_29750,N_29615,N_29613);
and U29751 (N_29751,N_29527,N_29545);
nor U29752 (N_29752,N_29539,N_29661);
or U29753 (N_29753,N_29556,N_29590);
xnor U29754 (N_29754,N_29506,N_29640);
and U29755 (N_29755,N_29658,N_29604);
xnor U29756 (N_29756,N_29690,N_29507);
nor U29757 (N_29757,N_29683,N_29738);
nand U29758 (N_29758,N_29559,N_29747);
nor U29759 (N_29759,N_29538,N_29575);
or U29760 (N_29760,N_29515,N_29706);
and U29761 (N_29761,N_29607,N_29555);
nand U29762 (N_29762,N_29655,N_29566);
xor U29763 (N_29763,N_29645,N_29509);
and U29764 (N_29764,N_29510,N_29584);
or U29765 (N_29765,N_29586,N_29562);
and U29766 (N_29766,N_29558,N_29668);
xnor U29767 (N_29767,N_29550,N_29730);
and U29768 (N_29768,N_29712,N_29621);
or U29769 (N_29769,N_29508,N_29720);
nor U29770 (N_29770,N_29696,N_29517);
nand U29771 (N_29771,N_29749,N_29564);
nor U29772 (N_29772,N_29600,N_29560);
nand U29773 (N_29773,N_29577,N_29744);
and U29774 (N_29774,N_29695,N_29561);
nand U29775 (N_29775,N_29525,N_29647);
nor U29776 (N_29776,N_29606,N_29500);
nor U29777 (N_29777,N_29589,N_29673);
nor U29778 (N_29778,N_29503,N_29609);
nand U29779 (N_29779,N_29588,N_29631);
or U29780 (N_29780,N_29724,N_29654);
nor U29781 (N_29781,N_29674,N_29521);
xor U29782 (N_29782,N_29578,N_29522);
and U29783 (N_29783,N_29530,N_29691);
or U29784 (N_29784,N_29568,N_29627);
nor U29785 (N_29785,N_29714,N_29628);
or U29786 (N_29786,N_29703,N_29697);
nand U29787 (N_29787,N_29701,N_29520);
nor U29788 (N_29788,N_29549,N_29667);
nor U29789 (N_29789,N_29599,N_29644);
xor U29790 (N_29790,N_29651,N_29502);
and U29791 (N_29791,N_29534,N_29659);
nand U29792 (N_29792,N_29572,N_29686);
nand U29793 (N_29793,N_29698,N_29685);
xor U29794 (N_29794,N_29597,N_29657);
xor U29795 (N_29795,N_29596,N_29618);
and U29796 (N_29796,N_29602,N_29633);
or U29797 (N_29797,N_29652,N_29543);
nor U29798 (N_29798,N_29565,N_29646);
nand U29799 (N_29799,N_29732,N_29595);
and U29800 (N_29800,N_29582,N_29721);
and U29801 (N_29801,N_29671,N_29605);
nor U29802 (N_29802,N_29725,N_29643);
or U29803 (N_29803,N_29684,N_29537);
nor U29804 (N_29804,N_29635,N_29514);
nand U29805 (N_29805,N_29603,N_29563);
nand U29806 (N_29806,N_29569,N_29501);
or U29807 (N_29807,N_29532,N_29663);
nor U29808 (N_29808,N_29580,N_29648);
nand U29809 (N_29809,N_29719,N_29629);
nor U29810 (N_29810,N_29702,N_29745);
or U29811 (N_29811,N_29601,N_29664);
xnor U29812 (N_29812,N_29634,N_29529);
nand U29813 (N_29813,N_29708,N_29662);
nand U29814 (N_29814,N_29598,N_29593);
nand U29815 (N_29815,N_29626,N_29611);
nor U29816 (N_29816,N_29675,N_29610);
or U29817 (N_29817,N_29710,N_29734);
nand U29818 (N_29818,N_29587,N_29666);
or U29819 (N_29819,N_29622,N_29672);
xnor U29820 (N_29820,N_29699,N_29669);
xor U29821 (N_29821,N_29709,N_29705);
nor U29822 (N_29822,N_29694,N_29692);
xnor U29823 (N_29823,N_29579,N_29625);
or U29824 (N_29824,N_29524,N_29612);
or U29825 (N_29825,N_29739,N_29670);
xor U29826 (N_29826,N_29638,N_29553);
nor U29827 (N_29827,N_29735,N_29642);
nand U29828 (N_29828,N_29571,N_29707);
nand U29829 (N_29829,N_29542,N_29729);
xor U29830 (N_29830,N_29704,N_29536);
nor U29831 (N_29831,N_29693,N_29742);
nor U29832 (N_29832,N_29570,N_29544);
and U29833 (N_29833,N_29726,N_29665);
or U29834 (N_29834,N_29504,N_29574);
xor U29835 (N_29835,N_29619,N_29741);
xor U29836 (N_29836,N_29614,N_29743);
nor U29837 (N_29837,N_29649,N_29608);
nor U29838 (N_29838,N_29722,N_29748);
nor U29839 (N_29839,N_29637,N_29678);
and U29840 (N_29840,N_29681,N_29513);
xor U29841 (N_29841,N_29576,N_29740);
xor U29842 (N_29842,N_29591,N_29526);
nand U29843 (N_29843,N_29523,N_29736);
xor U29844 (N_29844,N_29727,N_29528);
xor U29845 (N_29845,N_29567,N_29746);
and U29846 (N_29846,N_29656,N_29723);
xnor U29847 (N_29847,N_29592,N_29680);
and U29848 (N_29848,N_29676,N_29689);
and U29849 (N_29849,N_29511,N_29554);
nor U29850 (N_29850,N_29679,N_29541);
xor U29851 (N_29851,N_29639,N_29518);
nand U29852 (N_29852,N_29731,N_29713);
nor U29853 (N_29853,N_29733,N_29505);
or U29854 (N_29854,N_29546,N_29548);
or U29855 (N_29855,N_29630,N_29653);
and U29856 (N_29856,N_29716,N_29688);
xor U29857 (N_29857,N_29616,N_29516);
or U29858 (N_29858,N_29718,N_29583);
nor U29859 (N_29859,N_29519,N_29557);
or U29860 (N_29860,N_29677,N_29623);
nor U29861 (N_29861,N_29552,N_29641);
xor U29862 (N_29862,N_29594,N_29617);
or U29863 (N_29863,N_29547,N_29715);
and U29864 (N_29864,N_29700,N_29711);
nand U29865 (N_29865,N_29650,N_29531);
nor U29866 (N_29866,N_29687,N_29636);
xnor U29867 (N_29867,N_29551,N_29585);
nand U29868 (N_29868,N_29533,N_29728);
or U29869 (N_29869,N_29573,N_29632);
nor U29870 (N_29870,N_29512,N_29540);
and U29871 (N_29871,N_29535,N_29620);
nor U29872 (N_29872,N_29737,N_29660);
or U29873 (N_29873,N_29581,N_29624);
nor U29874 (N_29874,N_29682,N_29717);
nand U29875 (N_29875,N_29521,N_29628);
nand U29876 (N_29876,N_29652,N_29609);
and U29877 (N_29877,N_29671,N_29518);
nor U29878 (N_29878,N_29651,N_29711);
or U29879 (N_29879,N_29621,N_29706);
xnor U29880 (N_29880,N_29522,N_29628);
nand U29881 (N_29881,N_29663,N_29668);
nor U29882 (N_29882,N_29594,N_29504);
nand U29883 (N_29883,N_29744,N_29664);
xnor U29884 (N_29884,N_29611,N_29627);
and U29885 (N_29885,N_29688,N_29746);
nor U29886 (N_29886,N_29666,N_29737);
nor U29887 (N_29887,N_29527,N_29735);
and U29888 (N_29888,N_29613,N_29568);
and U29889 (N_29889,N_29664,N_29597);
nor U29890 (N_29890,N_29674,N_29682);
or U29891 (N_29891,N_29625,N_29732);
nand U29892 (N_29892,N_29528,N_29609);
nand U29893 (N_29893,N_29627,N_29692);
xnor U29894 (N_29894,N_29647,N_29539);
nor U29895 (N_29895,N_29743,N_29654);
and U29896 (N_29896,N_29554,N_29710);
nor U29897 (N_29897,N_29591,N_29679);
xor U29898 (N_29898,N_29735,N_29672);
nand U29899 (N_29899,N_29734,N_29671);
xor U29900 (N_29900,N_29587,N_29594);
nand U29901 (N_29901,N_29563,N_29697);
nand U29902 (N_29902,N_29560,N_29645);
and U29903 (N_29903,N_29614,N_29719);
or U29904 (N_29904,N_29538,N_29748);
nor U29905 (N_29905,N_29613,N_29690);
nand U29906 (N_29906,N_29698,N_29591);
or U29907 (N_29907,N_29641,N_29626);
and U29908 (N_29908,N_29723,N_29591);
or U29909 (N_29909,N_29665,N_29731);
nand U29910 (N_29910,N_29718,N_29621);
nand U29911 (N_29911,N_29504,N_29650);
nand U29912 (N_29912,N_29729,N_29725);
nand U29913 (N_29913,N_29712,N_29571);
and U29914 (N_29914,N_29599,N_29555);
or U29915 (N_29915,N_29728,N_29609);
and U29916 (N_29916,N_29573,N_29588);
nand U29917 (N_29917,N_29724,N_29678);
nor U29918 (N_29918,N_29621,N_29534);
or U29919 (N_29919,N_29635,N_29625);
or U29920 (N_29920,N_29530,N_29717);
nand U29921 (N_29921,N_29601,N_29617);
or U29922 (N_29922,N_29667,N_29671);
or U29923 (N_29923,N_29575,N_29582);
xor U29924 (N_29924,N_29721,N_29733);
and U29925 (N_29925,N_29548,N_29627);
and U29926 (N_29926,N_29709,N_29517);
nand U29927 (N_29927,N_29587,N_29726);
xnor U29928 (N_29928,N_29584,N_29733);
nor U29929 (N_29929,N_29560,N_29502);
or U29930 (N_29930,N_29624,N_29631);
nor U29931 (N_29931,N_29622,N_29682);
nor U29932 (N_29932,N_29683,N_29540);
nor U29933 (N_29933,N_29534,N_29718);
nor U29934 (N_29934,N_29739,N_29642);
and U29935 (N_29935,N_29611,N_29747);
nand U29936 (N_29936,N_29600,N_29530);
nand U29937 (N_29937,N_29598,N_29530);
xor U29938 (N_29938,N_29727,N_29601);
and U29939 (N_29939,N_29632,N_29617);
xor U29940 (N_29940,N_29736,N_29620);
nand U29941 (N_29941,N_29519,N_29500);
or U29942 (N_29942,N_29735,N_29573);
and U29943 (N_29943,N_29741,N_29563);
nand U29944 (N_29944,N_29628,N_29528);
nor U29945 (N_29945,N_29749,N_29583);
nand U29946 (N_29946,N_29657,N_29524);
nand U29947 (N_29947,N_29721,N_29511);
and U29948 (N_29948,N_29690,N_29691);
nand U29949 (N_29949,N_29545,N_29648);
nor U29950 (N_29950,N_29634,N_29647);
nor U29951 (N_29951,N_29665,N_29518);
nand U29952 (N_29952,N_29732,N_29654);
nand U29953 (N_29953,N_29634,N_29668);
nor U29954 (N_29954,N_29507,N_29524);
nand U29955 (N_29955,N_29686,N_29632);
xnor U29956 (N_29956,N_29678,N_29571);
nor U29957 (N_29957,N_29677,N_29551);
nand U29958 (N_29958,N_29641,N_29616);
nor U29959 (N_29959,N_29505,N_29509);
or U29960 (N_29960,N_29717,N_29616);
nand U29961 (N_29961,N_29574,N_29526);
nor U29962 (N_29962,N_29672,N_29634);
nor U29963 (N_29963,N_29746,N_29732);
nor U29964 (N_29964,N_29661,N_29700);
or U29965 (N_29965,N_29562,N_29589);
or U29966 (N_29966,N_29549,N_29640);
xor U29967 (N_29967,N_29732,N_29749);
and U29968 (N_29968,N_29578,N_29642);
xor U29969 (N_29969,N_29591,N_29596);
or U29970 (N_29970,N_29518,N_29675);
nor U29971 (N_29971,N_29603,N_29552);
nor U29972 (N_29972,N_29559,N_29711);
nor U29973 (N_29973,N_29559,N_29606);
or U29974 (N_29974,N_29540,N_29520);
xor U29975 (N_29975,N_29685,N_29513);
or U29976 (N_29976,N_29618,N_29569);
xnor U29977 (N_29977,N_29669,N_29665);
or U29978 (N_29978,N_29719,N_29630);
nand U29979 (N_29979,N_29601,N_29679);
and U29980 (N_29980,N_29730,N_29585);
xor U29981 (N_29981,N_29705,N_29702);
and U29982 (N_29982,N_29720,N_29648);
xor U29983 (N_29983,N_29589,N_29708);
xor U29984 (N_29984,N_29546,N_29575);
nand U29985 (N_29985,N_29637,N_29546);
xor U29986 (N_29986,N_29591,N_29554);
nand U29987 (N_29987,N_29644,N_29681);
or U29988 (N_29988,N_29605,N_29639);
xor U29989 (N_29989,N_29510,N_29536);
and U29990 (N_29990,N_29726,N_29580);
or U29991 (N_29991,N_29631,N_29748);
nor U29992 (N_29992,N_29726,N_29511);
nand U29993 (N_29993,N_29571,N_29565);
or U29994 (N_29994,N_29648,N_29588);
nand U29995 (N_29995,N_29578,N_29537);
nor U29996 (N_29996,N_29576,N_29516);
and U29997 (N_29997,N_29692,N_29535);
and U29998 (N_29998,N_29575,N_29674);
and U29999 (N_29999,N_29548,N_29551);
or U30000 (N_30000,N_29975,N_29953);
and U30001 (N_30001,N_29858,N_29819);
or U30002 (N_30002,N_29963,N_29883);
and U30003 (N_30003,N_29766,N_29967);
or U30004 (N_30004,N_29917,N_29802);
nor U30005 (N_30005,N_29801,N_29970);
and U30006 (N_30006,N_29811,N_29929);
and U30007 (N_30007,N_29979,N_29793);
nor U30008 (N_30008,N_29927,N_29770);
nor U30009 (N_30009,N_29895,N_29807);
and U30010 (N_30010,N_29789,N_29922);
nor U30011 (N_30011,N_29936,N_29836);
or U30012 (N_30012,N_29812,N_29885);
nand U30013 (N_30013,N_29792,N_29939);
nor U30014 (N_30014,N_29839,N_29956);
nor U30015 (N_30015,N_29901,N_29850);
xnor U30016 (N_30016,N_29930,N_29750);
nand U30017 (N_30017,N_29889,N_29938);
or U30018 (N_30018,N_29906,N_29842);
nand U30019 (N_30019,N_29997,N_29908);
xor U30020 (N_30020,N_29892,N_29940);
or U30021 (N_30021,N_29969,N_29759);
nand U30022 (N_30022,N_29968,N_29844);
nor U30023 (N_30023,N_29863,N_29871);
nand U30024 (N_30024,N_29809,N_29830);
and U30025 (N_30025,N_29952,N_29964);
or U30026 (N_30026,N_29757,N_29834);
xnor U30027 (N_30027,N_29902,N_29851);
and U30028 (N_30028,N_29904,N_29914);
nand U30029 (N_30029,N_29852,N_29794);
and U30030 (N_30030,N_29762,N_29881);
nor U30031 (N_30031,N_29983,N_29980);
or U30032 (N_30032,N_29974,N_29993);
xor U30033 (N_30033,N_29804,N_29905);
or U30034 (N_30034,N_29976,N_29783);
xor U30035 (N_30035,N_29767,N_29948);
nand U30036 (N_30036,N_29873,N_29884);
or U30037 (N_30037,N_29821,N_29788);
xor U30038 (N_30038,N_29806,N_29928);
nand U30039 (N_30039,N_29896,N_29916);
and U30040 (N_30040,N_29787,N_29826);
nor U30041 (N_30041,N_29808,N_29876);
and U30042 (N_30042,N_29995,N_29988);
nand U30043 (N_30043,N_29846,N_29986);
and U30044 (N_30044,N_29875,N_29822);
xor U30045 (N_30045,N_29773,N_29751);
nand U30046 (N_30046,N_29778,N_29814);
and U30047 (N_30047,N_29820,N_29756);
and U30048 (N_30048,N_29894,N_29942);
xnor U30049 (N_30049,N_29992,N_29944);
xor U30050 (N_30050,N_29754,N_29775);
nor U30051 (N_30051,N_29990,N_29903);
or U30052 (N_30052,N_29972,N_29998);
nor U30053 (N_30053,N_29941,N_29932);
nand U30054 (N_30054,N_29829,N_29860);
nor U30055 (N_30055,N_29982,N_29978);
xor U30056 (N_30056,N_29849,N_29973);
nor U30057 (N_30057,N_29769,N_29985);
and U30058 (N_30058,N_29877,N_29813);
nand U30059 (N_30059,N_29874,N_29843);
nand U30060 (N_30060,N_29961,N_29828);
xnor U30061 (N_30061,N_29818,N_29947);
and U30062 (N_30062,N_29845,N_29886);
and U30063 (N_30063,N_29795,N_29887);
nor U30064 (N_30064,N_29955,N_29785);
nor U30065 (N_30065,N_29933,N_29893);
xor U30066 (N_30066,N_29924,N_29923);
and U30067 (N_30067,N_29891,N_29919);
nor U30068 (N_30068,N_29921,N_29999);
xor U30069 (N_30069,N_29866,N_29833);
and U30070 (N_30070,N_29797,N_29780);
or U30071 (N_30071,N_29847,N_29774);
and U30072 (N_30072,N_29989,N_29925);
or U30073 (N_30073,N_29864,N_29765);
xor U30074 (N_30074,N_29880,N_29816);
and U30075 (N_30075,N_29915,N_29878);
nand U30076 (N_30076,N_29946,N_29817);
nand U30077 (N_30077,N_29782,N_29959);
nand U30078 (N_30078,N_29758,N_29753);
and U30079 (N_30079,N_29805,N_29958);
or U30080 (N_30080,N_29865,N_29779);
nand U30081 (N_30081,N_29838,N_29987);
xnor U30082 (N_30082,N_29768,N_29862);
nor U30083 (N_30083,N_29911,N_29869);
nor U30084 (N_30084,N_29771,N_29888);
or U30085 (N_30085,N_29790,N_29763);
nor U30086 (N_30086,N_29996,N_29784);
nor U30087 (N_30087,N_29832,N_29837);
or U30088 (N_30088,N_29831,N_29760);
and U30089 (N_30089,N_29912,N_29772);
nand U30090 (N_30090,N_29781,N_29854);
nand U30091 (N_30091,N_29800,N_29909);
xnor U30092 (N_30092,N_29823,N_29868);
xnor U30093 (N_30093,N_29841,N_29951);
xnor U30094 (N_30094,N_29994,N_29810);
or U30095 (N_30095,N_29950,N_29899);
nor U30096 (N_30096,N_29949,N_29848);
nand U30097 (N_30097,N_29957,N_29855);
nand U30098 (N_30098,N_29943,N_29977);
or U30099 (N_30099,N_29962,N_29752);
xnor U30100 (N_30100,N_29890,N_29966);
and U30101 (N_30101,N_29920,N_29861);
xnor U30102 (N_30102,N_29965,N_29761);
nand U30103 (N_30103,N_29825,N_29857);
or U30104 (N_30104,N_29776,N_29853);
nand U30105 (N_30105,N_29926,N_29799);
nand U30106 (N_30106,N_29897,N_29910);
nor U30107 (N_30107,N_29913,N_29918);
and U30108 (N_30108,N_29764,N_29945);
nand U30109 (N_30109,N_29824,N_29856);
xor U30110 (N_30110,N_29835,N_29900);
or U30111 (N_30111,N_29971,N_29867);
nor U30112 (N_30112,N_29879,N_29859);
nor U30113 (N_30113,N_29934,N_29907);
or U30114 (N_30114,N_29796,N_29755);
and U30115 (N_30115,N_29786,N_29803);
or U30116 (N_30116,N_29991,N_29870);
nand U30117 (N_30117,N_29827,N_29815);
or U30118 (N_30118,N_29840,N_29882);
and U30119 (N_30119,N_29954,N_29937);
nand U30120 (N_30120,N_29981,N_29935);
nor U30121 (N_30121,N_29777,N_29960);
or U30122 (N_30122,N_29872,N_29791);
or U30123 (N_30123,N_29798,N_29984);
and U30124 (N_30124,N_29898,N_29931);
nor U30125 (N_30125,N_29917,N_29852);
or U30126 (N_30126,N_29907,N_29939);
or U30127 (N_30127,N_29824,N_29872);
nor U30128 (N_30128,N_29755,N_29933);
nor U30129 (N_30129,N_29994,N_29879);
and U30130 (N_30130,N_29757,N_29915);
nor U30131 (N_30131,N_29978,N_29997);
or U30132 (N_30132,N_29772,N_29768);
nand U30133 (N_30133,N_29955,N_29908);
and U30134 (N_30134,N_29767,N_29772);
xnor U30135 (N_30135,N_29838,N_29844);
nand U30136 (N_30136,N_29941,N_29847);
xor U30137 (N_30137,N_29926,N_29987);
and U30138 (N_30138,N_29805,N_29926);
or U30139 (N_30139,N_29839,N_29875);
or U30140 (N_30140,N_29991,N_29776);
or U30141 (N_30141,N_29779,N_29879);
xnor U30142 (N_30142,N_29941,N_29978);
nor U30143 (N_30143,N_29927,N_29943);
xor U30144 (N_30144,N_29792,N_29762);
nand U30145 (N_30145,N_29857,N_29845);
xnor U30146 (N_30146,N_29897,N_29787);
or U30147 (N_30147,N_29758,N_29946);
and U30148 (N_30148,N_29868,N_29839);
nor U30149 (N_30149,N_29946,N_29914);
nand U30150 (N_30150,N_29879,N_29900);
or U30151 (N_30151,N_29988,N_29906);
and U30152 (N_30152,N_29917,N_29909);
xor U30153 (N_30153,N_29812,N_29974);
and U30154 (N_30154,N_29945,N_29750);
nand U30155 (N_30155,N_29922,N_29895);
nor U30156 (N_30156,N_29990,N_29849);
or U30157 (N_30157,N_29855,N_29755);
or U30158 (N_30158,N_29840,N_29816);
nor U30159 (N_30159,N_29813,N_29899);
nor U30160 (N_30160,N_29955,N_29753);
xnor U30161 (N_30161,N_29760,N_29964);
xor U30162 (N_30162,N_29880,N_29950);
and U30163 (N_30163,N_29851,N_29811);
nand U30164 (N_30164,N_29906,N_29882);
or U30165 (N_30165,N_29864,N_29900);
xnor U30166 (N_30166,N_29776,N_29967);
and U30167 (N_30167,N_29967,N_29894);
nor U30168 (N_30168,N_29808,N_29944);
xnor U30169 (N_30169,N_29903,N_29821);
or U30170 (N_30170,N_29928,N_29877);
nor U30171 (N_30171,N_29810,N_29959);
xnor U30172 (N_30172,N_29826,N_29857);
or U30173 (N_30173,N_29905,N_29943);
nand U30174 (N_30174,N_29979,N_29939);
and U30175 (N_30175,N_29791,N_29999);
and U30176 (N_30176,N_29909,N_29859);
xor U30177 (N_30177,N_29962,N_29972);
or U30178 (N_30178,N_29933,N_29786);
nand U30179 (N_30179,N_29858,N_29855);
nand U30180 (N_30180,N_29769,N_29868);
nor U30181 (N_30181,N_29842,N_29863);
nand U30182 (N_30182,N_29821,N_29840);
and U30183 (N_30183,N_29944,N_29854);
xnor U30184 (N_30184,N_29754,N_29941);
nor U30185 (N_30185,N_29971,N_29896);
xnor U30186 (N_30186,N_29909,N_29957);
or U30187 (N_30187,N_29982,N_29932);
and U30188 (N_30188,N_29971,N_29910);
or U30189 (N_30189,N_29934,N_29857);
nand U30190 (N_30190,N_29875,N_29838);
and U30191 (N_30191,N_29886,N_29753);
nor U30192 (N_30192,N_29879,N_29856);
and U30193 (N_30193,N_29764,N_29992);
or U30194 (N_30194,N_29815,N_29764);
nor U30195 (N_30195,N_29974,N_29912);
nand U30196 (N_30196,N_29910,N_29792);
xnor U30197 (N_30197,N_29769,N_29788);
and U30198 (N_30198,N_29860,N_29886);
nand U30199 (N_30199,N_29794,N_29890);
nand U30200 (N_30200,N_29767,N_29813);
or U30201 (N_30201,N_29900,N_29849);
nand U30202 (N_30202,N_29973,N_29791);
and U30203 (N_30203,N_29862,N_29857);
nand U30204 (N_30204,N_29967,N_29813);
and U30205 (N_30205,N_29792,N_29825);
nor U30206 (N_30206,N_29843,N_29969);
xnor U30207 (N_30207,N_29972,N_29752);
or U30208 (N_30208,N_29883,N_29755);
or U30209 (N_30209,N_29776,N_29832);
nand U30210 (N_30210,N_29958,N_29970);
or U30211 (N_30211,N_29783,N_29797);
and U30212 (N_30212,N_29917,N_29898);
nand U30213 (N_30213,N_29764,N_29872);
xor U30214 (N_30214,N_29990,N_29955);
or U30215 (N_30215,N_29755,N_29999);
nor U30216 (N_30216,N_29926,N_29911);
or U30217 (N_30217,N_29921,N_29967);
nor U30218 (N_30218,N_29750,N_29839);
and U30219 (N_30219,N_29862,N_29913);
nor U30220 (N_30220,N_29910,N_29977);
nand U30221 (N_30221,N_29831,N_29824);
nor U30222 (N_30222,N_29857,N_29793);
nor U30223 (N_30223,N_29951,N_29763);
or U30224 (N_30224,N_29892,N_29848);
or U30225 (N_30225,N_29822,N_29882);
nand U30226 (N_30226,N_29884,N_29988);
or U30227 (N_30227,N_29924,N_29864);
nor U30228 (N_30228,N_29886,N_29949);
or U30229 (N_30229,N_29866,N_29955);
nand U30230 (N_30230,N_29865,N_29910);
nor U30231 (N_30231,N_29845,N_29869);
and U30232 (N_30232,N_29838,N_29984);
nor U30233 (N_30233,N_29909,N_29780);
and U30234 (N_30234,N_29926,N_29915);
xnor U30235 (N_30235,N_29862,N_29840);
nand U30236 (N_30236,N_29982,N_29885);
or U30237 (N_30237,N_29842,N_29919);
and U30238 (N_30238,N_29759,N_29904);
nand U30239 (N_30239,N_29997,N_29790);
nor U30240 (N_30240,N_29754,N_29801);
nand U30241 (N_30241,N_29862,N_29836);
or U30242 (N_30242,N_29934,N_29779);
nand U30243 (N_30243,N_29973,N_29913);
xor U30244 (N_30244,N_29905,N_29913);
and U30245 (N_30245,N_29924,N_29951);
xor U30246 (N_30246,N_29810,N_29806);
or U30247 (N_30247,N_29978,N_29841);
nand U30248 (N_30248,N_29869,N_29865);
and U30249 (N_30249,N_29832,N_29958);
and U30250 (N_30250,N_30033,N_30003);
nor U30251 (N_30251,N_30098,N_30036);
xor U30252 (N_30252,N_30212,N_30215);
nor U30253 (N_30253,N_30184,N_30174);
nand U30254 (N_30254,N_30163,N_30247);
nand U30255 (N_30255,N_30234,N_30005);
and U30256 (N_30256,N_30012,N_30238);
nor U30257 (N_30257,N_30173,N_30084);
and U30258 (N_30258,N_30006,N_30194);
and U30259 (N_30259,N_30244,N_30082);
or U30260 (N_30260,N_30227,N_30079);
and U30261 (N_30261,N_30207,N_30156);
and U30262 (N_30262,N_30027,N_30050);
nor U30263 (N_30263,N_30111,N_30106);
xor U30264 (N_30264,N_30200,N_30043);
xor U30265 (N_30265,N_30135,N_30020);
xnor U30266 (N_30266,N_30028,N_30118);
and U30267 (N_30267,N_30225,N_30228);
or U30268 (N_30268,N_30047,N_30008);
or U30269 (N_30269,N_30113,N_30166);
nand U30270 (N_30270,N_30123,N_30051);
xnor U30271 (N_30271,N_30040,N_30096);
nor U30272 (N_30272,N_30158,N_30213);
and U30273 (N_30273,N_30042,N_30103);
or U30274 (N_30274,N_30101,N_30218);
nor U30275 (N_30275,N_30066,N_30133);
xnor U30276 (N_30276,N_30094,N_30143);
nor U30277 (N_30277,N_30139,N_30085);
nor U30278 (N_30278,N_30080,N_30186);
and U30279 (N_30279,N_30162,N_30242);
nor U30280 (N_30280,N_30109,N_30171);
and U30281 (N_30281,N_30180,N_30046);
or U30282 (N_30282,N_30010,N_30142);
nand U30283 (N_30283,N_30107,N_30165);
xor U30284 (N_30284,N_30019,N_30037);
or U30285 (N_30285,N_30235,N_30120);
xor U30286 (N_30286,N_30049,N_30059);
and U30287 (N_30287,N_30181,N_30151);
and U30288 (N_30288,N_30026,N_30065);
or U30289 (N_30289,N_30229,N_30009);
nor U30290 (N_30290,N_30187,N_30104);
nor U30291 (N_30291,N_30192,N_30152);
nor U30292 (N_30292,N_30102,N_30086);
nand U30293 (N_30293,N_30100,N_30190);
xor U30294 (N_30294,N_30205,N_30141);
nor U30295 (N_30295,N_30024,N_30063);
nand U30296 (N_30296,N_30221,N_30236);
nand U30297 (N_30297,N_30130,N_30057);
nand U30298 (N_30298,N_30074,N_30149);
and U30299 (N_30299,N_30185,N_30099);
and U30300 (N_30300,N_30054,N_30230);
xor U30301 (N_30301,N_30189,N_30155);
nand U30302 (N_30302,N_30092,N_30014);
and U30303 (N_30303,N_30147,N_30126);
nand U30304 (N_30304,N_30091,N_30011);
nor U30305 (N_30305,N_30191,N_30241);
nand U30306 (N_30306,N_30125,N_30144);
nand U30307 (N_30307,N_30249,N_30214);
nor U30308 (N_30308,N_30128,N_30004);
or U30309 (N_30309,N_30088,N_30197);
and U30310 (N_30310,N_30220,N_30140);
nand U30311 (N_30311,N_30219,N_30114);
xor U30312 (N_30312,N_30129,N_30052);
or U30313 (N_30313,N_30182,N_30035);
and U30314 (N_30314,N_30039,N_30044);
nand U30315 (N_30315,N_30206,N_30062);
or U30316 (N_30316,N_30041,N_30073);
and U30317 (N_30317,N_30222,N_30031);
nand U30318 (N_30318,N_30097,N_30217);
xor U30319 (N_30319,N_30022,N_30090);
or U30320 (N_30320,N_30132,N_30061);
or U30321 (N_30321,N_30030,N_30160);
xor U30322 (N_30322,N_30150,N_30021);
and U30323 (N_30323,N_30175,N_30245);
and U30324 (N_30324,N_30154,N_30069);
and U30325 (N_30325,N_30029,N_30053);
and U30326 (N_30326,N_30131,N_30095);
nand U30327 (N_30327,N_30170,N_30193);
xor U30328 (N_30328,N_30145,N_30216);
or U30329 (N_30329,N_30122,N_30110);
nand U30330 (N_30330,N_30167,N_30164);
nand U30331 (N_30331,N_30119,N_30112);
nor U30332 (N_30332,N_30183,N_30226);
and U30333 (N_30333,N_30209,N_30071);
nand U30334 (N_30334,N_30000,N_30153);
xnor U30335 (N_30335,N_30078,N_30016);
xor U30336 (N_30336,N_30083,N_30007);
nand U30337 (N_30337,N_30199,N_30202);
or U30338 (N_30338,N_30237,N_30048);
or U30339 (N_30339,N_30081,N_30121);
xnor U30340 (N_30340,N_30178,N_30060);
nor U30341 (N_30341,N_30023,N_30105);
and U30342 (N_30342,N_30068,N_30208);
or U30343 (N_30343,N_30204,N_30127);
nor U30344 (N_30344,N_30196,N_30056);
or U30345 (N_30345,N_30075,N_30233);
xnor U30346 (N_30346,N_30002,N_30211);
and U30347 (N_30347,N_30224,N_30067);
xnor U30348 (N_30348,N_30076,N_30177);
or U30349 (N_30349,N_30070,N_30243);
xnor U30350 (N_30350,N_30115,N_30134);
nand U30351 (N_30351,N_30055,N_30117);
nand U30352 (N_30352,N_30038,N_30198);
nor U30353 (N_30353,N_30240,N_30148);
nor U30354 (N_30354,N_30116,N_30124);
xor U30355 (N_30355,N_30045,N_30032);
or U30356 (N_30356,N_30168,N_30015);
or U30357 (N_30357,N_30179,N_30064);
xor U30358 (N_30358,N_30223,N_30025);
nand U30359 (N_30359,N_30188,N_30013);
nor U30360 (N_30360,N_30093,N_30136);
nor U30361 (N_30361,N_30248,N_30077);
nand U30362 (N_30362,N_30017,N_30201);
nand U30363 (N_30363,N_30001,N_30087);
nand U30364 (N_30364,N_30108,N_30146);
nor U30365 (N_30365,N_30034,N_30172);
or U30366 (N_30366,N_30239,N_30195);
nand U30367 (N_30367,N_30137,N_30018);
nor U30368 (N_30368,N_30058,N_30161);
nand U30369 (N_30369,N_30231,N_30246);
xor U30370 (N_30370,N_30169,N_30089);
xor U30371 (N_30371,N_30210,N_30157);
xnor U30372 (N_30372,N_30232,N_30176);
or U30373 (N_30373,N_30138,N_30159);
and U30374 (N_30374,N_30072,N_30203);
and U30375 (N_30375,N_30036,N_30112);
and U30376 (N_30376,N_30083,N_30086);
or U30377 (N_30377,N_30148,N_30238);
or U30378 (N_30378,N_30130,N_30187);
xor U30379 (N_30379,N_30135,N_30238);
nand U30380 (N_30380,N_30083,N_30008);
xnor U30381 (N_30381,N_30243,N_30163);
nor U30382 (N_30382,N_30199,N_30119);
nor U30383 (N_30383,N_30237,N_30188);
or U30384 (N_30384,N_30050,N_30014);
nand U30385 (N_30385,N_30203,N_30206);
nor U30386 (N_30386,N_30146,N_30041);
nand U30387 (N_30387,N_30004,N_30092);
xor U30388 (N_30388,N_30047,N_30179);
and U30389 (N_30389,N_30185,N_30006);
and U30390 (N_30390,N_30148,N_30105);
and U30391 (N_30391,N_30112,N_30126);
xor U30392 (N_30392,N_30012,N_30045);
xnor U30393 (N_30393,N_30202,N_30161);
or U30394 (N_30394,N_30178,N_30114);
and U30395 (N_30395,N_30086,N_30204);
or U30396 (N_30396,N_30060,N_30066);
xnor U30397 (N_30397,N_30166,N_30156);
xor U30398 (N_30398,N_30128,N_30085);
xnor U30399 (N_30399,N_30102,N_30234);
and U30400 (N_30400,N_30169,N_30241);
xnor U30401 (N_30401,N_30163,N_30072);
and U30402 (N_30402,N_30084,N_30183);
and U30403 (N_30403,N_30233,N_30153);
nand U30404 (N_30404,N_30106,N_30127);
xor U30405 (N_30405,N_30194,N_30218);
and U30406 (N_30406,N_30197,N_30232);
xnor U30407 (N_30407,N_30031,N_30114);
nand U30408 (N_30408,N_30178,N_30249);
and U30409 (N_30409,N_30005,N_30221);
or U30410 (N_30410,N_30112,N_30026);
and U30411 (N_30411,N_30075,N_30232);
xor U30412 (N_30412,N_30178,N_30204);
nor U30413 (N_30413,N_30192,N_30197);
or U30414 (N_30414,N_30219,N_30185);
nor U30415 (N_30415,N_30189,N_30013);
and U30416 (N_30416,N_30142,N_30070);
or U30417 (N_30417,N_30142,N_30185);
xor U30418 (N_30418,N_30216,N_30134);
and U30419 (N_30419,N_30065,N_30053);
and U30420 (N_30420,N_30205,N_30238);
xor U30421 (N_30421,N_30191,N_30098);
xnor U30422 (N_30422,N_30177,N_30078);
or U30423 (N_30423,N_30082,N_30172);
xor U30424 (N_30424,N_30022,N_30141);
or U30425 (N_30425,N_30202,N_30060);
or U30426 (N_30426,N_30013,N_30033);
nor U30427 (N_30427,N_30000,N_30080);
xor U30428 (N_30428,N_30074,N_30082);
or U30429 (N_30429,N_30101,N_30233);
or U30430 (N_30430,N_30161,N_30131);
nand U30431 (N_30431,N_30092,N_30052);
or U30432 (N_30432,N_30079,N_30226);
nor U30433 (N_30433,N_30059,N_30030);
and U30434 (N_30434,N_30081,N_30165);
nor U30435 (N_30435,N_30173,N_30246);
nor U30436 (N_30436,N_30049,N_30010);
or U30437 (N_30437,N_30001,N_30235);
nand U30438 (N_30438,N_30216,N_30123);
and U30439 (N_30439,N_30030,N_30236);
or U30440 (N_30440,N_30174,N_30030);
and U30441 (N_30441,N_30249,N_30094);
nand U30442 (N_30442,N_30000,N_30149);
or U30443 (N_30443,N_30030,N_30233);
nand U30444 (N_30444,N_30026,N_30067);
and U30445 (N_30445,N_30011,N_30186);
nor U30446 (N_30446,N_30233,N_30126);
nand U30447 (N_30447,N_30114,N_30057);
xor U30448 (N_30448,N_30148,N_30206);
xnor U30449 (N_30449,N_30158,N_30239);
or U30450 (N_30450,N_30037,N_30073);
and U30451 (N_30451,N_30151,N_30093);
xor U30452 (N_30452,N_30071,N_30120);
nor U30453 (N_30453,N_30226,N_30187);
and U30454 (N_30454,N_30237,N_30195);
nor U30455 (N_30455,N_30105,N_30043);
and U30456 (N_30456,N_30171,N_30201);
or U30457 (N_30457,N_30144,N_30016);
or U30458 (N_30458,N_30090,N_30079);
xnor U30459 (N_30459,N_30033,N_30081);
nor U30460 (N_30460,N_30164,N_30005);
nand U30461 (N_30461,N_30093,N_30024);
xor U30462 (N_30462,N_30022,N_30002);
xor U30463 (N_30463,N_30005,N_30133);
xor U30464 (N_30464,N_30054,N_30076);
or U30465 (N_30465,N_30224,N_30115);
and U30466 (N_30466,N_30058,N_30083);
or U30467 (N_30467,N_30156,N_30136);
and U30468 (N_30468,N_30156,N_30246);
and U30469 (N_30469,N_30091,N_30214);
or U30470 (N_30470,N_30240,N_30082);
nand U30471 (N_30471,N_30216,N_30109);
nor U30472 (N_30472,N_30015,N_30085);
xor U30473 (N_30473,N_30010,N_30125);
nand U30474 (N_30474,N_30119,N_30240);
xor U30475 (N_30475,N_30151,N_30076);
and U30476 (N_30476,N_30023,N_30209);
xor U30477 (N_30477,N_30071,N_30020);
and U30478 (N_30478,N_30236,N_30011);
nand U30479 (N_30479,N_30030,N_30004);
or U30480 (N_30480,N_30116,N_30238);
nor U30481 (N_30481,N_30224,N_30099);
and U30482 (N_30482,N_30002,N_30125);
nand U30483 (N_30483,N_30205,N_30232);
and U30484 (N_30484,N_30086,N_30174);
or U30485 (N_30485,N_30143,N_30004);
or U30486 (N_30486,N_30125,N_30185);
nand U30487 (N_30487,N_30136,N_30197);
nand U30488 (N_30488,N_30205,N_30115);
xor U30489 (N_30489,N_30128,N_30105);
and U30490 (N_30490,N_30092,N_30148);
and U30491 (N_30491,N_30117,N_30192);
nor U30492 (N_30492,N_30055,N_30126);
or U30493 (N_30493,N_30016,N_30080);
xor U30494 (N_30494,N_30170,N_30185);
nand U30495 (N_30495,N_30218,N_30249);
xor U30496 (N_30496,N_30175,N_30208);
xor U30497 (N_30497,N_30068,N_30167);
nor U30498 (N_30498,N_30147,N_30246);
and U30499 (N_30499,N_30081,N_30228);
xnor U30500 (N_30500,N_30293,N_30450);
and U30501 (N_30501,N_30284,N_30277);
xnor U30502 (N_30502,N_30495,N_30404);
nand U30503 (N_30503,N_30292,N_30347);
nor U30504 (N_30504,N_30322,N_30415);
and U30505 (N_30505,N_30275,N_30412);
xor U30506 (N_30506,N_30368,N_30289);
and U30507 (N_30507,N_30385,N_30261);
xnor U30508 (N_30508,N_30474,N_30315);
or U30509 (N_30509,N_30365,N_30464);
nand U30510 (N_30510,N_30471,N_30447);
nor U30511 (N_30511,N_30324,N_30256);
xnor U30512 (N_30512,N_30250,N_30346);
and U30513 (N_30513,N_30254,N_30420);
xor U30514 (N_30514,N_30453,N_30426);
or U30515 (N_30515,N_30396,N_30440);
nand U30516 (N_30516,N_30397,N_30483);
and U30517 (N_30517,N_30298,N_30395);
or U30518 (N_30518,N_30466,N_30452);
or U30519 (N_30519,N_30458,N_30372);
nor U30520 (N_30520,N_30306,N_30391);
nand U30521 (N_30521,N_30487,N_30427);
or U30522 (N_30522,N_30352,N_30449);
and U30523 (N_30523,N_30300,N_30311);
or U30524 (N_30524,N_30473,N_30366);
or U30525 (N_30525,N_30467,N_30363);
or U30526 (N_30526,N_30373,N_30438);
nand U30527 (N_30527,N_30288,N_30394);
xor U30528 (N_30528,N_30496,N_30357);
nor U30529 (N_30529,N_30402,N_30328);
and U30530 (N_30530,N_30341,N_30305);
nor U30531 (N_30531,N_30330,N_30258);
nor U30532 (N_30532,N_30334,N_30253);
nand U30533 (N_30533,N_30418,N_30419);
nand U30534 (N_30534,N_30273,N_30424);
or U30535 (N_30535,N_30428,N_30374);
or U30536 (N_30536,N_30403,N_30409);
nor U30537 (N_30537,N_30278,N_30484);
and U30538 (N_30538,N_30345,N_30490);
nand U30539 (N_30539,N_30414,N_30367);
nor U30540 (N_30540,N_30493,N_30462);
or U30541 (N_30541,N_30475,N_30400);
or U30542 (N_30542,N_30489,N_30333);
or U30543 (N_30543,N_30349,N_30316);
and U30544 (N_30544,N_30383,N_30413);
nand U30545 (N_30545,N_30459,N_30263);
xor U30546 (N_30546,N_30405,N_30327);
or U30547 (N_30547,N_30429,N_30406);
nor U30548 (N_30548,N_30451,N_30386);
nor U30549 (N_30549,N_30304,N_30353);
and U30550 (N_30550,N_30472,N_30361);
and U30551 (N_30551,N_30314,N_30431);
nor U30552 (N_30552,N_30332,N_30390);
nand U30553 (N_30553,N_30340,N_30302);
or U30554 (N_30554,N_30494,N_30287);
xnor U30555 (N_30555,N_30369,N_30355);
and U30556 (N_30556,N_30432,N_30380);
xor U30557 (N_30557,N_30468,N_30477);
or U30558 (N_30558,N_30262,N_30437);
or U30559 (N_30559,N_30470,N_30425);
xor U30560 (N_30560,N_30433,N_30269);
nor U30561 (N_30561,N_30444,N_30266);
and U30562 (N_30562,N_30388,N_30338);
and U30563 (N_30563,N_30382,N_30356);
or U30564 (N_30564,N_30303,N_30280);
or U30565 (N_30565,N_30497,N_30279);
nand U30566 (N_30566,N_30320,N_30401);
xnor U30567 (N_30567,N_30443,N_30498);
and U30568 (N_30568,N_30499,N_30370);
xnor U30569 (N_30569,N_30271,N_30491);
nor U30570 (N_30570,N_30375,N_30312);
and U30571 (N_30571,N_30407,N_30488);
nor U30572 (N_30572,N_30364,N_30252);
or U30573 (N_30573,N_30387,N_30448);
or U30574 (N_30574,N_30268,N_30329);
xnor U30575 (N_30575,N_30348,N_30393);
xnor U30576 (N_30576,N_30339,N_30389);
xnor U30577 (N_30577,N_30301,N_30461);
nor U30578 (N_30578,N_30325,N_30486);
nor U30579 (N_30579,N_30479,N_30318);
nand U30580 (N_30580,N_30259,N_30442);
and U30581 (N_30581,N_30456,N_30326);
or U30582 (N_30582,N_30478,N_30398);
nand U30583 (N_30583,N_30321,N_30342);
nand U30584 (N_30584,N_30331,N_30480);
nand U30585 (N_30585,N_30492,N_30358);
or U30586 (N_30586,N_30481,N_30317);
nor U30587 (N_30587,N_30465,N_30354);
and U30588 (N_30588,N_30344,N_30422);
and U30589 (N_30589,N_30445,N_30323);
or U30590 (N_30590,N_30392,N_30337);
xnor U30591 (N_30591,N_30408,N_30285);
nor U30592 (N_30592,N_30399,N_30282);
xnor U30593 (N_30593,N_30309,N_30371);
nor U30594 (N_30594,N_30310,N_30291);
nor U30595 (N_30595,N_30351,N_30307);
or U30596 (N_30596,N_30454,N_30421);
xor U30597 (N_30597,N_30423,N_30411);
and U30598 (N_30598,N_30485,N_30294);
and U30599 (N_30599,N_30299,N_30286);
nor U30600 (N_30600,N_30384,N_30297);
or U30601 (N_30601,N_30381,N_30257);
nand U30602 (N_30602,N_30343,N_30296);
or U30603 (N_30603,N_30290,N_30283);
nand U30604 (N_30604,N_30295,N_30272);
nand U30605 (N_30605,N_30417,N_30378);
xnor U30606 (N_30606,N_30335,N_30276);
xnor U30607 (N_30607,N_30455,N_30350);
xor U30608 (N_30608,N_30255,N_30410);
nor U30609 (N_30609,N_30313,N_30435);
and U30610 (N_30610,N_30430,N_30360);
nand U30611 (N_30611,N_30416,N_30439);
and U30612 (N_30612,N_30308,N_30270);
nor U30613 (N_30613,N_30436,N_30251);
or U30614 (N_30614,N_30359,N_30460);
and U30615 (N_30615,N_30260,N_30264);
and U30616 (N_30616,N_30362,N_30379);
and U30617 (N_30617,N_30446,N_30265);
and U30618 (N_30618,N_30457,N_30267);
nand U30619 (N_30619,N_30377,N_30434);
xnor U30620 (N_30620,N_30441,N_30482);
or U30621 (N_30621,N_30274,N_30319);
nand U30622 (N_30622,N_30336,N_30476);
nand U30623 (N_30623,N_30463,N_30469);
and U30624 (N_30624,N_30376,N_30281);
nor U30625 (N_30625,N_30274,N_30300);
and U30626 (N_30626,N_30446,N_30415);
xnor U30627 (N_30627,N_30400,N_30392);
nor U30628 (N_30628,N_30426,N_30465);
nand U30629 (N_30629,N_30258,N_30306);
and U30630 (N_30630,N_30357,N_30421);
nand U30631 (N_30631,N_30267,N_30368);
nor U30632 (N_30632,N_30344,N_30251);
and U30633 (N_30633,N_30374,N_30323);
and U30634 (N_30634,N_30496,N_30397);
or U30635 (N_30635,N_30276,N_30479);
nor U30636 (N_30636,N_30270,N_30290);
or U30637 (N_30637,N_30468,N_30430);
and U30638 (N_30638,N_30313,N_30481);
nand U30639 (N_30639,N_30250,N_30311);
xnor U30640 (N_30640,N_30376,N_30315);
nor U30641 (N_30641,N_30285,N_30420);
xnor U30642 (N_30642,N_30299,N_30330);
nand U30643 (N_30643,N_30440,N_30354);
nor U30644 (N_30644,N_30420,N_30456);
or U30645 (N_30645,N_30433,N_30485);
nor U30646 (N_30646,N_30456,N_30375);
nor U30647 (N_30647,N_30490,N_30255);
nor U30648 (N_30648,N_30288,N_30407);
and U30649 (N_30649,N_30362,N_30469);
nor U30650 (N_30650,N_30329,N_30373);
nor U30651 (N_30651,N_30340,N_30301);
or U30652 (N_30652,N_30316,N_30250);
and U30653 (N_30653,N_30428,N_30460);
nor U30654 (N_30654,N_30290,N_30434);
or U30655 (N_30655,N_30358,N_30453);
nor U30656 (N_30656,N_30464,N_30460);
or U30657 (N_30657,N_30441,N_30314);
nand U30658 (N_30658,N_30453,N_30447);
nor U30659 (N_30659,N_30267,N_30441);
xnor U30660 (N_30660,N_30386,N_30432);
and U30661 (N_30661,N_30460,N_30472);
or U30662 (N_30662,N_30407,N_30294);
nand U30663 (N_30663,N_30357,N_30488);
and U30664 (N_30664,N_30425,N_30307);
nor U30665 (N_30665,N_30288,N_30452);
or U30666 (N_30666,N_30472,N_30451);
and U30667 (N_30667,N_30468,N_30412);
and U30668 (N_30668,N_30388,N_30350);
xnor U30669 (N_30669,N_30251,N_30276);
xnor U30670 (N_30670,N_30271,N_30376);
nand U30671 (N_30671,N_30386,N_30269);
nand U30672 (N_30672,N_30303,N_30405);
xnor U30673 (N_30673,N_30451,N_30322);
and U30674 (N_30674,N_30351,N_30478);
or U30675 (N_30675,N_30457,N_30317);
nor U30676 (N_30676,N_30427,N_30390);
or U30677 (N_30677,N_30318,N_30348);
nand U30678 (N_30678,N_30398,N_30350);
or U30679 (N_30679,N_30301,N_30439);
nand U30680 (N_30680,N_30262,N_30359);
nor U30681 (N_30681,N_30432,N_30396);
and U30682 (N_30682,N_30355,N_30444);
nand U30683 (N_30683,N_30264,N_30362);
or U30684 (N_30684,N_30451,N_30463);
nand U30685 (N_30685,N_30468,N_30446);
or U30686 (N_30686,N_30485,N_30419);
xnor U30687 (N_30687,N_30335,N_30289);
xor U30688 (N_30688,N_30461,N_30458);
or U30689 (N_30689,N_30427,N_30259);
and U30690 (N_30690,N_30342,N_30258);
xor U30691 (N_30691,N_30393,N_30487);
nand U30692 (N_30692,N_30275,N_30468);
or U30693 (N_30693,N_30412,N_30472);
nor U30694 (N_30694,N_30400,N_30370);
xor U30695 (N_30695,N_30433,N_30439);
nor U30696 (N_30696,N_30478,N_30426);
nor U30697 (N_30697,N_30333,N_30339);
xnor U30698 (N_30698,N_30443,N_30274);
and U30699 (N_30699,N_30347,N_30461);
and U30700 (N_30700,N_30335,N_30313);
nand U30701 (N_30701,N_30336,N_30316);
or U30702 (N_30702,N_30436,N_30261);
xor U30703 (N_30703,N_30336,N_30479);
nor U30704 (N_30704,N_30499,N_30405);
or U30705 (N_30705,N_30371,N_30466);
xor U30706 (N_30706,N_30408,N_30452);
and U30707 (N_30707,N_30348,N_30440);
or U30708 (N_30708,N_30279,N_30444);
and U30709 (N_30709,N_30350,N_30411);
nand U30710 (N_30710,N_30406,N_30287);
xnor U30711 (N_30711,N_30351,N_30490);
and U30712 (N_30712,N_30456,N_30381);
nand U30713 (N_30713,N_30253,N_30279);
and U30714 (N_30714,N_30356,N_30268);
xor U30715 (N_30715,N_30400,N_30256);
and U30716 (N_30716,N_30316,N_30305);
and U30717 (N_30717,N_30451,N_30371);
or U30718 (N_30718,N_30343,N_30357);
xnor U30719 (N_30719,N_30379,N_30366);
xor U30720 (N_30720,N_30456,N_30413);
nor U30721 (N_30721,N_30309,N_30324);
xor U30722 (N_30722,N_30410,N_30485);
and U30723 (N_30723,N_30346,N_30479);
and U30724 (N_30724,N_30439,N_30487);
and U30725 (N_30725,N_30270,N_30489);
and U30726 (N_30726,N_30402,N_30384);
xor U30727 (N_30727,N_30394,N_30484);
xor U30728 (N_30728,N_30368,N_30397);
or U30729 (N_30729,N_30430,N_30310);
and U30730 (N_30730,N_30397,N_30352);
or U30731 (N_30731,N_30296,N_30469);
nor U30732 (N_30732,N_30407,N_30338);
nand U30733 (N_30733,N_30352,N_30420);
and U30734 (N_30734,N_30413,N_30395);
xnor U30735 (N_30735,N_30484,N_30414);
and U30736 (N_30736,N_30466,N_30346);
and U30737 (N_30737,N_30454,N_30477);
and U30738 (N_30738,N_30441,N_30493);
nor U30739 (N_30739,N_30363,N_30346);
xnor U30740 (N_30740,N_30303,N_30370);
and U30741 (N_30741,N_30264,N_30413);
nand U30742 (N_30742,N_30346,N_30298);
xnor U30743 (N_30743,N_30263,N_30455);
xnor U30744 (N_30744,N_30453,N_30423);
xor U30745 (N_30745,N_30264,N_30456);
nor U30746 (N_30746,N_30468,N_30254);
and U30747 (N_30747,N_30457,N_30463);
xor U30748 (N_30748,N_30426,N_30268);
or U30749 (N_30749,N_30310,N_30260);
or U30750 (N_30750,N_30695,N_30660);
nand U30751 (N_30751,N_30506,N_30526);
nor U30752 (N_30752,N_30607,N_30557);
and U30753 (N_30753,N_30540,N_30724);
xor U30754 (N_30754,N_30699,N_30718);
or U30755 (N_30755,N_30543,N_30636);
nor U30756 (N_30756,N_30617,N_30597);
or U30757 (N_30757,N_30561,N_30731);
and U30758 (N_30758,N_30656,N_30568);
nand U30759 (N_30759,N_30664,N_30562);
xor U30760 (N_30760,N_30517,N_30696);
or U30761 (N_30761,N_30675,N_30666);
or U30762 (N_30762,N_30602,N_30580);
and U30763 (N_30763,N_30501,N_30592);
nor U30764 (N_30764,N_30601,N_30548);
and U30765 (N_30765,N_30616,N_30577);
and U30766 (N_30766,N_30608,N_30658);
nor U30767 (N_30767,N_30653,N_30735);
nor U30768 (N_30768,N_30502,N_30504);
and U30769 (N_30769,N_30726,N_30746);
nor U30770 (N_30770,N_30667,N_30533);
xnor U30771 (N_30771,N_30575,N_30593);
xnor U30772 (N_30772,N_30670,N_30643);
or U30773 (N_30773,N_30522,N_30662);
and U30774 (N_30774,N_30518,N_30657);
nand U30775 (N_30775,N_30694,N_30711);
nand U30776 (N_30776,N_30537,N_30564);
nor U30777 (N_30777,N_30574,N_30744);
nand U30778 (N_30778,N_30685,N_30683);
and U30779 (N_30779,N_30606,N_30513);
nand U30780 (N_30780,N_30565,N_30661);
xor U30781 (N_30781,N_30578,N_30622);
and U30782 (N_30782,N_30638,N_30573);
or U30783 (N_30783,N_30560,N_30581);
or U30784 (N_30784,N_30740,N_30702);
nor U30785 (N_30785,N_30668,N_30716);
nand U30786 (N_30786,N_30613,N_30621);
and U30787 (N_30787,N_30516,N_30717);
or U30788 (N_30788,N_30598,N_30632);
nand U30789 (N_30789,N_30505,N_30651);
xor U30790 (N_30790,N_30549,N_30633);
xnor U30791 (N_30791,N_30538,N_30539);
or U30792 (N_30792,N_30611,N_30659);
nor U30793 (N_30793,N_30665,N_30747);
or U30794 (N_30794,N_30527,N_30691);
nand U30795 (N_30795,N_30722,N_30567);
xnor U30796 (N_30796,N_30693,N_30690);
xnor U30797 (N_30797,N_30584,N_30559);
and U30798 (N_30798,N_30737,N_30637);
or U30799 (N_30799,N_30544,N_30604);
nor U30800 (N_30800,N_30646,N_30595);
or U30801 (N_30801,N_30749,N_30509);
and U30802 (N_30802,N_30671,N_30588);
xor U30803 (N_30803,N_30647,N_30710);
and U30804 (N_30804,N_30729,N_30619);
and U30805 (N_30805,N_30500,N_30555);
or U30806 (N_30806,N_30728,N_30631);
nand U30807 (N_30807,N_30566,N_30640);
and U30808 (N_30808,N_30620,N_30576);
or U30809 (N_30809,N_30725,N_30645);
nor U30810 (N_30810,N_30589,N_30705);
or U30811 (N_30811,N_30748,N_30615);
or U30812 (N_30812,N_30676,N_30635);
nand U30813 (N_30813,N_30507,N_30547);
and U30814 (N_30814,N_30678,N_30569);
nand U30815 (N_30815,N_30596,N_30612);
nor U30816 (N_30816,N_30680,N_30603);
nand U30817 (N_30817,N_30599,N_30704);
nand U30818 (N_30818,N_30706,N_30623);
nor U30819 (N_30819,N_30508,N_30503);
nand U30820 (N_30820,N_30536,N_30655);
xor U30821 (N_30821,N_30663,N_30558);
and U30822 (N_30822,N_30650,N_30551);
xor U30823 (N_30823,N_30649,N_30625);
nand U30824 (N_30824,N_30515,N_30525);
xor U30825 (N_30825,N_30514,N_30738);
and U30826 (N_30826,N_30714,N_30552);
nand U30827 (N_30827,N_30707,N_30745);
nor U30828 (N_30828,N_30733,N_30634);
and U30829 (N_30829,N_30648,N_30532);
or U30830 (N_30830,N_30644,N_30654);
xor U30831 (N_30831,N_30519,N_30730);
or U30832 (N_30832,N_30600,N_30628);
nand U30833 (N_30833,N_30629,N_30624);
nor U30834 (N_30834,N_30542,N_30523);
xnor U30835 (N_30835,N_30579,N_30719);
or U30836 (N_30836,N_30688,N_30732);
nand U30837 (N_30837,N_30689,N_30639);
xor U30838 (N_30838,N_30642,N_30563);
nand U30839 (N_30839,N_30610,N_30550);
nor U30840 (N_30840,N_30734,N_30529);
xnor U30841 (N_30841,N_30524,N_30708);
nor U30842 (N_30842,N_30677,N_30556);
or U30843 (N_30843,N_30545,N_30701);
and U30844 (N_30844,N_30553,N_30679);
and U30845 (N_30845,N_30672,N_30586);
and U30846 (N_30846,N_30521,N_30571);
nand U30847 (N_30847,N_30585,N_30652);
nor U30848 (N_30848,N_30692,N_30741);
nor U30849 (N_30849,N_30520,N_30681);
and U30850 (N_30850,N_30534,N_30712);
or U30851 (N_30851,N_30554,N_30541);
and U30852 (N_30852,N_30512,N_30669);
nor U30853 (N_30853,N_30687,N_30739);
or U30854 (N_30854,N_30510,N_30703);
or U30855 (N_30855,N_30736,N_30626);
nand U30856 (N_30856,N_30720,N_30570);
or U30857 (N_30857,N_30594,N_30535);
nand U30858 (N_30858,N_30630,N_30684);
or U30859 (N_30859,N_30727,N_30528);
nand U30860 (N_30860,N_30700,N_30618);
nor U30861 (N_30861,N_30641,N_30673);
or U30862 (N_30862,N_30583,N_30682);
nand U30863 (N_30863,N_30723,N_30713);
or U30864 (N_30864,N_30627,N_30614);
nor U30865 (N_30865,N_30546,N_30742);
nor U30866 (N_30866,N_30609,N_30697);
nand U30867 (N_30867,N_30686,N_30591);
xor U30868 (N_30868,N_30674,N_30605);
xor U30869 (N_30869,N_30721,N_30582);
nand U30870 (N_30870,N_30590,N_30511);
and U30871 (N_30871,N_30530,N_30572);
and U30872 (N_30872,N_30531,N_30698);
xor U30873 (N_30873,N_30715,N_30743);
and U30874 (N_30874,N_30587,N_30709);
xnor U30875 (N_30875,N_30603,N_30675);
nand U30876 (N_30876,N_30743,N_30505);
nand U30877 (N_30877,N_30655,N_30621);
and U30878 (N_30878,N_30580,N_30684);
xor U30879 (N_30879,N_30500,N_30726);
nand U30880 (N_30880,N_30532,N_30602);
or U30881 (N_30881,N_30516,N_30554);
or U30882 (N_30882,N_30705,N_30704);
xor U30883 (N_30883,N_30687,N_30683);
nand U30884 (N_30884,N_30692,N_30688);
and U30885 (N_30885,N_30534,N_30686);
xnor U30886 (N_30886,N_30557,N_30654);
and U30887 (N_30887,N_30658,N_30641);
xor U30888 (N_30888,N_30737,N_30697);
nor U30889 (N_30889,N_30544,N_30579);
nand U30890 (N_30890,N_30613,N_30524);
and U30891 (N_30891,N_30645,N_30524);
nor U30892 (N_30892,N_30559,N_30632);
nand U30893 (N_30893,N_30687,N_30634);
nand U30894 (N_30894,N_30641,N_30689);
nor U30895 (N_30895,N_30588,N_30595);
nand U30896 (N_30896,N_30547,N_30743);
nor U30897 (N_30897,N_30568,N_30667);
or U30898 (N_30898,N_30714,N_30743);
nor U30899 (N_30899,N_30618,N_30624);
or U30900 (N_30900,N_30714,N_30670);
nor U30901 (N_30901,N_30748,N_30737);
nor U30902 (N_30902,N_30545,N_30731);
nand U30903 (N_30903,N_30566,N_30621);
nand U30904 (N_30904,N_30674,N_30576);
or U30905 (N_30905,N_30622,N_30671);
or U30906 (N_30906,N_30715,N_30508);
xor U30907 (N_30907,N_30691,N_30597);
xor U30908 (N_30908,N_30712,N_30609);
and U30909 (N_30909,N_30581,N_30580);
nand U30910 (N_30910,N_30699,N_30581);
nor U30911 (N_30911,N_30539,N_30714);
nand U30912 (N_30912,N_30554,N_30542);
nor U30913 (N_30913,N_30598,N_30568);
and U30914 (N_30914,N_30633,N_30660);
or U30915 (N_30915,N_30630,N_30535);
nand U30916 (N_30916,N_30608,N_30724);
nand U30917 (N_30917,N_30736,N_30737);
nand U30918 (N_30918,N_30727,N_30687);
and U30919 (N_30919,N_30619,N_30588);
and U30920 (N_30920,N_30556,N_30542);
xor U30921 (N_30921,N_30702,N_30656);
xnor U30922 (N_30922,N_30684,N_30727);
nor U30923 (N_30923,N_30561,N_30717);
or U30924 (N_30924,N_30517,N_30683);
nor U30925 (N_30925,N_30669,N_30707);
xnor U30926 (N_30926,N_30605,N_30687);
xnor U30927 (N_30927,N_30530,N_30520);
or U30928 (N_30928,N_30556,N_30705);
nor U30929 (N_30929,N_30570,N_30652);
xor U30930 (N_30930,N_30625,N_30710);
nor U30931 (N_30931,N_30623,N_30644);
xnor U30932 (N_30932,N_30731,N_30599);
nor U30933 (N_30933,N_30734,N_30599);
and U30934 (N_30934,N_30517,N_30602);
and U30935 (N_30935,N_30507,N_30677);
or U30936 (N_30936,N_30691,N_30659);
nand U30937 (N_30937,N_30526,N_30675);
nor U30938 (N_30938,N_30536,N_30621);
nor U30939 (N_30939,N_30527,N_30619);
or U30940 (N_30940,N_30599,N_30623);
nand U30941 (N_30941,N_30574,N_30514);
nor U30942 (N_30942,N_30663,N_30714);
or U30943 (N_30943,N_30661,N_30532);
or U30944 (N_30944,N_30501,N_30649);
xnor U30945 (N_30945,N_30534,N_30701);
xnor U30946 (N_30946,N_30690,N_30535);
nand U30947 (N_30947,N_30592,N_30737);
nor U30948 (N_30948,N_30693,N_30660);
nor U30949 (N_30949,N_30562,N_30600);
and U30950 (N_30950,N_30665,N_30746);
xor U30951 (N_30951,N_30621,N_30732);
xnor U30952 (N_30952,N_30563,N_30730);
nand U30953 (N_30953,N_30710,N_30652);
and U30954 (N_30954,N_30597,N_30748);
or U30955 (N_30955,N_30644,N_30736);
xor U30956 (N_30956,N_30712,N_30642);
and U30957 (N_30957,N_30612,N_30585);
or U30958 (N_30958,N_30715,N_30738);
nand U30959 (N_30959,N_30594,N_30635);
xnor U30960 (N_30960,N_30536,N_30743);
nand U30961 (N_30961,N_30520,N_30748);
nor U30962 (N_30962,N_30743,N_30534);
or U30963 (N_30963,N_30561,N_30549);
or U30964 (N_30964,N_30538,N_30563);
or U30965 (N_30965,N_30620,N_30710);
nand U30966 (N_30966,N_30539,N_30549);
nor U30967 (N_30967,N_30645,N_30610);
xor U30968 (N_30968,N_30683,N_30508);
xor U30969 (N_30969,N_30627,N_30501);
nand U30970 (N_30970,N_30685,N_30613);
nand U30971 (N_30971,N_30549,N_30651);
and U30972 (N_30972,N_30681,N_30507);
nand U30973 (N_30973,N_30535,N_30598);
or U30974 (N_30974,N_30535,N_30730);
or U30975 (N_30975,N_30749,N_30731);
nand U30976 (N_30976,N_30564,N_30678);
and U30977 (N_30977,N_30626,N_30725);
xnor U30978 (N_30978,N_30588,N_30688);
nand U30979 (N_30979,N_30526,N_30620);
and U30980 (N_30980,N_30526,N_30719);
and U30981 (N_30981,N_30639,N_30582);
nand U30982 (N_30982,N_30687,N_30586);
nand U30983 (N_30983,N_30570,N_30694);
xor U30984 (N_30984,N_30654,N_30539);
nor U30985 (N_30985,N_30540,N_30593);
nand U30986 (N_30986,N_30584,N_30548);
nand U30987 (N_30987,N_30747,N_30703);
and U30988 (N_30988,N_30745,N_30720);
or U30989 (N_30989,N_30557,N_30613);
nor U30990 (N_30990,N_30626,N_30654);
and U30991 (N_30991,N_30658,N_30515);
nand U30992 (N_30992,N_30568,N_30537);
nor U30993 (N_30993,N_30673,N_30579);
nand U30994 (N_30994,N_30671,N_30545);
or U30995 (N_30995,N_30707,N_30539);
xor U30996 (N_30996,N_30644,N_30549);
nor U30997 (N_30997,N_30607,N_30572);
or U30998 (N_30998,N_30698,N_30639);
and U30999 (N_30999,N_30566,N_30712);
or U31000 (N_31000,N_30885,N_30823);
or U31001 (N_31001,N_30751,N_30766);
or U31002 (N_31002,N_30995,N_30967);
and U31003 (N_31003,N_30847,N_30866);
nor U31004 (N_31004,N_30977,N_30852);
nor U31005 (N_31005,N_30806,N_30772);
xnor U31006 (N_31006,N_30870,N_30993);
or U31007 (N_31007,N_30889,N_30824);
xnor U31008 (N_31008,N_30802,N_30902);
nand U31009 (N_31009,N_30974,N_30907);
or U31010 (N_31010,N_30799,N_30937);
xnor U31011 (N_31011,N_30776,N_30930);
and U31012 (N_31012,N_30814,N_30787);
xnor U31013 (N_31013,N_30773,N_30928);
xnor U31014 (N_31014,N_30999,N_30884);
nand U31015 (N_31015,N_30841,N_30958);
nor U31016 (N_31016,N_30803,N_30826);
or U31017 (N_31017,N_30899,N_30813);
and U31018 (N_31018,N_30756,N_30941);
nor U31019 (N_31019,N_30956,N_30834);
or U31020 (N_31020,N_30949,N_30940);
nand U31021 (N_31021,N_30777,N_30860);
and U31022 (N_31022,N_30825,N_30779);
nand U31023 (N_31023,N_30938,N_30982);
nand U31024 (N_31024,N_30838,N_30843);
or U31025 (N_31025,N_30979,N_30904);
or U31026 (N_31026,N_30819,N_30831);
nor U31027 (N_31027,N_30768,N_30973);
nor U31028 (N_31028,N_30959,N_30997);
and U31029 (N_31029,N_30877,N_30848);
nor U31030 (N_31030,N_30984,N_30871);
nor U31031 (N_31031,N_30972,N_30818);
nand U31032 (N_31032,N_30898,N_30955);
and U31033 (N_31033,N_30857,N_30908);
xnor U31034 (N_31034,N_30916,N_30906);
or U31035 (N_31035,N_30820,N_30778);
xnor U31036 (N_31036,N_30755,N_30964);
xnor U31037 (N_31037,N_30983,N_30992);
nand U31038 (N_31038,N_30939,N_30792);
nor U31039 (N_31039,N_30853,N_30986);
nand U31040 (N_31040,N_30896,N_30835);
and U31041 (N_31041,N_30788,N_30762);
nand U31042 (N_31042,N_30822,N_30905);
xor U31043 (N_31043,N_30897,N_30796);
and U31044 (N_31044,N_30855,N_30919);
nand U31045 (N_31045,N_30886,N_30975);
or U31046 (N_31046,N_30829,N_30882);
xor U31047 (N_31047,N_30863,N_30791);
nand U31048 (N_31048,N_30929,N_30892);
or U31049 (N_31049,N_30913,N_30794);
and U31050 (N_31050,N_30854,N_30931);
nor U31051 (N_31051,N_30827,N_30933);
and U31052 (N_31052,N_30921,N_30873);
xnor U31053 (N_31053,N_30785,N_30932);
nor U31054 (N_31054,N_30985,N_30774);
or U31055 (N_31055,N_30798,N_30808);
xor U31056 (N_31056,N_30900,N_30832);
and U31057 (N_31057,N_30978,N_30811);
nand U31058 (N_31058,N_30888,N_30812);
and U31059 (N_31059,N_30951,N_30804);
nand U31060 (N_31060,N_30895,N_30864);
and U31061 (N_31061,N_30954,N_30966);
or U31062 (N_31062,N_30890,N_30948);
or U31063 (N_31063,N_30833,N_30800);
nor U31064 (N_31064,N_30943,N_30935);
and U31065 (N_31065,N_30849,N_30942);
nand U31066 (N_31066,N_30927,N_30754);
xnor U31067 (N_31067,N_30781,N_30909);
or U31068 (N_31068,N_30789,N_30965);
xor U31069 (N_31069,N_30780,N_30945);
nor U31070 (N_31070,N_30887,N_30809);
nor U31071 (N_31071,N_30946,N_30915);
xnor U31072 (N_31072,N_30934,N_30752);
nand U31073 (N_31073,N_30963,N_30981);
xnor U31074 (N_31074,N_30761,N_30994);
and U31075 (N_31075,N_30891,N_30878);
nor U31076 (N_31076,N_30944,N_30759);
and U31077 (N_31077,N_30880,N_30753);
nor U31078 (N_31078,N_30969,N_30790);
nor U31079 (N_31079,N_30947,N_30875);
nand U31080 (N_31080,N_30926,N_30828);
nand U31081 (N_31081,N_30980,N_30869);
and U31082 (N_31082,N_30971,N_30910);
nor U31083 (N_31083,N_30859,N_30840);
or U31084 (N_31084,N_30837,N_30758);
or U31085 (N_31085,N_30801,N_30805);
xor U31086 (N_31086,N_30770,N_30784);
xor U31087 (N_31087,N_30861,N_30912);
or U31088 (N_31088,N_30903,N_30953);
or U31089 (N_31089,N_30830,N_30783);
xor U31090 (N_31090,N_30987,N_30816);
nand U31091 (N_31091,N_30918,N_30865);
nor U31092 (N_31092,N_30996,N_30867);
and U31093 (N_31093,N_30998,N_30782);
and U31094 (N_31094,N_30872,N_30970);
xnor U31095 (N_31095,N_30936,N_30850);
nand U31096 (N_31096,N_30901,N_30962);
or U31097 (N_31097,N_30786,N_30815);
xnor U31098 (N_31098,N_30976,N_30883);
xnor U31099 (N_31099,N_30750,N_30968);
or U31100 (N_31100,N_30844,N_30960);
nor U31101 (N_31101,N_30950,N_30924);
and U31102 (N_31102,N_30925,N_30856);
nand U31103 (N_31103,N_30845,N_30757);
xor U31104 (N_31104,N_30989,N_30876);
and U31105 (N_31105,N_30894,N_30881);
xor U31106 (N_31106,N_30807,N_30760);
nor U31107 (N_31107,N_30879,N_30769);
and U31108 (N_31108,N_30868,N_30920);
nand U31109 (N_31109,N_30771,N_30952);
or U31110 (N_31110,N_30911,N_30842);
nor U31111 (N_31111,N_30957,N_30862);
nand U31112 (N_31112,N_30764,N_30961);
nor U31113 (N_31113,N_30817,N_30991);
and U31114 (N_31114,N_30836,N_30765);
nand U31115 (N_31115,N_30810,N_30793);
nand U31116 (N_31116,N_30795,N_30917);
nor U31117 (N_31117,N_30988,N_30821);
and U31118 (N_31118,N_30839,N_30893);
and U31119 (N_31119,N_30858,N_30914);
xor U31120 (N_31120,N_30846,N_30922);
nor U31121 (N_31121,N_30797,N_30990);
or U31122 (N_31122,N_30763,N_30874);
nor U31123 (N_31123,N_30923,N_30767);
nor U31124 (N_31124,N_30775,N_30851);
or U31125 (N_31125,N_30921,N_30941);
nand U31126 (N_31126,N_30760,N_30948);
nand U31127 (N_31127,N_30820,N_30828);
and U31128 (N_31128,N_30762,N_30860);
nand U31129 (N_31129,N_30977,N_30788);
nor U31130 (N_31130,N_30872,N_30958);
and U31131 (N_31131,N_30844,N_30955);
or U31132 (N_31132,N_30954,N_30968);
nand U31133 (N_31133,N_30899,N_30990);
nor U31134 (N_31134,N_30947,N_30754);
and U31135 (N_31135,N_30873,N_30798);
or U31136 (N_31136,N_30847,N_30767);
or U31137 (N_31137,N_30974,N_30917);
or U31138 (N_31138,N_30787,N_30777);
and U31139 (N_31139,N_30805,N_30847);
nor U31140 (N_31140,N_30843,N_30891);
or U31141 (N_31141,N_30884,N_30998);
and U31142 (N_31142,N_30981,N_30914);
nor U31143 (N_31143,N_30900,N_30926);
and U31144 (N_31144,N_30852,N_30851);
or U31145 (N_31145,N_30958,N_30837);
xor U31146 (N_31146,N_30906,N_30839);
nand U31147 (N_31147,N_30817,N_30882);
or U31148 (N_31148,N_30787,N_30973);
and U31149 (N_31149,N_30912,N_30813);
nor U31150 (N_31150,N_30851,N_30979);
and U31151 (N_31151,N_30767,N_30792);
nor U31152 (N_31152,N_30986,N_30799);
nor U31153 (N_31153,N_30836,N_30992);
or U31154 (N_31154,N_30786,N_30885);
xnor U31155 (N_31155,N_30873,N_30864);
xnor U31156 (N_31156,N_30755,N_30864);
or U31157 (N_31157,N_30956,N_30960);
xor U31158 (N_31158,N_30792,N_30914);
or U31159 (N_31159,N_30815,N_30841);
nor U31160 (N_31160,N_30833,N_30784);
xnor U31161 (N_31161,N_30831,N_30846);
xnor U31162 (N_31162,N_30997,N_30872);
nand U31163 (N_31163,N_30979,N_30930);
nand U31164 (N_31164,N_30900,N_30932);
xnor U31165 (N_31165,N_30933,N_30846);
nand U31166 (N_31166,N_30938,N_30839);
nor U31167 (N_31167,N_30836,N_30999);
and U31168 (N_31168,N_30775,N_30965);
or U31169 (N_31169,N_30933,N_30879);
or U31170 (N_31170,N_30832,N_30845);
nor U31171 (N_31171,N_30958,N_30953);
xor U31172 (N_31172,N_30974,N_30756);
and U31173 (N_31173,N_30962,N_30906);
xor U31174 (N_31174,N_30785,N_30892);
or U31175 (N_31175,N_30814,N_30971);
xor U31176 (N_31176,N_30940,N_30802);
nand U31177 (N_31177,N_30929,N_30827);
or U31178 (N_31178,N_30835,N_30751);
xor U31179 (N_31179,N_30964,N_30914);
xnor U31180 (N_31180,N_30786,N_30856);
nand U31181 (N_31181,N_30959,N_30991);
and U31182 (N_31182,N_30953,N_30766);
xor U31183 (N_31183,N_30816,N_30899);
xor U31184 (N_31184,N_30777,N_30868);
nand U31185 (N_31185,N_30764,N_30979);
nand U31186 (N_31186,N_30974,N_30839);
nand U31187 (N_31187,N_30846,N_30900);
nand U31188 (N_31188,N_30978,N_30808);
and U31189 (N_31189,N_30878,N_30955);
xnor U31190 (N_31190,N_30881,N_30819);
nor U31191 (N_31191,N_30910,N_30792);
xor U31192 (N_31192,N_30981,N_30802);
nor U31193 (N_31193,N_30871,N_30857);
xnor U31194 (N_31194,N_30839,N_30957);
xnor U31195 (N_31195,N_30829,N_30944);
nand U31196 (N_31196,N_30966,N_30755);
nand U31197 (N_31197,N_30876,N_30865);
and U31198 (N_31198,N_30782,N_30935);
or U31199 (N_31199,N_30976,N_30958);
nand U31200 (N_31200,N_30884,N_30978);
nand U31201 (N_31201,N_30986,N_30850);
and U31202 (N_31202,N_30781,N_30845);
or U31203 (N_31203,N_30955,N_30947);
nand U31204 (N_31204,N_30918,N_30936);
nor U31205 (N_31205,N_30867,N_30985);
xnor U31206 (N_31206,N_30970,N_30757);
and U31207 (N_31207,N_30929,N_30856);
nor U31208 (N_31208,N_30954,N_30823);
xnor U31209 (N_31209,N_30888,N_30861);
and U31210 (N_31210,N_30835,N_30821);
nor U31211 (N_31211,N_30898,N_30786);
nor U31212 (N_31212,N_30995,N_30846);
nand U31213 (N_31213,N_30992,N_30880);
or U31214 (N_31214,N_30918,N_30816);
nor U31215 (N_31215,N_30781,N_30824);
and U31216 (N_31216,N_30806,N_30898);
nor U31217 (N_31217,N_30851,N_30815);
nor U31218 (N_31218,N_30771,N_30758);
or U31219 (N_31219,N_30757,N_30893);
or U31220 (N_31220,N_30971,N_30788);
nor U31221 (N_31221,N_30939,N_30795);
xor U31222 (N_31222,N_30904,N_30827);
nor U31223 (N_31223,N_30761,N_30755);
and U31224 (N_31224,N_30859,N_30880);
nand U31225 (N_31225,N_30786,N_30876);
and U31226 (N_31226,N_30971,N_30810);
nor U31227 (N_31227,N_30915,N_30949);
xnor U31228 (N_31228,N_30798,N_30910);
nand U31229 (N_31229,N_30793,N_30826);
nor U31230 (N_31230,N_30867,N_30966);
xnor U31231 (N_31231,N_30859,N_30792);
xor U31232 (N_31232,N_30993,N_30858);
xnor U31233 (N_31233,N_30998,N_30818);
xor U31234 (N_31234,N_30914,N_30921);
nand U31235 (N_31235,N_30937,N_30814);
xnor U31236 (N_31236,N_30840,N_30851);
or U31237 (N_31237,N_30787,N_30997);
and U31238 (N_31238,N_30871,N_30932);
and U31239 (N_31239,N_30800,N_30896);
nand U31240 (N_31240,N_30789,N_30926);
nand U31241 (N_31241,N_30949,N_30869);
nor U31242 (N_31242,N_30917,N_30966);
and U31243 (N_31243,N_30821,N_30788);
or U31244 (N_31244,N_30757,N_30991);
and U31245 (N_31245,N_30812,N_30790);
and U31246 (N_31246,N_30936,N_30964);
and U31247 (N_31247,N_30903,N_30760);
and U31248 (N_31248,N_30855,N_30885);
nand U31249 (N_31249,N_30878,N_30806);
and U31250 (N_31250,N_31122,N_31203);
xor U31251 (N_31251,N_31103,N_31009);
and U31252 (N_31252,N_31075,N_31044);
xnor U31253 (N_31253,N_31143,N_31020);
nand U31254 (N_31254,N_31029,N_31144);
nand U31255 (N_31255,N_31006,N_31025);
xor U31256 (N_31256,N_31083,N_31120);
nand U31257 (N_31257,N_31134,N_31207);
or U31258 (N_31258,N_31107,N_31224);
and U31259 (N_31259,N_31171,N_31165);
or U31260 (N_31260,N_31152,N_31186);
and U31261 (N_31261,N_31128,N_31149);
and U31262 (N_31262,N_31169,N_31185);
xnor U31263 (N_31263,N_31038,N_31012);
and U31264 (N_31264,N_31223,N_31115);
nand U31265 (N_31265,N_31225,N_31201);
nor U31266 (N_31266,N_31102,N_31013);
nand U31267 (N_31267,N_31050,N_31153);
nand U31268 (N_31268,N_31190,N_31004);
xnor U31269 (N_31269,N_31008,N_31162);
nand U31270 (N_31270,N_31125,N_31051);
xor U31271 (N_31271,N_31059,N_31123);
nor U31272 (N_31272,N_31068,N_31133);
and U31273 (N_31273,N_31121,N_31174);
and U31274 (N_31274,N_31178,N_31187);
xor U31275 (N_31275,N_31217,N_31064);
xor U31276 (N_31276,N_31236,N_31100);
nor U31277 (N_31277,N_31147,N_31140);
or U31278 (N_31278,N_31243,N_31049);
xor U31279 (N_31279,N_31196,N_31156);
or U31280 (N_31280,N_31076,N_31124);
nand U31281 (N_31281,N_31231,N_31112);
and U31282 (N_31282,N_31092,N_31234);
xor U31283 (N_31283,N_31226,N_31090);
and U31284 (N_31284,N_31109,N_31206);
and U31285 (N_31285,N_31007,N_31130);
xnor U31286 (N_31286,N_31011,N_31015);
xor U31287 (N_31287,N_31198,N_31213);
or U31288 (N_31288,N_31010,N_31105);
xnor U31289 (N_31289,N_31063,N_31175);
xnor U31290 (N_31290,N_31228,N_31245);
nor U31291 (N_31291,N_31166,N_31071);
nand U31292 (N_31292,N_31096,N_31235);
xor U31293 (N_31293,N_31084,N_31035);
or U31294 (N_31294,N_31003,N_31210);
xor U31295 (N_31295,N_31205,N_31212);
nor U31296 (N_31296,N_31157,N_31214);
or U31297 (N_31297,N_31135,N_31104);
nand U31298 (N_31298,N_31114,N_31097);
nor U31299 (N_31299,N_31229,N_31047);
xnor U31300 (N_31300,N_31057,N_31237);
or U31301 (N_31301,N_31145,N_31054);
nor U31302 (N_31302,N_31098,N_31200);
nor U31303 (N_31303,N_31118,N_31070);
nand U31304 (N_31304,N_31161,N_31242);
nor U31305 (N_31305,N_31194,N_31034);
and U31306 (N_31306,N_31085,N_31027);
or U31307 (N_31307,N_31040,N_31209);
nor U31308 (N_31308,N_31093,N_31222);
and U31309 (N_31309,N_31126,N_31017);
xor U31310 (N_31310,N_31033,N_31046);
nand U31311 (N_31311,N_31042,N_31131);
xor U31312 (N_31312,N_31148,N_31208);
nand U31313 (N_31313,N_31142,N_31014);
nand U31314 (N_31314,N_31106,N_31066);
nor U31315 (N_31315,N_31030,N_31246);
xor U31316 (N_31316,N_31036,N_31220);
xnor U31317 (N_31317,N_31219,N_31216);
or U31318 (N_31318,N_31058,N_31164);
or U31319 (N_31319,N_31177,N_31053);
nor U31320 (N_31320,N_31158,N_31155);
or U31321 (N_31321,N_31037,N_31127);
nand U31322 (N_31322,N_31211,N_31019);
nor U31323 (N_31323,N_31154,N_31141);
nand U31324 (N_31324,N_31056,N_31089);
nand U31325 (N_31325,N_31146,N_31167);
xnor U31326 (N_31326,N_31002,N_31091);
nor U31327 (N_31327,N_31111,N_31000);
and U31328 (N_31328,N_31215,N_31024);
xor U31329 (N_31329,N_31176,N_31132);
nor U31330 (N_31330,N_31168,N_31241);
or U31331 (N_31331,N_31173,N_31060);
nor U31332 (N_31332,N_31067,N_31119);
nor U31333 (N_31333,N_31077,N_31110);
and U31334 (N_31334,N_31117,N_31136);
or U31335 (N_31335,N_31137,N_31026);
nand U31336 (N_31336,N_31065,N_31184);
and U31337 (N_31337,N_31081,N_31052);
xor U31338 (N_31338,N_31192,N_31073);
xor U31339 (N_31339,N_31193,N_31016);
and U31340 (N_31340,N_31022,N_31095);
nor U31341 (N_31341,N_31218,N_31099);
and U31342 (N_31342,N_31001,N_31195);
nand U31343 (N_31343,N_31101,N_31159);
and U31344 (N_31344,N_31163,N_31202);
nand U31345 (N_31345,N_31247,N_31032);
xnor U31346 (N_31346,N_31080,N_31041);
nor U31347 (N_31347,N_31072,N_31079);
xnor U31348 (N_31348,N_31023,N_31086);
nand U31349 (N_31349,N_31069,N_31039);
or U31350 (N_31350,N_31238,N_31055);
nand U31351 (N_31351,N_31074,N_31230);
nand U31352 (N_31352,N_31151,N_31031);
xnor U31353 (N_31353,N_31018,N_31244);
or U31354 (N_31354,N_31249,N_31233);
nor U31355 (N_31355,N_31062,N_31005);
or U31356 (N_31356,N_31139,N_31172);
and U31357 (N_31357,N_31232,N_31150);
nor U31358 (N_31358,N_31191,N_31204);
nor U31359 (N_31359,N_31078,N_31181);
nand U31360 (N_31360,N_31138,N_31113);
and U31361 (N_31361,N_31028,N_31129);
xnor U31362 (N_31362,N_31248,N_31197);
nor U31363 (N_31363,N_31045,N_31088);
or U31364 (N_31364,N_31170,N_31021);
or U31365 (N_31365,N_31189,N_31082);
nor U31366 (N_31366,N_31043,N_31179);
or U31367 (N_31367,N_31094,N_31188);
nor U31368 (N_31368,N_31180,N_31108);
nor U31369 (N_31369,N_31160,N_31227);
and U31370 (N_31370,N_31199,N_31182);
nand U31371 (N_31371,N_31240,N_31061);
nand U31372 (N_31372,N_31116,N_31048);
xnor U31373 (N_31373,N_31221,N_31183);
nor U31374 (N_31374,N_31087,N_31239);
and U31375 (N_31375,N_31028,N_31215);
or U31376 (N_31376,N_31183,N_31239);
or U31377 (N_31377,N_31242,N_31102);
or U31378 (N_31378,N_31056,N_31220);
xnor U31379 (N_31379,N_31022,N_31014);
nand U31380 (N_31380,N_31059,N_31144);
nand U31381 (N_31381,N_31041,N_31181);
xnor U31382 (N_31382,N_31002,N_31034);
and U31383 (N_31383,N_31068,N_31236);
or U31384 (N_31384,N_31240,N_31082);
or U31385 (N_31385,N_31051,N_31007);
or U31386 (N_31386,N_31135,N_31180);
nand U31387 (N_31387,N_31229,N_31144);
and U31388 (N_31388,N_31218,N_31031);
and U31389 (N_31389,N_31201,N_31188);
or U31390 (N_31390,N_31114,N_31070);
nand U31391 (N_31391,N_31190,N_31193);
and U31392 (N_31392,N_31087,N_31246);
xnor U31393 (N_31393,N_31022,N_31216);
nor U31394 (N_31394,N_31057,N_31080);
xnor U31395 (N_31395,N_31113,N_31240);
or U31396 (N_31396,N_31041,N_31125);
and U31397 (N_31397,N_31185,N_31202);
nor U31398 (N_31398,N_31133,N_31007);
nand U31399 (N_31399,N_31011,N_31103);
nand U31400 (N_31400,N_31226,N_31171);
or U31401 (N_31401,N_31207,N_31061);
and U31402 (N_31402,N_31085,N_31230);
nor U31403 (N_31403,N_31049,N_31236);
nand U31404 (N_31404,N_31201,N_31117);
or U31405 (N_31405,N_31153,N_31176);
and U31406 (N_31406,N_31108,N_31126);
or U31407 (N_31407,N_31242,N_31086);
nor U31408 (N_31408,N_31009,N_31201);
or U31409 (N_31409,N_31134,N_31190);
xor U31410 (N_31410,N_31031,N_31039);
xor U31411 (N_31411,N_31052,N_31126);
and U31412 (N_31412,N_31229,N_31166);
xnor U31413 (N_31413,N_31024,N_31046);
or U31414 (N_31414,N_31053,N_31091);
and U31415 (N_31415,N_31104,N_31231);
nand U31416 (N_31416,N_31068,N_31087);
xnor U31417 (N_31417,N_31094,N_31165);
and U31418 (N_31418,N_31072,N_31018);
xor U31419 (N_31419,N_31032,N_31071);
or U31420 (N_31420,N_31060,N_31025);
nand U31421 (N_31421,N_31129,N_31078);
xnor U31422 (N_31422,N_31134,N_31009);
nand U31423 (N_31423,N_31190,N_31070);
nor U31424 (N_31424,N_31157,N_31033);
xor U31425 (N_31425,N_31231,N_31232);
and U31426 (N_31426,N_31056,N_31032);
xor U31427 (N_31427,N_31000,N_31162);
nor U31428 (N_31428,N_31000,N_31044);
or U31429 (N_31429,N_31188,N_31235);
nand U31430 (N_31430,N_31169,N_31202);
xnor U31431 (N_31431,N_31119,N_31059);
or U31432 (N_31432,N_31026,N_31191);
nor U31433 (N_31433,N_31069,N_31000);
and U31434 (N_31434,N_31047,N_31162);
nand U31435 (N_31435,N_31221,N_31025);
nor U31436 (N_31436,N_31051,N_31010);
or U31437 (N_31437,N_31149,N_31087);
or U31438 (N_31438,N_31030,N_31007);
nand U31439 (N_31439,N_31178,N_31095);
nor U31440 (N_31440,N_31002,N_31198);
nand U31441 (N_31441,N_31088,N_31023);
or U31442 (N_31442,N_31058,N_31182);
xnor U31443 (N_31443,N_31213,N_31236);
and U31444 (N_31444,N_31130,N_31195);
xor U31445 (N_31445,N_31085,N_31195);
nor U31446 (N_31446,N_31032,N_31095);
and U31447 (N_31447,N_31030,N_31210);
nand U31448 (N_31448,N_31044,N_31038);
and U31449 (N_31449,N_31147,N_31168);
xor U31450 (N_31450,N_31059,N_31033);
xor U31451 (N_31451,N_31023,N_31246);
nand U31452 (N_31452,N_31139,N_31129);
or U31453 (N_31453,N_31016,N_31154);
nand U31454 (N_31454,N_31241,N_31243);
nand U31455 (N_31455,N_31037,N_31239);
xnor U31456 (N_31456,N_31034,N_31029);
xor U31457 (N_31457,N_31118,N_31134);
or U31458 (N_31458,N_31231,N_31163);
and U31459 (N_31459,N_31033,N_31211);
and U31460 (N_31460,N_31088,N_31158);
or U31461 (N_31461,N_31054,N_31037);
or U31462 (N_31462,N_31010,N_31060);
and U31463 (N_31463,N_31168,N_31177);
or U31464 (N_31464,N_31014,N_31170);
xnor U31465 (N_31465,N_31009,N_31246);
and U31466 (N_31466,N_31005,N_31217);
nor U31467 (N_31467,N_31203,N_31002);
nand U31468 (N_31468,N_31153,N_31083);
xor U31469 (N_31469,N_31221,N_31023);
nand U31470 (N_31470,N_31120,N_31238);
or U31471 (N_31471,N_31052,N_31020);
nor U31472 (N_31472,N_31223,N_31099);
and U31473 (N_31473,N_31222,N_31201);
or U31474 (N_31474,N_31201,N_31150);
nand U31475 (N_31475,N_31112,N_31201);
xor U31476 (N_31476,N_31182,N_31085);
or U31477 (N_31477,N_31149,N_31187);
and U31478 (N_31478,N_31069,N_31092);
or U31479 (N_31479,N_31001,N_31005);
xnor U31480 (N_31480,N_31133,N_31064);
xor U31481 (N_31481,N_31120,N_31056);
or U31482 (N_31482,N_31023,N_31004);
xor U31483 (N_31483,N_31229,N_31039);
nor U31484 (N_31484,N_31158,N_31130);
or U31485 (N_31485,N_31053,N_31067);
nor U31486 (N_31486,N_31167,N_31223);
nand U31487 (N_31487,N_31025,N_31216);
xor U31488 (N_31488,N_31113,N_31195);
or U31489 (N_31489,N_31048,N_31129);
and U31490 (N_31490,N_31201,N_31191);
and U31491 (N_31491,N_31069,N_31167);
and U31492 (N_31492,N_31049,N_31247);
and U31493 (N_31493,N_31179,N_31039);
or U31494 (N_31494,N_31048,N_31218);
nor U31495 (N_31495,N_31216,N_31249);
nor U31496 (N_31496,N_31242,N_31133);
nor U31497 (N_31497,N_31165,N_31015);
and U31498 (N_31498,N_31201,N_31174);
or U31499 (N_31499,N_31145,N_31216);
or U31500 (N_31500,N_31269,N_31475);
nor U31501 (N_31501,N_31290,N_31317);
nand U31502 (N_31502,N_31486,N_31407);
xnor U31503 (N_31503,N_31494,N_31427);
xnor U31504 (N_31504,N_31313,N_31418);
and U31505 (N_31505,N_31264,N_31390);
and U31506 (N_31506,N_31280,N_31399);
nand U31507 (N_31507,N_31455,N_31309);
nand U31508 (N_31508,N_31318,N_31391);
and U31509 (N_31509,N_31428,N_31379);
and U31510 (N_31510,N_31493,N_31302);
xor U31511 (N_31511,N_31471,N_31373);
nand U31512 (N_31512,N_31378,N_31343);
or U31513 (N_31513,N_31351,N_31294);
xnor U31514 (N_31514,N_31439,N_31325);
and U31515 (N_31515,N_31276,N_31452);
and U31516 (N_31516,N_31476,N_31329);
xor U31517 (N_31517,N_31437,N_31337);
or U31518 (N_31518,N_31497,N_31487);
nand U31519 (N_31519,N_31385,N_31334);
and U31520 (N_31520,N_31319,N_31388);
and U31521 (N_31521,N_31308,N_31404);
nor U31522 (N_31522,N_31331,N_31430);
nand U31523 (N_31523,N_31441,N_31321);
nand U31524 (N_31524,N_31425,N_31456);
nand U31525 (N_31525,N_31490,N_31267);
nand U31526 (N_31526,N_31307,N_31292);
nor U31527 (N_31527,N_31466,N_31473);
or U31528 (N_31528,N_31414,N_31339);
xor U31529 (N_31529,N_31448,N_31401);
nand U31530 (N_31530,N_31374,N_31433);
xnor U31531 (N_31531,N_31410,N_31350);
nor U31532 (N_31532,N_31396,N_31324);
nand U31533 (N_31533,N_31261,N_31303);
and U31534 (N_31534,N_31316,N_31352);
nor U31535 (N_31535,N_31434,N_31345);
and U31536 (N_31536,N_31499,N_31451);
xnor U31537 (N_31537,N_31336,N_31330);
or U31538 (N_31538,N_31250,N_31484);
or U31539 (N_31539,N_31394,N_31420);
nor U31540 (N_31540,N_31299,N_31263);
or U31541 (N_31541,N_31479,N_31365);
or U31542 (N_31542,N_31323,N_31279);
nand U31543 (N_31543,N_31393,N_31477);
nor U31544 (N_31544,N_31462,N_31300);
or U31545 (N_31545,N_31492,N_31413);
xor U31546 (N_31546,N_31296,N_31354);
or U31547 (N_31547,N_31429,N_31282);
and U31548 (N_31548,N_31363,N_31253);
xnor U31549 (N_31549,N_31366,N_31277);
xor U31550 (N_31550,N_31400,N_31470);
nor U31551 (N_31551,N_31454,N_31436);
and U31552 (N_31552,N_31412,N_31335);
and U31553 (N_31553,N_31310,N_31364);
nor U31554 (N_31554,N_31328,N_31252);
xor U31555 (N_31555,N_31445,N_31417);
or U31556 (N_31556,N_31361,N_31370);
and U31557 (N_31557,N_31338,N_31332);
xnor U31558 (N_31558,N_31450,N_31457);
xor U31559 (N_31559,N_31389,N_31369);
nand U31560 (N_31560,N_31432,N_31453);
and U31561 (N_31561,N_31295,N_31371);
or U31562 (N_31562,N_31356,N_31293);
xnor U31563 (N_31563,N_31440,N_31362);
nor U31564 (N_31564,N_31483,N_31386);
nand U31565 (N_31565,N_31259,N_31358);
and U31566 (N_31566,N_31387,N_31395);
and U31567 (N_31567,N_31382,N_31273);
and U31568 (N_31568,N_31344,N_31372);
and U31569 (N_31569,N_31489,N_31415);
xnor U31570 (N_31570,N_31284,N_31392);
or U31571 (N_31571,N_31459,N_31355);
or U31572 (N_31572,N_31272,N_31341);
nor U31573 (N_31573,N_31384,N_31397);
and U31574 (N_31574,N_31262,N_31256);
and U31575 (N_31575,N_31266,N_31346);
and U31576 (N_31576,N_31260,N_31405);
or U31577 (N_31577,N_31289,N_31357);
or U31578 (N_31578,N_31291,N_31411);
xor U31579 (N_31579,N_31301,N_31314);
nor U31580 (N_31580,N_31408,N_31333);
or U31581 (N_31581,N_31375,N_31340);
nand U31582 (N_31582,N_31426,N_31422);
nor U31583 (N_31583,N_31469,N_31446);
xor U31584 (N_31584,N_31305,N_31419);
nor U31585 (N_31585,N_31353,N_31327);
nand U31586 (N_31586,N_31349,N_31480);
nand U31587 (N_31587,N_31381,N_31322);
xor U31588 (N_31588,N_31442,N_31286);
nor U31589 (N_31589,N_31270,N_31311);
nor U31590 (N_31590,N_31406,N_31464);
nand U31591 (N_31591,N_31359,N_31347);
and U31592 (N_31592,N_31431,N_31495);
nor U31593 (N_31593,N_31271,N_31447);
nor U31594 (N_31594,N_31278,N_31306);
and U31595 (N_31595,N_31403,N_31496);
xor U31596 (N_31596,N_31444,N_31255);
or U31597 (N_31597,N_31482,N_31254);
nor U31598 (N_31598,N_31265,N_31257);
xnor U31599 (N_31599,N_31380,N_31288);
nor U31600 (N_31600,N_31376,N_31467);
or U31601 (N_31601,N_31481,N_31258);
nor U31602 (N_31602,N_31463,N_31438);
xnor U31603 (N_31603,N_31298,N_31485);
or U31604 (N_31604,N_31320,N_31283);
xnor U31605 (N_31605,N_31367,N_31416);
nor U31606 (N_31606,N_31326,N_31460);
or U31607 (N_31607,N_31297,N_31423);
nand U31608 (N_31608,N_31461,N_31275);
and U31609 (N_31609,N_31474,N_31368);
xor U31610 (N_31610,N_31443,N_31398);
nand U31611 (N_31611,N_31342,N_31274);
nor U31612 (N_31612,N_31348,N_31424);
and U31613 (N_31613,N_31251,N_31287);
and U31614 (N_31614,N_31449,N_31409);
xor U31615 (N_31615,N_31488,N_31383);
nor U31616 (N_31616,N_31468,N_31285);
or U31617 (N_31617,N_31498,N_31360);
xor U31618 (N_31618,N_31472,N_31304);
nor U31619 (N_31619,N_31491,N_31421);
xor U31620 (N_31620,N_31478,N_31281);
xor U31621 (N_31621,N_31458,N_31402);
or U31622 (N_31622,N_31315,N_31312);
xnor U31623 (N_31623,N_31435,N_31377);
xnor U31624 (N_31624,N_31465,N_31268);
nand U31625 (N_31625,N_31437,N_31345);
or U31626 (N_31626,N_31440,N_31297);
nand U31627 (N_31627,N_31339,N_31426);
xnor U31628 (N_31628,N_31347,N_31370);
xnor U31629 (N_31629,N_31391,N_31435);
and U31630 (N_31630,N_31350,N_31341);
or U31631 (N_31631,N_31313,N_31349);
nor U31632 (N_31632,N_31300,N_31415);
nor U31633 (N_31633,N_31463,N_31497);
nor U31634 (N_31634,N_31293,N_31435);
nor U31635 (N_31635,N_31320,N_31354);
or U31636 (N_31636,N_31359,N_31486);
and U31637 (N_31637,N_31378,N_31465);
or U31638 (N_31638,N_31287,N_31270);
and U31639 (N_31639,N_31250,N_31337);
and U31640 (N_31640,N_31366,N_31269);
nand U31641 (N_31641,N_31358,N_31436);
and U31642 (N_31642,N_31474,N_31383);
and U31643 (N_31643,N_31489,N_31375);
nand U31644 (N_31644,N_31396,N_31394);
or U31645 (N_31645,N_31322,N_31431);
or U31646 (N_31646,N_31395,N_31263);
and U31647 (N_31647,N_31330,N_31325);
xor U31648 (N_31648,N_31420,N_31288);
nand U31649 (N_31649,N_31384,N_31411);
nor U31650 (N_31650,N_31366,N_31330);
and U31651 (N_31651,N_31406,N_31293);
or U31652 (N_31652,N_31312,N_31272);
nand U31653 (N_31653,N_31443,N_31454);
xor U31654 (N_31654,N_31359,N_31378);
xor U31655 (N_31655,N_31326,N_31381);
xnor U31656 (N_31656,N_31429,N_31287);
nand U31657 (N_31657,N_31349,N_31434);
or U31658 (N_31658,N_31385,N_31474);
and U31659 (N_31659,N_31480,N_31371);
nand U31660 (N_31660,N_31473,N_31268);
and U31661 (N_31661,N_31492,N_31325);
and U31662 (N_31662,N_31384,N_31429);
xnor U31663 (N_31663,N_31295,N_31459);
or U31664 (N_31664,N_31462,N_31484);
nand U31665 (N_31665,N_31490,N_31348);
nand U31666 (N_31666,N_31353,N_31385);
and U31667 (N_31667,N_31450,N_31430);
or U31668 (N_31668,N_31489,N_31354);
nand U31669 (N_31669,N_31349,N_31323);
nand U31670 (N_31670,N_31255,N_31279);
xnor U31671 (N_31671,N_31454,N_31309);
nand U31672 (N_31672,N_31373,N_31412);
nand U31673 (N_31673,N_31383,N_31496);
xnor U31674 (N_31674,N_31418,N_31255);
xnor U31675 (N_31675,N_31452,N_31375);
and U31676 (N_31676,N_31293,N_31307);
nand U31677 (N_31677,N_31292,N_31328);
nor U31678 (N_31678,N_31294,N_31378);
or U31679 (N_31679,N_31292,N_31351);
or U31680 (N_31680,N_31445,N_31358);
and U31681 (N_31681,N_31410,N_31417);
or U31682 (N_31682,N_31339,N_31460);
nand U31683 (N_31683,N_31368,N_31402);
and U31684 (N_31684,N_31330,N_31482);
xnor U31685 (N_31685,N_31469,N_31287);
nor U31686 (N_31686,N_31442,N_31465);
nand U31687 (N_31687,N_31383,N_31319);
nor U31688 (N_31688,N_31400,N_31338);
nand U31689 (N_31689,N_31392,N_31477);
nand U31690 (N_31690,N_31288,N_31411);
and U31691 (N_31691,N_31392,N_31340);
or U31692 (N_31692,N_31491,N_31496);
nor U31693 (N_31693,N_31427,N_31364);
nor U31694 (N_31694,N_31433,N_31301);
and U31695 (N_31695,N_31290,N_31402);
nor U31696 (N_31696,N_31323,N_31359);
or U31697 (N_31697,N_31470,N_31409);
and U31698 (N_31698,N_31430,N_31309);
nor U31699 (N_31699,N_31341,N_31320);
or U31700 (N_31700,N_31480,N_31440);
nand U31701 (N_31701,N_31338,N_31377);
xnor U31702 (N_31702,N_31308,N_31337);
xnor U31703 (N_31703,N_31313,N_31425);
or U31704 (N_31704,N_31348,N_31353);
xnor U31705 (N_31705,N_31485,N_31494);
nand U31706 (N_31706,N_31385,N_31279);
nor U31707 (N_31707,N_31346,N_31321);
nand U31708 (N_31708,N_31262,N_31409);
nand U31709 (N_31709,N_31337,N_31471);
or U31710 (N_31710,N_31411,N_31383);
or U31711 (N_31711,N_31330,N_31353);
nor U31712 (N_31712,N_31356,N_31252);
xor U31713 (N_31713,N_31323,N_31302);
nor U31714 (N_31714,N_31499,N_31378);
nand U31715 (N_31715,N_31306,N_31300);
or U31716 (N_31716,N_31377,N_31493);
or U31717 (N_31717,N_31317,N_31282);
or U31718 (N_31718,N_31301,N_31396);
and U31719 (N_31719,N_31496,N_31382);
nand U31720 (N_31720,N_31280,N_31381);
nor U31721 (N_31721,N_31289,N_31419);
nor U31722 (N_31722,N_31370,N_31425);
and U31723 (N_31723,N_31351,N_31302);
nand U31724 (N_31724,N_31445,N_31292);
or U31725 (N_31725,N_31403,N_31392);
nand U31726 (N_31726,N_31359,N_31357);
nor U31727 (N_31727,N_31388,N_31430);
nor U31728 (N_31728,N_31463,N_31267);
nand U31729 (N_31729,N_31373,N_31469);
xor U31730 (N_31730,N_31345,N_31499);
or U31731 (N_31731,N_31393,N_31495);
and U31732 (N_31732,N_31401,N_31403);
or U31733 (N_31733,N_31408,N_31358);
and U31734 (N_31734,N_31287,N_31488);
xor U31735 (N_31735,N_31466,N_31342);
xor U31736 (N_31736,N_31390,N_31326);
and U31737 (N_31737,N_31304,N_31277);
nand U31738 (N_31738,N_31372,N_31474);
nand U31739 (N_31739,N_31489,N_31358);
nor U31740 (N_31740,N_31372,N_31382);
nor U31741 (N_31741,N_31457,N_31336);
xor U31742 (N_31742,N_31308,N_31422);
nor U31743 (N_31743,N_31253,N_31409);
xor U31744 (N_31744,N_31369,N_31326);
xor U31745 (N_31745,N_31263,N_31297);
nand U31746 (N_31746,N_31460,N_31432);
xor U31747 (N_31747,N_31329,N_31463);
xor U31748 (N_31748,N_31476,N_31260);
nand U31749 (N_31749,N_31265,N_31458);
nor U31750 (N_31750,N_31567,N_31617);
and U31751 (N_31751,N_31651,N_31687);
nor U31752 (N_31752,N_31717,N_31581);
or U31753 (N_31753,N_31749,N_31718);
and U31754 (N_31754,N_31643,N_31723);
and U31755 (N_31755,N_31621,N_31601);
xnor U31756 (N_31756,N_31678,N_31665);
nor U31757 (N_31757,N_31624,N_31611);
or U31758 (N_31758,N_31696,N_31725);
nor U31759 (N_31759,N_31571,N_31721);
and U31760 (N_31760,N_31736,N_31686);
nor U31761 (N_31761,N_31518,N_31582);
nor U31762 (N_31762,N_31684,N_31610);
or U31763 (N_31763,N_31585,N_31535);
and U31764 (N_31764,N_31530,N_31598);
and U31765 (N_31765,N_31555,N_31644);
or U31766 (N_31766,N_31680,N_31603);
nor U31767 (N_31767,N_31536,N_31501);
and U31768 (N_31768,N_31633,N_31515);
and U31769 (N_31769,N_31682,N_31600);
or U31770 (N_31770,N_31742,N_31513);
xnor U31771 (N_31771,N_31589,N_31511);
or U31772 (N_31772,N_31538,N_31689);
and U31773 (N_31773,N_31658,N_31645);
and U31774 (N_31774,N_31584,N_31668);
nor U31775 (N_31775,N_31550,N_31710);
nor U31776 (N_31776,N_31639,N_31500);
nand U31777 (N_31777,N_31542,N_31634);
nand U31778 (N_31778,N_31619,N_31580);
nor U31779 (N_31779,N_31572,N_31745);
xnor U31780 (N_31780,N_31510,N_31508);
xor U31781 (N_31781,N_31588,N_31591);
and U31782 (N_31782,N_31529,N_31618);
and U31783 (N_31783,N_31656,N_31583);
nand U31784 (N_31784,N_31666,N_31597);
xor U31785 (N_31785,N_31740,N_31677);
xor U31786 (N_31786,N_31626,N_31671);
nor U31787 (N_31787,N_31704,N_31635);
or U31788 (N_31788,N_31661,N_31596);
nor U31789 (N_31789,N_31594,N_31657);
nor U31790 (N_31790,N_31659,N_31506);
and U31791 (N_31791,N_31568,N_31629);
nor U31792 (N_31792,N_31539,N_31612);
nand U31793 (N_31793,N_31531,N_31632);
or U31794 (N_31794,N_31625,N_31565);
or U31795 (N_31795,N_31509,N_31650);
or U31796 (N_31796,N_31517,N_31747);
and U31797 (N_31797,N_31700,N_31524);
xnor U31798 (N_31798,N_31560,N_31637);
xnor U31799 (N_31799,N_31595,N_31613);
xnor U31800 (N_31800,N_31602,N_31738);
xnor U31801 (N_31801,N_31520,N_31732);
and U31802 (N_31802,N_31512,N_31711);
xnor U31803 (N_31803,N_31514,N_31590);
and U31804 (N_31804,N_31566,N_31712);
or U31805 (N_31805,N_31559,N_31607);
xor U31806 (N_31806,N_31586,N_31553);
nor U31807 (N_31807,N_31574,N_31527);
or U31808 (N_31808,N_31516,N_31748);
nor U31809 (N_31809,N_31642,N_31675);
xnor U31810 (N_31810,N_31739,N_31690);
or U31811 (N_31811,N_31576,N_31698);
nand U31812 (N_31812,N_31622,N_31699);
xor U31813 (N_31813,N_31681,N_31627);
nor U31814 (N_31814,N_31557,N_31662);
xnor U31815 (N_31815,N_31703,N_31743);
nand U31816 (N_31816,N_31693,N_31620);
and U31817 (N_31817,N_31664,N_31521);
nor U31818 (N_31818,N_31691,N_31606);
and U31819 (N_31819,N_31551,N_31545);
xnor U31820 (N_31820,N_31528,N_31706);
and U31821 (N_31821,N_31556,N_31578);
and U31822 (N_31822,N_31573,N_31720);
nor U31823 (N_31823,N_31523,N_31663);
nor U31824 (N_31824,N_31705,N_31562);
nor U31825 (N_31825,N_31605,N_31672);
or U31826 (N_31826,N_31541,N_31652);
nor U31827 (N_31827,N_31615,N_31604);
nand U31828 (N_31828,N_31667,N_31579);
nor U31829 (N_31829,N_31729,N_31636);
nor U31830 (N_31830,N_31653,N_31697);
and U31831 (N_31831,N_31676,N_31537);
and U31832 (N_31832,N_31505,N_31549);
nand U31833 (N_31833,N_31592,N_31731);
and U31834 (N_31834,N_31519,N_31587);
nor U31835 (N_31835,N_31713,N_31546);
xor U31836 (N_31836,N_31575,N_31730);
nor U31837 (N_31837,N_31654,N_31599);
nor U31838 (N_31838,N_31694,N_31544);
nor U31839 (N_31839,N_31669,N_31688);
xnor U31840 (N_31840,N_31641,N_31623);
xnor U31841 (N_31841,N_31532,N_31734);
xnor U31842 (N_31842,N_31577,N_31640);
and U31843 (N_31843,N_31695,N_31504);
nand U31844 (N_31844,N_31503,N_31707);
nor U31845 (N_31845,N_31719,N_31628);
nand U31846 (N_31846,N_31507,N_31737);
nor U31847 (N_31847,N_31522,N_31655);
and U31848 (N_31848,N_31569,N_31540);
and U31849 (N_31849,N_31552,N_31570);
nand U31850 (N_31850,N_31631,N_31733);
nand U31851 (N_31851,N_31670,N_31608);
xnor U31852 (N_31852,N_31616,N_31674);
and U31853 (N_31853,N_31744,N_31741);
xor U31854 (N_31854,N_31722,N_31548);
and U31855 (N_31855,N_31746,N_31716);
or U31856 (N_31856,N_31502,N_31563);
nand U31857 (N_31857,N_31673,N_31525);
nand U31858 (N_31858,N_31593,N_31683);
or U31859 (N_31859,N_31724,N_31649);
nand U31860 (N_31860,N_31679,N_31708);
nand U31861 (N_31861,N_31564,N_31709);
and U31862 (N_31862,N_31726,N_31533);
or U31863 (N_31863,N_31554,N_31702);
and U31864 (N_31864,N_31547,N_31543);
xor U31865 (N_31865,N_31701,N_31660);
nand U31866 (N_31866,N_31714,N_31526);
xor U31867 (N_31867,N_31630,N_31638);
or U31868 (N_31868,N_31561,N_31727);
nand U31869 (N_31869,N_31735,N_31614);
or U31870 (N_31870,N_31685,N_31728);
nand U31871 (N_31871,N_31648,N_31715);
nor U31872 (N_31872,N_31558,N_31646);
xnor U31873 (N_31873,N_31647,N_31534);
xor U31874 (N_31874,N_31609,N_31692);
nand U31875 (N_31875,N_31694,N_31554);
or U31876 (N_31876,N_31673,N_31633);
xnor U31877 (N_31877,N_31741,N_31635);
or U31878 (N_31878,N_31679,N_31666);
xor U31879 (N_31879,N_31521,N_31675);
xor U31880 (N_31880,N_31620,N_31653);
xor U31881 (N_31881,N_31720,N_31701);
nor U31882 (N_31882,N_31547,N_31579);
nor U31883 (N_31883,N_31583,N_31652);
nand U31884 (N_31884,N_31519,N_31561);
and U31885 (N_31885,N_31706,N_31733);
and U31886 (N_31886,N_31694,N_31550);
nand U31887 (N_31887,N_31688,N_31652);
or U31888 (N_31888,N_31621,N_31614);
nor U31889 (N_31889,N_31681,N_31674);
and U31890 (N_31890,N_31636,N_31674);
nand U31891 (N_31891,N_31688,N_31606);
or U31892 (N_31892,N_31728,N_31530);
and U31893 (N_31893,N_31591,N_31717);
or U31894 (N_31894,N_31603,N_31515);
xor U31895 (N_31895,N_31572,N_31581);
or U31896 (N_31896,N_31666,N_31658);
nor U31897 (N_31897,N_31657,N_31534);
nor U31898 (N_31898,N_31721,N_31627);
nor U31899 (N_31899,N_31712,N_31622);
nor U31900 (N_31900,N_31677,N_31587);
xor U31901 (N_31901,N_31560,N_31513);
xor U31902 (N_31902,N_31501,N_31745);
nor U31903 (N_31903,N_31641,N_31602);
xor U31904 (N_31904,N_31536,N_31722);
nor U31905 (N_31905,N_31586,N_31639);
nor U31906 (N_31906,N_31536,N_31568);
nand U31907 (N_31907,N_31693,N_31559);
and U31908 (N_31908,N_31609,N_31631);
xor U31909 (N_31909,N_31731,N_31610);
nor U31910 (N_31910,N_31532,N_31630);
or U31911 (N_31911,N_31679,N_31638);
nand U31912 (N_31912,N_31589,N_31729);
and U31913 (N_31913,N_31733,N_31721);
or U31914 (N_31914,N_31671,N_31555);
or U31915 (N_31915,N_31694,N_31696);
nor U31916 (N_31916,N_31682,N_31510);
and U31917 (N_31917,N_31581,N_31694);
nor U31918 (N_31918,N_31505,N_31558);
and U31919 (N_31919,N_31650,N_31501);
and U31920 (N_31920,N_31707,N_31560);
nor U31921 (N_31921,N_31502,N_31661);
nor U31922 (N_31922,N_31664,N_31652);
xor U31923 (N_31923,N_31521,N_31509);
or U31924 (N_31924,N_31677,N_31645);
xnor U31925 (N_31925,N_31510,N_31524);
xnor U31926 (N_31926,N_31524,N_31706);
and U31927 (N_31927,N_31626,N_31686);
nand U31928 (N_31928,N_31700,N_31589);
and U31929 (N_31929,N_31599,N_31732);
xor U31930 (N_31930,N_31617,N_31552);
nand U31931 (N_31931,N_31673,N_31694);
nor U31932 (N_31932,N_31571,N_31524);
or U31933 (N_31933,N_31541,N_31740);
xor U31934 (N_31934,N_31712,N_31679);
and U31935 (N_31935,N_31524,N_31593);
or U31936 (N_31936,N_31658,N_31577);
or U31937 (N_31937,N_31733,N_31699);
nand U31938 (N_31938,N_31646,N_31599);
and U31939 (N_31939,N_31588,N_31552);
or U31940 (N_31940,N_31518,N_31501);
or U31941 (N_31941,N_31547,N_31677);
and U31942 (N_31942,N_31595,N_31662);
and U31943 (N_31943,N_31613,N_31681);
or U31944 (N_31944,N_31669,N_31604);
xnor U31945 (N_31945,N_31708,N_31594);
or U31946 (N_31946,N_31538,N_31583);
or U31947 (N_31947,N_31550,N_31662);
nor U31948 (N_31948,N_31523,N_31608);
xnor U31949 (N_31949,N_31630,N_31644);
or U31950 (N_31950,N_31500,N_31535);
nand U31951 (N_31951,N_31573,N_31551);
nor U31952 (N_31952,N_31537,N_31636);
xor U31953 (N_31953,N_31597,N_31611);
and U31954 (N_31954,N_31601,N_31548);
or U31955 (N_31955,N_31717,N_31691);
nand U31956 (N_31956,N_31614,N_31559);
nor U31957 (N_31957,N_31526,N_31556);
nor U31958 (N_31958,N_31738,N_31633);
and U31959 (N_31959,N_31689,N_31525);
or U31960 (N_31960,N_31566,N_31691);
nand U31961 (N_31961,N_31708,N_31619);
nand U31962 (N_31962,N_31561,N_31655);
nor U31963 (N_31963,N_31612,N_31619);
and U31964 (N_31964,N_31696,N_31699);
xnor U31965 (N_31965,N_31709,N_31721);
or U31966 (N_31966,N_31577,N_31632);
nand U31967 (N_31967,N_31635,N_31674);
xor U31968 (N_31968,N_31587,N_31513);
nor U31969 (N_31969,N_31658,N_31552);
nor U31970 (N_31970,N_31561,N_31740);
nor U31971 (N_31971,N_31566,N_31551);
xnor U31972 (N_31972,N_31675,N_31628);
or U31973 (N_31973,N_31555,N_31550);
xor U31974 (N_31974,N_31659,N_31589);
or U31975 (N_31975,N_31546,N_31726);
and U31976 (N_31976,N_31613,N_31635);
and U31977 (N_31977,N_31594,N_31696);
xnor U31978 (N_31978,N_31718,N_31502);
nor U31979 (N_31979,N_31675,N_31727);
nand U31980 (N_31980,N_31615,N_31505);
nor U31981 (N_31981,N_31604,N_31598);
nand U31982 (N_31982,N_31554,N_31599);
nand U31983 (N_31983,N_31612,N_31731);
xor U31984 (N_31984,N_31517,N_31597);
xor U31985 (N_31985,N_31644,N_31661);
or U31986 (N_31986,N_31674,N_31699);
or U31987 (N_31987,N_31637,N_31690);
xor U31988 (N_31988,N_31649,N_31546);
nor U31989 (N_31989,N_31567,N_31561);
or U31990 (N_31990,N_31536,N_31642);
nor U31991 (N_31991,N_31733,N_31679);
xor U31992 (N_31992,N_31712,N_31591);
or U31993 (N_31993,N_31552,N_31576);
nor U31994 (N_31994,N_31745,N_31718);
and U31995 (N_31995,N_31719,N_31613);
nand U31996 (N_31996,N_31610,N_31518);
nand U31997 (N_31997,N_31746,N_31551);
or U31998 (N_31998,N_31514,N_31652);
nand U31999 (N_31999,N_31590,N_31700);
nor U32000 (N_32000,N_31814,N_31949);
nor U32001 (N_32001,N_31756,N_31805);
nand U32002 (N_32002,N_31889,N_31755);
nand U32003 (N_32003,N_31882,N_31914);
and U32004 (N_32004,N_31987,N_31894);
nor U32005 (N_32005,N_31907,N_31820);
xnor U32006 (N_32006,N_31818,N_31846);
and U32007 (N_32007,N_31992,N_31845);
nand U32008 (N_32008,N_31969,N_31993);
xnor U32009 (N_32009,N_31765,N_31997);
nand U32010 (N_32010,N_31826,N_31788);
or U32011 (N_32011,N_31841,N_31859);
and U32012 (N_32012,N_31954,N_31804);
xnor U32013 (N_32013,N_31860,N_31924);
xnor U32014 (N_32014,N_31848,N_31878);
xor U32015 (N_32015,N_31861,N_31800);
xnor U32016 (N_32016,N_31831,N_31994);
and U32017 (N_32017,N_31785,N_31783);
nand U32018 (N_32018,N_31919,N_31928);
nor U32019 (N_32019,N_31975,N_31821);
nand U32020 (N_32020,N_31927,N_31921);
nor U32021 (N_32021,N_31854,N_31835);
or U32022 (N_32022,N_31798,N_31869);
and U32023 (N_32023,N_31867,N_31839);
or U32024 (N_32024,N_31998,N_31908);
xor U32025 (N_32025,N_31901,N_31829);
and U32026 (N_32026,N_31779,N_31970);
and U32027 (N_32027,N_31881,N_31767);
and U32028 (N_32028,N_31912,N_31776);
xnor U32029 (N_32029,N_31838,N_31811);
and U32030 (N_32030,N_31792,N_31855);
or U32031 (N_32031,N_31906,N_31795);
nor U32032 (N_32032,N_31934,N_31898);
nand U32033 (N_32033,N_31982,N_31833);
or U32034 (N_32034,N_31762,N_31989);
xor U32035 (N_32035,N_31948,N_31752);
or U32036 (N_32036,N_31922,N_31813);
xor U32037 (N_32037,N_31761,N_31942);
and U32038 (N_32038,N_31957,N_31790);
or U32039 (N_32039,N_31893,N_31817);
nand U32040 (N_32040,N_31771,N_31777);
or U32041 (N_32041,N_31849,N_31976);
xnor U32042 (N_32042,N_31923,N_31754);
nand U32043 (N_32043,N_31981,N_31900);
nand U32044 (N_32044,N_31773,N_31874);
nand U32045 (N_32045,N_31902,N_31772);
or U32046 (N_32046,N_31910,N_31809);
nand U32047 (N_32047,N_31815,N_31905);
and U32048 (N_32048,N_31953,N_31827);
and U32049 (N_32049,N_31796,N_31963);
or U32050 (N_32050,N_31886,N_31778);
or U32051 (N_32051,N_31959,N_31842);
or U32052 (N_32052,N_31844,N_31918);
or U32053 (N_32053,N_31995,N_31939);
xor U32054 (N_32054,N_31864,N_31808);
or U32055 (N_32055,N_31896,N_31757);
xnor U32056 (N_32056,N_31965,N_31787);
xor U32057 (N_32057,N_31973,N_31843);
xor U32058 (N_32058,N_31875,N_31780);
or U32059 (N_32059,N_31759,N_31840);
and U32060 (N_32060,N_31943,N_31760);
and U32061 (N_32061,N_31911,N_31824);
or U32062 (N_32062,N_31819,N_31823);
nor U32063 (N_32063,N_31852,N_31916);
or U32064 (N_32064,N_31950,N_31917);
nor U32065 (N_32065,N_31784,N_31979);
nand U32066 (N_32066,N_31863,N_31937);
nand U32067 (N_32067,N_31877,N_31847);
or U32068 (N_32068,N_31816,N_31974);
nor U32069 (N_32069,N_31883,N_31884);
xnor U32070 (N_32070,N_31888,N_31850);
and U32071 (N_32071,N_31946,N_31880);
xor U32072 (N_32072,N_31944,N_31920);
nand U32073 (N_32073,N_31865,N_31885);
nand U32074 (N_32074,N_31853,N_31764);
and U32075 (N_32075,N_31909,N_31897);
or U32076 (N_32076,N_31988,N_31890);
and U32077 (N_32077,N_31806,N_31830);
nand U32078 (N_32078,N_31951,N_31887);
or U32079 (N_32079,N_31892,N_31828);
nand U32080 (N_32080,N_31899,N_31807);
or U32081 (N_32081,N_31810,N_31904);
xor U32082 (N_32082,N_31933,N_31936);
or U32083 (N_32083,N_31856,N_31832);
and U32084 (N_32084,N_31915,N_31945);
nand U32085 (N_32085,N_31967,N_31774);
nor U32086 (N_32086,N_31868,N_31930);
nand U32087 (N_32087,N_31985,N_31822);
or U32088 (N_32088,N_31990,N_31781);
nand U32089 (N_32089,N_31931,N_31782);
nor U32090 (N_32090,N_31879,N_31960);
nand U32091 (N_32091,N_31895,N_31977);
nand U32092 (N_32092,N_31966,N_31968);
or U32093 (N_32093,N_31870,N_31753);
xor U32094 (N_32094,N_31961,N_31789);
nor U32095 (N_32095,N_31851,N_31812);
nor U32096 (N_32096,N_31956,N_31866);
and U32097 (N_32097,N_31962,N_31872);
nor U32098 (N_32098,N_31964,N_31834);
xor U32099 (N_32099,N_31802,N_31972);
and U32100 (N_32100,N_31769,N_31941);
or U32101 (N_32101,N_31986,N_31825);
xor U32102 (N_32102,N_31797,N_31903);
nor U32103 (N_32103,N_31768,N_31958);
and U32104 (N_32104,N_31871,N_31955);
xor U32105 (N_32105,N_31758,N_31793);
and U32106 (N_32106,N_31926,N_31836);
nand U32107 (N_32107,N_31873,N_31837);
and U32108 (N_32108,N_31940,N_31803);
xnor U32109 (N_32109,N_31862,N_31876);
nand U32110 (N_32110,N_31786,N_31766);
nor U32111 (N_32111,N_31983,N_31858);
or U32112 (N_32112,N_31999,N_31938);
xnor U32113 (N_32113,N_31935,N_31984);
xnor U32114 (N_32114,N_31991,N_31952);
xor U32115 (N_32115,N_31947,N_31857);
xnor U32116 (N_32116,N_31971,N_31799);
or U32117 (N_32117,N_31794,N_31913);
or U32118 (N_32118,N_31932,N_31770);
xnor U32119 (N_32119,N_31763,N_31980);
nand U32120 (N_32120,N_31978,N_31891);
nand U32121 (N_32121,N_31996,N_31925);
xor U32122 (N_32122,N_31791,N_31929);
xor U32123 (N_32123,N_31750,N_31801);
nand U32124 (N_32124,N_31751,N_31775);
xor U32125 (N_32125,N_31856,N_31802);
nor U32126 (N_32126,N_31778,N_31779);
xnor U32127 (N_32127,N_31939,N_31988);
nand U32128 (N_32128,N_31887,N_31764);
nor U32129 (N_32129,N_31884,N_31876);
nand U32130 (N_32130,N_31753,N_31897);
nand U32131 (N_32131,N_31978,N_31781);
nand U32132 (N_32132,N_31935,N_31793);
nor U32133 (N_32133,N_31772,N_31929);
and U32134 (N_32134,N_31769,N_31952);
nor U32135 (N_32135,N_31811,N_31876);
nor U32136 (N_32136,N_31841,N_31761);
nand U32137 (N_32137,N_31915,N_31968);
xnor U32138 (N_32138,N_31978,N_31964);
and U32139 (N_32139,N_31841,N_31981);
xnor U32140 (N_32140,N_31826,N_31793);
or U32141 (N_32141,N_31855,N_31933);
nor U32142 (N_32142,N_31889,N_31761);
and U32143 (N_32143,N_31868,N_31864);
nor U32144 (N_32144,N_31795,N_31982);
and U32145 (N_32145,N_31956,N_31981);
and U32146 (N_32146,N_31905,N_31837);
nor U32147 (N_32147,N_31786,N_31819);
or U32148 (N_32148,N_31810,N_31798);
and U32149 (N_32149,N_31827,N_31967);
nand U32150 (N_32150,N_31914,N_31834);
xnor U32151 (N_32151,N_31787,N_31792);
nand U32152 (N_32152,N_31983,N_31770);
xor U32153 (N_32153,N_31892,N_31836);
and U32154 (N_32154,N_31906,N_31977);
or U32155 (N_32155,N_31954,N_31971);
nor U32156 (N_32156,N_31913,N_31848);
nand U32157 (N_32157,N_31813,N_31852);
or U32158 (N_32158,N_31805,N_31885);
nand U32159 (N_32159,N_31919,N_31915);
nor U32160 (N_32160,N_31960,N_31781);
and U32161 (N_32161,N_31937,N_31878);
nor U32162 (N_32162,N_31829,N_31824);
nor U32163 (N_32163,N_31782,N_31914);
nand U32164 (N_32164,N_31937,N_31761);
and U32165 (N_32165,N_31808,N_31750);
nor U32166 (N_32166,N_31803,N_31750);
and U32167 (N_32167,N_31865,N_31913);
nor U32168 (N_32168,N_31928,N_31750);
nor U32169 (N_32169,N_31996,N_31921);
nand U32170 (N_32170,N_31858,N_31945);
or U32171 (N_32171,N_31769,N_31857);
nor U32172 (N_32172,N_31795,N_31848);
xnor U32173 (N_32173,N_31764,N_31971);
nand U32174 (N_32174,N_31814,N_31964);
nor U32175 (N_32175,N_31850,N_31984);
and U32176 (N_32176,N_31777,N_31901);
xor U32177 (N_32177,N_31969,N_31994);
xnor U32178 (N_32178,N_31821,N_31987);
nor U32179 (N_32179,N_31766,N_31875);
nor U32180 (N_32180,N_31810,N_31919);
nor U32181 (N_32181,N_31893,N_31833);
xnor U32182 (N_32182,N_31824,N_31757);
nand U32183 (N_32183,N_31864,N_31996);
and U32184 (N_32184,N_31838,N_31833);
nor U32185 (N_32185,N_31775,N_31930);
or U32186 (N_32186,N_31793,N_31895);
and U32187 (N_32187,N_31854,N_31991);
and U32188 (N_32188,N_31788,N_31808);
or U32189 (N_32189,N_31978,N_31801);
or U32190 (N_32190,N_31992,N_31849);
and U32191 (N_32191,N_31892,N_31883);
and U32192 (N_32192,N_31861,N_31753);
or U32193 (N_32193,N_31903,N_31920);
or U32194 (N_32194,N_31884,N_31860);
nand U32195 (N_32195,N_31952,N_31993);
nor U32196 (N_32196,N_31920,N_31756);
and U32197 (N_32197,N_31807,N_31953);
nor U32198 (N_32198,N_31787,N_31786);
nor U32199 (N_32199,N_31941,N_31989);
and U32200 (N_32200,N_31752,N_31808);
and U32201 (N_32201,N_31789,N_31759);
and U32202 (N_32202,N_31871,N_31791);
xnor U32203 (N_32203,N_31776,N_31885);
xor U32204 (N_32204,N_31917,N_31802);
or U32205 (N_32205,N_31774,N_31893);
nand U32206 (N_32206,N_31823,N_31781);
nand U32207 (N_32207,N_31974,N_31944);
or U32208 (N_32208,N_31961,N_31989);
nor U32209 (N_32209,N_31846,N_31923);
nor U32210 (N_32210,N_31751,N_31887);
nor U32211 (N_32211,N_31793,N_31803);
and U32212 (N_32212,N_31796,N_31906);
nor U32213 (N_32213,N_31978,N_31961);
nor U32214 (N_32214,N_31897,N_31800);
or U32215 (N_32215,N_31793,N_31913);
or U32216 (N_32216,N_31956,N_31756);
xnor U32217 (N_32217,N_31926,N_31798);
xor U32218 (N_32218,N_31989,N_31872);
or U32219 (N_32219,N_31787,N_31906);
and U32220 (N_32220,N_31967,N_31862);
and U32221 (N_32221,N_31830,N_31770);
and U32222 (N_32222,N_31829,N_31963);
nand U32223 (N_32223,N_31994,N_31766);
or U32224 (N_32224,N_31982,N_31972);
nand U32225 (N_32225,N_31893,N_31830);
or U32226 (N_32226,N_31995,N_31879);
nor U32227 (N_32227,N_31779,N_31990);
xnor U32228 (N_32228,N_31758,N_31921);
or U32229 (N_32229,N_31761,N_31850);
and U32230 (N_32230,N_31862,N_31885);
nand U32231 (N_32231,N_31967,N_31982);
or U32232 (N_32232,N_31985,N_31942);
or U32233 (N_32233,N_31904,N_31804);
nand U32234 (N_32234,N_31901,N_31997);
xor U32235 (N_32235,N_31864,N_31907);
or U32236 (N_32236,N_31986,N_31945);
and U32237 (N_32237,N_31796,N_31962);
nand U32238 (N_32238,N_31950,N_31918);
or U32239 (N_32239,N_31795,N_31944);
xor U32240 (N_32240,N_31916,N_31892);
or U32241 (N_32241,N_31752,N_31819);
nor U32242 (N_32242,N_31871,N_31836);
xor U32243 (N_32243,N_31938,N_31923);
xnor U32244 (N_32244,N_31926,N_31998);
and U32245 (N_32245,N_31842,N_31786);
xor U32246 (N_32246,N_31888,N_31755);
nand U32247 (N_32247,N_31817,N_31913);
nor U32248 (N_32248,N_31795,N_31782);
and U32249 (N_32249,N_31906,N_31833);
xor U32250 (N_32250,N_32061,N_32074);
xnor U32251 (N_32251,N_32131,N_32245);
nor U32252 (N_32252,N_32102,N_32030);
nor U32253 (N_32253,N_32123,N_32012);
and U32254 (N_32254,N_32170,N_32140);
xnor U32255 (N_32255,N_32180,N_32191);
xnor U32256 (N_32256,N_32053,N_32160);
and U32257 (N_32257,N_32081,N_32147);
nor U32258 (N_32258,N_32019,N_32073);
and U32259 (N_32259,N_32178,N_32117);
nand U32260 (N_32260,N_32168,N_32068);
or U32261 (N_32261,N_32247,N_32138);
xnor U32262 (N_32262,N_32060,N_32210);
or U32263 (N_32263,N_32221,N_32018);
and U32264 (N_32264,N_32033,N_32201);
and U32265 (N_32265,N_32200,N_32148);
xnor U32266 (N_32266,N_32126,N_32046);
or U32267 (N_32267,N_32152,N_32241);
and U32268 (N_32268,N_32238,N_32041);
xor U32269 (N_32269,N_32037,N_32101);
nor U32270 (N_32270,N_32194,N_32144);
and U32271 (N_32271,N_32009,N_32179);
nand U32272 (N_32272,N_32136,N_32235);
nor U32273 (N_32273,N_32202,N_32242);
nand U32274 (N_32274,N_32153,N_32005);
and U32275 (N_32275,N_32198,N_32130);
xnor U32276 (N_32276,N_32139,N_32055);
xnor U32277 (N_32277,N_32090,N_32013);
and U32278 (N_32278,N_32133,N_32026);
nor U32279 (N_32279,N_32028,N_32063);
and U32280 (N_32280,N_32038,N_32087);
xor U32281 (N_32281,N_32067,N_32181);
or U32282 (N_32282,N_32159,N_32157);
nand U32283 (N_32283,N_32092,N_32014);
nand U32284 (N_32284,N_32010,N_32127);
and U32285 (N_32285,N_32187,N_32118);
nand U32286 (N_32286,N_32069,N_32015);
nand U32287 (N_32287,N_32212,N_32007);
nand U32288 (N_32288,N_32171,N_32079);
xnor U32289 (N_32289,N_32035,N_32225);
nand U32290 (N_32290,N_32048,N_32184);
nand U32291 (N_32291,N_32166,N_32045);
nand U32292 (N_32292,N_32040,N_32236);
nor U32293 (N_32293,N_32229,N_32158);
nand U32294 (N_32294,N_32219,N_32192);
nand U32295 (N_32295,N_32151,N_32218);
and U32296 (N_32296,N_32155,N_32149);
and U32297 (N_32297,N_32039,N_32052);
or U32298 (N_32298,N_32084,N_32057);
nor U32299 (N_32299,N_32216,N_32188);
and U32300 (N_32300,N_32064,N_32124);
nor U32301 (N_32301,N_32213,N_32112);
nor U32302 (N_32302,N_32141,N_32116);
and U32303 (N_32303,N_32204,N_32240);
xnor U32304 (N_32304,N_32162,N_32075);
and U32305 (N_32305,N_32146,N_32108);
nor U32306 (N_32306,N_32121,N_32190);
and U32307 (N_32307,N_32020,N_32077);
xor U32308 (N_32308,N_32165,N_32056);
nor U32309 (N_32309,N_32243,N_32000);
or U32310 (N_32310,N_32177,N_32089);
or U32311 (N_32311,N_32017,N_32215);
and U32312 (N_32312,N_32095,N_32244);
or U32313 (N_32313,N_32071,N_32011);
xnor U32314 (N_32314,N_32206,N_32143);
nand U32315 (N_32315,N_32109,N_32163);
nand U32316 (N_32316,N_32232,N_32186);
nand U32317 (N_32317,N_32167,N_32226);
nand U32318 (N_32318,N_32085,N_32111);
and U32319 (N_32319,N_32249,N_32237);
or U32320 (N_32320,N_32208,N_32097);
and U32321 (N_32321,N_32128,N_32096);
nor U32322 (N_32322,N_32105,N_32199);
nand U32323 (N_32323,N_32022,N_32049);
xnor U32324 (N_32324,N_32025,N_32217);
xnor U32325 (N_32325,N_32161,N_32066);
nand U32326 (N_32326,N_32006,N_32003);
nor U32327 (N_32327,N_32134,N_32076);
nand U32328 (N_32328,N_32032,N_32093);
xnor U32329 (N_32329,N_32182,N_32233);
and U32330 (N_32330,N_32072,N_32195);
nand U32331 (N_32331,N_32175,N_32104);
and U32332 (N_32332,N_32172,N_32044);
and U32333 (N_32333,N_32125,N_32021);
xor U32334 (N_32334,N_32058,N_32246);
nor U32335 (N_32335,N_32135,N_32042);
xnor U32336 (N_32336,N_32114,N_32036);
and U32337 (N_32337,N_32034,N_32174);
or U32338 (N_32338,N_32164,N_32083);
xor U32339 (N_32339,N_32001,N_32004);
and U32340 (N_32340,N_32110,N_32016);
nand U32341 (N_32341,N_32065,N_32115);
nor U32342 (N_32342,N_32091,N_32086);
or U32343 (N_32343,N_32207,N_32142);
nor U32344 (N_32344,N_32024,N_32154);
nand U32345 (N_32345,N_32082,N_32231);
xnor U32346 (N_32346,N_32047,N_32119);
nor U32347 (N_32347,N_32228,N_32222);
xor U32348 (N_32348,N_32230,N_32107);
nor U32349 (N_32349,N_32197,N_32220);
nor U32350 (N_32350,N_32078,N_32088);
nor U32351 (N_32351,N_32080,N_32234);
nor U32352 (N_32352,N_32008,N_32203);
or U32353 (N_32353,N_32193,N_32027);
nor U32354 (N_32354,N_32223,N_32248);
and U32355 (N_32355,N_32137,N_32051);
xnor U32356 (N_32356,N_32050,N_32031);
nand U32357 (N_32357,N_32169,N_32224);
xor U32358 (N_32358,N_32099,N_32062);
nor U32359 (N_32359,N_32227,N_32002);
xor U32360 (N_32360,N_32145,N_32029);
nor U32361 (N_32361,N_32120,N_32054);
nor U32362 (N_32362,N_32129,N_32211);
and U32363 (N_32363,N_32132,N_32103);
and U32364 (N_32364,N_32122,N_32239);
nand U32365 (N_32365,N_32023,N_32100);
or U32366 (N_32366,N_32205,N_32176);
nor U32367 (N_32367,N_32214,N_32173);
and U32368 (N_32368,N_32183,N_32150);
xnor U32369 (N_32369,N_32196,N_32185);
or U32370 (N_32370,N_32098,N_32043);
and U32371 (N_32371,N_32094,N_32209);
xor U32372 (N_32372,N_32106,N_32156);
or U32373 (N_32373,N_32070,N_32113);
and U32374 (N_32374,N_32059,N_32189);
and U32375 (N_32375,N_32037,N_32144);
and U32376 (N_32376,N_32246,N_32122);
nand U32377 (N_32377,N_32014,N_32030);
xor U32378 (N_32378,N_32063,N_32110);
xor U32379 (N_32379,N_32186,N_32246);
and U32380 (N_32380,N_32163,N_32091);
and U32381 (N_32381,N_32138,N_32015);
nand U32382 (N_32382,N_32026,N_32168);
xor U32383 (N_32383,N_32080,N_32055);
or U32384 (N_32384,N_32079,N_32141);
nor U32385 (N_32385,N_32247,N_32106);
nand U32386 (N_32386,N_32198,N_32172);
or U32387 (N_32387,N_32179,N_32154);
or U32388 (N_32388,N_32069,N_32096);
xor U32389 (N_32389,N_32228,N_32051);
and U32390 (N_32390,N_32110,N_32156);
or U32391 (N_32391,N_32209,N_32026);
xor U32392 (N_32392,N_32103,N_32131);
nand U32393 (N_32393,N_32084,N_32063);
nor U32394 (N_32394,N_32026,N_32188);
nor U32395 (N_32395,N_32021,N_32109);
and U32396 (N_32396,N_32070,N_32181);
or U32397 (N_32397,N_32137,N_32190);
nor U32398 (N_32398,N_32235,N_32014);
or U32399 (N_32399,N_32228,N_32198);
nor U32400 (N_32400,N_32199,N_32092);
xnor U32401 (N_32401,N_32178,N_32112);
xor U32402 (N_32402,N_32206,N_32112);
and U32403 (N_32403,N_32184,N_32010);
nand U32404 (N_32404,N_32042,N_32228);
nand U32405 (N_32405,N_32234,N_32232);
and U32406 (N_32406,N_32168,N_32137);
and U32407 (N_32407,N_32072,N_32013);
and U32408 (N_32408,N_32131,N_32104);
or U32409 (N_32409,N_32172,N_32025);
nand U32410 (N_32410,N_32249,N_32231);
nand U32411 (N_32411,N_32081,N_32141);
xor U32412 (N_32412,N_32233,N_32175);
nor U32413 (N_32413,N_32019,N_32142);
xnor U32414 (N_32414,N_32213,N_32011);
xnor U32415 (N_32415,N_32006,N_32162);
and U32416 (N_32416,N_32076,N_32009);
or U32417 (N_32417,N_32020,N_32166);
xnor U32418 (N_32418,N_32140,N_32238);
or U32419 (N_32419,N_32029,N_32238);
nor U32420 (N_32420,N_32241,N_32058);
xnor U32421 (N_32421,N_32206,N_32085);
nand U32422 (N_32422,N_32021,N_32120);
nand U32423 (N_32423,N_32214,N_32092);
or U32424 (N_32424,N_32110,N_32026);
nand U32425 (N_32425,N_32159,N_32130);
or U32426 (N_32426,N_32229,N_32023);
or U32427 (N_32427,N_32007,N_32100);
or U32428 (N_32428,N_32057,N_32247);
or U32429 (N_32429,N_32137,N_32125);
and U32430 (N_32430,N_32244,N_32100);
or U32431 (N_32431,N_32213,N_32127);
nor U32432 (N_32432,N_32177,N_32070);
nor U32433 (N_32433,N_32209,N_32076);
nor U32434 (N_32434,N_32159,N_32200);
nor U32435 (N_32435,N_32108,N_32084);
xnor U32436 (N_32436,N_32151,N_32133);
xor U32437 (N_32437,N_32135,N_32152);
or U32438 (N_32438,N_32245,N_32018);
nand U32439 (N_32439,N_32049,N_32183);
nor U32440 (N_32440,N_32195,N_32111);
nor U32441 (N_32441,N_32229,N_32233);
or U32442 (N_32442,N_32105,N_32163);
or U32443 (N_32443,N_32021,N_32055);
and U32444 (N_32444,N_32028,N_32140);
xnor U32445 (N_32445,N_32071,N_32028);
nor U32446 (N_32446,N_32183,N_32109);
nand U32447 (N_32447,N_32010,N_32239);
nor U32448 (N_32448,N_32060,N_32032);
and U32449 (N_32449,N_32019,N_32065);
or U32450 (N_32450,N_32138,N_32060);
nand U32451 (N_32451,N_32172,N_32048);
nand U32452 (N_32452,N_32006,N_32013);
or U32453 (N_32453,N_32012,N_32007);
and U32454 (N_32454,N_32223,N_32061);
nor U32455 (N_32455,N_32123,N_32031);
or U32456 (N_32456,N_32236,N_32155);
or U32457 (N_32457,N_32076,N_32114);
and U32458 (N_32458,N_32130,N_32002);
and U32459 (N_32459,N_32000,N_32077);
nand U32460 (N_32460,N_32071,N_32018);
xnor U32461 (N_32461,N_32210,N_32224);
xor U32462 (N_32462,N_32014,N_32142);
nor U32463 (N_32463,N_32106,N_32020);
nor U32464 (N_32464,N_32057,N_32167);
xnor U32465 (N_32465,N_32170,N_32016);
or U32466 (N_32466,N_32062,N_32203);
or U32467 (N_32467,N_32064,N_32025);
nand U32468 (N_32468,N_32085,N_32080);
xor U32469 (N_32469,N_32006,N_32137);
nand U32470 (N_32470,N_32221,N_32138);
or U32471 (N_32471,N_32247,N_32077);
and U32472 (N_32472,N_32186,N_32071);
xnor U32473 (N_32473,N_32050,N_32181);
nor U32474 (N_32474,N_32118,N_32032);
nor U32475 (N_32475,N_32231,N_32233);
nor U32476 (N_32476,N_32179,N_32189);
or U32477 (N_32477,N_32161,N_32145);
xor U32478 (N_32478,N_32182,N_32027);
and U32479 (N_32479,N_32037,N_32202);
and U32480 (N_32480,N_32166,N_32010);
nand U32481 (N_32481,N_32109,N_32081);
nand U32482 (N_32482,N_32021,N_32064);
nor U32483 (N_32483,N_32106,N_32048);
and U32484 (N_32484,N_32204,N_32127);
and U32485 (N_32485,N_32053,N_32069);
xor U32486 (N_32486,N_32045,N_32198);
xor U32487 (N_32487,N_32159,N_32057);
nor U32488 (N_32488,N_32057,N_32015);
and U32489 (N_32489,N_32112,N_32192);
nand U32490 (N_32490,N_32237,N_32234);
and U32491 (N_32491,N_32208,N_32146);
or U32492 (N_32492,N_32004,N_32029);
and U32493 (N_32493,N_32200,N_32047);
nand U32494 (N_32494,N_32215,N_32043);
or U32495 (N_32495,N_32184,N_32106);
and U32496 (N_32496,N_32203,N_32054);
and U32497 (N_32497,N_32145,N_32051);
nand U32498 (N_32498,N_32065,N_32164);
nand U32499 (N_32499,N_32092,N_32115);
nor U32500 (N_32500,N_32410,N_32267);
or U32501 (N_32501,N_32304,N_32305);
xnor U32502 (N_32502,N_32395,N_32332);
nor U32503 (N_32503,N_32470,N_32336);
and U32504 (N_32504,N_32432,N_32442);
nor U32505 (N_32505,N_32309,N_32359);
or U32506 (N_32506,N_32375,N_32486);
xnor U32507 (N_32507,N_32427,N_32352);
or U32508 (N_32508,N_32421,N_32324);
nor U32509 (N_32509,N_32483,N_32406);
nor U32510 (N_32510,N_32268,N_32314);
nand U32511 (N_32511,N_32413,N_32398);
nor U32512 (N_32512,N_32482,N_32255);
and U32513 (N_32513,N_32489,N_32487);
and U32514 (N_32514,N_32298,N_32380);
and U32515 (N_32515,N_32257,N_32390);
and U32516 (N_32516,N_32274,N_32408);
or U32517 (N_32517,N_32308,N_32460);
or U32518 (N_32518,N_32364,N_32490);
or U32519 (N_32519,N_32402,N_32423);
nor U32520 (N_32520,N_32358,N_32383);
and U32521 (N_32521,N_32291,N_32493);
nor U32522 (N_32522,N_32295,N_32450);
and U32523 (N_32523,N_32347,N_32430);
or U32524 (N_32524,N_32447,N_32429);
and U32525 (N_32525,N_32376,N_32286);
and U32526 (N_32526,N_32302,N_32277);
xor U32527 (N_32527,N_32435,N_32259);
and U32528 (N_32528,N_32338,N_32321);
nor U32529 (N_32529,N_32272,N_32443);
nor U32530 (N_32530,N_32253,N_32307);
nand U32531 (N_32531,N_32265,N_32288);
nand U32532 (N_32532,N_32351,N_32373);
xnor U32533 (N_32533,N_32488,N_32439);
or U32534 (N_32534,N_32287,N_32475);
nor U32535 (N_32535,N_32451,N_32329);
nor U32536 (N_32536,N_32280,N_32312);
xnor U32537 (N_32537,N_32294,N_32454);
nor U32538 (N_32538,N_32340,N_32261);
nand U32539 (N_32539,N_32455,N_32326);
nand U32540 (N_32540,N_32392,N_32260);
or U32541 (N_32541,N_32252,N_32330);
nand U32542 (N_32542,N_32316,N_32419);
nor U32543 (N_32543,N_32285,N_32424);
or U32544 (N_32544,N_32317,N_32471);
and U32545 (N_32545,N_32325,N_32420);
or U32546 (N_32546,N_32296,N_32355);
nor U32547 (N_32547,N_32356,N_32446);
nor U32548 (N_32548,N_32464,N_32499);
or U32549 (N_32549,N_32496,N_32431);
nand U32550 (N_32550,N_32281,N_32331);
or U32551 (N_32551,N_32284,N_32414);
xor U32552 (N_32552,N_32441,N_32494);
nor U32553 (N_32553,N_32337,N_32485);
nor U32554 (N_32554,N_32382,N_32365);
or U32555 (N_32555,N_32399,N_32251);
xnor U32556 (N_32556,N_32405,N_32346);
xnor U32557 (N_32557,N_32467,N_32264);
and U32558 (N_32558,N_32480,N_32306);
nor U32559 (N_32559,N_32437,N_32387);
xnor U32560 (N_32560,N_32403,N_32492);
and U32561 (N_32561,N_32448,N_32457);
xnor U32562 (N_32562,N_32449,N_32444);
and U32563 (N_32563,N_32293,N_32456);
nor U32564 (N_32564,N_32438,N_32472);
or U32565 (N_32565,N_32458,N_32354);
nand U32566 (N_32566,N_32400,N_32436);
or U32567 (N_32567,N_32301,N_32303);
xor U32568 (N_32568,N_32391,N_32319);
xnor U32569 (N_32569,N_32478,N_32341);
and U32570 (N_32570,N_32310,N_32323);
nand U32571 (N_32571,N_32378,N_32369);
nand U32572 (N_32572,N_32381,N_32466);
xor U32573 (N_32573,N_32385,N_32275);
nand U32574 (N_32574,N_32290,N_32327);
or U32575 (N_32575,N_32320,N_32394);
and U32576 (N_32576,N_32418,N_32269);
xnor U32577 (N_32577,N_32425,N_32254);
and U32578 (N_32578,N_32463,N_32256);
nand U32579 (N_32579,N_32417,N_32271);
nor U32580 (N_32580,N_32292,N_32397);
and U32581 (N_32581,N_32426,N_32416);
or U32582 (N_32582,N_32297,N_32453);
xnor U32583 (N_32583,N_32318,N_32481);
nand U32584 (N_32584,N_32282,N_32357);
nand U32585 (N_32585,N_32388,N_32434);
nand U32586 (N_32586,N_32322,N_32283);
xor U32587 (N_32587,N_32404,N_32445);
xnor U32588 (N_32588,N_32299,N_32409);
and U32589 (N_32589,N_32333,N_32345);
or U32590 (N_32590,N_32495,N_32279);
nor U32591 (N_32591,N_32393,N_32497);
nand U32592 (N_32592,N_32343,N_32350);
nor U32593 (N_32593,N_32368,N_32384);
nand U32594 (N_32594,N_32367,N_32353);
xor U32595 (N_32595,N_32372,N_32311);
and U32596 (N_32596,N_32468,N_32411);
or U32597 (N_32597,N_32362,N_32349);
nand U32598 (N_32598,N_32379,N_32498);
nor U32599 (N_32599,N_32491,N_32263);
and U32600 (N_32600,N_32270,N_32377);
nor U32601 (N_32601,N_32289,N_32396);
nand U32602 (N_32602,N_32334,N_32469);
or U32603 (N_32603,N_32250,N_32370);
or U32604 (N_32604,N_32407,N_32262);
xnor U32605 (N_32605,N_32278,N_32452);
or U32606 (N_32606,N_32273,N_32276);
nand U32607 (N_32607,N_32371,N_32348);
xor U32608 (N_32608,N_32465,N_32374);
and U32609 (N_32609,N_32428,N_32461);
and U32610 (N_32610,N_32361,N_32258);
nand U32611 (N_32611,N_32328,N_32474);
nand U32612 (N_32612,N_32479,N_32433);
nor U32613 (N_32613,N_32363,N_32266);
and U32614 (N_32614,N_32440,N_32484);
and U32615 (N_32615,N_32389,N_32477);
or U32616 (N_32616,N_32342,N_32415);
and U32617 (N_32617,N_32300,N_32422);
or U32618 (N_32618,N_32366,N_32386);
nor U32619 (N_32619,N_32473,N_32360);
or U32620 (N_32620,N_32335,N_32401);
xnor U32621 (N_32621,N_32344,N_32315);
or U32622 (N_32622,N_32339,N_32462);
or U32623 (N_32623,N_32459,N_32412);
or U32624 (N_32624,N_32476,N_32313);
xnor U32625 (N_32625,N_32269,N_32463);
or U32626 (N_32626,N_32354,N_32323);
xor U32627 (N_32627,N_32327,N_32337);
nor U32628 (N_32628,N_32445,N_32391);
xnor U32629 (N_32629,N_32363,N_32312);
nand U32630 (N_32630,N_32315,N_32484);
and U32631 (N_32631,N_32379,N_32273);
nand U32632 (N_32632,N_32293,N_32467);
or U32633 (N_32633,N_32327,N_32495);
xnor U32634 (N_32634,N_32309,N_32455);
and U32635 (N_32635,N_32419,N_32435);
nand U32636 (N_32636,N_32378,N_32298);
xor U32637 (N_32637,N_32472,N_32331);
nand U32638 (N_32638,N_32283,N_32361);
and U32639 (N_32639,N_32290,N_32497);
nor U32640 (N_32640,N_32405,N_32461);
and U32641 (N_32641,N_32484,N_32434);
or U32642 (N_32642,N_32294,N_32365);
nand U32643 (N_32643,N_32392,N_32326);
nor U32644 (N_32644,N_32297,N_32423);
and U32645 (N_32645,N_32365,N_32360);
and U32646 (N_32646,N_32439,N_32338);
and U32647 (N_32647,N_32348,N_32369);
nand U32648 (N_32648,N_32270,N_32492);
nor U32649 (N_32649,N_32396,N_32335);
or U32650 (N_32650,N_32295,N_32473);
nand U32651 (N_32651,N_32408,N_32451);
or U32652 (N_32652,N_32427,N_32472);
and U32653 (N_32653,N_32281,N_32344);
or U32654 (N_32654,N_32426,N_32287);
nand U32655 (N_32655,N_32391,N_32464);
xnor U32656 (N_32656,N_32429,N_32414);
nor U32657 (N_32657,N_32379,N_32324);
nor U32658 (N_32658,N_32468,N_32408);
xor U32659 (N_32659,N_32280,N_32469);
xor U32660 (N_32660,N_32469,N_32331);
nand U32661 (N_32661,N_32392,N_32410);
nand U32662 (N_32662,N_32475,N_32497);
nor U32663 (N_32663,N_32445,N_32440);
xor U32664 (N_32664,N_32449,N_32481);
and U32665 (N_32665,N_32333,N_32466);
or U32666 (N_32666,N_32345,N_32417);
and U32667 (N_32667,N_32496,N_32294);
or U32668 (N_32668,N_32357,N_32304);
and U32669 (N_32669,N_32399,N_32477);
or U32670 (N_32670,N_32395,N_32338);
xor U32671 (N_32671,N_32441,N_32424);
nand U32672 (N_32672,N_32445,N_32420);
and U32673 (N_32673,N_32278,N_32331);
xor U32674 (N_32674,N_32316,N_32384);
nand U32675 (N_32675,N_32426,N_32403);
xor U32676 (N_32676,N_32343,N_32451);
or U32677 (N_32677,N_32399,N_32390);
and U32678 (N_32678,N_32435,N_32327);
or U32679 (N_32679,N_32281,N_32394);
or U32680 (N_32680,N_32452,N_32305);
nand U32681 (N_32681,N_32401,N_32321);
nand U32682 (N_32682,N_32487,N_32361);
or U32683 (N_32683,N_32327,N_32391);
or U32684 (N_32684,N_32328,N_32294);
or U32685 (N_32685,N_32451,N_32446);
and U32686 (N_32686,N_32420,N_32322);
nand U32687 (N_32687,N_32293,N_32264);
xor U32688 (N_32688,N_32316,N_32275);
xor U32689 (N_32689,N_32411,N_32307);
nand U32690 (N_32690,N_32353,N_32403);
nor U32691 (N_32691,N_32328,N_32440);
nand U32692 (N_32692,N_32383,N_32360);
or U32693 (N_32693,N_32411,N_32467);
nand U32694 (N_32694,N_32456,N_32423);
or U32695 (N_32695,N_32381,N_32342);
or U32696 (N_32696,N_32328,N_32333);
and U32697 (N_32697,N_32396,N_32337);
nor U32698 (N_32698,N_32403,N_32297);
xnor U32699 (N_32699,N_32318,N_32419);
nand U32700 (N_32700,N_32373,N_32384);
and U32701 (N_32701,N_32284,N_32425);
and U32702 (N_32702,N_32266,N_32367);
nor U32703 (N_32703,N_32466,N_32287);
nor U32704 (N_32704,N_32296,N_32278);
nor U32705 (N_32705,N_32306,N_32330);
xnor U32706 (N_32706,N_32426,N_32496);
nor U32707 (N_32707,N_32322,N_32363);
or U32708 (N_32708,N_32330,N_32270);
nand U32709 (N_32709,N_32322,N_32344);
nand U32710 (N_32710,N_32448,N_32388);
and U32711 (N_32711,N_32404,N_32365);
nand U32712 (N_32712,N_32373,N_32447);
nor U32713 (N_32713,N_32402,N_32259);
and U32714 (N_32714,N_32472,N_32400);
nand U32715 (N_32715,N_32419,N_32406);
nand U32716 (N_32716,N_32402,N_32351);
xnor U32717 (N_32717,N_32483,N_32359);
xor U32718 (N_32718,N_32280,N_32281);
nor U32719 (N_32719,N_32353,N_32268);
nor U32720 (N_32720,N_32257,N_32256);
nor U32721 (N_32721,N_32297,N_32355);
nor U32722 (N_32722,N_32422,N_32323);
or U32723 (N_32723,N_32380,N_32324);
or U32724 (N_32724,N_32256,N_32258);
xor U32725 (N_32725,N_32296,N_32426);
and U32726 (N_32726,N_32460,N_32453);
xor U32727 (N_32727,N_32478,N_32274);
or U32728 (N_32728,N_32446,N_32425);
xor U32729 (N_32729,N_32403,N_32376);
nand U32730 (N_32730,N_32419,N_32434);
xor U32731 (N_32731,N_32405,N_32310);
and U32732 (N_32732,N_32395,N_32471);
or U32733 (N_32733,N_32379,N_32286);
or U32734 (N_32734,N_32275,N_32330);
xor U32735 (N_32735,N_32423,N_32274);
nor U32736 (N_32736,N_32486,N_32293);
nand U32737 (N_32737,N_32444,N_32349);
or U32738 (N_32738,N_32287,N_32349);
nand U32739 (N_32739,N_32492,N_32468);
nand U32740 (N_32740,N_32277,N_32438);
nor U32741 (N_32741,N_32379,N_32302);
nand U32742 (N_32742,N_32394,N_32442);
nand U32743 (N_32743,N_32493,N_32489);
and U32744 (N_32744,N_32296,N_32300);
xnor U32745 (N_32745,N_32251,N_32358);
and U32746 (N_32746,N_32347,N_32463);
and U32747 (N_32747,N_32331,N_32335);
xor U32748 (N_32748,N_32435,N_32274);
or U32749 (N_32749,N_32452,N_32431);
nand U32750 (N_32750,N_32506,N_32540);
nand U32751 (N_32751,N_32590,N_32505);
and U32752 (N_32752,N_32558,N_32502);
or U32753 (N_32753,N_32651,N_32567);
nand U32754 (N_32754,N_32745,N_32622);
or U32755 (N_32755,N_32693,N_32671);
nor U32756 (N_32756,N_32726,N_32638);
xor U32757 (N_32757,N_32549,N_32574);
xor U32758 (N_32758,N_32737,N_32668);
or U32759 (N_32759,N_32636,N_32727);
xor U32760 (N_32760,N_32521,N_32542);
or U32761 (N_32761,N_32621,N_32679);
xor U32762 (N_32762,N_32717,N_32695);
or U32763 (N_32763,N_32568,N_32701);
nor U32764 (N_32764,N_32708,N_32605);
and U32765 (N_32765,N_32665,N_32612);
nand U32766 (N_32766,N_32527,N_32699);
nand U32767 (N_32767,N_32631,N_32584);
nand U32768 (N_32768,N_32735,N_32704);
or U32769 (N_32769,N_32738,N_32697);
nor U32770 (N_32770,N_32732,N_32640);
or U32771 (N_32771,N_32518,N_32620);
or U32772 (N_32772,N_32610,N_32741);
and U32773 (N_32773,N_32661,N_32734);
and U32774 (N_32774,N_32560,N_32725);
nor U32775 (N_32775,N_32513,N_32552);
or U32776 (N_32776,N_32592,N_32746);
or U32777 (N_32777,N_32654,N_32594);
nand U32778 (N_32778,N_32722,N_32642);
nor U32779 (N_32779,N_32575,N_32660);
nand U32780 (N_32780,N_32511,N_32514);
or U32781 (N_32781,N_32517,N_32707);
and U32782 (N_32782,N_32503,N_32559);
and U32783 (N_32783,N_32625,N_32616);
nor U32784 (N_32784,N_32563,N_32565);
nor U32785 (N_32785,N_32507,N_32510);
nand U32786 (N_32786,N_32623,N_32687);
xnor U32787 (N_32787,N_32535,N_32644);
nor U32788 (N_32788,N_32652,N_32508);
or U32789 (N_32789,N_32674,N_32710);
or U32790 (N_32790,N_32730,N_32677);
or U32791 (N_32791,N_32706,N_32676);
and U32792 (N_32792,N_32711,N_32599);
and U32793 (N_32793,N_32553,N_32615);
and U32794 (N_32794,N_32541,N_32512);
nand U32795 (N_32795,N_32709,N_32650);
nand U32796 (N_32796,N_32723,N_32538);
and U32797 (N_32797,N_32606,N_32600);
or U32798 (N_32798,N_32694,N_32739);
and U32799 (N_32799,N_32587,N_32536);
or U32800 (N_32800,N_32597,N_32678);
nand U32801 (N_32801,N_32686,N_32670);
nor U32802 (N_32802,N_32532,N_32653);
and U32803 (N_32803,N_32613,N_32509);
xor U32804 (N_32804,N_32595,N_32525);
nand U32805 (N_32805,N_32718,N_32534);
and U32806 (N_32806,N_32596,N_32672);
or U32807 (N_32807,N_32635,N_32626);
and U32808 (N_32808,N_32608,N_32659);
or U32809 (N_32809,N_32747,N_32529);
xnor U32810 (N_32810,N_32682,N_32743);
nand U32811 (N_32811,N_32641,N_32580);
and U32812 (N_32812,N_32680,N_32664);
nand U32813 (N_32813,N_32729,N_32548);
nand U32814 (N_32814,N_32602,N_32705);
and U32815 (N_32815,N_32689,N_32688);
xnor U32816 (N_32816,N_32572,N_32633);
xor U32817 (N_32817,N_32581,N_32551);
and U32818 (N_32818,N_32658,N_32524);
nor U32819 (N_32819,N_32649,N_32618);
nand U32820 (N_32820,N_32673,N_32576);
nand U32821 (N_32821,N_32571,N_32564);
and U32822 (N_32822,N_32691,N_32634);
or U32823 (N_32823,N_32582,N_32583);
xnor U32824 (N_32824,N_32639,N_32562);
nor U32825 (N_32825,N_32528,N_32632);
nor U32826 (N_32826,N_32555,N_32539);
nand U32827 (N_32827,N_32504,N_32585);
nand U32828 (N_32828,N_32724,N_32611);
or U32829 (N_32829,N_32619,N_32692);
nor U32830 (N_32830,N_32557,N_32545);
xnor U32831 (N_32831,N_32713,N_32591);
nand U32832 (N_32832,N_32593,N_32515);
and U32833 (N_32833,N_32603,N_32744);
or U32834 (N_32834,N_32643,N_32614);
xor U32835 (N_32835,N_32516,N_32533);
and U32836 (N_32836,N_32749,N_32566);
nor U32837 (N_32837,N_32685,N_32712);
and U32838 (N_32838,N_32628,N_32501);
and U32839 (N_32839,N_32667,N_32531);
nand U32840 (N_32840,N_32655,N_32681);
nand U32841 (N_32841,N_32609,N_32646);
nor U32842 (N_32842,N_32648,N_32579);
and U32843 (N_32843,N_32696,N_32662);
nand U32844 (N_32844,N_32526,N_32637);
and U32845 (N_32845,N_32720,N_32546);
or U32846 (N_32846,N_32588,N_32740);
xnor U32847 (N_32847,N_32573,N_32543);
and U32848 (N_32848,N_32537,N_32684);
nor U32849 (N_32849,N_32715,N_32666);
nand U32850 (N_32850,N_32647,N_32577);
or U32851 (N_32851,N_32663,N_32656);
xor U32852 (N_32852,N_32547,N_32522);
or U32853 (N_32853,N_32731,N_32561);
and U32854 (N_32854,N_32624,N_32570);
and U32855 (N_32855,N_32554,N_32748);
or U32856 (N_32856,N_32530,N_32657);
xor U32857 (N_32857,N_32721,N_32728);
nor U32858 (N_32858,N_32607,N_32742);
nand U32859 (N_32859,N_32716,N_32589);
nand U32860 (N_32860,N_32569,N_32578);
nand U32861 (N_32861,N_32675,N_32520);
or U32862 (N_32862,N_32519,N_32586);
nand U32863 (N_32863,N_32736,N_32703);
and U32864 (N_32864,N_32698,N_32645);
nor U32865 (N_32865,N_32630,N_32702);
nand U32866 (N_32866,N_32719,N_32669);
xor U32867 (N_32867,N_32550,N_32700);
nor U32868 (N_32868,N_32556,N_32629);
nor U32869 (N_32869,N_32544,N_32604);
or U32870 (N_32870,N_32714,N_32598);
nand U32871 (N_32871,N_32601,N_32690);
or U32872 (N_32872,N_32683,N_32523);
nor U32873 (N_32873,N_32500,N_32733);
or U32874 (N_32874,N_32627,N_32617);
nor U32875 (N_32875,N_32641,N_32664);
nand U32876 (N_32876,N_32647,N_32507);
and U32877 (N_32877,N_32649,N_32611);
xor U32878 (N_32878,N_32649,N_32520);
or U32879 (N_32879,N_32723,N_32711);
or U32880 (N_32880,N_32519,N_32587);
nor U32881 (N_32881,N_32699,N_32563);
and U32882 (N_32882,N_32671,N_32597);
and U32883 (N_32883,N_32710,N_32568);
and U32884 (N_32884,N_32657,N_32593);
nand U32885 (N_32885,N_32521,N_32544);
and U32886 (N_32886,N_32579,N_32675);
nor U32887 (N_32887,N_32715,N_32585);
xnor U32888 (N_32888,N_32737,N_32617);
xnor U32889 (N_32889,N_32545,N_32601);
xor U32890 (N_32890,N_32534,N_32529);
xnor U32891 (N_32891,N_32623,N_32502);
xnor U32892 (N_32892,N_32576,N_32719);
or U32893 (N_32893,N_32684,N_32699);
nand U32894 (N_32894,N_32692,N_32614);
nor U32895 (N_32895,N_32571,N_32685);
nor U32896 (N_32896,N_32746,N_32672);
or U32897 (N_32897,N_32736,N_32593);
nor U32898 (N_32898,N_32571,N_32554);
and U32899 (N_32899,N_32646,N_32736);
nor U32900 (N_32900,N_32575,N_32553);
nor U32901 (N_32901,N_32742,N_32553);
xnor U32902 (N_32902,N_32508,N_32540);
xor U32903 (N_32903,N_32621,N_32615);
xor U32904 (N_32904,N_32542,N_32554);
nand U32905 (N_32905,N_32650,N_32510);
or U32906 (N_32906,N_32564,N_32581);
nor U32907 (N_32907,N_32569,N_32730);
nand U32908 (N_32908,N_32720,N_32539);
nor U32909 (N_32909,N_32726,N_32639);
nor U32910 (N_32910,N_32532,N_32585);
nor U32911 (N_32911,N_32616,N_32628);
nand U32912 (N_32912,N_32545,N_32510);
or U32913 (N_32913,N_32507,N_32522);
or U32914 (N_32914,N_32718,N_32694);
and U32915 (N_32915,N_32527,N_32577);
nor U32916 (N_32916,N_32729,N_32688);
or U32917 (N_32917,N_32665,N_32562);
or U32918 (N_32918,N_32583,N_32632);
nor U32919 (N_32919,N_32737,N_32604);
nor U32920 (N_32920,N_32533,N_32687);
nand U32921 (N_32921,N_32714,N_32620);
or U32922 (N_32922,N_32723,N_32664);
nor U32923 (N_32923,N_32522,N_32700);
or U32924 (N_32924,N_32614,N_32506);
or U32925 (N_32925,N_32600,N_32583);
nand U32926 (N_32926,N_32739,N_32519);
nor U32927 (N_32927,N_32638,N_32690);
or U32928 (N_32928,N_32675,N_32576);
nor U32929 (N_32929,N_32523,N_32564);
and U32930 (N_32930,N_32504,N_32534);
nand U32931 (N_32931,N_32628,N_32595);
xor U32932 (N_32932,N_32700,N_32653);
nor U32933 (N_32933,N_32678,N_32742);
and U32934 (N_32934,N_32501,N_32648);
and U32935 (N_32935,N_32616,N_32647);
nor U32936 (N_32936,N_32745,N_32747);
nor U32937 (N_32937,N_32537,N_32717);
nor U32938 (N_32938,N_32708,N_32603);
xor U32939 (N_32939,N_32607,N_32745);
nand U32940 (N_32940,N_32573,N_32715);
nand U32941 (N_32941,N_32748,N_32747);
and U32942 (N_32942,N_32662,N_32741);
nor U32943 (N_32943,N_32595,N_32510);
and U32944 (N_32944,N_32704,N_32553);
nor U32945 (N_32945,N_32508,N_32519);
xor U32946 (N_32946,N_32614,N_32629);
or U32947 (N_32947,N_32621,N_32673);
nand U32948 (N_32948,N_32535,N_32519);
nand U32949 (N_32949,N_32712,N_32723);
xor U32950 (N_32950,N_32732,N_32598);
or U32951 (N_32951,N_32530,N_32676);
and U32952 (N_32952,N_32673,N_32701);
nand U32953 (N_32953,N_32614,N_32579);
or U32954 (N_32954,N_32745,N_32718);
or U32955 (N_32955,N_32692,N_32645);
nand U32956 (N_32956,N_32544,N_32560);
nor U32957 (N_32957,N_32530,N_32709);
xnor U32958 (N_32958,N_32568,N_32655);
nand U32959 (N_32959,N_32503,N_32514);
nand U32960 (N_32960,N_32616,N_32578);
or U32961 (N_32961,N_32673,N_32584);
nor U32962 (N_32962,N_32624,N_32562);
nor U32963 (N_32963,N_32578,N_32592);
xnor U32964 (N_32964,N_32630,N_32586);
nor U32965 (N_32965,N_32663,N_32518);
xor U32966 (N_32966,N_32539,N_32679);
xor U32967 (N_32967,N_32619,N_32647);
nand U32968 (N_32968,N_32525,N_32603);
and U32969 (N_32969,N_32660,N_32738);
nor U32970 (N_32970,N_32520,N_32692);
nor U32971 (N_32971,N_32664,N_32615);
xnor U32972 (N_32972,N_32550,N_32721);
and U32973 (N_32973,N_32707,N_32560);
xor U32974 (N_32974,N_32537,N_32715);
or U32975 (N_32975,N_32687,N_32578);
nor U32976 (N_32976,N_32713,N_32680);
nor U32977 (N_32977,N_32532,N_32694);
xnor U32978 (N_32978,N_32535,N_32609);
xor U32979 (N_32979,N_32606,N_32691);
nor U32980 (N_32980,N_32533,N_32588);
and U32981 (N_32981,N_32586,N_32729);
xor U32982 (N_32982,N_32730,N_32610);
nand U32983 (N_32983,N_32717,N_32611);
nand U32984 (N_32984,N_32745,N_32501);
xnor U32985 (N_32985,N_32744,N_32604);
nor U32986 (N_32986,N_32506,N_32558);
nand U32987 (N_32987,N_32606,N_32622);
and U32988 (N_32988,N_32550,N_32675);
nor U32989 (N_32989,N_32612,N_32686);
and U32990 (N_32990,N_32578,N_32583);
nor U32991 (N_32991,N_32536,N_32599);
and U32992 (N_32992,N_32556,N_32596);
xor U32993 (N_32993,N_32717,N_32737);
and U32994 (N_32994,N_32708,N_32575);
and U32995 (N_32995,N_32697,N_32663);
and U32996 (N_32996,N_32524,N_32701);
xor U32997 (N_32997,N_32664,N_32650);
and U32998 (N_32998,N_32729,N_32668);
or U32999 (N_32999,N_32584,N_32640);
xor U33000 (N_33000,N_32999,N_32817);
and U33001 (N_33001,N_32782,N_32783);
nand U33002 (N_33002,N_32830,N_32771);
or U33003 (N_33003,N_32810,N_32892);
nor U33004 (N_33004,N_32889,N_32964);
and U33005 (N_33005,N_32870,N_32957);
nor U33006 (N_33006,N_32805,N_32822);
and U33007 (N_33007,N_32881,N_32750);
nor U33008 (N_33008,N_32751,N_32812);
and U33009 (N_33009,N_32928,N_32987);
nand U33010 (N_33010,N_32818,N_32958);
nand U33011 (N_33011,N_32918,N_32763);
or U33012 (N_33012,N_32843,N_32895);
or U33013 (N_33013,N_32922,N_32886);
or U33014 (N_33014,N_32894,N_32756);
nand U33015 (N_33015,N_32953,N_32914);
nor U33016 (N_33016,N_32754,N_32753);
nor U33017 (N_33017,N_32997,N_32982);
nand U33018 (N_33018,N_32853,N_32841);
and U33019 (N_33019,N_32758,N_32855);
or U33020 (N_33020,N_32992,N_32806);
nand U33021 (N_33021,N_32963,N_32814);
or U33022 (N_33022,N_32784,N_32905);
nand U33023 (N_33023,N_32872,N_32973);
xor U33024 (N_33024,N_32926,N_32901);
and U33025 (N_33025,N_32865,N_32773);
xnor U33026 (N_33026,N_32891,N_32885);
nor U33027 (N_33027,N_32854,N_32815);
nor U33028 (N_33028,N_32788,N_32775);
nand U33029 (N_33029,N_32835,N_32868);
xnor U33030 (N_33030,N_32799,N_32871);
and U33031 (N_33031,N_32764,N_32893);
nor U33032 (N_33032,N_32800,N_32789);
nor U33033 (N_33033,N_32794,N_32925);
and U33034 (N_33034,N_32755,N_32832);
and U33035 (N_33035,N_32796,N_32777);
nor U33036 (N_33036,N_32945,N_32920);
and U33037 (N_33037,N_32867,N_32828);
nand U33038 (N_33038,N_32848,N_32765);
or U33039 (N_33039,N_32911,N_32898);
and U33040 (N_33040,N_32908,N_32974);
or U33041 (N_33041,N_32803,N_32860);
or U33042 (N_33042,N_32962,N_32966);
nor U33043 (N_33043,N_32847,N_32787);
nand U33044 (N_33044,N_32846,N_32781);
xor U33045 (N_33045,N_32861,N_32790);
and U33046 (N_33046,N_32996,N_32932);
xnor U33047 (N_33047,N_32952,N_32995);
and U33048 (N_33048,N_32943,N_32998);
or U33049 (N_33049,N_32831,N_32917);
nand U33050 (N_33050,N_32845,N_32804);
or U33051 (N_33051,N_32821,N_32791);
and U33052 (N_33052,N_32864,N_32772);
xnor U33053 (N_33053,N_32856,N_32769);
xnor U33054 (N_33054,N_32915,N_32874);
nor U33055 (N_33055,N_32850,N_32933);
xor U33056 (N_33056,N_32948,N_32882);
xor U33057 (N_33057,N_32942,N_32972);
nor U33058 (N_33058,N_32959,N_32976);
xnor U33059 (N_33059,N_32807,N_32971);
nand U33060 (N_33060,N_32852,N_32904);
and U33061 (N_33061,N_32968,N_32927);
xnor U33062 (N_33062,N_32813,N_32809);
nand U33063 (N_33063,N_32938,N_32916);
and U33064 (N_33064,N_32879,N_32836);
xnor U33065 (N_33065,N_32906,N_32876);
and U33066 (N_33066,N_32940,N_32949);
or U33067 (N_33067,N_32980,N_32859);
or U33068 (N_33068,N_32839,N_32984);
and U33069 (N_33069,N_32986,N_32902);
nand U33070 (N_33070,N_32887,N_32862);
and U33071 (N_33071,N_32798,N_32875);
or U33072 (N_33072,N_32955,N_32767);
and U33073 (N_33073,N_32858,N_32977);
or U33074 (N_33074,N_32951,N_32770);
nor U33075 (N_33075,N_32969,N_32827);
and U33076 (N_33076,N_32909,N_32840);
nand U33077 (N_33077,N_32936,N_32752);
xor U33078 (N_33078,N_32919,N_32978);
nor U33079 (N_33079,N_32760,N_32981);
nand U33080 (N_33080,N_32899,N_32990);
and U33081 (N_33081,N_32857,N_32989);
and U33082 (N_33082,N_32946,N_32961);
or U33083 (N_33083,N_32826,N_32866);
nor U33084 (N_33084,N_32816,N_32792);
nand U33085 (N_33085,N_32965,N_32947);
nor U33086 (N_33086,N_32896,N_32954);
nand U33087 (N_33087,N_32762,N_32930);
and U33088 (N_33088,N_32913,N_32994);
nor U33089 (N_33089,N_32829,N_32975);
or U33090 (N_33090,N_32802,N_32960);
xor U33091 (N_33091,N_32825,N_32811);
xor U33092 (N_33092,N_32795,N_32884);
or U33093 (N_33093,N_32849,N_32941);
nand U33094 (N_33094,N_32937,N_32837);
xnor U33095 (N_33095,N_32935,N_32912);
xnor U33096 (N_33096,N_32779,N_32985);
nand U33097 (N_33097,N_32851,N_32890);
or U33098 (N_33098,N_32967,N_32786);
nor U33099 (N_33099,N_32907,N_32903);
xor U33100 (N_33100,N_32877,N_32950);
xnor U33101 (N_33101,N_32863,N_32785);
nor U33102 (N_33102,N_32983,N_32834);
nand U33103 (N_33103,N_32844,N_32761);
nand U33104 (N_33104,N_32808,N_32873);
nor U33105 (N_33105,N_32757,N_32923);
and U33106 (N_33106,N_32824,N_32833);
nand U33107 (N_33107,N_32801,N_32778);
or U33108 (N_33108,N_32797,N_32934);
or U33109 (N_33109,N_32897,N_32820);
nor U33110 (N_33110,N_32939,N_32768);
xnor U33111 (N_33111,N_32774,N_32759);
or U33112 (N_33112,N_32929,N_32910);
nand U33113 (N_33113,N_32842,N_32776);
xor U33114 (N_33114,N_32988,N_32793);
and U33115 (N_33115,N_32979,N_32880);
and U33116 (N_33116,N_32823,N_32766);
nor U33117 (N_33117,N_32900,N_32970);
xnor U33118 (N_33118,N_32931,N_32924);
and U33119 (N_33119,N_32944,N_32956);
xor U33120 (N_33120,N_32991,N_32869);
and U33121 (N_33121,N_32883,N_32780);
xor U33122 (N_33122,N_32838,N_32921);
nor U33123 (N_33123,N_32878,N_32888);
and U33124 (N_33124,N_32993,N_32819);
nor U33125 (N_33125,N_32850,N_32947);
nor U33126 (N_33126,N_32764,N_32768);
and U33127 (N_33127,N_32847,N_32980);
and U33128 (N_33128,N_32963,N_32889);
nand U33129 (N_33129,N_32966,N_32791);
and U33130 (N_33130,N_32897,N_32967);
nand U33131 (N_33131,N_32868,N_32926);
nand U33132 (N_33132,N_32864,N_32898);
nand U33133 (N_33133,N_32901,N_32808);
xnor U33134 (N_33134,N_32904,N_32997);
nor U33135 (N_33135,N_32873,N_32876);
and U33136 (N_33136,N_32765,N_32983);
xor U33137 (N_33137,N_32786,N_32751);
nor U33138 (N_33138,N_32758,N_32825);
nor U33139 (N_33139,N_32968,N_32830);
xnor U33140 (N_33140,N_32864,N_32787);
nand U33141 (N_33141,N_32910,N_32943);
or U33142 (N_33142,N_32946,N_32786);
nand U33143 (N_33143,N_32932,N_32934);
nand U33144 (N_33144,N_32777,N_32947);
nor U33145 (N_33145,N_32886,N_32818);
and U33146 (N_33146,N_32889,N_32986);
nor U33147 (N_33147,N_32967,N_32829);
and U33148 (N_33148,N_32761,N_32885);
nor U33149 (N_33149,N_32836,N_32818);
nand U33150 (N_33150,N_32793,N_32794);
nor U33151 (N_33151,N_32832,N_32816);
nor U33152 (N_33152,N_32844,N_32762);
or U33153 (N_33153,N_32826,N_32778);
xnor U33154 (N_33154,N_32873,N_32778);
nor U33155 (N_33155,N_32868,N_32866);
and U33156 (N_33156,N_32937,N_32874);
nand U33157 (N_33157,N_32780,N_32971);
xnor U33158 (N_33158,N_32778,N_32881);
nor U33159 (N_33159,N_32809,N_32764);
and U33160 (N_33160,N_32770,N_32966);
nor U33161 (N_33161,N_32956,N_32794);
and U33162 (N_33162,N_32843,N_32899);
or U33163 (N_33163,N_32843,N_32824);
nand U33164 (N_33164,N_32878,N_32807);
nor U33165 (N_33165,N_32980,N_32807);
and U33166 (N_33166,N_32786,N_32982);
or U33167 (N_33167,N_32942,N_32878);
and U33168 (N_33168,N_32957,N_32889);
nand U33169 (N_33169,N_32841,N_32899);
nor U33170 (N_33170,N_32936,N_32796);
or U33171 (N_33171,N_32777,N_32849);
xor U33172 (N_33172,N_32987,N_32781);
nor U33173 (N_33173,N_32997,N_32999);
nor U33174 (N_33174,N_32820,N_32867);
nor U33175 (N_33175,N_32804,N_32775);
and U33176 (N_33176,N_32759,N_32756);
and U33177 (N_33177,N_32825,N_32937);
and U33178 (N_33178,N_32947,N_32889);
nand U33179 (N_33179,N_32964,N_32963);
xnor U33180 (N_33180,N_32920,N_32972);
and U33181 (N_33181,N_32988,N_32954);
or U33182 (N_33182,N_32838,N_32967);
or U33183 (N_33183,N_32931,N_32778);
xnor U33184 (N_33184,N_32774,N_32938);
xor U33185 (N_33185,N_32790,N_32758);
nor U33186 (N_33186,N_32798,N_32786);
nor U33187 (N_33187,N_32784,N_32931);
xor U33188 (N_33188,N_32950,N_32816);
nor U33189 (N_33189,N_32981,N_32938);
or U33190 (N_33190,N_32935,N_32987);
and U33191 (N_33191,N_32972,N_32867);
or U33192 (N_33192,N_32915,N_32843);
nand U33193 (N_33193,N_32899,N_32809);
xnor U33194 (N_33194,N_32818,N_32975);
and U33195 (N_33195,N_32823,N_32891);
nand U33196 (N_33196,N_32786,N_32934);
nand U33197 (N_33197,N_32998,N_32885);
or U33198 (N_33198,N_32952,N_32803);
nor U33199 (N_33199,N_32967,N_32869);
and U33200 (N_33200,N_32987,N_32963);
or U33201 (N_33201,N_32864,N_32803);
nor U33202 (N_33202,N_32873,N_32837);
and U33203 (N_33203,N_32791,N_32954);
xnor U33204 (N_33204,N_32862,N_32870);
nor U33205 (N_33205,N_32952,N_32958);
nor U33206 (N_33206,N_32857,N_32892);
xor U33207 (N_33207,N_32812,N_32965);
xnor U33208 (N_33208,N_32834,N_32817);
nor U33209 (N_33209,N_32795,N_32899);
nor U33210 (N_33210,N_32952,N_32904);
or U33211 (N_33211,N_32757,N_32891);
xor U33212 (N_33212,N_32891,N_32927);
and U33213 (N_33213,N_32923,N_32884);
xnor U33214 (N_33214,N_32849,N_32762);
nor U33215 (N_33215,N_32850,N_32839);
and U33216 (N_33216,N_32941,N_32875);
nor U33217 (N_33217,N_32992,N_32946);
nand U33218 (N_33218,N_32936,N_32970);
nor U33219 (N_33219,N_32873,N_32819);
and U33220 (N_33220,N_32889,N_32918);
nand U33221 (N_33221,N_32903,N_32966);
xor U33222 (N_33222,N_32902,N_32841);
nor U33223 (N_33223,N_32780,N_32822);
nor U33224 (N_33224,N_32770,N_32848);
and U33225 (N_33225,N_32823,N_32767);
xor U33226 (N_33226,N_32910,N_32983);
nand U33227 (N_33227,N_32916,N_32805);
xnor U33228 (N_33228,N_32841,N_32766);
and U33229 (N_33229,N_32864,N_32837);
or U33230 (N_33230,N_32768,N_32895);
or U33231 (N_33231,N_32798,N_32792);
or U33232 (N_33232,N_32906,N_32795);
nor U33233 (N_33233,N_32807,N_32989);
nor U33234 (N_33234,N_32884,N_32943);
or U33235 (N_33235,N_32819,N_32870);
nand U33236 (N_33236,N_32969,N_32767);
nand U33237 (N_33237,N_32885,N_32864);
nand U33238 (N_33238,N_32981,N_32752);
and U33239 (N_33239,N_32890,N_32964);
and U33240 (N_33240,N_32907,N_32815);
or U33241 (N_33241,N_32953,N_32753);
and U33242 (N_33242,N_32861,N_32902);
and U33243 (N_33243,N_32982,N_32752);
and U33244 (N_33244,N_32784,N_32980);
or U33245 (N_33245,N_32803,N_32780);
and U33246 (N_33246,N_32880,N_32822);
or U33247 (N_33247,N_32853,N_32902);
nand U33248 (N_33248,N_32932,N_32855);
xor U33249 (N_33249,N_32790,N_32945);
and U33250 (N_33250,N_33220,N_33015);
nand U33251 (N_33251,N_33129,N_33070);
and U33252 (N_33252,N_33026,N_33172);
and U33253 (N_33253,N_33068,N_33152);
nor U33254 (N_33254,N_33155,N_33144);
nand U33255 (N_33255,N_33004,N_33241);
nor U33256 (N_33256,N_33117,N_33197);
or U33257 (N_33257,N_33067,N_33120);
and U33258 (N_33258,N_33227,N_33249);
xor U33259 (N_33259,N_33066,N_33083);
or U33260 (N_33260,N_33166,N_33033);
and U33261 (N_33261,N_33069,N_33239);
xnor U33262 (N_33262,N_33211,N_33053);
nor U33263 (N_33263,N_33058,N_33023);
nand U33264 (N_33264,N_33100,N_33046);
and U33265 (N_33265,N_33128,N_33114);
nand U33266 (N_33266,N_33240,N_33022);
xor U33267 (N_33267,N_33073,N_33086);
nand U33268 (N_33268,N_33064,N_33163);
and U33269 (N_33269,N_33052,N_33008);
and U33270 (N_33270,N_33124,N_33168);
xor U33271 (N_33271,N_33158,N_33138);
and U33272 (N_33272,N_33121,N_33179);
nor U33273 (N_33273,N_33061,N_33057);
and U33274 (N_33274,N_33012,N_33071);
xor U33275 (N_33275,N_33036,N_33130);
xnor U33276 (N_33276,N_33242,N_33159);
and U33277 (N_33277,N_33146,N_33000);
xnor U33278 (N_33278,N_33009,N_33029);
xor U33279 (N_33279,N_33038,N_33021);
or U33280 (N_33280,N_33154,N_33233);
nor U33281 (N_33281,N_33176,N_33207);
and U33282 (N_33282,N_33181,N_33035);
xnor U33283 (N_33283,N_33018,N_33190);
nor U33284 (N_33284,N_33200,N_33082);
nand U33285 (N_33285,N_33056,N_33236);
nand U33286 (N_33286,N_33010,N_33132);
nand U33287 (N_33287,N_33119,N_33123);
xor U33288 (N_33288,N_33189,N_33145);
xor U33289 (N_33289,N_33001,N_33059);
nor U33290 (N_33290,N_33076,N_33054);
nor U33291 (N_33291,N_33186,N_33079);
xor U33292 (N_33292,N_33042,N_33125);
nor U33293 (N_33293,N_33131,N_33014);
or U33294 (N_33294,N_33135,N_33148);
nand U33295 (N_33295,N_33212,N_33112);
nand U33296 (N_33296,N_33103,N_33080);
nand U33297 (N_33297,N_33230,N_33216);
or U33298 (N_33298,N_33013,N_33043);
nand U33299 (N_33299,N_33143,N_33037);
and U33300 (N_33300,N_33045,N_33049);
or U33301 (N_33301,N_33183,N_33185);
xor U33302 (N_33302,N_33111,N_33137);
nand U33303 (N_33303,N_33127,N_33020);
and U33304 (N_33304,N_33167,N_33217);
or U33305 (N_33305,N_33244,N_33027);
nand U33306 (N_33306,N_33208,N_33213);
nand U33307 (N_33307,N_33133,N_33201);
nor U33308 (N_33308,N_33024,N_33170);
nand U33309 (N_33309,N_33002,N_33075);
nand U33310 (N_33310,N_33234,N_33205);
or U33311 (N_33311,N_33175,N_33245);
and U33312 (N_33312,N_33060,N_33174);
nor U33313 (N_33313,N_33202,N_33243);
xnor U33314 (N_33314,N_33184,N_33224);
nand U33315 (N_33315,N_33098,N_33198);
xnor U33316 (N_33316,N_33106,N_33116);
or U33317 (N_33317,N_33169,N_33248);
or U33318 (N_33318,N_33164,N_33044);
nor U33319 (N_33319,N_33084,N_33160);
and U33320 (N_33320,N_33063,N_33085);
nor U33321 (N_33321,N_33161,N_33108);
and U33322 (N_33322,N_33142,N_33007);
and U33323 (N_33323,N_33047,N_33048);
or U33324 (N_33324,N_33065,N_33055);
nor U33325 (N_33325,N_33150,N_33182);
nand U33326 (N_33326,N_33077,N_33187);
nor U33327 (N_33327,N_33147,N_33232);
nor U33328 (N_33328,N_33003,N_33081);
xor U33329 (N_33329,N_33094,N_33203);
nand U33330 (N_33330,N_33221,N_33102);
xnor U33331 (N_33331,N_33034,N_33223);
or U33332 (N_33332,N_33180,N_33199);
xor U33333 (N_33333,N_33193,N_33011);
nor U33334 (N_33334,N_33088,N_33247);
and U33335 (N_33335,N_33099,N_33237);
or U33336 (N_33336,N_33188,N_33210);
nor U33337 (N_33337,N_33177,N_33017);
and U33338 (N_33338,N_33226,N_33238);
and U33339 (N_33339,N_33204,N_33228);
nand U33340 (N_33340,N_33115,N_33196);
nor U33341 (N_33341,N_33156,N_33104);
nor U33342 (N_33342,N_33222,N_33101);
nor U33343 (N_33343,N_33050,N_33157);
nand U33344 (N_33344,N_33136,N_33096);
nand U33345 (N_33345,N_33195,N_33231);
nor U33346 (N_33346,N_33041,N_33074);
or U33347 (N_33347,N_33040,N_33141);
xor U33348 (N_33348,N_33093,N_33235);
nand U33349 (N_33349,N_33118,N_33246);
or U33350 (N_33350,N_33192,N_33215);
nand U33351 (N_33351,N_33051,N_33113);
or U33352 (N_33352,N_33209,N_33090);
nor U33353 (N_33353,N_33091,N_33032);
and U33354 (N_33354,N_33139,N_33219);
nor U33355 (N_33355,N_33153,N_33025);
nand U33356 (N_33356,N_33110,N_33028);
and U33357 (N_33357,N_33092,N_33107);
nor U33358 (N_33358,N_33229,N_33126);
nand U33359 (N_33359,N_33109,N_33095);
and U33360 (N_33360,N_33105,N_33218);
or U33361 (N_33361,N_33122,N_33173);
or U33362 (N_33362,N_33072,N_33149);
nand U33363 (N_33363,N_33162,N_33151);
and U33364 (N_33364,N_33225,N_33171);
nand U33365 (N_33365,N_33006,N_33016);
and U33366 (N_33366,N_33140,N_33087);
xnor U33367 (N_33367,N_33078,N_33062);
nand U33368 (N_33368,N_33194,N_33206);
nor U33369 (N_33369,N_33089,N_33039);
nor U33370 (N_33370,N_33019,N_33031);
nor U33371 (N_33371,N_33030,N_33165);
or U33372 (N_33372,N_33214,N_33134);
nand U33373 (N_33373,N_33005,N_33191);
or U33374 (N_33374,N_33097,N_33178);
xnor U33375 (N_33375,N_33238,N_33148);
or U33376 (N_33376,N_33114,N_33202);
and U33377 (N_33377,N_33100,N_33061);
xor U33378 (N_33378,N_33115,N_33090);
nor U33379 (N_33379,N_33202,N_33197);
xor U33380 (N_33380,N_33093,N_33193);
nor U33381 (N_33381,N_33080,N_33221);
and U33382 (N_33382,N_33023,N_33211);
nor U33383 (N_33383,N_33076,N_33016);
nand U33384 (N_33384,N_33156,N_33217);
nor U33385 (N_33385,N_33219,N_33070);
and U33386 (N_33386,N_33060,N_33036);
or U33387 (N_33387,N_33016,N_33240);
nor U33388 (N_33388,N_33122,N_33159);
nand U33389 (N_33389,N_33066,N_33007);
and U33390 (N_33390,N_33226,N_33177);
or U33391 (N_33391,N_33033,N_33003);
nand U33392 (N_33392,N_33199,N_33005);
or U33393 (N_33393,N_33230,N_33242);
or U33394 (N_33394,N_33162,N_33012);
and U33395 (N_33395,N_33051,N_33091);
and U33396 (N_33396,N_33225,N_33135);
nand U33397 (N_33397,N_33021,N_33127);
nand U33398 (N_33398,N_33158,N_33242);
nand U33399 (N_33399,N_33068,N_33106);
xnor U33400 (N_33400,N_33201,N_33003);
nand U33401 (N_33401,N_33162,N_33216);
and U33402 (N_33402,N_33113,N_33232);
or U33403 (N_33403,N_33087,N_33246);
nor U33404 (N_33404,N_33099,N_33105);
nor U33405 (N_33405,N_33201,N_33011);
or U33406 (N_33406,N_33168,N_33196);
nor U33407 (N_33407,N_33149,N_33245);
and U33408 (N_33408,N_33003,N_33237);
xor U33409 (N_33409,N_33096,N_33135);
and U33410 (N_33410,N_33156,N_33018);
or U33411 (N_33411,N_33230,N_33233);
nor U33412 (N_33412,N_33132,N_33178);
and U33413 (N_33413,N_33146,N_33108);
or U33414 (N_33414,N_33010,N_33121);
nand U33415 (N_33415,N_33019,N_33094);
and U33416 (N_33416,N_33234,N_33088);
or U33417 (N_33417,N_33066,N_33075);
nor U33418 (N_33418,N_33223,N_33095);
and U33419 (N_33419,N_33207,N_33028);
nand U33420 (N_33420,N_33062,N_33040);
xnor U33421 (N_33421,N_33013,N_33049);
nand U33422 (N_33422,N_33210,N_33207);
nand U33423 (N_33423,N_33229,N_33189);
nand U33424 (N_33424,N_33249,N_33005);
or U33425 (N_33425,N_33167,N_33043);
xor U33426 (N_33426,N_33107,N_33133);
or U33427 (N_33427,N_33227,N_33136);
nand U33428 (N_33428,N_33088,N_33239);
or U33429 (N_33429,N_33010,N_33179);
nor U33430 (N_33430,N_33136,N_33052);
and U33431 (N_33431,N_33159,N_33063);
xnor U33432 (N_33432,N_33003,N_33031);
and U33433 (N_33433,N_33230,N_33134);
or U33434 (N_33434,N_33057,N_33178);
xor U33435 (N_33435,N_33161,N_33199);
xor U33436 (N_33436,N_33176,N_33067);
xor U33437 (N_33437,N_33024,N_33076);
nand U33438 (N_33438,N_33161,N_33072);
and U33439 (N_33439,N_33049,N_33204);
or U33440 (N_33440,N_33231,N_33239);
or U33441 (N_33441,N_33168,N_33216);
or U33442 (N_33442,N_33186,N_33102);
nor U33443 (N_33443,N_33115,N_33064);
or U33444 (N_33444,N_33227,N_33082);
or U33445 (N_33445,N_33245,N_33085);
xnor U33446 (N_33446,N_33114,N_33107);
or U33447 (N_33447,N_33224,N_33058);
xor U33448 (N_33448,N_33075,N_33024);
or U33449 (N_33449,N_33241,N_33169);
or U33450 (N_33450,N_33074,N_33005);
xor U33451 (N_33451,N_33106,N_33238);
and U33452 (N_33452,N_33163,N_33221);
xnor U33453 (N_33453,N_33064,N_33036);
nand U33454 (N_33454,N_33146,N_33022);
nor U33455 (N_33455,N_33090,N_33081);
or U33456 (N_33456,N_33110,N_33046);
nand U33457 (N_33457,N_33122,N_33178);
xor U33458 (N_33458,N_33131,N_33072);
xor U33459 (N_33459,N_33023,N_33245);
nor U33460 (N_33460,N_33159,N_33089);
nor U33461 (N_33461,N_33002,N_33058);
and U33462 (N_33462,N_33151,N_33042);
and U33463 (N_33463,N_33037,N_33078);
or U33464 (N_33464,N_33134,N_33002);
and U33465 (N_33465,N_33208,N_33002);
nand U33466 (N_33466,N_33173,N_33228);
or U33467 (N_33467,N_33199,N_33035);
nand U33468 (N_33468,N_33138,N_33153);
nand U33469 (N_33469,N_33126,N_33052);
xor U33470 (N_33470,N_33130,N_33033);
xnor U33471 (N_33471,N_33175,N_33132);
nor U33472 (N_33472,N_33127,N_33067);
or U33473 (N_33473,N_33044,N_33248);
or U33474 (N_33474,N_33076,N_33138);
nand U33475 (N_33475,N_33138,N_33145);
nand U33476 (N_33476,N_33141,N_33052);
and U33477 (N_33477,N_33059,N_33127);
nand U33478 (N_33478,N_33019,N_33248);
or U33479 (N_33479,N_33192,N_33222);
or U33480 (N_33480,N_33023,N_33197);
and U33481 (N_33481,N_33096,N_33062);
nor U33482 (N_33482,N_33174,N_33229);
or U33483 (N_33483,N_33118,N_33068);
nand U33484 (N_33484,N_33140,N_33153);
or U33485 (N_33485,N_33207,N_33165);
xor U33486 (N_33486,N_33129,N_33144);
or U33487 (N_33487,N_33014,N_33071);
xor U33488 (N_33488,N_33243,N_33216);
and U33489 (N_33489,N_33224,N_33091);
and U33490 (N_33490,N_33139,N_33071);
nor U33491 (N_33491,N_33022,N_33041);
nand U33492 (N_33492,N_33019,N_33241);
or U33493 (N_33493,N_33153,N_33018);
nand U33494 (N_33494,N_33092,N_33053);
or U33495 (N_33495,N_33071,N_33241);
and U33496 (N_33496,N_33233,N_33200);
or U33497 (N_33497,N_33216,N_33108);
nor U33498 (N_33498,N_33166,N_33022);
xnor U33499 (N_33499,N_33170,N_33130);
nand U33500 (N_33500,N_33307,N_33329);
and U33501 (N_33501,N_33299,N_33409);
nor U33502 (N_33502,N_33411,N_33331);
xor U33503 (N_33503,N_33278,N_33443);
nand U33504 (N_33504,N_33470,N_33496);
and U33505 (N_33505,N_33358,N_33476);
xor U33506 (N_33506,N_33371,N_33455);
or U33507 (N_33507,N_33494,N_33427);
or U33508 (N_33508,N_33321,N_33268);
nand U33509 (N_33509,N_33316,N_33353);
nor U33510 (N_33510,N_33432,N_33308);
and U33511 (N_33511,N_33349,N_33407);
and U33512 (N_33512,N_33356,N_33343);
nor U33513 (N_33513,N_33254,N_33294);
nand U33514 (N_33514,N_33287,N_33415);
xor U33515 (N_33515,N_33477,N_33489);
xnor U33516 (N_33516,N_33456,N_33383);
xor U33517 (N_33517,N_33313,N_33460);
and U33518 (N_33518,N_33352,N_33304);
xor U33519 (N_33519,N_33255,N_33387);
or U33520 (N_33520,N_33417,N_33271);
nor U33521 (N_33521,N_33341,N_33306);
or U33522 (N_33522,N_33291,N_33499);
xor U33523 (N_33523,N_33333,N_33274);
or U33524 (N_33524,N_33437,N_33327);
nor U33525 (N_33525,N_33478,N_33376);
xor U33526 (N_33526,N_33487,N_33326);
or U33527 (N_33527,N_33257,N_33338);
or U33528 (N_33528,N_33280,N_33282);
nor U33529 (N_33529,N_33416,N_33450);
xnor U33530 (N_33530,N_33467,N_33302);
nor U33531 (N_33531,N_33453,N_33264);
xor U33532 (N_33532,N_33422,N_33441);
or U33533 (N_33533,N_33317,N_33377);
xnor U33534 (N_33534,N_33462,N_33355);
nand U33535 (N_33535,N_33449,N_33429);
or U33536 (N_33536,N_33366,N_33297);
and U33537 (N_33537,N_33335,N_33281);
nor U33538 (N_33538,N_33310,N_33466);
nor U33539 (N_33539,N_33418,N_33479);
xnor U33540 (N_33540,N_33279,N_33347);
or U33541 (N_33541,N_33272,N_33368);
nand U33542 (N_33542,N_33360,N_33348);
nand U33543 (N_33543,N_33433,N_33459);
and U33544 (N_33544,N_33445,N_33448);
nor U33545 (N_33545,N_33270,N_33324);
and U33546 (N_33546,N_33364,N_33414);
nor U33547 (N_33547,N_33398,N_33259);
nor U33548 (N_33548,N_33488,N_33471);
nor U33549 (N_33549,N_33498,N_33258);
or U33550 (N_33550,N_33406,N_33284);
and U33551 (N_33551,N_33252,N_33421);
xor U33552 (N_33552,N_33400,N_33286);
or U33553 (N_33553,N_33266,N_33401);
or U33554 (N_33554,N_33410,N_33357);
or U33555 (N_33555,N_33413,N_33375);
xnor U33556 (N_33556,N_33295,N_33379);
and U33557 (N_33557,N_33388,N_33367);
or U33558 (N_33558,N_33438,N_33277);
nor U33559 (N_33559,N_33293,N_33283);
and U33560 (N_33560,N_33384,N_33262);
or U33561 (N_33561,N_33336,N_33273);
or U33562 (N_33562,N_33276,N_33373);
and U33563 (N_33563,N_33267,N_33454);
nor U33564 (N_33564,N_33396,N_33369);
xnor U33565 (N_33565,N_33346,N_33303);
nor U33566 (N_33566,N_33334,N_33399);
nor U33567 (N_33567,N_33380,N_33391);
xnor U33568 (N_33568,N_33397,N_33473);
xor U33569 (N_33569,N_33469,N_33419);
and U33570 (N_33570,N_33362,N_33440);
xnor U33571 (N_33571,N_33439,N_33318);
nor U33572 (N_33572,N_33285,N_33374);
and U33573 (N_33573,N_33428,N_33394);
and U33574 (N_33574,N_33344,N_33386);
nand U33575 (N_33575,N_33392,N_33385);
nor U33576 (N_33576,N_33461,N_33463);
or U33577 (N_33577,N_33464,N_33492);
and U33578 (N_33578,N_33393,N_33468);
or U33579 (N_33579,N_33482,N_33404);
nand U33580 (N_33580,N_33480,N_33296);
nor U33581 (N_33581,N_33465,N_33350);
xor U33582 (N_33582,N_33430,N_33381);
or U33583 (N_33583,N_33497,N_33351);
xnor U33584 (N_33584,N_33444,N_33265);
nor U33585 (N_33585,N_33378,N_33251);
or U33586 (N_33586,N_33301,N_33442);
nand U33587 (N_33587,N_33314,N_33423);
or U33588 (N_33588,N_33493,N_33484);
or U33589 (N_33589,N_33402,N_33483);
nand U33590 (N_33590,N_33370,N_33345);
nor U33591 (N_33591,N_33485,N_33447);
nor U33592 (N_33592,N_33390,N_33290);
and U33593 (N_33593,N_33474,N_33361);
nor U33594 (N_33594,N_33261,N_33424);
xor U33595 (N_33595,N_33495,N_33395);
nand U33596 (N_33596,N_33315,N_33337);
nor U33597 (N_33597,N_33320,N_33451);
or U33598 (N_33598,N_33405,N_33426);
nor U33599 (N_33599,N_33363,N_33481);
or U33600 (N_33600,N_33305,N_33275);
nand U33601 (N_33601,N_33260,N_33490);
xnor U33602 (N_33602,N_33332,N_33312);
nor U33603 (N_33603,N_33389,N_33269);
nor U33604 (N_33604,N_33298,N_33311);
nor U33605 (N_33605,N_33309,N_33365);
xnor U33606 (N_33606,N_33412,N_33446);
or U33607 (N_33607,N_33452,N_33263);
nor U33608 (N_33608,N_33431,N_33322);
nand U33609 (N_33609,N_33420,N_33475);
or U33610 (N_33610,N_33354,N_33435);
nor U33611 (N_33611,N_33359,N_33330);
and U33612 (N_33612,N_33256,N_33289);
and U33613 (N_33613,N_33403,N_33408);
xnor U33614 (N_33614,N_33436,N_33472);
or U33615 (N_33615,N_33382,N_33339);
or U33616 (N_33616,N_33458,N_33425);
xor U33617 (N_33617,N_33340,N_33434);
or U33618 (N_33618,N_33328,N_33486);
and U33619 (N_33619,N_33457,N_33491);
and U33620 (N_33620,N_33325,N_33323);
and U33621 (N_33621,N_33288,N_33250);
xor U33622 (N_33622,N_33292,N_33342);
and U33623 (N_33623,N_33319,N_33300);
xor U33624 (N_33624,N_33253,N_33372);
nand U33625 (N_33625,N_33373,N_33317);
nand U33626 (N_33626,N_33450,N_33495);
and U33627 (N_33627,N_33488,N_33482);
or U33628 (N_33628,N_33431,N_33303);
or U33629 (N_33629,N_33401,N_33255);
or U33630 (N_33630,N_33418,N_33475);
or U33631 (N_33631,N_33427,N_33387);
nand U33632 (N_33632,N_33495,N_33252);
and U33633 (N_33633,N_33297,N_33428);
nand U33634 (N_33634,N_33313,N_33359);
nand U33635 (N_33635,N_33424,N_33291);
nor U33636 (N_33636,N_33473,N_33321);
xor U33637 (N_33637,N_33277,N_33304);
xnor U33638 (N_33638,N_33482,N_33335);
nor U33639 (N_33639,N_33346,N_33338);
and U33640 (N_33640,N_33414,N_33313);
and U33641 (N_33641,N_33453,N_33351);
nor U33642 (N_33642,N_33312,N_33294);
nor U33643 (N_33643,N_33418,N_33404);
and U33644 (N_33644,N_33371,N_33379);
and U33645 (N_33645,N_33461,N_33303);
and U33646 (N_33646,N_33320,N_33499);
nor U33647 (N_33647,N_33399,N_33305);
and U33648 (N_33648,N_33324,N_33309);
and U33649 (N_33649,N_33317,N_33412);
or U33650 (N_33650,N_33335,N_33254);
nor U33651 (N_33651,N_33263,N_33360);
xnor U33652 (N_33652,N_33455,N_33363);
xnor U33653 (N_33653,N_33283,N_33250);
or U33654 (N_33654,N_33288,N_33477);
and U33655 (N_33655,N_33323,N_33413);
nor U33656 (N_33656,N_33363,N_33365);
nand U33657 (N_33657,N_33344,N_33456);
xnor U33658 (N_33658,N_33381,N_33294);
nand U33659 (N_33659,N_33468,N_33429);
and U33660 (N_33660,N_33448,N_33425);
or U33661 (N_33661,N_33468,N_33254);
nor U33662 (N_33662,N_33448,N_33310);
and U33663 (N_33663,N_33327,N_33400);
nor U33664 (N_33664,N_33291,N_33395);
or U33665 (N_33665,N_33490,N_33285);
nand U33666 (N_33666,N_33458,N_33260);
or U33667 (N_33667,N_33391,N_33255);
xnor U33668 (N_33668,N_33397,N_33474);
nor U33669 (N_33669,N_33460,N_33466);
xor U33670 (N_33670,N_33291,N_33412);
nand U33671 (N_33671,N_33405,N_33470);
xnor U33672 (N_33672,N_33471,N_33325);
nor U33673 (N_33673,N_33297,N_33257);
and U33674 (N_33674,N_33317,N_33358);
or U33675 (N_33675,N_33369,N_33255);
xor U33676 (N_33676,N_33301,N_33483);
nor U33677 (N_33677,N_33376,N_33380);
or U33678 (N_33678,N_33329,N_33469);
or U33679 (N_33679,N_33250,N_33389);
and U33680 (N_33680,N_33477,N_33393);
nand U33681 (N_33681,N_33354,N_33383);
nand U33682 (N_33682,N_33484,N_33401);
nor U33683 (N_33683,N_33351,N_33489);
or U33684 (N_33684,N_33409,N_33382);
nand U33685 (N_33685,N_33288,N_33272);
xnor U33686 (N_33686,N_33306,N_33425);
xor U33687 (N_33687,N_33297,N_33436);
nand U33688 (N_33688,N_33432,N_33410);
nor U33689 (N_33689,N_33292,N_33410);
xor U33690 (N_33690,N_33271,N_33469);
or U33691 (N_33691,N_33326,N_33417);
and U33692 (N_33692,N_33340,N_33321);
and U33693 (N_33693,N_33433,N_33391);
or U33694 (N_33694,N_33279,N_33264);
nor U33695 (N_33695,N_33341,N_33386);
xnor U33696 (N_33696,N_33362,N_33321);
nor U33697 (N_33697,N_33276,N_33366);
nor U33698 (N_33698,N_33426,N_33492);
or U33699 (N_33699,N_33343,N_33424);
nand U33700 (N_33700,N_33298,N_33385);
nor U33701 (N_33701,N_33441,N_33299);
and U33702 (N_33702,N_33468,N_33414);
and U33703 (N_33703,N_33457,N_33311);
or U33704 (N_33704,N_33251,N_33454);
nand U33705 (N_33705,N_33297,N_33291);
nor U33706 (N_33706,N_33449,N_33279);
and U33707 (N_33707,N_33376,N_33290);
xnor U33708 (N_33708,N_33387,N_33335);
nor U33709 (N_33709,N_33340,N_33378);
nor U33710 (N_33710,N_33346,N_33418);
and U33711 (N_33711,N_33278,N_33450);
or U33712 (N_33712,N_33409,N_33350);
and U33713 (N_33713,N_33269,N_33299);
and U33714 (N_33714,N_33398,N_33442);
xnor U33715 (N_33715,N_33370,N_33390);
and U33716 (N_33716,N_33345,N_33346);
nor U33717 (N_33717,N_33426,N_33281);
xnor U33718 (N_33718,N_33462,N_33455);
nor U33719 (N_33719,N_33491,N_33404);
and U33720 (N_33720,N_33346,N_33498);
or U33721 (N_33721,N_33396,N_33453);
xnor U33722 (N_33722,N_33399,N_33446);
nand U33723 (N_33723,N_33256,N_33491);
or U33724 (N_33724,N_33335,N_33498);
nor U33725 (N_33725,N_33365,N_33327);
nor U33726 (N_33726,N_33273,N_33274);
nor U33727 (N_33727,N_33279,N_33328);
nor U33728 (N_33728,N_33389,N_33321);
nand U33729 (N_33729,N_33382,N_33461);
nand U33730 (N_33730,N_33326,N_33373);
nand U33731 (N_33731,N_33409,N_33304);
or U33732 (N_33732,N_33463,N_33476);
nand U33733 (N_33733,N_33385,N_33460);
xnor U33734 (N_33734,N_33320,N_33306);
or U33735 (N_33735,N_33254,N_33330);
nand U33736 (N_33736,N_33334,N_33383);
nor U33737 (N_33737,N_33486,N_33421);
nor U33738 (N_33738,N_33460,N_33495);
and U33739 (N_33739,N_33366,N_33431);
nor U33740 (N_33740,N_33313,N_33415);
nor U33741 (N_33741,N_33375,N_33422);
nor U33742 (N_33742,N_33330,N_33404);
and U33743 (N_33743,N_33455,N_33387);
or U33744 (N_33744,N_33261,N_33442);
nor U33745 (N_33745,N_33397,N_33419);
nor U33746 (N_33746,N_33454,N_33499);
nor U33747 (N_33747,N_33332,N_33474);
xor U33748 (N_33748,N_33264,N_33298);
and U33749 (N_33749,N_33381,N_33299);
nand U33750 (N_33750,N_33610,N_33745);
and U33751 (N_33751,N_33601,N_33617);
or U33752 (N_33752,N_33500,N_33725);
or U33753 (N_33753,N_33523,N_33568);
nand U33754 (N_33754,N_33672,N_33660);
and U33755 (N_33755,N_33653,N_33737);
xor U33756 (N_33756,N_33507,N_33532);
xnor U33757 (N_33757,N_33675,N_33692);
nand U33758 (N_33758,N_33722,N_33713);
or U33759 (N_33759,N_33519,N_33721);
and U33760 (N_33760,N_33749,N_33593);
or U33761 (N_33761,N_33676,N_33540);
xnor U33762 (N_33762,N_33585,N_33548);
nor U33763 (N_33763,N_33586,N_33525);
and U33764 (N_33764,N_33556,N_33543);
and U33765 (N_33765,N_33613,N_33553);
or U33766 (N_33766,N_33592,N_33643);
xnor U33767 (N_33767,N_33572,N_33719);
nand U33768 (N_33768,N_33612,N_33580);
xnor U33769 (N_33769,N_33689,N_33521);
nand U33770 (N_33770,N_33642,N_33697);
nor U33771 (N_33771,N_33724,N_33703);
and U33772 (N_33772,N_33607,N_33618);
xor U33773 (N_33773,N_33638,N_33527);
nand U33774 (N_33774,N_33656,N_33723);
or U33775 (N_33775,N_33736,N_33684);
or U33776 (N_33776,N_33664,N_33545);
nor U33777 (N_33777,N_33668,N_33730);
or U33778 (N_33778,N_33503,N_33663);
and U33779 (N_33779,N_33590,N_33597);
nor U33780 (N_33780,N_33706,N_33620);
nand U33781 (N_33781,N_33558,N_33603);
or U33782 (N_33782,N_33625,N_33515);
and U33783 (N_33783,N_33670,N_33528);
xor U33784 (N_33784,N_33667,N_33526);
and U33785 (N_33785,N_33657,N_33627);
nand U33786 (N_33786,N_33596,N_33655);
and U33787 (N_33787,N_33598,N_33741);
and U33788 (N_33788,N_33662,N_33728);
nor U33789 (N_33789,N_33533,N_33693);
and U33790 (N_33790,N_33536,N_33648);
nor U33791 (N_33791,N_33560,N_33748);
xnor U33792 (N_33792,N_33674,N_33551);
and U33793 (N_33793,N_33554,N_33649);
and U33794 (N_33794,N_33661,N_33566);
nand U33795 (N_33795,N_33567,N_33505);
and U33796 (N_33796,N_33504,N_33608);
nand U33797 (N_33797,N_33632,N_33726);
xnor U33798 (N_33798,N_33744,N_33520);
nand U33799 (N_33799,N_33534,N_33733);
nor U33800 (N_33800,N_33501,N_33575);
nor U33801 (N_33801,N_33633,N_33552);
xor U33802 (N_33802,N_33683,N_33563);
xor U33803 (N_33803,N_33747,N_33579);
xor U33804 (N_33804,N_33509,N_33604);
and U33805 (N_33805,N_33559,N_33619);
or U33806 (N_33806,N_33712,N_33517);
and U33807 (N_33807,N_33637,N_33651);
or U33808 (N_33808,N_33680,N_33530);
and U33809 (N_33809,N_33647,N_33628);
xnor U33810 (N_33810,N_33577,N_33701);
xnor U33811 (N_33811,N_33547,N_33702);
xor U33812 (N_33812,N_33688,N_33666);
and U33813 (N_33813,N_33639,N_33609);
nand U33814 (N_33814,N_33587,N_33738);
nor U33815 (N_33815,N_33705,N_33681);
and U33816 (N_33816,N_33569,N_33582);
and U33817 (N_33817,N_33690,N_33695);
and U33818 (N_33818,N_33731,N_33699);
nand U33819 (N_33819,N_33574,N_33570);
nand U33820 (N_33820,N_33640,N_33518);
xor U33821 (N_33821,N_33600,N_33606);
xnor U33822 (N_33822,N_33658,N_33740);
or U33823 (N_33823,N_33571,N_33623);
nor U33824 (N_33824,N_33615,N_33541);
nand U33825 (N_33825,N_33652,N_33591);
nor U33826 (N_33826,N_33624,N_33546);
and U33827 (N_33827,N_33707,N_33594);
and U33828 (N_33828,N_33709,N_33514);
nor U33829 (N_33829,N_33679,N_33516);
or U33830 (N_33830,N_33644,N_33673);
or U33831 (N_33831,N_33573,N_33614);
and U33832 (N_33832,N_33700,N_33634);
and U33833 (N_33833,N_33659,N_33641);
nor U33834 (N_33834,N_33715,N_33711);
nor U33835 (N_33835,N_33696,N_33734);
or U33836 (N_33836,N_33549,N_33669);
or U33837 (N_33837,N_33529,N_33665);
nand U33838 (N_33838,N_33621,N_33616);
xor U33839 (N_33839,N_33502,N_33589);
and U33840 (N_33840,N_33583,N_33650);
nand U33841 (N_33841,N_33561,N_33704);
nor U33842 (N_33842,N_33602,N_33508);
or U33843 (N_33843,N_33524,N_33510);
xnor U33844 (N_33844,N_33742,N_33513);
xnor U33845 (N_33845,N_33631,N_33544);
nand U33846 (N_33846,N_33605,N_33743);
and U33847 (N_33847,N_33708,N_33645);
nor U33848 (N_33848,N_33710,N_33542);
xnor U33849 (N_33849,N_33646,N_33691);
xor U33850 (N_33850,N_33694,N_33511);
xor U33851 (N_33851,N_33584,N_33562);
nand U33852 (N_33852,N_33739,N_33581);
xor U33853 (N_33853,N_33729,N_33537);
nor U33854 (N_33854,N_33630,N_33718);
xnor U33855 (N_33855,N_33599,N_33538);
and U33856 (N_33856,N_33716,N_33746);
xor U33857 (N_33857,N_33564,N_33682);
and U33858 (N_33858,N_33727,N_33539);
nor U33859 (N_33859,N_33611,N_33636);
and U33860 (N_33860,N_33578,N_33717);
or U33861 (N_33861,N_33735,N_33522);
nand U33862 (N_33862,N_33565,N_33595);
nor U33863 (N_33863,N_33685,N_33576);
xor U33864 (N_33864,N_33622,N_33550);
or U33865 (N_33865,N_33714,N_33686);
nand U33866 (N_33866,N_33588,N_33531);
xnor U33867 (N_33867,N_33678,N_33626);
nor U33868 (N_33868,N_33698,N_33555);
nor U33869 (N_33869,N_33687,N_33720);
or U33870 (N_33870,N_33654,N_33506);
nor U33871 (N_33871,N_33732,N_33629);
and U33872 (N_33872,N_33512,N_33557);
xor U33873 (N_33873,N_33635,N_33535);
xnor U33874 (N_33874,N_33671,N_33677);
and U33875 (N_33875,N_33645,N_33654);
or U33876 (N_33876,N_33634,N_33744);
xnor U33877 (N_33877,N_33574,N_33592);
or U33878 (N_33878,N_33694,N_33608);
or U33879 (N_33879,N_33546,N_33573);
or U33880 (N_33880,N_33667,N_33716);
and U33881 (N_33881,N_33649,N_33683);
xor U33882 (N_33882,N_33735,N_33625);
or U33883 (N_33883,N_33588,N_33563);
nor U33884 (N_33884,N_33516,N_33630);
nor U33885 (N_33885,N_33709,N_33690);
nor U33886 (N_33886,N_33642,N_33723);
and U33887 (N_33887,N_33676,N_33685);
xnor U33888 (N_33888,N_33716,N_33732);
nor U33889 (N_33889,N_33645,N_33734);
nand U33890 (N_33890,N_33521,N_33694);
nand U33891 (N_33891,N_33667,N_33699);
and U33892 (N_33892,N_33507,N_33674);
nor U33893 (N_33893,N_33595,N_33627);
or U33894 (N_33894,N_33732,N_33648);
and U33895 (N_33895,N_33670,N_33728);
nand U33896 (N_33896,N_33606,N_33535);
nand U33897 (N_33897,N_33632,N_33500);
nand U33898 (N_33898,N_33539,N_33682);
nand U33899 (N_33899,N_33713,N_33600);
xnor U33900 (N_33900,N_33522,N_33638);
nor U33901 (N_33901,N_33632,N_33565);
nand U33902 (N_33902,N_33511,N_33576);
nor U33903 (N_33903,N_33610,N_33708);
or U33904 (N_33904,N_33731,N_33630);
and U33905 (N_33905,N_33605,N_33590);
xor U33906 (N_33906,N_33680,N_33738);
nand U33907 (N_33907,N_33727,N_33652);
nor U33908 (N_33908,N_33642,N_33665);
nand U33909 (N_33909,N_33697,N_33537);
nand U33910 (N_33910,N_33547,N_33713);
or U33911 (N_33911,N_33710,N_33733);
nor U33912 (N_33912,N_33600,N_33704);
or U33913 (N_33913,N_33711,N_33639);
nand U33914 (N_33914,N_33545,N_33568);
xnor U33915 (N_33915,N_33558,N_33568);
nor U33916 (N_33916,N_33715,N_33587);
xor U33917 (N_33917,N_33673,N_33572);
nor U33918 (N_33918,N_33572,N_33694);
nor U33919 (N_33919,N_33697,N_33628);
nand U33920 (N_33920,N_33567,N_33562);
and U33921 (N_33921,N_33714,N_33546);
xnor U33922 (N_33922,N_33664,N_33724);
xnor U33923 (N_33923,N_33540,N_33634);
nor U33924 (N_33924,N_33637,N_33504);
nor U33925 (N_33925,N_33699,N_33736);
and U33926 (N_33926,N_33596,N_33563);
nor U33927 (N_33927,N_33694,N_33605);
or U33928 (N_33928,N_33504,N_33635);
xnor U33929 (N_33929,N_33549,N_33539);
nor U33930 (N_33930,N_33523,N_33578);
nor U33931 (N_33931,N_33667,N_33622);
or U33932 (N_33932,N_33588,N_33616);
or U33933 (N_33933,N_33725,N_33648);
or U33934 (N_33934,N_33626,N_33662);
or U33935 (N_33935,N_33585,N_33731);
nand U33936 (N_33936,N_33741,N_33540);
nor U33937 (N_33937,N_33644,N_33603);
or U33938 (N_33938,N_33511,N_33510);
xor U33939 (N_33939,N_33651,N_33669);
nand U33940 (N_33940,N_33673,N_33643);
xnor U33941 (N_33941,N_33537,N_33597);
nand U33942 (N_33942,N_33508,N_33691);
nand U33943 (N_33943,N_33637,N_33587);
nand U33944 (N_33944,N_33630,N_33552);
xnor U33945 (N_33945,N_33693,N_33644);
xnor U33946 (N_33946,N_33590,N_33738);
nand U33947 (N_33947,N_33677,N_33573);
xnor U33948 (N_33948,N_33587,N_33632);
nand U33949 (N_33949,N_33690,N_33716);
and U33950 (N_33950,N_33522,N_33579);
nand U33951 (N_33951,N_33609,N_33585);
nand U33952 (N_33952,N_33617,N_33519);
and U33953 (N_33953,N_33662,N_33606);
nand U33954 (N_33954,N_33590,N_33688);
nor U33955 (N_33955,N_33560,N_33589);
and U33956 (N_33956,N_33540,N_33655);
and U33957 (N_33957,N_33571,N_33671);
xor U33958 (N_33958,N_33746,N_33675);
or U33959 (N_33959,N_33640,N_33679);
nand U33960 (N_33960,N_33517,N_33523);
or U33961 (N_33961,N_33544,N_33716);
nand U33962 (N_33962,N_33524,N_33594);
nand U33963 (N_33963,N_33597,N_33566);
xnor U33964 (N_33964,N_33705,N_33519);
nor U33965 (N_33965,N_33701,N_33576);
or U33966 (N_33966,N_33592,N_33597);
xor U33967 (N_33967,N_33664,N_33610);
nand U33968 (N_33968,N_33746,N_33501);
nand U33969 (N_33969,N_33503,N_33578);
or U33970 (N_33970,N_33520,N_33644);
xor U33971 (N_33971,N_33619,N_33680);
and U33972 (N_33972,N_33653,N_33539);
xnor U33973 (N_33973,N_33555,N_33601);
nand U33974 (N_33974,N_33725,N_33624);
xnor U33975 (N_33975,N_33586,N_33572);
xor U33976 (N_33976,N_33538,N_33676);
nor U33977 (N_33977,N_33562,N_33532);
and U33978 (N_33978,N_33704,N_33544);
or U33979 (N_33979,N_33539,N_33638);
or U33980 (N_33980,N_33582,N_33542);
nor U33981 (N_33981,N_33733,N_33685);
nand U33982 (N_33982,N_33567,N_33725);
nand U33983 (N_33983,N_33699,N_33614);
nand U33984 (N_33984,N_33732,N_33513);
xnor U33985 (N_33985,N_33711,N_33603);
nor U33986 (N_33986,N_33590,N_33593);
xnor U33987 (N_33987,N_33553,N_33575);
nand U33988 (N_33988,N_33671,N_33568);
or U33989 (N_33989,N_33587,N_33579);
nand U33990 (N_33990,N_33744,N_33682);
xor U33991 (N_33991,N_33566,N_33569);
or U33992 (N_33992,N_33562,N_33565);
and U33993 (N_33993,N_33543,N_33590);
nand U33994 (N_33994,N_33500,N_33747);
nor U33995 (N_33995,N_33698,N_33697);
nor U33996 (N_33996,N_33722,N_33665);
nor U33997 (N_33997,N_33586,N_33643);
nor U33998 (N_33998,N_33713,N_33502);
nor U33999 (N_33999,N_33502,N_33570);
xor U34000 (N_34000,N_33768,N_33944);
xor U34001 (N_34001,N_33756,N_33853);
and U34002 (N_34002,N_33986,N_33927);
or U34003 (N_34003,N_33760,N_33793);
and U34004 (N_34004,N_33751,N_33913);
xnor U34005 (N_34005,N_33750,N_33818);
xnor U34006 (N_34006,N_33849,N_33922);
and U34007 (N_34007,N_33786,N_33802);
nor U34008 (N_34008,N_33785,N_33804);
nor U34009 (N_34009,N_33953,N_33891);
nand U34010 (N_34010,N_33884,N_33993);
nand U34011 (N_34011,N_33822,N_33905);
and U34012 (N_34012,N_33771,N_33835);
xor U34013 (N_34013,N_33803,N_33916);
xor U34014 (N_34014,N_33873,N_33964);
or U34015 (N_34015,N_33865,N_33954);
nand U34016 (N_34016,N_33859,N_33805);
nand U34017 (N_34017,N_33808,N_33777);
nor U34018 (N_34018,N_33758,N_33992);
nand U34019 (N_34019,N_33796,N_33856);
or U34020 (N_34020,N_33995,N_33938);
xor U34021 (N_34021,N_33860,N_33962);
and U34022 (N_34022,N_33904,N_33985);
nor U34023 (N_34023,N_33979,N_33915);
or U34024 (N_34024,N_33893,N_33923);
nand U34025 (N_34025,N_33861,N_33824);
and U34026 (N_34026,N_33975,N_33817);
or U34027 (N_34027,N_33929,N_33752);
xnor U34028 (N_34028,N_33984,N_33887);
or U34029 (N_34029,N_33779,N_33902);
xor U34030 (N_34030,N_33882,N_33982);
and U34031 (N_34031,N_33857,N_33945);
nor U34032 (N_34032,N_33978,N_33754);
or U34033 (N_34033,N_33942,N_33903);
and U34034 (N_34034,N_33762,N_33920);
xnor U34035 (N_34035,N_33811,N_33981);
and U34036 (N_34036,N_33968,N_33937);
nand U34037 (N_34037,N_33926,N_33901);
nor U34038 (N_34038,N_33976,N_33827);
xor U34039 (N_34039,N_33838,N_33991);
or U34040 (N_34040,N_33983,N_33814);
nor U34041 (N_34041,N_33775,N_33888);
nor U34042 (N_34042,N_33850,N_33950);
nor U34043 (N_34043,N_33876,N_33909);
or U34044 (N_34044,N_33969,N_33897);
nor U34045 (N_34045,N_33855,N_33878);
nand U34046 (N_34046,N_33911,N_33772);
nand U34047 (N_34047,N_33840,N_33987);
nor U34048 (N_34048,N_33990,N_33880);
nand U34049 (N_34049,N_33858,N_33948);
xor U34050 (N_34050,N_33932,N_33947);
nor U34051 (N_34051,N_33955,N_33765);
or U34052 (N_34052,N_33966,N_33815);
xnor U34053 (N_34053,N_33764,N_33820);
xnor U34054 (N_34054,N_33924,N_33939);
xor U34055 (N_34055,N_33801,N_33997);
nor U34056 (N_34056,N_33946,N_33914);
or U34057 (N_34057,N_33892,N_33951);
xnor U34058 (N_34058,N_33843,N_33918);
and U34059 (N_34059,N_33896,N_33836);
nand U34060 (N_34060,N_33988,N_33797);
or U34061 (N_34061,N_33770,N_33807);
and U34062 (N_34062,N_33883,N_33753);
xnor U34063 (N_34063,N_33907,N_33956);
nor U34064 (N_34064,N_33921,N_33973);
nor U34065 (N_34065,N_33959,N_33763);
and U34066 (N_34066,N_33931,N_33800);
xnor U34067 (N_34067,N_33996,N_33999);
and U34068 (N_34068,N_33841,N_33940);
nor U34069 (N_34069,N_33839,N_33972);
and U34070 (N_34070,N_33898,N_33813);
nor U34071 (N_34071,N_33848,N_33980);
and U34072 (N_34072,N_33812,N_33773);
nand U34073 (N_34073,N_33952,N_33766);
nand U34074 (N_34074,N_33780,N_33790);
or U34075 (N_34075,N_33906,N_33963);
and U34076 (N_34076,N_33894,N_33816);
nor U34077 (N_34077,N_33837,N_33810);
nor U34078 (N_34078,N_33871,N_33847);
or U34079 (N_34079,N_33957,N_33788);
nand U34080 (N_34080,N_33776,N_33823);
nor U34081 (N_34081,N_33899,N_33792);
nand U34082 (N_34082,N_33821,N_33833);
and U34083 (N_34083,N_33829,N_33787);
xor U34084 (N_34084,N_33806,N_33809);
and U34085 (N_34085,N_33885,N_33778);
nor U34086 (N_34086,N_33872,N_33879);
nor U34087 (N_34087,N_33933,N_33890);
nand U34088 (N_34088,N_33757,N_33769);
and U34089 (N_34089,N_33934,N_33834);
nand U34090 (N_34090,N_33774,N_33895);
nand U34091 (N_34091,N_33935,N_33900);
or U34092 (N_34092,N_33886,N_33917);
nand U34093 (N_34093,N_33869,N_33974);
and U34094 (N_34094,N_33994,N_33759);
or U34095 (N_34095,N_33862,N_33881);
nor U34096 (N_34096,N_33889,N_33989);
and U34097 (N_34097,N_33870,N_33867);
xor U34098 (N_34098,N_33791,N_33863);
xnor U34099 (N_34099,N_33961,N_33761);
and U34100 (N_34100,N_33874,N_33868);
nand U34101 (N_34101,N_33798,N_33844);
or U34102 (N_34102,N_33908,N_33970);
and U34103 (N_34103,N_33819,N_33910);
xor U34104 (N_34104,N_33767,N_33925);
xnor U34105 (N_34105,N_33795,N_33936);
xor U34106 (N_34106,N_33877,N_33875);
nor U34107 (N_34107,N_33799,N_33977);
xnor U34108 (N_34108,N_33864,N_33971);
nor U34109 (N_34109,N_33943,N_33912);
nor U34110 (N_34110,N_33852,N_33941);
and U34111 (N_34111,N_33866,N_33854);
nor U34112 (N_34112,N_33825,N_33781);
nor U34113 (N_34113,N_33830,N_33832);
nand U34114 (N_34114,N_33783,N_33794);
and U34115 (N_34115,N_33755,N_33998);
xor U34116 (N_34116,N_33846,N_33782);
or U34117 (N_34117,N_33826,N_33928);
nor U34118 (N_34118,N_33919,N_33845);
xnor U34119 (N_34119,N_33789,N_33842);
and U34120 (N_34120,N_33967,N_33831);
and U34121 (N_34121,N_33828,N_33851);
xnor U34122 (N_34122,N_33930,N_33949);
nand U34123 (N_34123,N_33958,N_33784);
and U34124 (N_34124,N_33960,N_33965);
and U34125 (N_34125,N_33841,N_33835);
xor U34126 (N_34126,N_33923,N_33777);
nor U34127 (N_34127,N_33870,N_33901);
nand U34128 (N_34128,N_33818,N_33836);
or U34129 (N_34129,N_33937,N_33909);
nand U34130 (N_34130,N_33939,N_33880);
and U34131 (N_34131,N_33768,N_33764);
nor U34132 (N_34132,N_33994,N_33921);
nand U34133 (N_34133,N_33957,N_33828);
and U34134 (N_34134,N_33902,N_33966);
nand U34135 (N_34135,N_33946,N_33891);
nand U34136 (N_34136,N_33813,N_33965);
nand U34137 (N_34137,N_33827,N_33778);
or U34138 (N_34138,N_33866,N_33761);
nor U34139 (N_34139,N_33801,N_33967);
xor U34140 (N_34140,N_33927,N_33903);
and U34141 (N_34141,N_33873,N_33775);
and U34142 (N_34142,N_33984,N_33823);
and U34143 (N_34143,N_33862,N_33939);
and U34144 (N_34144,N_33971,N_33914);
or U34145 (N_34145,N_33887,N_33794);
nand U34146 (N_34146,N_33945,N_33765);
or U34147 (N_34147,N_33844,N_33758);
xor U34148 (N_34148,N_33887,N_33817);
nand U34149 (N_34149,N_33952,N_33885);
and U34150 (N_34150,N_33867,N_33806);
nor U34151 (N_34151,N_33886,N_33754);
xnor U34152 (N_34152,N_33751,N_33840);
and U34153 (N_34153,N_33921,N_33862);
and U34154 (N_34154,N_33948,N_33951);
nand U34155 (N_34155,N_33884,N_33823);
and U34156 (N_34156,N_33994,N_33791);
nand U34157 (N_34157,N_33925,N_33977);
and U34158 (N_34158,N_33948,N_33792);
nand U34159 (N_34159,N_33843,N_33855);
nand U34160 (N_34160,N_33936,N_33935);
nand U34161 (N_34161,N_33837,N_33787);
or U34162 (N_34162,N_33891,N_33999);
nand U34163 (N_34163,N_33951,N_33779);
xor U34164 (N_34164,N_33802,N_33840);
nand U34165 (N_34165,N_33861,N_33905);
nand U34166 (N_34166,N_33879,N_33976);
or U34167 (N_34167,N_33928,N_33948);
or U34168 (N_34168,N_33966,N_33961);
xor U34169 (N_34169,N_33955,N_33811);
or U34170 (N_34170,N_33801,N_33963);
xnor U34171 (N_34171,N_33852,N_33905);
or U34172 (N_34172,N_33988,N_33855);
nor U34173 (N_34173,N_33787,N_33970);
xor U34174 (N_34174,N_33757,N_33965);
or U34175 (N_34175,N_33953,N_33990);
xnor U34176 (N_34176,N_33936,N_33760);
and U34177 (N_34177,N_33825,N_33879);
xnor U34178 (N_34178,N_33815,N_33808);
and U34179 (N_34179,N_33796,N_33942);
nor U34180 (N_34180,N_33909,N_33960);
or U34181 (N_34181,N_33902,N_33810);
or U34182 (N_34182,N_33957,N_33875);
nand U34183 (N_34183,N_33833,N_33849);
nor U34184 (N_34184,N_33988,N_33925);
nor U34185 (N_34185,N_33839,N_33907);
nand U34186 (N_34186,N_33951,N_33826);
or U34187 (N_34187,N_33845,N_33819);
or U34188 (N_34188,N_33750,N_33875);
nand U34189 (N_34189,N_33855,N_33924);
and U34190 (N_34190,N_33828,N_33789);
nand U34191 (N_34191,N_33942,N_33990);
or U34192 (N_34192,N_33807,N_33829);
and U34193 (N_34193,N_33926,N_33945);
or U34194 (N_34194,N_33977,N_33897);
or U34195 (N_34195,N_33945,N_33804);
nand U34196 (N_34196,N_33849,N_33800);
nor U34197 (N_34197,N_33753,N_33940);
xnor U34198 (N_34198,N_33869,N_33898);
nor U34199 (N_34199,N_33827,N_33899);
and U34200 (N_34200,N_33952,N_33765);
and U34201 (N_34201,N_33823,N_33946);
nand U34202 (N_34202,N_33977,N_33774);
xor U34203 (N_34203,N_33929,N_33842);
xor U34204 (N_34204,N_33931,N_33954);
nor U34205 (N_34205,N_33867,N_33979);
xor U34206 (N_34206,N_33890,N_33926);
or U34207 (N_34207,N_33763,N_33871);
xor U34208 (N_34208,N_33942,N_33914);
and U34209 (N_34209,N_33989,N_33847);
and U34210 (N_34210,N_33998,N_33885);
nor U34211 (N_34211,N_33950,N_33765);
or U34212 (N_34212,N_33981,N_33827);
or U34213 (N_34213,N_33918,N_33920);
xor U34214 (N_34214,N_33852,N_33798);
nor U34215 (N_34215,N_33998,N_33784);
nand U34216 (N_34216,N_33959,N_33817);
or U34217 (N_34217,N_33788,N_33763);
nand U34218 (N_34218,N_33752,N_33982);
nor U34219 (N_34219,N_33870,N_33779);
and U34220 (N_34220,N_33807,N_33964);
xnor U34221 (N_34221,N_33914,N_33929);
xor U34222 (N_34222,N_33774,N_33998);
nand U34223 (N_34223,N_33913,N_33821);
or U34224 (N_34224,N_33968,N_33796);
nor U34225 (N_34225,N_33952,N_33974);
and U34226 (N_34226,N_33979,N_33762);
and U34227 (N_34227,N_33814,N_33785);
and U34228 (N_34228,N_33888,N_33904);
and U34229 (N_34229,N_33843,N_33964);
and U34230 (N_34230,N_33960,N_33941);
xnor U34231 (N_34231,N_33853,N_33979);
or U34232 (N_34232,N_33844,N_33871);
nand U34233 (N_34233,N_33967,N_33804);
nand U34234 (N_34234,N_33791,N_33839);
and U34235 (N_34235,N_33957,N_33765);
nor U34236 (N_34236,N_33944,N_33974);
or U34237 (N_34237,N_33912,N_33881);
xnor U34238 (N_34238,N_33982,N_33896);
or U34239 (N_34239,N_33773,N_33976);
nand U34240 (N_34240,N_33867,N_33967);
or U34241 (N_34241,N_33984,N_33755);
nand U34242 (N_34242,N_33930,N_33926);
and U34243 (N_34243,N_33942,N_33895);
nand U34244 (N_34244,N_33929,N_33801);
or U34245 (N_34245,N_33945,N_33808);
nand U34246 (N_34246,N_33857,N_33776);
or U34247 (N_34247,N_33942,N_33776);
and U34248 (N_34248,N_33754,N_33891);
nor U34249 (N_34249,N_33751,N_33903);
xnor U34250 (N_34250,N_34198,N_34044);
nor U34251 (N_34251,N_34134,N_34187);
nand U34252 (N_34252,N_34233,N_34113);
or U34253 (N_34253,N_34138,N_34118);
nand U34254 (N_34254,N_34078,N_34057);
and U34255 (N_34255,N_34099,N_34071);
nand U34256 (N_34256,N_34043,N_34175);
xnor U34257 (N_34257,N_34114,N_34086);
or U34258 (N_34258,N_34238,N_34201);
and U34259 (N_34259,N_34240,N_34056);
or U34260 (N_34260,N_34145,N_34003);
xnor U34261 (N_34261,N_34096,N_34139);
nand U34262 (N_34262,N_34136,N_34149);
nor U34263 (N_34263,N_34017,N_34102);
nor U34264 (N_34264,N_34068,N_34129);
xnor U34265 (N_34265,N_34235,N_34179);
xnor U34266 (N_34266,N_34019,N_34212);
xnor U34267 (N_34267,N_34048,N_34074);
xor U34268 (N_34268,N_34177,N_34084);
nor U34269 (N_34269,N_34182,N_34122);
xor U34270 (N_34270,N_34224,N_34242);
nand U34271 (N_34271,N_34217,N_34010);
xnor U34272 (N_34272,N_34152,N_34249);
xor U34273 (N_34273,N_34008,N_34091);
nand U34274 (N_34274,N_34246,N_34062);
xnor U34275 (N_34275,N_34181,N_34028);
xnor U34276 (N_34276,N_34237,N_34137);
nor U34277 (N_34277,N_34222,N_34047);
xor U34278 (N_34278,N_34040,N_34070);
nor U34279 (N_34279,N_34117,N_34041);
nor U34280 (N_34280,N_34075,N_34241);
or U34281 (N_34281,N_34190,N_34006);
xor U34282 (N_34282,N_34020,N_34061);
or U34283 (N_34283,N_34065,N_34083);
nand U34284 (N_34284,N_34239,N_34215);
nand U34285 (N_34285,N_34077,N_34227);
xnor U34286 (N_34286,N_34150,N_34144);
and U34287 (N_34287,N_34130,N_34104);
or U34288 (N_34288,N_34123,N_34112);
and U34289 (N_34289,N_34169,N_34206);
nor U34290 (N_34290,N_34115,N_34004);
and U34291 (N_34291,N_34024,N_34166);
nor U34292 (N_34292,N_34165,N_34023);
and U34293 (N_34293,N_34053,N_34002);
and U34294 (N_34294,N_34103,N_34033);
and U34295 (N_34295,N_34140,N_34230);
xor U34296 (N_34296,N_34058,N_34178);
xor U34297 (N_34297,N_34200,N_34049);
or U34298 (N_34298,N_34111,N_34228);
xnor U34299 (N_34299,N_34073,N_34219);
nand U34300 (N_34300,N_34066,N_34045);
or U34301 (N_34301,N_34171,N_34121);
and U34302 (N_34302,N_34155,N_34089);
or U34303 (N_34303,N_34176,N_34164);
and U34304 (N_34304,N_34243,N_34097);
or U34305 (N_34305,N_34059,N_34054);
nor U34306 (N_34306,N_34223,N_34157);
and U34307 (N_34307,N_34159,N_34210);
and U34308 (N_34308,N_34080,N_34147);
nand U34309 (N_34309,N_34030,N_34093);
nand U34310 (N_34310,N_34188,N_34052);
xor U34311 (N_34311,N_34192,N_34090);
xor U34312 (N_34312,N_34076,N_34209);
or U34313 (N_34313,N_34234,N_34055);
nand U34314 (N_34314,N_34214,N_34173);
nand U34315 (N_34315,N_34088,N_34193);
or U34316 (N_34316,N_34127,N_34146);
xor U34317 (N_34317,N_34029,N_34162);
nor U34318 (N_34318,N_34027,N_34072);
nor U34319 (N_34319,N_34189,N_34244);
nand U34320 (N_34320,N_34092,N_34202);
or U34321 (N_34321,N_34079,N_34016);
or U34322 (N_34322,N_34185,N_34095);
xor U34323 (N_34323,N_34110,N_34225);
nand U34324 (N_34324,N_34180,N_34194);
or U34325 (N_34325,N_34184,N_34207);
nor U34326 (N_34326,N_34142,N_34131);
nor U34327 (N_34327,N_34218,N_34100);
nand U34328 (N_34328,N_34160,N_34120);
or U34329 (N_34329,N_34015,N_34151);
or U34330 (N_34330,N_34183,N_34216);
xor U34331 (N_34331,N_34213,N_34000);
nand U34332 (N_34332,N_34018,N_34153);
or U34333 (N_34333,N_34126,N_34148);
or U34334 (N_34334,N_34063,N_34098);
nand U34335 (N_34335,N_34101,N_34132);
xnor U34336 (N_34336,N_34128,N_34005);
nor U34337 (N_34337,N_34143,N_34022);
xor U34338 (N_34338,N_34032,N_34245);
or U34339 (N_34339,N_34087,N_34085);
xnor U34340 (N_34340,N_34026,N_34141);
xor U34341 (N_34341,N_34031,N_34221);
nand U34342 (N_34342,N_34034,N_34226);
xor U34343 (N_34343,N_34025,N_34236);
xor U34344 (N_34344,N_34174,N_34211);
xor U34345 (N_34345,N_34081,N_34011);
and U34346 (N_34346,N_34229,N_34037);
nor U34347 (N_34347,N_34196,N_34069);
nor U34348 (N_34348,N_34163,N_34197);
xnor U34349 (N_34349,N_34124,N_34248);
or U34350 (N_34350,N_34105,N_34231);
nand U34351 (N_34351,N_34001,N_34007);
and U34352 (N_34352,N_34108,N_34186);
and U34353 (N_34353,N_34154,N_34067);
or U34354 (N_34354,N_34060,N_34051);
nand U34355 (N_34355,N_34082,N_34014);
nand U34356 (N_34356,N_34161,N_34168);
nand U34357 (N_34357,N_34042,N_34247);
nor U34358 (N_34358,N_34107,N_34050);
nor U34359 (N_34359,N_34125,N_34013);
nand U34360 (N_34360,N_34036,N_34172);
xnor U34361 (N_34361,N_34094,N_34039);
nand U34362 (N_34362,N_34009,N_34133);
or U34363 (N_34363,N_34208,N_34135);
nand U34364 (N_34364,N_34203,N_34156);
nand U34365 (N_34365,N_34064,N_34038);
or U34366 (N_34366,N_34035,N_34232);
nor U34367 (N_34367,N_34167,N_34046);
and U34368 (N_34368,N_34170,N_34195);
nand U34369 (N_34369,N_34012,N_34116);
and U34370 (N_34370,N_34119,N_34199);
nor U34371 (N_34371,N_34220,N_34204);
nor U34372 (N_34372,N_34109,N_34021);
or U34373 (N_34373,N_34191,N_34158);
or U34374 (N_34374,N_34205,N_34106);
nand U34375 (N_34375,N_34139,N_34243);
nor U34376 (N_34376,N_34181,N_34147);
or U34377 (N_34377,N_34223,N_34243);
nor U34378 (N_34378,N_34242,N_34178);
and U34379 (N_34379,N_34177,N_34212);
nor U34380 (N_34380,N_34218,N_34224);
nand U34381 (N_34381,N_34139,N_34195);
nor U34382 (N_34382,N_34229,N_34022);
xnor U34383 (N_34383,N_34120,N_34005);
xor U34384 (N_34384,N_34084,N_34105);
nor U34385 (N_34385,N_34110,N_34074);
nand U34386 (N_34386,N_34016,N_34113);
or U34387 (N_34387,N_34243,N_34132);
xnor U34388 (N_34388,N_34034,N_34198);
nand U34389 (N_34389,N_34078,N_34003);
nand U34390 (N_34390,N_34235,N_34212);
or U34391 (N_34391,N_34146,N_34006);
and U34392 (N_34392,N_34014,N_34208);
nand U34393 (N_34393,N_34038,N_34195);
xnor U34394 (N_34394,N_34117,N_34089);
nor U34395 (N_34395,N_34090,N_34145);
or U34396 (N_34396,N_34107,N_34141);
xor U34397 (N_34397,N_34107,N_34065);
nor U34398 (N_34398,N_34106,N_34211);
nor U34399 (N_34399,N_34154,N_34049);
nand U34400 (N_34400,N_34057,N_34023);
nor U34401 (N_34401,N_34102,N_34088);
or U34402 (N_34402,N_34124,N_34227);
nand U34403 (N_34403,N_34190,N_34045);
or U34404 (N_34404,N_34029,N_34158);
xnor U34405 (N_34405,N_34144,N_34201);
nor U34406 (N_34406,N_34034,N_34174);
nand U34407 (N_34407,N_34196,N_34052);
xnor U34408 (N_34408,N_34052,N_34099);
nor U34409 (N_34409,N_34210,N_34208);
nor U34410 (N_34410,N_34050,N_34183);
nand U34411 (N_34411,N_34111,N_34056);
nand U34412 (N_34412,N_34225,N_34050);
and U34413 (N_34413,N_34188,N_34058);
nor U34414 (N_34414,N_34222,N_34086);
or U34415 (N_34415,N_34176,N_34064);
nor U34416 (N_34416,N_34246,N_34061);
nand U34417 (N_34417,N_34114,N_34079);
and U34418 (N_34418,N_34169,N_34002);
or U34419 (N_34419,N_34035,N_34103);
and U34420 (N_34420,N_34189,N_34185);
nand U34421 (N_34421,N_34126,N_34177);
xnor U34422 (N_34422,N_34183,N_34213);
and U34423 (N_34423,N_34013,N_34149);
and U34424 (N_34424,N_34044,N_34213);
and U34425 (N_34425,N_34021,N_34036);
or U34426 (N_34426,N_34175,N_34077);
xor U34427 (N_34427,N_34160,N_34084);
or U34428 (N_34428,N_34110,N_34019);
nor U34429 (N_34429,N_34111,N_34030);
xnor U34430 (N_34430,N_34025,N_34011);
and U34431 (N_34431,N_34127,N_34094);
xnor U34432 (N_34432,N_34167,N_34094);
nor U34433 (N_34433,N_34172,N_34140);
nor U34434 (N_34434,N_34172,N_34086);
or U34435 (N_34435,N_34012,N_34112);
or U34436 (N_34436,N_34158,N_34101);
xnor U34437 (N_34437,N_34105,N_34242);
and U34438 (N_34438,N_34184,N_34092);
nor U34439 (N_34439,N_34025,N_34074);
xor U34440 (N_34440,N_34212,N_34154);
and U34441 (N_34441,N_34228,N_34119);
and U34442 (N_34442,N_34170,N_34232);
xor U34443 (N_34443,N_34148,N_34230);
or U34444 (N_34444,N_34175,N_34060);
nand U34445 (N_34445,N_34205,N_34244);
nor U34446 (N_34446,N_34090,N_34212);
and U34447 (N_34447,N_34168,N_34055);
nand U34448 (N_34448,N_34064,N_34207);
or U34449 (N_34449,N_34192,N_34067);
nor U34450 (N_34450,N_34120,N_34041);
or U34451 (N_34451,N_34128,N_34241);
xor U34452 (N_34452,N_34219,N_34124);
xor U34453 (N_34453,N_34240,N_34219);
and U34454 (N_34454,N_34083,N_34214);
and U34455 (N_34455,N_34216,N_34074);
or U34456 (N_34456,N_34085,N_34028);
nand U34457 (N_34457,N_34074,N_34242);
and U34458 (N_34458,N_34112,N_34195);
nor U34459 (N_34459,N_34021,N_34153);
xnor U34460 (N_34460,N_34200,N_34022);
nor U34461 (N_34461,N_34075,N_34103);
and U34462 (N_34462,N_34114,N_34228);
and U34463 (N_34463,N_34244,N_34179);
nor U34464 (N_34464,N_34077,N_34068);
or U34465 (N_34465,N_34158,N_34086);
nor U34466 (N_34466,N_34087,N_34015);
xor U34467 (N_34467,N_34144,N_34139);
xor U34468 (N_34468,N_34168,N_34144);
or U34469 (N_34469,N_34041,N_34089);
nor U34470 (N_34470,N_34042,N_34018);
nor U34471 (N_34471,N_34189,N_34091);
or U34472 (N_34472,N_34220,N_34203);
nand U34473 (N_34473,N_34016,N_34025);
nand U34474 (N_34474,N_34032,N_34086);
or U34475 (N_34475,N_34208,N_34180);
nor U34476 (N_34476,N_34092,N_34199);
nand U34477 (N_34477,N_34239,N_34136);
or U34478 (N_34478,N_34000,N_34185);
nand U34479 (N_34479,N_34169,N_34070);
xnor U34480 (N_34480,N_34181,N_34043);
nor U34481 (N_34481,N_34115,N_34185);
nor U34482 (N_34482,N_34054,N_34199);
and U34483 (N_34483,N_34105,N_34158);
nor U34484 (N_34484,N_34023,N_34207);
and U34485 (N_34485,N_34059,N_34239);
or U34486 (N_34486,N_34087,N_34221);
nand U34487 (N_34487,N_34242,N_34039);
and U34488 (N_34488,N_34148,N_34249);
nand U34489 (N_34489,N_34004,N_34207);
nand U34490 (N_34490,N_34216,N_34147);
nor U34491 (N_34491,N_34072,N_34144);
xor U34492 (N_34492,N_34016,N_34067);
or U34493 (N_34493,N_34047,N_34203);
and U34494 (N_34494,N_34037,N_34126);
nor U34495 (N_34495,N_34029,N_34163);
or U34496 (N_34496,N_34091,N_34211);
nand U34497 (N_34497,N_34087,N_34092);
and U34498 (N_34498,N_34008,N_34162);
nand U34499 (N_34499,N_34089,N_34227);
nor U34500 (N_34500,N_34268,N_34289);
xor U34501 (N_34501,N_34489,N_34362);
nor U34502 (N_34502,N_34294,N_34275);
xor U34503 (N_34503,N_34363,N_34478);
xor U34504 (N_34504,N_34364,N_34269);
or U34505 (N_34505,N_34428,N_34284);
nor U34506 (N_34506,N_34400,N_34256);
or U34507 (N_34507,N_34344,N_34448);
nand U34508 (N_34508,N_34437,N_34305);
or U34509 (N_34509,N_34271,N_34323);
nand U34510 (N_34510,N_34393,N_34450);
nand U34511 (N_34511,N_34250,N_34286);
nand U34512 (N_34512,N_34471,N_34310);
nand U34513 (N_34513,N_34388,N_34343);
and U34514 (N_34514,N_34272,N_34409);
nor U34515 (N_34515,N_34464,N_34446);
nand U34516 (N_34516,N_34261,N_34325);
nor U34517 (N_34517,N_34341,N_34487);
xor U34518 (N_34518,N_34259,N_34380);
or U34519 (N_34519,N_34290,N_34279);
or U34520 (N_34520,N_34273,N_34350);
xnor U34521 (N_34521,N_34386,N_34408);
xor U34522 (N_34522,N_34338,N_34353);
nand U34523 (N_34523,N_34327,N_34361);
nor U34524 (N_34524,N_34413,N_34266);
nand U34525 (N_34525,N_34307,N_34451);
and U34526 (N_34526,N_34333,N_34348);
xnor U34527 (N_34527,N_34398,N_34382);
and U34528 (N_34528,N_34420,N_34383);
or U34529 (N_34529,N_34312,N_34292);
nor U34530 (N_34530,N_34476,N_34372);
or U34531 (N_34531,N_34337,N_34480);
and U34532 (N_34532,N_34440,N_34472);
xor U34533 (N_34533,N_34295,N_34412);
and U34534 (N_34534,N_34457,N_34314);
xnor U34535 (N_34535,N_34373,N_34481);
nand U34536 (N_34536,N_34418,N_34411);
or U34537 (N_34537,N_34298,N_34479);
or U34538 (N_34538,N_34253,N_34278);
or U34539 (N_34539,N_34465,N_34477);
or U34540 (N_34540,N_34374,N_34391);
or U34541 (N_34541,N_34425,N_34280);
xor U34542 (N_34542,N_34475,N_34387);
nand U34543 (N_34543,N_34316,N_34311);
and U34544 (N_34544,N_34324,N_34328);
nand U34545 (N_34545,N_34433,N_34300);
nor U34546 (N_34546,N_34330,N_34376);
xnor U34547 (N_34547,N_34329,N_34371);
nor U34548 (N_34548,N_34454,N_34389);
xor U34549 (N_34549,N_34319,N_34375);
xnor U34550 (N_34550,N_34499,N_34392);
nand U34551 (N_34551,N_34442,N_34384);
xor U34552 (N_34552,N_34331,N_34491);
nand U34553 (N_34553,N_34474,N_34493);
xor U34554 (N_34554,N_34320,N_34262);
nand U34555 (N_34555,N_34449,N_34459);
or U34556 (N_34556,N_34385,N_34297);
and U34557 (N_34557,N_34417,N_34264);
nand U34558 (N_34558,N_34378,N_34470);
nand U34559 (N_34559,N_34357,N_34463);
or U34560 (N_34560,N_34263,N_34497);
nand U34561 (N_34561,N_34274,N_34365);
nand U34562 (N_34562,N_34293,N_34315);
nand U34563 (N_34563,N_34435,N_34347);
xor U34564 (N_34564,N_34453,N_34462);
or U34565 (N_34565,N_34354,N_34434);
xor U34566 (N_34566,N_34429,N_34441);
xor U34567 (N_34567,N_34490,N_34318);
nor U34568 (N_34568,N_34469,N_34349);
nand U34569 (N_34569,N_34445,N_34415);
nor U34570 (N_34570,N_34456,N_34317);
xor U34571 (N_34571,N_34302,N_34460);
xor U34572 (N_34572,N_34342,N_34260);
xor U34573 (N_34573,N_34397,N_34467);
and U34574 (N_34574,N_34345,N_34301);
or U34575 (N_34575,N_34498,N_34282);
or U34576 (N_34576,N_34339,N_34281);
or U34577 (N_34577,N_34287,N_34495);
and U34578 (N_34578,N_34356,N_34367);
or U34579 (N_34579,N_34422,N_34458);
or U34580 (N_34580,N_34359,N_34326);
nor U34581 (N_34581,N_34405,N_34304);
nor U34582 (N_34582,N_34431,N_34270);
nand U34583 (N_34583,N_34473,N_34351);
and U34584 (N_34584,N_34277,N_34399);
xor U34585 (N_34585,N_34436,N_34452);
nor U34586 (N_34586,N_34402,N_34395);
or U34587 (N_34587,N_34484,N_34254);
nor U34588 (N_34588,N_34255,N_34352);
xnor U34589 (N_34589,N_34407,N_34482);
and U34590 (N_34590,N_34358,N_34336);
nor U34591 (N_34591,N_34252,N_34321);
xnor U34592 (N_34592,N_34265,N_34416);
or U34593 (N_34593,N_34370,N_34468);
or U34594 (N_34594,N_34483,N_34340);
xnor U34595 (N_34595,N_34251,N_34466);
nand U34596 (N_34596,N_34439,N_34396);
nand U34597 (N_34597,N_34313,N_34303);
nor U34598 (N_34598,N_34369,N_34443);
or U34599 (N_34599,N_34401,N_34288);
and U34600 (N_34600,N_34403,N_34332);
nor U34601 (N_34601,N_34404,N_34447);
or U34602 (N_34602,N_34419,N_34368);
or U34603 (N_34603,N_34296,N_34486);
nand U34604 (N_34604,N_34299,N_34424);
or U34605 (N_34605,N_34494,N_34309);
nand U34606 (N_34606,N_34258,N_34377);
nor U34607 (N_34607,N_34366,N_34308);
xor U34608 (N_34608,N_34276,N_34355);
and U34609 (N_34609,N_34379,N_34455);
or U34610 (N_34610,N_34423,N_34285);
nor U34611 (N_34611,N_34394,N_34421);
nor U34612 (N_34612,N_34306,N_34257);
or U34613 (N_34613,N_34427,N_34430);
or U34614 (N_34614,N_34444,N_34492);
nor U34615 (N_34615,N_34426,N_34283);
or U34616 (N_34616,N_34291,N_34485);
or U34617 (N_34617,N_34461,N_34496);
and U34618 (N_34618,N_34432,N_34267);
or U34619 (N_34619,N_34414,N_34390);
or U34620 (N_34620,N_34346,N_34488);
nand U34621 (N_34621,N_34410,N_34334);
nor U34622 (N_34622,N_34335,N_34438);
or U34623 (N_34623,N_34406,N_34322);
nor U34624 (N_34624,N_34381,N_34360);
nand U34625 (N_34625,N_34306,N_34277);
and U34626 (N_34626,N_34428,N_34286);
nor U34627 (N_34627,N_34461,N_34370);
nand U34628 (N_34628,N_34497,N_34394);
and U34629 (N_34629,N_34382,N_34319);
nand U34630 (N_34630,N_34446,N_34482);
xnor U34631 (N_34631,N_34446,N_34490);
nor U34632 (N_34632,N_34319,N_34274);
and U34633 (N_34633,N_34251,N_34477);
or U34634 (N_34634,N_34437,N_34339);
nor U34635 (N_34635,N_34480,N_34445);
or U34636 (N_34636,N_34261,N_34442);
xor U34637 (N_34637,N_34283,N_34371);
nand U34638 (N_34638,N_34279,N_34409);
and U34639 (N_34639,N_34458,N_34444);
and U34640 (N_34640,N_34413,N_34422);
or U34641 (N_34641,N_34396,N_34449);
or U34642 (N_34642,N_34368,N_34430);
nand U34643 (N_34643,N_34347,N_34339);
or U34644 (N_34644,N_34352,N_34374);
nand U34645 (N_34645,N_34306,N_34456);
xor U34646 (N_34646,N_34413,N_34370);
nand U34647 (N_34647,N_34454,N_34443);
and U34648 (N_34648,N_34380,N_34386);
nand U34649 (N_34649,N_34401,N_34384);
nor U34650 (N_34650,N_34341,N_34477);
and U34651 (N_34651,N_34398,N_34319);
nand U34652 (N_34652,N_34439,N_34455);
nand U34653 (N_34653,N_34435,N_34452);
and U34654 (N_34654,N_34461,N_34408);
or U34655 (N_34655,N_34401,N_34457);
xnor U34656 (N_34656,N_34363,N_34309);
or U34657 (N_34657,N_34444,N_34441);
nor U34658 (N_34658,N_34446,N_34412);
or U34659 (N_34659,N_34412,N_34484);
nand U34660 (N_34660,N_34362,N_34385);
nor U34661 (N_34661,N_34494,N_34270);
xor U34662 (N_34662,N_34376,N_34309);
nor U34663 (N_34663,N_34487,N_34395);
nand U34664 (N_34664,N_34438,N_34358);
nor U34665 (N_34665,N_34404,N_34250);
nand U34666 (N_34666,N_34250,N_34385);
nand U34667 (N_34667,N_34387,N_34276);
nor U34668 (N_34668,N_34497,N_34460);
or U34669 (N_34669,N_34251,N_34431);
nand U34670 (N_34670,N_34383,N_34489);
and U34671 (N_34671,N_34496,N_34377);
nor U34672 (N_34672,N_34368,N_34388);
and U34673 (N_34673,N_34393,N_34257);
xnor U34674 (N_34674,N_34405,N_34420);
nand U34675 (N_34675,N_34486,N_34291);
xor U34676 (N_34676,N_34432,N_34331);
and U34677 (N_34677,N_34351,N_34287);
or U34678 (N_34678,N_34352,N_34487);
nor U34679 (N_34679,N_34261,N_34371);
xor U34680 (N_34680,N_34498,N_34331);
nand U34681 (N_34681,N_34405,N_34380);
and U34682 (N_34682,N_34318,N_34349);
nand U34683 (N_34683,N_34482,N_34272);
nor U34684 (N_34684,N_34374,N_34439);
and U34685 (N_34685,N_34474,N_34261);
nand U34686 (N_34686,N_34394,N_34254);
or U34687 (N_34687,N_34379,N_34476);
nor U34688 (N_34688,N_34335,N_34453);
and U34689 (N_34689,N_34401,N_34458);
nor U34690 (N_34690,N_34371,N_34320);
nand U34691 (N_34691,N_34378,N_34493);
or U34692 (N_34692,N_34286,N_34318);
or U34693 (N_34693,N_34362,N_34368);
nor U34694 (N_34694,N_34369,N_34490);
or U34695 (N_34695,N_34369,N_34458);
and U34696 (N_34696,N_34262,N_34417);
nand U34697 (N_34697,N_34496,N_34353);
and U34698 (N_34698,N_34367,N_34498);
xnor U34699 (N_34699,N_34387,N_34264);
nand U34700 (N_34700,N_34330,N_34469);
xor U34701 (N_34701,N_34340,N_34314);
and U34702 (N_34702,N_34393,N_34274);
nand U34703 (N_34703,N_34469,N_34375);
nand U34704 (N_34704,N_34351,N_34310);
and U34705 (N_34705,N_34416,N_34378);
and U34706 (N_34706,N_34380,N_34439);
nor U34707 (N_34707,N_34393,N_34497);
nor U34708 (N_34708,N_34471,N_34467);
nor U34709 (N_34709,N_34276,N_34440);
xor U34710 (N_34710,N_34310,N_34279);
nor U34711 (N_34711,N_34438,N_34466);
nand U34712 (N_34712,N_34393,N_34396);
xor U34713 (N_34713,N_34390,N_34372);
nand U34714 (N_34714,N_34281,N_34296);
nand U34715 (N_34715,N_34496,N_34271);
nand U34716 (N_34716,N_34495,N_34340);
nor U34717 (N_34717,N_34283,N_34303);
nor U34718 (N_34718,N_34344,N_34498);
or U34719 (N_34719,N_34316,N_34434);
nor U34720 (N_34720,N_34417,N_34253);
or U34721 (N_34721,N_34252,N_34351);
nor U34722 (N_34722,N_34272,N_34310);
xor U34723 (N_34723,N_34318,N_34357);
and U34724 (N_34724,N_34386,N_34447);
or U34725 (N_34725,N_34351,N_34389);
or U34726 (N_34726,N_34405,N_34257);
nand U34727 (N_34727,N_34383,N_34275);
xor U34728 (N_34728,N_34354,N_34269);
or U34729 (N_34729,N_34477,N_34280);
and U34730 (N_34730,N_34457,N_34385);
xor U34731 (N_34731,N_34388,N_34473);
and U34732 (N_34732,N_34330,N_34259);
nand U34733 (N_34733,N_34433,N_34310);
and U34734 (N_34734,N_34411,N_34341);
xor U34735 (N_34735,N_34414,N_34412);
nor U34736 (N_34736,N_34493,N_34384);
nor U34737 (N_34737,N_34470,N_34305);
xnor U34738 (N_34738,N_34370,N_34489);
xor U34739 (N_34739,N_34363,N_34268);
nor U34740 (N_34740,N_34258,N_34465);
nand U34741 (N_34741,N_34323,N_34299);
nor U34742 (N_34742,N_34289,N_34275);
or U34743 (N_34743,N_34291,N_34396);
or U34744 (N_34744,N_34334,N_34370);
or U34745 (N_34745,N_34408,N_34441);
nand U34746 (N_34746,N_34359,N_34285);
nor U34747 (N_34747,N_34477,N_34269);
nand U34748 (N_34748,N_34433,N_34420);
or U34749 (N_34749,N_34439,N_34377);
nand U34750 (N_34750,N_34718,N_34631);
and U34751 (N_34751,N_34744,N_34679);
or U34752 (N_34752,N_34522,N_34530);
nor U34753 (N_34753,N_34720,N_34674);
or U34754 (N_34754,N_34587,N_34616);
nor U34755 (N_34755,N_34512,N_34698);
nand U34756 (N_34756,N_34584,N_34683);
nor U34757 (N_34757,N_34639,N_34517);
nor U34758 (N_34758,N_34513,N_34702);
nand U34759 (N_34759,N_34736,N_34693);
or U34760 (N_34760,N_34543,N_34711);
and U34761 (N_34761,N_34562,N_34690);
nand U34762 (N_34762,N_34538,N_34594);
xor U34763 (N_34763,N_34546,N_34723);
and U34764 (N_34764,N_34629,N_34595);
nor U34765 (N_34765,N_34531,N_34633);
or U34766 (N_34766,N_34678,N_34554);
nor U34767 (N_34767,N_34550,N_34710);
xnor U34768 (N_34768,N_34727,N_34614);
xor U34769 (N_34769,N_34511,N_34516);
nor U34770 (N_34770,N_34600,N_34520);
xnor U34771 (N_34771,N_34724,N_34505);
and U34772 (N_34772,N_34689,N_34604);
and U34773 (N_34773,N_34568,N_34721);
nor U34774 (N_34774,N_34575,N_34592);
and U34775 (N_34775,N_34561,N_34636);
or U34776 (N_34776,N_34749,N_34502);
xor U34777 (N_34777,N_34738,N_34688);
and U34778 (N_34778,N_34691,N_34703);
nor U34779 (N_34779,N_34729,N_34672);
nand U34780 (N_34780,N_34588,N_34748);
or U34781 (N_34781,N_34700,N_34500);
xor U34782 (N_34782,N_34529,N_34535);
xnor U34783 (N_34783,N_34685,N_34556);
or U34784 (N_34784,N_34746,N_34667);
or U34785 (N_34785,N_34548,N_34743);
and U34786 (N_34786,N_34694,N_34552);
xor U34787 (N_34787,N_34663,N_34670);
nor U34788 (N_34788,N_34553,N_34589);
or U34789 (N_34789,N_34585,N_34508);
or U34790 (N_34790,N_34571,N_34640);
or U34791 (N_34791,N_34622,N_34653);
xnor U34792 (N_34792,N_34591,N_34608);
nor U34793 (N_34793,N_34716,N_34652);
or U34794 (N_34794,N_34547,N_34647);
nor U34795 (N_34795,N_34687,N_34655);
and U34796 (N_34796,N_34680,N_34654);
nor U34797 (N_34797,N_34603,N_34573);
nor U34798 (N_34798,N_34740,N_34747);
and U34799 (N_34799,N_34545,N_34593);
and U34800 (N_34800,N_34521,N_34551);
and U34801 (N_34801,N_34705,N_34650);
nor U34802 (N_34802,N_34501,N_34659);
and U34803 (N_34803,N_34665,N_34628);
and U34804 (N_34804,N_34620,N_34519);
nor U34805 (N_34805,N_34596,N_34638);
and U34806 (N_34806,N_34684,N_34671);
and U34807 (N_34807,N_34560,N_34514);
and U34808 (N_34808,N_34737,N_34742);
and U34809 (N_34809,N_34506,N_34523);
nor U34810 (N_34810,N_34578,N_34612);
and U34811 (N_34811,N_34621,N_34722);
xnor U34812 (N_34812,N_34725,N_34527);
nor U34813 (N_34813,N_34615,N_34668);
nand U34814 (N_34814,N_34706,N_34682);
or U34815 (N_34815,N_34664,N_34701);
and U34816 (N_34816,N_34719,N_34731);
or U34817 (N_34817,N_34507,N_34569);
xor U34818 (N_34818,N_34558,N_34518);
or U34819 (N_34819,N_34717,N_34630);
nor U34820 (N_34820,N_34539,N_34657);
nor U34821 (N_34821,N_34632,N_34637);
or U34822 (N_34822,N_34576,N_34675);
nor U34823 (N_34823,N_34745,N_34618);
or U34824 (N_34824,N_34741,N_34651);
and U34825 (N_34825,N_34735,N_34697);
and U34826 (N_34826,N_34734,N_34607);
and U34827 (N_34827,N_34599,N_34601);
or U34828 (N_34828,N_34565,N_34714);
nor U34829 (N_34829,N_34732,N_34676);
nand U34830 (N_34830,N_34726,N_34627);
or U34831 (N_34831,N_34623,N_34634);
nand U34832 (N_34832,N_34686,N_34559);
or U34833 (N_34833,N_34515,N_34526);
nor U34834 (N_34834,N_34619,N_34577);
xor U34835 (N_34835,N_34524,N_34509);
nand U34836 (N_34836,N_34583,N_34606);
and U34837 (N_34837,N_34617,N_34555);
nor U34838 (N_34838,N_34635,N_34712);
and U34839 (N_34839,N_34549,N_34566);
or U34840 (N_34840,N_34626,N_34642);
xor U34841 (N_34841,N_34641,N_34673);
nand U34842 (N_34842,N_34537,N_34649);
or U34843 (N_34843,N_34610,N_34624);
nand U34844 (N_34844,N_34669,N_34536);
xor U34845 (N_34845,N_34658,N_34597);
and U34846 (N_34846,N_34661,N_34570);
xor U34847 (N_34847,N_34598,N_34681);
nand U34848 (N_34848,N_34580,N_34709);
and U34849 (N_34849,N_34542,N_34510);
nor U34850 (N_34850,N_34660,N_34544);
nand U34851 (N_34851,N_34704,N_34533);
xnor U34852 (N_34852,N_34730,N_34605);
or U34853 (N_34853,N_34564,N_34613);
nand U34854 (N_34854,N_34574,N_34567);
nor U34855 (N_34855,N_34609,N_34715);
nor U34856 (N_34856,N_34699,N_34586);
nand U34857 (N_34857,N_34534,N_34666);
and U34858 (N_34858,N_34611,N_34662);
nand U34859 (N_34859,N_34582,N_34503);
nor U34860 (N_34860,N_34728,N_34646);
xor U34861 (N_34861,N_34643,N_34528);
and U34862 (N_34862,N_34504,N_34645);
nor U34863 (N_34863,N_34625,N_34540);
or U34864 (N_34864,N_34532,N_34695);
nand U34865 (N_34865,N_34563,N_34656);
and U34866 (N_34866,N_34733,N_34677);
or U34867 (N_34867,N_34692,N_34541);
nand U34868 (N_34868,N_34708,N_34572);
xor U34869 (N_34869,N_34590,N_34739);
nor U34870 (N_34870,N_34579,N_34713);
nor U34871 (N_34871,N_34581,N_34707);
and U34872 (N_34872,N_34696,N_34644);
or U34873 (N_34873,N_34648,N_34525);
nand U34874 (N_34874,N_34602,N_34557);
xor U34875 (N_34875,N_34616,N_34631);
nor U34876 (N_34876,N_34734,N_34645);
and U34877 (N_34877,N_34584,N_34667);
nand U34878 (N_34878,N_34729,N_34503);
xor U34879 (N_34879,N_34626,N_34621);
nor U34880 (N_34880,N_34746,N_34539);
nand U34881 (N_34881,N_34647,N_34667);
or U34882 (N_34882,N_34509,N_34659);
nand U34883 (N_34883,N_34525,N_34719);
and U34884 (N_34884,N_34677,N_34657);
xnor U34885 (N_34885,N_34535,N_34742);
and U34886 (N_34886,N_34564,N_34632);
xnor U34887 (N_34887,N_34729,N_34566);
nand U34888 (N_34888,N_34653,N_34747);
nor U34889 (N_34889,N_34547,N_34686);
or U34890 (N_34890,N_34734,N_34739);
and U34891 (N_34891,N_34579,N_34691);
nor U34892 (N_34892,N_34536,N_34687);
xnor U34893 (N_34893,N_34690,N_34746);
and U34894 (N_34894,N_34585,N_34729);
nand U34895 (N_34895,N_34554,N_34694);
or U34896 (N_34896,N_34680,N_34524);
and U34897 (N_34897,N_34720,N_34560);
xor U34898 (N_34898,N_34562,N_34506);
or U34899 (N_34899,N_34585,N_34639);
nand U34900 (N_34900,N_34703,N_34585);
nor U34901 (N_34901,N_34523,N_34712);
nor U34902 (N_34902,N_34742,N_34515);
or U34903 (N_34903,N_34516,N_34529);
xor U34904 (N_34904,N_34576,N_34650);
nand U34905 (N_34905,N_34692,N_34527);
and U34906 (N_34906,N_34587,N_34636);
xnor U34907 (N_34907,N_34718,N_34501);
xor U34908 (N_34908,N_34731,N_34675);
nand U34909 (N_34909,N_34736,N_34566);
or U34910 (N_34910,N_34715,N_34653);
nor U34911 (N_34911,N_34564,N_34667);
and U34912 (N_34912,N_34629,N_34563);
nor U34913 (N_34913,N_34699,N_34742);
nor U34914 (N_34914,N_34555,N_34709);
or U34915 (N_34915,N_34587,N_34650);
or U34916 (N_34916,N_34738,N_34578);
and U34917 (N_34917,N_34545,N_34600);
nand U34918 (N_34918,N_34607,N_34534);
or U34919 (N_34919,N_34664,N_34601);
xor U34920 (N_34920,N_34626,N_34724);
xnor U34921 (N_34921,N_34679,N_34524);
nand U34922 (N_34922,N_34694,N_34680);
and U34923 (N_34923,N_34538,N_34730);
xnor U34924 (N_34924,N_34677,N_34739);
and U34925 (N_34925,N_34745,N_34638);
or U34926 (N_34926,N_34606,N_34582);
and U34927 (N_34927,N_34573,N_34514);
and U34928 (N_34928,N_34572,N_34698);
and U34929 (N_34929,N_34562,N_34718);
xnor U34930 (N_34930,N_34600,N_34681);
xnor U34931 (N_34931,N_34740,N_34509);
xnor U34932 (N_34932,N_34713,N_34582);
xor U34933 (N_34933,N_34620,N_34529);
nor U34934 (N_34934,N_34626,N_34674);
nand U34935 (N_34935,N_34743,N_34515);
nor U34936 (N_34936,N_34545,N_34653);
or U34937 (N_34937,N_34514,N_34603);
and U34938 (N_34938,N_34565,N_34553);
or U34939 (N_34939,N_34556,N_34716);
xor U34940 (N_34940,N_34541,N_34510);
xnor U34941 (N_34941,N_34663,N_34745);
nand U34942 (N_34942,N_34619,N_34676);
or U34943 (N_34943,N_34549,N_34741);
and U34944 (N_34944,N_34680,N_34636);
nor U34945 (N_34945,N_34683,N_34525);
xnor U34946 (N_34946,N_34531,N_34527);
nand U34947 (N_34947,N_34585,N_34646);
xnor U34948 (N_34948,N_34667,N_34631);
nor U34949 (N_34949,N_34697,N_34724);
nand U34950 (N_34950,N_34714,N_34511);
or U34951 (N_34951,N_34525,N_34559);
nand U34952 (N_34952,N_34647,N_34555);
or U34953 (N_34953,N_34629,N_34655);
nand U34954 (N_34954,N_34540,N_34552);
nand U34955 (N_34955,N_34649,N_34654);
or U34956 (N_34956,N_34732,N_34729);
nand U34957 (N_34957,N_34507,N_34710);
nand U34958 (N_34958,N_34564,N_34513);
nor U34959 (N_34959,N_34571,N_34501);
and U34960 (N_34960,N_34651,N_34642);
or U34961 (N_34961,N_34671,N_34590);
nor U34962 (N_34962,N_34749,N_34554);
and U34963 (N_34963,N_34648,N_34592);
nor U34964 (N_34964,N_34566,N_34653);
and U34965 (N_34965,N_34645,N_34724);
nand U34966 (N_34966,N_34510,N_34745);
nor U34967 (N_34967,N_34522,N_34646);
nor U34968 (N_34968,N_34703,N_34629);
nand U34969 (N_34969,N_34587,N_34535);
nor U34970 (N_34970,N_34559,N_34505);
xor U34971 (N_34971,N_34732,N_34733);
and U34972 (N_34972,N_34617,N_34718);
nand U34973 (N_34973,N_34533,N_34599);
xnor U34974 (N_34974,N_34650,N_34704);
nand U34975 (N_34975,N_34527,N_34632);
or U34976 (N_34976,N_34711,N_34560);
nor U34977 (N_34977,N_34638,N_34542);
xor U34978 (N_34978,N_34738,N_34500);
xnor U34979 (N_34979,N_34648,N_34614);
xor U34980 (N_34980,N_34621,N_34693);
or U34981 (N_34981,N_34631,N_34670);
and U34982 (N_34982,N_34582,N_34570);
xnor U34983 (N_34983,N_34710,N_34654);
and U34984 (N_34984,N_34715,N_34701);
xor U34985 (N_34985,N_34556,N_34597);
xor U34986 (N_34986,N_34643,N_34525);
xor U34987 (N_34987,N_34632,N_34580);
nand U34988 (N_34988,N_34590,N_34527);
nor U34989 (N_34989,N_34508,N_34738);
xor U34990 (N_34990,N_34745,N_34681);
nor U34991 (N_34991,N_34590,N_34651);
and U34992 (N_34992,N_34532,N_34674);
nand U34993 (N_34993,N_34509,N_34571);
and U34994 (N_34994,N_34713,N_34659);
nor U34995 (N_34995,N_34680,N_34677);
xnor U34996 (N_34996,N_34748,N_34680);
or U34997 (N_34997,N_34574,N_34519);
and U34998 (N_34998,N_34725,N_34561);
nand U34999 (N_34999,N_34620,N_34601);
nand U35000 (N_35000,N_34835,N_34883);
and U35001 (N_35001,N_34855,N_34892);
nor U35002 (N_35002,N_34980,N_34757);
nand U35003 (N_35003,N_34838,N_34863);
nand U35004 (N_35004,N_34888,N_34988);
nor U35005 (N_35005,N_34955,N_34813);
xor U35006 (N_35006,N_34793,N_34913);
and U35007 (N_35007,N_34925,N_34958);
xor U35008 (N_35008,N_34931,N_34805);
xor U35009 (N_35009,N_34930,N_34882);
nand U35010 (N_35010,N_34798,N_34964);
xnor U35011 (N_35011,N_34810,N_34845);
or U35012 (N_35012,N_34756,N_34830);
nor U35013 (N_35013,N_34812,N_34897);
nor U35014 (N_35014,N_34859,N_34962);
xnor U35015 (N_35015,N_34750,N_34939);
and U35016 (N_35016,N_34824,N_34850);
nand U35017 (N_35017,N_34954,N_34784);
or U35018 (N_35018,N_34848,N_34790);
xor U35019 (N_35019,N_34814,N_34949);
and U35020 (N_35020,N_34936,N_34841);
and U35021 (N_35021,N_34817,N_34942);
nor U35022 (N_35022,N_34754,N_34804);
or U35023 (N_35023,N_34788,N_34950);
or U35024 (N_35024,N_34986,N_34898);
xor U35025 (N_35025,N_34891,N_34965);
nor U35026 (N_35026,N_34865,N_34929);
xor U35027 (N_35027,N_34818,N_34956);
nand U35028 (N_35028,N_34975,N_34774);
xnor U35029 (N_35029,N_34787,N_34919);
or U35030 (N_35030,N_34806,N_34826);
nor U35031 (N_35031,N_34911,N_34844);
or U35032 (N_35032,N_34753,N_34775);
xnor U35033 (N_35033,N_34864,N_34760);
nand U35034 (N_35034,N_34837,N_34996);
xor U35035 (N_35035,N_34809,N_34857);
and U35036 (N_35036,N_34998,N_34991);
and U35037 (N_35037,N_34921,N_34825);
xnor U35038 (N_35038,N_34854,N_34785);
nand U35039 (N_35039,N_34764,N_34761);
nand U35040 (N_35040,N_34758,N_34786);
nand U35041 (N_35041,N_34867,N_34769);
or U35042 (N_35042,N_34852,N_34999);
nor U35043 (N_35043,N_34997,N_34872);
and U35044 (N_35044,N_34781,N_34895);
nand U35045 (N_35045,N_34928,N_34799);
xor U35046 (N_35046,N_34816,N_34934);
nand U35047 (N_35047,N_34943,N_34994);
or U35048 (N_35048,N_34766,N_34899);
and U35049 (N_35049,N_34952,N_34961);
xnor U35050 (N_35050,N_34778,N_34987);
nor U35051 (N_35051,N_34968,N_34909);
xor U35052 (N_35052,N_34861,N_34944);
or U35053 (N_35053,N_34796,N_34772);
and U35054 (N_35054,N_34941,N_34780);
and U35055 (N_35055,N_34822,N_34795);
and U35056 (N_35056,N_34908,N_34910);
and U35057 (N_35057,N_34840,N_34977);
xor U35058 (N_35058,N_34789,N_34992);
and U35059 (N_35059,N_34959,N_34896);
and U35060 (N_35060,N_34917,N_34920);
and U35061 (N_35061,N_34776,N_34937);
xnor U35062 (N_35062,N_34808,N_34759);
xor U35063 (N_35063,N_34971,N_34963);
and U35064 (N_35064,N_34792,N_34894);
or U35065 (N_35065,N_34948,N_34933);
xor U35066 (N_35066,N_34907,N_34803);
nand U35067 (N_35067,N_34960,N_34811);
xnor U35068 (N_35068,N_34981,N_34871);
xor U35069 (N_35069,N_34797,N_34983);
and U35070 (N_35070,N_34762,N_34938);
xor U35071 (N_35071,N_34771,N_34947);
or U35072 (N_35072,N_34881,N_34889);
nand U35073 (N_35073,N_34815,N_34833);
or U35074 (N_35074,N_34879,N_34755);
nand U35075 (N_35075,N_34945,N_34877);
nand U35076 (N_35076,N_34820,N_34885);
nor U35077 (N_35077,N_34970,N_34957);
xor U35078 (N_35078,N_34849,N_34801);
nor U35079 (N_35079,N_34876,N_34976);
nor U35080 (N_35080,N_34829,N_34782);
nor U35081 (N_35081,N_34884,N_34995);
nor U35082 (N_35082,N_34974,N_34869);
and U35083 (N_35083,N_34843,N_34924);
nor U35084 (N_35084,N_34777,N_34862);
xor U35085 (N_35085,N_34900,N_34873);
nor U35086 (N_35086,N_34993,N_34870);
nor U35087 (N_35087,N_34856,N_34779);
nand U35088 (N_35088,N_34946,N_34927);
xnor U35089 (N_35089,N_34767,N_34783);
nor U35090 (N_35090,N_34923,N_34972);
xnor U35091 (N_35091,N_34874,N_34800);
xnor U35092 (N_35092,N_34836,N_34973);
nand U35093 (N_35093,N_34878,N_34912);
nor U35094 (N_35094,N_34979,N_34906);
xor U35095 (N_35095,N_34773,N_34989);
and U35096 (N_35096,N_34967,N_34794);
or U35097 (N_35097,N_34860,N_34851);
nand U35098 (N_35098,N_34834,N_34922);
nor U35099 (N_35099,N_34802,N_34827);
and U35100 (N_35100,N_34880,N_34842);
xnor U35101 (N_35101,N_34831,N_34847);
nor U35102 (N_35102,N_34951,N_34770);
xnor U35103 (N_35103,N_34832,N_34904);
xnor U35104 (N_35104,N_34887,N_34953);
or U35105 (N_35105,N_34985,N_34763);
or U35106 (N_35106,N_34918,N_34875);
or U35107 (N_35107,N_34823,N_34940);
and U35108 (N_35108,N_34866,N_34768);
or U35109 (N_35109,N_34765,N_34752);
xnor U35110 (N_35110,N_34868,N_34926);
or U35111 (N_35111,N_34846,N_34902);
and U35112 (N_35112,N_34978,N_34966);
and U35113 (N_35113,N_34893,N_34935);
nor U35114 (N_35114,N_34828,N_34890);
or U35115 (N_35115,N_34916,N_34982);
nand U35116 (N_35116,N_34807,N_34751);
nand U35117 (N_35117,N_34791,N_34839);
or U35118 (N_35118,N_34901,N_34914);
nand U35119 (N_35119,N_34905,N_34903);
nor U35120 (N_35120,N_34853,N_34821);
xnor U35121 (N_35121,N_34932,N_34990);
xor U35122 (N_35122,N_34969,N_34984);
and U35123 (N_35123,N_34858,N_34915);
xnor U35124 (N_35124,N_34819,N_34886);
nor U35125 (N_35125,N_34811,N_34987);
xnor U35126 (N_35126,N_34896,N_34751);
nor U35127 (N_35127,N_34975,N_34914);
nor U35128 (N_35128,N_34962,N_34872);
nor U35129 (N_35129,N_34777,N_34880);
and U35130 (N_35130,N_34781,N_34765);
and U35131 (N_35131,N_34821,N_34817);
or U35132 (N_35132,N_34857,N_34877);
xor U35133 (N_35133,N_34916,N_34907);
nand U35134 (N_35134,N_34864,N_34841);
and U35135 (N_35135,N_34942,N_34982);
and U35136 (N_35136,N_34883,N_34957);
xor U35137 (N_35137,N_34752,N_34878);
xnor U35138 (N_35138,N_34791,N_34872);
or U35139 (N_35139,N_34762,N_34828);
or U35140 (N_35140,N_34802,N_34928);
xnor U35141 (N_35141,N_34840,N_34965);
or U35142 (N_35142,N_34831,N_34824);
or U35143 (N_35143,N_34984,N_34912);
nand U35144 (N_35144,N_34808,N_34859);
or U35145 (N_35145,N_34944,N_34910);
or U35146 (N_35146,N_34866,N_34880);
xnor U35147 (N_35147,N_34957,N_34800);
nor U35148 (N_35148,N_34826,N_34761);
nand U35149 (N_35149,N_34833,N_34926);
or U35150 (N_35150,N_34874,N_34944);
nor U35151 (N_35151,N_34980,N_34803);
and U35152 (N_35152,N_34777,N_34849);
xor U35153 (N_35153,N_34823,N_34838);
xnor U35154 (N_35154,N_34817,N_34939);
nor U35155 (N_35155,N_34965,N_34967);
nor U35156 (N_35156,N_34838,N_34980);
and U35157 (N_35157,N_34803,N_34759);
or U35158 (N_35158,N_34894,N_34753);
nor U35159 (N_35159,N_34943,N_34776);
or U35160 (N_35160,N_34897,N_34851);
and U35161 (N_35161,N_34760,N_34953);
and U35162 (N_35162,N_34902,N_34833);
nor U35163 (N_35163,N_34876,N_34806);
nor U35164 (N_35164,N_34991,N_34827);
and U35165 (N_35165,N_34926,N_34965);
nor U35166 (N_35166,N_34961,N_34975);
nand U35167 (N_35167,N_34818,N_34936);
xnor U35168 (N_35168,N_34809,N_34957);
xnor U35169 (N_35169,N_34998,N_34878);
and U35170 (N_35170,N_34955,N_34782);
and U35171 (N_35171,N_34842,N_34969);
nor U35172 (N_35172,N_34971,N_34881);
or U35173 (N_35173,N_34867,N_34923);
or U35174 (N_35174,N_34776,N_34849);
or U35175 (N_35175,N_34777,N_34963);
nand U35176 (N_35176,N_34876,N_34999);
nand U35177 (N_35177,N_34841,N_34995);
nand U35178 (N_35178,N_34804,N_34823);
or U35179 (N_35179,N_34887,N_34963);
nand U35180 (N_35180,N_34970,N_34912);
nor U35181 (N_35181,N_34784,N_34807);
nand U35182 (N_35182,N_34939,N_34959);
nand U35183 (N_35183,N_34870,N_34772);
and U35184 (N_35184,N_34776,N_34795);
or U35185 (N_35185,N_34900,N_34928);
or U35186 (N_35186,N_34800,N_34888);
or U35187 (N_35187,N_34935,N_34986);
nor U35188 (N_35188,N_34823,N_34917);
nor U35189 (N_35189,N_34975,N_34862);
nor U35190 (N_35190,N_34779,N_34877);
and U35191 (N_35191,N_34780,N_34862);
and U35192 (N_35192,N_34826,N_34913);
xor U35193 (N_35193,N_34808,N_34933);
or U35194 (N_35194,N_34917,N_34996);
and U35195 (N_35195,N_34866,N_34895);
nand U35196 (N_35196,N_34920,N_34763);
and U35197 (N_35197,N_34963,N_34793);
xnor U35198 (N_35198,N_34918,N_34871);
nor U35199 (N_35199,N_34797,N_34828);
or U35200 (N_35200,N_34951,N_34994);
nand U35201 (N_35201,N_34861,N_34995);
or U35202 (N_35202,N_34767,N_34983);
or U35203 (N_35203,N_34978,N_34912);
and U35204 (N_35204,N_34783,N_34992);
xnor U35205 (N_35205,N_34848,N_34778);
and U35206 (N_35206,N_34856,N_34818);
nand U35207 (N_35207,N_34823,N_34782);
and U35208 (N_35208,N_34851,N_34945);
nor U35209 (N_35209,N_34866,N_34835);
or U35210 (N_35210,N_34830,N_34910);
nand U35211 (N_35211,N_34895,N_34934);
or U35212 (N_35212,N_34846,N_34774);
or U35213 (N_35213,N_34963,N_34950);
nand U35214 (N_35214,N_34948,N_34800);
xor U35215 (N_35215,N_34847,N_34939);
nand U35216 (N_35216,N_34848,N_34958);
and U35217 (N_35217,N_34995,N_34989);
nor U35218 (N_35218,N_34940,N_34871);
nand U35219 (N_35219,N_34766,N_34758);
nand U35220 (N_35220,N_34778,N_34888);
xnor U35221 (N_35221,N_34750,N_34888);
and U35222 (N_35222,N_34811,N_34893);
xnor U35223 (N_35223,N_34821,N_34774);
xor U35224 (N_35224,N_34902,N_34884);
xor U35225 (N_35225,N_34836,N_34954);
nand U35226 (N_35226,N_34990,N_34808);
nand U35227 (N_35227,N_34885,N_34938);
and U35228 (N_35228,N_34873,N_34912);
nor U35229 (N_35229,N_34896,N_34866);
xnor U35230 (N_35230,N_34883,N_34968);
nor U35231 (N_35231,N_34847,N_34856);
and U35232 (N_35232,N_34790,N_34828);
xor U35233 (N_35233,N_34802,N_34838);
nand U35234 (N_35234,N_34996,N_34806);
xor U35235 (N_35235,N_34977,N_34752);
and U35236 (N_35236,N_34994,N_34816);
xor U35237 (N_35237,N_34949,N_34966);
and U35238 (N_35238,N_34905,N_34886);
nor U35239 (N_35239,N_34962,N_34835);
or U35240 (N_35240,N_34878,N_34947);
or U35241 (N_35241,N_34945,N_34951);
or U35242 (N_35242,N_34875,N_34883);
and U35243 (N_35243,N_34997,N_34766);
and U35244 (N_35244,N_34781,N_34930);
nand U35245 (N_35245,N_34835,N_34990);
and U35246 (N_35246,N_34960,N_34866);
or U35247 (N_35247,N_34765,N_34764);
nor U35248 (N_35248,N_34785,N_34914);
nand U35249 (N_35249,N_34862,N_34831);
xnor U35250 (N_35250,N_35154,N_35056);
nand U35251 (N_35251,N_35152,N_35137);
nor U35252 (N_35252,N_35170,N_35248);
nor U35253 (N_35253,N_35153,N_35197);
or U35254 (N_35254,N_35209,N_35242);
xnor U35255 (N_35255,N_35157,N_35091);
and U35256 (N_35256,N_35129,N_35050);
and U35257 (N_35257,N_35193,N_35133);
nor U35258 (N_35258,N_35236,N_35127);
and U35259 (N_35259,N_35076,N_35090);
and U35260 (N_35260,N_35169,N_35247);
nor U35261 (N_35261,N_35113,N_35034);
or U35262 (N_35262,N_35052,N_35245);
and U35263 (N_35263,N_35072,N_35223);
xor U35264 (N_35264,N_35174,N_35240);
nand U35265 (N_35265,N_35087,N_35118);
nor U35266 (N_35266,N_35032,N_35180);
xnor U35267 (N_35267,N_35017,N_35008);
nand U35268 (N_35268,N_35028,N_35198);
or U35269 (N_35269,N_35046,N_35201);
and U35270 (N_35270,N_35199,N_35016);
or U35271 (N_35271,N_35030,N_35018);
nand U35272 (N_35272,N_35234,N_35105);
and U35273 (N_35273,N_35196,N_35057);
or U35274 (N_35274,N_35039,N_35071);
nand U35275 (N_35275,N_35027,N_35086);
and U35276 (N_35276,N_35191,N_35235);
nand U35277 (N_35277,N_35121,N_35211);
xor U35278 (N_35278,N_35204,N_35115);
or U35279 (N_35279,N_35144,N_35213);
nand U35280 (N_35280,N_35110,N_35156);
nor U35281 (N_35281,N_35162,N_35000);
xnor U35282 (N_35282,N_35177,N_35062);
and U35283 (N_35283,N_35014,N_35058);
xnor U35284 (N_35284,N_35140,N_35094);
nor U35285 (N_35285,N_35220,N_35024);
nor U35286 (N_35286,N_35088,N_35120);
and U35287 (N_35287,N_35190,N_35045);
and U35288 (N_35288,N_35066,N_35098);
and U35289 (N_35289,N_35095,N_35015);
or U35290 (N_35290,N_35184,N_35202);
xnor U35291 (N_35291,N_35012,N_35188);
and U35292 (N_35292,N_35093,N_35044);
xnor U35293 (N_35293,N_35084,N_35216);
or U35294 (N_35294,N_35054,N_35228);
and U35295 (N_35295,N_35224,N_35053);
and U35296 (N_35296,N_35007,N_35033);
nand U35297 (N_35297,N_35059,N_35179);
nand U35298 (N_35298,N_35243,N_35219);
xnor U35299 (N_35299,N_35131,N_35151);
xnor U35300 (N_35300,N_35143,N_35205);
nand U35301 (N_35301,N_35080,N_35134);
nand U35302 (N_35302,N_35222,N_35023);
or U35303 (N_35303,N_35231,N_35172);
or U35304 (N_35304,N_35003,N_35020);
or U35305 (N_35305,N_35109,N_35155);
nand U35306 (N_35306,N_35117,N_35029);
nor U35307 (N_35307,N_35004,N_35005);
nand U35308 (N_35308,N_35065,N_35009);
nand U35309 (N_35309,N_35048,N_35025);
xnor U35310 (N_35310,N_35183,N_35064);
xor U35311 (N_35311,N_35145,N_35089);
and U35312 (N_35312,N_35161,N_35195);
nor U35313 (N_35313,N_35233,N_35103);
nor U35314 (N_35314,N_35073,N_35119);
or U35315 (N_35315,N_35104,N_35239);
and U35316 (N_35316,N_35075,N_35107);
and U35317 (N_35317,N_35002,N_35101);
xor U35318 (N_35318,N_35022,N_35112);
or U35319 (N_35319,N_35124,N_35100);
or U35320 (N_35320,N_35130,N_35167);
and U35321 (N_35321,N_35106,N_35141);
and U35322 (N_35322,N_35108,N_35189);
nand U35323 (N_35323,N_35206,N_35078);
nand U35324 (N_35324,N_35010,N_35001);
and U35325 (N_35325,N_35042,N_35159);
xnor U35326 (N_35326,N_35132,N_35122);
nand U35327 (N_35327,N_35246,N_35135);
nand U35328 (N_35328,N_35031,N_35125);
nor U35329 (N_35329,N_35229,N_35210);
nor U35330 (N_35330,N_35111,N_35081);
nand U35331 (N_35331,N_35035,N_35136);
or U35332 (N_35332,N_35043,N_35214);
xor U35333 (N_35333,N_35178,N_35067);
and U35334 (N_35334,N_35187,N_35225);
xnor U35335 (N_35335,N_35069,N_35102);
nand U35336 (N_35336,N_35051,N_35139);
and U35337 (N_35337,N_35194,N_35237);
nand U35338 (N_35338,N_35186,N_35068);
and U35339 (N_35339,N_35049,N_35181);
xnor U35340 (N_35340,N_35192,N_35146);
xor U35341 (N_35341,N_35083,N_35218);
or U35342 (N_35342,N_35176,N_35126);
nand U35343 (N_35343,N_35036,N_35166);
nand U35344 (N_35344,N_35160,N_35021);
and U35345 (N_35345,N_35226,N_35232);
or U35346 (N_35346,N_35182,N_35085);
and U35347 (N_35347,N_35055,N_35092);
or U35348 (N_35348,N_35038,N_35149);
or U35349 (N_35349,N_35171,N_35070);
nor U35350 (N_35350,N_35047,N_35215);
or U35351 (N_35351,N_35230,N_35173);
or U35352 (N_35352,N_35203,N_35150);
nor U35353 (N_35353,N_35099,N_35185);
nor U35354 (N_35354,N_35040,N_35168);
or U35355 (N_35355,N_35006,N_35019);
nand U35356 (N_35356,N_35096,N_35013);
or U35357 (N_35357,N_35165,N_35116);
and U35358 (N_35358,N_35074,N_35163);
or U35359 (N_35359,N_35241,N_35207);
xor U35360 (N_35360,N_35244,N_35227);
nor U35361 (N_35361,N_35063,N_35249);
nand U35362 (N_35362,N_35158,N_35097);
and U35363 (N_35363,N_35221,N_35208);
nand U35364 (N_35364,N_35148,N_35128);
or U35365 (N_35365,N_35200,N_35114);
nor U35366 (N_35366,N_35061,N_35123);
nor U35367 (N_35367,N_35082,N_35142);
xnor U35368 (N_35368,N_35079,N_35026);
nand U35369 (N_35369,N_35217,N_35011);
nand U35370 (N_35370,N_35238,N_35164);
and U35371 (N_35371,N_35060,N_35212);
nand U35372 (N_35372,N_35147,N_35138);
nand U35373 (N_35373,N_35041,N_35175);
or U35374 (N_35374,N_35077,N_35037);
or U35375 (N_35375,N_35213,N_35097);
nor U35376 (N_35376,N_35055,N_35180);
nor U35377 (N_35377,N_35183,N_35069);
nor U35378 (N_35378,N_35145,N_35131);
or U35379 (N_35379,N_35131,N_35019);
nand U35380 (N_35380,N_35110,N_35143);
xnor U35381 (N_35381,N_35115,N_35038);
xnor U35382 (N_35382,N_35169,N_35163);
or U35383 (N_35383,N_35130,N_35190);
xor U35384 (N_35384,N_35098,N_35015);
xnor U35385 (N_35385,N_35170,N_35024);
nor U35386 (N_35386,N_35224,N_35026);
nand U35387 (N_35387,N_35200,N_35001);
nor U35388 (N_35388,N_35171,N_35140);
nor U35389 (N_35389,N_35172,N_35080);
nor U35390 (N_35390,N_35175,N_35205);
or U35391 (N_35391,N_35089,N_35204);
xnor U35392 (N_35392,N_35151,N_35246);
nand U35393 (N_35393,N_35057,N_35129);
or U35394 (N_35394,N_35099,N_35186);
nand U35395 (N_35395,N_35169,N_35227);
nand U35396 (N_35396,N_35007,N_35123);
nand U35397 (N_35397,N_35235,N_35125);
or U35398 (N_35398,N_35029,N_35210);
xnor U35399 (N_35399,N_35161,N_35007);
nand U35400 (N_35400,N_35154,N_35087);
nand U35401 (N_35401,N_35114,N_35024);
nor U35402 (N_35402,N_35026,N_35033);
or U35403 (N_35403,N_35081,N_35233);
or U35404 (N_35404,N_35047,N_35115);
and U35405 (N_35405,N_35056,N_35010);
and U35406 (N_35406,N_35031,N_35200);
and U35407 (N_35407,N_35105,N_35163);
and U35408 (N_35408,N_35144,N_35001);
nor U35409 (N_35409,N_35128,N_35013);
or U35410 (N_35410,N_35214,N_35100);
nand U35411 (N_35411,N_35085,N_35140);
xnor U35412 (N_35412,N_35171,N_35075);
nand U35413 (N_35413,N_35068,N_35132);
and U35414 (N_35414,N_35207,N_35195);
nand U35415 (N_35415,N_35242,N_35205);
nor U35416 (N_35416,N_35103,N_35017);
nand U35417 (N_35417,N_35248,N_35007);
nand U35418 (N_35418,N_35031,N_35181);
and U35419 (N_35419,N_35011,N_35149);
nand U35420 (N_35420,N_35025,N_35143);
and U35421 (N_35421,N_35198,N_35116);
nor U35422 (N_35422,N_35141,N_35026);
and U35423 (N_35423,N_35003,N_35079);
xor U35424 (N_35424,N_35089,N_35149);
nand U35425 (N_35425,N_35185,N_35097);
and U35426 (N_35426,N_35026,N_35115);
nand U35427 (N_35427,N_35027,N_35196);
and U35428 (N_35428,N_35106,N_35073);
xnor U35429 (N_35429,N_35225,N_35012);
xnor U35430 (N_35430,N_35150,N_35097);
or U35431 (N_35431,N_35069,N_35208);
or U35432 (N_35432,N_35211,N_35153);
and U35433 (N_35433,N_35148,N_35124);
and U35434 (N_35434,N_35111,N_35096);
nor U35435 (N_35435,N_35007,N_35059);
or U35436 (N_35436,N_35013,N_35216);
xnor U35437 (N_35437,N_35235,N_35221);
nand U35438 (N_35438,N_35217,N_35080);
or U35439 (N_35439,N_35017,N_35180);
nor U35440 (N_35440,N_35019,N_35072);
xor U35441 (N_35441,N_35220,N_35187);
or U35442 (N_35442,N_35236,N_35104);
nor U35443 (N_35443,N_35235,N_35151);
or U35444 (N_35444,N_35050,N_35166);
nor U35445 (N_35445,N_35081,N_35180);
nor U35446 (N_35446,N_35209,N_35197);
xnor U35447 (N_35447,N_35167,N_35207);
nand U35448 (N_35448,N_35046,N_35044);
and U35449 (N_35449,N_35040,N_35220);
nor U35450 (N_35450,N_35057,N_35063);
and U35451 (N_35451,N_35236,N_35242);
xor U35452 (N_35452,N_35206,N_35199);
or U35453 (N_35453,N_35152,N_35134);
or U35454 (N_35454,N_35180,N_35021);
nand U35455 (N_35455,N_35202,N_35010);
nor U35456 (N_35456,N_35017,N_35211);
or U35457 (N_35457,N_35138,N_35208);
and U35458 (N_35458,N_35155,N_35119);
nor U35459 (N_35459,N_35099,N_35205);
and U35460 (N_35460,N_35149,N_35067);
and U35461 (N_35461,N_35212,N_35247);
or U35462 (N_35462,N_35012,N_35151);
nand U35463 (N_35463,N_35122,N_35184);
or U35464 (N_35464,N_35073,N_35055);
and U35465 (N_35465,N_35026,N_35219);
xnor U35466 (N_35466,N_35237,N_35116);
xnor U35467 (N_35467,N_35036,N_35081);
xor U35468 (N_35468,N_35100,N_35099);
nor U35469 (N_35469,N_35119,N_35015);
xor U35470 (N_35470,N_35092,N_35235);
or U35471 (N_35471,N_35118,N_35061);
xnor U35472 (N_35472,N_35198,N_35207);
nor U35473 (N_35473,N_35111,N_35057);
nor U35474 (N_35474,N_35241,N_35118);
and U35475 (N_35475,N_35183,N_35180);
nor U35476 (N_35476,N_35196,N_35003);
nor U35477 (N_35477,N_35073,N_35237);
nor U35478 (N_35478,N_35031,N_35168);
or U35479 (N_35479,N_35114,N_35069);
nand U35480 (N_35480,N_35155,N_35168);
and U35481 (N_35481,N_35150,N_35042);
nor U35482 (N_35482,N_35006,N_35192);
or U35483 (N_35483,N_35086,N_35233);
or U35484 (N_35484,N_35126,N_35232);
nor U35485 (N_35485,N_35121,N_35079);
nor U35486 (N_35486,N_35155,N_35103);
or U35487 (N_35487,N_35024,N_35203);
xor U35488 (N_35488,N_35078,N_35243);
xor U35489 (N_35489,N_35116,N_35069);
nand U35490 (N_35490,N_35035,N_35169);
or U35491 (N_35491,N_35038,N_35083);
nand U35492 (N_35492,N_35142,N_35109);
xnor U35493 (N_35493,N_35248,N_35091);
or U35494 (N_35494,N_35142,N_35080);
nand U35495 (N_35495,N_35088,N_35117);
and U35496 (N_35496,N_35232,N_35006);
or U35497 (N_35497,N_35090,N_35153);
xnor U35498 (N_35498,N_35049,N_35141);
nand U35499 (N_35499,N_35204,N_35194);
xnor U35500 (N_35500,N_35408,N_35393);
or U35501 (N_35501,N_35278,N_35392);
nand U35502 (N_35502,N_35475,N_35373);
and U35503 (N_35503,N_35411,N_35365);
and U35504 (N_35504,N_35439,N_35391);
nand U35505 (N_35505,N_35368,N_35428);
or U35506 (N_35506,N_35402,N_35495);
xor U35507 (N_35507,N_35390,N_35324);
xnor U35508 (N_35508,N_35294,N_35447);
or U35509 (N_35509,N_35273,N_35378);
and U35510 (N_35510,N_35289,N_35497);
and U35511 (N_35511,N_35277,N_35491);
and U35512 (N_35512,N_35425,N_35412);
nand U35513 (N_35513,N_35427,N_35356);
nand U35514 (N_35514,N_35317,N_35464);
nand U35515 (N_35515,N_35473,N_35271);
nor U35516 (N_35516,N_35252,N_35421);
xor U35517 (N_35517,N_35329,N_35337);
nor U35518 (N_35518,N_35265,N_35496);
xor U35519 (N_35519,N_35340,N_35443);
nor U35520 (N_35520,N_35266,N_35384);
and U35521 (N_35521,N_35326,N_35431);
xor U35522 (N_35522,N_35472,N_35469);
or U35523 (N_35523,N_35298,N_35311);
xnor U35524 (N_35524,N_35465,N_35344);
and U35525 (N_35525,N_35334,N_35293);
or U35526 (N_35526,N_35323,N_35260);
or U35527 (N_35527,N_35409,N_35254);
or U35528 (N_35528,N_35330,N_35463);
nand U35529 (N_35529,N_35314,N_35452);
xor U35530 (N_35530,N_35355,N_35436);
nand U35531 (N_35531,N_35288,N_35297);
nand U35532 (N_35532,N_35383,N_35492);
or U35533 (N_35533,N_35380,N_35397);
and U35534 (N_35534,N_35274,N_35370);
xor U35535 (N_35535,N_35299,N_35480);
or U35536 (N_35536,N_35419,N_35313);
and U35537 (N_35537,N_35435,N_35262);
or U35538 (N_35538,N_35346,N_35270);
or U35539 (N_35539,N_35461,N_35433);
xor U35540 (N_35540,N_35479,N_35400);
xnor U35541 (N_35541,N_35287,N_35424);
nand U35542 (N_35542,N_35338,N_35302);
nand U35543 (N_35543,N_35332,N_35386);
and U35544 (N_35544,N_35498,N_35410);
or U35545 (N_35545,N_35394,N_35426);
and U35546 (N_35546,N_35372,N_35375);
or U35547 (N_35547,N_35450,N_35485);
xor U35548 (N_35548,N_35458,N_35335);
or U35549 (N_35549,N_35477,N_35321);
nand U35550 (N_35550,N_35462,N_35490);
xor U35551 (N_35551,N_35357,N_35320);
and U35552 (N_35552,N_35445,N_35367);
or U35553 (N_35553,N_35369,N_35363);
and U35554 (N_35554,N_35381,N_35301);
and U35555 (N_35555,N_35296,N_35403);
nand U35556 (N_35556,N_35455,N_35251);
or U35557 (N_35557,N_35256,N_35449);
xor U35558 (N_35558,N_35257,N_35336);
nor U35559 (N_35559,N_35434,N_35347);
or U35560 (N_35560,N_35417,N_35269);
nand U35561 (N_35561,N_35290,N_35432);
and U35562 (N_35562,N_35413,N_35267);
and U35563 (N_35563,N_35395,N_35282);
or U35564 (N_35564,N_35328,N_35487);
nor U35565 (N_35565,N_35295,N_35483);
nand U35566 (N_35566,N_35429,N_35351);
xnor U35567 (N_35567,N_35376,N_35300);
xnor U35568 (N_35568,N_35468,N_35414);
and U35569 (N_35569,N_35339,N_35359);
and U35570 (N_35570,N_35404,N_35259);
and U35571 (N_35571,N_35308,N_35352);
xnor U35572 (N_35572,N_35307,N_35454);
nand U35573 (N_35573,N_35305,N_35283);
nor U35574 (N_35574,N_35258,N_35276);
and U35575 (N_35575,N_35250,N_35405);
and U35576 (N_35576,N_35399,N_35327);
or U35577 (N_35577,N_35420,N_35292);
nand U35578 (N_35578,N_35345,N_35440);
and U35579 (N_35579,N_35389,N_35291);
nand U35580 (N_35580,N_35488,N_35418);
or U35581 (N_35581,N_35309,N_35422);
xor U35582 (N_35582,N_35255,N_35285);
and U35583 (N_35583,N_35353,N_35319);
nor U35584 (N_35584,N_35310,N_35438);
and U35585 (N_35585,N_35437,N_35444);
nand U35586 (N_35586,N_35361,N_35358);
xor U35587 (N_35587,N_35481,N_35460);
or U35588 (N_35588,N_35261,N_35371);
nand U35589 (N_35589,N_35322,N_35388);
or U35590 (N_35590,N_35441,N_35448);
nor U35591 (N_35591,N_35489,N_35306);
and U35592 (N_35592,N_35467,N_35451);
or U35593 (N_35593,N_35423,N_35484);
and U35594 (N_35594,N_35430,N_35272);
nor U35595 (N_35595,N_35325,N_35348);
and U35596 (N_35596,N_35268,N_35398);
xor U35597 (N_35597,N_35407,N_35387);
xor U35598 (N_35598,N_35264,N_35478);
and U35599 (N_35599,N_35476,N_35280);
or U35600 (N_35600,N_35360,N_35362);
nand U35601 (N_35601,N_35456,N_35406);
nor U35602 (N_35602,N_35303,N_35499);
and U35603 (N_35603,N_35446,N_35415);
nand U35604 (N_35604,N_35316,N_35396);
or U35605 (N_35605,N_35284,N_35401);
and U35606 (N_35606,N_35341,N_35349);
and U35607 (N_35607,N_35364,N_35279);
nor U35608 (N_35608,N_35342,N_35482);
and U35609 (N_35609,N_35382,N_35333);
or U35610 (N_35610,N_35486,N_35474);
and U35611 (N_35611,N_35281,N_35493);
nand U35612 (N_35612,N_35416,N_35312);
and U35613 (N_35613,N_35315,N_35457);
and U35614 (N_35614,N_35354,N_35466);
and U35615 (N_35615,N_35374,N_35459);
or U35616 (N_35616,N_35379,N_35275);
or U35617 (N_35617,N_35350,N_35343);
or U35618 (N_35618,N_35286,N_35385);
nor U35619 (N_35619,N_35331,N_35442);
or U35620 (N_35620,N_35318,N_35253);
and U35621 (N_35621,N_35494,N_35470);
nor U35622 (N_35622,N_35377,N_35263);
xor U35623 (N_35623,N_35366,N_35471);
nand U35624 (N_35624,N_35453,N_35304);
nand U35625 (N_35625,N_35449,N_35318);
xor U35626 (N_35626,N_35289,N_35288);
or U35627 (N_35627,N_35418,N_35473);
or U35628 (N_35628,N_35318,N_35251);
nand U35629 (N_35629,N_35422,N_35310);
xor U35630 (N_35630,N_35446,N_35400);
or U35631 (N_35631,N_35475,N_35478);
nor U35632 (N_35632,N_35394,N_35346);
and U35633 (N_35633,N_35323,N_35392);
nor U35634 (N_35634,N_35401,N_35280);
nand U35635 (N_35635,N_35299,N_35340);
or U35636 (N_35636,N_35433,N_35280);
or U35637 (N_35637,N_35392,N_35452);
nor U35638 (N_35638,N_35450,N_35331);
xnor U35639 (N_35639,N_35377,N_35413);
nor U35640 (N_35640,N_35254,N_35333);
and U35641 (N_35641,N_35348,N_35456);
xor U35642 (N_35642,N_35449,N_35464);
nand U35643 (N_35643,N_35355,N_35494);
nand U35644 (N_35644,N_35442,N_35398);
nor U35645 (N_35645,N_35399,N_35445);
or U35646 (N_35646,N_35397,N_35477);
nand U35647 (N_35647,N_35339,N_35395);
nand U35648 (N_35648,N_35255,N_35313);
or U35649 (N_35649,N_35301,N_35264);
nor U35650 (N_35650,N_35275,N_35257);
or U35651 (N_35651,N_35431,N_35356);
or U35652 (N_35652,N_35307,N_35342);
and U35653 (N_35653,N_35254,N_35404);
nand U35654 (N_35654,N_35298,N_35379);
or U35655 (N_35655,N_35312,N_35283);
nand U35656 (N_35656,N_35354,N_35326);
or U35657 (N_35657,N_35390,N_35467);
nand U35658 (N_35658,N_35461,N_35431);
and U35659 (N_35659,N_35268,N_35390);
xnor U35660 (N_35660,N_35442,N_35496);
nand U35661 (N_35661,N_35254,N_35329);
and U35662 (N_35662,N_35361,N_35256);
nor U35663 (N_35663,N_35488,N_35305);
or U35664 (N_35664,N_35421,N_35402);
or U35665 (N_35665,N_35353,N_35347);
xnor U35666 (N_35666,N_35323,N_35432);
nand U35667 (N_35667,N_35465,N_35292);
or U35668 (N_35668,N_35292,N_35344);
nand U35669 (N_35669,N_35366,N_35258);
or U35670 (N_35670,N_35355,N_35377);
and U35671 (N_35671,N_35383,N_35264);
xnor U35672 (N_35672,N_35266,N_35396);
or U35673 (N_35673,N_35437,N_35421);
and U35674 (N_35674,N_35411,N_35308);
nor U35675 (N_35675,N_35358,N_35256);
and U35676 (N_35676,N_35467,N_35279);
nor U35677 (N_35677,N_35470,N_35259);
nor U35678 (N_35678,N_35376,N_35385);
or U35679 (N_35679,N_35459,N_35475);
or U35680 (N_35680,N_35277,N_35483);
nand U35681 (N_35681,N_35348,N_35362);
nand U35682 (N_35682,N_35324,N_35418);
nor U35683 (N_35683,N_35354,N_35433);
or U35684 (N_35684,N_35265,N_35464);
nor U35685 (N_35685,N_35450,N_35426);
nand U35686 (N_35686,N_35345,N_35402);
xnor U35687 (N_35687,N_35414,N_35412);
nor U35688 (N_35688,N_35498,N_35496);
xor U35689 (N_35689,N_35327,N_35460);
xor U35690 (N_35690,N_35481,N_35419);
nand U35691 (N_35691,N_35335,N_35319);
and U35692 (N_35692,N_35367,N_35360);
and U35693 (N_35693,N_35489,N_35260);
nand U35694 (N_35694,N_35361,N_35306);
nand U35695 (N_35695,N_35357,N_35267);
nor U35696 (N_35696,N_35324,N_35401);
nand U35697 (N_35697,N_35351,N_35404);
nand U35698 (N_35698,N_35348,N_35462);
or U35699 (N_35699,N_35269,N_35257);
xor U35700 (N_35700,N_35476,N_35468);
xor U35701 (N_35701,N_35298,N_35280);
xnor U35702 (N_35702,N_35406,N_35480);
nand U35703 (N_35703,N_35329,N_35456);
nor U35704 (N_35704,N_35342,N_35272);
or U35705 (N_35705,N_35477,N_35476);
nand U35706 (N_35706,N_35382,N_35319);
and U35707 (N_35707,N_35487,N_35466);
nand U35708 (N_35708,N_35449,N_35436);
nand U35709 (N_35709,N_35256,N_35338);
or U35710 (N_35710,N_35495,N_35376);
and U35711 (N_35711,N_35393,N_35454);
xor U35712 (N_35712,N_35462,N_35344);
and U35713 (N_35713,N_35398,N_35495);
nor U35714 (N_35714,N_35250,N_35450);
nor U35715 (N_35715,N_35429,N_35416);
nor U35716 (N_35716,N_35363,N_35387);
xnor U35717 (N_35717,N_35319,N_35380);
and U35718 (N_35718,N_35290,N_35396);
nand U35719 (N_35719,N_35387,N_35257);
and U35720 (N_35720,N_35456,N_35475);
and U35721 (N_35721,N_35414,N_35435);
or U35722 (N_35722,N_35376,N_35383);
xnor U35723 (N_35723,N_35277,N_35284);
nand U35724 (N_35724,N_35435,N_35264);
xnor U35725 (N_35725,N_35483,N_35467);
xnor U35726 (N_35726,N_35492,N_35483);
nor U35727 (N_35727,N_35393,N_35478);
or U35728 (N_35728,N_35345,N_35331);
nand U35729 (N_35729,N_35453,N_35477);
nor U35730 (N_35730,N_35343,N_35353);
nor U35731 (N_35731,N_35463,N_35398);
xor U35732 (N_35732,N_35449,N_35438);
nand U35733 (N_35733,N_35438,N_35422);
nor U35734 (N_35734,N_35327,N_35484);
nand U35735 (N_35735,N_35346,N_35340);
or U35736 (N_35736,N_35344,N_35351);
nor U35737 (N_35737,N_35487,N_35336);
nand U35738 (N_35738,N_35314,N_35481);
nand U35739 (N_35739,N_35416,N_35379);
and U35740 (N_35740,N_35296,N_35311);
xor U35741 (N_35741,N_35271,N_35445);
and U35742 (N_35742,N_35384,N_35334);
nor U35743 (N_35743,N_35313,N_35420);
nor U35744 (N_35744,N_35384,N_35474);
or U35745 (N_35745,N_35441,N_35488);
or U35746 (N_35746,N_35410,N_35353);
and U35747 (N_35747,N_35297,N_35277);
nor U35748 (N_35748,N_35274,N_35288);
nand U35749 (N_35749,N_35273,N_35463);
or U35750 (N_35750,N_35712,N_35665);
nand U35751 (N_35751,N_35554,N_35510);
nor U35752 (N_35752,N_35650,N_35562);
nor U35753 (N_35753,N_35611,N_35570);
or U35754 (N_35754,N_35578,N_35607);
and U35755 (N_35755,N_35672,N_35616);
nor U35756 (N_35756,N_35713,N_35580);
xor U35757 (N_35757,N_35559,N_35663);
and U35758 (N_35758,N_35660,N_35637);
nor U35759 (N_35759,N_35536,N_35626);
nor U35760 (N_35760,N_35649,N_35747);
xor U35761 (N_35761,N_35614,N_35659);
nand U35762 (N_35762,N_35549,N_35568);
xnor U35763 (N_35763,N_35593,N_35629);
and U35764 (N_35764,N_35581,N_35598);
or U35765 (N_35765,N_35688,N_35633);
xnor U35766 (N_35766,N_35682,N_35661);
and U35767 (N_35767,N_35675,N_35502);
or U35768 (N_35768,N_35621,N_35680);
nand U35769 (N_35769,N_35583,N_35622);
and U35770 (N_35770,N_35654,N_35523);
nand U35771 (N_35771,N_35511,N_35708);
nand U35772 (N_35772,N_35744,N_35571);
nand U35773 (N_35773,N_35695,N_35743);
nand U35774 (N_35774,N_35624,N_35513);
nor U35775 (N_35775,N_35730,N_35518);
or U35776 (N_35776,N_35636,N_35556);
nor U35777 (N_35777,N_35666,N_35699);
nor U35778 (N_35778,N_35718,N_35560);
nor U35779 (N_35779,N_35577,N_35534);
nor U35780 (N_35780,N_35725,N_35734);
nand U35781 (N_35781,N_35669,N_35603);
nand U35782 (N_35782,N_35528,N_35738);
or U35783 (N_35783,N_35612,N_35509);
nor U35784 (N_35784,N_35692,N_35646);
nor U35785 (N_35785,N_35749,N_35740);
xor U35786 (N_35786,N_35564,N_35574);
nor U35787 (N_35787,N_35613,N_35716);
nor U35788 (N_35788,N_35604,N_35671);
nor U35789 (N_35789,N_35670,N_35652);
or U35790 (N_35790,N_35573,N_35698);
nor U35791 (N_35791,N_35674,N_35679);
xnor U35792 (N_35792,N_35686,N_35543);
xnor U35793 (N_35793,N_35522,N_35504);
or U35794 (N_35794,N_35693,N_35736);
xnor U35795 (N_35795,N_35532,N_35507);
and U35796 (N_35796,N_35732,N_35569);
xnor U35797 (N_35797,N_35694,N_35677);
or U35798 (N_35798,N_35587,N_35628);
and U35799 (N_35799,N_35687,N_35605);
or U35800 (N_35800,N_35582,N_35527);
or U35801 (N_35801,N_35704,N_35703);
xnor U35802 (N_35802,N_35627,N_35602);
and U35803 (N_35803,N_35745,N_35741);
nand U35804 (N_35804,N_35617,N_35722);
nand U35805 (N_35805,N_35739,N_35707);
nor U35806 (N_35806,N_35702,N_35684);
or U35807 (N_35807,N_35538,N_35634);
nand U35808 (N_35808,N_35685,N_35592);
and U35809 (N_35809,N_35644,N_35548);
and U35810 (N_35810,N_35517,N_35653);
nand U35811 (N_35811,N_35563,N_35668);
nor U35812 (N_35812,N_35643,N_35726);
or U35813 (N_35813,N_35586,N_35589);
and U35814 (N_35814,N_35676,N_35552);
xnor U35815 (N_35815,N_35729,N_35544);
or U35816 (N_35816,N_35557,N_35706);
and U35817 (N_35817,N_35512,N_35508);
or U35818 (N_35818,N_35639,N_35608);
or U35819 (N_35819,N_35642,N_35524);
nand U35820 (N_35820,N_35535,N_35594);
or U35821 (N_35821,N_35638,N_35724);
and U35822 (N_35822,N_35648,N_35551);
nand U35823 (N_35823,N_35651,N_35678);
nand U35824 (N_35824,N_35742,N_35606);
xor U35825 (N_35825,N_35565,N_35516);
or U35826 (N_35826,N_35715,N_35541);
nor U35827 (N_35827,N_35727,N_35505);
nand U35828 (N_35828,N_35664,N_35537);
and U35829 (N_35829,N_35500,N_35545);
and U35830 (N_35830,N_35721,N_35585);
xor U35831 (N_35831,N_35689,N_35709);
and U35832 (N_35832,N_35667,N_35632);
nand U35833 (N_35833,N_35641,N_35540);
or U35834 (N_35834,N_35657,N_35719);
nand U35835 (N_35835,N_35596,N_35655);
or U35836 (N_35836,N_35572,N_35520);
and U35837 (N_35837,N_35550,N_35542);
xnor U35838 (N_35838,N_35600,N_35640);
nor U35839 (N_35839,N_35588,N_35601);
nor U35840 (N_35840,N_35717,N_35555);
nor U35841 (N_35841,N_35615,N_35690);
xor U35842 (N_35842,N_35701,N_35623);
and U35843 (N_35843,N_35566,N_35519);
nand U35844 (N_35844,N_35558,N_35567);
nand U35845 (N_35845,N_35561,N_35631);
nor U35846 (N_35846,N_35506,N_35590);
xnor U35847 (N_35847,N_35683,N_35625);
xor U35848 (N_35848,N_35515,N_35503);
and U35849 (N_35849,N_35501,N_35635);
or U35850 (N_35850,N_35620,N_35673);
and U35851 (N_35851,N_35526,N_35662);
or U35852 (N_35852,N_35746,N_35584);
or U35853 (N_35853,N_35647,N_35609);
nor U35854 (N_35854,N_35525,N_35539);
nor U35855 (N_35855,N_35546,N_35723);
nor U35856 (N_35856,N_35711,N_35514);
nand U35857 (N_35857,N_35530,N_35720);
or U35858 (N_35858,N_35710,N_35728);
or U35859 (N_35859,N_35656,N_35599);
or U35860 (N_35860,N_35591,N_35705);
nor U35861 (N_35861,N_35700,N_35533);
xor U35862 (N_35862,N_35521,N_35576);
xnor U35863 (N_35863,N_35553,N_35658);
nor U35864 (N_35864,N_35691,N_35531);
and U35865 (N_35865,N_35696,N_35733);
and U35866 (N_35866,N_35579,N_35748);
xor U35867 (N_35867,N_35681,N_35610);
nand U35868 (N_35868,N_35735,N_35714);
xnor U35869 (N_35869,N_35618,N_35547);
nand U35870 (N_35870,N_35697,N_35597);
nand U35871 (N_35871,N_35575,N_35595);
nand U35872 (N_35872,N_35529,N_35619);
xnor U35873 (N_35873,N_35630,N_35737);
and U35874 (N_35874,N_35731,N_35645);
and U35875 (N_35875,N_35524,N_35733);
xnor U35876 (N_35876,N_35735,N_35504);
nor U35877 (N_35877,N_35677,N_35533);
and U35878 (N_35878,N_35511,N_35744);
xor U35879 (N_35879,N_35748,N_35646);
nand U35880 (N_35880,N_35628,N_35749);
or U35881 (N_35881,N_35512,N_35509);
nor U35882 (N_35882,N_35523,N_35510);
nor U35883 (N_35883,N_35666,N_35644);
nand U35884 (N_35884,N_35550,N_35712);
nand U35885 (N_35885,N_35604,N_35599);
nand U35886 (N_35886,N_35582,N_35633);
nand U35887 (N_35887,N_35515,N_35719);
nand U35888 (N_35888,N_35702,N_35573);
or U35889 (N_35889,N_35650,N_35689);
nor U35890 (N_35890,N_35580,N_35639);
xor U35891 (N_35891,N_35685,N_35657);
or U35892 (N_35892,N_35671,N_35503);
xor U35893 (N_35893,N_35630,N_35746);
nor U35894 (N_35894,N_35625,N_35648);
nand U35895 (N_35895,N_35518,N_35561);
xor U35896 (N_35896,N_35614,N_35601);
nor U35897 (N_35897,N_35696,N_35612);
xnor U35898 (N_35898,N_35534,N_35646);
and U35899 (N_35899,N_35702,N_35691);
nand U35900 (N_35900,N_35515,N_35660);
and U35901 (N_35901,N_35722,N_35732);
or U35902 (N_35902,N_35732,N_35522);
and U35903 (N_35903,N_35717,N_35679);
and U35904 (N_35904,N_35726,N_35513);
nor U35905 (N_35905,N_35648,N_35521);
xor U35906 (N_35906,N_35734,N_35574);
or U35907 (N_35907,N_35694,N_35652);
and U35908 (N_35908,N_35515,N_35748);
nand U35909 (N_35909,N_35545,N_35721);
or U35910 (N_35910,N_35741,N_35518);
and U35911 (N_35911,N_35725,N_35723);
nor U35912 (N_35912,N_35696,N_35617);
nand U35913 (N_35913,N_35653,N_35730);
or U35914 (N_35914,N_35564,N_35643);
nand U35915 (N_35915,N_35706,N_35573);
xnor U35916 (N_35916,N_35569,N_35501);
and U35917 (N_35917,N_35731,N_35714);
xor U35918 (N_35918,N_35686,N_35619);
or U35919 (N_35919,N_35633,N_35689);
nand U35920 (N_35920,N_35580,N_35600);
xor U35921 (N_35921,N_35586,N_35537);
nor U35922 (N_35922,N_35590,N_35746);
nor U35923 (N_35923,N_35605,N_35586);
or U35924 (N_35924,N_35628,N_35542);
or U35925 (N_35925,N_35534,N_35720);
and U35926 (N_35926,N_35680,N_35564);
nand U35927 (N_35927,N_35642,N_35671);
or U35928 (N_35928,N_35523,N_35603);
nor U35929 (N_35929,N_35558,N_35675);
or U35930 (N_35930,N_35719,N_35705);
nor U35931 (N_35931,N_35513,N_35553);
or U35932 (N_35932,N_35585,N_35727);
or U35933 (N_35933,N_35522,N_35512);
or U35934 (N_35934,N_35669,N_35545);
nor U35935 (N_35935,N_35688,N_35505);
and U35936 (N_35936,N_35648,N_35526);
nand U35937 (N_35937,N_35590,N_35607);
and U35938 (N_35938,N_35603,N_35582);
nor U35939 (N_35939,N_35715,N_35727);
nand U35940 (N_35940,N_35607,N_35576);
nor U35941 (N_35941,N_35540,N_35609);
xor U35942 (N_35942,N_35614,N_35576);
xnor U35943 (N_35943,N_35713,N_35742);
xor U35944 (N_35944,N_35741,N_35734);
nand U35945 (N_35945,N_35696,N_35635);
or U35946 (N_35946,N_35576,N_35644);
or U35947 (N_35947,N_35640,N_35693);
xor U35948 (N_35948,N_35514,N_35748);
and U35949 (N_35949,N_35501,N_35652);
nor U35950 (N_35950,N_35527,N_35517);
nand U35951 (N_35951,N_35707,N_35559);
and U35952 (N_35952,N_35514,N_35592);
xnor U35953 (N_35953,N_35679,N_35599);
nand U35954 (N_35954,N_35707,N_35742);
nand U35955 (N_35955,N_35534,N_35728);
nor U35956 (N_35956,N_35624,N_35526);
nor U35957 (N_35957,N_35739,N_35656);
nor U35958 (N_35958,N_35534,N_35634);
nor U35959 (N_35959,N_35507,N_35634);
and U35960 (N_35960,N_35610,N_35636);
xor U35961 (N_35961,N_35532,N_35643);
and U35962 (N_35962,N_35590,N_35742);
nor U35963 (N_35963,N_35685,N_35531);
or U35964 (N_35964,N_35722,N_35645);
xor U35965 (N_35965,N_35685,N_35725);
xor U35966 (N_35966,N_35601,N_35700);
nor U35967 (N_35967,N_35721,N_35549);
nor U35968 (N_35968,N_35728,N_35621);
and U35969 (N_35969,N_35514,N_35557);
and U35970 (N_35970,N_35508,N_35665);
or U35971 (N_35971,N_35657,N_35593);
nand U35972 (N_35972,N_35551,N_35631);
nand U35973 (N_35973,N_35676,N_35658);
or U35974 (N_35974,N_35535,N_35700);
xnor U35975 (N_35975,N_35554,N_35519);
nand U35976 (N_35976,N_35649,N_35510);
xnor U35977 (N_35977,N_35512,N_35694);
xnor U35978 (N_35978,N_35748,N_35731);
or U35979 (N_35979,N_35701,N_35569);
and U35980 (N_35980,N_35659,N_35612);
nor U35981 (N_35981,N_35586,N_35625);
and U35982 (N_35982,N_35611,N_35520);
nor U35983 (N_35983,N_35662,N_35509);
nand U35984 (N_35984,N_35614,N_35632);
or U35985 (N_35985,N_35601,N_35507);
or U35986 (N_35986,N_35678,N_35674);
nor U35987 (N_35987,N_35674,N_35666);
nor U35988 (N_35988,N_35512,N_35727);
nor U35989 (N_35989,N_35734,N_35645);
or U35990 (N_35990,N_35583,N_35510);
nand U35991 (N_35991,N_35725,N_35650);
and U35992 (N_35992,N_35694,N_35598);
xnor U35993 (N_35993,N_35650,N_35736);
or U35994 (N_35994,N_35505,N_35622);
and U35995 (N_35995,N_35669,N_35544);
nand U35996 (N_35996,N_35525,N_35617);
nand U35997 (N_35997,N_35683,N_35724);
and U35998 (N_35998,N_35664,N_35731);
or U35999 (N_35999,N_35501,N_35725);
and U36000 (N_36000,N_35906,N_35861);
nand U36001 (N_36001,N_35859,N_35858);
nor U36002 (N_36002,N_35989,N_35759);
xor U36003 (N_36003,N_35843,N_35915);
xnor U36004 (N_36004,N_35812,N_35913);
and U36005 (N_36005,N_35959,N_35925);
nand U36006 (N_36006,N_35967,N_35780);
nand U36007 (N_36007,N_35831,N_35886);
nor U36008 (N_36008,N_35771,N_35995);
and U36009 (N_36009,N_35778,N_35969);
xor U36010 (N_36010,N_35908,N_35930);
nand U36011 (N_36011,N_35900,N_35945);
or U36012 (N_36012,N_35924,N_35835);
nor U36013 (N_36013,N_35820,N_35784);
xnor U36014 (N_36014,N_35755,N_35997);
nand U36015 (N_36015,N_35776,N_35871);
or U36016 (N_36016,N_35903,N_35762);
xnor U36017 (N_36017,N_35801,N_35792);
nor U36018 (N_36018,N_35754,N_35875);
xnor U36019 (N_36019,N_35993,N_35873);
xor U36020 (N_36020,N_35988,N_35898);
and U36021 (N_36021,N_35775,N_35793);
nand U36022 (N_36022,N_35788,N_35795);
and U36023 (N_36023,N_35847,N_35802);
nor U36024 (N_36024,N_35757,N_35981);
nand U36025 (N_36025,N_35951,N_35910);
and U36026 (N_36026,N_35880,N_35862);
xor U36027 (N_36027,N_35916,N_35773);
nor U36028 (N_36028,N_35899,N_35934);
and U36029 (N_36029,N_35881,N_35949);
or U36030 (N_36030,N_35817,N_35810);
or U36031 (N_36031,N_35994,N_35936);
and U36032 (N_36032,N_35944,N_35971);
xor U36033 (N_36033,N_35763,N_35987);
and U36034 (N_36034,N_35984,N_35955);
nand U36035 (N_36035,N_35846,N_35825);
or U36036 (N_36036,N_35766,N_35927);
xor U36037 (N_36037,N_35961,N_35806);
xnor U36038 (N_36038,N_35917,N_35853);
nor U36039 (N_36039,N_35956,N_35790);
nand U36040 (N_36040,N_35932,N_35937);
nor U36041 (N_36041,N_35824,N_35895);
and U36042 (N_36042,N_35879,N_35946);
or U36043 (N_36043,N_35919,N_35901);
and U36044 (N_36044,N_35756,N_35896);
or U36045 (N_36045,N_35912,N_35920);
and U36046 (N_36046,N_35844,N_35941);
nand U36047 (N_36047,N_35842,N_35797);
and U36048 (N_36048,N_35939,N_35863);
or U36049 (N_36049,N_35870,N_35933);
and U36050 (N_36050,N_35851,N_35772);
xnor U36051 (N_36051,N_35996,N_35965);
nor U36052 (N_36052,N_35891,N_35791);
or U36053 (N_36053,N_35991,N_35970);
or U36054 (N_36054,N_35992,N_35874);
and U36055 (N_36055,N_35911,N_35902);
nand U36056 (N_36056,N_35830,N_35809);
and U36057 (N_36057,N_35958,N_35882);
or U36058 (N_36058,N_35964,N_35781);
nand U36059 (N_36059,N_35977,N_35815);
nor U36060 (N_36060,N_35905,N_35926);
and U36061 (N_36061,N_35938,N_35867);
nand U36062 (N_36062,N_35856,N_35888);
or U36063 (N_36063,N_35887,N_35866);
xor U36064 (N_36064,N_35834,N_35808);
or U36065 (N_36065,N_35803,N_35990);
xnor U36066 (N_36066,N_35818,N_35782);
and U36067 (N_36067,N_35783,N_35811);
nor U36068 (N_36068,N_35804,N_35768);
or U36069 (N_36069,N_35962,N_35752);
or U36070 (N_36070,N_35979,N_35957);
xnor U36071 (N_36071,N_35904,N_35998);
nand U36072 (N_36072,N_35893,N_35827);
or U36073 (N_36073,N_35785,N_35884);
nor U36074 (N_36074,N_35897,N_35935);
nor U36075 (N_36075,N_35798,N_35805);
or U36076 (N_36076,N_35890,N_35813);
xor U36077 (N_36077,N_35889,N_35796);
nand U36078 (N_36078,N_35975,N_35950);
nand U36079 (N_36079,N_35865,N_35953);
nor U36080 (N_36080,N_35982,N_35857);
xnor U36081 (N_36081,N_35770,N_35814);
nand U36082 (N_36082,N_35828,N_35832);
or U36083 (N_36083,N_35860,N_35787);
xor U36084 (N_36084,N_35838,N_35850);
xor U36085 (N_36085,N_35909,N_35942);
or U36086 (N_36086,N_35819,N_35750);
nor U36087 (N_36087,N_35761,N_35878);
or U36088 (N_36088,N_35789,N_35940);
nand U36089 (N_36089,N_35849,N_35760);
nand U36090 (N_36090,N_35823,N_35929);
or U36091 (N_36091,N_35985,N_35877);
nand U36092 (N_36092,N_35931,N_35769);
xnor U36093 (N_36093,N_35826,N_35868);
and U36094 (N_36094,N_35972,N_35885);
and U36095 (N_36095,N_35751,N_35999);
xnor U36096 (N_36096,N_35774,N_35800);
nand U36097 (N_36097,N_35807,N_35883);
xnor U36098 (N_36098,N_35864,N_35777);
and U36099 (N_36099,N_35779,N_35845);
or U36100 (N_36100,N_35841,N_35952);
nor U36101 (N_36101,N_35869,N_35833);
nand U36102 (N_36102,N_35758,N_35764);
or U36103 (N_36103,N_35765,N_35923);
and U36104 (N_36104,N_35960,N_35974);
nor U36105 (N_36105,N_35907,N_35976);
nand U36106 (N_36106,N_35854,N_35892);
nor U36107 (N_36107,N_35839,N_35966);
xor U36108 (N_36108,N_35829,N_35799);
and U36109 (N_36109,N_35852,N_35821);
and U36110 (N_36110,N_35983,N_35978);
xnor U36111 (N_36111,N_35872,N_35963);
nor U36112 (N_36112,N_35921,N_35948);
or U36113 (N_36113,N_35918,N_35914);
nor U36114 (N_36114,N_35855,N_35922);
xor U36115 (N_36115,N_35943,N_35848);
nor U36116 (N_36116,N_35837,N_35954);
nand U36117 (N_36117,N_35836,N_35986);
or U36118 (N_36118,N_35973,N_35894);
nand U36119 (N_36119,N_35928,N_35840);
nor U36120 (N_36120,N_35794,N_35822);
xor U36121 (N_36121,N_35947,N_35753);
or U36122 (N_36122,N_35786,N_35767);
and U36123 (N_36123,N_35876,N_35968);
and U36124 (N_36124,N_35980,N_35816);
xor U36125 (N_36125,N_35992,N_35869);
nand U36126 (N_36126,N_35842,N_35845);
xnor U36127 (N_36127,N_35926,N_35955);
or U36128 (N_36128,N_35936,N_35758);
xnor U36129 (N_36129,N_35943,N_35998);
xor U36130 (N_36130,N_35797,N_35845);
xnor U36131 (N_36131,N_35988,N_35805);
nand U36132 (N_36132,N_35830,N_35919);
nand U36133 (N_36133,N_35862,N_35885);
xnor U36134 (N_36134,N_35862,N_35845);
or U36135 (N_36135,N_35750,N_35943);
xnor U36136 (N_36136,N_35926,N_35767);
nand U36137 (N_36137,N_35890,N_35968);
nor U36138 (N_36138,N_35898,N_35836);
or U36139 (N_36139,N_35912,N_35995);
nor U36140 (N_36140,N_35856,N_35900);
or U36141 (N_36141,N_35915,N_35919);
xor U36142 (N_36142,N_35811,N_35962);
and U36143 (N_36143,N_35754,N_35902);
nor U36144 (N_36144,N_35870,N_35817);
nand U36145 (N_36145,N_35959,N_35899);
or U36146 (N_36146,N_35786,N_35814);
or U36147 (N_36147,N_35758,N_35970);
xor U36148 (N_36148,N_35936,N_35785);
xor U36149 (N_36149,N_35894,N_35925);
nand U36150 (N_36150,N_35830,N_35994);
and U36151 (N_36151,N_35790,N_35980);
and U36152 (N_36152,N_35973,N_35802);
and U36153 (N_36153,N_35782,N_35849);
xor U36154 (N_36154,N_35898,N_35941);
nor U36155 (N_36155,N_35806,N_35878);
nand U36156 (N_36156,N_35772,N_35767);
nand U36157 (N_36157,N_35828,N_35980);
or U36158 (N_36158,N_35924,N_35948);
xnor U36159 (N_36159,N_35941,N_35996);
and U36160 (N_36160,N_35917,N_35875);
xor U36161 (N_36161,N_35951,N_35952);
xnor U36162 (N_36162,N_35788,N_35840);
nor U36163 (N_36163,N_35943,N_35810);
and U36164 (N_36164,N_35967,N_35912);
or U36165 (N_36165,N_35958,N_35808);
xor U36166 (N_36166,N_35914,N_35795);
or U36167 (N_36167,N_35922,N_35936);
nand U36168 (N_36168,N_35834,N_35752);
nand U36169 (N_36169,N_35908,N_35987);
xnor U36170 (N_36170,N_35919,N_35859);
and U36171 (N_36171,N_35973,N_35839);
nor U36172 (N_36172,N_35766,N_35844);
xor U36173 (N_36173,N_35948,N_35897);
or U36174 (N_36174,N_35958,N_35771);
nor U36175 (N_36175,N_35847,N_35868);
xnor U36176 (N_36176,N_35837,N_35982);
xnor U36177 (N_36177,N_35971,N_35992);
or U36178 (N_36178,N_35869,N_35947);
and U36179 (N_36179,N_35757,N_35943);
or U36180 (N_36180,N_35939,N_35891);
xor U36181 (N_36181,N_35794,N_35997);
or U36182 (N_36182,N_35895,N_35751);
xnor U36183 (N_36183,N_35791,N_35930);
and U36184 (N_36184,N_35870,N_35912);
nand U36185 (N_36185,N_35775,N_35901);
nor U36186 (N_36186,N_35953,N_35945);
and U36187 (N_36187,N_35918,N_35980);
and U36188 (N_36188,N_35916,N_35995);
xor U36189 (N_36189,N_35921,N_35961);
xnor U36190 (N_36190,N_35903,N_35996);
nor U36191 (N_36191,N_35839,N_35885);
and U36192 (N_36192,N_35858,N_35785);
or U36193 (N_36193,N_35893,N_35830);
nand U36194 (N_36194,N_35842,N_35941);
nor U36195 (N_36195,N_35988,N_35879);
or U36196 (N_36196,N_35780,N_35827);
and U36197 (N_36197,N_35998,N_35991);
nor U36198 (N_36198,N_35840,N_35768);
and U36199 (N_36199,N_35752,N_35860);
xor U36200 (N_36200,N_35770,N_35799);
and U36201 (N_36201,N_35760,N_35973);
and U36202 (N_36202,N_35890,N_35895);
nand U36203 (N_36203,N_35953,N_35818);
nor U36204 (N_36204,N_35897,N_35927);
or U36205 (N_36205,N_35878,N_35853);
nand U36206 (N_36206,N_35933,N_35901);
nor U36207 (N_36207,N_35930,N_35953);
or U36208 (N_36208,N_35776,N_35889);
and U36209 (N_36209,N_35934,N_35957);
nand U36210 (N_36210,N_35771,N_35942);
nor U36211 (N_36211,N_35863,N_35874);
or U36212 (N_36212,N_35966,N_35990);
nor U36213 (N_36213,N_35983,N_35779);
xor U36214 (N_36214,N_35837,N_35928);
and U36215 (N_36215,N_35878,N_35889);
nor U36216 (N_36216,N_35903,N_35975);
and U36217 (N_36217,N_35779,N_35920);
xor U36218 (N_36218,N_35910,N_35787);
and U36219 (N_36219,N_35838,N_35928);
and U36220 (N_36220,N_35768,N_35893);
xnor U36221 (N_36221,N_35814,N_35993);
nor U36222 (N_36222,N_35879,N_35933);
and U36223 (N_36223,N_35770,N_35754);
nand U36224 (N_36224,N_35938,N_35814);
nand U36225 (N_36225,N_35840,N_35920);
nand U36226 (N_36226,N_35822,N_35931);
or U36227 (N_36227,N_35793,N_35866);
nor U36228 (N_36228,N_35863,N_35836);
nand U36229 (N_36229,N_35810,N_35813);
nor U36230 (N_36230,N_35973,N_35886);
and U36231 (N_36231,N_35813,N_35872);
xnor U36232 (N_36232,N_35914,N_35850);
nor U36233 (N_36233,N_35763,N_35774);
or U36234 (N_36234,N_35776,N_35977);
nor U36235 (N_36235,N_35947,N_35940);
and U36236 (N_36236,N_35926,N_35833);
and U36237 (N_36237,N_35847,N_35877);
xor U36238 (N_36238,N_35924,N_35996);
and U36239 (N_36239,N_35850,N_35763);
nor U36240 (N_36240,N_35850,N_35946);
nor U36241 (N_36241,N_35827,N_35873);
nor U36242 (N_36242,N_35899,N_35816);
xor U36243 (N_36243,N_35798,N_35953);
nor U36244 (N_36244,N_35834,N_35987);
nor U36245 (N_36245,N_35816,N_35788);
nand U36246 (N_36246,N_35992,N_35832);
xnor U36247 (N_36247,N_35881,N_35966);
xnor U36248 (N_36248,N_35973,N_35963);
and U36249 (N_36249,N_35884,N_35780);
xor U36250 (N_36250,N_36116,N_36184);
or U36251 (N_36251,N_36245,N_36053);
or U36252 (N_36252,N_36020,N_36092);
nand U36253 (N_36253,N_36118,N_36067);
xor U36254 (N_36254,N_36002,N_36177);
or U36255 (N_36255,N_36080,N_36015);
or U36256 (N_36256,N_36155,N_36142);
nand U36257 (N_36257,N_36230,N_36145);
nand U36258 (N_36258,N_36138,N_36097);
nor U36259 (N_36259,N_36223,N_36041);
nor U36260 (N_36260,N_36115,N_36217);
xor U36261 (N_36261,N_36112,N_36072);
and U36262 (N_36262,N_36059,N_36058);
xor U36263 (N_36263,N_36218,N_36180);
or U36264 (N_36264,N_36154,N_36036);
nand U36265 (N_36265,N_36128,N_36068);
xnor U36266 (N_36266,N_36098,N_36205);
xor U36267 (N_36267,N_36091,N_36240);
or U36268 (N_36268,N_36221,N_36111);
and U36269 (N_36269,N_36212,N_36135);
xor U36270 (N_36270,N_36216,N_36214);
xnor U36271 (N_36271,N_36076,N_36123);
nand U36272 (N_36272,N_36120,N_36073);
xor U36273 (N_36273,N_36066,N_36191);
nor U36274 (N_36274,N_36082,N_36193);
nand U36275 (N_36275,N_36189,N_36083);
xnor U36276 (N_36276,N_36071,N_36108);
nand U36277 (N_36277,N_36125,N_36023);
nor U36278 (N_36278,N_36009,N_36074);
nor U36279 (N_36279,N_36011,N_36161);
nand U36280 (N_36280,N_36147,N_36045);
xor U36281 (N_36281,N_36163,N_36150);
and U36282 (N_36282,N_36236,N_36046);
or U36283 (N_36283,N_36167,N_36192);
or U36284 (N_36284,N_36124,N_36114);
and U36285 (N_36285,N_36033,N_36090);
xnor U36286 (N_36286,N_36085,N_36153);
nor U36287 (N_36287,N_36182,N_36219);
or U36288 (N_36288,N_36117,N_36172);
nor U36289 (N_36289,N_36007,N_36235);
xor U36290 (N_36290,N_36201,N_36141);
nand U36291 (N_36291,N_36113,N_36047);
nand U36292 (N_36292,N_36237,N_36086);
and U36293 (N_36293,N_36151,N_36241);
nand U36294 (N_36294,N_36137,N_36244);
or U36295 (N_36295,N_36231,N_36133);
nand U36296 (N_36296,N_36204,N_36040);
and U36297 (N_36297,N_36211,N_36243);
and U36298 (N_36298,N_36207,N_36035);
or U36299 (N_36299,N_36190,N_36144);
xnor U36300 (N_36300,N_36202,N_36065);
nand U36301 (N_36301,N_36158,N_36210);
xor U36302 (N_36302,N_36032,N_36100);
and U36303 (N_36303,N_36064,N_36176);
or U36304 (N_36304,N_36175,N_36183);
or U36305 (N_36305,N_36110,N_36042);
or U36306 (N_36306,N_36208,N_36044);
xnor U36307 (N_36307,N_36012,N_36061);
xor U36308 (N_36308,N_36018,N_36234);
and U36309 (N_36309,N_36198,N_36054);
nand U36310 (N_36310,N_36229,N_36103);
and U36311 (N_36311,N_36197,N_36186);
and U36312 (N_36312,N_36209,N_36049);
nand U36313 (N_36313,N_36050,N_36028);
or U36314 (N_36314,N_36052,N_36031);
or U36315 (N_36315,N_36140,N_36017);
nor U36316 (N_36316,N_36029,N_36179);
nand U36317 (N_36317,N_36106,N_36089);
nor U36318 (N_36318,N_36159,N_36087);
or U36319 (N_36319,N_36043,N_36199);
and U36320 (N_36320,N_36134,N_36078);
nor U36321 (N_36321,N_36019,N_36014);
nand U36322 (N_36322,N_36139,N_36121);
or U36323 (N_36323,N_36232,N_36249);
nand U36324 (N_36324,N_36056,N_36101);
nor U36325 (N_36325,N_36174,N_36149);
and U36326 (N_36326,N_36143,N_36195);
nand U36327 (N_36327,N_36006,N_36194);
nand U36328 (N_36328,N_36119,N_36130);
and U36329 (N_36329,N_36005,N_36132);
xnor U36330 (N_36330,N_36247,N_36157);
nor U36331 (N_36331,N_36156,N_36055);
xnor U36332 (N_36332,N_36099,N_36122);
or U36333 (N_36333,N_36181,N_36013);
nor U36334 (N_36334,N_36069,N_36025);
nor U36335 (N_36335,N_36060,N_36026);
nor U36336 (N_36336,N_36148,N_36188);
or U36337 (N_36337,N_36164,N_36173);
or U36338 (N_36338,N_36213,N_36004);
xnor U36339 (N_36339,N_36200,N_36169);
and U36340 (N_36340,N_36196,N_36062);
and U36341 (N_36341,N_36105,N_36070);
nand U36342 (N_36342,N_36129,N_36051);
and U36343 (N_36343,N_36246,N_36024);
nand U36344 (N_36344,N_36224,N_36206);
xor U36345 (N_36345,N_36225,N_36168);
and U36346 (N_36346,N_36010,N_36162);
and U36347 (N_36347,N_36003,N_36037);
and U36348 (N_36348,N_36242,N_36094);
or U36349 (N_36349,N_36170,N_36203);
xnor U36350 (N_36350,N_36187,N_36160);
nand U36351 (N_36351,N_36001,N_36222);
nand U36352 (N_36352,N_36022,N_36136);
and U36353 (N_36353,N_36081,N_36178);
and U36354 (N_36354,N_36107,N_36146);
and U36355 (N_36355,N_36126,N_36131);
or U36356 (N_36356,N_36021,N_36077);
nand U36357 (N_36357,N_36034,N_36008);
nand U36358 (N_36358,N_36096,N_36079);
and U36359 (N_36359,N_36084,N_36027);
xor U36360 (N_36360,N_36127,N_36063);
xnor U36361 (N_36361,N_36039,N_36233);
and U36362 (N_36362,N_36030,N_36088);
nand U36363 (N_36363,N_36248,N_36166);
and U36364 (N_36364,N_36220,N_36227);
or U36365 (N_36365,N_36239,N_36226);
nor U36366 (N_36366,N_36185,N_36109);
nor U36367 (N_36367,N_36171,N_36228);
or U36368 (N_36368,N_36095,N_36057);
or U36369 (N_36369,N_36038,N_36048);
and U36370 (N_36370,N_36000,N_36016);
or U36371 (N_36371,N_36104,N_36093);
nor U36372 (N_36372,N_36215,N_36238);
nand U36373 (N_36373,N_36102,N_36165);
or U36374 (N_36374,N_36075,N_36152);
nor U36375 (N_36375,N_36004,N_36098);
xnor U36376 (N_36376,N_36043,N_36141);
nand U36377 (N_36377,N_36122,N_36009);
nor U36378 (N_36378,N_36097,N_36135);
or U36379 (N_36379,N_36060,N_36115);
and U36380 (N_36380,N_36186,N_36127);
or U36381 (N_36381,N_36038,N_36213);
xnor U36382 (N_36382,N_36014,N_36163);
xor U36383 (N_36383,N_36098,N_36044);
or U36384 (N_36384,N_36023,N_36026);
nor U36385 (N_36385,N_36125,N_36088);
nor U36386 (N_36386,N_36183,N_36063);
nand U36387 (N_36387,N_36024,N_36213);
and U36388 (N_36388,N_36076,N_36024);
nor U36389 (N_36389,N_36056,N_36092);
nor U36390 (N_36390,N_36091,N_36078);
nor U36391 (N_36391,N_36222,N_36058);
xor U36392 (N_36392,N_36133,N_36068);
nand U36393 (N_36393,N_36231,N_36082);
xnor U36394 (N_36394,N_36001,N_36047);
nor U36395 (N_36395,N_36124,N_36031);
and U36396 (N_36396,N_36043,N_36068);
nor U36397 (N_36397,N_36208,N_36115);
and U36398 (N_36398,N_36180,N_36192);
and U36399 (N_36399,N_36062,N_36158);
nand U36400 (N_36400,N_36038,N_36104);
nor U36401 (N_36401,N_36180,N_36019);
nor U36402 (N_36402,N_36056,N_36244);
nor U36403 (N_36403,N_36078,N_36158);
or U36404 (N_36404,N_36022,N_36054);
nand U36405 (N_36405,N_36179,N_36075);
or U36406 (N_36406,N_36223,N_36200);
xor U36407 (N_36407,N_36181,N_36071);
nor U36408 (N_36408,N_36131,N_36245);
or U36409 (N_36409,N_36229,N_36153);
nor U36410 (N_36410,N_36113,N_36086);
nor U36411 (N_36411,N_36241,N_36231);
xor U36412 (N_36412,N_36159,N_36138);
nor U36413 (N_36413,N_36244,N_36027);
nand U36414 (N_36414,N_36127,N_36134);
nor U36415 (N_36415,N_36141,N_36033);
nor U36416 (N_36416,N_36181,N_36067);
xnor U36417 (N_36417,N_36104,N_36242);
and U36418 (N_36418,N_36236,N_36038);
or U36419 (N_36419,N_36003,N_36183);
xnor U36420 (N_36420,N_36132,N_36016);
nand U36421 (N_36421,N_36094,N_36123);
nor U36422 (N_36422,N_36157,N_36109);
xor U36423 (N_36423,N_36229,N_36127);
nand U36424 (N_36424,N_36189,N_36015);
and U36425 (N_36425,N_36035,N_36039);
nor U36426 (N_36426,N_36166,N_36180);
nand U36427 (N_36427,N_36113,N_36080);
nor U36428 (N_36428,N_36070,N_36249);
nor U36429 (N_36429,N_36215,N_36087);
nor U36430 (N_36430,N_36160,N_36054);
or U36431 (N_36431,N_36055,N_36062);
nor U36432 (N_36432,N_36056,N_36235);
nor U36433 (N_36433,N_36141,N_36016);
and U36434 (N_36434,N_36002,N_36246);
nor U36435 (N_36435,N_36228,N_36066);
xnor U36436 (N_36436,N_36240,N_36026);
and U36437 (N_36437,N_36196,N_36065);
nand U36438 (N_36438,N_36169,N_36189);
nor U36439 (N_36439,N_36183,N_36121);
and U36440 (N_36440,N_36214,N_36227);
nand U36441 (N_36441,N_36129,N_36152);
nand U36442 (N_36442,N_36111,N_36211);
or U36443 (N_36443,N_36104,N_36219);
and U36444 (N_36444,N_36063,N_36094);
and U36445 (N_36445,N_36000,N_36068);
and U36446 (N_36446,N_36171,N_36131);
nor U36447 (N_36447,N_36081,N_36233);
nand U36448 (N_36448,N_36064,N_36245);
and U36449 (N_36449,N_36044,N_36084);
nand U36450 (N_36450,N_36034,N_36070);
and U36451 (N_36451,N_36088,N_36047);
nor U36452 (N_36452,N_36152,N_36165);
or U36453 (N_36453,N_36173,N_36143);
xnor U36454 (N_36454,N_36228,N_36189);
nand U36455 (N_36455,N_36193,N_36234);
or U36456 (N_36456,N_36103,N_36075);
xnor U36457 (N_36457,N_36006,N_36187);
and U36458 (N_36458,N_36208,N_36079);
or U36459 (N_36459,N_36081,N_36232);
and U36460 (N_36460,N_36177,N_36180);
xnor U36461 (N_36461,N_36004,N_36220);
nand U36462 (N_36462,N_36194,N_36055);
or U36463 (N_36463,N_36221,N_36119);
or U36464 (N_36464,N_36087,N_36151);
nor U36465 (N_36465,N_36085,N_36125);
and U36466 (N_36466,N_36065,N_36217);
nand U36467 (N_36467,N_36075,N_36230);
and U36468 (N_36468,N_36048,N_36114);
xnor U36469 (N_36469,N_36141,N_36143);
and U36470 (N_36470,N_36015,N_36214);
nand U36471 (N_36471,N_36026,N_36052);
and U36472 (N_36472,N_36155,N_36214);
or U36473 (N_36473,N_36038,N_36154);
or U36474 (N_36474,N_36073,N_36067);
and U36475 (N_36475,N_36090,N_36217);
and U36476 (N_36476,N_36011,N_36074);
nor U36477 (N_36477,N_36222,N_36168);
or U36478 (N_36478,N_36039,N_36133);
xnor U36479 (N_36479,N_36008,N_36220);
nand U36480 (N_36480,N_36094,N_36084);
nor U36481 (N_36481,N_36154,N_36143);
or U36482 (N_36482,N_36069,N_36238);
nor U36483 (N_36483,N_36048,N_36191);
nand U36484 (N_36484,N_36021,N_36062);
xor U36485 (N_36485,N_36222,N_36093);
nand U36486 (N_36486,N_36240,N_36059);
nand U36487 (N_36487,N_36129,N_36066);
nor U36488 (N_36488,N_36137,N_36181);
and U36489 (N_36489,N_36244,N_36155);
nand U36490 (N_36490,N_36157,N_36015);
xnor U36491 (N_36491,N_36201,N_36146);
nor U36492 (N_36492,N_36013,N_36134);
or U36493 (N_36493,N_36070,N_36066);
xnor U36494 (N_36494,N_36155,N_36245);
or U36495 (N_36495,N_36033,N_36140);
nand U36496 (N_36496,N_36211,N_36150);
and U36497 (N_36497,N_36128,N_36211);
xnor U36498 (N_36498,N_36090,N_36242);
nor U36499 (N_36499,N_36091,N_36022);
or U36500 (N_36500,N_36438,N_36457);
or U36501 (N_36501,N_36308,N_36404);
or U36502 (N_36502,N_36327,N_36403);
and U36503 (N_36503,N_36332,N_36264);
xor U36504 (N_36504,N_36482,N_36448);
xnor U36505 (N_36505,N_36340,N_36333);
nand U36506 (N_36506,N_36278,N_36365);
and U36507 (N_36507,N_36255,N_36396);
nand U36508 (N_36508,N_36446,N_36271);
or U36509 (N_36509,N_36280,N_36428);
or U36510 (N_36510,N_36445,N_36490);
xor U36511 (N_36511,N_36319,N_36392);
xnor U36512 (N_36512,N_36492,N_36459);
and U36513 (N_36513,N_36330,N_36461);
nand U36514 (N_36514,N_36312,N_36373);
nand U36515 (N_36515,N_36410,N_36498);
nor U36516 (N_36516,N_36260,N_36393);
nor U36517 (N_36517,N_36353,N_36262);
nand U36518 (N_36518,N_36479,N_36360);
or U36519 (N_36519,N_36497,N_36417);
or U36520 (N_36520,N_36272,N_36366);
nor U36521 (N_36521,N_36345,N_36287);
nand U36522 (N_36522,N_36299,N_36383);
or U36523 (N_36523,N_36491,N_36375);
or U36524 (N_36524,N_36359,N_36306);
or U36525 (N_36525,N_36437,N_36391);
xnor U36526 (N_36526,N_36303,N_36368);
nand U36527 (N_36527,N_36488,N_36374);
xnor U36528 (N_36528,N_36313,N_36251);
and U36529 (N_36529,N_36415,N_36485);
nand U36530 (N_36530,N_36263,N_36290);
nor U36531 (N_36531,N_36371,N_36413);
or U36532 (N_36532,N_36387,N_36355);
nor U36533 (N_36533,N_36493,N_36378);
or U36534 (N_36534,N_36307,N_36351);
nand U36535 (N_36535,N_36289,N_36377);
nand U36536 (N_36536,N_36385,N_36369);
and U36537 (N_36537,N_36300,N_36380);
or U36538 (N_36538,N_36376,N_36399);
xor U36539 (N_36539,N_36442,N_36402);
or U36540 (N_36540,N_36476,N_36483);
nand U36541 (N_36541,N_36452,N_36274);
or U36542 (N_36542,N_36389,N_36397);
and U36543 (N_36543,N_36495,N_36408);
and U36544 (N_36544,N_36337,N_36462);
or U36545 (N_36545,N_36418,N_36284);
or U36546 (N_36546,N_36258,N_36394);
xor U36547 (N_36547,N_36296,N_36382);
and U36548 (N_36548,N_36405,N_36434);
nand U36549 (N_36549,N_36411,N_36325);
xnor U36550 (N_36550,N_36338,N_36266);
nand U36551 (N_36551,N_36322,N_36423);
nor U36552 (N_36552,N_36257,N_36460);
nand U36553 (N_36553,N_36318,N_36412);
and U36554 (N_36554,N_36270,N_36297);
nand U36555 (N_36555,N_36426,N_36254);
nor U36556 (N_36556,N_36265,N_36354);
xnor U36557 (N_36557,N_36269,N_36348);
or U36558 (N_36558,N_36499,N_36343);
nand U36559 (N_36559,N_36424,N_36283);
nand U36560 (N_36560,N_36430,N_36473);
nand U36561 (N_36561,N_36432,N_36304);
or U36562 (N_36562,N_36364,N_36294);
nand U36563 (N_36563,N_36302,N_36352);
and U36564 (N_36564,N_36349,N_36362);
xor U36565 (N_36565,N_36401,N_36468);
and U36566 (N_36566,N_36455,N_36346);
and U36567 (N_36567,N_36471,N_36475);
xnor U36568 (N_36568,N_36400,N_36470);
and U36569 (N_36569,N_36431,N_36358);
nor U36570 (N_36570,N_36441,N_36328);
xor U36571 (N_36571,N_36253,N_36489);
or U36572 (N_36572,N_36487,N_36316);
nor U36573 (N_36573,N_36429,N_36276);
nor U36574 (N_36574,N_36259,N_36285);
nor U36575 (N_36575,N_36494,N_36252);
or U36576 (N_36576,N_36464,N_36458);
and U36577 (N_36577,N_36291,N_36466);
nor U36578 (N_36578,N_36305,N_36469);
and U36579 (N_36579,N_36480,N_36261);
or U36580 (N_36580,N_36409,N_36453);
or U36581 (N_36581,N_36463,N_36425);
and U36582 (N_36582,N_36478,N_36422);
nand U36583 (N_36583,N_36277,N_36321);
nor U36584 (N_36584,N_36395,N_36406);
nor U36585 (N_36585,N_36449,N_36344);
and U36586 (N_36586,N_36314,N_36329);
or U36587 (N_36587,N_36384,N_36331);
or U36588 (N_36588,N_36496,N_36407);
xnor U36589 (N_36589,N_36367,N_36363);
nor U36590 (N_36590,N_36273,N_36436);
and U36591 (N_36591,N_36281,N_36390);
nor U36592 (N_36592,N_36311,N_36472);
nor U36593 (N_36593,N_36419,N_36372);
and U36594 (N_36594,N_36484,N_36323);
nor U36595 (N_36595,N_36465,N_36347);
xor U36596 (N_36596,N_36477,N_36456);
nand U36597 (N_36597,N_36467,N_36339);
nand U36598 (N_36598,N_36286,N_36326);
nor U36599 (N_36599,N_36298,N_36279);
xor U36600 (N_36600,N_36379,N_36310);
or U36601 (N_36601,N_36386,N_36335);
nand U36602 (N_36602,N_36342,N_36320);
and U36603 (N_36603,N_36268,N_36256);
or U36604 (N_36604,N_36435,N_36474);
nand U36605 (N_36605,N_36444,N_36288);
xor U36606 (N_36606,N_36443,N_36315);
nand U36607 (N_36607,N_36440,N_36454);
xor U36608 (N_36608,N_36293,N_36398);
or U36609 (N_36609,N_36450,N_36317);
and U36610 (N_36610,N_36421,N_36336);
and U36611 (N_36611,N_36414,N_36433);
nand U36612 (N_36612,N_36250,N_36481);
nor U36613 (N_36613,N_36295,N_36439);
nor U36614 (N_36614,N_36341,N_36334);
nor U36615 (N_36615,N_36356,N_36350);
xnor U36616 (N_36616,N_36267,N_36282);
or U36617 (N_36617,N_36486,N_36447);
nand U36618 (N_36618,N_36427,N_36416);
nor U36619 (N_36619,N_36292,N_36357);
nand U36620 (N_36620,N_36275,N_36361);
xnor U36621 (N_36621,N_36451,N_36301);
or U36622 (N_36622,N_36309,N_36388);
and U36623 (N_36623,N_36420,N_36370);
or U36624 (N_36624,N_36324,N_36381);
nor U36625 (N_36625,N_36450,N_36287);
and U36626 (N_36626,N_36416,N_36298);
and U36627 (N_36627,N_36340,N_36382);
xor U36628 (N_36628,N_36312,N_36328);
and U36629 (N_36629,N_36290,N_36348);
or U36630 (N_36630,N_36466,N_36386);
nand U36631 (N_36631,N_36262,N_36351);
nand U36632 (N_36632,N_36302,N_36309);
and U36633 (N_36633,N_36402,N_36405);
and U36634 (N_36634,N_36376,N_36353);
and U36635 (N_36635,N_36314,N_36303);
and U36636 (N_36636,N_36317,N_36292);
or U36637 (N_36637,N_36475,N_36384);
and U36638 (N_36638,N_36282,N_36481);
xnor U36639 (N_36639,N_36440,N_36348);
and U36640 (N_36640,N_36376,N_36395);
nor U36641 (N_36641,N_36456,N_36258);
or U36642 (N_36642,N_36451,N_36386);
or U36643 (N_36643,N_36357,N_36385);
nand U36644 (N_36644,N_36362,N_36339);
nor U36645 (N_36645,N_36412,N_36285);
nor U36646 (N_36646,N_36472,N_36267);
or U36647 (N_36647,N_36396,N_36439);
or U36648 (N_36648,N_36391,N_36485);
nor U36649 (N_36649,N_36278,N_36413);
nand U36650 (N_36650,N_36350,N_36318);
nor U36651 (N_36651,N_36426,N_36283);
and U36652 (N_36652,N_36316,N_36284);
nand U36653 (N_36653,N_36343,N_36432);
nand U36654 (N_36654,N_36361,N_36472);
and U36655 (N_36655,N_36333,N_36394);
and U36656 (N_36656,N_36410,N_36373);
xnor U36657 (N_36657,N_36463,N_36335);
and U36658 (N_36658,N_36491,N_36269);
or U36659 (N_36659,N_36423,N_36301);
nor U36660 (N_36660,N_36390,N_36371);
and U36661 (N_36661,N_36277,N_36324);
or U36662 (N_36662,N_36273,N_36252);
xnor U36663 (N_36663,N_36376,N_36277);
nor U36664 (N_36664,N_36380,N_36255);
nand U36665 (N_36665,N_36477,N_36304);
nand U36666 (N_36666,N_36297,N_36493);
nor U36667 (N_36667,N_36375,N_36465);
nor U36668 (N_36668,N_36314,N_36420);
nor U36669 (N_36669,N_36254,N_36485);
and U36670 (N_36670,N_36251,N_36364);
nor U36671 (N_36671,N_36492,N_36397);
nand U36672 (N_36672,N_36320,N_36457);
or U36673 (N_36673,N_36297,N_36278);
nand U36674 (N_36674,N_36405,N_36272);
xnor U36675 (N_36675,N_36428,N_36360);
nand U36676 (N_36676,N_36384,N_36419);
nand U36677 (N_36677,N_36427,N_36415);
or U36678 (N_36678,N_36420,N_36337);
nand U36679 (N_36679,N_36331,N_36254);
nand U36680 (N_36680,N_36394,N_36470);
nand U36681 (N_36681,N_36315,N_36415);
nand U36682 (N_36682,N_36291,N_36392);
nor U36683 (N_36683,N_36321,N_36452);
nand U36684 (N_36684,N_36305,N_36451);
or U36685 (N_36685,N_36414,N_36458);
or U36686 (N_36686,N_36349,N_36265);
nand U36687 (N_36687,N_36330,N_36362);
nand U36688 (N_36688,N_36304,N_36381);
nor U36689 (N_36689,N_36497,N_36334);
or U36690 (N_36690,N_36465,N_36259);
and U36691 (N_36691,N_36452,N_36430);
nor U36692 (N_36692,N_36260,N_36442);
nor U36693 (N_36693,N_36254,N_36359);
nor U36694 (N_36694,N_36311,N_36482);
or U36695 (N_36695,N_36419,N_36438);
or U36696 (N_36696,N_36326,N_36360);
nand U36697 (N_36697,N_36472,N_36265);
xnor U36698 (N_36698,N_36278,N_36367);
or U36699 (N_36699,N_36418,N_36276);
nor U36700 (N_36700,N_36268,N_36281);
nor U36701 (N_36701,N_36298,N_36442);
or U36702 (N_36702,N_36298,N_36294);
nor U36703 (N_36703,N_36464,N_36251);
or U36704 (N_36704,N_36341,N_36304);
nor U36705 (N_36705,N_36397,N_36445);
xor U36706 (N_36706,N_36331,N_36484);
and U36707 (N_36707,N_36348,N_36316);
and U36708 (N_36708,N_36274,N_36347);
nand U36709 (N_36709,N_36407,N_36477);
xnor U36710 (N_36710,N_36352,N_36437);
nor U36711 (N_36711,N_36314,N_36441);
nand U36712 (N_36712,N_36424,N_36346);
nor U36713 (N_36713,N_36482,N_36390);
and U36714 (N_36714,N_36417,N_36368);
or U36715 (N_36715,N_36441,N_36330);
and U36716 (N_36716,N_36395,N_36480);
or U36717 (N_36717,N_36453,N_36359);
and U36718 (N_36718,N_36442,N_36374);
nor U36719 (N_36719,N_36333,N_36356);
nor U36720 (N_36720,N_36281,N_36459);
nor U36721 (N_36721,N_36493,N_36446);
and U36722 (N_36722,N_36333,N_36294);
and U36723 (N_36723,N_36330,N_36414);
nand U36724 (N_36724,N_36342,N_36387);
nand U36725 (N_36725,N_36312,N_36341);
and U36726 (N_36726,N_36254,N_36475);
xor U36727 (N_36727,N_36288,N_36446);
and U36728 (N_36728,N_36455,N_36474);
xnor U36729 (N_36729,N_36415,N_36408);
xor U36730 (N_36730,N_36486,N_36408);
nand U36731 (N_36731,N_36308,N_36463);
xnor U36732 (N_36732,N_36327,N_36318);
xor U36733 (N_36733,N_36310,N_36360);
xnor U36734 (N_36734,N_36342,N_36424);
nor U36735 (N_36735,N_36475,N_36379);
and U36736 (N_36736,N_36458,N_36255);
xnor U36737 (N_36737,N_36305,N_36474);
nor U36738 (N_36738,N_36497,N_36255);
or U36739 (N_36739,N_36330,N_36374);
xor U36740 (N_36740,N_36418,N_36358);
or U36741 (N_36741,N_36368,N_36418);
and U36742 (N_36742,N_36324,N_36320);
or U36743 (N_36743,N_36352,N_36312);
nand U36744 (N_36744,N_36477,N_36495);
nand U36745 (N_36745,N_36376,N_36252);
and U36746 (N_36746,N_36323,N_36277);
xnor U36747 (N_36747,N_36339,N_36493);
nand U36748 (N_36748,N_36388,N_36451);
and U36749 (N_36749,N_36378,N_36454);
nand U36750 (N_36750,N_36655,N_36580);
nor U36751 (N_36751,N_36611,N_36579);
xor U36752 (N_36752,N_36624,N_36744);
or U36753 (N_36753,N_36646,N_36673);
nor U36754 (N_36754,N_36612,N_36657);
nand U36755 (N_36755,N_36535,N_36648);
xor U36756 (N_36756,N_36514,N_36537);
and U36757 (N_36757,N_36699,N_36576);
or U36758 (N_36758,N_36713,N_36630);
and U36759 (N_36759,N_36735,N_36543);
or U36760 (N_36760,N_36637,N_36678);
nor U36761 (N_36761,N_36723,N_36586);
nor U36762 (N_36762,N_36725,N_36668);
or U36763 (N_36763,N_36741,N_36683);
nor U36764 (N_36764,N_36531,N_36519);
xor U36765 (N_36765,N_36704,N_36603);
nand U36766 (N_36766,N_36548,N_36726);
xor U36767 (N_36767,N_36712,N_36555);
nor U36768 (N_36768,N_36598,N_36690);
and U36769 (N_36769,N_36584,N_36564);
xor U36770 (N_36770,N_36567,N_36529);
and U36771 (N_36771,N_36572,N_36560);
and U36772 (N_36772,N_36626,N_36717);
nand U36773 (N_36773,N_36512,N_36595);
or U36774 (N_36774,N_36643,N_36628);
or U36775 (N_36775,N_36711,N_36731);
or U36776 (N_36776,N_36588,N_36621);
and U36777 (N_36777,N_36502,N_36620);
nand U36778 (N_36778,N_36720,N_36739);
nand U36779 (N_36779,N_36634,N_36526);
nand U36780 (N_36780,N_36728,N_36700);
and U36781 (N_36781,N_36594,N_36672);
xnor U36782 (N_36782,N_36654,N_36638);
and U36783 (N_36783,N_36604,N_36610);
xnor U36784 (N_36784,N_36695,N_36600);
nand U36785 (N_36785,N_36517,N_36568);
nor U36786 (N_36786,N_36671,N_36685);
nor U36787 (N_36787,N_36591,N_36633);
nand U36788 (N_36788,N_36684,N_36550);
and U36789 (N_36789,N_36544,N_36736);
and U36790 (N_36790,N_36571,N_36602);
or U36791 (N_36791,N_36641,N_36619);
nand U36792 (N_36792,N_36734,N_36748);
and U36793 (N_36793,N_36592,N_36737);
xor U36794 (N_36794,N_36709,N_36599);
nor U36795 (N_36795,N_36503,N_36509);
and U36796 (N_36796,N_36623,N_36651);
and U36797 (N_36797,N_36719,N_36642);
nor U36798 (N_36798,N_36631,N_36557);
or U36799 (N_36799,N_36528,N_36504);
and U36800 (N_36800,N_36727,N_36636);
xor U36801 (N_36801,N_36746,N_36617);
xnor U36802 (N_36802,N_36570,N_36689);
xor U36803 (N_36803,N_36688,N_36694);
nand U36804 (N_36804,N_36582,N_36743);
nor U36805 (N_36805,N_36670,N_36687);
nor U36806 (N_36806,N_36587,N_36625);
nand U36807 (N_36807,N_36506,N_36547);
nor U36808 (N_36808,N_36664,N_36534);
nand U36809 (N_36809,N_36615,N_36697);
xor U36810 (N_36810,N_36682,N_36705);
or U36811 (N_36811,N_36540,N_36585);
or U36812 (N_36812,N_36500,N_36613);
or U36813 (N_36813,N_36703,N_36573);
and U36814 (N_36814,N_36522,N_36561);
nor U36815 (N_36815,N_36606,N_36562);
xnor U36816 (N_36816,N_36663,N_36674);
nand U36817 (N_36817,N_36702,N_36549);
nor U36818 (N_36818,N_36732,N_36590);
or U36819 (N_36819,N_36541,N_36618);
nor U36820 (N_36820,N_36733,N_36523);
nor U36821 (N_36821,N_36644,N_36607);
or U36822 (N_36822,N_36552,N_36505);
or U36823 (N_36823,N_36533,N_36647);
nand U36824 (N_36824,N_36658,N_36708);
nor U36825 (N_36825,N_36559,N_36577);
xnor U36826 (N_36826,N_36681,N_36539);
and U36827 (N_36827,N_36551,N_36578);
and U36828 (N_36828,N_36738,N_36546);
nor U36829 (N_36829,N_36536,N_36721);
or U36830 (N_36830,N_36525,N_36652);
and U36831 (N_36831,N_36501,N_36740);
xnor U36832 (N_36832,N_36521,N_36558);
nor U36833 (N_36833,N_36718,N_36622);
nand U36834 (N_36834,N_36605,N_36710);
xnor U36835 (N_36835,N_36507,N_36542);
or U36836 (N_36836,N_36608,N_36589);
nor U36837 (N_36837,N_36632,N_36575);
and U36838 (N_36838,N_36563,N_36715);
nor U36839 (N_36839,N_36698,N_36722);
xnor U36840 (N_36840,N_36516,N_36554);
nor U36841 (N_36841,N_36569,N_36706);
and U36842 (N_36842,N_36749,N_36692);
nand U36843 (N_36843,N_36675,N_36538);
or U36844 (N_36844,N_36532,N_36614);
nand U36845 (N_36845,N_36601,N_36686);
or U36846 (N_36846,N_36639,N_36530);
xnor U36847 (N_36847,N_36691,N_36665);
nand U36848 (N_36848,N_36680,N_36742);
nor U36849 (N_36849,N_36716,N_36724);
and U36850 (N_36850,N_36645,N_36565);
nor U36851 (N_36851,N_36520,N_36729);
nor U36852 (N_36852,N_36635,N_36661);
nor U36853 (N_36853,N_36609,N_36696);
nor U36854 (N_36854,N_36640,N_36574);
and U36855 (N_36855,N_36662,N_36747);
or U36856 (N_36856,N_36745,N_36597);
nand U36857 (N_36857,N_36656,N_36508);
and U36858 (N_36858,N_36524,N_36596);
nor U36859 (N_36859,N_36593,N_36545);
or U36860 (N_36860,N_36616,N_36566);
or U36861 (N_36861,N_36627,N_36511);
nor U36862 (N_36862,N_36730,N_36556);
nor U36863 (N_36863,N_36653,N_36581);
nand U36864 (N_36864,N_36679,N_36553);
and U36865 (N_36865,N_36714,N_36583);
nor U36866 (N_36866,N_36513,N_36666);
or U36867 (N_36867,N_36667,N_36650);
nand U36868 (N_36868,N_36660,N_36518);
nor U36869 (N_36869,N_36693,N_36707);
xnor U36870 (N_36870,N_36649,N_36510);
and U36871 (N_36871,N_36676,N_36515);
nor U36872 (N_36872,N_36669,N_36659);
nor U36873 (N_36873,N_36701,N_36629);
or U36874 (N_36874,N_36677,N_36527);
and U36875 (N_36875,N_36595,N_36714);
nand U36876 (N_36876,N_36502,N_36628);
nor U36877 (N_36877,N_36561,N_36681);
or U36878 (N_36878,N_36607,N_36566);
or U36879 (N_36879,N_36594,N_36512);
nor U36880 (N_36880,N_36601,N_36679);
nand U36881 (N_36881,N_36603,N_36732);
and U36882 (N_36882,N_36656,N_36689);
or U36883 (N_36883,N_36580,N_36712);
or U36884 (N_36884,N_36555,N_36583);
or U36885 (N_36885,N_36565,N_36700);
xnor U36886 (N_36886,N_36664,N_36639);
and U36887 (N_36887,N_36708,N_36635);
xor U36888 (N_36888,N_36684,N_36706);
nor U36889 (N_36889,N_36605,N_36729);
xnor U36890 (N_36890,N_36687,N_36714);
or U36891 (N_36891,N_36619,N_36540);
nand U36892 (N_36892,N_36578,N_36686);
or U36893 (N_36893,N_36613,N_36666);
and U36894 (N_36894,N_36586,N_36743);
or U36895 (N_36895,N_36692,N_36687);
xor U36896 (N_36896,N_36703,N_36501);
and U36897 (N_36897,N_36555,N_36648);
nor U36898 (N_36898,N_36666,N_36640);
or U36899 (N_36899,N_36584,N_36693);
xnor U36900 (N_36900,N_36708,N_36744);
and U36901 (N_36901,N_36522,N_36568);
or U36902 (N_36902,N_36667,N_36520);
or U36903 (N_36903,N_36712,N_36538);
and U36904 (N_36904,N_36668,N_36529);
xnor U36905 (N_36905,N_36630,N_36569);
xor U36906 (N_36906,N_36630,N_36507);
xor U36907 (N_36907,N_36577,N_36522);
xnor U36908 (N_36908,N_36718,N_36613);
and U36909 (N_36909,N_36614,N_36580);
and U36910 (N_36910,N_36506,N_36560);
nand U36911 (N_36911,N_36743,N_36520);
nor U36912 (N_36912,N_36597,N_36680);
nand U36913 (N_36913,N_36734,N_36551);
nand U36914 (N_36914,N_36611,N_36628);
nor U36915 (N_36915,N_36686,N_36747);
or U36916 (N_36916,N_36557,N_36740);
xnor U36917 (N_36917,N_36702,N_36628);
and U36918 (N_36918,N_36636,N_36645);
xnor U36919 (N_36919,N_36723,N_36526);
nand U36920 (N_36920,N_36731,N_36709);
or U36921 (N_36921,N_36650,N_36579);
and U36922 (N_36922,N_36575,N_36582);
and U36923 (N_36923,N_36685,N_36584);
or U36924 (N_36924,N_36538,N_36595);
nor U36925 (N_36925,N_36666,N_36560);
or U36926 (N_36926,N_36686,N_36571);
and U36927 (N_36927,N_36692,N_36612);
nor U36928 (N_36928,N_36693,N_36536);
and U36929 (N_36929,N_36606,N_36514);
xnor U36930 (N_36930,N_36511,N_36645);
and U36931 (N_36931,N_36662,N_36504);
nand U36932 (N_36932,N_36647,N_36652);
nor U36933 (N_36933,N_36742,N_36650);
and U36934 (N_36934,N_36697,N_36630);
nor U36935 (N_36935,N_36706,N_36663);
or U36936 (N_36936,N_36683,N_36541);
and U36937 (N_36937,N_36654,N_36644);
xnor U36938 (N_36938,N_36727,N_36744);
or U36939 (N_36939,N_36657,N_36735);
nand U36940 (N_36940,N_36508,N_36650);
nand U36941 (N_36941,N_36666,N_36664);
and U36942 (N_36942,N_36725,N_36634);
and U36943 (N_36943,N_36626,N_36566);
xnor U36944 (N_36944,N_36616,N_36610);
nand U36945 (N_36945,N_36671,N_36536);
nand U36946 (N_36946,N_36686,N_36732);
and U36947 (N_36947,N_36557,N_36735);
xor U36948 (N_36948,N_36512,N_36672);
xnor U36949 (N_36949,N_36576,N_36729);
xor U36950 (N_36950,N_36520,N_36542);
xor U36951 (N_36951,N_36634,N_36589);
or U36952 (N_36952,N_36622,N_36570);
and U36953 (N_36953,N_36573,N_36693);
or U36954 (N_36954,N_36567,N_36676);
and U36955 (N_36955,N_36626,N_36652);
or U36956 (N_36956,N_36675,N_36599);
or U36957 (N_36957,N_36560,N_36644);
or U36958 (N_36958,N_36588,N_36601);
and U36959 (N_36959,N_36740,N_36615);
xnor U36960 (N_36960,N_36543,N_36502);
nor U36961 (N_36961,N_36618,N_36505);
nand U36962 (N_36962,N_36656,N_36733);
nor U36963 (N_36963,N_36532,N_36649);
xor U36964 (N_36964,N_36662,N_36581);
nor U36965 (N_36965,N_36622,N_36585);
and U36966 (N_36966,N_36613,N_36655);
and U36967 (N_36967,N_36523,N_36736);
xor U36968 (N_36968,N_36536,N_36670);
and U36969 (N_36969,N_36694,N_36567);
nor U36970 (N_36970,N_36615,N_36743);
nand U36971 (N_36971,N_36703,N_36579);
and U36972 (N_36972,N_36581,N_36625);
nor U36973 (N_36973,N_36733,N_36596);
nor U36974 (N_36974,N_36556,N_36651);
nor U36975 (N_36975,N_36591,N_36514);
or U36976 (N_36976,N_36709,N_36677);
and U36977 (N_36977,N_36668,N_36609);
nor U36978 (N_36978,N_36683,N_36746);
and U36979 (N_36979,N_36674,N_36702);
or U36980 (N_36980,N_36711,N_36568);
and U36981 (N_36981,N_36679,N_36723);
or U36982 (N_36982,N_36709,N_36650);
nor U36983 (N_36983,N_36704,N_36544);
nand U36984 (N_36984,N_36513,N_36699);
nor U36985 (N_36985,N_36637,N_36671);
xor U36986 (N_36986,N_36609,N_36728);
and U36987 (N_36987,N_36516,N_36627);
nand U36988 (N_36988,N_36694,N_36587);
xor U36989 (N_36989,N_36531,N_36627);
or U36990 (N_36990,N_36659,N_36627);
or U36991 (N_36991,N_36581,N_36652);
nor U36992 (N_36992,N_36646,N_36617);
or U36993 (N_36993,N_36562,N_36644);
nor U36994 (N_36994,N_36670,N_36697);
xnor U36995 (N_36995,N_36504,N_36670);
nor U36996 (N_36996,N_36534,N_36680);
nand U36997 (N_36997,N_36741,N_36623);
and U36998 (N_36998,N_36562,N_36563);
and U36999 (N_36999,N_36588,N_36709);
or U37000 (N_37000,N_36783,N_36818);
nand U37001 (N_37001,N_36808,N_36835);
nand U37002 (N_37002,N_36995,N_36825);
and U37003 (N_37003,N_36877,N_36785);
or U37004 (N_37004,N_36916,N_36888);
or U37005 (N_37005,N_36895,N_36985);
and U37006 (N_37006,N_36816,N_36983);
nor U37007 (N_37007,N_36991,N_36942);
xor U37008 (N_37008,N_36950,N_36860);
nand U37009 (N_37009,N_36922,N_36798);
and U37010 (N_37010,N_36973,N_36960);
nor U37011 (N_37011,N_36897,N_36750);
nor U37012 (N_37012,N_36886,N_36866);
nand U37013 (N_37013,N_36878,N_36924);
nor U37014 (N_37014,N_36794,N_36815);
nor U37015 (N_37015,N_36787,N_36752);
nand U37016 (N_37016,N_36976,N_36863);
nand U37017 (N_37017,N_36887,N_36817);
nand U37018 (N_37018,N_36765,N_36837);
or U37019 (N_37019,N_36993,N_36826);
and U37020 (N_37020,N_36987,N_36846);
nand U37021 (N_37021,N_36864,N_36780);
xnor U37022 (N_37022,N_36795,N_36968);
xnor U37023 (N_37023,N_36900,N_36961);
or U37024 (N_37024,N_36937,N_36777);
xnor U37025 (N_37025,N_36938,N_36756);
xnor U37026 (N_37026,N_36881,N_36963);
or U37027 (N_37027,N_36905,N_36824);
xnor U37028 (N_37028,N_36933,N_36941);
or U37029 (N_37029,N_36969,N_36977);
or U37030 (N_37030,N_36940,N_36834);
nand U37031 (N_37031,N_36909,N_36885);
and U37032 (N_37032,N_36774,N_36845);
or U37033 (N_37033,N_36989,N_36844);
nor U37034 (N_37034,N_36978,N_36855);
nor U37035 (N_37035,N_36988,N_36853);
and U37036 (N_37036,N_36776,N_36788);
nand U37037 (N_37037,N_36904,N_36974);
nand U37038 (N_37038,N_36936,N_36962);
or U37039 (N_37039,N_36859,N_36896);
nor U37040 (N_37040,N_36959,N_36838);
xor U37041 (N_37041,N_36869,N_36791);
or U37042 (N_37042,N_36994,N_36934);
xor U37043 (N_37043,N_36814,N_36753);
or U37044 (N_37044,N_36832,N_36767);
nor U37045 (N_37045,N_36759,N_36918);
and U37046 (N_37046,N_36883,N_36819);
xnor U37047 (N_37047,N_36910,N_36899);
nor U37048 (N_37048,N_36872,N_36912);
nor U37049 (N_37049,N_36944,N_36884);
and U37050 (N_37050,N_36840,N_36958);
nor U37051 (N_37051,N_36820,N_36980);
or U37052 (N_37052,N_36799,N_36992);
nor U37053 (N_37053,N_36921,N_36984);
and U37054 (N_37054,N_36957,N_36971);
nor U37055 (N_37055,N_36928,N_36823);
nand U37056 (N_37056,N_36805,N_36813);
or U37057 (N_37057,N_36754,N_36821);
xor U37058 (N_37058,N_36998,N_36906);
or U37059 (N_37059,N_36914,N_36882);
and U37060 (N_37060,N_36943,N_36803);
nor U37061 (N_37061,N_36781,N_36953);
nand U37062 (N_37062,N_36806,N_36778);
nand U37063 (N_37063,N_36852,N_36925);
or U37064 (N_37064,N_36898,N_36854);
and U37065 (N_37065,N_36861,N_36804);
xnor U37066 (N_37066,N_36842,N_36792);
xnor U37067 (N_37067,N_36875,N_36893);
and U37068 (N_37068,N_36831,N_36800);
or U37069 (N_37069,N_36789,N_36929);
nor U37070 (N_37070,N_36876,N_36927);
nor U37071 (N_37071,N_36945,N_36847);
nor U37072 (N_37072,N_36862,N_36784);
xor U37073 (N_37073,N_36986,N_36811);
nor U37074 (N_37074,N_36851,N_36757);
and U37075 (N_37075,N_36982,N_36903);
xor U37076 (N_37076,N_36873,N_36979);
nand U37077 (N_37077,N_36894,N_36919);
or U37078 (N_37078,N_36907,N_36843);
and U37079 (N_37079,N_36920,N_36771);
and U37080 (N_37080,N_36935,N_36809);
nor U37081 (N_37081,N_36871,N_36901);
and U37082 (N_37082,N_36758,N_36828);
nand U37083 (N_37083,N_36967,N_36972);
or U37084 (N_37084,N_36890,N_36892);
nand U37085 (N_37085,N_36779,N_36850);
or U37086 (N_37086,N_36797,N_36849);
nor U37087 (N_37087,N_36913,N_36915);
nand U37088 (N_37088,N_36996,N_36891);
or U37089 (N_37089,N_36930,N_36833);
nand U37090 (N_37090,N_36923,N_36926);
xor U37091 (N_37091,N_36812,N_36829);
nand U37092 (N_37092,N_36790,N_36793);
nor U37093 (N_37093,N_36951,N_36755);
nand U37094 (N_37094,N_36908,N_36956);
nor U37095 (N_37095,N_36911,N_36902);
and U37096 (N_37096,N_36997,N_36955);
nor U37097 (N_37097,N_36839,N_36954);
xnor U37098 (N_37098,N_36932,N_36772);
nand U37099 (N_37099,N_36827,N_36773);
nand U37100 (N_37100,N_36868,N_36762);
and U37101 (N_37101,N_36966,N_36865);
xnor U37102 (N_37102,N_36880,N_36760);
xnor U37103 (N_37103,N_36949,N_36981);
and U37104 (N_37104,N_36917,N_36879);
xor U37105 (N_37105,N_36802,N_36939);
xnor U37106 (N_37106,N_36830,N_36889);
xor U37107 (N_37107,N_36782,N_36975);
xnor U37108 (N_37108,N_36768,N_36990);
xnor U37109 (N_37109,N_36948,N_36858);
nand U37110 (N_37110,N_36796,N_36810);
and U37111 (N_37111,N_36952,N_36766);
or U37112 (N_37112,N_36764,N_36999);
nand U37113 (N_37113,N_36856,N_36770);
nor U37114 (N_37114,N_36857,N_36841);
or U37115 (N_37115,N_36946,N_36769);
and U37116 (N_37116,N_36931,N_36822);
or U37117 (N_37117,N_36867,N_36947);
and U37118 (N_37118,N_36965,N_36874);
or U37119 (N_37119,N_36761,N_36848);
nand U37120 (N_37120,N_36970,N_36775);
nor U37121 (N_37121,N_36801,N_36836);
or U37122 (N_37122,N_36751,N_36786);
or U37123 (N_37123,N_36807,N_36870);
nor U37124 (N_37124,N_36964,N_36763);
nor U37125 (N_37125,N_36992,N_36751);
nand U37126 (N_37126,N_36817,N_36763);
nor U37127 (N_37127,N_36931,N_36932);
xor U37128 (N_37128,N_36806,N_36997);
xnor U37129 (N_37129,N_36948,N_36836);
or U37130 (N_37130,N_36967,N_36780);
xnor U37131 (N_37131,N_36892,N_36820);
and U37132 (N_37132,N_36900,N_36987);
nand U37133 (N_37133,N_36895,N_36759);
or U37134 (N_37134,N_36850,N_36797);
nor U37135 (N_37135,N_36758,N_36964);
nor U37136 (N_37136,N_36995,N_36866);
xnor U37137 (N_37137,N_36911,N_36775);
nand U37138 (N_37138,N_36857,N_36916);
nand U37139 (N_37139,N_36818,N_36813);
or U37140 (N_37140,N_36904,N_36823);
or U37141 (N_37141,N_36834,N_36910);
xor U37142 (N_37142,N_36921,N_36882);
xnor U37143 (N_37143,N_36844,N_36882);
nor U37144 (N_37144,N_36874,N_36897);
nand U37145 (N_37145,N_36937,N_36898);
nand U37146 (N_37146,N_36853,N_36816);
nor U37147 (N_37147,N_36793,N_36945);
and U37148 (N_37148,N_36904,N_36947);
nand U37149 (N_37149,N_36770,N_36769);
nor U37150 (N_37150,N_36858,N_36958);
xor U37151 (N_37151,N_36973,N_36834);
xor U37152 (N_37152,N_36996,N_36890);
and U37153 (N_37153,N_36962,N_36754);
nand U37154 (N_37154,N_36851,N_36830);
nor U37155 (N_37155,N_36790,N_36846);
xor U37156 (N_37156,N_36761,N_36933);
xor U37157 (N_37157,N_36769,N_36798);
nand U37158 (N_37158,N_36878,N_36936);
and U37159 (N_37159,N_36865,N_36910);
or U37160 (N_37160,N_36757,N_36824);
nor U37161 (N_37161,N_36902,N_36875);
or U37162 (N_37162,N_36895,N_36947);
and U37163 (N_37163,N_36808,N_36975);
and U37164 (N_37164,N_36867,N_36963);
and U37165 (N_37165,N_36752,N_36871);
nand U37166 (N_37166,N_36839,N_36914);
nor U37167 (N_37167,N_36949,N_36986);
nor U37168 (N_37168,N_36916,N_36754);
nand U37169 (N_37169,N_36955,N_36809);
nor U37170 (N_37170,N_36907,N_36756);
and U37171 (N_37171,N_36755,N_36991);
nand U37172 (N_37172,N_36833,N_36851);
nor U37173 (N_37173,N_36798,N_36941);
nor U37174 (N_37174,N_36844,N_36991);
and U37175 (N_37175,N_36766,N_36759);
xor U37176 (N_37176,N_36808,N_36909);
nor U37177 (N_37177,N_36876,N_36895);
or U37178 (N_37178,N_36854,N_36998);
or U37179 (N_37179,N_36990,N_36978);
nand U37180 (N_37180,N_36814,N_36885);
nor U37181 (N_37181,N_36764,N_36822);
nor U37182 (N_37182,N_36898,N_36873);
xor U37183 (N_37183,N_36876,N_36753);
nand U37184 (N_37184,N_36983,N_36865);
nor U37185 (N_37185,N_36757,N_36778);
and U37186 (N_37186,N_36947,N_36957);
xnor U37187 (N_37187,N_36973,N_36846);
xnor U37188 (N_37188,N_36931,N_36831);
xor U37189 (N_37189,N_36814,N_36757);
xnor U37190 (N_37190,N_36750,N_36851);
xnor U37191 (N_37191,N_36996,N_36924);
xor U37192 (N_37192,N_36878,N_36955);
xor U37193 (N_37193,N_36821,N_36849);
and U37194 (N_37194,N_36832,N_36862);
nor U37195 (N_37195,N_36934,N_36914);
or U37196 (N_37196,N_36998,N_36959);
or U37197 (N_37197,N_36914,N_36848);
or U37198 (N_37198,N_36927,N_36934);
nor U37199 (N_37199,N_36761,N_36949);
nor U37200 (N_37200,N_36984,N_36970);
and U37201 (N_37201,N_36980,N_36826);
xor U37202 (N_37202,N_36872,N_36919);
or U37203 (N_37203,N_36776,N_36965);
and U37204 (N_37204,N_36849,N_36869);
nor U37205 (N_37205,N_36840,N_36962);
and U37206 (N_37206,N_36884,N_36989);
xnor U37207 (N_37207,N_36935,N_36922);
nor U37208 (N_37208,N_36939,N_36888);
xor U37209 (N_37209,N_36782,N_36762);
xnor U37210 (N_37210,N_36949,N_36859);
nand U37211 (N_37211,N_36949,N_36970);
nor U37212 (N_37212,N_36964,N_36777);
nand U37213 (N_37213,N_36838,N_36778);
xnor U37214 (N_37214,N_36796,N_36853);
xor U37215 (N_37215,N_36850,N_36916);
nand U37216 (N_37216,N_36807,N_36842);
nand U37217 (N_37217,N_36755,N_36896);
or U37218 (N_37218,N_36850,N_36982);
nand U37219 (N_37219,N_36795,N_36777);
and U37220 (N_37220,N_36753,N_36917);
nor U37221 (N_37221,N_36868,N_36878);
and U37222 (N_37222,N_36797,N_36832);
or U37223 (N_37223,N_36859,N_36818);
xnor U37224 (N_37224,N_36929,N_36953);
nor U37225 (N_37225,N_36914,N_36915);
nor U37226 (N_37226,N_36756,N_36819);
xor U37227 (N_37227,N_36970,N_36803);
and U37228 (N_37228,N_36848,N_36760);
and U37229 (N_37229,N_36769,N_36991);
xnor U37230 (N_37230,N_36999,N_36987);
xnor U37231 (N_37231,N_36970,N_36988);
xnor U37232 (N_37232,N_36965,N_36959);
and U37233 (N_37233,N_36832,N_36769);
and U37234 (N_37234,N_36869,N_36978);
or U37235 (N_37235,N_36921,N_36797);
or U37236 (N_37236,N_36820,N_36835);
nand U37237 (N_37237,N_36855,N_36756);
nand U37238 (N_37238,N_36797,N_36990);
and U37239 (N_37239,N_36930,N_36787);
nor U37240 (N_37240,N_36804,N_36957);
and U37241 (N_37241,N_36785,N_36953);
xor U37242 (N_37242,N_36804,N_36874);
and U37243 (N_37243,N_36907,N_36776);
nor U37244 (N_37244,N_36905,N_36902);
nand U37245 (N_37245,N_36845,N_36752);
and U37246 (N_37246,N_36867,N_36862);
xnor U37247 (N_37247,N_36839,N_36887);
nor U37248 (N_37248,N_36836,N_36953);
or U37249 (N_37249,N_36788,N_36862);
or U37250 (N_37250,N_37070,N_37056);
xor U37251 (N_37251,N_37100,N_37052);
nor U37252 (N_37252,N_37242,N_37075);
xor U37253 (N_37253,N_37117,N_37144);
or U37254 (N_37254,N_37103,N_37164);
or U37255 (N_37255,N_37219,N_37235);
nand U37256 (N_37256,N_37028,N_37087);
nand U37257 (N_37257,N_37107,N_37138);
or U37258 (N_37258,N_37233,N_37132);
and U37259 (N_37259,N_37048,N_37083);
or U37260 (N_37260,N_37158,N_37031);
nand U37261 (N_37261,N_37029,N_37224);
and U37262 (N_37262,N_37163,N_37039);
xor U37263 (N_37263,N_37012,N_37054);
xor U37264 (N_37264,N_37035,N_37215);
or U37265 (N_37265,N_37025,N_37232);
and U37266 (N_37266,N_37033,N_37049);
and U37267 (N_37267,N_37245,N_37106);
nand U37268 (N_37268,N_37178,N_37135);
and U37269 (N_37269,N_37032,N_37124);
nor U37270 (N_37270,N_37131,N_37184);
nand U37271 (N_37271,N_37197,N_37244);
and U37272 (N_37272,N_37228,N_37162);
and U37273 (N_37273,N_37059,N_37072);
nand U37274 (N_37274,N_37222,N_37081);
nand U37275 (N_37275,N_37129,N_37113);
and U37276 (N_37276,N_37071,N_37088);
and U37277 (N_37277,N_37201,N_37002);
nor U37278 (N_37278,N_37140,N_37217);
xnor U37279 (N_37279,N_37120,N_37213);
xor U37280 (N_37280,N_37154,N_37016);
xor U37281 (N_37281,N_37202,N_37063);
nor U37282 (N_37282,N_37209,N_37148);
nand U37283 (N_37283,N_37168,N_37125);
nor U37284 (N_37284,N_37171,N_37069);
nor U37285 (N_37285,N_37000,N_37192);
nand U37286 (N_37286,N_37108,N_37210);
xor U37287 (N_37287,N_37142,N_37079);
xor U37288 (N_37288,N_37119,N_37118);
and U37289 (N_37289,N_37018,N_37225);
xnor U37290 (N_37290,N_37045,N_37150);
nor U37291 (N_37291,N_37001,N_37145);
and U37292 (N_37292,N_37247,N_37127);
nor U37293 (N_37293,N_37173,N_37064);
and U37294 (N_37294,N_37169,N_37157);
and U37295 (N_37295,N_37199,N_37237);
nor U37296 (N_37296,N_37159,N_37006);
nor U37297 (N_37297,N_37166,N_37139);
nand U37298 (N_37298,N_37037,N_37080);
nor U37299 (N_37299,N_37076,N_37165);
xor U37300 (N_37300,N_37229,N_37218);
nor U37301 (N_37301,N_37023,N_37122);
xnor U37302 (N_37302,N_37147,N_37126);
nor U37303 (N_37303,N_37022,N_37236);
xor U37304 (N_37304,N_37114,N_37143);
nor U37305 (N_37305,N_37011,N_37067);
xnor U37306 (N_37306,N_37065,N_37151);
nor U37307 (N_37307,N_37093,N_37047);
nand U37308 (N_37308,N_37051,N_37026);
and U37309 (N_37309,N_37085,N_37249);
nand U37310 (N_37310,N_37188,N_37130);
nand U37311 (N_37311,N_37152,N_37221);
or U37312 (N_37312,N_37111,N_37013);
nor U37313 (N_37313,N_37073,N_37161);
nor U37314 (N_37314,N_37090,N_37094);
xor U37315 (N_37315,N_37101,N_37053);
and U37316 (N_37316,N_37041,N_37021);
and U37317 (N_37317,N_37238,N_37212);
xor U37318 (N_37318,N_37243,N_37050);
nor U37319 (N_37319,N_37102,N_37226);
xor U37320 (N_37320,N_37077,N_37198);
xor U37321 (N_37321,N_37007,N_37057);
nor U37322 (N_37322,N_37177,N_37099);
and U37323 (N_37323,N_37089,N_37155);
nand U37324 (N_37324,N_37128,N_37206);
xnor U37325 (N_37325,N_37084,N_37030);
and U37326 (N_37326,N_37167,N_37172);
or U37327 (N_37327,N_37149,N_37146);
and U37328 (N_37328,N_37020,N_37234);
nand U37329 (N_37329,N_37193,N_37156);
nor U37330 (N_37330,N_37121,N_37066);
and U37331 (N_37331,N_37204,N_37207);
nand U37332 (N_37332,N_37136,N_37082);
nand U37333 (N_37333,N_37019,N_37104);
or U37334 (N_37334,N_37017,N_37185);
xor U37335 (N_37335,N_37015,N_37086);
or U37336 (N_37336,N_37196,N_37174);
and U37337 (N_37337,N_37240,N_37134);
nand U37338 (N_37338,N_37061,N_37110);
nor U37339 (N_37339,N_37040,N_37211);
xor U37340 (N_37340,N_37034,N_37068);
or U37341 (N_37341,N_37182,N_37008);
nand U37342 (N_37342,N_37180,N_37055);
nand U37343 (N_37343,N_37176,N_37208);
and U37344 (N_37344,N_37246,N_37115);
and U37345 (N_37345,N_37241,N_37004);
nand U37346 (N_37346,N_37230,N_37187);
or U37347 (N_37347,N_37060,N_37074);
nand U37348 (N_37348,N_37248,N_37205);
and U37349 (N_37349,N_37014,N_37186);
or U37350 (N_37350,N_37191,N_37195);
xnor U37351 (N_37351,N_37046,N_37098);
xor U37352 (N_37352,N_37216,N_37058);
nor U37353 (N_37353,N_37181,N_37116);
nand U37354 (N_37354,N_37096,N_37189);
nand U37355 (N_37355,N_37123,N_37231);
nor U37356 (N_37356,N_37112,N_37179);
nand U37357 (N_37357,N_37036,N_37062);
nor U37358 (N_37358,N_37009,N_37097);
nand U37359 (N_37359,N_37170,N_37109);
xor U37360 (N_37360,N_37137,N_37175);
or U37361 (N_37361,N_37078,N_37003);
nor U37362 (N_37362,N_37044,N_37141);
and U37363 (N_37363,N_37153,N_37223);
and U37364 (N_37364,N_37214,N_37095);
and U37365 (N_37365,N_37227,N_37194);
or U37366 (N_37366,N_37203,N_37010);
nand U37367 (N_37367,N_37005,N_37105);
xor U37368 (N_37368,N_37092,N_37239);
xor U37369 (N_37369,N_37200,N_37183);
xor U37370 (N_37370,N_37133,N_37160);
nor U37371 (N_37371,N_37190,N_37043);
nor U37372 (N_37372,N_37042,N_37027);
xor U37373 (N_37373,N_37220,N_37024);
and U37374 (N_37374,N_37038,N_37091);
nor U37375 (N_37375,N_37236,N_37187);
and U37376 (N_37376,N_37155,N_37000);
or U37377 (N_37377,N_37170,N_37180);
and U37378 (N_37378,N_37200,N_37213);
nor U37379 (N_37379,N_37023,N_37149);
nand U37380 (N_37380,N_37099,N_37164);
xnor U37381 (N_37381,N_37041,N_37122);
nand U37382 (N_37382,N_37232,N_37242);
or U37383 (N_37383,N_37057,N_37245);
and U37384 (N_37384,N_37124,N_37197);
or U37385 (N_37385,N_37154,N_37096);
xor U37386 (N_37386,N_37160,N_37140);
xor U37387 (N_37387,N_37226,N_37113);
nand U37388 (N_37388,N_37148,N_37201);
nand U37389 (N_37389,N_37006,N_37099);
and U37390 (N_37390,N_37162,N_37201);
or U37391 (N_37391,N_37015,N_37143);
and U37392 (N_37392,N_37185,N_37060);
nand U37393 (N_37393,N_37024,N_37014);
or U37394 (N_37394,N_37166,N_37220);
nor U37395 (N_37395,N_37180,N_37203);
nand U37396 (N_37396,N_37190,N_37224);
or U37397 (N_37397,N_37241,N_37172);
nor U37398 (N_37398,N_37246,N_37043);
nand U37399 (N_37399,N_37114,N_37195);
or U37400 (N_37400,N_37152,N_37000);
or U37401 (N_37401,N_37240,N_37064);
and U37402 (N_37402,N_37191,N_37219);
nor U37403 (N_37403,N_37191,N_37152);
nor U37404 (N_37404,N_37137,N_37214);
nand U37405 (N_37405,N_37246,N_37207);
xnor U37406 (N_37406,N_37015,N_37002);
xnor U37407 (N_37407,N_37046,N_37107);
xnor U37408 (N_37408,N_37064,N_37202);
and U37409 (N_37409,N_37129,N_37016);
and U37410 (N_37410,N_37129,N_37026);
nor U37411 (N_37411,N_37120,N_37018);
nor U37412 (N_37412,N_37004,N_37016);
xnor U37413 (N_37413,N_37241,N_37097);
nor U37414 (N_37414,N_37081,N_37243);
and U37415 (N_37415,N_37024,N_37093);
and U37416 (N_37416,N_37242,N_37191);
nand U37417 (N_37417,N_37025,N_37151);
nand U37418 (N_37418,N_37192,N_37138);
and U37419 (N_37419,N_37088,N_37213);
nor U37420 (N_37420,N_37052,N_37049);
nand U37421 (N_37421,N_37062,N_37087);
or U37422 (N_37422,N_37034,N_37222);
or U37423 (N_37423,N_37117,N_37035);
xor U37424 (N_37424,N_37071,N_37019);
xor U37425 (N_37425,N_37167,N_37033);
xnor U37426 (N_37426,N_37077,N_37188);
xor U37427 (N_37427,N_37007,N_37019);
nand U37428 (N_37428,N_37117,N_37053);
and U37429 (N_37429,N_37198,N_37236);
nor U37430 (N_37430,N_37111,N_37238);
nand U37431 (N_37431,N_37234,N_37105);
nand U37432 (N_37432,N_37144,N_37098);
or U37433 (N_37433,N_37045,N_37194);
or U37434 (N_37434,N_37242,N_37205);
and U37435 (N_37435,N_37045,N_37073);
nor U37436 (N_37436,N_37249,N_37164);
xor U37437 (N_37437,N_37185,N_37069);
nand U37438 (N_37438,N_37016,N_37003);
nor U37439 (N_37439,N_37006,N_37038);
or U37440 (N_37440,N_37023,N_37093);
and U37441 (N_37441,N_37146,N_37001);
and U37442 (N_37442,N_37127,N_37082);
or U37443 (N_37443,N_37241,N_37134);
or U37444 (N_37444,N_37030,N_37249);
and U37445 (N_37445,N_37099,N_37102);
or U37446 (N_37446,N_37194,N_37027);
and U37447 (N_37447,N_37192,N_37145);
nand U37448 (N_37448,N_37191,N_37001);
nand U37449 (N_37449,N_37245,N_37054);
nor U37450 (N_37450,N_37063,N_37114);
nand U37451 (N_37451,N_37065,N_37059);
xnor U37452 (N_37452,N_37109,N_37110);
or U37453 (N_37453,N_37123,N_37184);
or U37454 (N_37454,N_37068,N_37060);
and U37455 (N_37455,N_37014,N_37190);
nor U37456 (N_37456,N_37140,N_37075);
or U37457 (N_37457,N_37212,N_37243);
or U37458 (N_37458,N_37201,N_37070);
nand U37459 (N_37459,N_37012,N_37177);
or U37460 (N_37460,N_37163,N_37159);
nor U37461 (N_37461,N_37243,N_37113);
nand U37462 (N_37462,N_37189,N_37190);
nor U37463 (N_37463,N_37086,N_37210);
nand U37464 (N_37464,N_37194,N_37225);
nand U37465 (N_37465,N_37199,N_37221);
xor U37466 (N_37466,N_37144,N_37243);
nand U37467 (N_37467,N_37085,N_37033);
and U37468 (N_37468,N_37098,N_37167);
and U37469 (N_37469,N_37121,N_37207);
nor U37470 (N_37470,N_37225,N_37165);
nand U37471 (N_37471,N_37056,N_37125);
nand U37472 (N_37472,N_37073,N_37007);
xor U37473 (N_37473,N_37161,N_37177);
nand U37474 (N_37474,N_37062,N_37064);
or U37475 (N_37475,N_37125,N_37030);
nor U37476 (N_37476,N_37148,N_37089);
and U37477 (N_37477,N_37026,N_37180);
or U37478 (N_37478,N_37050,N_37127);
or U37479 (N_37479,N_37095,N_37161);
xor U37480 (N_37480,N_37035,N_37012);
nor U37481 (N_37481,N_37180,N_37161);
nor U37482 (N_37482,N_37094,N_37133);
and U37483 (N_37483,N_37107,N_37170);
and U37484 (N_37484,N_37074,N_37216);
xnor U37485 (N_37485,N_37048,N_37061);
nand U37486 (N_37486,N_37138,N_37244);
xor U37487 (N_37487,N_37166,N_37188);
and U37488 (N_37488,N_37030,N_37208);
nand U37489 (N_37489,N_37087,N_37060);
nand U37490 (N_37490,N_37134,N_37158);
or U37491 (N_37491,N_37202,N_37086);
xor U37492 (N_37492,N_37183,N_37054);
and U37493 (N_37493,N_37155,N_37238);
and U37494 (N_37494,N_37189,N_37126);
xor U37495 (N_37495,N_37036,N_37181);
xor U37496 (N_37496,N_37090,N_37074);
nand U37497 (N_37497,N_37245,N_37182);
and U37498 (N_37498,N_37210,N_37127);
and U37499 (N_37499,N_37129,N_37230);
nand U37500 (N_37500,N_37375,N_37455);
xnor U37501 (N_37501,N_37328,N_37495);
and U37502 (N_37502,N_37301,N_37361);
nor U37503 (N_37503,N_37349,N_37331);
nor U37504 (N_37504,N_37496,N_37400);
xor U37505 (N_37505,N_37329,N_37364);
or U37506 (N_37506,N_37406,N_37438);
or U37507 (N_37507,N_37293,N_37326);
or U37508 (N_37508,N_37482,N_37353);
and U37509 (N_37509,N_37294,N_37436);
or U37510 (N_37510,N_37378,N_37255);
and U37511 (N_37511,N_37466,N_37464);
or U37512 (N_37512,N_37412,N_37467);
nor U37513 (N_37513,N_37420,N_37333);
nand U37514 (N_37514,N_37262,N_37315);
xnor U37515 (N_37515,N_37290,N_37252);
and U37516 (N_37516,N_37368,N_37308);
nand U37517 (N_37517,N_37469,N_37471);
nand U37518 (N_37518,N_37377,N_37426);
or U37519 (N_37519,N_37254,N_37295);
nor U37520 (N_37520,N_37320,N_37384);
or U37521 (N_37521,N_37306,N_37338);
nor U37522 (N_37522,N_37260,N_37419);
nor U37523 (N_37523,N_37473,N_37323);
xor U37524 (N_37524,N_37360,N_37451);
and U37525 (N_37525,N_37437,N_37314);
and U37526 (N_37526,N_37444,N_37448);
nand U37527 (N_37527,N_37282,N_37281);
xnor U37528 (N_37528,N_37393,N_37433);
nand U37529 (N_37529,N_37459,N_37408);
or U37530 (N_37530,N_37413,N_37371);
nor U37531 (N_37531,N_37257,N_37457);
nand U37532 (N_37532,N_37407,N_37280);
nand U37533 (N_37533,N_37454,N_37379);
nor U37534 (N_37534,N_37449,N_37380);
nor U37535 (N_37535,N_37298,N_37267);
or U37536 (N_37536,N_37268,N_37477);
xnor U37537 (N_37537,N_37345,N_37374);
xnor U37538 (N_37538,N_37428,N_37472);
nand U37539 (N_37539,N_37296,N_37358);
nor U37540 (N_37540,N_37327,N_37346);
nand U37541 (N_37541,N_37418,N_37264);
and U37542 (N_37542,N_37283,N_37404);
nor U37543 (N_37543,N_37439,N_37499);
nor U37544 (N_37544,N_37305,N_37410);
nand U37545 (N_37545,N_37429,N_37337);
nand U37546 (N_37546,N_37387,N_37250);
nand U37547 (N_37547,N_37494,N_37480);
nand U37548 (N_37548,N_37271,N_37340);
nand U37549 (N_37549,N_37299,N_37417);
nor U37550 (N_37550,N_37334,N_37415);
xor U37551 (N_37551,N_37251,N_37356);
or U37552 (N_37552,N_37311,N_37497);
nor U37553 (N_37553,N_37365,N_37392);
nand U37554 (N_37554,N_37395,N_37276);
xor U37555 (N_37555,N_37288,N_37265);
nand U37556 (N_37556,N_37493,N_37475);
nor U37557 (N_37557,N_37352,N_37285);
or U37558 (N_37558,N_37273,N_37453);
and U37559 (N_37559,N_37432,N_37287);
xor U37560 (N_37560,N_37302,N_37350);
nor U37561 (N_37561,N_37339,N_37385);
nand U37562 (N_37562,N_37431,N_37391);
and U37563 (N_37563,N_37357,N_37401);
nand U37564 (N_37564,N_37492,N_37484);
or U37565 (N_37565,N_37304,N_37458);
xnor U37566 (N_37566,N_37351,N_37373);
nor U37567 (N_37567,N_37465,N_37354);
or U37568 (N_37568,N_37403,N_37479);
or U37569 (N_37569,N_37263,N_37489);
and U37570 (N_37570,N_37383,N_37394);
xnor U37571 (N_37571,N_37388,N_37313);
and U37572 (N_37572,N_37303,N_37452);
or U37573 (N_37573,N_37463,N_37409);
nor U37574 (N_37574,N_37261,N_37474);
or U37575 (N_37575,N_37319,N_37462);
or U37576 (N_37576,N_37427,N_37456);
or U37577 (N_37577,N_37485,N_37416);
and U37578 (N_37578,N_37498,N_37275);
and U37579 (N_37579,N_37366,N_37470);
or U37580 (N_37580,N_37289,N_37478);
nor U37581 (N_37581,N_37277,N_37317);
xor U37582 (N_37582,N_37381,N_37335);
or U37583 (N_37583,N_37341,N_37443);
and U37584 (N_37584,N_37310,N_37291);
nand U37585 (N_37585,N_37256,N_37272);
and U37586 (N_37586,N_37278,N_37445);
and U37587 (N_37587,N_37367,N_37397);
nor U37588 (N_37588,N_37336,N_37423);
nand U37589 (N_37589,N_37363,N_37425);
or U37590 (N_37590,N_37396,N_37332);
nand U37591 (N_37591,N_37434,N_37279);
xor U37592 (N_37592,N_37269,N_37390);
xnor U37593 (N_37593,N_37405,N_37370);
or U37594 (N_37594,N_37322,N_37481);
nor U37595 (N_37595,N_37316,N_37490);
xnor U37596 (N_37596,N_37258,N_37421);
or U37597 (N_37597,N_37372,N_37292);
nand U37598 (N_37598,N_37286,N_37422);
nand U37599 (N_37599,N_37330,N_37284);
xor U37600 (N_37600,N_37460,N_37450);
and U37601 (N_37601,N_37430,N_37446);
nand U37602 (N_37602,N_37348,N_37487);
nand U37603 (N_37603,N_37447,N_37362);
nand U37604 (N_37604,N_37398,N_37325);
and U37605 (N_37605,N_37355,N_37376);
or U37606 (N_37606,N_37347,N_37491);
or U37607 (N_37607,N_37386,N_37402);
xnor U37608 (N_37608,N_37435,N_37369);
nor U37609 (N_37609,N_37344,N_37440);
or U37610 (N_37610,N_37461,N_37476);
xor U37611 (N_37611,N_37342,N_37259);
nand U37612 (N_37612,N_37266,N_37324);
and U37613 (N_37613,N_37442,N_37488);
or U37614 (N_37614,N_37486,N_37270);
nand U37615 (N_37615,N_37321,N_37441);
and U37616 (N_37616,N_37318,N_37297);
nand U37617 (N_37617,N_37389,N_37411);
and U37618 (N_37618,N_37382,N_37414);
nand U37619 (N_37619,N_37253,N_37307);
nor U37620 (N_37620,N_37312,N_37300);
xor U37621 (N_37621,N_37399,N_37343);
and U37622 (N_37622,N_37309,N_37468);
or U37623 (N_37623,N_37424,N_37359);
nor U37624 (N_37624,N_37274,N_37483);
or U37625 (N_37625,N_37329,N_37432);
and U37626 (N_37626,N_37491,N_37355);
nand U37627 (N_37627,N_37334,N_37314);
or U37628 (N_37628,N_37383,N_37333);
nand U37629 (N_37629,N_37496,N_37267);
or U37630 (N_37630,N_37450,N_37486);
xnor U37631 (N_37631,N_37429,N_37433);
nor U37632 (N_37632,N_37383,N_37389);
nor U37633 (N_37633,N_37254,N_37414);
xnor U37634 (N_37634,N_37268,N_37464);
and U37635 (N_37635,N_37463,N_37475);
and U37636 (N_37636,N_37389,N_37452);
or U37637 (N_37637,N_37270,N_37481);
or U37638 (N_37638,N_37472,N_37371);
xor U37639 (N_37639,N_37454,N_37425);
xor U37640 (N_37640,N_37290,N_37378);
xnor U37641 (N_37641,N_37490,N_37499);
nand U37642 (N_37642,N_37437,N_37495);
nor U37643 (N_37643,N_37343,N_37494);
or U37644 (N_37644,N_37415,N_37389);
nor U37645 (N_37645,N_37429,N_37346);
nor U37646 (N_37646,N_37384,N_37460);
and U37647 (N_37647,N_37311,N_37436);
xnor U37648 (N_37648,N_37339,N_37250);
and U37649 (N_37649,N_37327,N_37382);
nand U37650 (N_37650,N_37430,N_37331);
nand U37651 (N_37651,N_37378,N_37431);
or U37652 (N_37652,N_37397,N_37361);
and U37653 (N_37653,N_37480,N_37342);
nand U37654 (N_37654,N_37335,N_37256);
nand U37655 (N_37655,N_37301,N_37378);
nand U37656 (N_37656,N_37356,N_37299);
nor U37657 (N_37657,N_37422,N_37434);
and U37658 (N_37658,N_37310,N_37280);
nor U37659 (N_37659,N_37464,N_37294);
and U37660 (N_37660,N_37251,N_37282);
or U37661 (N_37661,N_37375,N_37298);
or U37662 (N_37662,N_37275,N_37370);
and U37663 (N_37663,N_37389,N_37356);
and U37664 (N_37664,N_37268,N_37379);
nor U37665 (N_37665,N_37466,N_37499);
nand U37666 (N_37666,N_37250,N_37400);
and U37667 (N_37667,N_37368,N_37465);
xor U37668 (N_37668,N_37443,N_37253);
nand U37669 (N_37669,N_37264,N_37490);
or U37670 (N_37670,N_37448,N_37301);
and U37671 (N_37671,N_37452,N_37349);
xor U37672 (N_37672,N_37463,N_37359);
nand U37673 (N_37673,N_37326,N_37496);
or U37674 (N_37674,N_37274,N_37337);
nor U37675 (N_37675,N_37450,N_37359);
or U37676 (N_37676,N_37253,N_37457);
nor U37677 (N_37677,N_37390,N_37332);
or U37678 (N_37678,N_37354,N_37455);
or U37679 (N_37679,N_37417,N_37454);
xor U37680 (N_37680,N_37356,N_37454);
or U37681 (N_37681,N_37250,N_37472);
or U37682 (N_37682,N_37462,N_37266);
or U37683 (N_37683,N_37301,N_37475);
nand U37684 (N_37684,N_37498,N_37465);
or U37685 (N_37685,N_37280,N_37413);
xor U37686 (N_37686,N_37412,N_37464);
or U37687 (N_37687,N_37397,N_37434);
xnor U37688 (N_37688,N_37463,N_37295);
nor U37689 (N_37689,N_37489,N_37476);
nor U37690 (N_37690,N_37300,N_37486);
nor U37691 (N_37691,N_37415,N_37395);
or U37692 (N_37692,N_37298,N_37401);
xor U37693 (N_37693,N_37350,N_37282);
and U37694 (N_37694,N_37325,N_37344);
xor U37695 (N_37695,N_37493,N_37435);
or U37696 (N_37696,N_37309,N_37338);
xnor U37697 (N_37697,N_37330,N_37261);
nor U37698 (N_37698,N_37393,N_37289);
xnor U37699 (N_37699,N_37345,N_37297);
nand U37700 (N_37700,N_37313,N_37422);
and U37701 (N_37701,N_37499,N_37401);
nor U37702 (N_37702,N_37424,N_37356);
and U37703 (N_37703,N_37444,N_37362);
or U37704 (N_37704,N_37368,N_37437);
nor U37705 (N_37705,N_37355,N_37368);
or U37706 (N_37706,N_37263,N_37271);
or U37707 (N_37707,N_37374,N_37389);
or U37708 (N_37708,N_37489,N_37340);
xor U37709 (N_37709,N_37491,N_37340);
or U37710 (N_37710,N_37306,N_37274);
or U37711 (N_37711,N_37324,N_37485);
or U37712 (N_37712,N_37299,N_37272);
and U37713 (N_37713,N_37261,N_37419);
nand U37714 (N_37714,N_37346,N_37303);
xnor U37715 (N_37715,N_37373,N_37496);
nor U37716 (N_37716,N_37319,N_37373);
or U37717 (N_37717,N_37367,N_37338);
nand U37718 (N_37718,N_37266,N_37489);
or U37719 (N_37719,N_37475,N_37497);
xnor U37720 (N_37720,N_37324,N_37429);
xnor U37721 (N_37721,N_37377,N_37360);
and U37722 (N_37722,N_37335,N_37333);
and U37723 (N_37723,N_37319,N_37445);
nor U37724 (N_37724,N_37498,N_37329);
nand U37725 (N_37725,N_37485,N_37418);
xnor U37726 (N_37726,N_37493,N_37469);
and U37727 (N_37727,N_37412,N_37455);
nor U37728 (N_37728,N_37271,N_37261);
or U37729 (N_37729,N_37251,N_37441);
nor U37730 (N_37730,N_37396,N_37417);
nand U37731 (N_37731,N_37374,N_37356);
or U37732 (N_37732,N_37409,N_37334);
and U37733 (N_37733,N_37485,N_37356);
and U37734 (N_37734,N_37354,N_37261);
nand U37735 (N_37735,N_37470,N_37298);
and U37736 (N_37736,N_37285,N_37355);
nand U37737 (N_37737,N_37472,N_37410);
xor U37738 (N_37738,N_37398,N_37452);
and U37739 (N_37739,N_37495,N_37459);
nand U37740 (N_37740,N_37374,N_37299);
xnor U37741 (N_37741,N_37307,N_37314);
xor U37742 (N_37742,N_37394,N_37389);
nor U37743 (N_37743,N_37478,N_37376);
xnor U37744 (N_37744,N_37467,N_37317);
nand U37745 (N_37745,N_37307,N_37468);
and U37746 (N_37746,N_37376,N_37405);
or U37747 (N_37747,N_37266,N_37356);
nor U37748 (N_37748,N_37455,N_37268);
nor U37749 (N_37749,N_37353,N_37362);
or U37750 (N_37750,N_37636,N_37582);
and U37751 (N_37751,N_37691,N_37700);
nand U37752 (N_37752,N_37514,N_37697);
nor U37753 (N_37753,N_37508,N_37506);
xnor U37754 (N_37754,N_37567,N_37629);
and U37755 (N_37755,N_37686,N_37673);
xnor U37756 (N_37756,N_37647,N_37665);
or U37757 (N_37757,N_37648,N_37724);
xnor U37758 (N_37758,N_37618,N_37745);
or U37759 (N_37759,N_37694,N_37692);
xnor U37760 (N_37760,N_37736,N_37573);
nand U37761 (N_37761,N_37703,N_37596);
and U37762 (N_37762,N_37619,N_37728);
and U37763 (N_37763,N_37502,N_37590);
or U37764 (N_37764,N_37706,N_37599);
or U37765 (N_37765,N_37655,N_37680);
or U37766 (N_37766,N_37747,N_37537);
nand U37767 (N_37767,N_37646,N_37543);
and U37768 (N_37768,N_37575,N_37683);
nand U37769 (N_37769,N_37589,N_37504);
and U37770 (N_37770,N_37663,N_37632);
nor U37771 (N_37771,N_37684,N_37524);
nor U37772 (N_37772,N_37592,N_37718);
nand U37773 (N_37773,N_37723,N_37733);
and U37774 (N_37774,N_37546,N_37651);
or U37775 (N_37775,N_37642,N_37563);
nand U37776 (N_37776,N_37610,N_37695);
and U37777 (N_37777,N_37679,N_37612);
or U37778 (N_37778,N_37699,N_37607);
xnor U37779 (N_37779,N_37572,N_37539);
or U37780 (N_37780,N_37501,N_37657);
xnor U37781 (N_37781,N_37737,N_37523);
xnor U37782 (N_37782,N_37507,N_37581);
and U37783 (N_37783,N_37637,N_37743);
nand U37784 (N_37784,N_37711,N_37565);
nand U37785 (N_37785,N_37740,N_37656);
xor U37786 (N_37786,N_37661,N_37588);
xor U37787 (N_37787,N_37533,N_37583);
nand U37788 (N_37788,N_37513,N_37519);
nor U37789 (N_37789,N_37571,N_37535);
xnor U37790 (N_37790,N_37649,N_37662);
or U37791 (N_37791,N_37639,N_37542);
or U37792 (N_37792,N_37585,N_37698);
or U37793 (N_37793,N_37515,N_37666);
nor U37794 (N_37794,N_37731,N_37749);
nor U37795 (N_37795,N_37628,N_37682);
xor U37796 (N_37796,N_37712,N_37630);
or U37797 (N_37797,N_37652,N_37702);
xor U37798 (N_37798,N_37552,N_37744);
or U37799 (N_37799,N_37742,N_37602);
nand U37800 (N_37800,N_37569,N_37560);
xor U37801 (N_37801,N_37709,N_37633);
or U37802 (N_37802,N_37503,N_37584);
nor U37803 (N_37803,N_37708,N_37696);
and U37804 (N_37804,N_37739,N_37681);
xor U37805 (N_37805,N_37600,N_37645);
or U37806 (N_37806,N_37517,N_37556);
nand U37807 (N_37807,N_37644,N_37601);
or U37808 (N_37808,N_37704,N_37500);
nand U37809 (N_37809,N_37613,N_37541);
or U37810 (N_37810,N_37561,N_37606);
nor U37811 (N_37811,N_37605,N_37677);
nand U37812 (N_37812,N_37748,N_37604);
or U37813 (N_37813,N_37641,N_37593);
or U37814 (N_37814,N_37650,N_37669);
nand U37815 (N_37815,N_37532,N_37623);
xnor U37816 (N_37816,N_37522,N_37531);
and U37817 (N_37817,N_37653,N_37530);
and U37818 (N_37818,N_37550,N_37527);
nand U37819 (N_37819,N_37621,N_37591);
nand U37820 (N_37820,N_37576,N_37587);
and U37821 (N_37821,N_37689,N_37638);
nand U37822 (N_37822,N_37511,N_37735);
and U37823 (N_37823,N_37518,N_37544);
nor U37824 (N_37824,N_37741,N_37634);
nand U37825 (N_37825,N_37617,N_37554);
nor U37826 (N_37826,N_37658,N_37719);
xor U37827 (N_37827,N_37597,N_37526);
or U37828 (N_37828,N_37534,N_37667);
xnor U37829 (N_37829,N_37727,N_37670);
or U37830 (N_37830,N_37674,N_37562);
xnor U37831 (N_37831,N_37675,N_37640);
xnor U37832 (N_37832,N_37643,N_37722);
and U37833 (N_37833,N_37580,N_37510);
nor U37834 (N_37834,N_37609,N_37668);
or U37835 (N_37835,N_37525,N_37624);
and U37836 (N_37836,N_37688,N_37734);
or U37837 (N_37837,N_37577,N_37707);
or U37838 (N_37838,N_37520,N_37659);
nand U37839 (N_37839,N_37713,N_37529);
nor U37840 (N_37840,N_37627,N_37586);
nand U37841 (N_37841,N_37557,N_37678);
xnor U37842 (N_37842,N_37553,N_37660);
and U37843 (N_37843,N_37614,N_37559);
or U37844 (N_37844,N_37615,N_37690);
nor U37845 (N_37845,N_37693,N_37732);
nand U37846 (N_37846,N_37616,N_37578);
and U37847 (N_37847,N_37714,N_37516);
nand U37848 (N_37848,N_37625,N_37595);
or U37849 (N_37849,N_37631,N_37512);
nor U37850 (N_37850,N_37555,N_37536);
nor U37851 (N_37851,N_37672,N_37685);
nand U37852 (N_37852,N_37594,N_37608);
or U37853 (N_37853,N_37548,N_37676);
or U37854 (N_37854,N_37620,N_37505);
nor U37855 (N_37855,N_37720,N_37671);
nand U37856 (N_37856,N_37726,N_37710);
or U37857 (N_37857,N_37551,N_37738);
nand U37858 (N_37858,N_37538,N_37570);
xnor U37859 (N_37859,N_37746,N_37566);
and U37860 (N_37860,N_37664,N_37725);
or U37861 (N_37861,N_37558,N_37716);
nor U37862 (N_37862,N_37622,N_37549);
or U37863 (N_37863,N_37701,N_37626);
and U37864 (N_37864,N_37568,N_37730);
xnor U37865 (N_37865,N_37654,N_37687);
xnor U37866 (N_37866,N_37729,N_37579);
or U37867 (N_37867,N_37717,N_37564);
nor U37868 (N_37868,N_37545,N_37721);
or U37869 (N_37869,N_37509,N_37715);
nor U37870 (N_37870,N_37705,N_37598);
or U37871 (N_37871,N_37611,N_37528);
nor U37872 (N_37872,N_37540,N_37547);
nand U37873 (N_37873,N_37635,N_37521);
nor U37874 (N_37874,N_37574,N_37603);
xor U37875 (N_37875,N_37743,N_37629);
and U37876 (N_37876,N_37586,N_37651);
nor U37877 (N_37877,N_37575,N_37519);
and U37878 (N_37878,N_37718,N_37609);
and U37879 (N_37879,N_37506,N_37533);
xnor U37880 (N_37880,N_37747,N_37648);
or U37881 (N_37881,N_37592,N_37633);
nand U37882 (N_37882,N_37566,N_37700);
or U37883 (N_37883,N_37689,N_37540);
xnor U37884 (N_37884,N_37529,N_37575);
and U37885 (N_37885,N_37581,N_37535);
and U37886 (N_37886,N_37566,N_37552);
nand U37887 (N_37887,N_37549,N_37532);
nor U37888 (N_37888,N_37522,N_37647);
nand U37889 (N_37889,N_37687,N_37725);
and U37890 (N_37890,N_37582,N_37536);
nor U37891 (N_37891,N_37609,N_37623);
and U37892 (N_37892,N_37694,N_37627);
xor U37893 (N_37893,N_37616,N_37727);
and U37894 (N_37894,N_37596,N_37539);
and U37895 (N_37895,N_37729,N_37688);
and U37896 (N_37896,N_37605,N_37509);
nand U37897 (N_37897,N_37672,N_37678);
nor U37898 (N_37898,N_37618,N_37718);
and U37899 (N_37899,N_37702,N_37561);
nor U37900 (N_37900,N_37608,N_37655);
or U37901 (N_37901,N_37536,N_37696);
nand U37902 (N_37902,N_37552,N_37694);
nand U37903 (N_37903,N_37583,N_37513);
xnor U37904 (N_37904,N_37742,N_37586);
or U37905 (N_37905,N_37679,N_37666);
nor U37906 (N_37906,N_37556,N_37583);
nand U37907 (N_37907,N_37536,N_37716);
nor U37908 (N_37908,N_37739,N_37682);
or U37909 (N_37909,N_37503,N_37518);
nand U37910 (N_37910,N_37671,N_37512);
xnor U37911 (N_37911,N_37720,N_37666);
xor U37912 (N_37912,N_37683,N_37694);
xor U37913 (N_37913,N_37557,N_37576);
nand U37914 (N_37914,N_37671,N_37674);
nand U37915 (N_37915,N_37515,N_37563);
or U37916 (N_37916,N_37737,N_37526);
nand U37917 (N_37917,N_37677,N_37502);
nand U37918 (N_37918,N_37682,N_37512);
nor U37919 (N_37919,N_37568,N_37549);
nand U37920 (N_37920,N_37652,N_37608);
nor U37921 (N_37921,N_37637,N_37551);
or U37922 (N_37922,N_37589,N_37678);
nand U37923 (N_37923,N_37569,N_37593);
and U37924 (N_37924,N_37681,N_37511);
xnor U37925 (N_37925,N_37672,N_37525);
or U37926 (N_37926,N_37741,N_37714);
or U37927 (N_37927,N_37522,N_37527);
xor U37928 (N_37928,N_37711,N_37666);
nand U37929 (N_37929,N_37722,N_37500);
nand U37930 (N_37930,N_37684,N_37583);
and U37931 (N_37931,N_37578,N_37744);
and U37932 (N_37932,N_37508,N_37626);
nand U37933 (N_37933,N_37504,N_37695);
and U37934 (N_37934,N_37564,N_37634);
xnor U37935 (N_37935,N_37746,N_37622);
nor U37936 (N_37936,N_37605,N_37674);
nand U37937 (N_37937,N_37643,N_37623);
or U37938 (N_37938,N_37599,N_37528);
or U37939 (N_37939,N_37640,N_37704);
or U37940 (N_37940,N_37686,N_37560);
nand U37941 (N_37941,N_37719,N_37691);
xnor U37942 (N_37942,N_37665,N_37701);
nor U37943 (N_37943,N_37723,N_37612);
or U37944 (N_37944,N_37661,N_37550);
or U37945 (N_37945,N_37736,N_37550);
nor U37946 (N_37946,N_37551,N_37627);
xnor U37947 (N_37947,N_37581,N_37714);
xor U37948 (N_37948,N_37729,N_37744);
and U37949 (N_37949,N_37586,N_37663);
xnor U37950 (N_37950,N_37597,N_37555);
nor U37951 (N_37951,N_37577,N_37556);
and U37952 (N_37952,N_37666,N_37680);
nor U37953 (N_37953,N_37687,N_37733);
and U37954 (N_37954,N_37727,N_37587);
nand U37955 (N_37955,N_37675,N_37736);
xor U37956 (N_37956,N_37627,N_37695);
nor U37957 (N_37957,N_37619,N_37639);
and U37958 (N_37958,N_37545,N_37561);
and U37959 (N_37959,N_37744,N_37649);
xor U37960 (N_37960,N_37503,N_37673);
and U37961 (N_37961,N_37571,N_37723);
nor U37962 (N_37962,N_37605,N_37538);
nand U37963 (N_37963,N_37679,N_37649);
nor U37964 (N_37964,N_37688,N_37672);
xor U37965 (N_37965,N_37532,N_37602);
or U37966 (N_37966,N_37523,N_37607);
nand U37967 (N_37967,N_37579,N_37601);
and U37968 (N_37968,N_37675,N_37681);
and U37969 (N_37969,N_37615,N_37565);
nand U37970 (N_37970,N_37532,N_37714);
nand U37971 (N_37971,N_37589,N_37567);
nor U37972 (N_37972,N_37682,N_37712);
and U37973 (N_37973,N_37559,N_37732);
nand U37974 (N_37974,N_37712,N_37662);
nor U37975 (N_37975,N_37633,N_37561);
nand U37976 (N_37976,N_37678,N_37677);
nand U37977 (N_37977,N_37540,N_37602);
nand U37978 (N_37978,N_37674,N_37670);
nor U37979 (N_37979,N_37592,N_37749);
xor U37980 (N_37980,N_37719,N_37742);
nand U37981 (N_37981,N_37537,N_37704);
or U37982 (N_37982,N_37662,N_37594);
nor U37983 (N_37983,N_37551,N_37715);
nand U37984 (N_37984,N_37615,N_37739);
and U37985 (N_37985,N_37605,N_37534);
or U37986 (N_37986,N_37517,N_37660);
nor U37987 (N_37987,N_37747,N_37658);
or U37988 (N_37988,N_37650,N_37654);
xnor U37989 (N_37989,N_37614,N_37686);
nand U37990 (N_37990,N_37641,N_37712);
nand U37991 (N_37991,N_37505,N_37700);
nand U37992 (N_37992,N_37603,N_37506);
or U37993 (N_37993,N_37524,N_37646);
and U37994 (N_37994,N_37719,N_37576);
and U37995 (N_37995,N_37657,N_37727);
nor U37996 (N_37996,N_37644,N_37665);
xor U37997 (N_37997,N_37632,N_37630);
xor U37998 (N_37998,N_37554,N_37650);
and U37999 (N_37999,N_37610,N_37678);
xnor U38000 (N_38000,N_37954,N_37902);
nand U38001 (N_38001,N_37776,N_37769);
nand U38002 (N_38002,N_37854,N_37812);
xnor U38003 (N_38003,N_37939,N_37916);
xor U38004 (N_38004,N_37774,N_37777);
nand U38005 (N_38005,N_37980,N_37845);
or U38006 (N_38006,N_37846,N_37792);
nand U38007 (N_38007,N_37835,N_37829);
and U38008 (N_38008,N_37999,N_37831);
nor U38009 (N_38009,N_37915,N_37797);
and U38010 (N_38010,N_37768,N_37978);
nand U38011 (N_38011,N_37799,N_37907);
nand U38012 (N_38012,N_37942,N_37901);
nor U38013 (N_38013,N_37826,N_37844);
nand U38014 (N_38014,N_37906,N_37969);
nand U38015 (N_38015,N_37856,N_37802);
or U38016 (N_38016,N_37933,N_37991);
or U38017 (N_38017,N_37806,N_37823);
xnor U38018 (N_38018,N_37897,N_37838);
nand U38019 (N_38019,N_37995,N_37919);
nor U38020 (N_38020,N_37819,N_37920);
nor U38021 (N_38021,N_37773,N_37898);
and U38022 (N_38022,N_37782,N_37968);
and U38023 (N_38023,N_37926,N_37816);
xnor U38024 (N_38024,N_37945,N_37890);
nor U38025 (N_38025,N_37783,N_37869);
nand U38026 (N_38026,N_37830,N_37953);
nor U38027 (N_38027,N_37785,N_37859);
xor U38028 (N_38028,N_37765,N_37763);
and U38029 (N_38029,N_37781,N_37853);
xnor U38030 (N_38030,N_37934,N_37943);
and U38031 (N_38031,N_37866,N_37895);
nor U38032 (N_38032,N_37810,N_37848);
nor U38033 (N_38033,N_37972,N_37904);
and U38034 (N_38034,N_37755,N_37805);
xnor U38035 (N_38035,N_37923,N_37917);
and U38036 (N_38036,N_37849,N_37825);
nand U38037 (N_38037,N_37770,N_37903);
nand U38038 (N_38038,N_37871,N_37753);
xnor U38039 (N_38039,N_37852,N_37918);
and U38040 (N_38040,N_37973,N_37964);
or U38041 (N_38041,N_37882,N_37985);
nor U38042 (N_38042,N_37790,N_37905);
nor U38043 (N_38043,N_37780,N_37861);
nand U38044 (N_38044,N_37837,N_37757);
or U38045 (N_38045,N_37894,N_37807);
nand U38046 (N_38046,N_37824,N_37883);
nand U38047 (N_38047,N_37789,N_37970);
and U38048 (N_38048,N_37908,N_37868);
xnor U38049 (N_38049,N_37767,N_37922);
nor U38050 (N_38050,N_37752,N_37850);
xnor U38051 (N_38051,N_37959,N_37966);
nand U38052 (N_38052,N_37779,N_37937);
nand U38053 (N_38053,N_37857,N_37936);
nand U38054 (N_38054,N_37888,N_37865);
xor U38055 (N_38055,N_37935,N_37815);
nor U38056 (N_38056,N_37965,N_37821);
or U38057 (N_38057,N_37863,N_37875);
and U38058 (N_38058,N_37950,N_37988);
nand U38059 (N_38059,N_37836,N_37791);
and U38060 (N_38060,N_37941,N_37803);
or U38061 (N_38061,N_37833,N_37958);
or U38062 (N_38062,N_37762,N_37794);
and U38063 (N_38063,N_37771,N_37884);
nor U38064 (N_38064,N_37944,N_37967);
xnor U38065 (N_38065,N_37960,N_37987);
and U38066 (N_38066,N_37977,N_37788);
or U38067 (N_38067,N_37998,N_37855);
and U38068 (N_38068,N_37962,N_37778);
nand U38069 (N_38069,N_37860,N_37842);
xor U38070 (N_38070,N_37843,N_37913);
and U38071 (N_38071,N_37760,N_37910);
nand U38072 (N_38072,N_37952,N_37879);
xnor U38073 (N_38073,N_37867,N_37928);
xnor U38074 (N_38074,N_37840,N_37834);
nor U38075 (N_38075,N_37956,N_37759);
xor U38076 (N_38076,N_37921,N_37955);
nor U38077 (N_38077,N_37775,N_37881);
xnor U38078 (N_38078,N_37847,N_37761);
or U38079 (N_38079,N_37951,N_37974);
nor U38080 (N_38080,N_37864,N_37784);
or U38081 (N_38081,N_37912,N_37754);
xnor U38082 (N_38082,N_37798,N_37931);
or U38083 (N_38083,N_37874,N_37756);
xnor U38084 (N_38084,N_37811,N_37986);
and U38085 (N_38085,N_37993,N_37996);
nand U38086 (N_38086,N_37885,N_37975);
or U38087 (N_38087,N_37766,N_37909);
nand U38088 (N_38088,N_37899,N_37801);
xnor U38089 (N_38089,N_37929,N_37880);
and U38090 (N_38090,N_37795,N_37981);
nand U38091 (N_38091,N_37813,N_37971);
nand U38092 (N_38092,N_37946,N_37827);
nand U38093 (N_38093,N_37961,N_37911);
nor U38094 (N_38094,N_37873,N_37924);
xor U38095 (N_38095,N_37820,N_37994);
xor U38096 (N_38096,N_37793,N_37896);
and U38097 (N_38097,N_37893,N_37822);
and U38098 (N_38098,N_37886,N_37957);
nor U38099 (N_38099,N_37858,N_37989);
xnor U38100 (N_38100,N_37751,N_37979);
nor U38101 (N_38101,N_37984,N_37990);
nand U38102 (N_38102,N_37930,N_37818);
and U38103 (N_38103,N_37949,N_37870);
nor U38104 (N_38104,N_37832,N_37814);
or U38105 (N_38105,N_37877,N_37796);
and U38106 (N_38106,N_37925,N_37983);
or U38107 (N_38107,N_37892,N_37914);
nand U38108 (N_38108,N_37800,N_37938);
xor U38109 (N_38109,N_37887,N_37891);
nand U38110 (N_38110,N_37927,N_37872);
or U38111 (N_38111,N_37841,N_37876);
and U38112 (N_38112,N_37804,N_37947);
or U38113 (N_38113,N_37889,N_37787);
nand U38114 (N_38114,N_37878,N_37764);
nor U38115 (N_38115,N_37839,N_37948);
nor U38116 (N_38116,N_37828,N_37940);
xnor U38117 (N_38117,N_37900,N_37750);
nor U38118 (N_38118,N_37932,N_37997);
nor U38119 (N_38119,N_37976,N_37963);
or U38120 (N_38120,N_37851,N_37862);
or U38121 (N_38121,N_37786,N_37772);
nor U38122 (N_38122,N_37808,N_37758);
nor U38123 (N_38123,N_37982,N_37809);
nor U38124 (N_38124,N_37817,N_37992);
or U38125 (N_38125,N_37889,N_37786);
and U38126 (N_38126,N_37995,N_37820);
or U38127 (N_38127,N_37860,N_37984);
xor U38128 (N_38128,N_37811,N_37795);
nand U38129 (N_38129,N_37988,N_37827);
nor U38130 (N_38130,N_37885,N_37814);
and U38131 (N_38131,N_37960,N_37953);
xnor U38132 (N_38132,N_37927,N_37836);
or U38133 (N_38133,N_37790,N_37751);
or U38134 (N_38134,N_37868,N_37914);
or U38135 (N_38135,N_37950,N_37784);
xnor U38136 (N_38136,N_37924,N_37767);
xnor U38137 (N_38137,N_37786,N_37925);
nand U38138 (N_38138,N_37775,N_37909);
xnor U38139 (N_38139,N_37750,N_37969);
xnor U38140 (N_38140,N_37967,N_37750);
and U38141 (N_38141,N_37887,N_37833);
xor U38142 (N_38142,N_37907,N_37897);
nand U38143 (N_38143,N_37962,N_37940);
xnor U38144 (N_38144,N_37982,N_37763);
and U38145 (N_38145,N_37892,N_37970);
or U38146 (N_38146,N_37951,N_37887);
nor U38147 (N_38147,N_37753,N_37785);
and U38148 (N_38148,N_37780,N_37978);
xnor U38149 (N_38149,N_37949,N_37923);
and U38150 (N_38150,N_37924,N_37880);
nor U38151 (N_38151,N_37811,N_37755);
nor U38152 (N_38152,N_37952,N_37967);
or U38153 (N_38153,N_37833,N_37871);
and U38154 (N_38154,N_37916,N_37849);
nand U38155 (N_38155,N_37990,N_37853);
or U38156 (N_38156,N_37880,N_37907);
nand U38157 (N_38157,N_37833,N_37846);
nand U38158 (N_38158,N_37960,N_37890);
or U38159 (N_38159,N_37820,N_37952);
nand U38160 (N_38160,N_37903,N_37801);
and U38161 (N_38161,N_37966,N_37886);
or U38162 (N_38162,N_37991,N_37989);
and U38163 (N_38163,N_37989,N_37850);
nand U38164 (N_38164,N_37818,N_37931);
xnor U38165 (N_38165,N_37974,N_37865);
and U38166 (N_38166,N_37808,N_37810);
nand U38167 (N_38167,N_37847,N_37921);
nand U38168 (N_38168,N_37937,N_37870);
xor U38169 (N_38169,N_37870,N_37938);
and U38170 (N_38170,N_37923,N_37782);
xnor U38171 (N_38171,N_37809,N_37834);
or U38172 (N_38172,N_37892,N_37907);
nor U38173 (N_38173,N_37962,N_37843);
nor U38174 (N_38174,N_37758,N_37806);
nor U38175 (N_38175,N_37891,N_37814);
or U38176 (N_38176,N_37902,N_37930);
nand U38177 (N_38177,N_37892,N_37810);
or U38178 (N_38178,N_37897,N_37820);
xor U38179 (N_38179,N_37917,N_37804);
nand U38180 (N_38180,N_37986,N_37800);
and U38181 (N_38181,N_37765,N_37761);
and U38182 (N_38182,N_37826,N_37986);
xor U38183 (N_38183,N_37935,N_37873);
or U38184 (N_38184,N_37944,N_37804);
xor U38185 (N_38185,N_37769,N_37984);
or U38186 (N_38186,N_37857,N_37872);
nand U38187 (N_38187,N_37976,N_37771);
and U38188 (N_38188,N_37993,N_37947);
nand U38189 (N_38189,N_37868,N_37803);
nor U38190 (N_38190,N_37820,N_37946);
and U38191 (N_38191,N_37999,N_37963);
nand U38192 (N_38192,N_37852,N_37878);
and U38193 (N_38193,N_37850,N_37810);
and U38194 (N_38194,N_37867,N_37920);
and U38195 (N_38195,N_37861,N_37869);
and U38196 (N_38196,N_37951,N_37895);
and U38197 (N_38197,N_37939,N_37963);
or U38198 (N_38198,N_37786,N_37918);
nand U38199 (N_38199,N_37823,N_37795);
nor U38200 (N_38200,N_37894,N_37937);
xor U38201 (N_38201,N_37775,N_37832);
nand U38202 (N_38202,N_37788,N_37958);
nand U38203 (N_38203,N_37976,N_37893);
nand U38204 (N_38204,N_37798,N_37943);
nor U38205 (N_38205,N_37812,N_37763);
nor U38206 (N_38206,N_37872,N_37856);
nor U38207 (N_38207,N_37842,N_37762);
nand U38208 (N_38208,N_37779,N_37856);
nand U38209 (N_38209,N_37854,N_37952);
xnor U38210 (N_38210,N_37944,N_37895);
or U38211 (N_38211,N_37971,N_37889);
nor U38212 (N_38212,N_37966,N_37822);
and U38213 (N_38213,N_37988,N_37772);
nor U38214 (N_38214,N_37943,N_37963);
or U38215 (N_38215,N_37858,N_37944);
or U38216 (N_38216,N_37870,N_37894);
nor U38217 (N_38217,N_37979,N_37975);
nand U38218 (N_38218,N_37783,N_37997);
nand U38219 (N_38219,N_37910,N_37884);
and U38220 (N_38220,N_37855,N_37895);
xnor U38221 (N_38221,N_37986,N_37861);
xor U38222 (N_38222,N_37983,N_37883);
or U38223 (N_38223,N_37785,N_37758);
or U38224 (N_38224,N_37864,N_37826);
xnor U38225 (N_38225,N_37762,N_37989);
and U38226 (N_38226,N_37797,N_37853);
or U38227 (N_38227,N_37896,N_37772);
xnor U38228 (N_38228,N_37850,N_37795);
nor U38229 (N_38229,N_37816,N_37879);
nand U38230 (N_38230,N_37993,N_37750);
xnor U38231 (N_38231,N_37937,N_37883);
nor U38232 (N_38232,N_37760,N_37994);
or U38233 (N_38233,N_37914,N_37927);
xor U38234 (N_38234,N_37858,N_37927);
xor U38235 (N_38235,N_37860,N_37949);
or U38236 (N_38236,N_37858,N_37919);
and U38237 (N_38237,N_37969,N_37820);
nand U38238 (N_38238,N_37855,N_37976);
nand U38239 (N_38239,N_37815,N_37785);
xnor U38240 (N_38240,N_37977,N_37757);
and U38241 (N_38241,N_37922,N_37938);
nand U38242 (N_38242,N_37797,N_37906);
xnor U38243 (N_38243,N_37800,N_37787);
nor U38244 (N_38244,N_37792,N_37799);
or U38245 (N_38245,N_37849,N_37750);
xnor U38246 (N_38246,N_37887,N_37884);
or U38247 (N_38247,N_37773,N_37818);
xnor U38248 (N_38248,N_37948,N_37871);
xnor U38249 (N_38249,N_37832,N_37882);
xor U38250 (N_38250,N_38226,N_38075);
and U38251 (N_38251,N_38041,N_38191);
nor U38252 (N_38252,N_38229,N_38003);
xor U38253 (N_38253,N_38043,N_38158);
nand U38254 (N_38254,N_38239,N_38004);
and U38255 (N_38255,N_38100,N_38073);
nor U38256 (N_38256,N_38001,N_38152);
xor U38257 (N_38257,N_38164,N_38110);
and U38258 (N_38258,N_38130,N_38161);
xnor U38259 (N_38259,N_38085,N_38209);
nor U38260 (N_38260,N_38079,N_38205);
xnor U38261 (N_38261,N_38201,N_38248);
or U38262 (N_38262,N_38056,N_38242);
xnor U38263 (N_38263,N_38218,N_38121);
or U38264 (N_38264,N_38195,N_38063);
nand U38265 (N_38265,N_38145,N_38114);
and U38266 (N_38266,N_38120,N_38159);
xnor U38267 (N_38267,N_38113,N_38142);
and U38268 (N_38268,N_38123,N_38156);
nand U38269 (N_38269,N_38125,N_38091);
and U38270 (N_38270,N_38240,N_38017);
nand U38271 (N_38271,N_38206,N_38211);
or U38272 (N_38272,N_38122,N_38208);
or U38273 (N_38273,N_38066,N_38144);
nand U38274 (N_38274,N_38234,N_38000);
nand U38275 (N_38275,N_38002,N_38105);
or U38276 (N_38276,N_38135,N_38098);
xor U38277 (N_38277,N_38057,N_38138);
and U38278 (N_38278,N_38081,N_38177);
xnor U38279 (N_38279,N_38112,N_38102);
nand U38280 (N_38280,N_38035,N_38050);
nand U38281 (N_38281,N_38092,N_38162);
nor U38282 (N_38282,N_38046,N_38154);
xor U38283 (N_38283,N_38048,N_38187);
xor U38284 (N_38284,N_38180,N_38243);
and U38285 (N_38285,N_38019,N_38228);
and U38286 (N_38286,N_38055,N_38015);
and U38287 (N_38287,N_38225,N_38064);
nor U38288 (N_38288,N_38101,N_38054);
nand U38289 (N_38289,N_38053,N_38246);
xnor U38290 (N_38290,N_38222,N_38196);
xor U38291 (N_38291,N_38087,N_38132);
nor U38292 (N_38292,N_38089,N_38137);
or U38293 (N_38293,N_38096,N_38020);
xnor U38294 (N_38294,N_38155,N_38038);
or U38295 (N_38295,N_38065,N_38029);
and U38296 (N_38296,N_38127,N_38249);
xor U38297 (N_38297,N_38178,N_38190);
nand U38298 (N_38298,N_38223,N_38028);
or U38299 (N_38299,N_38067,N_38082);
and U38300 (N_38300,N_38151,N_38212);
and U38301 (N_38301,N_38045,N_38059);
nor U38302 (N_38302,N_38213,N_38099);
and U38303 (N_38303,N_38016,N_38174);
or U38304 (N_38304,N_38047,N_38024);
or U38305 (N_38305,N_38094,N_38188);
xnor U38306 (N_38306,N_38183,N_38039);
xnor U38307 (N_38307,N_38236,N_38088);
nand U38308 (N_38308,N_38058,N_38148);
or U38309 (N_38309,N_38012,N_38136);
nand U38310 (N_38310,N_38171,N_38026);
and U38311 (N_38311,N_38128,N_38042);
and U38312 (N_38312,N_38005,N_38068);
or U38313 (N_38313,N_38097,N_38077);
xnor U38314 (N_38314,N_38049,N_38106);
nor U38315 (N_38315,N_38146,N_38032);
xnor U38316 (N_38316,N_38008,N_38072);
and U38317 (N_38317,N_38023,N_38103);
nand U38318 (N_38318,N_38198,N_38084);
nor U38319 (N_38319,N_38233,N_38062);
xnor U38320 (N_38320,N_38227,N_38104);
or U38321 (N_38321,N_38182,N_38160);
or U38322 (N_38322,N_38051,N_38149);
nor U38323 (N_38323,N_38207,N_38245);
and U38324 (N_38324,N_38216,N_38095);
nor U38325 (N_38325,N_38247,N_38139);
xor U38326 (N_38326,N_38157,N_38090);
and U38327 (N_38327,N_38111,N_38013);
nor U38328 (N_38328,N_38117,N_38166);
xor U38329 (N_38329,N_38086,N_38129);
or U38330 (N_38330,N_38124,N_38034);
nor U38331 (N_38331,N_38014,N_38169);
or U38332 (N_38332,N_38022,N_38184);
or U38333 (N_38333,N_38217,N_38214);
or U38334 (N_38334,N_38170,N_38031);
or U38335 (N_38335,N_38133,N_38021);
or U38336 (N_38336,N_38036,N_38194);
xnor U38337 (N_38337,N_38027,N_38060);
nor U38338 (N_38338,N_38224,N_38052);
nor U38339 (N_38339,N_38009,N_38199);
or U38340 (N_38340,N_38176,N_38197);
nor U38341 (N_38341,N_38109,N_38074);
and U38342 (N_38342,N_38107,N_38167);
xnor U38343 (N_38343,N_38069,N_38230);
nor U38344 (N_38344,N_38175,N_38141);
nor U38345 (N_38345,N_38078,N_38018);
or U38346 (N_38346,N_38203,N_38219);
and U38347 (N_38347,N_38126,N_38220);
nand U38348 (N_38348,N_38116,N_38037);
nor U38349 (N_38349,N_38192,N_38185);
nor U38350 (N_38350,N_38231,N_38010);
xor U38351 (N_38351,N_38025,N_38215);
nand U38352 (N_38352,N_38118,N_38030);
or U38353 (N_38353,N_38011,N_38061);
xnor U38354 (N_38354,N_38083,N_38076);
nand U38355 (N_38355,N_38033,N_38210);
or U38356 (N_38356,N_38235,N_38200);
or U38357 (N_38357,N_38189,N_38044);
nand U38358 (N_38358,N_38119,N_38221);
nand U38359 (N_38359,N_38232,N_38172);
xor U38360 (N_38360,N_38093,N_38165);
and U38361 (N_38361,N_38071,N_38202);
xor U38362 (N_38362,N_38108,N_38241);
and U38363 (N_38363,N_38147,N_38237);
and U38364 (N_38364,N_38238,N_38140);
xor U38365 (N_38365,N_38153,N_38040);
xor U38366 (N_38366,N_38179,N_38163);
nor U38367 (N_38367,N_38244,N_38115);
nor U38368 (N_38368,N_38193,N_38168);
and U38369 (N_38369,N_38134,N_38007);
xnor U38370 (N_38370,N_38204,N_38006);
xnor U38371 (N_38371,N_38150,N_38070);
xor U38372 (N_38372,N_38186,N_38173);
xor U38373 (N_38373,N_38181,N_38080);
and U38374 (N_38374,N_38131,N_38143);
or U38375 (N_38375,N_38160,N_38025);
or U38376 (N_38376,N_38205,N_38234);
or U38377 (N_38377,N_38099,N_38107);
or U38378 (N_38378,N_38020,N_38097);
and U38379 (N_38379,N_38116,N_38015);
nand U38380 (N_38380,N_38092,N_38035);
nand U38381 (N_38381,N_38154,N_38030);
xor U38382 (N_38382,N_38230,N_38228);
xnor U38383 (N_38383,N_38097,N_38157);
or U38384 (N_38384,N_38064,N_38234);
or U38385 (N_38385,N_38102,N_38021);
nor U38386 (N_38386,N_38163,N_38047);
nand U38387 (N_38387,N_38172,N_38123);
nand U38388 (N_38388,N_38174,N_38071);
nand U38389 (N_38389,N_38069,N_38150);
nand U38390 (N_38390,N_38044,N_38040);
or U38391 (N_38391,N_38204,N_38166);
nand U38392 (N_38392,N_38051,N_38044);
nor U38393 (N_38393,N_38206,N_38012);
or U38394 (N_38394,N_38244,N_38101);
nor U38395 (N_38395,N_38160,N_38241);
nand U38396 (N_38396,N_38118,N_38166);
or U38397 (N_38397,N_38050,N_38195);
nand U38398 (N_38398,N_38106,N_38018);
and U38399 (N_38399,N_38087,N_38060);
nor U38400 (N_38400,N_38212,N_38215);
nand U38401 (N_38401,N_38017,N_38132);
nand U38402 (N_38402,N_38083,N_38175);
and U38403 (N_38403,N_38000,N_38178);
nor U38404 (N_38404,N_38038,N_38078);
nand U38405 (N_38405,N_38117,N_38042);
xor U38406 (N_38406,N_38135,N_38101);
nor U38407 (N_38407,N_38208,N_38140);
or U38408 (N_38408,N_38101,N_38092);
nand U38409 (N_38409,N_38052,N_38136);
or U38410 (N_38410,N_38007,N_38158);
nand U38411 (N_38411,N_38096,N_38203);
or U38412 (N_38412,N_38176,N_38211);
or U38413 (N_38413,N_38105,N_38011);
or U38414 (N_38414,N_38191,N_38222);
and U38415 (N_38415,N_38036,N_38002);
nor U38416 (N_38416,N_38001,N_38205);
or U38417 (N_38417,N_38176,N_38078);
and U38418 (N_38418,N_38195,N_38145);
or U38419 (N_38419,N_38016,N_38168);
xor U38420 (N_38420,N_38145,N_38149);
xor U38421 (N_38421,N_38061,N_38184);
nand U38422 (N_38422,N_38108,N_38161);
nor U38423 (N_38423,N_38036,N_38037);
nand U38424 (N_38424,N_38249,N_38167);
and U38425 (N_38425,N_38088,N_38172);
nor U38426 (N_38426,N_38142,N_38231);
and U38427 (N_38427,N_38032,N_38019);
nor U38428 (N_38428,N_38234,N_38004);
and U38429 (N_38429,N_38222,N_38162);
or U38430 (N_38430,N_38243,N_38083);
and U38431 (N_38431,N_38168,N_38233);
nand U38432 (N_38432,N_38013,N_38043);
nor U38433 (N_38433,N_38105,N_38214);
nor U38434 (N_38434,N_38030,N_38248);
nor U38435 (N_38435,N_38067,N_38211);
nor U38436 (N_38436,N_38174,N_38209);
xnor U38437 (N_38437,N_38034,N_38149);
or U38438 (N_38438,N_38003,N_38096);
nand U38439 (N_38439,N_38039,N_38016);
and U38440 (N_38440,N_38174,N_38223);
nand U38441 (N_38441,N_38071,N_38170);
nor U38442 (N_38442,N_38057,N_38180);
or U38443 (N_38443,N_38245,N_38013);
and U38444 (N_38444,N_38136,N_38177);
nor U38445 (N_38445,N_38030,N_38165);
and U38446 (N_38446,N_38040,N_38001);
nor U38447 (N_38447,N_38057,N_38208);
or U38448 (N_38448,N_38132,N_38211);
xnor U38449 (N_38449,N_38178,N_38148);
xor U38450 (N_38450,N_38230,N_38152);
nor U38451 (N_38451,N_38125,N_38187);
and U38452 (N_38452,N_38151,N_38236);
and U38453 (N_38453,N_38214,N_38014);
and U38454 (N_38454,N_38142,N_38139);
or U38455 (N_38455,N_38050,N_38108);
xnor U38456 (N_38456,N_38061,N_38113);
nor U38457 (N_38457,N_38157,N_38091);
nand U38458 (N_38458,N_38041,N_38217);
xor U38459 (N_38459,N_38025,N_38106);
or U38460 (N_38460,N_38147,N_38121);
and U38461 (N_38461,N_38197,N_38152);
or U38462 (N_38462,N_38123,N_38134);
xor U38463 (N_38463,N_38137,N_38040);
and U38464 (N_38464,N_38019,N_38079);
or U38465 (N_38465,N_38051,N_38009);
or U38466 (N_38466,N_38089,N_38134);
nor U38467 (N_38467,N_38079,N_38229);
or U38468 (N_38468,N_38022,N_38151);
xor U38469 (N_38469,N_38170,N_38183);
and U38470 (N_38470,N_38090,N_38143);
nor U38471 (N_38471,N_38135,N_38146);
and U38472 (N_38472,N_38109,N_38003);
or U38473 (N_38473,N_38153,N_38239);
and U38474 (N_38474,N_38004,N_38068);
xor U38475 (N_38475,N_38216,N_38014);
and U38476 (N_38476,N_38158,N_38233);
nand U38477 (N_38477,N_38211,N_38113);
nand U38478 (N_38478,N_38052,N_38024);
nor U38479 (N_38479,N_38073,N_38006);
and U38480 (N_38480,N_38065,N_38082);
nand U38481 (N_38481,N_38208,N_38111);
or U38482 (N_38482,N_38078,N_38232);
and U38483 (N_38483,N_38196,N_38234);
nand U38484 (N_38484,N_38052,N_38006);
nor U38485 (N_38485,N_38241,N_38094);
and U38486 (N_38486,N_38044,N_38036);
and U38487 (N_38487,N_38041,N_38158);
nand U38488 (N_38488,N_38207,N_38202);
xor U38489 (N_38489,N_38025,N_38126);
xnor U38490 (N_38490,N_38100,N_38108);
nor U38491 (N_38491,N_38162,N_38063);
xnor U38492 (N_38492,N_38219,N_38045);
or U38493 (N_38493,N_38241,N_38206);
nor U38494 (N_38494,N_38008,N_38144);
nor U38495 (N_38495,N_38153,N_38230);
nor U38496 (N_38496,N_38120,N_38075);
and U38497 (N_38497,N_38135,N_38132);
nor U38498 (N_38498,N_38069,N_38032);
nor U38499 (N_38499,N_38066,N_38176);
nand U38500 (N_38500,N_38416,N_38402);
or U38501 (N_38501,N_38485,N_38400);
or U38502 (N_38502,N_38381,N_38286);
nor U38503 (N_38503,N_38496,N_38395);
nor U38504 (N_38504,N_38494,N_38462);
nand U38505 (N_38505,N_38391,N_38482);
xor U38506 (N_38506,N_38479,N_38401);
or U38507 (N_38507,N_38302,N_38307);
xnor U38508 (N_38508,N_38281,N_38461);
nand U38509 (N_38509,N_38480,N_38315);
nor U38510 (N_38510,N_38426,N_38303);
xor U38511 (N_38511,N_38396,N_38475);
and U38512 (N_38512,N_38367,N_38291);
xor U38513 (N_38513,N_38347,N_38487);
xnor U38514 (N_38514,N_38254,N_38257);
or U38515 (N_38515,N_38456,N_38273);
xor U38516 (N_38516,N_38417,N_38352);
nand U38517 (N_38517,N_38350,N_38411);
xor U38518 (N_38518,N_38343,N_38305);
and U38519 (N_38519,N_38375,N_38448);
or U38520 (N_38520,N_38441,N_38285);
and U38521 (N_38521,N_38477,N_38328);
nor U38522 (N_38522,N_38326,N_38360);
xor U38523 (N_38523,N_38435,N_38331);
or U38524 (N_38524,N_38329,N_38333);
nand U38525 (N_38525,N_38301,N_38459);
nand U38526 (N_38526,N_38432,N_38358);
xnor U38527 (N_38527,N_38310,N_38324);
or U38528 (N_38528,N_38420,N_38457);
and U38529 (N_38529,N_38450,N_38412);
xnor U38530 (N_38530,N_38268,N_38334);
nand U38531 (N_38531,N_38425,N_38455);
xnor U38532 (N_38532,N_38260,N_38481);
xnor U38533 (N_38533,N_38357,N_38321);
nor U38534 (N_38534,N_38282,N_38405);
xor U38535 (N_38535,N_38436,N_38262);
and U38536 (N_38536,N_38369,N_38362);
xor U38537 (N_38537,N_38403,N_38445);
nor U38538 (N_38538,N_38446,N_38337);
xor U38539 (N_38539,N_38255,N_38449);
nand U38540 (N_38540,N_38332,N_38299);
and U38541 (N_38541,N_38492,N_38320);
and U38542 (N_38542,N_38382,N_38486);
xor U38543 (N_38543,N_38390,N_38271);
and U38544 (N_38544,N_38258,N_38460);
nor U38545 (N_38545,N_38311,N_38344);
nor U38546 (N_38546,N_38309,N_38251);
or U38547 (N_38547,N_38438,N_38387);
and U38548 (N_38548,N_38313,N_38341);
nand U38549 (N_38549,N_38434,N_38284);
nand U38550 (N_38550,N_38379,N_38270);
xnor U38551 (N_38551,N_38444,N_38389);
nor U38552 (N_38552,N_38470,N_38272);
or U38553 (N_38553,N_38296,N_38419);
nor U38554 (N_38554,N_38484,N_38276);
xnor U38555 (N_38555,N_38308,N_38306);
and U38556 (N_38556,N_38415,N_38407);
nand U38557 (N_38557,N_38316,N_38290);
or U38558 (N_38558,N_38364,N_38322);
and U38559 (N_38559,N_38274,N_38263);
or U38560 (N_38560,N_38266,N_38256);
or U38561 (N_38561,N_38314,N_38312);
nand U38562 (N_38562,N_38261,N_38427);
nand U38563 (N_38563,N_38287,N_38410);
or U38564 (N_38564,N_38280,N_38476);
nor U38565 (N_38565,N_38372,N_38397);
and U38566 (N_38566,N_38464,N_38466);
xor U38567 (N_38567,N_38418,N_38253);
and U38568 (N_38568,N_38392,N_38378);
xor U38569 (N_38569,N_38269,N_38277);
or U38570 (N_38570,N_38264,N_38409);
nand U38571 (N_38571,N_38451,N_38495);
and U38572 (N_38572,N_38353,N_38458);
nor U38573 (N_38573,N_38442,N_38423);
nor U38574 (N_38574,N_38267,N_38295);
xnor U38575 (N_38575,N_38499,N_38393);
nand U38576 (N_38576,N_38298,N_38363);
xnor U38577 (N_38577,N_38356,N_38483);
and U38578 (N_38578,N_38454,N_38366);
nand U38579 (N_38579,N_38428,N_38383);
xnor U38580 (N_38580,N_38437,N_38351);
nand U38581 (N_38581,N_38283,N_38491);
nor U38582 (N_38582,N_38408,N_38497);
or U38583 (N_38583,N_38463,N_38292);
xor U38584 (N_38584,N_38346,N_38430);
xor U38585 (N_38585,N_38359,N_38465);
xnor U38586 (N_38586,N_38404,N_38288);
xor U38587 (N_38587,N_38474,N_38338);
nand U38588 (N_38588,N_38293,N_38443);
nand U38589 (N_38589,N_38473,N_38394);
nor U38590 (N_38590,N_38275,N_38398);
nand U38591 (N_38591,N_38453,N_38317);
nor U38592 (N_38592,N_38385,N_38349);
or U38593 (N_38593,N_38406,N_38354);
xor U38594 (N_38594,N_38414,N_38376);
and U38595 (N_38595,N_38325,N_38319);
or U38596 (N_38596,N_38252,N_38318);
nand U38597 (N_38597,N_38384,N_38265);
nor U38598 (N_38598,N_38439,N_38433);
nor U38599 (N_38599,N_38327,N_38447);
and U38600 (N_38600,N_38468,N_38339);
or U38601 (N_38601,N_38348,N_38469);
xor U38602 (N_38602,N_38471,N_38452);
or U38603 (N_38603,N_38467,N_38388);
and U38604 (N_38604,N_38294,N_38498);
or U38605 (N_38605,N_38493,N_38377);
xnor U38606 (N_38606,N_38490,N_38250);
and U38607 (N_38607,N_38440,N_38330);
or U38608 (N_38608,N_38297,N_38380);
xor U38609 (N_38609,N_38431,N_38361);
nand U38610 (N_38610,N_38365,N_38472);
and U38611 (N_38611,N_38342,N_38413);
nor U38612 (N_38612,N_38488,N_38300);
or U38613 (N_38613,N_38371,N_38279);
nor U38614 (N_38614,N_38478,N_38489);
and U38615 (N_38615,N_38340,N_38374);
and U38616 (N_38616,N_38289,N_38386);
nor U38617 (N_38617,N_38304,N_38373);
xnor U38618 (N_38618,N_38355,N_38335);
nand U38619 (N_38619,N_38259,N_38422);
nor U38620 (N_38620,N_38421,N_38399);
xnor U38621 (N_38621,N_38345,N_38429);
nand U38622 (N_38622,N_38424,N_38368);
or U38623 (N_38623,N_38370,N_38323);
nand U38624 (N_38624,N_38336,N_38278);
nor U38625 (N_38625,N_38493,N_38323);
or U38626 (N_38626,N_38391,N_38483);
xnor U38627 (N_38627,N_38387,N_38374);
or U38628 (N_38628,N_38453,N_38337);
nor U38629 (N_38629,N_38443,N_38472);
and U38630 (N_38630,N_38252,N_38436);
and U38631 (N_38631,N_38337,N_38276);
nand U38632 (N_38632,N_38383,N_38265);
nand U38633 (N_38633,N_38255,N_38467);
and U38634 (N_38634,N_38444,N_38457);
xor U38635 (N_38635,N_38267,N_38485);
nor U38636 (N_38636,N_38409,N_38355);
xor U38637 (N_38637,N_38442,N_38263);
xor U38638 (N_38638,N_38495,N_38441);
nand U38639 (N_38639,N_38390,N_38452);
nand U38640 (N_38640,N_38312,N_38281);
and U38641 (N_38641,N_38391,N_38325);
or U38642 (N_38642,N_38345,N_38251);
or U38643 (N_38643,N_38294,N_38363);
nor U38644 (N_38644,N_38386,N_38336);
and U38645 (N_38645,N_38394,N_38326);
nor U38646 (N_38646,N_38417,N_38457);
and U38647 (N_38647,N_38296,N_38376);
xnor U38648 (N_38648,N_38299,N_38421);
and U38649 (N_38649,N_38267,N_38440);
nor U38650 (N_38650,N_38316,N_38450);
and U38651 (N_38651,N_38264,N_38446);
and U38652 (N_38652,N_38469,N_38389);
xor U38653 (N_38653,N_38275,N_38484);
or U38654 (N_38654,N_38265,N_38339);
xor U38655 (N_38655,N_38348,N_38405);
xnor U38656 (N_38656,N_38311,N_38458);
xnor U38657 (N_38657,N_38486,N_38361);
nand U38658 (N_38658,N_38463,N_38428);
nand U38659 (N_38659,N_38352,N_38389);
nor U38660 (N_38660,N_38499,N_38383);
nor U38661 (N_38661,N_38431,N_38490);
nor U38662 (N_38662,N_38390,N_38458);
nor U38663 (N_38663,N_38330,N_38452);
and U38664 (N_38664,N_38486,N_38491);
xor U38665 (N_38665,N_38406,N_38317);
and U38666 (N_38666,N_38357,N_38305);
xor U38667 (N_38667,N_38278,N_38328);
nand U38668 (N_38668,N_38385,N_38420);
and U38669 (N_38669,N_38376,N_38254);
xnor U38670 (N_38670,N_38386,N_38301);
and U38671 (N_38671,N_38342,N_38276);
xnor U38672 (N_38672,N_38331,N_38315);
nor U38673 (N_38673,N_38317,N_38441);
nand U38674 (N_38674,N_38256,N_38312);
xor U38675 (N_38675,N_38424,N_38363);
nor U38676 (N_38676,N_38417,N_38287);
nand U38677 (N_38677,N_38461,N_38455);
and U38678 (N_38678,N_38321,N_38410);
nand U38679 (N_38679,N_38253,N_38365);
nor U38680 (N_38680,N_38268,N_38335);
nor U38681 (N_38681,N_38435,N_38439);
and U38682 (N_38682,N_38395,N_38440);
or U38683 (N_38683,N_38374,N_38343);
or U38684 (N_38684,N_38364,N_38403);
xor U38685 (N_38685,N_38263,N_38371);
xor U38686 (N_38686,N_38327,N_38338);
or U38687 (N_38687,N_38400,N_38404);
or U38688 (N_38688,N_38368,N_38342);
nor U38689 (N_38689,N_38416,N_38262);
and U38690 (N_38690,N_38378,N_38410);
nor U38691 (N_38691,N_38289,N_38360);
or U38692 (N_38692,N_38327,N_38448);
nor U38693 (N_38693,N_38496,N_38444);
nor U38694 (N_38694,N_38260,N_38285);
xnor U38695 (N_38695,N_38489,N_38305);
and U38696 (N_38696,N_38266,N_38433);
nor U38697 (N_38697,N_38474,N_38499);
and U38698 (N_38698,N_38338,N_38321);
and U38699 (N_38699,N_38381,N_38272);
xnor U38700 (N_38700,N_38431,N_38266);
or U38701 (N_38701,N_38303,N_38396);
xor U38702 (N_38702,N_38389,N_38344);
nor U38703 (N_38703,N_38446,N_38256);
xor U38704 (N_38704,N_38482,N_38253);
and U38705 (N_38705,N_38493,N_38440);
nor U38706 (N_38706,N_38324,N_38344);
nor U38707 (N_38707,N_38375,N_38302);
and U38708 (N_38708,N_38288,N_38365);
or U38709 (N_38709,N_38451,N_38471);
and U38710 (N_38710,N_38449,N_38450);
nand U38711 (N_38711,N_38422,N_38404);
nand U38712 (N_38712,N_38307,N_38411);
and U38713 (N_38713,N_38467,N_38333);
and U38714 (N_38714,N_38254,N_38280);
and U38715 (N_38715,N_38323,N_38253);
or U38716 (N_38716,N_38493,N_38463);
or U38717 (N_38717,N_38434,N_38449);
xor U38718 (N_38718,N_38293,N_38426);
and U38719 (N_38719,N_38276,N_38457);
or U38720 (N_38720,N_38420,N_38404);
or U38721 (N_38721,N_38368,N_38289);
xnor U38722 (N_38722,N_38300,N_38360);
xor U38723 (N_38723,N_38414,N_38313);
nor U38724 (N_38724,N_38256,N_38298);
or U38725 (N_38725,N_38398,N_38252);
xor U38726 (N_38726,N_38349,N_38424);
or U38727 (N_38727,N_38347,N_38476);
or U38728 (N_38728,N_38444,N_38298);
nand U38729 (N_38729,N_38373,N_38404);
nand U38730 (N_38730,N_38268,N_38326);
or U38731 (N_38731,N_38454,N_38427);
xor U38732 (N_38732,N_38315,N_38356);
nor U38733 (N_38733,N_38354,N_38393);
or U38734 (N_38734,N_38260,N_38368);
or U38735 (N_38735,N_38253,N_38343);
and U38736 (N_38736,N_38459,N_38367);
nor U38737 (N_38737,N_38396,N_38290);
and U38738 (N_38738,N_38392,N_38301);
nor U38739 (N_38739,N_38260,N_38315);
nand U38740 (N_38740,N_38373,N_38397);
nor U38741 (N_38741,N_38301,N_38400);
nor U38742 (N_38742,N_38499,N_38451);
nor U38743 (N_38743,N_38447,N_38276);
nand U38744 (N_38744,N_38371,N_38304);
or U38745 (N_38745,N_38304,N_38385);
and U38746 (N_38746,N_38448,N_38376);
nand U38747 (N_38747,N_38411,N_38294);
xnor U38748 (N_38748,N_38453,N_38339);
and U38749 (N_38749,N_38285,N_38415);
and U38750 (N_38750,N_38532,N_38738);
xnor U38751 (N_38751,N_38719,N_38507);
or U38752 (N_38752,N_38638,N_38525);
nand U38753 (N_38753,N_38724,N_38655);
nor U38754 (N_38754,N_38708,N_38650);
and U38755 (N_38755,N_38583,N_38611);
xnor U38756 (N_38756,N_38653,N_38615);
nand U38757 (N_38757,N_38586,N_38558);
xor U38758 (N_38758,N_38718,N_38517);
nand U38759 (N_38759,N_38502,N_38610);
nand U38760 (N_38760,N_38590,N_38698);
xor U38761 (N_38761,N_38622,N_38559);
or U38762 (N_38762,N_38690,N_38671);
nor U38763 (N_38763,N_38736,N_38699);
and U38764 (N_38764,N_38514,N_38619);
and U38765 (N_38765,N_38733,N_38585);
and U38766 (N_38766,N_38601,N_38503);
nor U38767 (N_38767,N_38509,N_38549);
nand U38768 (N_38768,N_38598,N_38554);
nor U38769 (N_38769,N_38665,N_38526);
or U38770 (N_38770,N_38578,N_38540);
nor U38771 (N_38771,N_38702,N_38714);
nor U38772 (N_38772,N_38537,N_38542);
nor U38773 (N_38773,N_38621,N_38584);
xor U38774 (N_38774,N_38544,N_38745);
and U38775 (N_38775,N_38734,N_38508);
nor U38776 (N_38776,N_38592,N_38591);
or U38777 (N_38777,N_38685,N_38747);
and U38778 (N_38778,N_38669,N_38641);
xnor U38779 (N_38779,N_38528,N_38726);
or U38780 (N_38780,N_38630,N_38723);
nor U38781 (N_38781,N_38531,N_38553);
xor U38782 (N_38782,N_38575,N_38687);
nor U38783 (N_38783,N_38634,N_38717);
xor U38784 (N_38784,N_38709,N_38602);
and U38785 (N_38785,N_38577,N_38651);
nor U38786 (N_38786,N_38605,N_38694);
or U38787 (N_38787,N_38656,N_38614);
xor U38788 (N_38788,N_38612,N_38649);
and U38789 (N_38789,N_38692,N_38530);
nor U38790 (N_38790,N_38710,N_38574);
or U38791 (N_38791,N_38555,N_38548);
nand U38792 (N_38792,N_38659,N_38712);
nand U38793 (N_38793,N_38501,N_38588);
nand U38794 (N_38794,N_38551,N_38679);
nand U38795 (N_38795,N_38515,N_38565);
nand U38796 (N_38796,N_38620,N_38654);
nor U38797 (N_38797,N_38676,N_38682);
and U38798 (N_38798,N_38701,N_38737);
or U38799 (N_38799,N_38607,N_38599);
nor U38800 (N_38800,N_38730,N_38552);
xnor U38801 (N_38801,N_38557,N_38568);
nor U38802 (N_38802,N_38686,N_38522);
and U38803 (N_38803,N_38543,N_38510);
nor U38804 (N_38804,N_38604,N_38563);
nand U38805 (N_38805,N_38561,N_38697);
nand U38806 (N_38806,N_38681,N_38519);
xor U38807 (N_38807,N_38729,N_38623);
nor U38808 (N_38808,N_38600,N_38646);
and U38809 (N_38809,N_38547,N_38504);
nand U38810 (N_38810,N_38579,N_38617);
nand U38811 (N_38811,N_38633,N_38707);
nor U38812 (N_38812,N_38523,N_38550);
nor U38813 (N_38813,N_38739,N_38566);
nor U38814 (N_38814,N_38742,N_38720);
or U38815 (N_38815,N_38713,N_38541);
or U38816 (N_38816,N_38748,N_38673);
or U38817 (N_38817,N_38564,N_38683);
nor U38818 (N_38818,N_38597,N_38658);
nand U38819 (N_38819,N_38631,N_38722);
nand U38820 (N_38820,N_38688,N_38652);
or U38821 (N_38821,N_38596,N_38572);
xor U38822 (N_38822,N_38516,N_38664);
xnor U38823 (N_38823,N_38626,N_38663);
or U38824 (N_38824,N_38520,N_38589);
and U38825 (N_38825,N_38594,N_38632);
nor U38826 (N_38826,N_38741,N_38715);
nand U38827 (N_38827,N_38538,N_38573);
nor U38828 (N_38828,N_38533,N_38666);
and U38829 (N_38829,N_38524,N_38735);
nand U38830 (N_38830,N_38582,N_38672);
and U38831 (N_38831,N_38642,N_38529);
or U38832 (N_38832,N_38645,N_38731);
and U38833 (N_38833,N_38680,N_38625);
nor U38834 (N_38834,N_38567,N_38576);
nor U38835 (N_38835,N_38647,N_38521);
nor U38836 (N_38836,N_38661,N_38662);
xnor U38837 (N_38837,N_38624,N_38640);
nand U38838 (N_38838,N_38580,N_38744);
nand U38839 (N_38839,N_38500,N_38616);
and U38840 (N_38840,N_38581,N_38684);
nand U38841 (N_38841,N_38705,N_38570);
nor U38842 (N_38842,N_38637,N_38693);
xor U38843 (N_38843,N_38506,N_38691);
nor U38844 (N_38844,N_38536,N_38546);
nor U38845 (N_38845,N_38706,N_38534);
and U38846 (N_38846,N_38527,N_38556);
and U38847 (N_38847,N_38535,N_38603);
and U38848 (N_38848,N_38657,N_38696);
nor U38849 (N_38849,N_38667,N_38518);
nor U38850 (N_38850,N_38749,N_38618);
nand U38851 (N_38851,N_38727,N_38593);
and U38852 (N_38852,N_38716,N_38677);
nor U38853 (N_38853,N_38627,N_38613);
nor U38854 (N_38854,N_38595,N_38700);
xor U38855 (N_38855,N_38704,N_38674);
or U38856 (N_38856,N_38608,N_38636);
or U38857 (N_38857,N_38628,N_38629);
or U38858 (N_38858,N_38703,N_38511);
and U38859 (N_38859,N_38689,N_38505);
or U38860 (N_38860,N_38635,N_38675);
nand U38861 (N_38861,N_38644,N_38639);
or U38862 (N_38862,N_38678,N_38660);
and U38863 (N_38863,N_38569,N_38670);
nor U38864 (N_38864,N_38740,N_38513);
or U38865 (N_38865,N_38562,N_38721);
nand U38866 (N_38866,N_38606,N_38609);
nor U38867 (N_38867,N_38725,N_38587);
nand U38868 (N_38868,N_38539,N_38746);
nand U38869 (N_38869,N_38711,N_38648);
and U38870 (N_38870,N_38512,N_38571);
or U38871 (N_38871,N_38643,N_38668);
xor U38872 (N_38872,N_38743,N_38545);
and U38873 (N_38873,N_38728,N_38695);
nand U38874 (N_38874,N_38732,N_38560);
or U38875 (N_38875,N_38605,N_38581);
nor U38876 (N_38876,N_38728,N_38503);
nor U38877 (N_38877,N_38677,N_38523);
and U38878 (N_38878,N_38569,N_38553);
nand U38879 (N_38879,N_38712,N_38685);
or U38880 (N_38880,N_38733,N_38617);
nand U38881 (N_38881,N_38740,N_38542);
xor U38882 (N_38882,N_38705,N_38547);
nor U38883 (N_38883,N_38735,N_38538);
nor U38884 (N_38884,N_38708,N_38586);
xnor U38885 (N_38885,N_38700,N_38648);
xnor U38886 (N_38886,N_38601,N_38659);
xor U38887 (N_38887,N_38730,N_38684);
nand U38888 (N_38888,N_38515,N_38649);
xor U38889 (N_38889,N_38561,N_38589);
and U38890 (N_38890,N_38642,N_38744);
nand U38891 (N_38891,N_38576,N_38748);
and U38892 (N_38892,N_38528,N_38567);
xnor U38893 (N_38893,N_38588,N_38631);
nand U38894 (N_38894,N_38593,N_38709);
nor U38895 (N_38895,N_38704,N_38517);
xnor U38896 (N_38896,N_38568,N_38587);
xor U38897 (N_38897,N_38703,N_38563);
xor U38898 (N_38898,N_38581,N_38693);
or U38899 (N_38899,N_38602,N_38685);
nor U38900 (N_38900,N_38729,N_38563);
nor U38901 (N_38901,N_38513,N_38682);
nand U38902 (N_38902,N_38548,N_38716);
xor U38903 (N_38903,N_38663,N_38711);
and U38904 (N_38904,N_38537,N_38627);
nor U38905 (N_38905,N_38718,N_38567);
nor U38906 (N_38906,N_38598,N_38550);
nor U38907 (N_38907,N_38709,N_38557);
nor U38908 (N_38908,N_38571,N_38646);
nand U38909 (N_38909,N_38670,N_38627);
nor U38910 (N_38910,N_38686,N_38534);
xor U38911 (N_38911,N_38628,N_38501);
xor U38912 (N_38912,N_38511,N_38628);
xor U38913 (N_38913,N_38643,N_38594);
nand U38914 (N_38914,N_38596,N_38542);
or U38915 (N_38915,N_38727,N_38573);
xnor U38916 (N_38916,N_38635,N_38620);
and U38917 (N_38917,N_38507,N_38724);
or U38918 (N_38918,N_38548,N_38543);
or U38919 (N_38919,N_38507,N_38632);
nor U38920 (N_38920,N_38633,N_38567);
xor U38921 (N_38921,N_38542,N_38509);
xor U38922 (N_38922,N_38636,N_38683);
and U38923 (N_38923,N_38588,N_38636);
nand U38924 (N_38924,N_38746,N_38723);
xnor U38925 (N_38925,N_38541,N_38630);
or U38926 (N_38926,N_38647,N_38666);
xnor U38927 (N_38927,N_38716,N_38730);
xnor U38928 (N_38928,N_38513,N_38748);
or U38929 (N_38929,N_38521,N_38628);
or U38930 (N_38930,N_38571,N_38740);
or U38931 (N_38931,N_38725,N_38562);
or U38932 (N_38932,N_38617,N_38687);
nand U38933 (N_38933,N_38727,N_38650);
nand U38934 (N_38934,N_38588,N_38598);
or U38935 (N_38935,N_38747,N_38642);
or U38936 (N_38936,N_38526,N_38668);
and U38937 (N_38937,N_38725,N_38583);
nor U38938 (N_38938,N_38629,N_38610);
nor U38939 (N_38939,N_38557,N_38573);
nor U38940 (N_38940,N_38530,N_38696);
or U38941 (N_38941,N_38585,N_38607);
nor U38942 (N_38942,N_38646,N_38533);
nor U38943 (N_38943,N_38522,N_38572);
or U38944 (N_38944,N_38625,N_38645);
nor U38945 (N_38945,N_38642,N_38663);
and U38946 (N_38946,N_38647,N_38551);
nand U38947 (N_38947,N_38676,N_38610);
xnor U38948 (N_38948,N_38560,N_38568);
xor U38949 (N_38949,N_38579,N_38650);
or U38950 (N_38950,N_38522,N_38550);
xnor U38951 (N_38951,N_38523,N_38538);
xor U38952 (N_38952,N_38678,N_38545);
xnor U38953 (N_38953,N_38691,N_38724);
xnor U38954 (N_38954,N_38699,N_38663);
or U38955 (N_38955,N_38563,N_38662);
nor U38956 (N_38956,N_38583,N_38737);
nand U38957 (N_38957,N_38553,N_38716);
or U38958 (N_38958,N_38613,N_38586);
and U38959 (N_38959,N_38698,N_38568);
xor U38960 (N_38960,N_38631,N_38653);
nand U38961 (N_38961,N_38521,N_38575);
nand U38962 (N_38962,N_38589,N_38636);
or U38963 (N_38963,N_38630,N_38687);
xnor U38964 (N_38964,N_38727,N_38685);
and U38965 (N_38965,N_38512,N_38537);
nor U38966 (N_38966,N_38732,N_38566);
nor U38967 (N_38967,N_38594,N_38576);
and U38968 (N_38968,N_38689,N_38532);
nor U38969 (N_38969,N_38730,N_38572);
xnor U38970 (N_38970,N_38676,N_38586);
xnor U38971 (N_38971,N_38585,N_38667);
or U38972 (N_38972,N_38524,N_38514);
xor U38973 (N_38973,N_38644,N_38731);
nand U38974 (N_38974,N_38557,N_38676);
xnor U38975 (N_38975,N_38567,N_38601);
xnor U38976 (N_38976,N_38699,N_38550);
nor U38977 (N_38977,N_38675,N_38608);
or U38978 (N_38978,N_38714,N_38616);
nand U38979 (N_38979,N_38674,N_38691);
nand U38980 (N_38980,N_38549,N_38696);
xor U38981 (N_38981,N_38679,N_38714);
nand U38982 (N_38982,N_38637,N_38741);
nor U38983 (N_38983,N_38564,N_38638);
nor U38984 (N_38984,N_38554,N_38664);
or U38985 (N_38985,N_38701,N_38514);
nor U38986 (N_38986,N_38700,N_38592);
xnor U38987 (N_38987,N_38637,N_38690);
xnor U38988 (N_38988,N_38706,N_38547);
or U38989 (N_38989,N_38704,N_38513);
and U38990 (N_38990,N_38747,N_38635);
and U38991 (N_38991,N_38600,N_38599);
nand U38992 (N_38992,N_38560,N_38657);
nand U38993 (N_38993,N_38580,N_38625);
nand U38994 (N_38994,N_38571,N_38620);
nor U38995 (N_38995,N_38665,N_38535);
nor U38996 (N_38996,N_38696,N_38601);
and U38997 (N_38997,N_38739,N_38672);
or U38998 (N_38998,N_38595,N_38663);
xor U38999 (N_38999,N_38538,N_38724);
or U39000 (N_39000,N_38965,N_38906);
and U39001 (N_39001,N_38971,N_38954);
nand U39002 (N_39002,N_38836,N_38960);
or U39003 (N_39003,N_38966,N_38963);
xor U39004 (N_39004,N_38808,N_38886);
xnor U39005 (N_39005,N_38818,N_38896);
nand U39006 (N_39006,N_38926,N_38988);
or U39007 (N_39007,N_38782,N_38761);
or U39008 (N_39008,N_38832,N_38880);
and U39009 (N_39009,N_38807,N_38969);
xor U39010 (N_39010,N_38957,N_38859);
xnor U39011 (N_39011,N_38820,N_38786);
and U39012 (N_39012,N_38947,N_38869);
xor U39013 (N_39013,N_38752,N_38772);
nand U39014 (N_39014,N_38823,N_38849);
or U39015 (N_39015,N_38821,N_38903);
nor U39016 (N_39016,N_38958,N_38937);
or U39017 (N_39017,N_38834,N_38941);
or U39018 (N_39018,N_38791,N_38853);
and U39019 (N_39019,N_38809,N_38845);
nand U39020 (N_39020,N_38928,N_38998);
or U39021 (N_39021,N_38975,N_38867);
nor U39022 (N_39022,N_38800,N_38798);
xnor U39023 (N_39023,N_38802,N_38861);
nor U39024 (N_39024,N_38992,N_38828);
xnor U39025 (N_39025,N_38913,N_38968);
and U39026 (N_39026,N_38917,N_38779);
nand U39027 (N_39027,N_38826,N_38907);
nor U39028 (N_39028,N_38938,N_38789);
xor U39029 (N_39029,N_38959,N_38863);
nor U39030 (N_39030,N_38881,N_38882);
nor U39031 (N_39031,N_38830,N_38788);
nor U39032 (N_39032,N_38945,N_38827);
xor U39033 (N_39033,N_38989,N_38891);
or U39034 (N_39034,N_38783,N_38961);
and U39035 (N_39035,N_38984,N_38936);
xor U39036 (N_39036,N_38773,N_38899);
and U39037 (N_39037,N_38905,N_38868);
and U39038 (N_39038,N_38795,N_38995);
or U39039 (N_39039,N_38805,N_38953);
or U39040 (N_39040,N_38885,N_38762);
or U39041 (N_39041,N_38876,N_38775);
and U39042 (N_39042,N_38933,N_38894);
nand U39043 (N_39043,N_38974,N_38967);
or U39044 (N_39044,N_38873,N_38750);
or U39045 (N_39045,N_38864,N_38768);
nor U39046 (N_39046,N_38996,N_38982);
or U39047 (N_39047,N_38923,N_38833);
nand U39048 (N_39048,N_38977,N_38790);
xor U39049 (N_39049,N_38858,N_38939);
and U39050 (N_39050,N_38983,N_38893);
xnor U39051 (N_39051,N_38962,N_38854);
nor U39052 (N_39052,N_38751,N_38910);
nand U39053 (N_39053,N_38878,N_38895);
xor U39054 (N_39054,N_38870,N_38806);
or U39055 (N_39055,N_38857,N_38888);
or U39056 (N_39056,N_38985,N_38892);
xor U39057 (N_39057,N_38986,N_38991);
nand U39058 (N_39058,N_38799,N_38850);
xnor U39059 (N_39059,N_38931,N_38787);
nand U39060 (N_39060,N_38980,N_38979);
nand U39061 (N_39061,N_38889,N_38897);
and U39062 (N_39062,N_38824,N_38829);
and U39063 (N_39063,N_38842,N_38841);
or U39064 (N_39064,N_38911,N_38948);
nor U39065 (N_39065,N_38813,N_38754);
xnor U39066 (N_39066,N_38976,N_38874);
nor U39067 (N_39067,N_38921,N_38908);
nand U39068 (N_39068,N_38901,N_38978);
or U39069 (N_39069,N_38848,N_38796);
xor U39070 (N_39070,N_38765,N_38835);
xnor U39071 (N_39071,N_38843,N_38943);
or U39072 (N_39072,N_38839,N_38778);
nand U39073 (N_39073,N_38914,N_38898);
and U39074 (N_39074,N_38924,N_38930);
nand U39075 (N_39075,N_38973,N_38753);
nor U39076 (N_39076,N_38970,N_38755);
or U39077 (N_39077,N_38952,N_38856);
xnor U39078 (N_39078,N_38774,N_38865);
or U39079 (N_39079,N_38797,N_38935);
nand U39080 (N_39080,N_38890,N_38916);
nand U39081 (N_39081,N_38822,N_38919);
and U39082 (N_39082,N_38776,N_38847);
or U39083 (N_39083,N_38780,N_38825);
nand U39084 (N_39084,N_38990,N_38769);
nor U39085 (N_39085,N_38883,N_38887);
nor U39086 (N_39086,N_38994,N_38840);
and U39087 (N_39087,N_38815,N_38942);
or U39088 (N_39088,N_38771,N_38844);
nand U39089 (N_39089,N_38816,N_38792);
and U39090 (N_39090,N_38758,N_38875);
nand U39091 (N_39091,N_38904,N_38920);
or U39092 (N_39092,N_38810,N_38987);
xnor U39093 (N_39093,N_38803,N_38909);
xor U39094 (N_39094,N_38794,N_38927);
nor U39095 (N_39095,N_38872,N_38918);
and U39096 (N_39096,N_38767,N_38946);
xor U39097 (N_39097,N_38756,N_38837);
nor U39098 (N_39098,N_38950,N_38932);
nor U39099 (N_39099,N_38766,N_38801);
nor U39100 (N_39100,N_38811,N_38871);
nand U39101 (N_39101,N_38993,N_38831);
nand U39102 (N_39102,N_38956,N_38866);
and U39103 (N_39103,N_38972,N_38862);
nor U39104 (N_39104,N_38804,N_38793);
and U39105 (N_39105,N_38934,N_38877);
or U39106 (N_39106,N_38940,N_38955);
and U39107 (N_39107,N_38912,N_38981);
or U39108 (N_39108,N_38785,N_38852);
and U39109 (N_39109,N_38925,N_38781);
or U39110 (N_39110,N_38879,N_38884);
and U39111 (N_39111,N_38929,N_38902);
nor U39112 (N_39112,N_38949,N_38763);
nor U39113 (N_39113,N_38951,N_38760);
xnor U39114 (N_39114,N_38997,N_38819);
nand U39115 (N_39115,N_38817,N_38855);
nand U39116 (N_39116,N_38944,N_38812);
nor U39117 (N_39117,N_38846,N_38757);
or U39118 (N_39118,N_38814,N_38851);
or U39119 (N_39119,N_38999,N_38860);
or U39120 (N_39120,N_38770,N_38900);
nor U39121 (N_39121,N_38764,N_38922);
nand U39122 (N_39122,N_38838,N_38964);
xor U39123 (N_39123,N_38777,N_38759);
nor U39124 (N_39124,N_38784,N_38915);
or U39125 (N_39125,N_38941,N_38826);
nand U39126 (N_39126,N_38992,N_38759);
nand U39127 (N_39127,N_38756,N_38945);
and U39128 (N_39128,N_38846,N_38781);
nor U39129 (N_39129,N_38793,N_38918);
and U39130 (N_39130,N_38884,N_38820);
nor U39131 (N_39131,N_38843,N_38785);
nor U39132 (N_39132,N_38759,N_38882);
and U39133 (N_39133,N_38782,N_38827);
and U39134 (N_39134,N_38777,N_38951);
nand U39135 (N_39135,N_38784,N_38813);
or U39136 (N_39136,N_38759,N_38972);
and U39137 (N_39137,N_38935,N_38760);
nor U39138 (N_39138,N_38900,N_38788);
xor U39139 (N_39139,N_38776,N_38874);
and U39140 (N_39140,N_38944,N_38843);
and U39141 (N_39141,N_38999,N_38903);
and U39142 (N_39142,N_38988,N_38833);
nor U39143 (N_39143,N_38985,N_38914);
xor U39144 (N_39144,N_38772,N_38967);
and U39145 (N_39145,N_38979,N_38916);
nand U39146 (N_39146,N_38762,N_38781);
nand U39147 (N_39147,N_38898,N_38969);
or U39148 (N_39148,N_38997,N_38974);
nand U39149 (N_39149,N_38896,N_38948);
or U39150 (N_39150,N_38773,N_38822);
xnor U39151 (N_39151,N_38978,N_38810);
nand U39152 (N_39152,N_38785,N_38871);
nor U39153 (N_39153,N_38787,N_38975);
nor U39154 (N_39154,N_38909,N_38767);
nand U39155 (N_39155,N_38761,N_38807);
nor U39156 (N_39156,N_38867,N_38862);
or U39157 (N_39157,N_38886,N_38993);
nand U39158 (N_39158,N_38811,N_38755);
xnor U39159 (N_39159,N_38863,N_38967);
and U39160 (N_39160,N_38869,N_38910);
nor U39161 (N_39161,N_38975,N_38941);
or U39162 (N_39162,N_38939,N_38877);
xor U39163 (N_39163,N_38838,N_38772);
nand U39164 (N_39164,N_38930,N_38858);
or U39165 (N_39165,N_38990,N_38881);
nor U39166 (N_39166,N_38914,N_38875);
xnor U39167 (N_39167,N_38768,N_38805);
xnor U39168 (N_39168,N_38785,N_38798);
nand U39169 (N_39169,N_38849,N_38984);
or U39170 (N_39170,N_38862,N_38894);
or U39171 (N_39171,N_38853,N_38769);
xor U39172 (N_39172,N_38782,N_38992);
nor U39173 (N_39173,N_38871,N_38836);
nor U39174 (N_39174,N_38971,N_38920);
or U39175 (N_39175,N_38839,N_38755);
nand U39176 (N_39176,N_38962,N_38804);
or U39177 (N_39177,N_38897,N_38826);
nand U39178 (N_39178,N_38769,N_38852);
xor U39179 (N_39179,N_38894,N_38826);
nor U39180 (N_39180,N_38840,N_38784);
and U39181 (N_39181,N_38781,N_38993);
xor U39182 (N_39182,N_38923,N_38870);
nor U39183 (N_39183,N_38879,N_38943);
nor U39184 (N_39184,N_38973,N_38852);
or U39185 (N_39185,N_38863,N_38818);
nor U39186 (N_39186,N_38819,N_38845);
xnor U39187 (N_39187,N_38800,N_38899);
xnor U39188 (N_39188,N_38900,N_38815);
xnor U39189 (N_39189,N_38794,N_38857);
and U39190 (N_39190,N_38822,N_38802);
xor U39191 (N_39191,N_38869,N_38763);
or U39192 (N_39192,N_38754,N_38818);
or U39193 (N_39193,N_38827,N_38882);
nor U39194 (N_39194,N_38796,N_38934);
nor U39195 (N_39195,N_38825,N_38776);
nand U39196 (N_39196,N_38878,N_38811);
xor U39197 (N_39197,N_38967,N_38812);
nand U39198 (N_39198,N_38971,N_38772);
or U39199 (N_39199,N_38758,N_38833);
xor U39200 (N_39200,N_38781,N_38878);
nand U39201 (N_39201,N_38818,N_38884);
or U39202 (N_39202,N_38877,N_38881);
or U39203 (N_39203,N_38977,N_38842);
or U39204 (N_39204,N_38804,N_38945);
xnor U39205 (N_39205,N_38930,N_38995);
nor U39206 (N_39206,N_38982,N_38986);
nand U39207 (N_39207,N_38777,N_38809);
or U39208 (N_39208,N_38923,N_38753);
and U39209 (N_39209,N_38944,N_38873);
or U39210 (N_39210,N_38959,N_38864);
and U39211 (N_39211,N_38864,N_38809);
nor U39212 (N_39212,N_38978,N_38984);
and U39213 (N_39213,N_38982,N_38845);
xor U39214 (N_39214,N_38865,N_38832);
and U39215 (N_39215,N_38875,N_38865);
nand U39216 (N_39216,N_38959,N_38907);
nand U39217 (N_39217,N_38890,N_38935);
xor U39218 (N_39218,N_38770,N_38842);
and U39219 (N_39219,N_38823,N_38884);
and U39220 (N_39220,N_38805,N_38846);
nor U39221 (N_39221,N_38935,N_38958);
nor U39222 (N_39222,N_38976,N_38937);
nor U39223 (N_39223,N_38793,N_38895);
xor U39224 (N_39224,N_38820,N_38844);
and U39225 (N_39225,N_38955,N_38902);
nor U39226 (N_39226,N_38846,N_38933);
or U39227 (N_39227,N_38855,N_38791);
xnor U39228 (N_39228,N_38973,N_38995);
xor U39229 (N_39229,N_38830,N_38941);
nand U39230 (N_39230,N_38814,N_38773);
or U39231 (N_39231,N_38990,N_38883);
xor U39232 (N_39232,N_38791,N_38816);
nand U39233 (N_39233,N_38802,N_38767);
or U39234 (N_39234,N_38776,N_38906);
and U39235 (N_39235,N_38987,N_38819);
or U39236 (N_39236,N_38984,N_38769);
nand U39237 (N_39237,N_38998,N_38973);
or U39238 (N_39238,N_38855,N_38823);
nand U39239 (N_39239,N_38850,N_38789);
xnor U39240 (N_39240,N_38776,N_38974);
nand U39241 (N_39241,N_38842,N_38822);
nor U39242 (N_39242,N_38815,N_38831);
xor U39243 (N_39243,N_38885,N_38777);
or U39244 (N_39244,N_38830,N_38969);
or U39245 (N_39245,N_38786,N_38764);
nand U39246 (N_39246,N_38778,N_38991);
xnor U39247 (N_39247,N_38942,N_38852);
nor U39248 (N_39248,N_38953,N_38978);
or U39249 (N_39249,N_38963,N_38930);
and U39250 (N_39250,N_39018,N_39119);
nand U39251 (N_39251,N_39003,N_39170);
xor U39252 (N_39252,N_39110,N_39057);
and U39253 (N_39253,N_39117,N_39077);
xor U39254 (N_39254,N_39213,N_39235);
xnor U39255 (N_39255,N_39061,N_39001);
nand U39256 (N_39256,N_39104,N_39016);
xnor U39257 (N_39257,N_39132,N_39115);
xnor U39258 (N_39258,N_39042,N_39010);
xor U39259 (N_39259,N_39015,N_39140);
and U39260 (N_39260,N_39126,N_39118);
xnor U39261 (N_39261,N_39175,N_39208);
or U39262 (N_39262,N_39070,N_39066);
nor U39263 (N_39263,N_39187,N_39091);
nand U39264 (N_39264,N_39123,N_39093);
nand U39265 (N_39265,N_39095,N_39108);
xnor U39266 (N_39266,N_39114,N_39034);
xor U39267 (N_39267,N_39197,N_39186);
nor U39268 (N_39268,N_39172,N_39142);
or U39269 (N_39269,N_39190,N_39098);
nand U39270 (N_39270,N_39072,N_39151);
xnor U39271 (N_39271,N_39153,N_39165);
and U39272 (N_39272,N_39136,N_39158);
nand U39273 (N_39273,N_39162,N_39031);
and U39274 (N_39274,N_39097,N_39074);
nand U39275 (N_39275,N_39244,N_39124);
and U39276 (N_39276,N_39221,N_39207);
nand U39277 (N_39277,N_39234,N_39183);
or U39278 (N_39278,N_39032,N_39089);
and U39279 (N_39279,N_39028,N_39182);
xor U39280 (N_39280,N_39169,N_39176);
or U39281 (N_39281,N_39198,N_39164);
xnor U39282 (N_39282,N_39026,N_39071);
xor U39283 (N_39283,N_39203,N_39243);
nor U39284 (N_39284,N_39025,N_39065);
nor U39285 (N_39285,N_39000,N_39079);
nand U39286 (N_39286,N_39080,N_39191);
nand U39287 (N_39287,N_39086,N_39111);
or U39288 (N_39288,N_39146,N_39092);
nor U39289 (N_39289,N_39109,N_39017);
and U39290 (N_39290,N_39129,N_39180);
nor U39291 (N_39291,N_39055,N_39178);
nand U39292 (N_39292,N_39037,N_39006);
xor U39293 (N_39293,N_39100,N_39116);
nand U39294 (N_39294,N_39033,N_39036);
xnor U39295 (N_39295,N_39241,N_39168);
nand U39296 (N_39296,N_39240,N_39131);
and U39297 (N_39297,N_39143,N_39013);
or U39298 (N_39298,N_39210,N_39189);
xnor U39299 (N_39299,N_39149,N_39035);
and U39300 (N_39300,N_39053,N_39029);
nor U39301 (N_39301,N_39027,N_39075);
or U39302 (N_39302,N_39192,N_39030);
and U39303 (N_39303,N_39051,N_39023);
nor U39304 (N_39304,N_39247,N_39159);
xor U39305 (N_39305,N_39217,N_39148);
and U39306 (N_39306,N_39007,N_39046);
nand U39307 (N_39307,N_39056,N_39204);
nand U39308 (N_39308,N_39139,N_39201);
nand U39309 (N_39309,N_39248,N_39096);
xnor U39310 (N_39310,N_39008,N_39113);
and U39311 (N_39311,N_39038,N_39084);
xnor U39312 (N_39312,N_39069,N_39009);
and U39313 (N_39313,N_39060,N_39152);
nand U39314 (N_39314,N_39102,N_39232);
and U39315 (N_39315,N_39237,N_39068);
and U39316 (N_39316,N_39157,N_39233);
nand U39317 (N_39317,N_39228,N_39177);
xnor U39318 (N_39318,N_39230,N_39044);
and U39319 (N_39319,N_39231,N_39181);
and U39320 (N_39320,N_39019,N_39155);
xnor U39321 (N_39321,N_39206,N_39141);
nand U39322 (N_39322,N_39128,N_39227);
and U39323 (N_39323,N_39112,N_39054);
nand U39324 (N_39324,N_39021,N_39225);
nor U39325 (N_39325,N_39052,N_39099);
or U39326 (N_39326,N_39200,N_39076);
and U39327 (N_39327,N_39196,N_39226);
nand U39328 (N_39328,N_39211,N_39167);
nor U39329 (N_39329,N_39024,N_39082);
nor U39330 (N_39330,N_39238,N_39105);
nor U39331 (N_39331,N_39045,N_39064);
xnor U39332 (N_39332,N_39094,N_39249);
and U39333 (N_39333,N_39004,N_39145);
xnor U39334 (N_39334,N_39050,N_39067);
and U39335 (N_39335,N_39011,N_39125);
and U39336 (N_39336,N_39216,N_39135);
nand U39337 (N_39337,N_39043,N_39088);
nand U39338 (N_39338,N_39107,N_39040);
and U39339 (N_39339,N_39130,N_39202);
or U39340 (N_39340,N_39085,N_39188);
xor U39341 (N_39341,N_39002,N_39224);
or U39342 (N_39342,N_39138,N_39209);
or U39343 (N_39343,N_39222,N_39184);
and U39344 (N_39344,N_39242,N_39144);
xor U39345 (N_39345,N_39012,N_39121);
or U39346 (N_39346,N_39205,N_39137);
and U39347 (N_39347,N_39062,N_39020);
nor U39348 (N_39348,N_39150,N_39087);
nor U39349 (N_39349,N_39049,N_39171);
and U39350 (N_39350,N_39101,N_39236);
nand U39351 (N_39351,N_39134,N_39154);
xnor U39352 (N_39352,N_39223,N_39173);
or U39353 (N_39353,N_39185,N_39147);
xnor U39354 (N_39354,N_39199,N_39058);
or U39355 (N_39355,N_39106,N_39219);
nor U39356 (N_39356,N_39047,N_39078);
xor U39357 (N_39357,N_39127,N_39059);
or U39358 (N_39358,N_39161,N_39103);
xnor U39359 (N_39359,N_39220,N_39214);
nor U39360 (N_39360,N_39212,N_39041);
and U39361 (N_39361,N_39179,N_39083);
and U39362 (N_39362,N_39156,N_39193);
xor U39363 (N_39363,N_39039,N_39081);
or U39364 (N_39364,N_39215,N_39120);
or U39365 (N_39365,N_39133,N_39163);
or U39366 (N_39366,N_39229,N_39073);
and U39367 (N_39367,N_39014,N_39245);
nor U39368 (N_39368,N_39090,N_39005);
nand U39369 (N_39369,N_39174,N_39239);
nand U39370 (N_39370,N_39022,N_39195);
nor U39371 (N_39371,N_39246,N_39048);
or U39372 (N_39372,N_39063,N_39218);
xor U39373 (N_39373,N_39194,N_39122);
and U39374 (N_39374,N_39166,N_39160);
xor U39375 (N_39375,N_39046,N_39131);
and U39376 (N_39376,N_39141,N_39026);
nor U39377 (N_39377,N_39228,N_39236);
or U39378 (N_39378,N_39087,N_39202);
and U39379 (N_39379,N_39109,N_39181);
nand U39380 (N_39380,N_39002,N_39142);
xnor U39381 (N_39381,N_39238,N_39107);
and U39382 (N_39382,N_39106,N_39063);
nand U39383 (N_39383,N_39181,N_39087);
or U39384 (N_39384,N_39141,N_39005);
nor U39385 (N_39385,N_39122,N_39111);
xnor U39386 (N_39386,N_39026,N_39010);
and U39387 (N_39387,N_39024,N_39140);
or U39388 (N_39388,N_39005,N_39162);
nand U39389 (N_39389,N_39026,N_39074);
or U39390 (N_39390,N_39036,N_39235);
nor U39391 (N_39391,N_39211,N_39094);
or U39392 (N_39392,N_39003,N_39156);
nor U39393 (N_39393,N_39239,N_39237);
xnor U39394 (N_39394,N_39124,N_39064);
nor U39395 (N_39395,N_39184,N_39175);
nand U39396 (N_39396,N_39064,N_39178);
nor U39397 (N_39397,N_39055,N_39023);
nor U39398 (N_39398,N_39243,N_39210);
or U39399 (N_39399,N_39026,N_39100);
or U39400 (N_39400,N_39104,N_39207);
or U39401 (N_39401,N_39235,N_39216);
nor U39402 (N_39402,N_39233,N_39215);
nand U39403 (N_39403,N_39201,N_39174);
xor U39404 (N_39404,N_39213,N_39224);
nor U39405 (N_39405,N_39247,N_39108);
xor U39406 (N_39406,N_39148,N_39031);
or U39407 (N_39407,N_39079,N_39248);
or U39408 (N_39408,N_39177,N_39049);
nand U39409 (N_39409,N_39040,N_39080);
or U39410 (N_39410,N_39081,N_39095);
nand U39411 (N_39411,N_39093,N_39133);
or U39412 (N_39412,N_39073,N_39131);
or U39413 (N_39413,N_39176,N_39139);
or U39414 (N_39414,N_39156,N_39061);
and U39415 (N_39415,N_39151,N_39057);
or U39416 (N_39416,N_39190,N_39249);
nand U39417 (N_39417,N_39240,N_39072);
nor U39418 (N_39418,N_39149,N_39008);
nand U39419 (N_39419,N_39156,N_39098);
nor U39420 (N_39420,N_39241,N_39210);
or U39421 (N_39421,N_39070,N_39118);
xor U39422 (N_39422,N_39030,N_39013);
or U39423 (N_39423,N_39216,N_39212);
xnor U39424 (N_39424,N_39181,N_39005);
nor U39425 (N_39425,N_39027,N_39193);
or U39426 (N_39426,N_39226,N_39028);
xnor U39427 (N_39427,N_39041,N_39106);
xnor U39428 (N_39428,N_39248,N_39054);
xnor U39429 (N_39429,N_39198,N_39244);
xor U39430 (N_39430,N_39070,N_39041);
nand U39431 (N_39431,N_39143,N_39133);
nor U39432 (N_39432,N_39195,N_39245);
or U39433 (N_39433,N_39209,N_39059);
or U39434 (N_39434,N_39017,N_39082);
or U39435 (N_39435,N_39004,N_39168);
nor U39436 (N_39436,N_39091,N_39046);
and U39437 (N_39437,N_39094,N_39028);
nand U39438 (N_39438,N_39182,N_39134);
nand U39439 (N_39439,N_39046,N_39064);
or U39440 (N_39440,N_39062,N_39016);
xnor U39441 (N_39441,N_39142,N_39071);
and U39442 (N_39442,N_39096,N_39040);
xnor U39443 (N_39443,N_39136,N_39170);
nand U39444 (N_39444,N_39035,N_39027);
xor U39445 (N_39445,N_39116,N_39180);
nand U39446 (N_39446,N_39082,N_39145);
or U39447 (N_39447,N_39080,N_39136);
nor U39448 (N_39448,N_39227,N_39147);
nor U39449 (N_39449,N_39098,N_39149);
nor U39450 (N_39450,N_39143,N_39166);
nand U39451 (N_39451,N_39166,N_39211);
and U39452 (N_39452,N_39079,N_39216);
nand U39453 (N_39453,N_39222,N_39204);
xnor U39454 (N_39454,N_39022,N_39172);
nand U39455 (N_39455,N_39017,N_39105);
or U39456 (N_39456,N_39016,N_39095);
nor U39457 (N_39457,N_39238,N_39078);
or U39458 (N_39458,N_39177,N_39111);
xor U39459 (N_39459,N_39143,N_39208);
or U39460 (N_39460,N_39022,N_39207);
and U39461 (N_39461,N_39040,N_39115);
or U39462 (N_39462,N_39128,N_39087);
and U39463 (N_39463,N_39186,N_39118);
xnor U39464 (N_39464,N_39189,N_39233);
nor U39465 (N_39465,N_39112,N_39219);
xor U39466 (N_39466,N_39124,N_39174);
xnor U39467 (N_39467,N_39127,N_39056);
nand U39468 (N_39468,N_39088,N_39079);
xnor U39469 (N_39469,N_39041,N_39125);
or U39470 (N_39470,N_39090,N_39214);
nor U39471 (N_39471,N_39225,N_39001);
xnor U39472 (N_39472,N_39121,N_39073);
nand U39473 (N_39473,N_39222,N_39121);
or U39474 (N_39474,N_39139,N_39110);
xnor U39475 (N_39475,N_39112,N_39151);
or U39476 (N_39476,N_39051,N_39208);
nand U39477 (N_39477,N_39028,N_39106);
nand U39478 (N_39478,N_39055,N_39088);
nor U39479 (N_39479,N_39195,N_39115);
xnor U39480 (N_39480,N_39163,N_39148);
or U39481 (N_39481,N_39152,N_39173);
xor U39482 (N_39482,N_39109,N_39227);
nand U39483 (N_39483,N_39239,N_39155);
nand U39484 (N_39484,N_39224,N_39123);
or U39485 (N_39485,N_39152,N_39020);
xnor U39486 (N_39486,N_39174,N_39209);
and U39487 (N_39487,N_39019,N_39005);
or U39488 (N_39488,N_39075,N_39195);
nand U39489 (N_39489,N_39061,N_39106);
xnor U39490 (N_39490,N_39130,N_39148);
nor U39491 (N_39491,N_39058,N_39231);
xnor U39492 (N_39492,N_39179,N_39113);
nor U39493 (N_39493,N_39016,N_39140);
nor U39494 (N_39494,N_39225,N_39149);
and U39495 (N_39495,N_39134,N_39060);
and U39496 (N_39496,N_39192,N_39068);
or U39497 (N_39497,N_39090,N_39247);
xor U39498 (N_39498,N_39064,N_39207);
and U39499 (N_39499,N_39103,N_39211);
or U39500 (N_39500,N_39265,N_39417);
nand U39501 (N_39501,N_39342,N_39469);
nand U39502 (N_39502,N_39382,N_39365);
nand U39503 (N_39503,N_39482,N_39363);
nor U39504 (N_39504,N_39443,N_39270);
xnor U39505 (N_39505,N_39376,N_39485);
nand U39506 (N_39506,N_39385,N_39471);
xnor U39507 (N_39507,N_39291,N_39466);
nor U39508 (N_39508,N_39435,N_39352);
xor U39509 (N_39509,N_39445,N_39425);
xnor U39510 (N_39510,N_39413,N_39487);
nand U39511 (N_39511,N_39398,N_39331);
nor U39512 (N_39512,N_39250,N_39344);
or U39513 (N_39513,N_39271,N_39338);
nor U39514 (N_39514,N_39419,N_39440);
xnor U39515 (N_39515,N_39492,N_39333);
nor U39516 (N_39516,N_39326,N_39493);
and U39517 (N_39517,N_39298,N_39348);
nor U39518 (N_39518,N_39422,N_39397);
and U39519 (N_39519,N_39456,N_39486);
or U39520 (N_39520,N_39438,N_39278);
xor U39521 (N_39521,N_39450,N_39394);
nand U39522 (N_39522,N_39310,N_39252);
or U39523 (N_39523,N_39304,N_39358);
and U39524 (N_39524,N_39465,N_39444);
xor U39525 (N_39525,N_39454,N_39286);
and U39526 (N_39526,N_39468,N_39288);
or U39527 (N_39527,N_39457,N_39290);
nand U39528 (N_39528,N_39459,N_39478);
or U39529 (N_39529,N_39403,N_39378);
or U39530 (N_39530,N_39476,N_39427);
nand U39531 (N_39531,N_39367,N_39295);
nor U39532 (N_39532,N_39254,N_39392);
xor U39533 (N_39533,N_39455,N_39421);
and U39534 (N_39534,N_39389,N_39449);
or U39535 (N_39535,N_39437,N_39351);
and U39536 (N_39536,N_39384,N_39386);
xor U39537 (N_39537,N_39416,N_39373);
nand U39538 (N_39538,N_39302,N_39369);
nand U39539 (N_39539,N_39280,N_39483);
nor U39540 (N_39540,N_39318,N_39350);
nor U39541 (N_39541,N_39391,N_39301);
xnor U39542 (N_39542,N_39317,N_39300);
nor U39543 (N_39543,N_39259,N_39412);
and U39544 (N_39544,N_39479,N_39266);
nor U39545 (N_39545,N_39495,N_39274);
and U39546 (N_39546,N_39383,N_39402);
xor U39547 (N_39547,N_39395,N_39433);
or U39548 (N_39548,N_39463,N_39467);
nor U39549 (N_39549,N_39251,N_39263);
or U39550 (N_39550,N_39441,N_39400);
and U39551 (N_39551,N_39299,N_39436);
xnor U39552 (N_39552,N_39303,N_39294);
or U39553 (N_39553,N_39341,N_39293);
and U39554 (N_39554,N_39349,N_39474);
nor U39555 (N_39555,N_39361,N_39289);
nor U39556 (N_39556,N_39292,N_39356);
and U39557 (N_39557,N_39374,N_39393);
xor U39558 (N_39558,N_39306,N_39336);
xor U39559 (N_39559,N_39267,N_39275);
nand U39560 (N_39560,N_39409,N_39281);
nand U39561 (N_39561,N_39264,N_39404);
xor U39562 (N_39562,N_39377,N_39327);
or U39563 (N_39563,N_39329,N_39432);
nor U39564 (N_39564,N_39381,N_39347);
xnor U39565 (N_39565,N_39484,N_39323);
or U39566 (N_39566,N_39339,N_39481);
and U39567 (N_39567,N_39460,N_39480);
and U39568 (N_39568,N_39488,N_39401);
and U39569 (N_39569,N_39362,N_39447);
or U39570 (N_39570,N_39489,N_39498);
xnor U39571 (N_39571,N_39337,N_39268);
nand U39572 (N_39572,N_39255,N_39340);
nand U39573 (N_39573,N_39388,N_39497);
nor U39574 (N_39574,N_39285,N_39313);
and U39575 (N_39575,N_39418,N_39257);
nor U39576 (N_39576,N_39330,N_39322);
or U39577 (N_39577,N_39472,N_39320);
nand U39578 (N_39578,N_39324,N_39451);
nor U39579 (N_39579,N_39387,N_39359);
and U39580 (N_39580,N_39311,N_39379);
nor U39581 (N_39581,N_39399,N_39282);
xor U39582 (N_39582,N_39496,N_39357);
or U39583 (N_39583,N_39253,N_39321);
or U39584 (N_39584,N_39284,N_39426);
nand U39585 (N_39585,N_39439,N_39410);
nand U39586 (N_39586,N_39368,N_39346);
xor U39587 (N_39587,N_39258,N_39473);
xor U39588 (N_39588,N_39325,N_39261);
and U39589 (N_39589,N_39332,N_39283);
nand U39590 (N_39590,N_39355,N_39423);
xor U39591 (N_39591,N_39434,N_39380);
and U39592 (N_39592,N_39334,N_39309);
xor U39593 (N_39593,N_39353,N_39366);
nand U39594 (N_39594,N_39354,N_39396);
nor U39595 (N_39595,N_39316,N_39272);
xnor U39596 (N_39596,N_39335,N_39328);
xnor U39597 (N_39597,N_39314,N_39370);
and U39598 (N_39598,N_39343,N_39411);
and U39599 (N_39599,N_39475,N_39319);
nor U39600 (N_39600,N_39287,N_39371);
xnor U39601 (N_39601,N_39453,N_39297);
xor U39602 (N_39602,N_39494,N_39405);
xor U39603 (N_39603,N_39452,N_39462);
and U39604 (N_39604,N_39420,N_39477);
nand U39605 (N_39605,N_39499,N_39256);
xnor U39606 (N_39606,N_39277,N_39305);
xor U39607 (N_39607,N_39407,N_39372);
nor U39608 (N_39608,N_39364,N_39260);
nand U39609 (N_39609,N_39429,N_39428);
xnor U39610 (N_39610,N_39269,N_39307);
nor U39611 (N_39611,N_39461,N_39431);
and U39612 (N_39612,N_39315,N_39308);
or U39613 (N_39613,N_39345,N_39446);
nor U39614 (N_39614,N_39279,N_39491);
nor U39615 (N_39615,N_39414,N_39458);
nand U39616 (N_39616,N_39262,N_39490);
or U39617 (N_39617,N_39312,N_39430);
nor U39618 (N_39618,N_39442,N_39390);
xnor U39619 (N_39619,N_39448,N_39424);
or U39620 (N_39620,N_39273,N_39375);
or U39621 (N_39621,N_39464,N_39415);
and U39622 (N_39622,N_39276,N_39296);
xor U39623 (N_39623,N_39406,N_39470);
and U39624 (N_39624,N_39360,N_39408);
nand U39625 (N_39625,N_39423,N_39418);
nor U39626 (N_39626,N_39364,N_39342);
nand U39627 (N_39627,N_39293,N_39357);
xnor U39628 (N_39628,N_39480,N_39266);
and U39629 (N_39629,N_39381,N_39393);
or U39630 (N_39630,N_39387,N_39280);
xor U39631 (N_39631,N_39381,N_39350);
and U39632 (N_39632,N_39369,N_39383);
xnor U39633 (N_39633,N_39441,N_39394);
or U39634 (N_39634,N_39394,N_39316);
xnor U39635 (N_39635,N_39354,N_39310);
and U39636 (N_39636,N_39372,N_39459);
nand U39637 (N_39637,N_39366,N_39418);
or U39638 (N_39638,N_39498,N_39412);
and U39639 (N_39639,N_39402,N_39328);
xor U39640 (N_39640,N_39453,N_39433);
and U39641 (N_39641,N_39354,N_39265);
and U39642 (N_39642,N_39331,N_39339);
or U39643 (N_39643,N_39317,N_39465);
nand U39644 (N_39644,N_39325,N_39327);
or U39645 (N_39645,N_39307,N_39306);
xnor U39646 (N_39646,N_39407,N_39375);
nand U39647 (N_39647,N_39499,N_39347);
nand U39648 (N_39648,N_39371,N_39383);
xor U39649 (N_39649,N_39360,N_39340);
nor U39650 (N_39650,N_39344,N_39326);
nor U39651 (N_39651,N_39328,N_39325);
nor U39652 (N_39652,N_39454,N_39346);
or U39653 (N_39653,N_39484,N_39378);
nor U39654 (N_39654,N_39409,N_39384);
xor U39655 (N_39655,N_39334,N_39257);
and U39656 (N_39656,N_39484,N_39277);
nor U39657 (N_39657,N_39302,N_39366);
xor U39658 (N_39658,N_39415,N_39277);
and U39659 (N_39659,N_39366,N_39326);
xnor U39660 (N_39660,N_39356,N_39362);
and U39661 (N_39661,N_39264,N_39498);
nand U39662 (N_39662,N_39261,N_39362);
and U39663 (N_39663,N_39267,N_39305);
nor U39664 (N_39664,N_39466,N_39467);
or U39665 (N_39665,N_39252,N_39479);
and U39666 (N_39666,N_39365,N_39395);
or U39667 (N_39667,N_39470,N_39419);
or U39668 (N_39668,N_39318,N_39287);
or U39669 (N_39669,N_39298,N_39427);
xor U39670 (N_39670,N_39279,N_39385);
and U39671 (N_39671,N_39481,N_39412);
and U39672 (N_39672,N_39433,N_39262);
and U39673 (N_39673,N_39460,N_39319);
nor U39674 (N_39674,N_39434,N_39455);
or U39675 (N_39675,N_39287,N_39445);
nor U39676 (N_39676,N_39441,N_39256);
xor U39677 (N_39677,N_39256,N_39399);
or U39678 (N_39678,N_39464,N_39413);
nand U39679 (N_39679,N_39289,N_39470);
or U39680 (N_39680,N_39280,N_39290);
and U39681 (N_39681,N_39317,N_39355);
xnor U39682 (N_39682,N_39270,N_39417);
or U39683 (N_39683,N_39428,N_39402);
or U39684 (N_39684,N_39288,N_39322);
nor U39685 (N_39685,N_39467,N_39371);
and U39686 (N_39686,N_39415,N_39298);
nor U39687 (N_39687,N_39462,N_39437);
or U39688 (N_39688,N_39332,N_39410);
or U39689 (N_39689,N_39401,N_39459);
xor U39690 (N_39690,N_39479,N_39443);
nand U39691 (N_39691,N_39380,N_39258);
and U39692 (N_39692,N_39462,N_39256);
or U39693 (N_39693,N_39465,N_39307);
or U39694 (N_39694,N_39350,N_39439);
nor U39695 (N_39695,N_39470,N_39254);
nor U39696 (N_39696,N_39288,N_39412);
nor U39697 (N_39697,N_39348,N_39326);
xor U39698 (N_39698,N_39286,N_39252);
xnor U39699 (N_39699,N_39317,N_39311);
xor U39700 (N_39700,N_39424,N_39431);
or U39701 (N_39701,N_39293,N_39345);
nor U39702 (N_39702,N_39374,N_39324);
or U39703 (N_39703,N_39345,N_39400);
or U39704 (N_39704,N_39497,N_39456);
xor U39705 (N_39705,N_39450,N_39405);
nand U39706 (N_39706,N_39496,N_39301);
and U39707 (N_39707,N_39343,N_39491);
nand U39708 (N_39708,N_39374,N_39301);
xor U39709 (N_39709,N_39398,N_39353);
nand U39710 (N_39710,N_39292,N_39481);
nand U39711 (N_39711,N_39450,N_39268);
xor U39712 (N_39712,N_39454,N_39447);
xor U39713 (N_39713,N_39252,N_39489);
xnor U39714 (N_39714,N_39480,N_39467);
or U39715 (N_39715,N_39364,N_39295);
and U39716 (N_39716,N_39453,N_39332);
nand U39717 (N_39717,N_39356,N_39297);
nand U39718 (N_39718,N_39427,N_39268);
xnor U39719 (N_39719,N_39379,N_39370);
xnor U39720 (N_39720,N_39427,N_39250);
nand U39721 (N_39721,N_39381,N_39466);
xnor U39722 (N_39722,N_39351,N_39377);
nor U39723 (N_39723,N_39336,N_39310);
xnor U39724 (N_39724,N_39411,N_39390);
and U39725 (N_39725,N_39365,N_39459);
xnor U39726 (N_39726,N_39318,N_39393);
nor U39727 (N_39727,N_39496,N_39447);
and U39728 (N_39728,N_39254,N_39361);
xor U39729 (N_39729,N_39257,N_39428);
nor U39730 (N_39730,N_39332,N_39261);
xnor U39731 (N_39731,N_39411,N_39256);
xor U39732 (N_39732,N_39361,N_39440);
or U39733 (N_39733,N_39470,N_39475);
nand U39734 (N_39734,N_39258,N_39318);
and U39735 (N_39735,N_39330,N_39286);
and U39736 (N_39736,N_39393,N_39348);
and U39737 (N_39737,N_39276,N_39378);
and U39738 (N_39738,N_39291,N_39449);
nor U39739 (N_39739,N_39297,N_39350);
or U39740 (N_39740,N_39462,N_39321);
nand U39741 (N_39741,N_39407,N_39432);
xor U39742 (N_39742,N_39392,N_39431);
nand U39743 (N_39743,N_39320,N_39398);
nand U39744 (N_39744,N_39265,N_39469);
or U39745 (N_39745,N_39487,N_39272);
and U39746 (N_39746,N_39290,N_39439);
or U39747 (N_39747,N_39368,N_39258);
or U39748 (N_39748,N_39487,N_39276);
nor U39749 (N_39749,N_39388,N_39462);
nand U39750 (N_39750,N_39719,N_39690);
nand U39751 (N_39751,N_39664,N_39706);
nor U39752 (N_39752,N_39588,N_39639);
or U39753 (N_39753,N_39655,N_39569);
xnor U39754 (N_39754,N_39711,N_39539);
and U39755 (N_39755,N_39714,N_39672);
or U39756 (N_39756,N_39651,N_39632);
xor U39757 (N_39757,N_39699,N_39529);
nand U39758 (N_39758,N_39570,N_39546);
nor U39759 (N_39759,N_39626,N_39614);
or U39760 (N_39760,N_39705,N_39702);
xnor U39761 (N_39761,N_39695,N_39741);
and U39762 (N_39762,N_39507,N_39520);
and U39763 (N_39763,N_39582,N_39662);
nand U39764 (N_39764,N_39501,N_39589);
and U39765 (N_39765,N_39506,N_39656);
nor U39766 (N_39766,N_39615,N_39528);
nor U39767 (N_39767,N_39748,N_39586);
nor U39768 (N_39768,N_39560,N_39619);
nor U39769 (N_39769,N_39658,N_39665);
nor U39770 (N_39770,N_39697,N_39727);
and U39771 (N_39771,N_39612,N_39737);
or U39772 (N_39772,N_39575,N_39647);
and U39773 (N_39773,N_39502,N_39540);
xor U39774 (N_39774,N_39683,N_39722);
nor U39775 (N_39775,N_39732,N_39542);
xnor U39776 (N_39776,N_39671,N_39530);
xnor U39777 (N_39777,N_39503,N_39668);
nand U39778 (N_39778,N_39686,N_39519);
and U39779 (N_39779,N_39624,N_39693);
xor U39780 (N_39780,N_39508,N_39500);
or U39781 (N_39781,N_39667,N_39543);
xor U39782 (N_39782,N_39680,N_39602);
and U39783 (N_39783,N_39703,N_39720);
and U39784 (N_39784,N_39553,N_39535);
or U39785 (N_39785,N_39708,N_39595);
nand U39786 (N_39786,N_39700,N_39573);
nand U39787 (N_39787,N_39733,N_39544);
and U39788 (N_39788,N_39601,N_39550);
nand U39789 (N_39789,N_39587,N_39734);
nor U39790 (N_39790,N_39710,N_39622);
nor U39791 (N_39791,N_39603,N_39666);
nor U39792 (N_39792,N_39523,N_39674);
nand U39793 (N_39793,N_39657,N_39524);
xor U39794 (N_39794,N_39628,N_39736);
or U39795 (N_39795,N_39561,N_39504);
nand U39796 (N_39796,N_39537,N_39649);
or U39797 (N_39797,N_39568,N_39558);
xor U39798 (N_39798,N_39648,N_39682);
and U39799 (N_39799,N_39675,N_39556);
xnor U39800 (N_39800,N_39670,N_39527);
xnor U39801 (N_39801,N_39522,N_39650);
nor U39802 (N_39802,N_39633,N_39597);
or U39803 (N_39803,N_39744,N_39571);
or U39804 (N_39804,N_39745,N_39634);
and U39805 (N_39805,N_39726,N_39646);
nor U39806 (N_39806,N_39557,N_39607);
nor U39807 (N_39807,N_39521,N_39735);
nand U39808 (N_39808,N_39746,N_39645);
nor U39809 (N_39809,N_39518,N_39511);
and U39810 (N_39810,N_39565,N_39514);
xnor U39811 (N_39811,N_39531,N_39599);
or U39812 (N_39812,N_39606,N_39669);
xor U39813 (N_39813,N_39684,N_39663);
or U39814 (N_39814,N_39562,N_39642);
nand U39815 (N_39815,N_39694,N_39564);
xnor U39816 (N_39816,N_39516,N_39638);
and U39817 (N_39817,N_39594,N_39525);
nor U39818 (N_39818,N_39563,N_39574);
or U39819 (N_39819,N_39729,N_39555);
and U39820 (N_39820,N_39712,N_39731);
and U39821 (N_39821,N_39610,N_39545);
nand U39822 (N_39822,N_39538,N_39692);
or U39823 (N_39823,N_39551,N_39704);
nor U39824 (N_39824,N_39660,N_39630);
or U39825 (N_39825,N_39631,N_39590);
nand U39826 (N_39826,N_39534,N_39554);
and U39827 (N_39827,N_39566,N_39512);
xor U39828 (N_39828,N_39696,N_39591);
nor U39829 (N_39829,N_39596,N_39629);
or U39830 (N_39830,N_39613,N_39513);
nor U39831 (N_39831,N_39559,N_39721);
or U39832 (N_39832,N_39641,N_39536);
and U39833 (N_39833,N_39583,N_39640);
nand U39834 (N_39834,N_39685,N_39617);
xnor U39835 (N_39835,N_39738,N_39698);
or U39836 (N_39836,N_39576,N_39673);
nand U39837 (N_39837,N_39749,N_39526);
xor U39838 (N_39838,N_39584,N_39585);
nand U39839 (N_39839,N_39598,N_39515);
xnor U39840 (N_39840,N_39747,N_39653);
xnor U39841 (N_39841,N_39579,N_39517);
nand U39842 (N_39842,N_39739,N_39743);
nor U39843 (N_39843,N_39567,N_39505);
nor U39844 (N_39844,N_39740,N_39679);
nand U39845 (N_39845,N_39510,N_39533);
nand U39846 (N_39846,N_39618,N_39621);
nand U39847 (N_39847,N_39688,N_39541);
xor U39848 (N_39848,N_39681,N_39580);
nand U39849 (N_39849,N_39644,N_39637);
or U39850 (N_39850,N_39723,N_39701);
and U39851 (N_39851,N_39549,N_39592);
nor U39852 (N_39852,N_39509,N_39713);
xor U39853 (N_39853,N_39659,N_39715);
or U39854 (N_39854,N_39643,N_39691);
nand U39855 (N_39855,N_39547,N_39687);
and U39856 (N_39856,N_39724,N_39600);
xor U39857 (N_39857,N_39548,N_39593);
nor U39858 (N_39858,N_39725,N_39709);
xnor U39859 (N_39859,N_39609,N_39728);
nand U39860 (N_39860,N_39652,N_39627);
nor U39861 (N_39861,N_39608,N_39678);
and U39862 (N_39862,N_39635,N_39578);
or U39863 (N_39863,N_39676,N_39605);
and U39864 (N_39864,N_39742,N_39654);
nor U39865 (N_39865,N_39572,N_39717);
nand U39866 (N_39866,N_39616,N_39623);
nor U39867 (N_39867,N_39625,N_39611);
and U39868 (N_39868,N_39552,N_39532);
nand U39869 (N_39869,N_39620,N_39707);
nand U39870 (N_39870,N_39604,N_39718);
and U39871 (N_39871,N_39730,N_39689);
and U39872 (N_39872,N_39577,N_39716);
nand U39873 (N_39873,N_39636,N_39661);
or U39874 (N_39874,N_39677,N_39581);
nor U39875 (N_39875,N_39721,N_39684);
nor U39876 (N_39876,N_39575,N_39715);
nor U39877 (N_39877,N_39599,N_39592);
nand U39878 (N_39878,N_39538,N_39702);
and U39879 (N_39879,N_39534,N_39709);
nor U39880 (N_39880,N_39518,N_39679);
xnor U39881 (N_39881,N_39677,N_39630);
and U39882 (N_39882,N_39600,N_39635);
xnor U39883 (N_39883,N_39711,N_39685);
and U39884 (N_39884,N_39615,N_39718);
nor U39885 (N_39885,N_39520,N_39542);
nor U39886 (N_39886,N_39576,N_39718);
and U39887 (N_39887,N_39742,N_39595);
and U39888 (N_39888,N_39616,N_39501);
or U39889 (N_39889,N_39565,N_39551);
or U39890 (N_39890,N_39501,N_39732);
or U39891 (N_39891,N_39543,N_39723);
xor U39892 (N_39892,N_39729,N_39575);
nor U39893 (N_39893,N_39554,N_39612);
nor U39894 (N_39894,N_39570,N_39624);
nand U39895 (N_39895,N_39578,N_39732);
nand U39896 (N_39896,N_39701,N_39717);
xor U39897 (N_39897,N_39666,N_39667);
or U39898 (N_39898,N_39550,N_39698);
and U39899 (N_39899,N_39505,N_39564);
xor U39900 (N_39900,N_39534,N_39741);
or U39901 (N_39901,N_39661,N_39545);
or U39902 (N_39902,N_39688,N_39690);
nand U39903 (N_39903,N_39672,N_39611);
and U39904 (N_39904,N_39668,N_39607);
or U39905 (N_39905,N_39581,N_39515);
xor U39906 (N_39906,N_39669,N_39683);
nor U39907 (N_39907,N_39711,N_39702);
nand U39908 (N_39908,N_39510,N_39684);
nor U39909 (N_39909,N_39507,N_39594);
nor U39910 (N_39910,N_39652,N_39700);
and U39911 (N_39911,N_39651,N_39640);
or U39912 (N_39912,N_39697,N_39694);
nor U39913 (N_39913,N_39550,N_39611);
xnor U39914 (N_39914,N_39537,N_39734);
and U39915 (N_39915,N_39520,N_39721);
or U39916 (N_39916,N_39522,N_39520);
xor U39917 (N_39917,N_39608,N_39668);
nand U39918 (N_39918,N_39672,N_39673);
nor U39919 (N_39919,N_39642,N_39609);
xor U39920 (N_39920,N_39524,N_39527);
xor U39921 (N_39921,N_39534,N_39525);
nor U39922 (N_39922,N_39630,N_39634);
nand U39923 (N_39923,N_39633,N_39550);
nor U39924 (N_39924,N_39510,N_39695);
or U39925 (N_39925,N_39611,N_39716);
or U39926 (N_39926,N_39744,N_39632);
xnor U39927 (N_39927,N_39725,N_39572);
nor U39928 (N_39928,N_39596,N_39597);
or U39929 (N_39929,N_39638,N_39644);
xnor U39930 (N_39930,N_39523,N_39508);
xnor U39931 (N_39931,N_39666,N_39514);
xor U39932 (N_39932,N_39663,N_39555);
nand U39933 (N_39933,N_39503,N_39549);
nand U39934 (N_39934,N_39572,N_39618);
or U39935 (N_39935,N_39620,N_39577);
xnor U39936 (N_39936,N_39675,N_39513);
and U39937 (N_39937,N_39676,N_39517);
or U39938 (N_39938,N_39598,N_39562);
xor U39939 (N_39939,N_39579,N_39582);
or U39940 (N_39940,N_39577,N_39695);
and U39941 (N_39941,N_39686,N_39730);
and U39942 (N_39942,N_39526,N_39657);
or U39943 (N_39943,N_39694,N_39719);
or U39944 (N_39944,N_39633,N_39501);
xor U39945 (N_39945,N_39595,N_39625);
nand U39946 (N_39946,N_39675,N_39555);
nand U39947 (N_39947,N_39648,N_39502);
nand U39948 (N_39948,N_39581,N_39725);
nor U39949 (N_39949,N_39615,N_39591);
xor U39950 (N_39950,N_39670,N_39723);
or U39951 (N_39951,N_39615,N_39629);
and U39952 (N_39952,N_39735,N_39713);
nand U39953 (N_39953,N_39567,N_39586);
nand U39954 (N_39954,N_39643,N_39662);
or U39955 (N_39955,N_39611,N_39577);
or U39956 (N_39956,N_39631,N_39550);
xnor U39957 (N_39957,N_39561,N_39729);
and U39958 (N_39958,N_39664,N_39737);
and U39959 (N_39959,N_39746,N_39709);
xor U39960 (N_39960,N_39522,N_39577);
xnor U39961 (N_39961,N_39657,N_39712);
nand U39962 (N_39962,N_39654,N_39658);
xor U39963 (N_39963,N_39637,N_39638);
nor U39964 (N_39964,N_39706,N_39574);
xnor U39965 (N_39965,N_39716,N_39672);
xnor U39966 (N_39966,N_39748,N_39709);
nor U39967 (N_39967,N_39518,N_39646);
and U39968 (N_39968,N_39625,N_39521);
nor U39969 (N_39969,N_39535,N_39546);
and U39970 (N_39970,N_39553,N_39691);
nand U39971 (N_39971,N_39648,N_39675);
and U39972 (N_39972,N_39556,N_39507);
nor U39973 (N_39973,N_39669,N_39672);
or U39974 (N_39974,N_39559,N_39664);
nor U39975 (N_39975,N_39608,N_39692);
or U39976 (N_39976,N_39723,N_39544);
nor U39977 (N_39977,N_39505,N_39634);
or U39978 (N_39978,N_39681,N_39704);
nand U39979 (N_39979,N_39701,N_39524);
nor U39980 (N_39980,N_39712,N_39662);
and U39981 (N_39981,N_39726,N_39593);
xnor U39982 (N_39982,N_39589,N_39571);
or U39983 (N_39983,N_39623,N_39531);
nor U39984 (N_39984,N_39645,N_39657);
or U39985 (N_39985,N_39595,N_39588);
and U39986 (N_39986,N_39666,N_39520);
nor U39987 (N_39987,N_39540,N_39713);
or U39988 (N_39988,N_39674,N_39551);
nand U39989 (N_39989,N_39674,N_39552);
nor U39990 (N_39990,N_39699,N_39722);
nor U39991 (N_39991,N_39631,N_39739);
xnor U39992 (N_39992,N_39549,N_39609);
xnor U39993 (N_39993,N_39526,N_39588);
nand U39994 (N_39994,N_39611,N_39569);
or U39995 (N_39995,N_39727,N_39569);
xnor U39996 (N_39996,N_39726,N_39627);
and U39997 (N_39997,N_39555,N_39652);
or U39998 (N_39998,N_39635,N_39516);
nand U39999 (N_39999,N_39579,N_39599);
nor U40000 (N_40000,N_39779,N_39781);
nand U40001 (N_40001,N_39849,N_39761);
and U40002 (N_40002,N_39825,N_39858);
nand U40003 (N_40003,N_39965,N_39992);
nand U40004 (N_40004,N_39802,N_39799);
and U40005 (N_40005,N_39998,N_39944);
and U40006 (N_40006,N_39787,N_39908);
and U40007 (N_40007,N_39986,N_39844);
nand U40008 (N_40008,N_39981,N_39996);
or U40009 (N_40009,N_39789,N_39791);
or U40010 (N_40010,N_39859,N_39780);
nor U40011 (N_40011,N_39970,N_39873);
xnor U40012 (N_40012,N_39978,N_39918);
nor U40013 (N_40013,N_39882,N_39903);
and U40014 (N_40014,N_39966,N_39980);
nand U40015 (N_40015,N_39968,N_39931);
nor U40016 (N_40016,N_39962,N_39995);
or U40017 (N_40017,N_39861,N_39866);
nand U40018 (N_40018,N_39775,N_39753);
or U40019 (N_40019,N_39940,N_39893);
nor U40020 (N_40020,N_39786,N_39875);
nor U40021 (N_40021,N_39897,N_39846);
nand U40022 (N_40022,N_39900,N_39892);
or U40023 (N_40023,N_39899,N_39788);
xnor U40024 (N_40024,N_39776,N_39993);
or U40025 (N_40025,N_39987,N_39848);
and U40026 (N_40026,N_39991,N_39759);
xnor U40027 (N_40027,N_39774,N_39826);
xnor U40028 (N_40028,N_39919,N_39763);
nand U40029 (N_40029,N_39878,N_39990);
or U40030 (N_40030,N_39905,N_39855);
nor U40031 (N_40031,N_39804,N_39762);
and U40032 (N_40032,N_39907,N_39796);
xor U40033 (N_40033,N_39988,N_39949);
xnor U40034 (N_40034,N_39979,N_39842);
nor U40035 (N_40035,N_39816,N_39857);
or U40036 (N_40036,N_39808,N_39831);
and U40037 (N_40037,N_39853,N_39818);
and U40038 (N_40038,N_39932,N_39889);
or U40039 (N_40039,N_39872,N_39963);
nand U40040 (N_40040,N_39792,N_39782);
xnor U40041 (N_40041,N_39894,N_39766);
and U40042 (N_40042,N_39954,N_39790);
or U40043 (N_40043,N_39922,N_39967);
nand U40044 (N_40044,N_39868,N_39943);
nor U40045 (N_40045,N_39915,N_39793);
xnor U40046 (N_40046,N_39864,N_39794);
nor U40047 (N_40047,N_39914,N_39895);
xor U40048 (N_40048,N_39834,N_39929);
xor U40049 (N_40049,N_39783,N_39916);
and U40050 (N_40050,N_39771,N_39810);
nand U40051 (N_40051,N_39896,N_39974);
and U40052 (N_40052,N_39960,N_39921);
and U40053 (N_40053,N_39942,N_39876);
nor U40054 (N_40054,N_39815,N_39933);
xnor U40055 (N_40055,N_39912,N_39837);
xor U40056 (N_40056,N_39983,N_39860);
nor U40057 (N_40057,N_39890,N_39851);
xnor U40058 (N_40058,N_39898,N_39755);
nand U40059 (N_40059,N_39977,N_39959);
nor U40060 (N_40060,N_39823,N_39847);
or U40061 (N_40061,N_39767,N_39854);
or U40062 (N_40062,N_39784,N_39862);
xnor U40063 (N_40063,N_39845,N_39817);
xor U40064 (N_40064,N_39874,N_39886);
nor U40065 (N_40065,N_39999,N_39982);
nand U40066 (N_40066,N_39984,N_39956);
xnor U40067 (N_40067,N_39805,N_39813);
or U40068 (N_40068,N_39777,N_39917);
or U40069 (N_40069,N_39936,N_39927);
nand U40070 (N_40070,N_39971,N_39839);
xnor U40071 (N_40071,N_39773,N_39928);
xnor U40072 (N_40072,N_39946,N_39833);
nand U40073 (N_40073,N_39871,N_39885);
and U40074 (N_40074,N_39953,N_39961);
xor U40075 (N_40075,N_39772,N_39865);
nand U40076 (N_40076,N_39923,N_39948);
nand U40077 (N_40077,N_39884,N_39795);
and U40078 (N_40078,N_39934,N_39830);
nor U40079 (N_40079,N_39840,N_39750);
or U40080 (N_40080,N_39972,N_39930);
or U40081 (N_40081,N_39957,N_39754);
or U40082 (N_40082,N_39945,N_39877);
or U40083 (N_40083,N_39939,N_39973);
and U40084 (N_40084,N_39937,N_39778);
and U40085 (N_40085,N_39798,N_39887);
xnor U40086 (N_40086,N_39801,N_39751);
nor U40087 (N_40087,N_39950,N_39926);
and U40088 (N_40088,N_39891,N_39832);
nor U40089 (N_40089,N_39768,N_39809);
nand U40090 (N_40090,N_39770,N_39800);
and U40091 (N_40091,N_39901,N_39824);
or U40092 (N_40092,N_39975,N_39947);
xor U40093 (N_40093,N_39850,N_39821);
and U40094 (N_40094,N_39812,N_39820);
xor U40095 (N_40095,N_39969,N_39976);
or U40096 (N_40096,N_39881,N_39752);
nor U40097 (N_40097,N_39964,N_39841);
and U40098 (N_40098,N_39951,N_39836);
nor U40099 (N_40099,N_39869,N_39806);
xor U40100 (N_40100,N_39909,N_39814);
xor U40101 (N_40101,N_39924,N_39910);
nand U40102 (N_40102,N_39765,N_39769);
xnor U40103 (N_40103,N_39838,N_39867);
and U40104 (N_40104,N_39756,N_39938);
nor U40105 (N_40105,N_39785,N_39920);
nor U40106 (N_40106,N_39803,N_39902);
xor U40107 (N_40107,N_39941,N_39994);
nand U40108 (N_40108,N_39958,N_39883);
nand U40109 (N_40109,N_39811,N_39906);
or U40110 (N_40110,N_39925,N_39955);
nand U40111 (N_40111,N_39997,N_39829);
nor U40112 (N_40112,N_39760,N_39807);
xor U40113 (N_40113,N_39880,N_39911);
nor U40114 (N_40114,N_39935,N_39952);
xor U40115 (N_40115,N_39822,N_39904);
and U40116 (N_40116,N_39852,N_39757);
nor U40117 (N_40117,N_39863,N_39985);
xor U40118 (N_40118,N_39856,N_39828);
or U40119 (N_40119,N_39913,N_39989);
and U40120 (N_40120,N_39827,N_39819);
nand U40121 (N_40121,N_39758,N_39888);
and U40122 (N_40122,N_39843,N_39870);
and U40123 (N_40123,N_39879,N_39835);
nand U40124 (N_40124,N_39797,N_39764);
nand U40125 (N_40125,N_39955,N_39900);
nand U40126 (N_40126,N_39812,N_39912);
or U40127 (N_40127,N_39997,N_39937);
nand U40128 (N_40128,N_39856,N_39958);
nor U40129 (N_40129,N_39840,N_39909);
nand U40130 (N_40130,N_39763,N_39994);
xor U40131 (N_40131,N_39983,N_39871);
nand U40132 (N_40132,N_39811,N_39938);
and U40133 (N_40133,N_39861,N_39966);
nor U40134 (N_40134,N_39913,N_39947);
nor U40135 (N_40135,N_39988,N_39816);
nand U40136 (N_40136,N_39947,N_39860);
nor U40137 (N_40137,N_39769,N_39891);
nand U40138 (N_40138,N_39794,N_39809);
and U40139 (N_40139,N_39851,N_39934);
nand U40140 (N_40140,N_39974,N_39805);
and U40141 (N_40141,N_39919,N_39940);
nor U40142 (N_40142,N_39938,N_39851);
xor U40143 (N_40143,N_39803,N_39975);
or U40144 (N_40144,N_39864,N_39913);
or U40145 (N_40145,N_39994,N_39785);
or U40146 (N_40146,N_39845,N_39814);
nand U40147 (N_40147,N_39867,N_39765);
or U40148 (N_40148,N_39828,N_39957);
xnor U40149 (N_40149,N_39983,N_39876);
and U40150 (N_40150,N_39878,N_39788);
nor U40151 (N_40151,N_39950,N_39887);
nor U40152 (N_40152,N_39963,N_39780);
or U40153 (N_40153,N_39965,N_39915);
nor U40154 (N_40154,N_39934,N_39869);
or U40155 (N_40155,N_39992,N_39926);
nand U40156 (N_40156,N_39810,N_39929);
nand U40157 (N_40157,N_39803,N_39766);
nor U40158 (N_40158,N_39866,N_39841);
nand U40159 (N_40159,N_39999,N_39768);
nand U40160 (N_40160,N_39767,N_39971);
nand U40161 (N_40161,N_39936,N_39987);
nor U40162 (N_40162,N_39771,N_39984);
or U40163 (N_40163,N_39875,N_39908);
or U40164 (N_40164,N_39931,N_39944);
or U40165 (N_40165,N_39883,N_39869);
nor U40166 (N_40166,N_39923,N_39757);
xor U40167 (N_40167,N_39808,N_39850);
and U40168 (N_40168,N_39823,N_39947);
nand U40169 (N_40169,N_39915,N_39918);
and U40170 (N_40170,N_39809,N_39822);
and U40171 (N_40171,N_39795,N_39842);
nand U40172 (N_40172,N_39754,N_39770);
nand U40173 (N_40173,N_39971,N_39858);
nand U40174 (N_40174,N_39972,N_39860);
xor U40175 (N_40175,N_39971,N_39788);
and U40176 (N_40176,N_39779,N_39955);
and U40177 (N_40177,N_39832,N_39870);
xnor U40178 (N_40178,N_39936,N_39966);
xor U40179 (N_40179,N_39814,N_39816);
nor U40180 (N_40180,N_39841,N_39991);
and U40181 (N_40181,N_39855,N_39965);
nand U40182 (N_40182,N_39845,N_39904);
or U40183 (N_40183,N_39987,N_39998);
or U40184 (N_40184,N_39927,N_39980);
xor U40185 (N_40185,N_39942,N_39891);
xnor U40186 (N_40186,N_39992,N_39838);
and U40187 (N_40187,N_39889,N_39840);
and U40188 (N_40188,N_39884,N_39921);
xnor U40189 (N_40189,N_39991,N_39780);
nand U40190 (N_40190,N_39815,N_39897);
xnor U40191 (N_40191,N_39794,N_39957);
xnor U40192 (N_40192,N_39866,N_39830);
xnor U40193 (N_40193,N_39926,N_39868);
or U40194 (N_40194,N_39806,N_39917);
nand U40195 (N_40195,N_39782,N_39866);
xnor U40196 (N_40196,N_39994,N_39916);
and U40197 (N_40197,N_39963,N_39806);
and U40198 (N_40198,N_39852,N_39955);
nand U40199 (N_40199,N_39858,N_39760);
nor U40200 (N_40200,N_39754,N_39904);
nor U40201 (N_40201,N_39922,N_39970);
and U40202 (N_40202,N_39799,N_39841);
and U40203 (N_40203,N_39818,N_39823);
or U40204 (N_40204,N_39840,N_39846);
or U40205 (N_40205,N_39941,N_39999);
xnor U40206 (N_40206,N_39825,N_39874);
or U40207 (N_40207,N_39831,N_39833);
nand U40208 (N_40208,N_39938,N_39848);
nor U40209 (N_40209,N_39951,N_39949);
nor U40210 (N_40210,N_39782,N_39835);
nor U40211 (N_40211,N_39820,N_39904);
and U40212 (N_40212,N_39872,N_39884);
and U40213 (N_40213,N_39819,N_39756);
and U40214 (N_40214,N_39897,N_39997);
xnor U40215 (N_40215,N_39965,N_39849);
xnor U40216 (N_40216,N_39814,N_39782);
nand U40217 (N_40217,N_39846,N_39945);
and U40218 (N_40218,N_39789,N_39861);
nand U40219 (N_40219,N_39947,N_39848);
nor U40220 (N_40220,N_39894,N_39777);
nand U40221 (N_40221,N_39924,N_39992);
or U40222 (N_40222,N_39901,N_39911);
xor U40223 (N_40223,N_39814,N_39801);
xnor U40224 (N_40224,N_39850,N_39865);
xnor U40225 (N_40225,N_39752,N_39829);
xor U40226 (N_40226,N_39833,N_39765);
nand U40227 (N_40227,N_39785,N_39765);
nor U40228 (N_40228,N_39765,N_39775);
nor U40229 (N_40229,N_39785,N_39795);
and U40230 (N_40230,N_39941,N_39789);
nor U40231 (N_40231,N_39826,N_39874);
xnor U40232 (N_40232,N_39780,N_39966);
nor U40233 (N_40233,N_39904,N_39979);
or U40234 (N_40234,N_39770,N_39784);
nor U40235 (N_40235,N_39956,N_39967);
xor U40236 (N_40236,N_39963,N_39815);
or U40237 (N_40237,N_39761,N_39935);
xnor U40238 (N_40238,N_39757,N_39969);
and U40239 (N_40239,N_39958,N_39779);
and U40240 (N_40240,N_39863,N_39975);
nor U40241 (N_40241,N_39982,N_39764);
or U40242 (N_40242,N_39998,N_39929);
xnor U40243 (N_40243,N_39949,N_39850);
and U40244 (N_40244,N_39942,N_39934);
nand U40245 (N_40245,N_39848,N_39992);
or U40246 (N_40246,N_39822,N_39761);
nand U40247 (N_40247,N_39761,N_39916);
nand U40248 (N_40248,N_39937,N_39859);
or U40249 (N_40249,N_39887,N_39767);
xnor U40250 (N_40250,N_40141,N_40120);
nand U40251 (N_40251,N_40110,N_40198);
and U40252 (N_40252,N_40187,N_40008);
nand U40253 (N_40253,N_40226,N_40124);
xnor U40254 (N_40254,N_40025,N_40174);
and U40255 (N_40255,N_40106,N_40007);
or U40256 (N_40256,N_40131,N_40233);
xor U40257 (N_40257,N_40005,N_40099);
nand U40258 (N_40258,N_40149,N_40011);
and U40259 (N_40259,N_40199,N_40053);
xnor U40260 (N_40260,N_40191,N_40098);
and U40261 (N_40261,N_40249,N_40242);
or U40262 (N_40262,N_40138,N_40221);
nand U40263 (N_40263,N_40091,N_40048);
and U40264 (N_40264,N_40216,N_40064);
nand U40265 (N_40265,N_40234,N_40229);
nand U40266 (N_40266,N_40070,N_40113);
and U40267 (N_40267,N_40243,N_40219);
nor U40268 (N_40268,N_40209,N_40122);
and U40269 (N_40269,N_40139,N_40118);
nand U40270 (N_40270,N_40235,N_40123);
and U40271 (N_40271,N_40157,N_40046);
xnor U40272 (N_40272,N_40237,N_40060);
and U40273 (N_40273,N_40093,N_40215);
nand U40274 (N_40274,N_40051,N_40127);
xor U40275 (N_40275,N_40115,N_40054);
or U40276 (N_40276,N_40193,N_40023);
nand U40277 (N_40277,N_40100,N_40044);
and U40278 (N_40278,N_40232,N_40004);
nand U40279 (N_40279,N_40196,N_40129);
nor U40280 (N_40280,N_40164,N_40205);
or U40281 (N_40281,N_40244,N_40069);
nor U40282 (N_40282,N_40200,N_40150);
nor U40283 (N_40283,N_40214,N_40081);
xor U40284 (N_40284,N_40059,N_40201);
nand U40285 (N_40285,N_40155,N_40089);
xor U40286 (N_40286,N_40076,N_40034);
nand U40287 (N_40287,N_40121,N_40086);
xnor U40288 (N_40288,N_40169,N_40063);
and U40289 (N_40289,N_40105,N_40185);
nand U40290 (N_40290,N_40208,N_40194);
xnor U40291 (N_40291,N_40217,N_40080);
xor U40292 (N_40292,N_40119,N_40167);
nor U40293 (N_40293,N_40236,N_40238);
nor U40294 (N_40294,N_40022,N_40017);
xor U40295 (N_40295,N_40135,N_40027);
and U40296 (N_40296,N_40188,N_40090);
nor U40297 (N_40297,N_40075,N_40225);
xor U40298 (N_40298,N_40112,N_40246);
and U40299 (N_40299,N_40016,N_40108);
and U40300 (N_40300,N_40001,N_40071);
xnor U40301 (N_40301,N_40211,N_40000);
nand U40302 (N_40302,N_40049,N_40074);
and U40303 (N_40303,N_40083,N_40009);
nor U40304 (N_40304,N_40125,N_40134);
nor U40305 (N_40305,N_40220,N_40186);
xnor U40306 (N_40306,N_40026,N_40223);
and U40307 (N_40307,N_40144,N_40172);
or U40308 (N_40308,N_40158,N_40183);
nor U40309 (N_40309,N_40203,N_40132);
nor U40310 (N_40310,N_40168,N_40133);
and U40311 (N_40311,N_40057,N_40037);
or U40312 (N_40312,N_40088,N_40042);
nand U40313 (N_40313,N_40154,N_40212);
xor U40314 (N_40314,N_40045,N_40239);
nor U40315 (N_40315,N_40160,N_40152);
nor U40316 (N_40316,N_40204,N_40095);
or U40317 (N_40317,N_40024,N_40068);
and U40318 (N_40318,N_40210,N_40010);
nor U40319 (N_40319,N_40029,N_40111);
nor U40320 (N_40320,N_40035,N_40202);
nor U40321 (N_40321,N_40116,N_40228);
xnor U40322 (N_40322,N_40230,N_40153);
nor U40323 (N_40323,N_40006,N_40078);
or U40324 (N_40324,N_40248,N_40207);
nand U40325 (N_40325,N_40173,N_40061);
and U40326 (N_40326,N_40107,N_40165);
nand U40327 (N_40327,N_40197,N_40030);
nor U40328 (N_40328,N_40047,N_40028);
and U40329 (N_40329,N_40072,N_40085);
xor U40330 (N_40330,N_40033,N_40103);
or U40331 (N_40331,N_40014,N_40140);
nand U40332 (N_40332,N_40087,N_40148);
xnor U40333 (N_40333,N_40181,N_40180);
xor U40334 (N_40334,N_40218,N_40021);
nor U40335 (N_40335,N_40067,N_40245);
xor U40336 (N_40336,N_40012,N_40136);
xor U40337 (N_40337,N_40247,N_40036);
and U40338 (N_40338,N_40020,N_40241);
and U40339 (N_40339,N_40032,N_40097);
or U40340 (N_40340,N_40192,N_40104);
xnor U40341 (N_40341,N_40195,N_40224);
nor U40342 (N_40342,N_40018,N_40092);
nand U40343 (N_40343,N_40213,N_40130);
xor U40344 (N_40344,N_40050,N_40142);
xor U40345 (N_40345,N_40062,N_40058);
or U40346 (N_40346,N_40137,N_40073);
xor U40347 (N_40347,N_40177,N_40052);
nand U40348 (N_40348,N_40231,N_40184);
xor U40349 (N_40349,N_40102,N_40189);
nor U40350 (N_40350,N_40182,N_40043);
xor U40351 (N_40351,N_40151,N_40179);
or U40352 (N_40352,N_40019,N_40190);
xor U40353 (N_40353,N_40162,N_40222);
and U40354 (N_40354,N_40206,N_40175);
and U40355 (N_40355,N_40147,N_40040);
nand U40356 (N_40356,N_40171,N_40163);
and U40357 (N_40357,N_40159,N_40146);
and U40358 (N_40358,N_40143,N_40082);
xor U40359 (N_40359,N_40056,N_40161);
or U40360 (N_40360,N_40039,N_40077);
nand U40361 (N_40361,N_40114,N_40079);
xnor U40362 (N_40362,N_40166,N_40227);
nand U40363 (N_40363,N_40128,N_40065);
nor U40364 (N_40364,N_40084,N_40126);
nor U40365 (N_40365,N_40055,N_40240);
or U40366 (N_40366,N_40178,N_40145);
nor U40367 (N_40367,N_40170,N_40003);
nand U40368 (N_40368,N_40002,N_40013);
or U40369 (N_40369,N_40096,N_40031);
nor U40370 (N_40370,N_40101,N_40094);
xor U40371 (N_40371,N_40041,N_40109);
or U40372 (N_40372,N_40015,N_40117);
or U40373 (N_40373,N_40066,N_40156);
nor U40374 (N_40374,N_40176,N_40038);
xor U40375 (N_40375,N_40196,N_40020);
and U40376 (N_40376,N_40004,N_40036);
nand U40377 (N_40377,N_40127,N_40214);
xnor U40378 (N_40378,N_40060,N_40138);
xnor U40379 (N_40379,N_40123,N_40013);
xnor U40380 (N_40380,N_40141,N_40148);
or U40381 (N_40381,N_40237,N_40139);
nor U40382 (N_40382,N_40205,N_40172);
or U40383 (N_40383,N_40157,N_40211);
nor U40384 (N_40384,N_40068,N_40103);
nor U40385 (N_40385,N_40180,N_40067);
nor U40386 (N_40386,N_40215,N_40131);
nor U40387 (N_40387,N_40029,N_40172);
and U40388 (N_40388,N_40229,N_40197);
xnor U40389 (N_40389,N_40000,N_40054);
nor U40390 (N_40390,N_40054,N_40155);
and U40391 (N_40391,N_40213,N_40030);
and U40392 (N_40392,N_40027,N_40051);
and U40393 (N_40393,N_40194,N_40209);
nand U40394 (N_40394,N_40039,N_40075);
xnor U40395 (N_40395,N_40030,N_40014);
or U40396 (N_40396,N_40223,N_40139);
and U40397 (N_40397,N_40051,N_40157);
nand U40398 (N_40398,N_40033,N_40097);
nand U40399 (N_40399,N_40212,N_40070);
nor U40400 (N_40400,N_40163,N_40146);
xnor U40401 (N_40401,N_40124,N_40145);
nor U40402 (N_40402,N_40174,N_40207);
or U40403 (N_40403,N_40125,N_40127);
and U40404 (N_40404,N_40162,N_40197);
and U40405 (N_40405,N_40128,N_40091);
xor U40406 (N_40406,N_40193,N_40033);
nand U40407 (N_40407,N_40190,N_40126);
nand U40408 (N_40408,N_40033,N_40073);
xnor U40409 (N_40409,N_40047,N_40192);
or U40410 (N_40410,N_40083,N_40230);
or U40411 (N_40411,N_40156,N_40018);
or U40412 (N_40412,N_40126,N_40146);
nand U40413 (N_40413,N_40153,N_40125);
nor U40414 (N_40414,N_40024,N_40011);
and U40415 (N_40415,N_40051,N_40220);
and U40416 (N_40416,N_40122,N_40212);
nand U40417 (N_40417,N_40102,N_40151);
nand U40418 (N_40418,N_40060,N_40211);
nand U40419 (N_40419,N_40097,N_40003);
nand U40420 (N_40420,N_40109,N_40180);
and U40421 (N_40421,N_40223,N_40215);
xnor U40422 (N_40422,N_40133,N_40197);
and U40423 (N_40423,N_40102,N_40178);
nand U40424 (N_40424,N_40229,N_40168);
or U40425 (N_40425,N_40014,N_40114);
nand U40426 (N_40426,N_40154,N_40130);
xnor U40427 (N_40427,N_40091,N_40163);
xor U40428 (N_40428,N_40101,N_40124);
or U40429 (N_40429,N_40207,N_40106);
or U40430 (N_40430,N_40164,N_40096);
nor U40431 (N_40431,N_40004,N_40026);
nor U40432 (N_40432,N_40155,N_40226);
nor U40433 (N_40433,N_40065,N_40112);
and U40434 (N_40434,N_40152,N_40015);
nand U40435 (N_40435,N_40153,N_40236);
or U40436 (N_40436,N_40050,N_40155);
nor U40437 (N_40437,N_40093,N_40003);
nor U40438 (N_40438,N_40040,N_40187);
xor U40439 (N_40439,N_40169,N_40203);
and U40440 (N_40440,N_40071,N_40201);
or U40441 (N_40441,N_40151,N_40046);
or U40442 (N_40442,N_40037,N_40239);
nor U40443 (N_40443,N_40154,N_40238);
xnor U40444 (N_40444,N_40027,N_40160);
nand U40445 (N_40445,N_40102,N_40065);
nor U40446 (N_40446,N_40087,N_40071);
and U40447 (N_40447,N_40179,N_40118);
nand U40448 (N_40448,N_40173,N_40214);
nor U40449 (N_40449,N_40096,N_40241);
and U40450 (N_40450,N_40086,N_40085);
or U40451 (N_40451,N_40054,N_40006);
xnor U40452 (N_40452,N_40152,N_40112);
nor U40453 (N_40453,N_40176,N_40228);
xnor U40454 (N_40454,N_40172,N_40120);
or U40455 (N_40455,N_40021,N_40145);
xnor U40456 (N_40456,N_40074,N_40220);
and U40457 (N_40457,N_40214,N_40130);
nand U40458 (N_40458,N_40182,N_40088);
nor U40459 (N_40459,N_40211,N_40071);
or U40460 (N_40460,N_40122,N_40196);
or U40461 (N_40461,N_40070,N_40086);
nand U40462 (N_40462,N_40186,N_40069);
and U40463 (N_40463,N_40173,N_40086);
or U40464 (N_40464,N_40162,N_40004);
or U40465 (N_40465,N_40008,N_40083);
and U40466 (N_40466,N_40171,N_40109);
xor U40467 (N_40467,N_40183,N_40074);
or U40468 (N_40468,N_40071,N_40059);
nor U40469 (N_40469,N_40229,N_40057);
and U40470 (N_40470,N_40243,N_40121);
and U40471 (N_40471,N_40026,N_40167);
nor U40472 (N_40472,N_40069,N_40010);
nand U40473 (N_40473,N_40029,N_40155);
nor U40474 (N_40474,N_40201,N_40118);
or U40475 (N_40475,N_40062,N_40123);
nor U40476 (N_40476,N_40199,N_40128);
xor U40477 (N_40477,N_40028,N_40072);
or U40478 (N_40478,N_40164,N_40054);
nor U40479 (N_40479,N_40125,N_40244);
and U40480 (N_40480,N_40197,N_40092);
nand U40481 (N_40481,N_40126,N_40188);
nor U40482 (N_40482,N_40136,N_40111);
xor U40483 (N_40483,N_40163,N_40175);
xnor U40484 (N_40484,N_40193,N_40190);
xor U40485 (N_40485,N_40077,N_40204);
nor U40486 (N_40486,N_40232,N_40043);
xor U40487 (N_40487,N_40137,N_40055);
nor U40488 (N_40488,N_40187,N_40071);
nor U40489 (N_40489,N_40010,N_40156);
nand U40490 (N_40490,N_40102,N_40155);
and U40491 (N_40491,N_40204,N_40177);
nand U40492 (N_40492,N_40161,N_40093);
and U40493 (N_40493,N_40148,N_40012);
and U40494 (N_40494,N_40097,N_40012);
nor U40495 (N_40495,N_40147,N_40206);
nor U40496 (N_40496,N_40151,N_40028);
and U40497 (N_40497,N_40242,N_40152);
nand U40498 (N_40498,N_40051,N_40231);
and U40499 (N_40499,N_40122,N_40189);
nor U40500 (N_40500,N_40314,N_40302);
nor U40501 (N_40501,N_40455,N_40264);
nor U40502 (N_40502,N_40418,N_40442);
nor U40503 (N_40503,N_40454,N_40433);
nand U40504 (N_40504,N_40465,N_40321);
nand U40505 (N_40505,N_40335,N_40430);
xor U40506 (N_40506,N_40356,N_40364);
nand U40507 (N_40507,N_40397,N_40429);
xor U40508 (N_40508,N_40289,N_40480);
nand U40509 (N_40509,N_40460,N_40408);
nand U40510 (N_40510,N_40471,N_40479);
or U40511 (N_40511,N_40478,N_40263);
nor U40512 (N_40512,N_40270,N_40309);
xor U40513 (N_40513,N_40492,N_40295);
xor U40514 (N_40514,N_40457,N_40343);
or U40515 (N_40515,N_40276,N_40463);
xnor U40516 (N_40516,N_40300,N_40412);
or U40517 (N_40517,N_40252,N_40251);
or U40518 (N_40518,N_40388,N_40481);
or U40519 (N_40519,N_40358,N_40307);
nor U40520 (N_40520,N_40474,N_40334);
and U40521 (N_40521,N_40486,N_40436);
nor U40522 (N_40522,N_40407,N_40472);
or U40523 (N_40523,N_40395,N_40280);
xnor U40524 (N_40524,N_40294,N_40473);
and U40525 (N_40525,N_40271,N_40275);
xor U40526 (N_40526,N_40490,N_40337);
xor U40527 (N_40527,N_40318,N_40425);
or U40528 (N_40528,N_40260,N_40353);
or U40529 (N_40529,N_40399,N_40391);
xnor U40530 (N_40530,N_40361,N_40417);
xnor U40531 (N_40531,N_40308,N_40447);
or U40532 (N_40532,N_40250,N_40446);
and U40533 (N_40533,N_40404,N_40402);
xor U40534 (N_40534,N_40434,N_40498);
nand U40535 (N_40535,N_40393,N_40444);
or U40536 (N_40536,N_40369,N_40466);
xnor U40537 (N_40537,N_40383,N_40256);
or U40538 (N_40538,N_40326,N_40296);
and U40539 (N_40539,N_40368,N_40421);
nand U40540 (N_40540,N_40427,N_40371);
nand U40541 (N_40541,N_40488,N_40386);
nand U40542 (N_40542,N_40445,N_40384);
nand U40543 (N_40543,N_40424,N_40458);
nor U40544 (N_40544,N_40400,N_40456);
nor U40545 (N_40545,N_40338,N_40420);
xnor U40546 (N_40546,N_40363,N_40435);
or U40547 (N_40547,N_40449,N_40290);
nand U40548 (N_40548,N_40331,N_40370);
nand U40549 (N_40549,N_40484,N_40414);
nor U40550 (N_40550,N_40413,N_40333);
nand U40551 (N_40551,N_40374,N_40366);
xor U40552 (N_40552,N_40459,N_40299);
xor U40553 (N_40553,N_40379,N_40350);
nor U40554 (N_40554,N_40362,N_40467);
xnor U40555 (N_40555,N_40390,N_40483);
nand U40556 (N_40556,N_40428,N_40272);
and U40557 (N_40557,N_40329,N_40265);
xnor U40558 (N_40558,N_40262,N_40423);
nand U40559 (N_40559,N_40415,N_40469);
and U40560 (N_40560,N_40382,N_40322);
or U40561 (N_40561,N_40281,N_40312);
nor U40562 (N_40562,N_40259,N_40257);
or U40563 (N_40563,N_40401,N_40266);
xor U40564 (N_40564,N_40340,N_40394);
nand U40565 (N_40565,N_40405,N_40306);
or U40566 (N_40566,N_40261,N_40293);
and U40567 (N_40567,N_40448,N_40323);
nand U40568 (N_40568,N_40438,N_40348);
nand U40569 (N_40569,N_40499,N_40311);
xnor U40570 (N_40570,N_40468,N_40389);
and U40571 (N_40571,N_40310,N_40432);
nor U40572 (N_40572,N_40327,N_40411);
nor U40573 (N_40573,N_40269,N_40439);
xor U40574 (N_40574,N_40441,N_40258);
nand U40575 (N_40575,N_40431,N_40332);
xnor U40576 (N_40576,N_40470,N_40283);
nand U40577 (N_40577,N_40381,N_40419);
and U40578 (N_40578,N_40301,N_40375);
nor U40579 (N_40579,N_40319,N_40336);
nor U40580 (N_40580,N_40380,N_40349);
or U40581 (N_40581,N_40376,N_40313);
nor U40582 (N_40582,N_40396,N_40268);
and U40583 (N_40583,N_40273,N_40387);
or U40584 (N_40584,N_40378,N_40373);
nor U40585 (N_40585,N_40324,N_40475);
nor U40586 (N_40586,N_40328,N_40285);
nor U40587 (N_40587,N_40482,N_40354);
xnor U40588 (N_40588,N_40494,N_40493);
and U40589 (N_40589,N_40437,N_40476);
nand U40590 (N_40590,N_40351,N_40330);
xor U40591 (N_40591,N_40410,N_40360);
nand U40592 (N_40592,N_40355,N_40464);
xor U40593 (N_40593,N_40392,N_40403);
and U40594 (N_40594,N_40303,N_40477);
xnor U40595 (N_40595,N_40286,N_40291);
and U40596 (N_40596,N_40344,N_40320);
or U40597 (N_40597,N_40385,N_40496);
or U40598 (N_40598,N_40352,N_40282);
xor U40599 (N_40599,N_40288,N_40497);
xor U40600 (N_40600,N_40409,N_40347);
nor U40601 (N_40601,N_40297,N_40416);
or U40602 (N_40602,N_40377,N_40254);
or U40603 (N_40603,N_40359,N_40315);
and U40604 (N_40604,N_40489,N_40316);
nand U40605 (N_40605,N_40339,N_40287);
or U40606 (N_40606,N_40422,N_40365);
nor U40607 (N_40607,N_40267,N_40495);
nand U40608 (N_40608,N_40341,N_40345);
or U40609 (N_40609,N_40406,N_40279);
nor U40610 (N_40610,N_40255,N_40342);
nor U40611 (N_40611,N_40298,N_40372);
nand U40612 (N_40612,N_40277,N_40453);
xnor U40613 (N_40613,N_40253,N_40304);
xnor U40614 (N_40614,N_40440,N_40305);
xor U40615 (N_40615,N_40278,N_40461);
and U40616 (N_40616,N_40450,N_40346);
nor U40617 (N_40617,N_40274,N_40284);
or U40618 (N_40618,N_40317,N_40487);
nand U40619 (N_40619,N_40491,N_40426);
and U40620 (N_40620,N_40452,N_40325);
nor U40621 (N_40621,N_40367,N_40451);
and U40622 (N_40622,N_40443,N_40462);
xor U40623 (N_40623,N_40292,N_40398);
xor U40624 (N_40624,N_40357,N_40485);
xnor U40625 (N_40625,N_40331,N_40440);
xnor U40626 (N_40626,N_40469,N_40338);
nand U40627 (N_40627,N_40302,N_40347);
nor U40628 (N_40628,N_40268,N_40256);
and U40629 (N_40629,N_40327,N_40325);
xnor U40630 (N_40630,N_40329,N_40383);
and U40631 (N_40631,N_40434,N_40426);
nand U40632 (N_40632,N_40349,N_40278);
nand U40633 (N_40633,N_40416,N_40317);
and U40634 (N_40634,N_40270,N_40414);
nor U40635 (N_40635,N_40330,N_40410);
or U40636 (N_40636,N_40400,N_40330);
nor U40637 (N_40637,N_40286,N_40342);
xor U40638 (N_40638,N_40281,N_40374);
and U40639 (N_40639,N_40374,N_40357);
and U40640 (N_40640,N_40269,N_40270);
nor U40641 (N_40641,N_40252,N_40469);
xor U40642 (N_40642,N_40331,N_40488);
or U40643 (N_40643,N_40425,N_40384);
or U40644 (N_40644,N_40332,N_40358);
and U40645 (N_40645,N_40327,N_40380);
nand U40646 (N_40646,N_40380,N_40282);
and U40647 (N_40647,N_40472,N_40270);
nor U40648 (N_40648,N_40374,N_40439);
and U40649 (N_40649,N_40414,N_40471);
or U40650 (N_40650,N_40367,N_40481);
nand U40651 (N_40651,N_40306,N_40265);
nand U40652 (N_40652,N_40427,N_40497);
nand U40653 (N_40653,N_40477,N_40456);
or U40654 (N_40654,N_40310,N_40366);
nor U40655 (N_40655,N_40365,N_40317);
and U40656 (N_40656,N_40298,N_40392);
or U40657 (N_40657,N_40477,N_40399);
nor U40658 (N_40658,N_40446,N_40367);
or U40659 (N_40659,N_40270,N_40288);
nor U40660 (N_40660,N_40463,N_40486);
xor U40661 (N_40661,N_40329,N_40391);
nor U40662 (N_40662,N_40429,N_40435);
and U40663 (N_40663,N_40417,N_40360);
and U40664 (N_40664,N_40297,N_40401);
xnor U40665 (N_40665,N_40287,N_40389);
xnor U40666 (N_40666,N_40406,N_40332);
nor U40667 (N_40667,N_40469,N_40363);
nor U40668 (N_40668,N_40357,N_40341);
nand U40669 (N_40669,N_40326,N_40434);
nand U40670 (N_40670,N_40440,N_40359);
nand U40671 (N_40671,N_40480,N_40406);
or U40672 (N_40672,N_40266,N_40472);
and U40673 (N_40673,N_40253,N_40329);
and U40674 (N_40674,N_40271,N_40429);
xnor U40675 (N_40675,N_40417,N_40416);
and U40676 (N_40676,N_40256,N_40443);
nand U40677 (N_40677,N_40333,N_40468);
xnor U40678 (N_40678,N_40365,N_40395);
nand U40679 (N_40679,N_40352,N_40448);
and U40680 (N_40680,N_40423,N_40425);
and U40681 (N_40681,N_40416,N_40427);
nor U40682 (N_40682,N_40419,N_40305);
and U40683 (N_40683,N_40262,N_40319);
xnor U40684 (N_40684,N_40349,N_40400);
or U40685 (N_40685,N_40389,N_40455);
nand U40686 (N_40686,N_40282,N_40400);
and U40687 (N_40687,N_40348,N_40323);
nor U40688 (N_40688,N_40401,N_40476);
nand U40689 (N_40689,N_40251,N_40460);
nand U40690 (N_40690,N_40478,N_40268);
and U40691 (N_40691,N_40282,N_40464);
nand U40692 (N_40692,N_40307,N_40460);
nor U40693 (N_40693,N_40491,N_40344);
xnor U40694 (N_40694,N_40344,N_40481);
or U40695 (N_40695,N_40320,N_40367);
nor U40696 (N_40696,N_40402,N_40348);
xnor U40697 (N_40697,N_40449,N_40358);
nor U40698 (N_40698,N_40419,N_40357);
nor U40699 (N_40699,N_40300,N_40342);
or U40700 (N_40700,N_40305,N_40284);
nand U40701 (N_40701,N_40416,N_40316);
and U40702 (N_40702,N_40254,N_40331);
xor U40703 (N_40703,N_40437,N_40330);
and U40704 (N_40704,N_40352,N_40301);
xor U40705 (N_40705,N_40448,N_40408);
nor U40706 (N_40706,N_40344,N_40386);
or U40707 (N_40707,N_40346,N_40479);
nor U40708 (N_40708,N_40359,N_40317);
or U40709 (N_40709,N_40363,N_40430);
and U40710 (N_40710,N_40488,N_40327);
nor U40711 (N_40711,N_40300,N_40411);
and U40712 (N_40712,N_40414,N_40479);
or U40713 (N_40713,N_40444,N_40492);
xor U40714 (N_40714,N_40250,N_40297);
nand U40715 (N_40715,N_40394,N_40479);
nand U40716 (N_40716,N_40311,N_40455);
xor U40717 (N_40717,N_40282,N_40340);
nand U40718 (N_40718,N_40481,N_40414);
or U40719 (N_40719,N_40495,N_40422);
nor U40720 (N_40720,N_40334,N_40269);
and U40721 (N_40721,N_40295,N_40422);
or U40722 (N_40722,N_40346,N_40323);
xor U40723 (N_40723,N_40360,N_40356);
nand U40724 (N_40724,N_40360,N_40358);
nand U40725 (N_40725,N_40422,N_40274);
nand U40726 (N_40726,N_40419,N_40430);
xor U40727 (N_40727,N_40374,N_40325);
xor U40728 (N_40728,N_40336,N_40367);
and U40729 (N_40729,N_40430,N_40403);
or U40730 (N_40730,N_40274,N_40335);
nand U40731 (N_40731,N_40292,N_40317);
xnor U40732 (N_40732,N_40409,N_40279);
and U40733 (N_40733,N_40321,N_40449);
xor U40734 (N_40734,N_40480,N_40301);
nor U40735 (N_40735,N_40360,N_40302);
and U40736 (N_40736,N_40324,N_40431);
and U40737 (N_40737,N_40416,N_40331);
nor U40738 (N_40738,N_40416,N_40471);
xnor U40739 (N_40739,N_40276,N_40304);
nand U40740 (N_40740,N_40448,N_40326);
xor U40741 (N_40741,N_40253,N_40388);
nor U40742 (N_40742,N_40445,N_40454);
nor U40743 (N_40743,N_40479,N_40484);
xor U40744 (N_40744,N_40331,N_40346);
or U40745 (N_40745,N_40269,N_40324);
nand U40746 (N_40746,N_40424,N_40380);
and U40747 (N_40747,N_40276,N_40412);
nor U40748 (N_40748,N_40277,N_40499);
or U40749 (N_40749,N_40390,N_40435);
nand U40750 (N_40750,N_40587,N_40511);
xnor U40751 (N_40751,N_40547,N_40623);
nand U40752 (N_40752,N_40531,N_40745);
or U40753 (N_40753,N_40685,N_40622);
or U40754 (N_40754,N_40570,N_40675);
nor U40755 (N_40755,N_40719,N_40615);
and U40756 (N_40756,N_40559,N_40695);
nor U40757 (N_40757,N_40680,N_40712);
nand U40758 (N_40758,N_40709,N_40744);
nand U40759 (N_40759,N_40542,N_40624);
or U40760 (N_40760,N_40640,N_40525);
xor U40761 (N_40761,N_40657,N_40549);
nand U40762 (N_40762,N_40618,N_40597);
xnor U40763 (N_40763,N_40605,N_40703);
nand U40764 (N_40764,N_40649,N_40563);
and U40765 (N_40765,N_40526,N_40513);
xor U40766 (N_40766,N_40591,N_40550);
xnor U40767 (N_40767,N_40704,N_40508);
or U40768 (N_40768,N_40644,N_40600);
nand U40769 (N_40769,N_40551,N_40669);
nand U40770 (N_40770,N_40598,N_40503);
and U40771 (N_40771,N_40647,N_40656);
nor U40772 (N_40772,N_40571,N_40522);
and U40773 (N_40773,N_40529,N_40552);
or U40774 (N_40774,N_40635,N_40518);
or U40775 (N_40775,N_40737,N_40608);
xnor U40776 (N_40776,N_40504,N_40725);
and U40777 (N_40777,N_40507,N_40642);
xnor U40778 (N_40778,N_40727,N_40683);
and U40779 (N_40779,N_40742,N_40509);
and U40780 (N_40780,N_40710,N_40747);
or U40781 (N_40781,N_40581,N_40662);
and U40782 (N_40782,N_40554,N_40620);
and U40783 (N_40783,N_40674,N_40583);
and U40784 (N_40784,N_40740,N_40735);
xnor U40785 (N_40785,N_40527,N_40702);
nand U40786 (N_40786,N_40588,N_40728);
and U40787 (N_40787,N_40612,N_40520);
or U40788 (N_40788,N_40731,N_40512);
nand U40789 (N_40789,N_40610,N_40564);
nand U40790 (N_40790,N_40652,N_40541);
nor U40791 (N_40791,N_40514,N_40660);
or U40792 (N_40792,N_40500,N_40720);
xor U40793 (N_40793,N_40540,N_40593);
nor U40794 (N_40794,N_40679,N_40546);
and U40795 (N_40795,N_40670,N_40641);
or U40796 (N_40796,N_40714,N_40510);
and U40797 (N_40797,N_40626,N_40700);
xor U40798 (N_40798,N_40613,N_40619);
nand U40799 (N_40799,N_40666,N_40694);
nand U40800 (N_40800,N_40579,N_40566);
xor U40801 (N_40801,N_40711,N_40708);
and U40802 (N_40802,N_40732,N_40736);
nand U40803 (N_40803,N_40734,N_40632);
or U40804 (N_40804,N_40705,N_40606);
or U40805 (N_40805,N_40659,N_40574);
or U40806 (N_40806,N_40722,N_40650);
nor U40807 (N_40807,N_40590,N_40533);
nor U40808 (N_40808,N_40592,N_40611);
and U40809 (N_40809,N_40524,N_40621);
and U40810 (N_40810,N_40603,N_40569);
or U40811 (N_40811,N_40543,N_40672);
nor U40812 (N_40812,N_40578,N_40627);
or U40813 (N_40813,N_40665,N_40690);
or U40814 (N_40814,N_40664,N_40561);
nor U40815 (N_40815,N_40743,N_40538);
xnor U40816 (N_40816,N_40638,N_40733);
nand U40817 (N_40817,N_40607,N_40654);
nand U40818 (N_40818,N_40661,N_40625);
nor U40819 (N_40819,N_40629,N_40609);
or U40820 (N_40820,N_40686,N_40604);
or U40821 (N_40821,N_40658,N_40537);
nand U40822 (N_40822,N_40575,N_40599);
nor U40823 (N_40823,N_40721,N_40730);
xor U40824 (N_40824,N_40678,N_40692);
or U40825 (N_40825,N_40637,N_40601);
xor U40826 (N_40826,N_40596,N_40548);
nor U40827 (N_40827,N_40673,N_40723);
nor U40828 (N_40828,N_40668,N_40651);
xor U40829 (N_40829,N_40653,N_40594);
nand U40830 (N_40830,N_40655,N_40572);
or U40831 (N_40831,N_40616,N_40576);
nand U40832 (N_40832,N_40691,N_40516);
nor U40833 (N_40833,N_40739,N_40687);
and U40834 (N_40834,N_40717,N_40628);
or U40835 (N_40835,N_40699,N_40568);
and U40836 (N_40836,N_40580,N_40681);
xor U40837 (N_40837,N_40617,N_40565);
nand U40838 (N_40838,N_40718,N_40697);
nand U40839 (N_40839,N_40577,N_40741);
xor U40840 (N_40840,N_40724,N_40631);
xnor U40841 (N_40841,N_40532,N_40521);
xor U40842 (N_40842,N_40682,N_40688);
nand U40843 (N_40843,N_40689,N_40636);
or U40844 (N_40844,N_40501,N_40536);
xnor U40845 (N_40845,N_40715,N_40589);
or U40846 (N_40846,N_40676,N_40746);
and U40847 (N_40847,N_40645,N_40584);
nand U40848 (N_40848,N_40671,N_40539);
or U40849 (N_40849,N_40716,N_40544);
or U40850 (N_40850,N_40535,N_40633);
xor U40851 (N_40851,N_40555,N_40560);
nor U40852 (N_40852,N_40582,N_40729);
or U40853 (N_40853,N_40677,N_40523);
nand U40854 (N_40854,N_40602,N_40667);
nor U40855 (N_40855,N_40558,N_40567);
nor U40856 (N_40856,N_40519,N_40562);
nor U40857 (N_40857,N_40634,N_40573);
nand U40858 (N_40858,N_40528,N_40585);
or U40859 (N_40859,N_40698,N_40557);
or U40860 (N_40860,N_40595,N_40696);
nand U40861 (N_40861,N_40713,N_40515);
nor U40862 (N_40862,N_40502,N_40738);
and U40863 (N_40863,N_40749,N_40545);
nor U40864 (N_40864,N_40534,N_40530);
and U40865 (N_40865,N_40684,N_40726);
and U40866 (N_40866,N_40646,N_40517);
nand U40867 (N_40867,N_40701,N_40505);
xor U40868 (N_40868,N_40586,N_40748);
or U40869 (N_40869,N_40639,N_40614);
or U40870 (N_40870,N_40707,N_40648);
xor U40871 (N_40871,N_40663,N_40506);
nor U40872 (N_40872,N_40556,N_40706);
nand U40873 (N_40873,N_40553,N_40643);
nor U40874 (N_40874,N_40693,N_40630);
nand U40875 (N_40875,N_40533,N_40615);
or U40876 (N_40876,N_40734,N_40699);
or U40877 (N_40877,N_40619,N_40720);
nor U40878 (N_40878,N_40654,N_40691);
or U40879 (N_40879,N_40707,N_40680);
nand U40880 (N_40880,N_40596,N_40661);
nand U40881 (N_40881,N_40727,N_40605);
or U40882 (N_40882,N_40669,N_40589);
nor U40883 (N_40883,N_40591,N_40553);
or U40884 (N_40884,N_40565,N_40551);
nor U40885 (N_40885,N_40523,N_40560);
nand U40886 (N_40886,N_40561,N_40623);
nor U40887 (N_40887,N_40595,N_40633);
nor U40888 (N_40888,N_40530,N_40659);
nor U40889 (N_40889,N_40646,N_40564);
nor U40890 (N_40890,N_40506,N_40505);
or U40891 (N_40891,N_40698,N_40748);
nor U40892 (N_40892,N_40512,N_40593);
xor U40893 (N_40893,N_40520,N_40615);
xor U40894 (N_40894,N_40613,N_40659);
and U40895 (N_40895,N_40690,N_40715);
xnor U40896 (N_40896,N_40670,N_40622);
nor U40897 (N_40897,N_40655,N_40659);
nand U40898 (N_40898,N_40665,N_40731);
or U40899 (N_40899,N_40508,N_40532);
nand U40900 (N_40900,N_40681,N_40529);
nor U40901 (N_40901,N_40699,N_40706);
xnor U40902 (N_40902,N_40722,N_40695);
and U40903 (N_40903,N_40528,N_40701);
or U40904 (N_40904,N_40722,N_40737);
xor U40905 (N_40905,N_40675,N_40637);
and U40906 (N_40906,N_40703,N_40527);
or U40907 (N_40907,N_40730,N_40637);
and U40908 (N_40908,N_40559,N_40645);
nor U40909 (N_40909,N_40659,N_40589);
nor U40910 (N_40910,N_40510,N_40684);
and U40911 (N_40911,N_40658,N_40618);
nor U40912 (N_40912,N_40660,N_40555);
nand U40913 (N_40913,N_40641,N_40558);
xnor U40914 (N_40914,N_40676,N_40745);
nand U40915 (N_40915,N_40673,N_40566);
or U40916 (N_40916,N_40540,N_40677);
and U40917 (N_40917,N_40564,N_40680);
or U40918 (N_40918,N_40578,N_40585);
and U40919 (N_40919,N_40691,N_40545);
or U40920 (N_40920,N_40709,N_40666);
xnor U40921 (N_40921,N_40568,N_40743);
nor U40922 (N_40922,N_40711,N_40528);
or U40923 (N_40923,N_40515,N_40717);
nor U40924 (N_40924,N_40621,N_40626);
and U40925 (N_40925,N_40654,N_40519);
and U40926 (N_40926,N_40578,N_40605);
xnor U40927 (N_40927,N_40582,N_40730);
nand U40928 (N_40928,N_40524,N_40556);
and U40929 (N_40929,N_40663,N_40551);
xnor U40930 (N_40930,N_40514,N_40681);
xnor U40931 (N_40931,N_40526,N_40618);
nand U40932 (N_40932,N_40746,N_40620);
nor U40933 (N_40933,N_40529,N_40541);
and U40934 (N_40934,N_40591,N_40613);
and U40935 (N_40935,N_40591,N_40694);
or U40936 (N_40936,N_40702,N_40612);
xnor U40937 (N_40937,N_40678,N_40704);
nand U40938 (N_40938,N_40611,N_40533);
xor U40939 (N_40939,N_40520,N_40531);
and U40940 (N_40940,N_40720,N_40628);
or U40941 (N_40941,N_40525,N_40537);
and U40942 (N_40942,N_40672,N_40696);
and U40943 (N_40943,N_40613,N_40594);
and U40944 (N_40944,N_40643,N_40538);
nor U40945 (N_40945,N_40626,N_40695);
nor U40946 (N_40946,N_40501,N_40700);
xnor U40947 (N_40947,N_40634,N_40524);
or U40948 (N_40948,N_40597,N_40528);
and U40949 (N_40949,N_40619,N_40682);
nand U40950 (N_40950,N_40705,N_40669);
or U40951 (N_40951,N_40711,N_40741);
and U40952 (N_40952,N_40539,N_40703);
nor U40953 (N_40953,N_40621,N_40619);
nand U40954 (N_40954,N_40532,N_40579);
or U40955 (N_40955,N_40708,N_40637);
or U40956 (N_40956,N_40685,N_40694);
nor U40957 (N_40957,N_40505,N_40685);
nor U40958 (N_40958,N_40672,N_40715);
nor U40959 (N_40959,N_40696,N_40631);
nand U40960 (N_40960,N_40732,N_40568);
and U40961 (N_40961,N_40560,N_40738);
or U40962 (N_40962,N_40694,N_40573);
nand U40963 (N_40963,N_40658,N_40570);
xor U40964 (N_40964,N_40657,N_40722);
and U40965 (N_40965,N_40516,N_40731);
or U40966 (N_40966,N_40740,N_40589);
xor U40967 (N_40967,N_40503,N_40586);
nand U40968 (N_40968,N_40573,N_40724);
and U40969 (N_40969,N_40647,N_40641);
nor U40970 (N_40970,N_40668,N_40634);
xnor U40971 (N_40971,N_40745,N_40553);
or U40972 (N_40972,N_40624,N_40650);
xor U40973 (N_40973,N_40594,N_40654);
nor U40974 (N_40974,N_40659,N_40546);
and U40975 (N_40975,N_40592,N_40659);
nor U40976 (N_40976,N_40737,N_40507);
nand U40977 (N_40977,N_40555,N_40607);
or U40978 (N_40978,N_40735,N_40719);
nand U40979 (N_40979,N_40690,N_40686);
nand U40980 (N_40980,N_40540,N_40577);
nor U40981 (N_40981,N_40611,N_40509);
nor U40982 (N_40982,N_40645,N_40596);
xor U40983 (N_40983,N_40626,N_40684);
nor U40984 (N_40984,N_40544,N_40711);
or U40985 (N_40985,N_40520,N_40572);
or U40986 (N_40986,N_40709,N_40718);
or U40987 (N_40987,N_40535,N_40524);
xnor U40988 (N_40988,N_40545,N_40611);
or U40989 (N_40989,N_40646,N_40645);
or U40990 (N_40990,N_40545,N_40610);
nor U40991 (N_40991,N_40713,N_40594);
nand U40992 (N_40992,N_40692,N_40669);
nor U40993 (N_40993,N_40582,N_40607);
and U40994 (N_40994,N_40705,N_40673);
nor U40995 (N_40995,N_40612,N_40530);
and U40996 (N_40996,N_40708,N_40645);
xor U40997 (N_40997,N_40517,N_40518);
nand U40998 (N_40998,N_40671,N_40674);
xor U40999 (N_40999,N_40689,N_40747);
nand U41000 (N_41000,N_40991,N_40859);
or U41001 (N_41001,N_40832,N_40845);
and U41002 (N_41002,N_40757,N_40969);
and U41003 (N_41003,N_40925,N_40872);
xnor U41004 (N_41004,N_40959,N_40971);
nor U41005 (N_41005,N_40780,N_40913);
and U41006 (N_41006,N_40985,N_40867);
nand U41007 (N_41007,N_40766,N_40905);
and U41008 (N_41008,N_40815,N_40956);
and U41009 (N_41009,N_40792,N_40906);
nor U41010 (N_41010,N_40822,N_40938);
and U41011 (N_41011,N_40789,N_40779);
nor U41012 (N_41012,N_40960,N_40941);
nor U41013 (N_41013,N_40948,N_40951);
nor U41014 (N_41014,N_40882,N_40890);
nor U41015 (N_41015,N_40806,N_40914);
or U41016 (N_41016,N_40785,N_40919);
nand U41017 (N_41017,N_40896,N_40894);
xor U41018 (N_41018,N_40835,N_40924);
or U41019 (N_41019,N_40920,N_40841);
nor U41020 (N_41020,N_40831,N_40870);
or U41021 (N_41021,N_40999,N_40825);
nand U41022 (N_41022,N_40937,N_40887);
and U41023 (N_41023,N_40970,N_40878);
and U41024 (N_41024,N_40860,N_40858);
and U41025 (N_41025,N_40814,N_40955);
or U41026 (N_41026,N_40935,N_40799);
nand U41027 (N_41027,N_40972,N_40989);
and U41028 (N_41028,N_40926,N_40994);
nand U41029 (N_41029,N_40921,N_40911);
or U41030 (N_41030,N_40877,N_40833);
and U41031 (N_41031,N_40864,N_40755);
or U41032 (N_41032,N_40945,N_40861);
nand U41033 (N_41033,N_40876,N_40988);
nand U41034 (N_41034,N_40897,N_40764);
xnor U41035 (N_41035,N_40866,N_40886);
or U41036 (N_41036,N_40895,N_40761);
and U41037 (N_41037,N_40852,N_40979);
nand U41038 (N_41038,N_40954,N_40770);
xor U41039 (N_41039,N_40790,N_40856);
xnor U41040 (N_41040,N_40889,N_40810);
nand U41041 (N_41041,N_40869,N_40899);
xor U41042 (N_41042,N_40939,N_40855);
or U41043 (N_41043,N_40928,N_40885);
or U41044 (N_41044,N_40962,N_40909);
xnor U41045 (N_41045,N_40808,N_40838);
nor U41046 (N_41046,N_40823,N_40978);
nand U41047 (N_41047,N_40943,N_40801);
nand U41048 (N_41048,N_40847,N_40908);
nor U41049 (N_41049,N_40863,N_40983);
nor U41050 (N_41050,N_40968,N_40849);
or U41051 (N_41051,N_40839,N_40763);
or U41052 (N_41052,N_40933,N_40884);
xor U41053 (N_41053,N_40756,N_40848);
xor U41054 (N_41054,N_40995,N_40751);
nor U41055 (N_41055,N_40797,N_40977);
and U41056 (N_41056,N_40793,N_40750);
or U41057 (N_41057,N_40944,N_40795);
xnor U41058 (N_41058,N_40987,N_40967);
or U41059 (N_41059,N_40805,N_40850);
nand U41060 (N_41060,N_40929,N_40993);
or U41061 (N_41061,N_40961,N_40986);
nor U41062 (N_41062,N_40786,N_40992);
and U41063 (N_41063,N_40901,N_40871);
nand U41064 (N_41064,N_40762,N_40821);
or U41065 (N_41065,N_40868,N_40932);
xor U41066 (N_41066,N_40875,N_40950);
and U41067 (N_41067,N_40923,N_40990);
and U41068 (N_41068,N_40903,N_40865);
nand U41069 (N_41069,N_40931,N_40794);
and U41070 (N_41070,N_40796,N_40836);
nand U41071 (N_41071,N_40771,N_40759);
nand U41072 (N_41072,N_40862,N_40984);
xnor U41073 (N_41073,N_40980,N_40846);
xor U41074 (N_41074,N_40777,N_40830);
or U41075 (N_41075,N_40964,N_40974);
nand U41076 (N_41076,N_40883,N_40898);
nor U41077 (N_41077,N_40998,N_40879);
xnor U41078 (N_41078,N_40829,N_40791);
and U41079 (N_41079,N_40982,N_40973);
nor U41080 (N_41080,N_40952,N_40840);
and U41081 (N_41081,N_40817,N_40774);
and U41082 (N_41082,N_40881,N_40784);
nor U41083 (N_41083,N_40783,N_40803);
nor U41084 (N_41084,N_40927,N_40853);
nand U41085 (N_41085,N_40843,N_40816);
and U41086 (N_41086,N_40753,N_40778);
nand U41087 (N_41087,N_40976,N_40802);
xnor U41088 (N_41088,N_40874,N_40824);
and U41089 (N_41089,N_40997,N_40891);
and U41090 (N_41090,N_40916,N_40904);
or U41091 (N_41091,N_40813,N_40754);
xor U41092 (N_41092,N_40776,N_40946);
xor U41093 (N_41093,N_40934,N_40775);
xor U41094 (N_41094,N_40782,N_40760);
or U41095 (N_41095,N_40957,N_40981);
or U41096 (N_41096,N_40765,N_40880);
xnor U41097 (N_41097,N_40953,N_40818);
xor U41098 (N_41098,N_40773,N_40918);
nand U41099 (N_41099,N_40902,N_40752);
nor U41100 (N_41100,N_40965,N_40947);
nand U41101 (N_41101,N_40807,N_40975);
nand U41102 (N_41102,N_40788,N_40958);
xor U41103 (N_41103,N_40772,N_40834);
nor U41104 (N_41104,N_40917,N_40893);
nand U41105 (N_41105,N_40963,N_40812);
xnor U41106 (N_41106,N_40851,N_40996);
nand U41107 (N_41107,N_40804,N_40966);
nand U41108 (N_41108,N_40767,N_40842);
nand U41109 (N_41109,N_40768,N_40811);
or U41110 (N_41110,N_40854,N_40907);
nor U41111 (N_41111,N_40857,N_40844);
nor U41112 (N_41112,N_40819,N_40912);
and U41113 (N_41113,N_40809,N_40798);
xnor U41114 (N_41114,N_40769,N_40826);
xnor U41115 (N_41115,N_40936,N_40837);
and U41116 (N_41116,N_40828,N_40942);
nand U41117 (N_41117,N_40888,N_40787);
and U41118 (N_41118,N_40949,N_40940);
and U41119 (N_41119,N_40873,N_40892);
or U41120 (N_41120,N_40910,N_40800);
nor U41121 (N_41121,N_40758,N_40781);
xor U41122 (N_41122,N_40915,N_40922);
xnor U41123 (N_41123,N_40827,N_40930);
nand U41124 (N_41124,N_40820,N_40900);
and U41125 (N_41125,N_40994,N_40948);
nand U41126 (N_41126,N_40932,N_40754);
or U41127 (N_41127,N_40825,N_40844);
and U41128 (N_41128,N_40805,N_40915);
or U41129 (N_41129,N_40769,N_40791);
nand U41130 (N_41130,N_40906,N_40770);
or U41131 (N_41131,N_40975,N_40886);
or U41132 (N_41132,N_40879,N_40994);
or U41133 (N_41133,N_40886,N_40810);
and U41134 (N_41134,N_40750,N_40998);
nand U41135 (N_41135,N_40936,N_40876);
and U41136 (N_41136,N_40753,N_40967);
and U41137 (N_41137,N_40874,N_40807);
nand U41138 (N_41138,N_40989,N_40889);
and U41139 (N_41139,N_40925,N_40808);
or U41140 (N_41140,N_40782,N_40819);
xnor U41141 (N_41141,N_40880,N_40976);
xor U41142 (N_41142,N_40753,N_40883);
and U41143 (N_41143,N_40827,N_40912);
xnor U41144 (N_41144,N_40927,N_40961);
nand U41145 (N_41145,N_40835,N_40935);
and U41146 (N_41146,N_40847,N_40895);
xor U41147 (N_41147,N_40866,N_40763);
nand U41148 (N_41148,N_40756,N_40858);
nor U41149 (N_41149,N_40772,N_40985);
and U41150 (N_41150,N_40788,N_40852);
or U41151 (N_41151,N_40992,N_40923);
or U41152 (N_41152,N_40929,N_40958);
nor U41153 (N_41153,N_40841,N_40881);
xor U41154 (N_41154,N_40859,N_40869);
xor U41155 (N_41155,N_40934,N_40843);
and U41156 (N_41156,N_40986,N_40926);
or U41157 (N_41157,N_40814,N_40889);
xor U41158 (N_41158,N_40989,N_40877);
xnor U41159 (N_41159,N_40865,N_40913);
nand U41160 (N_41160,N_40810,N_40870);
and U41161 (N_41161,N_40815,N_40977);
or U41162 (N_41162,N_40950,N_40907);
or U41163 (N_41163,N_40921,N_40835);
and U41164 (N_41164,N_40855,N_40940);
xor U41165 (N_41165,N_40885,N_40761);
nand U41166 (N_41166,N_40825,N_40880);
nor U41167 (N_41167,N_40915,N_40797);
xor U41168 (N_41168,N_40925,N_40866);
or U41169 (N_41169,N_40926,N_40801);
nor U41170 (N_41170,N_40848,N_40996);
nand U41171 (N_41171,N_40963,N_40784);
nor U41172 (N_41172,N_40790,N_40892);
xnor U41173 (N_41173,N_40831,N_40913);
nor U41174 (N_41174,N_40840,N_40787);
xor U41175 (N_41175,N_40813,N_40799);
nand U41176 (N_41176,N_40827,N_40943);
xnor U41177 (N_41177,N_40908,N_40799);
nand U41178 (N_41178,N_40952,N_40835);
nor U41179 (N_41179,N_40916,N_40999);
and U41180 (N_41180,N_40856,N_40900);
and U41181 (N_41181,N_40876,N_40859);
and U41182 (N_41182,N_40825,N_40874);
nor U41183 (N_41183,N_40772,N_40755);
or U41184 (N_41184,N_40909,N_40986);
nor U41185 (N_41185,N_40993,N_40915);
or U41186 (N_41186,N_40858,N_40896);
nand U41187 (N_41187,N_40927,N_40999);
xor U41188 (N_41188,N_40932,N_40762);
and U41189 (N_41189,N_40999,N_40861);
xor U41190 (N_41190,N_40905,N_40823);
or U41191 (N_41191,N_40845,N_40831);
and U41192 (N_41192,N_40886,N_40895);
nor U41193 (N_41193,N_40883,N_40878);
nor U41194 (N_41194,N_40937,N_40881);
nand U41195 (N_41195,N_40762,N_40827);
xor U41196 (N_41196,N_40830,N_40988);
nor U41197 (N_41197,N_40760,N_40990);
and U41198 (N_41198,N_40815,N_40847);
nand U41199 (N_41199,N_40932,N_40836);
nor U41200 (N_41200,N_40860,N_40978);
nor U41201 (N_41201,N_40959,N_40943);
nor U41202 (N_41202,N_40958,N_40939);
or U41203 (N_41203,N_40967,N_40804);
and U41204 (N_41204,N_40809,N_40767);
xnor U41205 (N_41205,N_40917,N_40973);
xor U41206 (N_41206,N_40856,N_40771);
xor U41207 (N_41207,N_40990,N_40882);
xor U41208 (N_41208,N_40985,N_40925);
nor U41209 (N_41209,N_40778,N_40834);
nand U41210 (N_41210,N_40951,N_40970);
nand U41211 (N_41211,N_40870,N_40992);
and U41212 (N_41212,N_40986,N_40964);
or U41213 (N_41213,N_40830,N_40955);
nor U41214 (N_41214,N_40760,N_40977);
xor U41215 (N_41215,N_40988,N_40996);
nand U41216 (N_41216,N_40931,N_40910);
or U41217 (N_41217,N_40975,N_40824);
nand U41218 (N_41218,N_40899,N_40753);
nor U41219 (N_41219,N_40910,N_40935);
nor U41220 (N_41220,N_40766,N_40762);
xor U41221 (N_41221,N_40981,N_40894);
nand U41222 (N_41222,N_40777,N_40835);
or U41223 (N_41223,N_40809,N_40816);
nand U41224 (N_41224,N_40762,N_40783);
nand U41225 (N_41225,N_40901,N_40976);
xor U41226 (N_41226,N_40956,N_40895);
nand U41227 (N_41227,N_40755,N_40879);
nand U41228 (N_41228,N_40752,N_40853);
nand U41229 (N_41229,N_40925,N_40951);
nor U41230 (N_41230,N_40908,N_40973);
nor U41231 (N_41231,N_40796,N_40855);
xnor U41232 (N_41232,N_40916,N_40970);
nand U41233 (N_41233,N_40947,N_40808);
and U41234 (N_41234,N_40958,N_40828);
xnor U41235 (N_41235,N_40858,N_40949);
or U41236 (N_41236,N_40938,N_40835);
and U41237 (N_41237,N_40804,N_40900);
and U41238 (N_41238,N_40771,N_40805);
nor U41239 (N_41239,N_40911,N_40773);
nand U41240 (N_41240,N_40877,N_40988);
and U41241 (N_41241,N_40875,N_40835);
xnor U41242 (N_41242,N_40905,N_40957);
nor U41243 (N_41243,N_40768,N_40860);
nor U41244 (N_41244,N_40760,N_40853);
and U41245 (N_41245,N_40968,N_40795);
nand U41246 (N_41246,N_40770,N_40871);
and U41247 (N_41247,N_40761,N_40829);
nand U41248 (N_41248,N_40847,N_40974);
or U41249 (N_41249,N_40852,N_40754);
xor U41250 (N_41250,N_41211,N_41066);
xor U41251 (N_41251,N_41031,N_41101);
and U41252 (N_41252,N_41103,N_41012);
xnor U41253 (N_41253,N_41200,N_41083);
nor U41254 (N_41254,N_41227,N_41069);
xor U41255 (N_41255,N_41023,N_41122);
and U41256 (N_41256,N_41198,N_41123);
xnor U41257 (N_41257,N_41051,N_41222);
or U41258 (N_41258,N_41099,N_41174);
nor U41259 (N_41259,N_41243,N_41040);
nand U41260 (N_41260,N_41048,N_41027);
nor U41261 (N_41261,N_41148,N_41055);
and U41262 (N_41262,N_41005,N_41004);
or U41263 (N_41263,N_41114,N_41249);
and U41264 (N_41264,N_41244,N_41079);
xor U41265 (N_41265,N_41229,N_41093);
or U41266 (N_41266,N_41224,N_41098);
or U41267 (N_41267,N_41176,N_41213);
xor U41268 (N_41268,N_41155,N_41000);
or U41269 (N_41269,N_41164,N_41014);
and U41270 (N_41270,N_41020,N_41100);
and U41271 (N_41271,N_41218,N_41199);
nand U41272 (N_41272,N_41158,N_41120);
and U41273 (N_41273,N_41003,N_41172);
nor U41274 (N_41274,N_41095,N_41248);
or U41275 (N_41275,N_41077,N_41130);
and U41276 (N_41276,N_41043,N_41065);
and U41277 (N_41277,N_41221,N_41135);
xnor U41278 (N_41278,N_41163,N_41235);
nand U41279 (N_41279,N_41226,N_41237);
or U41280 (N_41280,N_41220,N_41029);
and U41281 (N_41281,N_41178,N_41032);
nor U41282 (N_41282,N_41175,N_41133);
and U41283 (N_41283,N_41016,N_41245);
xor U41284 (N_41284,N_41106,N_41063);
nor U41285 (N_41285,N_41137,N_41088);
nand U41286 (N_41286,N_41109,N_41072);
xnor U41287 (N_41287,N_41052,N_41210);
xnor U41288 (N_41288,N_41037,N_41057);
nor U41289 (N_41289,N_41042,N_41017);
or U41290 (N_41290,N_41025,N_41024);
xnor U41291 (N_41291,N_41151,N_41149);
xor U41292 (N_41292,N_41215,N_41168);
or U41293 (N_41293,N_41097,N_41087);
nand U41294 (N_41294,N_41105,N_41108);
or U41295 (N_41295,N_41241,N_41019);
and U41296 (N_41296,N_41080,N_41177);
xnor U41297 (N_41297,N_41138,N_41026);
or U41298 (N_41298,N_41152,N_41081);
xor U41299 (N_41299,N_41143,N_41056);
xor U41300 (N_41300,N_41146,N_41038);
xor U41301 (N_41301,N_41184,N_41110);
nand U41302 (N_41302,N_41239,N_41188);
or U41303 (N_41303,N_41233,N_41159);
and U41304 (N_41304,N_41107,N_41113);
nor U41305 (N_41305,N_41228,N_41160);
and U41306 (N_41306,N_41161,N_41242);
nand U41307 (N_41307,N_41018,N_41115);
and U41308 (N_41308,N_41028,N_41201);
nor U41309 (N_41309,N_41092,N_41119);
nor U41310 (N_41310,N_41142,N_41231);
nand U41311 (N_41311,N_41207,N_41140);
nor U41312 (N_41312,N_41147,N_41185);
nor U41313 (N_41313,N_41195,N_41121);
nor U41314 (N_41314,N_41015,N_41202);
nand U41315 (N_41315,N_41154,N_41205);
xor U41316 (N_41316,N_41236,N_41167);
nor U41317 (N_41317,N_41219,N_41203);
nand U41318 (N_41318,N_41190,N_41011);
or U41319 (N_41319,N_41234,N_41086);
xor U41320 (N_41320,N_41127,N_41041);
and U41321 (N_41321,N_41094,N_41156);
or U41322 (N_41322,N_41125,N_41002);
or U41323 (N_41323,N_41145,N_41096);
and U41324 (N_41324,N_41010,N_41171);
nor U41325 (N_41325,N_41075,N_41084);
xnor U41326 (N_41326,N_41074,N_41071);
nor U41327 (N_41327,N_41208,N_41078);
or U41328 (N_41328,N_41197,N_41008);
and U41329 (N_41329,N_41194,N_41131);
nor U41330 (N_41330,N_41001,N_41036);
or U41331 (N_41331,N_41047,N_41021);
nor U41332 (N_41332,N_41247,N_41064);
or U41333 (N_41333,N_41013,N_41193);
and U41334 (N_41334,N_41166,N_41124);
xor U41335 (N_41335,N_41134,N_41223);
and U41336 (N_41336,N_41196,N_41091);
nor U41337 (N_41337,N_41090,N_41112);
nand U41338 (N_41338,N_41191,N_41181);
nand U41339 (N_41339,N_41116,N_41150);
nand U41340 (N_41340,N_41240,N_41053);
nor U41341 (N_41341,N_41006,N_41173);
or U41342 (N_41342,N_41232,N_41192);
xor U41343 (N_41343,N_41076,N_41157);
xor U41344 (N_41344,N_41165,N_41246);
and U41345 (N_41345,N_41111,N_41030);
xnor U41346 (N_41346,N_41186,N_41129);
or U41347 (N_41347,N_41007,N_41139);
nor U41348 (N_41348,N_41216,N_41126);
nand U41349 (N_41349,N_41070,N_41060);
nand U41350 (N_41350,N_41238,N_41034);
xor U41351 (N_41351,N_41180,N_41214);
nor U41352 (N_41352,N_41022,N_41204);
xnor U41353 (N_41353,N_41189,N_41049);
xor U41354 (N_41354,N_41061,N_41187);
nand U41355 (N_41355,N_41144,N_41054);
and U41356 (N_41356,N_41117,N_41044);
or U41357 (N_41357,N_41141,N_41118);
nor U41358 (N_41358,N_41104,N_41062);
or U41359 (N_41359,N_41089,N_41225);
xor U41360 (N_41360,N_41082,N_41183);
xnor U41361 (N_41361,N_41102,N_41073);
nor U41362 (N_41362,N_41179,N_41153);
and U41363 (N_41363,N_41067,N_41039);
and U41364 (N_41364,N_41136,N_41033);
xor U41365 (N_41365,N_41217,N_41182);
or U41366 (N_41366,N_41206,N_41230);
or U41367 (N_41367,N_41059,N_41128);
and U41368 (N_41368,N_41045,N_41132);
and U41369 (N_41369,N_41085,N_41058);
or U41370 (N_41370,N_41068,N_41046);
and U41371 (N_41371,N_41162,N_41170);
nor U41372 (N_41372,N_41209,N_41050);
and U41373 (N_41373,N_41009,N_41169);
and U41374 (N_41374,N_41212,N_41035);
nand U41375 (N_41375,N_41020,N_41103);
xnor U41376 (N_41376,N_41091,N_41051);
xnor U41377 (N_41377,N_41160,N_41152);
and U41378 (N_41378,N_41016,N_41051);
nor U41379 (N_41379,N_41098,N_41108);
or U41380 (N_41380,N_41169,N_41059);
nor U41381 (N_41381,N_41246,N_41040);
or U41382 (N_41382,N_41051,N_41180);
nand U41383 (N_41383,N_41133,N_41013);
or U41384 (N_41384,N_41075,N_41083);
or U41385 (N_41385,N_41242,N_41054);
xor U41386 (N_41386,N_41132,N_41122);
and U41387 (N_41387,N_41048,N_41241);
nor U41388 (N_41388,N_41002,N_41094);
nor U41389 (N_41389,N_41047,N_41098);
nor U41390 (N_41390,N_41224,N_41030);
xor U41391 (N_41391,N_41108,N_41134);
xnor U41392 (N_41392,N_41014,N_41171);
nand U41393 (N_41393,N_41144,N_41241);
or U41394 (N_41394,N_41232,N_41201);
nor U41395 (N_41395,N_41040,N_41135);
nand U41396 (N_41396,N_41129,N_41045);
xnor U41397 (N_41397,N_41238,N_41134);
and U41398 (N_41398,N_41171,N_41132);
nand U41399 (N_41399,N_41067,N_41115);
xnor U41400 (N_41400,N_41188,N_41090);
nor U41401 (N_41401,N_41142,N_41048);
xnor U41402 (N_41402,N_41108,N_41004);
and U41403 (N_41403,N_41156,N_41133);
or U41404 (N_41404,N_41045,N_41082);
nor U41405 (N_41405,N_41164,N_41027);
and U41406 (N_41406,N_41038,N_41132);
or U41407 (N_41407,N_41191,N_41201);
nand U41408 (N_41408,N_41081,N_41091);
xor U41409 (N_41409,N_41094,N_41226);
nand U41410 (N_41410,N_41126,N_41036);
nand U41411 (N_41411,N_41037,N_41165);
nand U41412 (N_41412,N_41109,N_41105);
and U41413 (N_41413,N_41188,N_41221);
xor U41414 (N_41414,N_41026,N_41160);
or U41415 (N_41415,N_41048,N_41189);
or U41416 (N_41416,N_41179,N_41057);
and U41417 (N_41417,N_41219,N_41239);
nand U41418 (N_41418,N_41093,N_41008);
or U41419 (N_41419,N_41048,N_41238);
nand U41420 (N_41420,N_41028,N_41157);
nor U41421 (N_41421,N_41119,N_41200);
xnor U41422 (N_41422,N_41187,N_41192);
and U41423 (N_41423,N_41051,N_41027);
nor U41424 (N_41424,N_41017,N_41077);
nor U41425 (N_41425,N_41011,N_41242);
or U41426 (N_41426,N_41067,N_41200);
and U41427 (N_41427,N_41050,N_41025);
and U41428 (N_41428,N_41235,N_41131);
xnor U41429 (N_41429,N_41183,N_41050);
or U41430 (N_41430,N_41212,N_41042);
nand U41431 (N_41431,N_41126,N_41218);
nor U41432 (N_41432,N_41038,N_41186);
or U41433 (N_41433,N_41197,N_41102);
and U41434 (N_41434,N_41241,N_41197);
xor U41435 (N_41435,N_41188,N_41037);
xor U41436 (N_41436,N_41235,N_41008);
and U41437 (N_41437,N_41136,N_41103);
and U41438 (N_41438,N_41221,N_41016);
or U41439 (N_41439,N_41005,N_41194);
nor U41440 (N_41440,N_41231,N_41160);
and U41441 (N_41441,N_41244,N_41234);
or U41442 (N_41442,N_41189,N_41106);
nor U41443 (N_41443,N_41082,N_41041);
and U41444 (N_41444,N_41014,N_41056);
xor U41445 (N_41445,N_41105,N_41244);
nor U41446 (N_41446,N_41222,N_41114);
and U41447 (N_41447,N_41021,N_41012);
xor U41448 (N_41448,N_41029,N_41089);
xor U41449 (N_41449,N_41081,N_41084);
nor U41450 (N_41450,N_41101,N_41214);
and U41451 (N_41451,N_41014,N_41197);
xor U41452 (N_41452,N_41117,N_41150);
and U41453 (N_41453,N_41076,N_41194);
and U41454 (N_41454,N_41026,N_41066);
or U41455 (N_41455,N_41091,N_41067);
and U41456 (N_41456,N_41070,N_41045);
nor U41457 (N_41457,N_41117,N_41079);
nand U41458 (N_41458,N_41046,N_41141);
and U41459 (N_41459,N_41134,N_41205);
and U41460 (N_41460,N_41193,N_41067);
or U41461 (N_41461,N_41156,N_41105);
nor U41462 (N_41462,N_41083,N_41177);
nor U41463 (N_41463,N_41237,N_41004);
xnor U41464 (N_41464,N_41203,N_41143);
or U41465 (N_41465,N_41245,N_41066);
or U41466 (N_41466,N_41079,N_41169);
nand U41467 (N_41467,N_41017,N_41192);
xor U41468 (N_41468,N_41033,N_41078);
nor U41469 (N_41469,N_41043,N_41201);
and U41470 (N_41470,N_41194,N_41191);
nor U41471 (N_41471,N_41058,N_41234);
nor U41472 (N_41472,N_41036,N_41077);
xnor U41473 (N_41473,N_41099,N_41143);
xor U41474 (N_41474,N_41165,N_41173);
and U41475 (N_41475,N_41225,N_41149);
or U41476 (N_41476,N_41017,N_41174);
and U41477 (N_41477,N_41146,N_41158);
and U41478 (N_41478,N_41225,N_41214);
nor U41479 (N_41479,N_41175,N_41030);
and U41480 (N_41480,N_41091,N_41039);
and U41481 (N_41481,N_41248,N_41070);
and U41482 (N_41482,N_41040,N_41095);
xor U41483 (N_41483,N_41131,N_41167);
xor U41484 (N_41484,N_41037,N_41031);
and U41485 (N_41485,N_41108,N_41028);
nor U41486 (N_41486,N_41237,N_41013);
nor U41487 (N_41487,N_41185,N_41015);
nor U41488 (N_41488,N_41190,N_41242);
and U41489 (N_41489,N_41052,N_41141);
nor U41490 (N_41490,N_41185,N_41191);
nor U41491 (N_41491,N_41013,N_41037);
xor U41492 (N_41492,N_41204,N_41207);
nand U41493 (N_41493,N_41162,N_41016);
or U41494 (N_41494,N_41033,N_41140);
or U41495 (N_41495,N_41173,N_41023);
xor U41496 (N_41496,N_41060,N_41072);
and U41497 (N_41497,N_41126,N_41073);
nor U41498 (N_41498,N_41054,N_41239);
and U41499 (N_41499,N_41150,N_41095);
nor U41500 (N_41500,N_41256,N_41339);
and U41501 (N_41501,N_41350,N_41309);
and U41502 (N_41502,N_41363,N_41406);
nand U41503 (N_41503,N_41462,N_41328);
and U41504 (N_41504,N_41314,N_41332);
or U41505 (N_41505,N_41496,N_41338);
or U41506 (N_41506,N_41492,N_41424);
and U41507 (N_41507,N_41478,N_41342);
xor U41508 (N_41508,N_41439,N_41284);
nand U41509 (N_41509,N_41355,N_41412);
xor U41510 (N_41510,N_41446,N_41413);
nor U41511 (N_41511,N_41428,N_41254);
or U41512 (N_41512,N_41469,N_41385);
or U41513 (N_41513,N_41408,N_41487);
nor U41514 (N_41514,N_41497,N_41366);
xor U41515 (N_41515,N_41384,N_41281);
and U41516 (N_41516,N_41357,N_41272);
nand U41517 (N_41517,N_41485,N_41300);
nand U41518 (N_41518,N_41321,N_41377);
and U41519 (N_41519,N_41333,N_41459);
nor U41520 (N_41520,N_41419,N_41450);
xor U41521 (N_41521,N_41489,N_41463);
nor U41522 (N_41522,N_41390,N_41398);
nor U41523 (N_41523,N_41343,N_41375);
nand U41524 (N_41524,N_41494,N_41417);
nand U41525 (N_41525,N_41451,N_41251);
nand U41526 (N_41526,N_41416,N_41275);
and U41527 (N_41527,N_41449,N_41286);
nand U41528 (N_41528,N_41486,N_41257);
or U41529 (N_41529,N_41381,N_41279);
and U41530 (N_41530,N_41336,N_41443);
nor U41531 (N_41531,N_41306,N_41269);
nor U41532 (N_41532,N_41358,N_41312);
nor U41533 (N_41533,N_41488,N_41456);
or U41534 (N_41534,N_41356,N_41368);
nor U41535 (N_41535,N_41442,N_41266);
or U41536 (N_41536,N_41397,N_41404);
nor U41537 (N_41537,N_41431,N_41430);
and U41538 (N_41538,N_41274,N_41411);
or U41539 (N_41539,N_41380,N_41340);
and U41540 (N_41540,N_41295,N_41301);
nor U41541 (N_41541,N_41460,N_41435);
or U41542 (N_41542,N_41308,N_41371);
or U41543 (N_41543,N_41317,N_41353);
and U41544 (N_41544,N_41255,N_41334);
or U41545 (N_41545,N_41327,N_41464);
xnor U41546 (N_41546,N_41493,N_41258);
or U41547 (N_41547,N_41311,N_41268);
nor U41548 (N_41548,N_41318,N_41396);
nor U41549 (N_41549,N_41283,N_41470);
nor U41550 (N_41550,N_41364,N_41369);
xor U41551 (N_41551,N_41346,N_41466);
or U41552 (N_41552,N_41252,N_41427);
or U41553 (N_41553,N_41289,N_41432);
or U41554 (N_41554,N_41293,N_41423);
and U41555 (N_41555,N_41324,N_41482);
and U41556 (N_41556,N_41323,N_41325);
nand U41557 (N_41557,N_41345,N_41278);
nand U41558 (N_41558,N_41326,N_41457);
or U41559 (N_41559,N_41331,N_41426);
nor U41560 (N_41560,N_41479,N_41480);
xnor U41561 (N_41561,N_41296,N_41445);
or U41562 (N_41562,N_41273,N_41261);
or U41563 (N_41563,N_41483,N_41316);
or U41564 (N_41564,N_41407,N_41448);
or U41565 (N_41565,N_41253,N_41382);
nand U41566 (N_41566,N_41472,N_41418);
xnor U41567 (N_41567,N_41389,N_41265);
nand U41568 (N_41568,N_41499,N_41474);
xnor U41569 (N_41569,N_41498,N_41458);
nor U41570 (N_41570,N_41271,N_41399);
nand U41571 (N_41571,N_41280,N_41490);
xor U41572 (N_41572,N_41402,N_41422);
nor U41573 (N_41573,N_41319,N_41374);
nor U41574 (N_41574,N_41467,N_41347);
and U41575 (N_41575,N_41436,N_41276);
xor U41576 (N_41576,N_41444,N_41387);
xor U41577 (N_41577,N_41259,N_41373);
or U41578 (N_41578,N_41378,N_41270);
nor U41579 (N_41579,N_41437,N_41414);
nand U41580 (N_41580,N_41393,N_41302);
xor U41581 (N_41581,N_41330,N_41433);
nor U41582 (N_41582,N_41349,N_41354);
nor U41583 (N_41583,N_41307,N_41425);
or U41584 (N_41584,N_41304,N_41298);
and U41585 (N_41585,N_41351,N_41322);
nand U41586 (N_41586,N_41484,N_41438);
and U41587 (N_41587,N_41415,N_41305);
nor U41588 (N_41588,N_41313,N_41361);
nand U41589 (N_41589,N_41344,N_41477);
xnor U41590 (N_41590,N_41491,N_41287);
and U41591 (N_41591,N_41352,N_41409);
and U41592 (N_41592,N_41453,N_41394);
or U41593 (N_41593,N_41359,N_41447);
xnor U41594 (N_41594,N_41495,N_41277);
and U41595 (N_41595,N_41370,N_41262);
nor U41596 (N_41596,N_41362,N_41383);
xnor U41597 (N_41597,N_41291,N_41476);
nor U41598 (N_41598,N_41454,N_41299);
or U41599 (N_41599,N_41310,N_41434);
or U41600 (N_41600,N_41282,N_41440);
and U41601 (N_41601,N_41263,N_41337);
and U41602 (N_41602,N_41303,N_41481);
or U41603 (N_41603,N_41391,N_41461);
and U41604 (N_41604,N_41379,N_41285);
nand U41605 (N_41605,N_41260,N_41267);
nor U41606 (N_41606,N_41441,N_41401);
xor U41607 (N_41607,N_41395,N_41315);
and U41608 (N_41608,N_41341,N_41360);
nand U41609 (N_41609,N_41335,N_41365);
or U41610 (N_41610,N_41367,N_41388);
nand U41611 (N_41611,N_41320,N_41372);
nand U41612 (N_41612,N_41386,N_41465);
xor U41613 (N_41613,N_41292,N_41329);
nor U41614 (N_41614,N_41455,N_41452);
xnor U41615 (N_41615,N_41475,N_41429);
xnor U41616 (N_41616,N_41421,N_41290);
or U41617 (N_41617,N_41348,N_41473);
or U41618 (N_41618,N_41376,N_41468);
xnor U41619 (N_41619,N_41250,N_41405);
nand U41620 (N_41620,N_41420,N_41403);
or U41621 (N_41621,N_41264,N_41294);
and U41622 (N_41622,N_41471,N_41392);
xor U41623 (N_41623,N_41288,N_41297);
and U41624 (N_41624,N_41400,N_41410);
xnor U41625 (N_41625,N_41309,N_41400);
xor U41626 (N_41626,N_41449,N_41388);
or U41627 (N_41627,N_41496,N_41483);
or U41628 (N_41628,N_41276,N_41444);
or U41629 (N_41629,N_41433,N_41445);
nor U41630 (N_41630,N_41451,N_41469);
or U41631 (N_41631,N_41394,N_41347);
or U41632 (N_41632,N_41386,N_41490);
and U41633 (N_41633,N_41477,N_41290);
nand U41634 (N_41634,N_41469,N_41389);
and U41635 (N_41635,N_41345,N_41374);
and U41636 (N_41636,N_41273,N_41264);
xnor U41637 (N_41637,N_41383,N_41418);
xor U41638 (N_41638,N_41453,N_41437);
nand U41639 (N_41639,N_41388,N_41431);
and U41640 (N_41640,N_41436,N_41260);
nand U41641 (N_41641,N_41278,N_41270);
xnor U41642 (N_41642,N_41496,N_41430);
xor U41643 (N_41643,N_41345,N_41454);
xor U41644 (N_41644,N_41485,N_41455);
nand U41645 (N_41645,N_41410,N_41490);
and U41646 (N_41646,N_41355,N_41288);
and U41647 (N_41647,N_41473,N_41360);
or U41648 (N_41648,N_41320,N_41365);
nor U41649 (N_41649,N_41330,N_41338);
xnor U41650 (N_41650,N_41489,N_41362);
xnor U41651 (N_41651,N_41310,N_41329);
nand U41652 (N_41652,N_41414,N_41349);
nand U41653 (N_41653,N_41290,N_41293);
nand U41654 (N_41654,N_41408,N_41343);
or U41655 (N_41655,N_41394,N_41465);
or U41656 (N_41656,N_41371,N_41394);
nand U41657 (N_41657,N_41375,N_41330);
nor U41658 (N_41658,N_41369,N_41415);
and U41659 (N_41659,N_41441,N_41446);
and U41660 (N_41660,N_41255,N_41343);
or U41661 (N_41661,N_41347,N_41405);
and U41662 (N_41662,N_41286,N_41259);
xnor U41663 (N_41663,N_41417,N_41305);
and U41664 (N_41664,N_41487,N_41442);
or U41665 (N_41665,N_41315,N_41365);
or U41666 (N_41666,N_41434,N_41353);
xor U41667 (N_41667,N_41346,N_41339);
or U41668 (N_41668,N_41286,N_41470);
and U41669 (N_41669,N_41269,N_41373);
xnor U41670 (N_41670,N_41401,N_41309);
nand U41671 (N_41671,N_41307,N_41457);
xor U41672 (N_41672,N_41377,N_41409);
or U41673 (N_41673,N_41326,N_41329);
nand U41674 (N_41674,N_41465,N_41320);
and U41675 (N_41675,N_41407,N_41475);
and U41676 (N_41676,N_41469,N_41443);
nand U41677 (N_41677,N_41413,N_41296);
nor U41678 (N_41678,N_41262,N_41269);
nor U41679 (N_41679,N_41389,N_41328);
nand U41680 (N_41680,N_41386,N_41385);
xor U41681 (N_41681,N_41386,N_41357);
xor U41682 (N_41682,N_41356,N_41497);
or U41683 (N_41683,N_41491,N_41291);
nor U41684 (N_41684,N_41312,N_41404);
nor U41685 (N_41685,N_41351,N_41380);
nand U41686 (N_41686,N_41363,N_41342);
nand U41687 (N_41687,N_41357,N_41483);
and U41688 (N_41688,N_41397,N_41484);
or U41689 (N_41689,N_41414,N_41415);
or U41690 (N_41690,N_41386,N_41369);
nor U41691 (N_41691,N_41257,N_41459);
and U41692 (N_41692,N_41448,N_41429);
nand U41693 (N_41693,N_41268,N_41493);
xnor U41694 (N_41694,N_41251,N_41414);
or U41695 (N_41695,N_41325,N_41400);
xnor U41696 (N_41696,N_41413,N_41265);
nand U41697 (N_41697,N_41427,N_41420);
and U41698 (N_41698,N_41416,N_41287);
nor U41699 (N_41699,N_41383,N_41320);
or U41700 (N_41700,N_41320,N_41337);
and U41701 (N_41701,N_41266,N_41260);
and U41702 (N_41702,N_41422,N_41348);
nor U41703 (N_41703,N_41302,N_41261);
and U41704 (N_41704,N_41453,N_41471);
xor U41705 (N_41705,N_41326,N_41303);
or U41706 (N_41706,N_41281,N_41250);
and U41707 (N_41707,N_41272,N_41297);
xor U41708 (N_41708,N_41420,N_41385);
nand U41709 (N_41709,N_41361,N_41271);
or U41710 (N_41710,N_41420,N_41475);
xnor U41711 (N_41711,N_41397,N_41363);
nand U41712 (N_41712,N_41290,N_41314);
and U41713 (N_41713,N_41476,N_41471);
nand U41714 (N_41714,N_41254,N_41321);
xnor U41715 (N_41715,N_41303,N_41486);
nor U41716 (N_41716,N_41375,N_41350);
nor U41717 (N_41717,N_41441,N_41431);
and U41718 (N_41718,N_41258,N_41291);
and U41719 (N_41719,N_41286,N_41388);
nand U41720 (N_41720,N_41271,N_41358);
or U41721 (N_41721,N_41363,N_41251);
nor U41722 (N_41722,N_41383,N_41465);
nor U41723 (N_41723,N_41490,N_41336);
and U41724 (N_41724,N_41297,N_41330);
and U41725 (N_41725,N_41385,N_41450);
or U41726 (N_41726,N_41310,N_41337);
xor U41727 (N_41727,N_41484,N_41481);
nor U41728 (N_41728,N_41340,N_41344);
or U41729 (N_41729,N_41435,N_41253);
xor U41730 (N_41730,N_41311,N_41451);
xnor U41731 (N_41731,N_41299,N_41253);
nor U41732 (N_41732,N_41496,N_41270);
xor U41733 (N_41733,N_41426,N_41364);
nor U41734 (N_41734,N_41262,N_41289);
xnor U41735 (N_41735,N_41313,N_41294);
xnor U41736 (N_41736,N_41441,N_41319);
or U41737 (N_41737,N_41322,N_41432);
xnor U41738 (N_41738,N_41461,N_41340);
nand U41739 (N_41739,N_41311,N_41302);
and U41740 (N_41740,N_41492,N_41250);
or U41741 (N_41741,N_41490,N_41392);
nand U41742 (N_41742,N_41491,N_41457);
xnor U41743 (N_41743,N_41330,N_41369);
and U41744 (N_41744,N_41399,N_41304);
and U41745 (N_41745,N_41321,N_41290);
xor U41746 (N_41746,N_41488,N_41310);
nand U41747 (N_41747,N_41460,N_41276);
and U41748 (N_41748,N_41482,N_41254);
xnor U41749 (N_41749,N_41303,N_41302);
nand U41750 (N_41750,N_41681,N_41602);
and U41751 (N_41751,N_41518,N_41568);
nand U41752 (N_41752,N_41668,N_41587);
or U41753 (N_41753,N_41590,N_41584);
nor U41754 (N_41754,N_41510,N_41674);
or U41755 (N_41755,N_41539,N_41549);
or U41756 (N_41756,N_41745,N_41593);
xnor U41757 (N_41757,N_41601,N_41582);
xnor U41758 (N_41758,N_41722,N_41702);
nand U41759 (N_41759,N_41511,N_41588);
or U41760 (N_41760,N_41527,N_41652);
and U41761 (N_41761,N_41565,N_41731);
nor U41762 (N_41762,N_41585,N_41739);
nand U41763 (N_41763,N_41547,N_41572);
nor U41764 (N_41764,N_41623,N_41642);
xnor U41765 (N_41765,N_41729,N_41621);
nor U41766 (N_41766,N_41727,N_41506);
or U41767 (N_41767,N_41573,N_41569);
nand U41768 (N_41768,N_41715,N_41699);
and U41769 (N_41769,N_41736,N_41649);
or U41770 (N_41770,N_41567,N_41686);
xnor U41771 (N_41771,N_41589,N_41576);
nand U41772 (N_41772,N_41720,N_41599);
or U41773 (N_41773,N_41716,N_41734);
nand U41774 (N_41774,N_41581,N_41579);
or U41775 (N_41775,N_41710,N_41563);
nor U41776 (N_41776,N_41651,N_41682);
nand U41777 (N_41777,N_41520,N_41524);
nand U41778 (N_41778,N_41586,N_41543);
xor U41779 (N_41779,N_41680,N_41546);
and U41780 (N_41780,N_41626,N_41619);
xor U41781 (N_41781,N_41502,N_41678);
nand U41782 (N_41782,N_41603,N_41500);
or U41783 (N_41783,N_41707,N_41612);
xor U41784 (N_41784,N_41558,N_41740);
or U41785 (N_41785,N_41662,N_41660);
or U41786 (N_41786,N_41654,N_41531);
xnor U41787 (N_41787,N_41639,N_41514);
or U41788 (N_41788,N_41718,N_41671);
xor U41789 (N_41789,N_41627,N_41548);
and U41790 (N_41790,N_41592,N_41737);
xor U41791 (N_41791,N_41560,N_41597);
nor U41792 (N_41792,N_41600,N_41638);
or U41793 (N_41793,N_41529,N_41705);
and U41794 (N_41794,N_41615,N_41617);
and U41795 (N_41795,N_41741,N_41607);
and U41796 (N_41796,N_41604,N_41550);
and U41797 (N_41797,N_41656,N_41606);
xnor U41798 (N_41798,N_41724,N_41570);
and U41799 (N_41799,N_41566,N_41732);
nand U41800 (N_41800,N_41684,N_41650);
nor U41801 (N_41801,N_41698,N_41536);
xor U41802 (N_41802,N_41669,N_41693);
nor U41803 (N_41803,N_41645,N_41622);
or U41804 (N_41804,N_41552,N_41706);
or U41805 (N_41805,N_41578,N_41577);
nand U41806 (N_41806,N_41685,N_41519);
or U41807 (N_41807,N_41551,N_41691);
nand U41808 (N_41808,N_41667,N_41528);
or U41809 (N_41809,N_41509,N_41687);
xnor U41810 (N_41810,N_41708,N_41700);
nand U41811 (N_41811,N_41555,N_41508);
xnor U41812 (N_41812,N_41744,N_41631);
nor U41813 (N_41813,N_41664,N_41513);
or U41814 (N_41814,N_41637,N_41618);
xor U41815 (N_41815,N_41512,N_41714);
nor U41816 (N_41816,N_41697,N_41561);
and U41817 (N_41817,N_41711,N_41624);
nand U41818 (N_41818,N_41663,N_41571);
and U41819 (N_41819,N_41525,N_41712);
xor U41820 (N_41820,N_41719,N_41505);
and U41821 (N_41821,N_41688,N_41703);
or U41822 (N_41822,N_41657,N_41683);
nor U41823 (N_41823,N_41672,N_41557);
xnor U41824 (N_41824,N_41613,N_41564);
nor U41825 (N_41825,N_41575,N_41709);
xnor U41826 (N_41826,N_41629,N_41689);
nand U41827 (N_41827,N_41696,N_41676);
xor U41828 (N_41828,N_41504,N_41742);
nand U41829 (N_41829,N_41634,N_41665);
nand U41830 (N_41830,N_41730,N_41628);
nand U41831 (N_41831,N_41659,N_41673);
or U41832 (N_41832,N_41533,N_41544);
nor U41833 (N_41833,N_41515,N_41503);
and U41834 (N_41834,N_41630,N_41692);
nor U41835 (N_41835,N_41553,N_41644);
nor U41836 (N_41836,N_41728,N_41526);
nor U41837 (N_41837,N_41609,N_41545);
nand U41838 (N_41838,N_41694,N_41614);
nand U41839 (N_41839,N_41632,N_41704);
and U41840 (N_41840,N_41556,N_41648);
and U41841 (N_41841,N_41647,N_41542);
xnor U41842 (N_41842,N_41735,N_41661);
and U41843 (N_41843,N_41641,N_41723);
or U41844 (N_41844,N_41616,N_41534);
or U41845 (N_41845,N_41598,N_41507);
or U41846 (N_41846,N_41583,N_41679);
or U41847 (N_41847,N_41748,N_41655);
and U41848 (N_41848,N_41636,N_41580);
nand U41849 (N_41849,N_41605,N_41670);
xnor U41850 (N_41850,N_41653,N_41743);
xor U41851 (N_41851,N_41521,N_41733);
or U41852 (N_41852,N_41532,N_41530);
and U41853 (N_41853,N_41620,N_41535);
nand U41854 (N_41854,N_41541,N_41725);
or U41855 (N_41855,N_41633,N_41610);
nor U41856 (N_41856,N_41516,N_41537);
and U41857 (N_41857,N_41749,N_41658);
or U41858 (N_41858,N_41690,N_41646);
xnor U41859 (N_41859,N_41611,N_41726);
xor U41860 (N_41860,N_41640,N_41523);
nand U41861 (N_41861,N_41594,N_41608);
nor U41862 (N_41862,N_41721,N_41501);
or U41863 (N_41863,N_41554,N_41677);
and U41864 (N_41864,N_41675,N_41738);
and U41865 (N_41865,N_41701,N_41713);
nand U41866 (N_41866,N_41746,N_41538);
or U41867 (N_41867,N_41643,N_41666);
nand U41868 (N_41868,N_41747,N_41517);
nand U41869 (N_41869,N_41540,N_41625);
and U41870 (N_41870,N_41574,N_41562);
nand U41871 (N_41871,N_41522,N_41596);
nor U41872 (N_41872,N_41559,N_41635);
xnor U41873 (N_41873,N_41591,N_41717);
xnor U41874 (N_41874,N_41695,N_41595);
or U41875 (N_41875,N_41737,N_41608);
nand U41876 (N_41876,N_41681,N_41735);
and U41877 (N_41877,N_41630,N_41608);
nor U41878 (N_41878,N_41632,N_41720);
nand U41879 (N_41879,N_41629,N_41555);
or U41880 (N_41880,N_41685,N_41666);
and U41881 (N_41881,N_41559,N_41704);
nand U41882 (N_41882,N_41602,N_41701);
and U41883 (N_41883,N_41641,N_41529);
and U41884 (N_41884,N_41595,N_41628);
and U41885 (N_41885,N_41676,N_41559);
nand U41886 (N_41886,N_41642,N_41608);
and U41887 (N_41887,N_41555,N_41665);
nand U41888 (N_41888,N_41667,N_41658);
nor U41889 (N_41889,N_41624,N_41513);
nor U41890 (N_41890,N_41675,N_41720);
xnor U41891 (N_41891,N_41608,N_41619);
or U41892 (N_41892,N_41700,N_41734);
nand U41893 (N_41893,N_41712,N_41559);
xor U41894 (N_41894,N_41618,N_41724);
or U41895 (N_41895,N_41702,N_41576);
and U41896 (N_41896,N_41520,N_41601);
and U41897 (N_41897,N_41699,N_41513);
nor U41898 (N_41898,N_41572,N_41534);
xnor U41899 (N_41899,N_41703,N_41547);
or U41900 (N_41900,N_41523,N_41565);
xor U41901 (N_41901,N_41588,N_41737);
nor U41902 (N_41902,N_41609,N_41592);
xnor U41903 (N_41903,N_41516,N_41543);
nor U41904 (N_41904,N_41719,N_41624);
xnor U41905 (N_41905,N_41622,N_41516);
xor U41906 (N_41906,N_41714,N_41553);
or U41907 (N_41907,N_41638,N_41506);
and U41908 (N_41908,N_41677,N_41715);
xnor U41909 (N_41909,N_41535,N_41507);
and U41910 (N_41910,N_41537,N_41742);
nor U41911 (N_41911,N_41620,N_41630);
nor U41912 (N_41912,N_41730,N_41723);
and U41913 (N_41913,N_41577,N_41580);
xor U41914 (N_41914,N_41533,N_41736);
nand U41915 (N_41915,N_41554,N_41614);
nand U41916 (N_41916,N_41610,N_41738);
nand U41917 (N_41917,N_41719,N_41537);
and U41918 (N_41918,N_41613,N_41556);
xor U41919 (N_41919,N_41674,N_41564);
or U41920 (N_41920,N_41530,N_41560);
nand U41921 (N_41921,N_41682,N_41658);
or U41922 (N_41922,N_41593,N_41645);
nand U41923 (N_41923,N_41591,N_41531);
or U41924 (N_41924,N_41691,N_41661);
nand U41925 (N_41925,N_41529,N_41502);
nor U41926 (N_41926,N_41519,N_41619);
and U41927 (N_41927,N_41628,N_41551);
xnor U41928 (N_41928,N_41711,N_41513);
or U41929 (N_41929,N_41682,N_41642);
xnor U41930 (N_41930,N_41731,N_41521);
nor U41931 (N_41931,N_41658,N_41641);
and U41932 (N_41932,N_41608,N_41680);
nand U41933 (N_41933,N_41576,N_41705);
and U41934 (N_41934,N_41649,N_41573);
nor U41935 (N_41935,N_41700,N_41737);
and U41936 (N_41936,N_41613,N_41514);
or U41937 (N_41937,N_41613,N_41737);
or U41938 (N_41938,N_41643,N_41535);
or U41939 (N_41939,N_41626,N_41677);
nor U41940 (N_41940,N_41730,N_41671);
or U41941 (N_41941,N_41583,N_41667);
xor U41942 (N_41942,N_41550,N_41613);
nor U41943 (N_41943,N_41729,N_41646);
nand U41944 (N_41944,N_41681,N_41559);
xor U41945 (N_41945,N_41500,N_41572);
nand U41946 (N_41946,N_41698,N_41644);
or U41947 (N_41947,N_41635,N_41625);
and U41948 (N_41948,N_41602,N_41557);
xor U41949 (N_41949,N_41653,N_41665);
or U41950 (N_41950,N_41580,N_41536);
xor U41951 (N_41951,N_41565,N_41581);
nor U41952 (N_41952,N_41571,N_41513);
nand U41953 (N_41953,N_41719,N_41611);
nand U41954 (N_41954,N_41515,N_41525);
nor U41955 (N_41955,N_41653,N_41649);
nor U41956 (N_41956,N_41689,N_41627);
xnor U41957 (N_41957,N_41595,N_41607);
xor U41958 (N_41958,N_41546,N_41598);
and U41959 (N_41959,N_41667,N_41670);
nand U41960 (N_41960,N_41547,N_41655);
nand U41961 (N_41961,N_41630,N_41555);
and U41962 (N_41962,N_41560,N_41536);
and U41963 (N_41963,N_41695,N_41749);
xnor U41964 (N_41964,N_41745,N_41502);
and U41965 (N_41965,N_41704,N_41544);
or U41966 (N_41966,N_41690,N_41624);
and U41967 (N_41967,N_41569,N_41733);
or U41968 (N_41968,N_41506,N_41672);
nor U41969 (N_41969,N_41594,N_41711);
or U41970 (N_41970,N_41578,N_41687);
xnor U41971 (N_41971,N_41582,N_41643);
or U41972 (N_41972,N_41619,N_41656);
nor U41973 (N_41973,N_41682,N_41724);
nor U41974 (N_41974,N_41564,N_41704);
xnor U41975 (N_41975,N_41676,N_41630);
xor U41976 (N_41976,N_41674,N_41610);
or U41977 (N_41977,N_41678,N_41573);
and U41978 (N_41978,N_41735,N_41590);
nor U41979 (N_41979,N_41518,N_41582);
nand U41980 (N_41980,N_41647,N_41600);
or U41981 (N_41981,N_41724,N_41679);
xnor U41982 (N_41982,N_41641,N_41522);
and U41983 (N_41983,N_41518,N_41600);
xnor U41984 (N_41984,N_41743,N_41730);
nand U41985 (N_41985,N_41592,N_41586);
and U41986 (N_41986,N_41545,N_41728);
nor U41987 (N_41987,N_41747,N_41604);
or U41988 (N_41988,N_41539,N_41543);
nand U41989 (N_41989,N_41690,N_41665);
xnor U41990 (N_41990,N_41706,N_41646);
nor U41991 (N_41991,N_41536,N_41680);
nor U41992 (N_41992,N_41718,N_41670);
xor U41993 (N_41993,N_41634,N_41666);
and U41994 (N_41994,N_41526,N_41735);
or U41995 (N_41995,N_41611,N_41672);
xnor U41996 (N_41996,N_41742,N_41510);
or U41997 (N_41997,N_41557,N_41526);
nor U41998 (N_41998,N_41553,N_41626);
and U41999 (N_41999,N_41602,N_41509);
xor U42000 (N_42000,N_41838,N_41810);
and U42001 (N_42001,N_41762,N_41833);
nor U42002 (N_42002,N_41817,N_41843);
or U42003 (N_42003,N_41768,N_41904);
xnor U42004 (N_42004,N_41992,N_41806);
or U42005 (N_42005,N_41830,N_41976);
nand U42006 (N_42006,N_41805,N_41880);
nor U42007 (N_42007,N_41867,N_41807);
or U42008 (N_42008,N_41942,N_41798);
and U42009 (N_42009,N_41821,N_41900);
or U42010 (N_42010,N_41896,N_41832);
nor U42011 (N_42011,N_41950,N_41919);
nand U42012 (N_42012,N_41765,N_41921);
xnor U42013 (N_42013,N_41909,N_41908);
nand U42014 (N_42014,N_41887,N_41915);
and U42015 (N_42015,N_41794,N_41845);
nor U42016 (N_42016,N_41967,N_41878);
xor U42017 (N_42017,N_41923,N_41809);
nand U42018 (N_42018,N_41780,N_41871);
and U42019 (N_42019,N_41934,N_41836);
nor U42020 (N_42020,N_41866,N_41960);
and U42021 (N_42021,N_41927,N_41995);
and U42022 (N_42022,N_41757,N_41857);
nand U42023 (N_42023,N_41940,N_41802);
nand U42024 (N_42024,N_41947,N_41982);
nand U42025 (N_42025,N_41933,N_41846);
xnor U42026 (N_42026,N_41784,N_41943);
nor U42027 (N_42027,N_41876,N_41891);
and U42028 (N_42028,N_41793,N_41850);
or U42029 (N_42029,N_41906,N_41782);
xor U42030 (N_42030,N_41861,N_41791);
xnor U42031 (N_42031,N_41851,N_41929);
nor U42032 (N_42032,N_41955,N_41824);
and U42033 (N_42033,N_41898,N_41840);
nor U42034 (N_42034,N_41973,N_41983);
or U42035 (N_42035,N_41972,N_41886);
xnor U42036 (N_42036,N_41970,N_41882);
xnor U42037 (N_42037,N_41987,N_41977);
or U42038 (N_42038,N_41792,N_41756);
or U42039 (N_42039,N_41914,N_41892);
nand U42040 (N_42040,N_41881,N_41889);
xor U42041 (N_42041,N_41854,N_41874);
nand U42042 (N_42042,N_41812,N_41831);
nor U42043 (N_42043,N_41764,N_41860);
nor U42044 (N_42044,N_41789,N_41799);
and U42045 (N_42045,N_41924,N_41971);
or U42046 (N_42046,N_41922,N_41752);
or U42047 (N_42047,N_41758,N_41912);
nand U42048 (N_42048,N_41979,N_41875);
nor U42049 (N_42049,N_41964,N_41993);
xnor U42050 (N_42050,N_41763,N_41963);
nor U42051 (N_42051,N_41974,N_41829);
xnor U42052 (N_42052,N_41796,N_41902);
or U42053 (N_42053,N_41781,N_41968);
and U42054 (N_42054,N_41911,N_41823);
and U42055 (N_42055,N_41958,N_41913);
xor U42056 (N_42056,N_41839,N_41771);
or U42057 (N_42057,N_41869,N_41819);
and U42058 (N_42058,N_41897,N_41920);
nor U42059 (N_42059,N_41965,N_41849);
or U42060 (N_42060,N_41828,N_41885);
or U42061 (N_42061,N_41951,N_41939);
nor U42062 (N_42062,N_41872,N_41918);
and U42063 (N_42063,N_41759,N_41984);
or U42064 (N_42064,N_41842,N_41801);
nor U42065 (N_42065,N_41814,N_41766);
or U42066 (N_42066,N_41873,N_41755);
nor U42067 (N_42067,N_41883,N_41853);
and U42068 (N_42068,N_41835,N_41879);
or U42069 (N_42069,N_41855,N_41877);
nand U42070 (N_42070,N_41953,N_41868);
and U42071 (N_42071,N_41962,N_41848);
or U42072 (N_42072,N_41797,N_41774);
nor U42073 (N_42073,N_41926,N_41767);
xor U42074 (N_42074,N_41916,N_41994);
xor U42075 (N_42075,N_41773,N_41804);
or U42076 (N_42076,N_41808,N_41760);
nand U42077 (N_42077,N_41899,N_41952);
and U42078 (N_42078,N_41790,N_41859);
nand U42079 (N_42079,N_41856,N_41775);
or U42080 (N_42080,N_41910,N_41750);
nand U42081 (N_42081,N_41925,N_41863);
nor U42082 (N_42082,N_41811,N_41816);
or U42083 (N_42083,N_41841,N_41936);
xor U42084 (N_42084,N_41844,N_41815);
and U42085 (N_42085,N_41776,N_41803);
or U42086 (N_42086,N_41751,N_41788);
xor U42087 (N_42087,N_41905,N_41818);
nand U42088 (N_42088,N_41949,N_41864);
nand U42089 (N_42089,N_41787,N_41954);
and U42090 (N_42090,N_41884,N_41827);
nor U42091 (N_42091,N_41825,N_41944);
nand U42092 (N_42092,N_41800,N_41989);
and U42093 (N_42093,N_41761,N_41837);
nand U42094 (N_42094,N_41938,N_41937);
nand U42095 (N_42095,N_41903,N_41858);
xor U42096 (N_42096,N_41893,N_41945);
xor U42097 (N_42097,N_41961,N_41998);
or U42098 (N_42098,N_41888,N_41847);
nand U42099 (N_42099,N_41770,N_41895);
nor U42100 (N_42100,N_41820,N_41978);
xor U42101 (N_42101,N_41997,N_41957);
xnor U42102 (N_42102,N_41772,N_41822);
nand U42103 (N_42103,N_41931,N_41990);
xor U42104 (N_42104,N_41779,N_41907);
and U42105 (N_42105,N_41980,N_41826);
xor U42106 (N_42106,N_41930,N_41991);
nor U42107 (N_42107,N_41941,N_41852);
or U42108 (N_42108,N_41865,N_41988);
xnor U42109 (N_42109,N_41917,N_41928);
or U42110 (N_42110,N_41777,N_41981);
nand U42111 (N_42111,N_41996,N_41948);
nand U42112 (N_42112,N_41946,N_41890);
nor U42113 (N_42113,N_41769,N_41862);
and U42114 (N_42114,N_41966,N_41894);
nand U42115 (N_42115,N_41999,N_41986);
and U42116 (N_42116,N_41969,N_41834);
nor U42117 (N_42117,N_41901,N_41795);
or U42118 (N_42118,N_41783,N_41956);
or U42119 (N_42119,N_41932,N_41870);
nor U42120 (N_42120,N_41778,N_41754);
or U42121 (N_42121,N_41985,N_41786);
or U42122 (N_42122,N_41935,N_41959);
or U42123 (N_42123,N_41753,N_41785);
and U42124 (N_42124,N_41813,N_41975);
xnor U42125 (N_42125,N_41863,N_41905);
and U42126 (N_42126,N_41850,N_41916);
nand U42127 (N_42127,N_41859,N_41807);
xnor U42128 (N_42128,N_41964,N_41872);
nand U42129 (N_42129,N_41948,N_41868);
xnor U42130 (N_42130,N_41916,N_41886);
nor U42131 (N_42131,N_41873,N_41917);
xor U42132 (N_42132,N_41983,N_41764);
and U42133 (N_42133,N_41983,N_41879);
nand U42134 (N_42134,N_41834,N_41802);
nor U42135 (N_42135,N_41818,N_41959);
xor U42136 (N_42136,N_41804,N_41757);
nand U42137 (N_42137,N_41927,N_41810);
nand U42138 (N_42138,N_41931,N_41982);
or U42139 (N_42139,N_41971,N_41927);
or U42140 (N_42140,N_41960,N_41843);
nor U42141 (N_42141,N_41762,N_41962);
or U42142 (N_42142,N_41929,N_41967);
and U42143 (N_42143,N_41900,N_41978);
and U42144 (N_42144,N_41974,N_41907);
nand U42145 (N_42145,N_41780,N_41867);
or U42146 (N_42146,N_41812,N_41818);
nand U42147 (N_42147,N_41792,N_41804);
nor U42148 (N_42148,N_41773,N_41815);
or U42149 (N_42149,N_41887,N_41820);
and U42150 (N_42150,N_41833,N_41785);
or U42151 (N_42151,N_41904,N_41908);
and U42152 (N_42152,N_41860,N_41847);
xnor U42153 (N_42153,N_41981,N_41954);
and U42154 (N_42154,N_41926,N_41909);
and U42155 (N_42155,N_41980,N_41931);
nand U42156 (N_42156,N_41939,N_41907);
nor U42157 (N_42157,N_41931,N_41965);
xnor U42158 (N_42158,N_41947,N_41793);
xnor U42159 (N_42159,N_41794,N_41859);
nand U42160 (N_42160,N_41891,N_41930);
and U42161 (N_42161,N_41839,N_41834);
xnor U42162 (N_42162,N_41953,N_41753);
xnor U42163 (N_42163,N_41798,N_41823);
and U42164 (N_42164,N_41956,N_41766);
xor U42165 (N_42165,N_41789,N_41845);
xor U42166 (N_42166,N_41791,N_41774);
nand U42167 (N_42167,N_41816,N_41847);
or U42168 (N_42168,N_41903,N_41874);
nor U42169 (N_42169,N_41772,N_41922);
nand U42170 (N_42170,N_41927,N_41957);
and U42171 (N_42171,N_41888,N_41910);
xor U42172 (N_42172,N_41794,N_41788);
or U42173 (N_42173,N_41996,N_41946);
and U42174 (N_42174,N_41803,N_41777);
and U42175 (N_42175,N_41763,N_41891);
nor U42176 (N_42176,N_41765,N_41769);
xnor U42177 (N_42177,N_41918,N_41764);
or U42178 (N_42178,N_41958,N_41851);
nor U42179 (N_42179,N_41845,N_41886);
or U42180 (N_42180,N_41837,N_41869);
or U42181 (N_42181,N_41926,N_41805);
or U42182 (N_42182,N_41978,N_41919);
nand U42183 (N_42183,N_41810,N_41859);
or U42184 (N_42184,N_41817,N_41902);
nand U42185 (N_42185,N_41899,N_41857);
nand U42186 (N_42186,N_41827,N_41833);
and U42187 (N_42187,N_41872,N_41897);
nor U42188 (N_42188,N_41787,N_41783);
or U42189 (N_42189,N_41803,N_41888);
or U42190 (N_42190,N_41984,N_41926);
nor U42191 (N_42191,N_41810,N_41857);
and U42192 (N_42192,N_41847,N_41981);
xnor U42193 (N_42193,N_41816,N_41892);
nor U42194 (N_42194,N_41887,N_41826);
xor U42195 (N_42195,N_41955,N_41946);
and U42196 (N_42196,N_41809,N_41799);
and U42197 (N_42197,N_41804,N_41866);
nor U42198 (N_42198,N_41994,N_41949);
or U42199 (N_42199,N_41963,N_41754);
nor U42200 (N_42200,N_41807,N_41965);
nor U42201 (N_42201,N_41937,N_41923);
nand U42202 (N_42202,N_41962,N_41965);
nor U42203 (N_42203,N_41864,N_41876);
xnor U42204 (N_42204,N_41902,N_41770);
nor U42205 (N_42205,N_41829,N_41758);
nor U42206 (N_42206,N_41751,N_41874);
xnor U42207 (N_42207,N_41767,N_41810);
nand U42208 (N_42208,N_41857,N_41914);
nand U42209 (N_42209,N_41799,N_41760);
xor U42210 (N_42210,N_41954,N_41779);
nand U42211 (N_42211,N_41948,N_41786);
and U42212 (N_42212,N_41790,N_41829);
or U42213 (N_42213,N_41912,N_41923);
xnor U42214 (N_42214,N_41987,N_41860);
or U42215 (N_42215,N_41907,N_41906);
nand U42216 (N_42216,N_41845,N_41853);
nand U42217 (N_42217,N_41959,N_41980);
nor U42218 (N_42218,N_41782,N_41795);
nor U42219 (N_42219,N_41927,N_41949);
nor U42220 (N_42220,N_41804,N_41919);
xnor U42221 (N_42221,N_41905,N_41791);
nor U42222 (N_42222,N_41962,N_41799);
and U42223 (N_42223,N_41800,N_41856);
and U42224 (N_42224,N_41863,N_41782);
and U42225 (N_42225,N_41890,N_41789);
nand U42226 (N_42226,N_41824,N_41766);
xnor U42227 (N_42227,N_41966,N_41887);
xor U42228 (N_42228,N_41802,N_41874);
xor U42229 (N_42229,N_41904,N_41920);
and U42230 (N_42230,N_41953,N_41818);
nor U42231 (N_42231,N_41910,N_41872);
or U42232 (N_42232,N_41753,N_41985);
nor U42233 (N_42233,N_41804,N_41966);
xnor U42234 (N_42234,N_41823,N_41917);
nand U42235 (N_42235,N_41812,N_41842);
xor U42236 (N_42236,N_41899,N_41901);
nand U42237 (N_42237,N_41958,N_41945);
and U42238 (N_42238,N_41765,N_41822);
nand U42239 (N_42239,N_41850,N_41832);
xnor U42240 (N_42240,N_41892,N_41933);
nand U42241 (N_42241,N_41877,N_41764);
nor U42242 (N_42242,N_41890,N_41850);
nand U42243 (N_42243,N_41999,N_41913);
or U42244 (N_42244,N_41904,N_41854);
and U42245 (N_42245,N_41915,N_41932);
and U42246 (N_42246,N_41826,N_41817);
nor U42247 (N_42247,N_41867,N_41763);
xor U42248 (N_42248,N_41821,N_41843);
xnor U42249 (N_42249,N_41898,N_41792);
nor U42250 (N_42250,N_42105,N_42045);
and U42251 (N_42251,N_42116,N_42174);
and U42252 (N_42252,N_42048,N_42097);
nor U42253 (N_42253,N_42099,N_42149);
xor U42254 (N_42254,N_42132,N_42220);
and U42255 (N_42255,N_42101,N_42061);
or U42256 (N_42256,N_42203,N_42021);
and U42257 (N_42257,N_42166,N_42169);
nor U42258 (N_42258,N_42131,N_42109);
and U42259 (N_42259,N_42197,N_42148);
nand U42260 (N_42260,N_42137,N_42065);
nor U42261 (N_42261,N_42163,N_42243);
and U42262 (N_42262,N_42117,N_42240);
and U42263 (N_42263,N_42112,N_42079);
nand U42264 (N_42264,N_42219,N_42086);
and U42265 (N_42265,N_42059,N_42182);
or U42266 (N_42266,N_42234,N_42189);
and U42267 (N_42267,N_42184,N_42227);
and U42268 (N_42268,N_42248,N_42145);
and U42269 (N_42269,N_42183,N_42102);
or U42270 (N_42270,N_42129,N_42010);
and U42271 (N_42271,N_42047,N_42110);
nand U42272 (N_42272,N_42027,N_42091);
or U42273 (N_42273,N_42067,N_42249);
xnor U42274 (N_42274,N_42009,N_42000);
xor U42275 (N_42275,N_42073,N_42108);
nor U42276 (N_42276,N_42039,N_42224);
xor U42277 (N_42277,N_42090,N_42029);
or U42278 (N_42278,N_42007,N_42168);
nor U42279 (N_42279,N_42094,N_42126);
xor U42280 (N_42280,N_42239,N_42153);
nor U42281 (N_42281,N_42241,N_42164);
nor U42282 (N_42282,N_42012,N_42150);
and U42283 (N_42283,N_42225,N_42171);
nand U42284 (N_42284,N_42071,N_42074);
and U42285 (N_42285,N_42032,N_42081);
nor U42286 (N_42286,N_42089,N_42207);
nand U42287 (N_42287,N_42191,N_42121);
xor U42288 (N_42288,N_42188,N_42209);
nand U42289 (N_42289,N_42177,N_42179);
and U42290 (N_42290,N_42068,N_42066);
or U42291 (N_42291,N_42172,N_42026);
nand U42292 (N_42292,N_42111,N_42057);
nand U42293 (N_42293,N_42056,N_42165);
nand U42294 (N_42294,N_42043,N_42155);
or U42295 (N_42295,N_42192,N_42142);
nor U42296 (N_42296,N_42022,N_42141);
and U42297 (N_42297,N_42233,N_42018);
nand U42298 (N_42298,N_42175,N_42005);
nor U42299 (N_42299,N_42031,N_42167);
and U42300 (N_42300,N_42223,N_42104);
and U42301 (N_42301,N_42041,N_42136);
nand U42302 (N_42302,N_42024,N_42014);
or U42303 (N_42303,N_42001,N_42211);
and U42304 (N_42304,N_42213,N_42135);
xnor U42305 (N_42305,N_42247,N_42127);
nor U42306 (N_42306,N_42013,N_42162);
or U42307 (N_42307,N_42038,N_42204);
nand U42308 (N_42308,N_42198,N_42237);
and U42309 (N_42309,N_42152,N_42100);
and U42310 (N_42310,N_42200,N_42222);
and U42311 (N_42311,N_42106,N_42082);
nand U42312 (N_42312,N_42186,N_42020);
nand U42313 (N_42313,N_42178,N_42064);
nor U42314 (N_42314,N_42235,N_42160);
nand U42315 (N_42315,N_42226,N_42113);
nor U42316 (N_42316,N_42208,N_42040);
and U42317 (N_42317,N_42015,N_42103);
or U42318 (N_42318,N_42072,N_42212);
and U42319 (N_42319,N_42122,N_42130);
or U42320 (N_42320,N_42221,N_42202);
xor U42321 (N_42321,N_42170,N_42217);
nand U42322 (N_42322,N_42232,N_42033);
and U42323 (N_42323,N_42181,N_42125);
xnor U42324 (N_42324,N_42210,N_42035);
nand U42325 (N_42325,N_42087,N_42143);
nand U42326 (N_42326,N_42036,N_42078);
xnor U42327 (N_42327,N_42025,N_42119);
or U42328 (N_42328,N_42216,N_42236);
xor U42329 (N_42329,N_42205,N_42124);
xor U42330 (N_42330,N_42214,N_42008);
or U42331 (N_42331,N_42176,N_42004);
or U42332 (N_42332,N_42157,N_42229);
nand U42333 (N_42333,N_42049,N_42120);
or U42334 (N_42334,N_42156,N_42096);
nor U42335 (N_42335,N_42083,N_42238);
or U42336 (N_42336,N_42070,N_42173);
nand U42337 (N_42337,N_42201,N_42140);
nor U42338 (N_42338,N_42093,N_42123);
xnor U42339 (N_42339,N_42054,N_42196);
xor U42340 (N_42340,N_42158,N_42060);
and U42341 (N_42341,N_42146,N_42244);
or U42342 (N_42342,N_42051,N_42134);
xor U42343 (N_42343,N_42088,N_42128);
nor U42344 (N_42344,N_42062,N_42245);
or U42345 (N_42345,N_42242,N_42114);
xor U42346 (N_42346,N_42095,N_42115);
nor U42347 (N_42347,N_42076,N_42080);
nor U42348 (N_42348,N_42159,N_42180);
and U42349 (N_42349,N_42199,N_42075);
and U42350 (N_42350,N_42006,N_42053);
and U42351 (N_42351,N_42194,N_42042);
nor U42352 (N_42352,N_42046,N_42228);
and U42353 (N_42353,N_42023,N_42133);
nand U42354 (N_42354,N_42003,N_42193);
or U42355 (N_42355,N_42077,N_42085);
nand U42356 (N_42356,N_42037,N_42139);
nand U42357 (N_42357,N_42019,N_42055);
nand U42358 (N_42358,N_42069,N_42187);
or U42359 (N_42359,N_42098,N_42092);
and U42360 (N_42360,N_42063,N_42058);
or U42361 (N_42361,N_42215,N_42034);
nor U42362 (N_42362,N_42195,N_42002);
xnor U42363 (N_42363,N_42050,N_42147);
and U42364 (N_42364,N_42044,N_42016);
xor U42365 (N_42365,N_42028,N_42118);
or U42366 (N_42366,N_42246,N_42144);
and U42367 (N_42367,N_42017,N_42231);
xor U42368 (N_42368,N_42011,N_42206);
nand U42369 (N_42369,N_42218,N_42138);
and U42370 (N_42370,N_42185,N_42084);
and U42371 (N_42371,N_42230,N_42052);
nor U42372 (N_42372,N_42030,N_42154);
xor U42373 (N_42373,N_42151,N_42161);
nor U42374 (N_42374,N_42107,N_42190);
or U42375 (N_42375,N_42103,N_42156);
or U42376 (N_42376,N_42113,N_42157);
nor U42377 (N_42377,N_42080,N_42023);
nand U42378 (N_42378,N_42145,N_42007);
nor U42379 (N_42379,N_42070,N_42163);
and U42380 (N_42380,N_42119,N_42029);
xnor U42381 (N_42381,N_42037,N_42091);
nor U42382 (N_42382,N_42130,N_42249);
and U42383 (N_42383,N_42109,N_42203);
xnor U42384 (N_42384,N_42018,N_42110);
and U42385 (N_42385,N_42012,N_42237);
nor U42386 (N_42386,N_42221,N_42035);
nor U42387 (N_42387,N_42113,N_42090);
xnor U42388 (N_42388,N_42240,N_42224);
or U42389 (N_42389,N_42053,N_42008);
xnor U42390 (N_42390,N_42197,N_42245);
xnor U42391 (N_42391,N_42069,N_42132);
nor U42392 (N_42392,N_42173,N_42149);
xnor U42393 (N_42393,N_42058,N_42057);
or U42394 (N_42394,N_42186,N_42071);
and U42395 (N_42395,N_42070,N_42199);
or U42396 (N_42396,N_42097,N_42196);
and U42397 (N_42397,N_42136,N_42004);
xor U42398 (N_42398,N_42116,N_42196);
and U42399 (N_42399,N_42136,N_42044);
nand U42400 (N_42400,N_42040,N_42226);
nor U42401 (N_42401,N_42114,N_42135);
and U42402 (N_42402,N_42170,N_42245);
nor U42403 (N_42403,N_42040,N_42117);
or U42404 (N_42404,N_42168,N_42043);
nor U42405 (N_42405,N_42017,N_42123);
and U42406 (N_42406,N_42183,N_42155);
nand U42407 (N_42407,N_42129,N_42038);
xor U42408 (N_42408,N_42237,N_42051);
nand U42409 (N_42409,N_42014,N_42206);
and U42410 (N_42410,N_42020,N_42113);
xor U42411 (N_42411,N_42154,N_42111);
xnor U42412 (N_42412,N_42041,N_42073);
or U42413 (N_42413,N_42049,N_42116);
and U42414 (N_42414,N_42057,N_42122);
nand U42415 (N_42415,N_42112,N_42205);
nor U42416 (N_42416,N_42150,N_42157);
and U42417 (N_42417,N_42132,N_42231);
xnor U42418 (N_42418,N_42072,N_42137);
nor U42419 (N_42419,N_42108,N_42136);
or U42420 (N_42420,N_42151,N_42023);
xor U42421 (N_42421,N_42199,N_42060);
xnor U42422 (N_42422,N_42173,N_42007);
or U42423 (N_42423,N_42116,N_42245);
and U42424 (N_42424,N_42062,N_42016);
or U42425 (N_42425,N_42126,N_42015);
nor U42426 (N_42426,N_42055,N_42036);
and U42427 (N_42427,N_42156,N_42141);
or U42428 (N_42428,N_42095,N_42120);
or U42429 (N_42429,N_42246,N_42061);
or U42430 (N_42430,N_42247,N_42058);
and U42431 (N_42431,N_42125,N_42154);
or U42432 (N_42432,N_42181,N_42179);
nand U42433 (N_42433,N_42081,N_42066);
nor U42434 (N_42434,N_42053,N_42242);
nor U42435 (N_42435,N_42130,N_42107);
xor U42436 (N_42436,N_42245,N_42076);
or U42437 (N_42437,N_42071,N_42170);
or U42438 (N_42438,N_42006,N_42062);
nand U42439 (N_42439,N_42077,N_42060);
xnor U42440 (N_42440,N_42074,N_42225);
or U42441 (N_42441,N_42198,N_42112);
nand U42442 (N_42442,N_42169,N_42039);
or U42443 (N_42443,N_42188,N_42116);
xor U42444 (N_42444,N_42032,N_42092);
nor U42445 (N_42445,N_42236,N_42168);
nand U42446 (N_42446,N_42080,N_42008);
nand U42447 (N_42447,N_42233,N_42092);
xor U42448 (N_42448,N_42078,N_42165);
nand U42449 (N_42449,N_42204,N_42217);
nor U42450 (N_42450,N_42214,N_42141);
nand U42451 (N_42451,N_42030,N_42148);
nor U42452 (N_42452,N_42014,N_42025);
xor U42453 (N_42453,N_42192,N_42176);
nand U42454 (N_42454,N_42178,N_42236);
nand U42455 (N_42455,N_42075,N_42232);
nand U42456 (N_42456,N_42137,N_42091);
and U42457 (N_42457,N_42087,N_42224);
and U42458 (N_42458,N_42030,N_42135);
nor U42459 (N_42459,N_42122,N_42217);
and U42460 (N_42460,N_42119,N_42071);
nor U42461 (N_42461,N_42158,N_42020);
xor U42462 (N_42462,N_42179,N_42187);
nand U42463 (N_42463,N_42215,N_42221);
nor U42464 (N_42464,N_42063,N_42011);
and U42465 (N_42465,N_42234,N_42175);
xor U42466 (N_42466,N_42243,N_42199);
nand U42467 (N_42467,N_42175,N_42184);
xor U42468 (N_42468,N_42222,N_42013);
xor U42469 (N_42469,N_42023,N_42128);
xor U42470 (N_42470,N_42046,N_42163);
and U42471 (N_42471,N_42146,N_42215);
and U42472 (N_42472,N_42038,N_42225);
nand U42473 (N_42473,N_42157,N_42061);
and U42474 (N_42474,N_42057,N_42175);
nand U42475 (N_42475,N_42108,N_42175);
nor U42476 (N_42476,N_42081,N_42072);
and U42477 (N_42477,N_42037,N_42161);
nand U42478 (N_42478,N_42039,N_42165);
xnor U42479 (N_42479,N_42113,N_42025);
nor U42480 (N_42480,N_42005,N_42043);
nand U42481 (N_42481,N_42186,N_42090);
nand U42482 (N_42482,N_42053,N_42195);
nand U42483 (N_42483,N_42146,N_42204);
and U42484 (N_42484,N_42146,N_42156);
nor U42485 (N_42485,N_42178,N_42078);
or U42486 (N_42486,N_42102,N_42018);
xnor U42487 (N_42487,N_42154,N_42020);
nor U42488 (N_42488,N_42001,N_42037);
and U42489 (N_42489,N_42241,N_42041);
nor U42490 (N_42490,N_42074,N_42096);
or U42491 (N_42491,N_42169,N_42015);
nand U42492 (N_42492,N_42087,N_42078);
xnor U42493 (N_42493,N_42240,N_42215);
and U42494 (N_42494,N_42228,N_42195);
xor U42495 (N_42495,N_42098,N_42119);
xor U42496 (N_42496,N_42001,N_42091);
and U42497 (N_42497,N_42116,N_42249);
nor U42498 (N_42498,N_42108,N_42052);
xor U42499 (N_42499,N_42216,N_42105);
and U42500 (N_42500,N_42480,N_42273);
or U42501 (N_42501,N_42255,N_42265);
and U42502 (N_42502,N_42397,N_42463);
nand U42503 (N_42503,N_42268,N_42444);
xor U42504 (N_42504,N_42317,N_42366);
nand U42505 (N_42505,N_42393,N_42484);
and U42506 (N_42506,N_42426,N_42263);
nor U42507 (N_42507,N_42460,N_42304);
xnor U42508 (N_42508,N_42462,N_42392);
xnor U42509 (N_42509,N_42468,N_42459);
nand U42510 (N_42510,N_42455,N_42274);
xnor U42511 (N_42511,N_42272,N_42422);
xor U42512 (N_42512,N_42355,N_42311);
nand U42513 (N_42513,N_42436,N_42325);
nor U42514 (N_42514,N_42312,N_42271);
and U42515 (N_42515,N_42405,N_42281);
xnor U42516 (N_42516,N_42384,N_42417);
xnor U42517 (N_42517,N_42406,N_42486);
xnor U42518 (N_42518,N_42357,N_42293);
nor U42519 (N_42519,N_42280,N_42286);
or U42520 (N_42520,N_42418,N_42431);
xor U42521 (N_42521,N_42421,N_42490);
and U42522 (N_42522,N_42439,N_42471);
nand U42523 (N_42523,N_42424,N_42327);
or U42524 (N_42524,N_42491,N_42361);
nand U42525 (N_42525,N_42448,N_42446);
xor U42526 (N_42526,N_42469,N_42302);
xor U42527 (N_42527,N_42282,N_42340);
nor U42528 (N_42528,N_42498,N_42332);
or U42529 (N_42529,N_42430,N_42464);
xor U42530 (N_42530,N_42432,N_42483);
or U42531 (N_42531,N_42359,N_42339);
xor U42532 (N_42532,N_42306,N_42258);
xnor U42533 (N_42533,N_42305,N_42434);
nand U42534 (N_42534,N_42379,N_42370);
nand U42535 (N_42535,N_42398,N_42334);
nand U42536 (N_42536,N_42453,N_42475);
or U42537 (N_42537,N_42308,N_42287);
nand U42538 (N_42538,N_42298,N_42284);
and U42539 (N_42539,N_42380,N_42467);
nor U42540 (N_42540,N_42289,N_42363);
nand U42541 (N_42541,N_42451,N_42429);
or U42542 (N_42542,N_42252,N_42378);
nand U42543 (N_42543,N_42326,N_42269);
nand U42544 (N_42544,N_42409,N_42313);
or U42545 (N_42545,N_42369,N_42320);
nor U42546 (N_42546,N_42300,N_42416);
and U42547 (N_42547,N_42443,N_42254);
xor U42548 (N_42548,N_42343,N_42351);
xor U42549 (N_42549,N_42388,N_42368);
xnor U42550 (N_42550,N_42387,N_42495);
nand U42551 (N_42551,N_42497,N_42479);
and U42552 (N_42552,N_42331,N_42303);
or U42553 (N_42553,N_42425,N_42295);
and U42554 (N_42554,N_42465,N_42382);
nor U42555 (N_42555,N_42261,N_42266);
and U42556 (N_42556,N_42437,N_42347);
xor U42557 (N_42557,N_42279,N_42338);
nand U42558 (N_42558,N_42333,N_42410);
nand U42559 (N_42559,N_42374,N_42315);
and U42560 (N_42560,N_42461,N_42458);
and U42561 (N_42561,N_42396,N_42411);
nor U42562 (N_42562,N_42401,N_42442);
xor U42563 (N_42563,N_42276,N_42342);
xor U42564 (N_42564,N_42358,N_42404);
xnor U42565 (N_42565,N_42264,N_42403);
or U42566 (N_42566,N_42447,N_42385);
or U42567 (N_42567,N_42481,N_42435);
nand U42568 (N_42568,N_42419,N_42323);
nor U42569 (N_42569,N_42292,N_42466);
nand U42570 (N_42570,N_42440,N_42329);
xor U42571 (N_42571,N_42307,N_42354);
nand U42572 (N_42572,N_42309,N_42341);
xnor U42573 (N_42573,N_42297,N_42407);
nand U42574 (N_42574,N_42413,N_42456);
or U42575 (N_42575,N_42372,N_42399);
and U42576 (N_42576,N_42260,N_42324);
and U42577 (N_42577,N_42328,N_42400);
xor U42578 (N_42578,N_42394,N_42408);
nand U42579 (N_42579,N_42485,N_42414);
nor U42580 (N_42580,N_42473,N_42322);
xnor U42581 (N_42581,N_42253,N_42415);
nand U42582 (N_42582,N_42373,N_42412);
and U42583 (N_42583,N_42344,N_42262);
xnor U42584 (N_42584,N_42499,N_42299);
or U42585 (N_42585,N_42376,N_42275);
nand U42586 (N_42586,N_42375,N_42423);
nand U42587 (N_42587,N_42310,N_42395);
and U42588 (N_42588,N_42428,N_42420);
xnor U42589 (N_42589,N_42301,N_42350);
nor U42590 (N_42590,N_42478,N_42438);
nor U42591 (N_42591,N_42348,N_42335);
xor U42592 (N_42592,N_42492,N_42296);
nand U42593 (N_42593,N_42318,N_42345);
xor U42594 (N_42594,N_42285,N_42474);
xnor U42595 (N_42595,N_42336,N_42433);
or U42596 (N_42596,N_42476,N_42250);
and U42597 (N_42597,N_42470,N_42267);
xnor U42598 (N_42598,N_42494,N_42441);
or U42599 (N_42599,N_42251,N_42450);
and U42600 (N_42600,N_42457,N_42314);
and U42601 (N_42601,N_42371,N_42477);
nor U42602 (N_42602,N_42283,N_42386);
xor U42603 (N_42603,N_42445,N_42488);
nand U42604 (N_42604,N_42482,N_42294);
and U42605 (N_42605,N_42330,N_42493);
or U42606 (N_42606,N_42391,N_42365);
or U42607 (N_42607,N_42349,N_42390);
nor U42608 (N_42608,N_42383,N_42256);
nand U42609 (N_42609,N_42316,N_42270);
and U42610 (N_42610,N_42291,N_42321);
nand U42611 (N_42611,N_42472,N_42364);
or U42612 (N_42612,N_42449,N_42337);
and U42613 (N_42613,N_42352,N_42389);
nand U42614 (N_42614,N_42259,N_42381);
and U42615 (N_42615,N_42360,N_42452);
or U42616 (N_42616,N_42353,N_42288);
nor U42617 (N_42617,N_42487,N_42377);
and U42618 (N_42618,N_42427,N_42362);
and U42619 (N_42619,N_42346,N_42290);
or U42620 (N_42620,N_42356,N_42367);
xor U42621 (N_42621,N_42257,N_42489);
or U42622 (N_42622,N_42402,N_42277);
nor U42623 (N_42623,N_42496,N_42454);
nor U42624 (N_42624,N_42278,N_42319);
and U42625 (N_42625,N_42380,N_42484);
or U42626 (N_42626,N_42393,N_42250);
nand U42627 (N_42627,N_42315,N_42324);
xnor U42628 (N_42628,N_42319,N_42253);
nand U42629 (N_42629,N_42284,N_42413);
and U42630 (N_42630,N_42372,N_42371);
xor U42631 (N_42631,N_42278,N_42307);
or U42632 (N_42632,N_42450,N_42274);
or U42633 (N_42633,N_42364,N_42306);
xnor U42634 (N_42634,N_42385,N_42289);
nand U42635 (N_42635,N_42305,N_42321);
nor U42636 (N_42636,N_42443,N_42275);
or U42637 (N_42637,N_42471,N_42425);
xor U42638 (N_42638,N_42261,N_42443);
and U42639 (N_42639,N_42397,N_42457);
or U42640 (N_42640,N_42254,N_42282);
or U42641 (N_42641,N_42294,N_42439);
nor U42642 (N_42642,N_42283,N_42307);
nand U42643 (N_42643,N_42408,N_42312);
nand U42644 (N_42644,N_42356,N_42438);
xnor U42645 (N_42645,N_42438,N_42467);
and U42646 (N_42646,N_42306,N_42478);
and U42647 (N_42647,N_42485,N_42279);
nand U42648 (N_42648,N_42451,N_42325);
xnor U42649 (N_42649,N_42362,N_42252);
nand U42650 (N_42650,N_42486,N_42485);
nand U42651 (N_42651,N_42438,N_42348);
xor U42652 (N_42652,N_42347,N_42407);
or U42653 (N_42653,N_42334,N_42340);
xor U42654 (N_42654,N_42345,N_42416);
xor U42655 (N_42655,N_42282,N_42461);
xor U42656 (N_42656,N_42435,N_42334);
and U42657 (N_42657,N_42340,N_42377);
and U42658 (N_42658,N_42323,N_42312);
or U42659 (N_42659,N_42258,N_42427);
or U42660 (N_42660,N_42451,N_42399);
or U42661 (N_42661,N_42323,N_42376);
or U42662 (N_42662,N_42493,N_42260);
nand U42663 (N_42663,N_42267,N_42336);
nand U42664 (N_42664,N_42345,N_42268);
nor U42665 (N_42665,N_42278,N_42266);
xor U42666 (N_42666,N_42308,N_42343);
nor U42667 (N_42667,N_42393,N_42303);
nor U42668 (N_42668,N_42337,N_42474);
or U42669 (N_42669,N_42444,N_42265);
xor U42670 (N_42670,N_42296,N_42314);
nor U42671 (N_42671,N_42451,N_42446);
or U42672 (N_42672,N_42359,N_42430);
and U42673 (N_42673,N_42288,N_42387);
nor U42674 (N_42674,N_42276,N_42405);
or U42675 (N_42675,N_42399,N_42405);
or U42676 (N_42676,N_42483,N_42291);
nand U42677 (N_42677,N_42278,N_42431);
xor U42678 (N_42678,N_42279,N_42256);
nor U42679 (N_42679,N_42305,N_42287);
nor U42680 (N_42680,N_42446,N_42278);
xor U42681 (N_42681,N_42405,N_42307);
and U42682 (N_42682,N_42391,N_42486);
and U42683 (N_42683,N_42338,N_42460);
or U42684 (N_42684,N_42363,N_42381);
nand U42685 (N_42685,N_42457,N_42448);
nor U42686 (N_42686,N_42425,N_42419);
nand U42687 (N_42687,N_42341,N_42464);
or U42688 (N_42688,N_42332,N_42281);
and U42689 (N_42689,N_42395,N_42334);
and U42690 (N_42690,N_42425,N_42276);
xor U42691 (N_42691,N_42385,N_42270);
or U42692 (N_42692,N_42263,N_42364);
nor U42693 (N_42693,N_42397,N_42455);
xnor U42694 (N_42694,N_42274,N_42427);
xnor U42695 (N_42695,N_42253,N_42348);
nand U42696 (N_42696,N_42303,N_42313);
nand U42697 (N_42697,N_42489,N_42331);
nand U42698 (N_42698,N_42479,N_42322);
and U42699 (N_42699,N_42491,N_42362);
nand U42700 (N_42700,N_42489,N_42314);
and U42701 (N_42701,N_42323,N_42382);
or U42702 (N_42702,N_42475,N_42370);
and U42703 (N_42703,N_42336,N_42328);
or U42704 (N_42704,N_42420,N_42289);
and U42705 (N_42705,N_42397,N_42298);
nand U42706 (N_42706,N_42431,N_42474);
nor U42707 (N_42707,N_42329,N_42441);
nor U42708 (N_42708,N_42404,N_42357);
nor U42709 (N_42709,N_42267,N_42271);
or U42710 (N_42710,N_42348,N_42409);
xnor U42711 (N_42711,N_42331,N_42266);
xnor U42712 (N_42712,N_42389,N_42318);
xor U42713 (N_42713,N_42442,N_42287);
nor U42714 (N_42714,N_42482,N_42290);
nand U42715 (N_42715,N_42299,N_42429);
nand U42716 (N_42716,N_42330,N_42425);
xnor U42717 (N_42717,N_42487,N_42264);
nor U42718 (N_42718,N_42348,N_42364);
nor U42719 (N_42719,N_42304,N_42415);
nor U42720 (N_42720,N_42427,N_42316);
and U42721 (N_42721,N_42429,N_42253);
or U42722 (N_42722,N_42395,N_42385);
nand U42723 (N_42723,N_42400,N_42358);
or U42724 (N_42724,N_42447,N_42295);
or U42725 (N_42725,N_42426,N_42463);
or U42726 (N_42726,N_42463,N_42303);
xor U42727 (N_42727,N_42463,N_42411);
xor U42728 (N_42728,N_42302,N_42353);
xnor U42729 (N_42729,N_42436,N_42355);
xnor U42730 (N_42730,N_42390,N_42287);
xor U42731 (N_42731,N_42283,N_42348);
and U42732 (N_42732,N_42360,N_42448);
or U42733 (N_42733,N_42271,N_42323);
and U42734 (N_42734,N_42315,N_42466);
nand U42735 (N_42735,N_42487,N_42491);
and U42736 (N_42736,N_42395,N_42493);
nand U42737 (N_42737,N_42394,N_42487);
nand U42738 (N_42738,N_42421,N_42384);
nor U42739 (N_42739,N_42384,N_42283);
and U42740 (N_42740,N_42450,N_42393);
nand U42741 (N_42741,N_42437,N_42291);
nand U42742 (N_42742,N_42292,N_42396);
xor U42743 (N_42743,N_42471,N_42390);
and U42744 (N_42744,N_42333,N_42408);
nand U42745 (N_42745,N_42396,N_42436);
nor U42746 (N_42746,N_42285,N_42376);
xor U42747 (N_42747,N_42496,N_42472);
or U42748 (N_42748,N_42474,N_42394);
or U42749 (N_42749,N_42359,N_42291);
or U42750 (N_42750,N_42609,N_42672);
and U42751 (N_42751,N_42733,N_42644);
nand U42752 (N_42752,N_42652,N_42532);
and U42753 (N_42753,N_42740,N_42696);
or U42754 (N_42754,N_42548,N_42725);
nand U42755 (N_42755,N_42688,N_42523);
and U42756 (N_42756,N_42570,N_42508);
and U42757 (N_42757,N_42573,N_42637);
and U42758 (N_42758,N_42514,N_42565);
nand U42759 (N_42759,N_42554,N_42675);
nor U42760 (N_42760,N_42651,N_42525);
nor U42761 (N_42761,N_42533,N_42623);
or U42762 (N_42762,N_42575,N_42661);
or U42763 (N_42763,N_42670,N_42539);
nand U42764 (N_42764,N_42530,N_42596);
nand U42765 (N_42765,N_42737,N_42543);
or U42766 (N_42766,N_42657,N_42723);
nor U42767 (N_42767,N_42622,N_42621);
and U42768 (N_42768,N_42580,N_42556);
nand U42769 (N_42769,N_42625,N_42536);
or U42770 (N_42770,N_42526,N_42615);
xor U42771 (N_42771,N_42607,N_42666);
nor U42772 (N_42772,N_42743,N_42597);
and U42773 (N_42773,N_42714,N_42674);
or U42774 (N_42774,N_42582,N_42600);
and U42775 (N_42775,N_42679,N_42531);
nor U42776 (N_42776,N_42519,N_42535);
nand U42777 (N_42777,N_42587,N_42728);
or U42778 (N_42778,N_42569,N_42617);
nor U42779 (N_42779,N_42738,N_42624);
nand U42780 (N_42780,N_42748,N_42640);
nor U42781 (N_42781,N_42683,N_42719);
and U42782 (N_42782,N_42520,N_42558);
xnor U42783 (N_42783,N_42638,N_42593);
xnor U42784 (N_42784,N_42694,N_42678);
or U42785 (N_42785,N_42635,N_42591);
nand U42786 (N_42786,N_42673,N_42668);
xnor U42787 (N_42787,N_42560,N_42549);
or U42788 (N_42788,N_42629,N_42701);
nor U42789 (N_42789,N_42524,N_42712);
or U42790 (N_42790,N_42703,N_42574);
or U42791 (N_42791,N_42538,N_42527);
nor U42792 (N_42792,N_42581,N_42730);
or U42793 (N_42793,N_42641,N_42613);
xnor U42794 (N_42794,N_42616,N_42620);
or U42795 (N_42795,N_42511,N_42653);
or U42796 (N_42796,N_42503,N_42612);
xnor U42797 (N_42797,N_42537,N_42687);
nor U42798 (N_42798,N_42685,N_42544);
nand U42799 (N_42799,N_42501,N_42542);
or U42800 (N_42800,N_42504,N_42708);
or U42801 (N_42801,N_42669,N_42643);
nand U42802 (N_42802,N_42695,N_42506);
nand U42803 (N_42803,N_42512,N_42577);
nand U42804 (N_42804,N_42516,N_42736);
xnor U42805 (N_42805,N_42734,N_42630);
nand U42806 (N_42806,N_42727,N_42572);
and U42807 (N_42807,N_42626,N_42718);
nor U42808 (N_42808,N_42729,N_42632);
and U42809 (N_42809,N_42715,N_42724);
xor U42810 (N_42810,N_42707,N_42744);
nand U42811 (N_42811,N_42717,N_42610);
nor U42812 (N_42812,N_42742,N_42557);
xor U42813 (N_42813,N_42713,N_42731);
xnor U42814 (N_42814,N_42601,N_42509);
xor U42815 (N_42815,N_42552,N_42513);
nor U42816 (N_42816,N_42576,N_42528);
nor U42817 (N_42817,N_42656,N_42691);
or U42818 (N_42818,N_42602,N_42721);
and U42819 (N_42819,N_42650,N_42749);
and U42820 (N_42820,N_42660,N_42633);
or U42821 (N_42821,N_42510,N_42655);
nand U42822 (N_42822,N_42711,N_42690);
nor U42823 (N_42823,N_42639,N_42561);
and U42824 (N_42824,N_42692,N_42568);
nand U42825 (N_42825,N_42704,N_42677);
nand U42826 (N_42826,N_42579,N_42592);
and U42827 (N_42827,N_42578,N_42540);
nor U42828 (N_42828,N_42664,N_42546);
or U42829 (N_42829,N_42746,N_42559);
nand U42830 (N_42830,N_42588,N_42710);
nand U42831 (N_42831,N_42706,N_42636);
nand U42832 (N_42832,N_42689,N_42505);
xnor U42833 (N_42833,N_42665,N_42619);
and U42834 (N_42834,N_42502,N_42646);
xnor U42835 (N_42835,N_42662,N_42699);
or U42836 (N_42836,N_42522,N_42605);
or U42837 (N_42837,N_42747,N_42534);
nor U42838 (N_42838,N_42603,N_42551);
or U42839 (N_42839,N_42604,N_42553);
or U42840 (N_42840,N_42698,N_42606);
nor U42841 (N_42841,N_42716,N_42590);
xnor U42842 (N_42842,N_42722,N_42697);
or U42843 (N_42843,N_42726,N_42667);
xnor U42844 (N_42844,N_42705,N_42529);
or U42845 (N_42845,N_42517,N_42628);
xnor U42846 (N_42846,N_42564,N_42709);
nand U42847 (N_42847,N_42595,N_42584);
xnor U42848 (N_42848,N_42693,N_42586);
nand U42849 (N_42849,N_42659,N_42634);
or U42850 (N_42850,N_42547,N_42594);
or U42851 (N_42851,N_42732,N_42589);
nand U42852 (N_42852,N_42648,N_42618);
xor U42853 (N_42853,N_42614,N_42562);
and U42854 (N_42854,N_42720,N_42663);
and U42855 (N_42855,N_42647,N_42507);
and U42856 (N_42856,N_42649,N_42563);
nand U42857 (N_42857,N_42745,N_42631);
nand U42858 (N_42858,N_42671,N_42599);
xor U42859 (N_42859,N_42571,N_42676);
nand U42860 (N_42860,N_42515,N_42566);
xor U42861 (N_42861,N_42684,N_42627);
nor U42862 (N_42862,N_42686,N_42681);
and U42863 (N_42863,N_42585,N_42682);
nor U42864 (N_42864,N_42541,N_42611);
xor U42865 (N_42865,N_42654,N_42680);
or U42866 (N_42866,N_42735,N_42550);
nand U42867 (N_42867,N_42545,N_42700);
and U42868 (N_42868,N_42658,N_42645);
or U42869 (N_42869,N_42739,N_42521);
or U42870 (N_42870,N_42598,N_42741);
nand U42871 (N_42871,N_42518,N_42702);
nor U42872 (N_42872,N_42500,N_42555);
nor U42873 (N_42873,N_42608,N_42583);
nand U42874 (N_42874,N_42567,N_42642);
xnor U42875 (N_42875,N_42569,N_42500);
nand U42876 (N_42876,N_42660,N_42604);
xnor U42877 (N_42877,N_42680,N_42581);
nand U42878 (N_42878,N_42681,N_42579);
nand U42879 (N_42879,N_42722,N_42577);
or U42880 (N_42880,N_42552,N_42591);
and U42881 (N_42881,N_42652,N_42633);
xnor U42882 (N_42882,N_42596,N_42681);
or U42883 (N_42883,N_42514,N_42575);
or U42884 (N_42884,N_42675,N_42546);
nor U42885 (N_42885,N_42600,N_42740);
nor U42886 (N_42886,N_42639,N_42677);
and U42887 (N_42887,N_42715,N_42557);
nand U42888 (N_42888,N_42706,N_42638);
nor U42889 (N_42889,N_42668,N_42628);
or U42890 (N_42890,N_42683,N_42532);
xnor U42891 (N_42891,N_42559,N_42680);
and U42892 (N_42892,N_42661,N_42539);
and U42893 (N_42893,N_42737,N_42638);
and U42894 (N_42894,N_42588,N_42640);
nand U42895 (N_42895,N_42615,N_42732);
nor U42896 (N_42896,N_42636,N_42660);
xor U42897 (N_42897,N_42716,N_42536);
nor U42898 (N_42898,N_42670,N_42505);
nand U42899 (N_42899,N_42584,N_42643);
nor U42900 (N_42900,N_42526,N_42660);
xor U42901 (N_42901,N_42638,N_42556);
nor U42902 (N_42902,N_42622,N_42668);
nand U42903 (N_42903,N_42564,N_42578);
nand U42904 (N_42904,N_42731,N_42590);
or U42905 (N_42905,N_42707,N_42657);
and U42906 (N_42906,N_42516,N_42652);
nor U42907 (N_42907,N_42690,N_42707);
and U42908 (N_42908,N_42665,N_42637);
and U42909 (N_42909,N_42688,N_42727);
xor U42910 (N_42910,N_42597,N_42675);
xor U42911 (N_42911,N_42656,N_42539);
or U42912 (N_42912,N_42695,N_42634);
and U42913 (N_42913,N_42669,N_42617);
nor U42914 (N_42914,N_42561,N_42668);
nor U42915 (N_42915,N_42578,N_42515);
nor U42916 (N_42916,N_42531,N_42701);
nand U42917 (N_42917,N_42714,N_42605);
nand U42918 (N_42918,N_42596,N_42688);
and U42919 (N_42919,N_42595,N_42577);
and U42920 (N_42920,N_42604,N_42518);
nor U42921 (N_42921,N_42704,N_42590);
or U42922 (N_42922,N_42627,N_42748);
or U42923 (N_42923,N_42507,N_42592);
xor U42924 (N_42924,N_42528,N_42629);
xor U42925 (N_42925,N_42584,N_42719);
xor U42926 (N_42926,N_42725,N_42636);
xor U42927 (N_42927,N_42583,N_42506);
or U42928 (N_42928,N_42597,N_42565);
and U42929 (N_42929,N_42668,N_42581);
or U42930 (N_42930,N_42600,N_42697);
nor U42931 (N_42931,N_42520,N_42671);
xnor U42932 (N_42932,N_42515,N_42724);
xnor U42933 (N_42933,N_42706,N_42662);
xnor U42934 (N_42934,N_42673,N_42676);
xor U42935 (N_42935,N_42609,N_42619);
or U42936 (N_42936,N_42579,N_42731);
xnor U42937 (N_42937,N_42701,N_42747);
or U42938 (N_42938,N_42551,N_42636);
nor U42939 (N_42939,N_42500,N_42675);
nand U42940 (N_42940,N_42659,N_42684);
nand U42941 (N_42941,N_42645,N_42522);
nand U42942 (N_42942,N_42695,N_42500);
and U42943 (N_42943,N_42536,N_42592);
xnor U42944 (N_42944,N_42714,N_42744);
xnor U42945 (N_42945,N_42618,N_42543);
or U42946 (N_42946,N_42665,N_42746);
nand U42947 (N_42947,N_42583,N_42549);
and U42948 (N_42948,N_42556,N_42612);
nand U42949 (N_42949,N_42672,N_42661);
and U42950 (N_42950,N_42671,N_42746);
or U42951 (N_42951,N_42687,N_42613);
nand U42952 (N_42952,N_42551,N_42617);
nor U42953 (N_42953,N_42738,N_42691);
xor U42954 (N_42954,N_42691,N_42665);
nor U42955 (N_42955,N_42684,N_42584);
nand U42956 (N_42956,N_42722,N_42748);
or U42957 (N_42957,N_42668,N_42528);
nand U42958 (N_42958,N_42655,N_42516);
xnor U42959 (N_42959,N_42658,N_42702);
nand U42960 (N_42960,N_42538,N_42692);
xor U42961 (N_42961,N_42555,N_42570);
and U42962 (N_42962,N_42689,N_42741);
nand U42963 (N_42963,N_42520,N_42596);
or U42964 (N_42964,N_42717,N_42671);
nand U42965 (N_42965,N_42600,N_42603);
nor U42966 (N_42966,N_42631,N_42536);
or U42967 (N_42967,N_42551,N_42591);
xor U42968 (N_42968,N_42514,N_42722);
xor U42969 (N_42969,N_42592,N_42550);
and U42970 (N_42970,N_42747,N_42586);
nor U42971 (N_42971,N_42733,N_42727);
nand U42972 (N_42972,N_42721,N_42644);
xor U42973 (N_42973,N_42599,N_42714);
nand U42974 (N_42974,N_42691,N_42517);
nand U42975 (N_42975,N_42654,N_42502);
and U42976 (N_42976,N_42531,N_42714);
xor U42977 (N_42977,N_42729,N_42537);
xor U42978 (N_42978,N_42697,N_42528);
and U42979 (N_42979,N_42563,N_42695);
and U42980 (N_42980,N_42643,N_42586);
nor U42981 (N_42981,N_42517,N_42608);
xnor U42982 (N_42982,N_42728,N_42661);
xnor U42983 (N_42983,N_42716,N_42622);
xnor U42984 (N_42984,N_42736,N_42631);
xor U42985 (N_42985,N_42706,N_42743);
nor U42986 (N_42986,N_42706,N_42654);
xor U42987 (N_42987,N_42609,N_42517);
or U42988 (N_42988,N_42570,N_42615);
nand U42989 (N_42989,N_42732,N_42586);
nor U42990 (N_42990,N_42584,N_42571);
nand U42991 (N_42991,N_42596,N_42556);
nor U42992 (N_42992,N_42524,N_42553);
or U42993 (N_42993,N_42746,N_42669);
nor U42994 (N_42994,N_42503,N_42708);
nand U42995 (N_42995,N_42713,N_42699);
nand U42996 (N_42996,N_42555,N_42629);
xor U42997 (N_42997,N_42709,N_42638);
nor U42998 (N_42998,N_42723,N_42598);
nand U42999 (N_42999,N_42504,N_42745);
nor U43000 (N_43000,N_42920,N_42960);
nor U43001 (N_43001,N_42848,N_42882);
nor U43002 (N_43002,N_42880,N_42790);
nand U43003 (N_43003,N_42964,N_42830);
nand U43004 (N_43004,N_42902,N_42860);
xor U43005 (N_43005,N_42835,N_42752);
or U43006 (N_43006,N_42912,N_42766);
or U43007 (N_43007,N_42973,N_42984);
or U43008 (N_43008,N_42893,N_42886);
nand U43009 (N_43009,N_42926,N_42769);
and U43010 (N_43010,N_42932,N_42821);
nor U43011 (N_43011,N_42846,N_42781);
nand U43012 (N_43012,N_42971,N_42887);
or U43013 (N_43013,N_42784,N_42833);
nor U43014 (N_43014,N_42849,N_42757);
and U43015 (N_43015,N_42888,N_42905);
or U43016 (N_43016,N_42758,N_42760);
and U43017 (N_43017,N_42844,N_42962);
nand U43018 (N_43018,N_42816,N_42797);
nor U43019 (N_43019,N_42947,N_42802);
nor U43020 (N_43020,N_42814,N_42901);
nand U43021 (N_43021,N_42904,N_42764);
and U43022 (N_43022,N_42870,N_42751);
xor U43023 (N_43023,N_42866,N_42909);
and U43024 (N_43024,N_42883,N_42968);
nand U43025 (N_43025,N_42896,N_42987);
xnor U43026 (N_43026,N_42859,N_42782);
nor U43027 (N_43027,N_42874,N_42818);
or U43028 (N_43028,N_42990,N_42765);
or U43029 (N_43029,N_42850,N_42789);
nor U43030 (N_43030,N_42998,N_42967);
nor U43031 (N_43031,N_42875,N_42950);
nand U43032 (N_43032,N_42956,N_42750);
or U43033 (N_43033,N_42899,N_42916);
xor U43034 (N_43034,N_42858,N_42953);
nor U43035 (N_43035,N_42892,N_42838);
nor U43036 (N_43036,N_42891,N_42890);
nand U43037 (N_43037,N_42805,N_42812);
xnor U43038 (N_43038,N_42770,N_42930);
nand U43039 (N_43039,N_42911,N_42780);
nand U43040 (N_43040,N_42785,N_42915);
nand U43041 (N_43041,N_42986,N_42929);
xor U43042 (N_43042,N_42980,N_42829);
nand U43043 (N_43043,N_42771,N_42863);
xor U43044 (N_43044,N_42940,N_42801);
xnor U43045 (N_43045,N_42997,N_42935);
and U43046 (N_43046,N_42753,N_42803);
or U43047 (N_43047,N_42871,N_42806);
or U43048 (N_43048,N_42857,N_42910);
nor U43049 (N_43049,N_42881,N_42832);
and U43050 (N_43050,N_42825,N_42921);
nand U43051 (N_43051,N_42991,N_42793);
or U43052 (N_43052,N_42869,N_42939);
and U43053 (N_43053,N_42836,N_42807);
nand U43054 (N_43054,N_42810,N_42800);
nand U43055 (N_43055,N_42755,N_42958);
or U43056 (N_43056,N_42925,N_42999);
xnor U43057 (N_43057,N_42970,N_42855);
and U43058 (N_43058,N_42817,N_42819);
and U43059 (N_43059,N_42954,N_42943);
nand U43060 (N_43060,N_42777,N_42783);
nor U43061 (N_43061,N_42982,N_42983);
nand U43062 (N_43062,N_42903,N_42972);
nand U43063 (N_43063,N_42878,N_42913);
and U43064 (N_43064,N_42897,N_42949);
and U43065 (N_43065,N_42876,N_42884);
and U43066 (N_43066,N_42772,N_42778);
or U43067 (N_43067,N_42839,N_42868);
xor U43068 (N_43068,N_42918,N_42872);
nand U43069 (N_43069,N_42865,N_42948);
or U43070 (N_43070,N_42952,N_42877);
and U43071 (N_43071,N_42774,N_42864);
or U43072 (N_43072,N_42754,N_42900);
and U43073 (N_43073,N_42792,N_42787);
xnor U43074 (N_43074,N_42831,N_42840);
or U43075 (N_43075,N_42873,N_42919);
nand U43076 (N_43076,N_42936,N_42989);
xor U43077 (N_43077,N_42898,N_42809);
nand U43078 (N_43078,N_42931,N_42908);
or U43079 (N_43079,N_42977,N_42826);
or U43080 (N_43080,N_42934,N_42854);
nor U43081 (N_43081,N_42756,N_42974);
and U43082 (N_43082,N_42853,N_42867);
nor U43083 (N_43083,N_42791,N_42815);
and U43084 (N_43084,N_42907,N_42963);
nor U43085 (N_43085,N_42852,N_42988);
and U43086 (N_43086,N_42773,N_42822);
nand U43087 (N_43087,N_42914,N_42922);
xor U43088 (N_43088,N_42862,N_42799);
nand U43089 (N_43089,N_42842,N_42996);
or U43090 (N_43090,N_42851,N_42834);
nor U43091 (N_43091,N_42927,N_42837);
nand U43092 (N_43092,N_42761,N_42767);
or U43093 (N_43093,N_42813,N_42856);
xnor U43094 (N_43094,N_42794,N_42944);
or U43095 (N_43095,N_42775,N_42768);
nor U43096 (N_43096,N_42917,N_42786);
and U43097 (N_43097,N_42879,N_42843);
nor U43098 (N_43098,N_42975,N_42796);
or U43099 (N_43099,N_42946,N_42795);
or U43100 (N_43100,N_42941,N_42961);
nand U43101 (N_43101,N_42951,N_42937);
and U43102 (N_43102,N_42965,N_42993);
nor U43103 (N_43103,N_42979,N_42847);
xor U43104 (N_43104,N_42994,N_42928);
nor U43105 (N_43105,N_42955,N_42824);
xor U43106 (N_43106,N_42959,N_42923);
nor U43107 (N_43107,N_42889,N_42804);
and U43108 (N_43108,N_42811,N_42779);
nor U43109 (N_43109,N_42828,N_42981);
and U43110 (N_43110,N_42841,N_42894);
nand U43111 (N_43111,N_42885,N_42942);
or U43112 (N_43112,N_42906,N_42995);
or U43113 (N_43113,N_42969,N_42845);
or U43114 (N_43114,N_42823,N_42978);
nor U43115 (N_43115,N_42966,N_42763);
xor U43116 (N_43116,N_42976,N_42895);
or U43117 (N_43117,N_42992,N_42776);
nor U43118 (N_43118,N_42933,N_42798);
or U43119 (N_43119,N_42985,N_42788);
and U43120 (N_43120,N_42924,N_42938);
xnor U43121 (N_43121,N_42957,N_42759);
or U43122 (N_43122,N_42762,N_42945);
xnor U43123 (N_43123,N_42827,N_42820);
nand U43124 (N_43124,N_42808,N_42861);
nor U43125 (N_43125,N_42803,N_42755);
nor U43126 (N_43126,N_42853,N_42799);
xnor U43127 (N_43127,N_42850,N_42853);
or U43128 (N_43128,N_42958,N_42976);
or U43129 (N_43129,N_42782,N_42910);
or U43130 (N_43130,N_42991,N_42760);
xnor U43131 (N_43131,N_42775,N_42853);
xnor U43132 (N_43132,N_42982,N_42800);
xor U43133 (N_43133,N_42995,N_42840);
or U43134 (N_43134,N_42859,N_42866);
and U43135 (N_43135,N_42772,N_42801);
nand U43136 (N_43136,N_42973,N_42909);
and U43137 (N_43137,N_42755,N_42925);
nand U43138 (N_43138,N_42856,N_42877);
or U43139 (N_43139,N_42751,N_42836);
nand U43140 (N_43140,N_42966,N_42847);
xor U43141 (N_43141,N_42996,N_42837);
xor U43142 (N_43142,N_42895,N_42931);
xor U43143 (N_43143,N_42858,N_42861);
nand U43144 (N_43144,N_42821,N_42992);
nand U43145 (N_43145,N_42916,N_42904);
or U43146 (N_43146,N_42950,N_42801);
nor U43147 (N_43147,N_42890,N_42924);
nor U43148 (N_43148,N_42914,N_42796);
or U43149 (N_43149,N_42816,N_42999);
nor U43150 (N_43150,N_42970,N_42820);
nor U43151 (N_43151,N_42803,N_42845);
and U43152 (N_43152,N_42811,N_42966);
nor U43153 (N_43153,N_42990,N_42900);
xor U43154 (N_43154,N_42816,N_42889);
or U43155 (N_43155,N_42927,N_42782);
nand U43156 (N_43156,N_42783,N_42999);
and U43157 (N_43157,N_42760,N_42753);
and U43158 (N_43158,N_42783,N_42836);
xor U43159 (N_43159,N_42963,N_42922);
nand U43160 (N_43160,N_42788,N_42778);
nor U43161 (N_43161,N_42834,N_42883);
and U43162 (N_43162,N_42796,N_42854);
or U43163 (N_43163,N_42846,N_42834);
nand U43164 (N_43164,N_42926,N_42970);
or U43165 (N_43165,N_42908,N_42872);
nand U43166 (N_43166,N_42756,N_42995);
nor U43167 (N_43167,N_42751,N_42977);
and U43168 (N_43168,N_42755,N_42860);
nor U43169 (N_43169,N_42870,N_42958);
nand U43170 (N_43170,N_42761,N_42820);
xor U43171 (N_43171,N_42929,N_42841);
nand U43172 (N_43172,N_42776,N_42853);
nand U43173 (N_43173,N_42994,N_42865);
nor U43174 (N_43174,N_42882,N_42782);
and U43175 (N_43175,N_42924,N_42858);
nand U43176 (N_43176,N_42833,N_42911);
nor U43177 (N_43177,N_42829,N_42814);
and U43178 (N_43178,N_42906,N_42862);
or U43179 (N_43179,N_42990,N_42951);
nand U43180 (N_43180,N_42788,N_42898);
nor U43181 (N_43181,N_42851,N_42901);
and U43182 (N_43182,N_42823,N_42976);
and U43183 (N_43183,N_42855,N_42870);
and U43184 (N_43184,N_42834,N_42874);
and U43185 (N_43185,N_42805,N_42776);
xnor U43186 (N_43186,N_42917,N_42873);
or U43187 (N_43187,N_42802,N_42813);
xor U43188 (N_43188,N_42782,N_42838);
xor U43189 (N_43189,N_42930,N_42913);
xor U43190 (N_43190,N_42950,N_42802);
xor U43191 (N_43191,N_42907,N_42914);
nor U43192 (N_43192,N_42899,N_42994);
or U43193 (N_43193,N_42983,N_42927);
nor U43194 (N_43194,N_42968,N_42890);
nand U43195 (N_43195,N_42848,N_42839);
or U43196 (N_43196,N_42770,N_42897);
nor U43197 (N_43197,N_42782,N_42993);
nand U43198 (N_43198,N_42800,N_42796);
nand U43199 (N_43199,N_42944,N_42942);
and U43200 (N_43200,N_42847,N_42753);
nor U43201 (N_43201,N_42938,N_42954);
xnor U43202 (N_43202,N_42752,N_42905);
nand U43203 (N_43203,N_42907,N_42811);
nor U43204 (N_43204,N_42804,N_42995);
nor U43205 (N_43205,N_42804,N_42831);
nor U43206 (N_43206,N_42995,N_42799);
nand U43207 (N_43207,N_42878,N_42923);
nand U43208 (N_43208,N_42970,N_42763);
nor U43209 (N_43209,N_42893,N_42763);
and U43210 (N_43210,N_42863,N_42951);
nor U43211 (N_43211,N_42999,N_42857);
nand U43212 (N_43212,N_42987,N_42844);
nor U43213 (N_43213,N_42855,N_42859);
nor U43214 (N_43214,N_42883,N_42958);
nand U43215 (N_43215,N_42805,N_42773);
nand U43216 (N_43216,N_42854,N_42771);
and U43217 (N_43217,N_42934,N_42937);
or U43218 (N_43218,N_42907,N_42820);
nor U43219 (N_43219,N_42927,N_42751);
and U43220 (N_43220,N_42908,N_42858);
nor U43221 (N_43221,N_42754,N_42828);
nand U43222 (N_43222,N_42961,N_42824);
nand U43223 (N_43223,N_42945,N_42861);
or U43224 (N_43224,N_42953,N_42871);
nand U43225 (N_43225,N_42987,N_42943);
xor U43226 (N_43226,N_42972,N_42921);
xor U43227 (N_43227,N_42880,N_42799);
xor U43228 (N_43228,N_42801,N_42878);
and U43229 (N_43229,N_42913,N_42836);
xor U43230 (N_43230,N_42900,N_42765);
and U43231 (N_43231,N_42944,N_42823);
nor U43232 (N_43232,N_42946,N_42819);
xor U43233 (N_43233,N_42872,N_42999);
or U43234 (N_43234,N_42752,N_42907);
nor U43235 (N_43235,N_42793,N_42825);
nor U43236 (N_43236,N_42938,N_42845);
or U43237 (N_43237,N_42843,N_42882);
nor U43238 (N_43238,N_42861,N_42881);
xor U43239 (N_43239,N_42873,N_42783);
and U43240 (N_43240,N_42900,N_42961);
or U43241 (N_43241,N_42822,N_42964);
and U43242 (N_43242,N_42776,N_42966);
nand U43243 (N_43243,N_42855,N_42802);
or U43244 (N_43244,N_42781,N_42944);
and U43245 (N_43245,N_42898,N_42971);
or U43246 (N_43246,N_42879,N_42787);
nand U43247 (N_43247,N_42976,N_42933);
xnor U43248 (N_43248,N_42786,N_42847);
or U43249 (N_43249,N_42944,N_42789);
nor U43250 (N_43250,N_43155,N_43066);
nand U43251 (N_43251,N_43178,N_43023);
and U43252 (N_43252,N_43226,N_43103);
xnor U43253 (N_43253,N_43236,N_43068);
or U43254 (N_43254,N_43051,N_43010);
nor U43255 (N_43255,N_43181,N_43119);
nand U43256 (N_43256,N_43197,N_43143);
or U43257 (N_43257,N_43011,N_43128);
nand U43258 (N_43258,N_43209,N_43002);
and U43259 (N_43259,N_43158,N_43164);
and U43260 (N_43260,N_43021,N_43201);
and U43261 (N_43261,N_43091,N_43049);
and U43262 (N_43262,N_43124,N_43136);
xor U43263 (N_43263,N_43229,N_43097);
and U43264 (N_43264,N_43216,N_43012);
or U43265 (N_43265,N_43234,N_43151);
and U43266 (N_43266,N_43227,N_43044);
nand U43267 (N_43267,N_43015,N_43099);
nor U43268 (N_43268,N_43083,N_43007);
nor U43269 (N_43269,N_43108,N_43195);
nor U43270 (N_43270,N_43064,N_43207);
nor U43271 (N_43271,N_43240,N_43038);
xnor U43272 (N_43272,N_43190,N_43067);
nand U43273 (N_43273,N_43019,N_43154);
or U43274 (N_43274,N_43070,N_43123);
and U43275 (N_43275,N_43183,N_43228);
or U43276 (N_43276,N_43187,N_43045);
or U43277 (N_43277,N_43213,N_43144);
nand U43278 (N_43278,N_43221,N_43041);
nand U43279 (N_43279,N_43173,N_43217);
nand U43280 (N_43280,N_43102,N_43107);
or U43281 (N_43281,N_43106,N_43192);
and U43282 (N_43282,N_43249,N_43105);
nand U43283 (N_43283,N_43057,N_43167);
nor U43284 (N_43284,N_43176,N_43037);
and U43285 (N_43285,N_43193,N_43239);
nor U43286 (N_43286,N_43206,N_43001);
xnor U43287 (N_43287,N_43118,N_43179);
and U43288 (N_43288,N_43157,N_43247);
nand U43289 (N_43289,N_43244,N_43082);
nand U43290 (N_43290,N_43222,N_43059);
nand U43291 (N_43291,N_43163,N_43086);
or U43292 (N_43292,N_43110,N_43026);
nand U43293 (N_43293,N_43036,N_43246);
or U43294 (N_43294,N_43203,N_43039);
nand U43295 (N_43295,N_43101,N_43077);
and U43296 (N_43296,N_43081,N_43138);
and U43297 (N_43297,N_43223,N_43235);
nand U43298 (N_43298,N_43120,N_43225);
nor U43299 (N_43299,N_43243,N_43000);
nor U43300 (N_43300,N_43146,N_43009);
or U43301 (N_43301,N_43104,N_43212);
nor U43302 (N_43302,N_43175,N_43072);
or U43303 (N_43303,N_43150,N_43092);
nor U43304 (N_43304,N_43126,N_43112);
or U43305 (N_43305,N_43109,N_43090);
nor U43306 (N_43306,N_43153,N_43141);
or U43307 (N_43307,N_43125,N_43199);
xnor U43308 (N_43308,N_43050,N_43028);
or U43309 (N_43309,N_43063,N_43020);
xor U43310 (N_43310,N_43029,N_43084);
and U43311 (N_43311,N_43114,N_43232);
xor U43312 (N_43312,N_43055,N_43152);
or U43313 (N_43313,N_43061,N_43230);
nor U43314 (N_43314,N_43211,N_43134);
nor U43315 (N_43315,N_43185,N_43191);
nor U43316 (N_43316,N_43162,N_43014);
nor U43317 (N_43317,N_43184,N_43115);
or U43318 (N_43318,N_43165,N_43169);
nor U43319 (N_43319,N_43048,N_43139);
nand U43320 (N_43320,N_43194,N_43046);
or U43321 (N_43321,N_43121,N_43135);
and U43322 (N_43322,N_43218,N_43075);
xnor U43323 (N_43323,N_43079,N_43030);
nand U43324 (N_43324,N_43111,N_43137);
nor U43325 (N_43325,N_43076,N_43188);
xor U43326 (N_43326,N_43204,N_43005);
nor U43327 (N_43327,N_43008,N_43168);
nor U43328 (N_43328,N_43022,N_43043);
nor U43329 (N_43329,N_43214,N_43034);
xnor U43330 (N_43330,N_43078,N_43042);
nand U43331 (N_43331,N_43215,N_43170);
or U43332 (N_43332,N_43241,N_43147);
or U43333 (N_43333,N_43127,N_43025);
nor U43334 (N_43334,N_43089,N_43027);
nor U43335 (N_43335,N_43189,N_43085);
and U43336 (N_43336,N_43210,N_43074);
or U43337 (N_43337,N_43117,N_43245);
nor U43338 (N_43338,N_43198,N_43177);
or U43339 (N_43339,N_43040,N_43033);
nand U43340 (N_43340,N_43208,N_43171);
xnor U43341 (N_43341,N_43205,N_43069);
and U43342 (N_43342,N_43047,N_43035);
nand U43343 (N_43343,N_43161,N_43156);
xor U43344 (N_43344,N_43238,N_43003);
nand U43345 (N_43345,N_43080,N_43174);
and U43346 (N_43346,N_43017,N_43095);
and U43347 (N_43347,N_43149,N_43142);
or U43348 (N_43348,N_43018,N_43013);
xor U43349 (N_43349,N_43133,N_43100);
nor U43350 (N_43350,N_43172,N_43098);
nor U43351 (N_43351,N_43006,N_43093);
nand U43352 (N_43352,N_43224,N_43159);
nor U43353 (N_43353,N_43096,N_43237);
or U43354 (N_43354,N_43056,N_43148);
or U43355 (N_43355,N_43132,N_43122);
and U43356 (N_43356,N_43032,N_43186);
and U43357 (N_43357,N_43231,N_43182);
nand U43358 (N_43358,N_43087,N_43062);
and U43359 (N_43359,N_43016,N_43088);
xor U43360 (N_43360,N_43145,N_43053);
xnor U43361 (N_43361,N_43140,N_43160);
or U43362 (N_43362,N_43166,N_43131);
nand U43363 (N_43363,N_43116,N_43065);
nand U43364 (N_43364,N_43073,N_43060);
xnor U43365 (N_43365,N_43071,N_43094);
or U43366 (N_43366,N_43052,N_43113);
xnor U43367 (N_43367,N_43004,N_43129);
nand U43368 (N_43368,N_43248,N_43054);
or U43369 (N_43369,N_43233,N_43130);
and U43370 (N_43370,N_43058,N_43202);
xor U43371 (N_43371,N_43031,N_43024);
xnor U43372 (N_43372,N_43220,N_43200);
nand U43373 (N_43373,N_43180,N_43242);
or U43374 (N_43374,N_43196,N_43219);
nand U43375 (N_43375,N_43230,N_43067);
xnor U43376 (N_43376,N_43016,N_43175);
nand U43377 (N_43377,N_43176,N_43177);
nor U43378 (N_43378,N_43145,N_43214);
nand U43379 (N_43379,N_43019,N_43144);
xnor U43380 (N_43380,N_43040,N_43182);
and U43381 (N_43381,N_43027,N_43185);
nor U43382 (N_43382,N_43150,N_43070);
nor U43383 (N_43383,N_43023,N_43217);
nor U43384 (N_43384,N_43108,N_43135);
and U43385 (N_43385,N_43121,N_43169);
and U43386 (N_43386,N_43158,N_43089);
nor U43387 (N_43387,N_43179,N_43054);
nand U43388 (N_43388,N_43006,N_43128);
and U43389 (N_43389,N_43132,N_43047);
or U43390 (N_43390,N_43033,N_43129);
and U43391 (N_43391,N_43052,N_43041);
nor U43392 (N_43392,N_43002,N_43105);
nor U43393 (N_43393,N_43093,N_43016);
and U43394 (N_43394,N_43003,N_43109);
or U43395 (N_43395,N_43084,N_43026);
nor U43396 (N_43396,N_43008,N_43229);
nor U43397 (N_43397,N_43173,N_43244);
nor U43398 (N_43398,N_43010,N_43005);
and U43399 (N_43399,N_43196,N_43032);
nand U43400 (N_43400,N_43147,N_43017);
nand U43401 (N_43401,N_43215,N_43120);
xor U43402 (N_43402,N_43062,N_43091);
xnor U43403 (N_43403,N_43031,N_43015);
nand U43404 (N_43404,N_43226,N_43200);
xor U43405 (N_43405,N_43040,N_43096);
or U43406 (N_43406,N_43120,N_43136);
nand U43407 (N_43407,N_43237,N_43230);
or U43408 (N_43408,N_43045,N_43171);
nor U43409 (N_43409,N_43155,N_43070);
or U43410 (N_43410,N_43038,N_43158);
xor U43411 (N_43411,N_43158,N_43049);
and U43412 (N_43412,N_43040,N_43043);
nor U43413 (N_43413,N_43013,N_43127);
or U43414 (N_43414,N_43192,N_43081);
or U43415 (N_43415,N_43190,N_43086);
nor U43416 (N_43416,N_43211,N_43190);
nor U43417 (N_43417,N_43042,N_43044);
nor U43418 (N_43418,N_43082,N_43067);
xnor U43419 (N_43419,N_43219,N_43171);
or U43420 (N_43420,N_43104,N_43008);
and U43421 (N_43421,N_43151,N_43146);
or U43422 (N_43422,N_43108,N_43119);
nand U43423 (N_43423,N_43070,N_43156);
xor U43424 (N_43424,N_43240,N_43022);
and U43425 (N_43425,N_43193,N_43181);
and U43426 (N_43426,N_43053,N_43207);
or U43427 (N_43427,N_43137,N_43103);
or U43428 (N_43428,N_43228,N_43137);
and U43429 (N_43429,N_43017,N_43001);
or U43430 (N_43430,N_43175,N_43079);
nor U43431 (N_43431,N_43000,N_43165);
nand U43432 (N_43432,N_43020,N_43239);
nand U43433 (N_43433,N_43016,N_43212);
nor U43434 (N_43434,N_43191,N_43081);
or U43435 (N_43435,N_43128,N_43180);
nand U43436 (N_43436,N_43160,N_43145);
nand U43437 (N_43437,N_43017,N_43013);
and U43438 (N_43438,N_43059,N_43193);
xor U43439 (N_43439,N_43060,N_43152);
xor U43440 (N_43440,N_43050,N_43225);
nor U43441 (N_43441,N_43000,N_43176);
nand U43442 (N_43442,N_43164,N_43005);
or U43443 (N_43443,N_43141,N_43211);
nor U43444 (N_43444,N_43139,N_43076);
nand U43445 (N_43445,N_43191,N_43220);
nand U43446 (N_43446,N_43158,N_43156);
or U43447 (N_43447,N_43131,N_43158);
xnor U43448 (N_43448,N_43063,N_43016);
nor U43449 (N_43449,N_43217,N_43126);
xnor U43450 (N_43450,N_43136,N_43176);
and U43451 (N_43451,N_43119,N_43063);
nand U43452 (N_43452,N_43113,N_43025);
nor U43453 (N_43453,N_43245,N_43193);
nand U43454 (N_43454,N_43029,N_43086);
nand U43455 (N_43455,N_43004,N_43234);
nor U43456 (N_43456,N_43093,N_43082);
and U43457 (N_43457,N_43242,N_43177);
nand U43458 (N_43458,N_43001,N_43173);
or U43459 (N_43459,N_43232,N_43007);
and U43460 (N_43460,N_43229,N_43126);
and U43461 (N_43461,N_43206,N_43039);
xor U43462 (N_43462,N_43168,N_43214);
or U43463 (N_43463,N_43233,N_43101);
xnor U43464 (N_43464,N_43026,N_43208);
nand U43465 (N_43465,N_43027,N_43187);
nand U43466 (N_43466,N_43209,N_43080);
and U43467 (N_43467,N_43225,N_43057);
and U43468 (N_43468,N_43176,N_43117);
and U43469 (N_43469,N_43052,N_43035);
or U43470 (N_43470,N_43247,N_43057);
or U43471 (N_43471,N_43232,N_43161);
or U43472 (N_43472,N_43222,N_43019);
and U43473 (N_43473,N_43176,N_43077);
nor U43474 (N_43474,N_43129,N_43166);
xor U43475 (N_43475,N_43231,N_43153);
nor U43476 (N_43476,N_43147,N_43104);
nor U43477 (N_43477,N_43192,N_43143);
nor U43478 (N_43478,N_43194,N_43105);
xor U43479 (N_43479,N_43036,N_43039);
nand U43480 (N_43480,N_43175,N_43076);
nand U43481 (N_43481,N_43026,N_43122);
and U43482 (N_43482,N_43089,N_43180);
nand U43483 (N_43483,N_43136,N_43019);
and U43484 (N_43484,N_43036,N_43195);
nand U43485 (N_43485,N_43161,N_43229);
nor U43486 (N_43486,N_43162,N_43010);
and U43487 (N_43487,N_43122,N_43149);
nand U43488 (N_43488,N_43022,N_43168);
xnor U43489 (N_43489,N_43063,N_43105);
or U43490 (N_43490,N_43002,N_43071);
nand U43491 (N_43491,N_43214,N_43070);
nand U43492 (N_43492,N_43084,N_43094);
nand U43493 (N_43493,N_43159,N_43067);
and U43494 (N_43494,N_43000,N_43068);
and U43495 (N_43495,N_43012,N_43167);
nand U43496 (N_43496,N_43059,N_43234);
or U43497 (N_43497,N_43172,N_43182);
nand U43498 (N_43498,N_43001,N_43053);
xnor U43499 (N_43499,N_43043,N_43080);
nand U43500 (N_43500,N_43293,N_43438);
and U43501 (N_43501,N_43326,N_43482);
xnor U43502 (N_43502,N_43493,N_43345);
nand U43503 (N_43503,N_43453,N_43404);
or U43504 (N_43504,N_43400,N_43408);
nor U43505 (N_43505,N_43369,N_43465);
and U43506 (N_43506,N_43339,N_43316);
nor U43507 (N_43507,N_43439,N_43486);
and U43508 (N_43508,N_43391,N_43458);
nor U43509 (N_43509,N_43376,N_43269);
or U43510 (N_43510,N_43450,N_43432);
nand U43511 (N_43511,N_43488,N_43427);
nand U43512 (N_43512,N_43347,N_43274);
nand U43513 (N_43513,N_43288,N_43324);
xor U43514 (N_43514,N_43462,N_43492);
nor U43515 (N_43515,N_43323,N_43401);
nand U43516 (N_43516,N_43412,N_43346);
and U43517 (N_43517,N_43307,N_43365);
and U43518 (N_43518,N_43416,N_43296);
nand U43519 (N_43519,N_43421,N_43280);
nor U43520 (N_43520,N_43305,N_43487);
nor U43521 (N_43521,N_43394,N_43437);
nor U43522 (N_43522,N_43255,N_43333);
xor U43523 (N_43523,N_43448,N_43371);
or U43524 (N_43524,N_43431,N_43409);
xor U43525 (N_43525,N_43382,N_43373);
nor U43526 (N_43526,N_43387,N_43452);
nor U43527 (N_43527,N_43484,N_43367);
nor U43528 (N_43528,N_43499,N_43395);
or U43529 (N_43529,N_43270,N_43260);
nand U43530 (N_43530,N_43429,N_43337);
and U43531 (N_43531,N_43297,N_43455);
nand U43532 (N_43532,N_43257,N_43348);
or U43533 (N_43533,N_43413,N_43322);
xor U43534 (N_43534,N_43298,N_43489);
xor U43535 (N_43535,N_43271,N_43361);
nand U43536 (N_43536,N_43428,N_43470);
nand U43537 (N_43537,N_43385,N_43299);
nand U43538 (N_43538,N_43352,N_43253);
and U43539 (N_43539,N_43362,N_43300);
nand U43540 (N_43540,N_43491,N_43366);
and U43541 (N_43541,N_43498,N_43254);
and U43542 (N_43542,N_43418,N_43423);
and U43543 (N_43543,N_43278,N_43328);
and U43544 (N_43544,N_43301,N_43321);
and U43545 (N_43545,N_43331,N_43363);
and U43546 (N_43546,N_43405,N_43436);
xor U43547 (N_43547,N_43327,N_43442);
nand U43548 (N_43548,N_43334,N_43368);
and U43549 (N_43549,N_43314,N_43351);
or U43550 (N_43550,N_43474,N_43310);
xnor U43551 (N_43551,N_43497,N_43434);
nand U43552 (N_43552,N_43258,N_43384);
nand U43553 (N_43553,N_43496,N_43287);
nor U43554 (N_43554,N_43479,N_43318);
nor U43555 (N_43555,N_43289,N_43342);
and U43556 (N_43556,N_43313,N_43317);
or U43557 (N_43557,N_43273,N_43360);
and U43558 (N_43558,N_43353,N_43381);
or U43559 (N_43559,N_43449,N_43294);
nor U43560 (N_43560,N_43256,N_43282);
or U43561 (N_43561,N_43349,N_43414);
and U43562 (N_43562,N_43295,N_43403);
and U43563 (N_43563,N_43378,N_43444);
xnor U43564 (N_43564,N_43315,N_43471);
xor U43565 (N_43565,N_43475,N_43311);
nor U43566 (N_43566,N_43467,N_43251);
nor U43567 (N_43567,N_43397,N_43302);
or U43568 (N_43568,N_43377,N_43263);
nor U43569 (N_43569,N_43374,N_43285);
nand U43570 (N_43570,N_43425,N_43386);
nor U43571 (N_43571,N_43341,N_43355);
and U43572 (N_43572,N_43398,N_43332);
nor U43573 (N_43573,N_43451,N_43252);
nand U43574 (N_43574,N_43494,N_43456);
nor U43575 (N_43575,N_43485,N_43424);
xnor U43576 (N_43576,N_43473,N_43461);
and U43577 (N_43577,N_43272,N_43459);
and U43578 (N_43578,N_43303,N_43276);
xnor U43579 (N_43579,N_43250,N_43354);
or U43580 (N_43580,N_43440,N_43283);
xnor U43581 (N_43581,N_43264,N_43343);
or U43582 (N_43582,N_43281,N_43261);
nand U43583 (N_43583,N_43441,N_43259);
or U43584 (N_43584,N_43284,N_43370);
or U43585 (N_43585,N_43290,N_43320);
nand U43586 (N_43586,N_43292,N_43364);
xnor U43587 (N_43587,N_43420,N_43447);
nor U43588 (N_43588,N_43306,N_43399);
and U43589 (N_43589,N_43344,N_43356);
nor U43590 (N_43590,N_43262,N_43350);
nand U43591 (N_43591,N_43309,N_43481);
or U43592 (N_43592,N_43319,N_43410);
or U43593 (N_43593,N_43433,N_43291);
and U43594 (N_43594,N_43335,N_43480);
xnor U43595 (N_43595,N_43422,N_43325);
nor U43596 (N_43596,N_43435,N_43469);
or U43597 (N_43597,N_43464,N_43393);
xnor U43598 (N_43598,N_43478,N_43457);
and U43599 (N_43599,N_43419,N_43426);
and U43600 (N_43600,N_43286,N_43468);
nand U43601 (N_43601,N_43329,N_43443);
and U43602 (N_43602,N_43340,N_43275);
or U43603 (N_43603,N_43312,N_43379);
xor U43604 (N_43604,N_43396,N_43454);
and U43605 (N_43605,N_43463,N_43338);
and U43606 (N_43606,N_43389,N_43445);
xnor U43607 (N_43607,N_43268,N_43402);
nor U43608 (N_43608,N_43388,N_43267);
xor U43609 (N_43609,N_43415,N_43460);
xnor U43610 (N_43610,N_43430,N_43477);
or U43611 (N_43611,N_43304,N_43359);
xor U43612 (N_43612,N_43372,N_43277);
xor U43613 (N_43613,N_43380,N_43336);
or U43614 (N_43614,N_43358,N_43495);
or U43615 (N_43615,N_43266,N_43265);
or U43616 (N_43616,N_43279,N_43406);
nor U43617 (N_43617,N_43383,N_43330);
nand U43618 (N_43618,N_43490,N_43476);
nand U43619 (N_43619,N_43375,N_43411);
nor U43620 (N_43620,N_43392,N_43390);
xnor U43621 (N_43621,N_43472,N_43417);
xor U43622 (N_43622,N_43308,N_43483);
nor U43623 (N_43623,N_43466,N_43407);
or U43624 (N_43624,N_43357,N_43446);
and U43625 (N_43625,N_43268,N_43321);
or U43626 (N_43626,N_43423,N_43348);
nor U43627 (N_43627,N_43460,N_43422);
and U43628 (N_43628,N_43366,N_43421);
or U43629 (N_43629,N_43437,N_43445);
xor U43630 (N_43630,N_43445,N_43462);
nor U43631 (N_43631,N_43350,N_43327);
nor U43632 (N_43632,N_43434,N_43403);
xnor U43633 (N_43633,N_43343,N_43433);
nor U43634 (N_43634,N_43338,N_43482);
and U43635 (N_43635,N_43252,N_43431);
nand U43636 (N_43636,N_43336,N_43365);
nor U43637 (N_43637,N_43293,N_43402);
nand U43638 (N_43638,N_43383,N_43343);
or U43639 (N_43639,N_43315,N_43332);
nand U43640 (N_43640,N_43492,N_43436);
nand U43641 (N_43641,N_43287,N_43452);
xnor U43642 (N_43642,N_43350,N_43294);
nand U43643 (N_43643,N_43360,N_43260);
nor U43644 (N_43644,N_43340,N_43478);
nor U43645 (N_43645,N_43306,N_43278);
xor U43646 (N_43646,N_43254,N_43261);
nand U43647 (N_43647,N_43480,N_43414);
or U43648 (N_43648,N_43255,N_43386);
nand U43649 (N_43649,N_43281,N_43296);
nor U43650 (N_43650,N_43338,N_43458);
and U43651 (N_43651,N_43403,N_43485);
nand U43652 (N_43652,N_43356,N_43351);
xor U43653 (N_43653,N_43465,N_43458);
nand U43654 (N_43654,N_43366,N_43367);
nor U43655 (N_43655,N_43484,N_43414);
or U43656 (N_43656,N_43317,N_43397);
xor U43657 (N_43657,N_43420,N_43340);
xor U43658 (N_43658,N_43283,N_43408);
nand U43659 (N_43659,N_43409,N_43351);
or U43660 (N_43660,N_43385,N_43485);
or U43661 (N_43661,N_43483,N_43320);
or U43662 (N_43662,N_43331,N_43497);
or U43663 (N_43663,N_43266,N_43317);
nand U43664 (N_43664,N_43494,N_43437);
or U43665 (N_43665,N_43432,N_43466);
nor U43666 (N_43666,N_43315,N_43423);
nand U43667 (N_43667,N_43481,N_43289);
or U43668 (N_43668,N_43447,N_43433);
nand U43669 (N_43669,N_43457,N_43298);
nand U43670 (N_43670,N_43332,N_43405);
nand U43671 (N_43671,N_43269,N_43422);
nand U43672 (N_43672,N_43415,N_43448);
nor U43673 (N_43673,N_43496,N_43448);
nand U43674 (N_43674,N_43297,N_43397);
and U43675 (N_43675,N_43333,N_43274);
or U43676 (N_43676,N_43455,N_43272);
and U43677 (N_43677,N_43495,N_43445);
nor U43678 (N_43678,N_43295,N_43369);
xor U43679 (N_43679,N_43416,N_43371);
and U43680 (N_43680,N_43485,N_43286);
nand U43681 (N_43681,N_43495,N_43349);
and U43682 (N_43682,N_43311,N_43328);
and U43683 (N_43683,N_43372,N_43308);
nand U43684 (N_43684,N_43279,N_43429);
xor U43685 (N_43685,N_43382,N_43330);
or U43686 (N_43686,N_43346,N_43409);
xnor U43687 (N_43687,N_43356,N_43308);
and U43688 (N_43688,N_43424,N_43428);
nor U43689 (N_43689,N_43279,N_43318);
xor U43690 (N_43690,N_43438,N_43403);
nor U43691 (N_43691,N_43483,N_43369);
xor U43692 (N_43692,N_43356,N_43477);
and U43693 (N_43693,N_43405,N_43451);
and U43694 (N_43694,N_43427,N_43328);
nand U43695 (N_43695,N_43377,N_43378);
or U43696 (N_43696,N_43481,N_43429);
and U43697 (N_43697,N_43489,N_43499);
and U43698 (N_43698,N_43489,N_43295);
or U43699 (N_43699,N_43473,N_43407);
nand U43700 (N_43700,N_43485,N_43250);
nor U43701 (N_43701,N_43377,N_43322);
xor U43702 (N_43702,N_43348,N_43448);
nor U43703 (N_43703,N_43330,N_43490);
or U43704 (N_43704,N_43486,N_43250);
nor U43705 (N_43705,N_43381,N_43415);
xnor U43706 (N_43706,N_43259,N_43498);
or U43707 (N_43707,N_43390,N_43433);
or U43708 (N_43708,N_43472,N_43391);
nor U43709 (N_43709,N_43331,N_43317);
or U43710 (N_43710,N_43274,N_43453);
xnor U43711 (N_43711,N_43376,N_43330);
nor U43712 (N_43712,N_43454,N_43327);
or U43713 (N_43713,N_43394,N_43461);
xnor U43714 (N_43714,N_43486,N_43264);
xnor U43715 (N_43715,N_43260,N_43376);
and U43716 (N_43716,N_43435,N_43340);
nor U43717 (N_43717,N_43268,N_43275);
nand U43718 (N_43718,N_43458,N_43450);
xnor U43719 (N_43719,N_43438,N_43381);
or U43720 (N_43720,N_43410,N_43465);
and U43721 (N_43721,N_43474,N_43404);
or U43722 (N_43722,N_43474,N_43358);
nand U43723 (N_43723,N_43439,N_43376);
nor U43724 (N_43724,N_43274,N_43441);
nand U43725 (N_43725,N_43315,N_43403);
nand U43726 (N_43726,N_43271,N_43490);
and U43727 (N_43727,N_43389,N_43439);
or U43728 (N_43728,N_43389,N_43421);
nor U43729 (N_43729,N_43391,N_43437);
nand U43730 (N_43730,N_43366,N_43302);
nand U43731 (N_43731,N_43289,N_43369);
nand U43732 (N_43732,N_43278,N_43324);
and U43733 (N_43733,N_43469,N_43423);
and U43734 (N_43734,N_43417,N_43436);
nor U43735 (N_43735,N_43485,N_43438);
or U43736 (N_43736,N_43352,N_43274);
nor U43737 (N_43737,N_43278,N_43485);
nand U43738 (N_43738,N_43406,N_43299);
nand U43739 (N_43739,N_43340,N_43334);
nor U43740 (N_43740,N_43430,N_43394);
nor U43741 (N_43741,N_43404,N_43451);
nand U43742 (N_43742,N_43488,N_43450);
and U43743 (N_43743,N_43408,N_43461);
or U43744 (N_43744,N_43347,N_43452);
and U43745 (N_43745,N_43301,N_43400);
nand U43746 (N_43746,N_43428,N_43335);
nand U43747 (N_43747,N_43441,N_43360);
nor U43748 (N_43748,N_43413,N_43496);
or U43749 (N_43749,N_43274,N_43346);
xor U43750 (N_43750,N_43699,N_43509);
nand U43751 (N_43751,N_43595,N_43714);
and U43752 (N_43752,N_43706,N_43626);
xor U43753 (N_43753,N_43746,N_43650);
or U43754 (N_43754,N_43539,N_43597);
or U43755 (N_43755,N_43716,N_43729);
and U43756 (N_43756,N_43683,N_43669);
and U43757 (N_43757,N_43549,N_43512);
or U43758 (N_43758,N_43567,N_43543);
xnor U43759 (N_43759,N_43631,N_43644);
or U43760 (N_43760,N_43585,N_43579);
nand U43761 (N_43761,N_43704,N_43628);
nand U43762 (N_43762,N_43518,N_43531);
xor U43763 (N_43763,N_43500,N_43682);
nand U43764 (N_43764,N_43608,N_43603);
and U43765 (N_43765,N_43604,N_43665);
or U43766 (N_43766,N_43725,N_43510);
or U43767 (N_43767,N_43587,N_43679);
or U43768 (N_43768,N_43647,N_43642);
nand U43769 (N_43769,N_43618,N_43694);
and U43770 (N_43770,N_43554,N_43533);
and U43771 (N_43771,N_43505,N_43556);
and U43772 (N_43772,N_43600,N_43660);
and U43773 (N_43773,N_43632,N_43697);
xnor U43774 (N_43774,N_43717,N_43561);
xor U43775 (N_43775,N_43610,N_43601);
nor U43776 (N_43776,N_43503,N_43573);
or U43777 (N_43777,N_43559,N_43745);
nand U43778 (N_43778,N_43507,N_43506);
nand U43779 (N_43779,N_43649,N_43728);
nor U43780 (N_43780,N_43615,N_43655);
nor U43781 (N_43781,N_43582,N_43749);
xnor U43782 (N_43782,N_43688,N_43698);
and U43783 (N_43783,N_43707,N_43741);
nor U43784 (N_43784,N_43508,N_43619);
nand U43785 (N_43785,N_43593,N_43544);
nand U43786 (N_43786,N_43691,N_43566);
xnor U43787 (N_43787,N_43629,N_43547);
or U43788 (N_43788,N_43592,N_43633);
and U43789 (N_43789,N_43536,N_43726);
nand U43790 (N_43790,N_43526,N_43641);
nor U43791 (N_43791,N_43534,N_43670);
nor U43792 (N_43792,N_43620,N_43524);
nor U43793 (N_43793,N_43738,N_43684);
and U43794 (N_43794,N_43550,N_43545);
nand U43795 (N_43795,N_43519,N_43520);
or U43796 (N_43796,N_43546,N_43611);
or U43797 (N_43797,N_43614,N_43734);
nand U43798 (N_43798,N_43637,N_43577);
nand U43799 (N_43799,N_43564,N_43596);
nor U43800 (N_43800,N_43576,N_43695);
nor U43801 (N_43801,N_43646,N_43692);
nor U43802 (N_43802,N_43586,N_43677);
or U43803 (N_43803,N_43722,N_43661);
nand U43804 (N_43804,N_43624,N_43532);
xor U43805 (N_43805,N_43735,N_43668);
nand U43806 (N_43806,N_43676,N_43671);
xor U43807 (N_43807,N_43652,N_43718);
nor U43808 (N_43808,N_43720,N_43541);
or U43809 (N_43809,N_43733,N_43640);
nand U43810 (N_43810,N_43590,N_43687);
nor U43811 (N_43811,N_43622,N_43709);
xnor U43812 (N_43812,N_43574,N_43594);
and U43813 (N_43813,N_43680,N_43602);
nand U43814 (N_43814,N_43588,N_43638);
or U43815 (N_43815,N_43723,N_43690);
nand U43816 (N_43816,N_43571,N_43731);
nand U43817 (N_43817,N_43643,N_43748);
xor U43818 (N_43818,N_43538,N_43696);
nand U43819 (N_43819,N_43719,N_43739);
and U43820 (N_43820,N_43705,N_43740);
or U43821 (N_43821,N_43516,N_43607);
and U43822 (N_43822,N_43711,N_43648);
nand U43823 (N_43823,N_43672,N_43674);
or U43824 (N_43824,N_43627,N_43525);
xor U43825 (N_43825,N_43528,N_43659);
nand U43826 (N_43826,N_43701,N_43732);
and U43827 (N_43827,N_43630,N_43552);
xnor U43828 (N_43828,N_43744,N_43617);
xnor U43829 (N_43829,N_43708,N_43609);
nand U43830 (N_43830,N_43517,N_43657);
nor U43831 (N_43831,N_43555,N_43551);
xnor U43832 (N_43832,N_43639,N_43681);
nand U43833 (N_43833,N_43742,N_43664);
xor U43834 (N_43834,N_43580,N_43558);
or U43835 (N_43835,N_43712,N_43502);
and U43836 (N_43836,N_43521,N_43658);
xnor U43837 (N_43837,N_43540,N_43542);
or U43838 (N_43838,N_43702,N_43654);
nor U43839 (N_43839,N_43736,N_43584);
nor U43840 (N_43840,N_43730,N_43514);
nand U43841 (N_43841,N_43635,N_43727);
and U43842 (N_43842,N_43673,N_43569);
and U43843 (N_43843,N_43553,N_43651);
nor U43844 (N_43844,N_43737,N_43656);
nand U43845 (N_43845,N_43636,N_43606);
xnor U43846 (N_43846,N_43613,N_43621);
xor U43847 (N_43847,N_43666,N_43589);
xor U43848 (N_43848,N_43678,N_43599);
or U43849 (N_43849,N_43667,N_43572);
nor U43850 (N_43850,N_43616,N_43703);
and U43851 (N_43851,N_43548,N_43523);
nand U43852 (N_43852,N_43530,N_43689);
xnor U43853 (N_43853,N_43686,N_43625);
nand U43854 (N_43854,N_43747,N_43535);
nand U43855 (N_43855,N_43575,N_43562);
nand U43856 (N_43856,N_43713,N_43653);
xnor U43857 (N_43857,N_43700,N_43721);
nand U43858 (N_43858,N_43710,N_43570);
or U43859 (N_43859,N_43515,N_43605);
or U43860 (N_43860,N_43557,N_43578);
nor U43861 (N_43861,N_43724,N_43560);
nand U43862 (N_43862,N_43715,N_43598);
and U43863 (N_43863,N_43662,N_43623);
xnor U43864 (N_43864,N_43537,N_43513);
nand U43865 (N_43865,N_43565,N_43501);
nand U43866 (N_43866,N_43743,N_43529);
nand U43867 (N_43867,N_43693,N_43504);
nor U43868 (N_43868,N_43568,N_43612);
nand U43869 (N_43869,N_43591,N_43563);
xnor U43870 (N_43870,N_43583,N_43511);
or U43871 (N_43871,N_43685,N_43663);
nor U43872 (N_43872,N_43522,N_43581);
or U43873 (N_43873,N_43634,N_43645);
nand U43874 (N_43874,N_43527,N_43675);
nand U43875 (N_43875,N_43703,N_43626);
xnor U43876 (N_43876,N_43500,N_43720);
xor U43877 (N_43877,N_43689,N_43695);
and U43878 (N_43878,N_43513,N_43697);
and U43879 (N_43879,N_43512,N_43653);
and U43880 (N_43880,N_43621,N_43609);
or U43881 (N_43881,N_43536,N_43675);
and U43882 (N_43882,N_43507,N_43534);
xnor U43883 (N_43883,N_43529,N_43578);
or U43884 (N_43884,N_43683,N_43749);
nand U43885 (N_43885,N_43660,N_43672);
xor U43886 (N_43886,N_43628,N_43739);
and U43887 (N_43887,N_43736,N_43634);
nand U43888 (N_43888,N_43632,N_43690);
nand U43889 (N_43889,N_43704,N_43515);
and U43890 (N_43890,N_43694,N_43541);
nor U43891 (N_43891,N_43547,N_43656);
nand U43892 (N_43892,N_43533,N_43521);
and U43893 (N_43893,N_43551,N_43627);
nand U43894 (N_43894,N_43623,N_43610);
nor U43895 (N_43895,N_43578,N_43547);
or U43896 (N_43896,N_43616,N_43688);
nand U43897 (N_43897,N_43637,N_43545);
or U43898 (N_43898,N_43590,N_43677);
nor U43899 (N_43899,N_43653,N_43632);
or U43900 (N_43900,N_43581,N_43669);
and U43901 (N_43901,N_43629,N_43596);
nand U43902 (N_43902,N_43607,N_43670);
or U43903 (N_43903,N_43633,N_43739);
nand U43904 (N_43904,N_43618,N_43500);
and U43905 (N_43905,N_43636,N_43653);
nor U43906 (N_43906,N_43735,N_43672);
nor U43907 (N_43907,N_43715,N_43741);
and U43908 (N_43908,N_43706,N_43538);
nor U43909 (N_43909,N_43685,N_43749);
nand U43910 (N_43910,N_43675,N_43568);
xor U43911 (N_43911,N_43727,N_43676);
or U43912 (N_43912,N_43504,N_43588);
and U43913 (N_43913,N_43700,N_43647);
nor U43914 (N_43914,N_43700,N_43749);
and U43915 (N_43915,N_43701,N_43573);
and U43916 (N_43916,N_43739,N_43638);
and U43917 (N_43917,N_43739,N_43590);
xor U43918 (N_43918,N_43593,N_43603);
or U43919 (N_43919,N_43717,N_43734);
or U43920 (N_43920,N_43713,N_43613);
nor U43921 (N_43921,N_43555,N_43527);
or U43922 (N_43922,N_43561,N_43633);
nand U43923 (N_43923,N_43512,N_43545);
and U43924 (N_43924,N_43548,N_43580);
nand U43925 (N_43925,N_43558,N_43629);
nand U43926 (N_43926,N_43727,N_43743);
and U43927 (N_43927,N_43728,N_43505);
nor U43928 (N_43928,N_43627,N_43617);
nor U43929 (N_43929,N_43550,N_43677);
nand U43930 (N_43930,N_43540,N_43721);
nand U43931 (N_43931,N_43648,N_43677);
xor U43932 (N_43932,N_43505,N_43625);
nor U43933 (N_43933,N_43673,N_43738);
or U43934 (N_43934,N_43694,N_43512);
or U43935 (N_43935,N_43726,N_43719);
xor U43936 (N_43936,N_43500,N_43511);
nor U43937 (N_43937,N_43598,N_43596);
or U43938 (N_43938,N_43502,N_43740);
and U43939 (N_43939,N_43599,N_43624);
nor U43940 (N_43940,N_43598,N_43580);
nor U43941 (N_43941,N_43610,N_43715);
nand U43942 (N_43942,N_43647,N_43519);
or U43943 (N_43943,N_43604,N_43575);
nand U43944 (N_43944,N_43556,N_43619);
nor U43945 (N_43945,N_43525,N_43717);
nand U43946 (N_43946,N_43526,N_43651);
nor U43947 (N_43947,N_43744,N_43552);
or U43948 (N_43948,N_43668,N_43597);
or U43949 (N_43949,N_43616,N_43737);
nor U43950 (N_43950,N_43681,N_43705);
nand U43951 (N_43951,N_43594,N_43530);
and U43952 (N_43952,N_43729,N_43685);
and U43953 (N_43953,N_43537,N_43629);
nor U43954 (N_43954,N_43697,N_43739);
nor U43955 (N_43955,N_43521,N_43528);
nand U43956 (N_43956,N_43678,N_43721);
and U43957 (N_43957,N_43555,N_43742);
nor U43958 (N_43958,N_43660,N_43594);
nand U43959 (N_43959,N_43530,N_43683);
and U43960 (N_43960,N_43688,N_43538);
or U43961 (N_43961,N_43624,N_43629);
or U43962 (N_43962,N_43633,N_43677);
xnor U43963 (N_43963,N_43588,N_43546);
nor U43964 (N_43964,N_43714,N_43706);
xnor U43965 (N_43965,N_43724,N_43687);
nand U43966 (N_43966,N_43574,N_43619);
xor U43967 (N_43967,N_43707,N_43663);
and U43968 (N_43968,N_43712,N_43641);
and U43969 (N_43969,N_43733,N_43612);
or U43970 (N_43970,N_43609,N_43636);
or U43971 (N_43971,N_43572,N_43657);
xor U43972 (N_43972,N_43740,N_43537);
or U43973 (N_43973,N_43643,N_43629);
nor U43974 (N_43974,N_43667,N_43742);
xor U43975 (N_43975,N_43641,N_43604);
or U43976 (N_43976,N_43733,N_43586);
xor U43977 (N_43977,N_43513,N_43729);
nand U43978 (N_43978,N_43656,N_43728);
xnor U43979 (N_43979,N_43696,N_43521);
nor U43980 (N_43980,N_43552,N_43655);
nor U43981 (N_43981,N_43556,N_43512);
and U43982 (N_43982,N_43540,N_43652);
or U43983 (N_43983,N_43521,N_43669);
or U43984 (N_43984,N_43653,N_43682);
nand U43985 (N_43985,N_43610,N_43712);
nor U43986 (N_43986,N_43714,N_43596);
and U43987 (N_43987,N_43608,N_43596);
nand U43988 (N_43988,N_43690,N_43616);
nand U43989 (N_43989,N_43514,N_43558);
xor U43990 (N_43990,N_43526,N_43625);
nor U43991 (N_43991,N_43618,N_43535);
nor U43992 (N_43992,N_43520,N_43503);
and U43993 (N_43993,N_43655,N_43651);
and U43994 (N_43994,N_43678,N_43705);
xnor U43995 (N_43995,N_43544,N_43693);
and U43996 (N_43996,N_43582,N_43738);
or U43997 (N_43997,N_43662,N_43678);
xor U43998 (N_43998,N_43744,N_43682);
xor U43999 (N_43999,N_43596,N_43679);
or U44000 (N_44000,N_43828,N_43847);
or U44001 (N_44001,N_43993,N_43875);
and U44002 (N_44002,N_43787,N_43768);
and U44003 (N_44003,N_43939,N_43871);
xor U44004 (N_44004,N_43891,N_43852);
or U44005 (N_44005,N_43784,N_43892);
xor U44006 (N_44006,N_43864,N_43980);
nand U44007 (N_44007,N_43782,N_43918);
and U44008 (N_44008,N_43886,N_43913);
and U44009 (N_44009,N_43879,N_43857);
or U44010 (N_44010,N_43963,N_43862);
or U44011 (N_44011,N_43932,N_43758);
xnor U44012 (N_44012,N_43845,N_43856);
nor U44013 (N_44013,N_43813,N_43934);
xor U44014 (N_44014,N_43773,N_43830);
nand U44015 (N_44015,N_43770,N_43849);
and U44016 (N_44016,N_43945,N_43797);
xor U44017 (N_44017,N_43915,N_43834);
or U44018 (N_44018,N_43824,N_43759);
nand U44019 (N_44019,N_43844,N_43983);
nor U44020 (N_44020,N_43969,N_43948);
or U44021 (N_44021,N_43867,N_43793);
nor U44022 (N_44022,N_43978,N_43767);
nand U44023 (N_44023,N_43977,N_43974);
and U44024 (N_44024,N_43912,N_43893);
or U44025 (N_44025,N_43803,N_43971);
nor U44026 (N_44026,N_43794,N_43946);
xnor U44027 (N_44027,N_43851,N_43878);
xor U44028 (N_44028,N_43829,N_43827);
xnor U44029 (N_44029,N_43801,N_43788);
nor U44030 (N_44030,N_43930,N_43861);
nor U44031 (N_44031,N_43938,N_43883);
and U44032 (N_44032,N_43858,N_43988);
nor U44033 (N_44033,N_43968,N_43804);
or U44034 (N_44034,N_43761,N_43752);
and U44035 (N_44035,N_43868,N_43955);
nand U44036 (N_44036,N_43917,N_43760);
xor U44037 (N_44037,N_43973,N_43853);
nand U44038 (N_44038,N_43769,N_43967);
or U44039 (N_44039,N_43766,N_43956);
and U44040 (N_44040,N_43994,N_43890);
and U44041 (N_44041,N_43846,N_43818);
nor U44042 (N_44042,N_43810,N_43869);
or U44043 (N_44043,N_43914,N_43757);
and U44044 (N_44044,N_43970,N_43928);
xnor U44045 (N_44045,N_43925,N_43774);
or U44046 (N_44046,N_43841,N_43923);
or U44047 (N_44047,N_43833,N_43835);
nor U44048 (N_44048,N_43838,N_43962);
nand U44049 (N_44049,N_43790,N_43753);
nor U44050 (N_44050,N_43947,N_43935);
nand U44051 (N_44051,N_43999,N_43802);
or U44052 (N_44052,N_43959,N_43795);
xnor U44053 (N_44053,N_43985,N_43855);
and U44054 (N_44054,N_43942,N_43836);
nor U44055 (N_44055,N_43863,N_43800);
nand U44056 (N_44056,N_43992,N_43894);
nor U44057 (N_44057,N_43763,N_43922);
or U44058 (N_44058,N_43850,N_43771);
nor U44059 (N_44059,N_43958,N_43907);
nand U44060 (N_44060,N_43811,N_43839);
xor U44061 (N_44061,N_43940,N_43895);
nand U44062 (N_44062,N_43979,N_43924);
nand U44063 (N_44063,N_43825,N_43887);
or U44064 (N_44064,N_43872,N_43859);
and U44065 (N_44065,N_43807,N_43885);
nor U44066 (N_44066,N_43989,N_43920);
nand U44067 (N_44067,N_43780,N_43966);
nand U44068 (N_44068,N_43908,N_43911);
nand U44069 (N_44069,N_43888,N_43902);
nand U44070 (N_44070,N_43822,N_43909);
nand U44071 (N_44071,N_43900,N_43951);
nand U44072 (N_44072,N_43873,N_43789);
nand U44073 (N_44073,N_43821,N_43816);
nand U44074 (N_44074,N_43982,N_43882);
nor U44075 (N_44075,N_43901,N_43750);
or U44076 (N_44076,N_43984,N_43943);
nand U44077 (N_44077,N_43832,N_43843);
xor U44078 (N_44078,N_43903,N_43756);
or U44079 (N_44079,N_43754,N_43840);
xnor U44080 (N_44080,N_43772,N_43899);
nor U44081 (N_44081,N_43792,N_43937);
nand U44082 (N_44082,N_43781,N_43866);
nand U44083 (N_44083,N_43817,N_43929);
and U44084 (N_44084,N_43799,N_43927);
and U44085 (N_44085,N_43905,N_43876);
and U44086 (N_44086,N_43949,N_43916);
nand U44087 (N_44087,N_43953,N_43944);
or U44088 (N_44088,N_43775,N_43936);
xor U44089 (N_44089,N_43921,N_43889);
nor U44090 (N_44090,N_43897,N_43933);
xor U44091 (N_44091,N_43941,N_43964);
nand U44092 (N_44092,N_43884,N_43981);
and U44093 (N_44093,N_43910,N_43854);
xnor U44094 (N_44094,N_43874,N_43842);
or U44095 (N_44095,N_43786,N_43791);
or U44096 (N_44096,N_43976,N_43954);
nor U44097 (N_44097,N_43785,N_43991);
xor U44098 (N_44098,N_43877,N_43865);
nor U44099 (N_44099,N_43919,N_43820);
nand U44100 (N_44100,N_43765,N_43952);
nor U44101 (N_44101,N_43960,N_43798);
nand U44102 (N_44102,N_43931,N_43975);
and U44103 (N_44103,N_43805,N_43814);
xnor U44104 (N_44104,N_43831,N_43812);
or U44105 (N_44105,N_43796,N_43961);
nor U44106 (N_44106,N_43764,N_43860);
xor U44107 (N_44107,N_43819,N_43906);
nor U44108 (N_44108,N_43996,N_43778);
or U44109 (N_44109,N_43776,N_43870);
or U44110 (N_44110,N_43808,N_43990);
or U44111 (N_44111,N_43998,N_43777);
nand U44112 (N_44112,N_43779,N_43751);
nand U44113 (N_44113,N_43880,N_43995);
or U44114 (N_44114,N_43904,N_43986);
nand U44115 (N_44115,N_43815,N_43826);
and U44116 (N_44116,N_43997,N_43783);
or U44117 (N_44117,N_43809,N_43957);
nor U44118 (N_44118,N_43972,N_43881);
and U44119 (N_44119,N_43823,N_43755);
nor U44120 (N_44120,N_43926,N_43837);
and U44121 (N_44121,N_43950,N_43762);
or U44122 (N_44122,N_43965,N_43987);
or U44123 (N_44123,N_43848,N_43896);
nand U44124 (N_44124,N_43898,N_43806);
or U44125 (N_44125,N_43788,N_43970);
xor U44126 (N_44126,N_43920,N_43838);
or U44127 (N_44127,N_43943,N_43780);
nor U44128 (N_44128,N_43892,N_43949);
and U44129 (N_44129,N_43843,N_43752);
xnor U44130 (N_44130,N_43893,N_43925);
nor U44131 (N_44131,N_43871,N_43807);
and U44132 (N_44132,N_43944,N_43960);
xor U44133 (N_44133,N_43792,N_43804);
nand U44134 (N_44134,N_43876,N_43888);
nand U44135 (N_44135,N_43963,N_43884);
xor U44136 (N_44136,N_43841,N_43977);
nor U44137 (N_44137,N_43959,N_43780);
xnor U44138 (N_44138,N_43973,N_43911);
nand U44139 (N_44139,N_43858,N_43955);
and U44140 (N_44140,N_43793,N_43978);
or U44141 (N_44141,N_43983,N_43857);
xnor U44142 (N_44142,N_43972,N_43777);
xnor U44143 (N_44143,N_43989,N_43981);
or U44144 (N_44144,N_43990,N_43978);
xnor U44145 (N_44145,N_43855,N_43771);
nand U44146 (N_44146,N_43750,N_43920);
nor U44147 (N_44147,N_43915,N_43838);
nand U44148 (N_44148,N_43942,N_43814);
or U44149 (N_44149,N_43798,N_43876);
xor U44150 (N_44150,N_43977,N_43759);
or U44151 (N_44151,N_43874,N_43805);
and U44152 (N_44152,N_43949,N_43978);
nor U44153 (N_44153,N_43952,N_43967);
nor U44154 (N_44154,N_43816,N_43842);
nor U44155 (N_44155,N_43806,N_43997);
xor U44156 (N_44156,N_43849,N_43909);
xnor U44157 (N_44157,N_43865,N_43950);
nor U44158 (N_44158,N_43901,N_43828);
and U44159 (N_44159,N_43867,N_43846);
nand U44160 (N_44160,N_43797,N_43967);
or U44161 (N_44161,N_43751,N_43843);
nor U44162 (N_44162,N_43866,N_43919);
and U44163 (N_44163,N_43885,N_43765);
nand U44164 (N_44164,N_43791,N_43800);
or U44165 (N_44165,N_43900,N_43947);
and U44166 (N_44166,N_43824,N_43812);
or U44167 (N_44167,N_43915,N_43946);
nor U44168 (N_44168,N_43806,N_43950);
nand U44169 (N_44169,N_43994,N_43915);
or U44170 (N_44170,N_43835,N_43955);
and U44171 (N_44171,N_43977,N_43760);
nand U44172 (N_44172,N_43765,N_43828);
or U44173 (N_44173,N_43759,N_43819);
or U44174 (N_44174,N_43861,N_43773);
xor U44175 (N_44175,N_43824,N_43822);
xnor U44176 (N_44176,N_43970,N_43964);
xnor U44177 (N_44177,N_43811,N_43771);
and U44178 (N_44178,N_43978,N_43769);
nor U44179 (N_44179,N_43804,N_43815);
xnor U44180 (N_44180,N_43755,N_43900);
and U44181 (N_44181,N_43798,N_43984);
or U44182 (N_44182,N_43941,N_43989);
and U44183 (N_44183,N_43934,N_43872);
nand U44184 (N_44184,N_43949,N_43824);
or U44185 (N_44185,N_43842,N_43954);
nand U44186 (N_44186,N_43765,N_43777);
nor U44187 (N_44187,N_43983,N_43770);
nand U44188 (N_44188,N_43797,N_43923);
nand U44189 (N_44189,N_43787,N_43777);
xor U44190 (N_44190,N_43965,N_43827);
nor U44191 (N_44191,N_43784,N_43753);
and U44192 (N_44192,N_43825,N_43998);
nand U44193 (N_44193,N_43797,N_43758);
nand U44194 (N_44194,N_43783,N_43757);
and U44195 (N_44195,N_43947,N_43877);
nand U44196 (N_44196,N_43907,N_43942);
and U44197 (N_44197,N_43815,N_43949);
and U44198 (N_44198,N_43935,N_43865);
and U44199 (N_44199,N_43795,N_43755);
xor U44200 (N_44200,N_43808,N_43854);
nand U44201 (N_44201,N_43807,N_43987);
and U44202 (N_44202,N_43861,N_43958);
or U44203 (N_44203,N_43973,N_43922);
nand U44204 (N_44204,N_43887,N_43964);
and U44205 (N_44205,N_43781,N_43994);
nor U44206 (N_44206,N_43992,N_43830);
xor U44207 (N_44207,N_43903,N_43914);
or U44208 (N_44208,N_43925,N_43783);
nand U44209 (N_44209,N_43891,N_43788);
and U44210 (N_44210,N_43775,N_43979);
nand U44211 (N_44211,N_43887,N_43784);
nand U44212 (N_44212,N_43839,N_43907);
or U44213 (N_44213,N_43971,N_43860);
or U44214 (N_44214,N_43812,N_43773);
or U44215 (N_44215,N_43951,N_43781);
and U44216 (N_44216,N_43937,N_43934);
or U44217 (N_44217,N_43983,N_43831);
nor U44218 (N_44218,N_43778,N_43907);
or U44219 (N_44219,N_43836,N_43849);
nand U44220 (N_44220,N_43925,N_43852);
and U44221 (N_44221,N_43891,N_43923);
nand U44222 (N_44222,N_43810,N_43988);
xnor U44223 (N_44223,N_43945,N_43920);
and U44224 (N_44224,N_43795,N_43923);
or U44225 (N_44225,N_43853,N_43830);
or U44226 (N_44226,N_43844,N_43887);
nand U44227 (N_44227,N_43793,N_43824);
and U44228 (N_44228,N_43906,N_43829);
nor U44229 (N_44229,N_43782,N_43768);
nand U44230 (N_44230,N_43923,N_43855);
nand U44231 (N_44231,N_43920,N_43998);
or U44232 (N_44232,N_43801,N_43805);
or U44233 (N_44233,N_43814,N_43874);
and U44234 (N_44234,N_43802,N_43974);
nand U44235 (N_44235,N_43768,N_43757);
xor U44236 (N_44236,N_43910,N_43759);
and U44237 (N_44237,N_43853,N_43826);
or U44238 (N_44238,N_43780,N_43795);
xor U44239 (N_44239,N_43926,N_43839);
and U44240 (N_44240,N_43769,N_43966);
and U44241 (N_44241,N_43839,N_43876);
nand U44242 (N_44242,N_43992,N_43903);
xnor U44243 (N_44243,N_43911,N_43762);
or U44244 (N_44244,N_43852,N_43887);
and U44245 (N_44245,N_43875,N_43984);
and U44246 (N_44246,N_43916,N_43989);
and U44247 (N_44247,N_43906,N_43976);
xnor U44248 (N_44248,N_43921,N_43958);
nand U44249 (N_44249,N_43996,N_43852);
nand U44250 (N_44250,N_44122,N_44095);
and U44251 (N_44251,N_44008,N_44137);
or U44252 (N_44252,N_44035,N_44036);
xnor U44253 (N_44253,N_44163,N_44094);
or U44254 (N_44254,N_44105,N_44099);
xnor U44255 (N_44255,N_44040,N_44150);
or U44256 (N_44256,N_44239,N_44144);
nand U44257 (N_44257,N_44199,N_44077);
nor U44258 (N_44258,N_44217,N_44173);
nor U44259 (N_44259,N_44056,N_44073);
nand U44260 (N_44260,N_44195,N_44228);
nor U44261 (N_44261,N_44044,N_44067);
or U44262 (N_44262,N_44240,N_44219);
xnor U44263 (N_44263,N_44134,N_44127);
nor U44264 (N_44264,N_44103,N_44086);
and U44265 (N_44265,N_44019,N_44189);
xnor U44266 (N_44266,N_44182,N_44154);
nor U44267 (N_44267,N_44213,N_44112);
or U44268 (N_44268,N_44041,N_44212);
nand U44269 (N_44269,N_44031,N_44072);
xnor U44270 (N_44270,N_44235,N_44117);
and U44271 (N_44271,N_44175,N_44087);
or U44272 (N_44272,N_44032,N_44026);
or U44273 (N_44273,N_44216,N_44069);
nand U44274 (N_44274,N_44227,N_44045);
nor U44275 (N_44275,N_44047,N_44151);
nor U44276 (N_44276,N_44160,N_44021);
nand U44277 (N_44277,N_44104,N_44043);
xor U44278 (N_44278,N_44162,N_44057);
nand U44279 (N_44279,N_44243,N_44037);
nand U44280 (N_44280,N_44200,N_44135);
and U44281 (N_44281,N_44100,N_44140);
nand U44282 (N_44282,N_44145,N_44014);
nor U44283 (N_44283,N_44190,N_44169);
nand U44284 (N_44284,N_44060,N_44229);
or U44285 (N_44285,N_44245,N_44198);
xnor U44286 (N_44286,N_44159,N_44223);
or U44287 (N_44287,N_44197,N_44185);
nor U44288 (N_44288,N_44034,N_44064);
nor U44289 (N_44289,N_44158,N_44241);
nand U44290 (N_44290,N_44209,N_44186);
nand U44291 (N_44291,N_44106,N_44093);
and U44292 (N_44292,N_44123,N_44215);
nor U44293 (N_44293,N_44242,N_44115);
and U44294 (N_44294,N_44167,N_44079);
xnor U44295 (N_44295,N_44029,N_44184);
or U44296 (N_44296,N_44234,N_44078);
xor U44297 (N_44297,N_44054,N_44211);
nand U44298 (N_44298,N_44138,N_44085);
xnor U44299 (N_44299,N_44232,N_44132);
or U44300 (N_44300,N_44204,N_44023);
nand U44301 (N_44301,N_44187,N_44165);
or U44302 (N_44302,N_44124,N_44025);
nor U44303 (N_44303,N_44089,N_44218);
or U44304 (N_44304,N_44136,N_44226);
xor U44305 (N_44305,N_44166,N_44013);
nor U44306 (N_44306,N_44061,N_44074);
and U44307 (N_44307,N_44155,N_44237);
and U44308 (N_44308,N_44075,N_44107);
nor U44309 (N_44309,N_44101,N_44142);
xor U44310 (N_44310,N_44076,N_44005);
or U44311 (N_44311,N_44033,N_44083);
xor U44312 (N_44312,N_44148,N_44178);
xnor U44313 (N_44313,N_44068,N_44121);
xor U44314 (N_44314,N_44238,N_44066);
nand U44315 (N_44315,N_44020,N_44096);
nor U44316 (N_44316,N_44233,N_44088);
or U44317 (N_44317,N_44090,N_44003);
nand U44318 (N_44318,N_44156,N_44181);
or U44319 (N_44319,N_44125,N_44249);
and U44320 (N_44320,N_44000,N_44007);
nor U44321 (N_44321,N_44052,N_44153);
nor U44322 (N_44322,N_44131,N_44006);
or U44323 (N_44323,N_44147,N_44179);
or U44324 (N_44324,N_44161,N_44203);
nand U44325 (N_44325,N_44236,N_44022);
nor U44326 (N_44326,N_44063,N_44247);
nand U44327 (N_44327,N_44141,N_44002);
and U44328 (N_44328,N_44059,N_44126);
xor U44329 (N_44329,N_44224,N_44018);
or U44330 (N_44330,N_44050,N_44171);
xnor U44331 (N_44331,N_44174,N_44152);
and U44332 (N_44332,N_44177,N_44016);
or U44333 (N_44333,N_44201,N_44062);
nand U44334 (N_44334,N_44102,N_44012);
and U44335 (N_44335,N_44164,N_44128);
nor U44336 (N_44336,N_44039,N_44113);
nand U44337 (N_44337,N_44053,N_44004);
and U44338 (N_44338,N_44048,N_44098);
xor U44339 (N_44339,N_44028,N_44214);
or U44340 (N_44340,N_44130,N_44194);
or U44341 (N_44341,N_44065,N_44110);
or U44342 (N_44342,N_44172,N_44183);
nor U44343 (N_44343,N_44191,N_44027);
or U44344 (N_44344,N_44192,N_44092);
nor U44345 (N_44345,N_44210,N_44225);
or U44346 (N_44346,N_44149,N_44120);
or U44347 (N_44347,N_44111,N_44084);
xor U44348 (N_44348,N_44206,N_44009);
or U44349 (N_44349,N_44222,N_44097);
xnor U44350 (N_44350,N_44193,N_44082);
or U44351 (N_44351,N_44188,N_44119);
nor U44352 (N_44352,N_44030,N_44139);
xor U44353 (N_44353,N_44011,N_44080);
nand U44354 (N_44354,N_44205,N_44042);
xnor U44355 (N_44355,N_44116,N_44015);
or U44356 (N_44356,N_44133,N_44220);
or U44357 (N_44357,N_44046,N_44208);
and U44358 (N_44358,N_44114,N_44244);
nor U44359 (N_44359,N_44168,N_44049);
nand U44360 (N_44360,N_44109,N_44058);
or U44361 (N_44361,N_44108,N_44196);
or U44362 (N_44362,N_44051,N_44221);
xor U44363 (N_44363,N_44157,N_44146);
nor U44364 (N_44364,N_44001,N_44176);
and U44365 (N_44365,N_44017,N_44118);
and U44366 (N_44366,N_44129,N_44246);
xnor U44367 (N_44367,N_44024,N_44143);
nor U44368 (N_44368,N_44055,N_44230);
nand U44369 (N_44369,N_44070,N_44038);
and U44370 (N_44370,N_44091,N_44180);
nand U44371 (N_44371,N_44248,N_44010);
nor U44372 (N_44372,N_44081,N_44071);
or U44373 (N_44373,N_44170,N_44202);
xor U44374 (N_44374,N_44207,N_44231);
and U44375 (N_44375,N_44145,N_44155);
nor U44376 (N_44376,N_44085,N_44173);
xor U44377 (N_44377,N_44072,N_44150);
nor U44378 (N_44378,N_44225,N_44053);
and U44379 (N_44379,N_44002,N_44223);
and U44380 (N_44380,N_44142,N_44229);
and U44381 (N_44381,N_44159,N_44206);
xnor U44382 (N_44382,N_44155,N_44105);
nand U44383 (N_44383,N_44114,N_44208);
nand U44384 (N_44384,N_44072,N_44205);
nand U44385 (N_44385,N_44045,N_44188);
and U44386 (N_44386,N_44135,N_44128);
nor U44387 (N_44387,N_44013,N_44220);
or U44388 (N_44388,N_44195,N_44077);
and U44389 (N_44389,N_44225,N_44129);
and U44390 (N_44390,N_44076,N_44196);
nor U44391 (N_44391,N_44047,N_44239);
nand U44392 (N_44392,N_44106,N_44053);
and U44393 (N_44393,N_44114,N_44129);
or U44394 (N_44394,N_44036,N_44060);
xnor U44395 (N_44395,N_44210,N_44053);
nor U44396 (N_44396,N_44224,N_44085);
xor U44397 (N_44397,N_44077,N_44171);
nor U44398 (N_44398,N_44189,N_44170);
nor U44399 (N_44399,N_44177,N_44134);
nor U44400 (N_44400,N_44127,N_44210);
or U44401 (N_44401,N_44189,N_44076);
xnor U44402 (N_44402,N_44025,N_44127);
nand U44403 (N_44403,N_44130,N_44086);
xor U44404 (N_44404,N_44169,N_44132);
xor U44405 (N_44405,N_44120,N_44234);
and U44406 (N_44406,N_44243,N_44216);
xor U44407 (N_44407,N_44073,N_44116);
or U44408 (N_44408,N_44079,N_44055);
nand U44409 (N_44409,N_44163,N_44104);
nand U44410 (N_44410,N_44103,N_44137);
nand U44411 (N_44411,N_44229,N_44126);
and U44412 (N_44412,N_44024,N_44045);
xor U44413 (N_44413,N_44042,N_44166);
nand U44414 (N_44414,N_44047,N_44031);
nor U44415 (N_44415,N_44049,N_44210);
xnor U44416 (N_44416,N_44054,N_44084);
nor U44417 (N_44417,N_44239,N_44195);
xnor U44418 (N_44418,N_44113,N_44065);
nand U44419 (N_44419,N_44091,N_44239);
and U44420 (N_44420,N_44113,N_44211);
or U44421 (N_44421,N_44052,N_44040);
nand U44422 (N_44422,N_44169,N_44199);
or U44423 (N_44423,N_44116,N_44146);
and U44424 (N_44424,N_44243,N_44142);
or U44425 (N_44425,N_44093,N_44006);
nor U44426 (N_44426,N_44111,N_44117);
xnor U44427 (N_44427,N_44132,N_44158);
nor U44428 (N_44428,N_44200,N_44120);
or U44429 (N_44429,N_44169,N_44194);
or U44430 (N_44430,N_44205,N_44146);
or U44431 (N_44431,N_44205,N_44235);
or U44432 (N_44432,N_44215,N_44210);
or U44433 (N_44433,N_44131,N_44233);
and U44434 (N_44434,N_44241,N_44059);
nand U44435 (N_44435,N_44078,N_44149);
xnor U44436 (N_44436,N_44199,N_44168);
and U44437 (N_44437,N_44025,N_44136);
nor U44438 (N_44438,N_44107,N_44072);
or U44439 (N_44439,N_44157,N_44096);
nand U44440 (N_44440,N_44103,N_44105);
and U44441 (N_44441,N_44127,N_44191);
or U44442 (N_44442,N_44233,N_44119);
or U44443 (N_44443,N_44224,N_44064);
nand U44444 (N_44444,N_44109,N_44014);
xnor U44445 (N_44445,N_44122,N_44072);
xor U44446 (N_44446,N_44138,N_44232);
xnor U44447 (N_44447,N_44063,N_44091);
or U44448 (N_44448,N_44196,N_44058);
xnor U44449 (N_44449,N_44194,N_44244);
nor U44450 (N_44450,N_44092,N_44178);
xnor U44451 (N_44451,N_44083,N_44175);
or U44452 (N_44452,N_44009,N_44236);
and U44453 (N_44453,N_44018,N_44101);
nand U44454 (N_44454,N_44172,N_44115);
and U44455 (N_44455,N_44145,N_44243);
nand U44456 (N_44456,N_44010,N_44110);
xor U44457 (N_44457,N_44011,N_44127);
nor U44458 (N_44458,N_44000,N_44231);
nor U44459 (N_44459,N_44033,N_44216);
or U44460 (N_44460,N_44178,N_44108);
nor U44461 (N_44461,N_44040,N_44079);
xnor U44462 (N_44462,N_44220,N_44068);
or U44463 (N_44463,N_44063,N_44087);
and U44464 (N_44464,N_44001,N_44047);
or U44465 (N_44465,N_44200,N_44004);
xnor U44466 (N_44466,N_44070,N_44104);
nor U44467 (N_44467,N_44096,N_44195);
nand U44468 (N_44468,N_44043,N_44236);
and U44469 (N_44469,N_44142,N_44012);
xnor U44470 (N_44470,N_44180,N_44104);
or U44471 (N_44471,N_44127,N_44054);
and U44472 (N_44472,N_44174,N_44154);
nor U44473 (N_44473,N_44042,N_44181);
nand U44474 (N_44474,N_44107,N_44014);
or U44475 (N_44475,N_44231,N_44045);
or U44476 (N_44476,N_44192,N_44184);
xnor U44477 (N_44477,N_44032,N_44002);
and U44478 (N_44478,N_44052,N_44152);
or U44479 (N_44479,N_44039,N_44103);
nand U44480 (N_44480,N_44062,N_44022);
or U44481 (N_44481,N_44179,N_44063);
and U44482 (N_44482,N_44049,N_44234);
xnor U44483 (N_44483,N_44103,N_44116);
nor U44484 (N_44484,N_44101,N_44115);
nand U44485 (N_44485,N_44053,N_44089);
nor U44486 (N_44486,N_44230,N_44115);
nand U44487 (N_44487,N_44167,N_44205);
and U44488 (N_44488,N_44087,N_44124);
nand U44489 (N_44489,N_44000,N_44157);
and U44490 (N_44490,N_44014,N_44030);
and U44491 (N_44491,N_44232,N_44071);
and U44492 (N_44492,N_44049,N_44056);
nor U44493 (N_44493,N_44200,N_44091);
and U44494 (N_44494,N_44183,N_44180);
nor U44495 (N_44495,N_44035,N_44208);
nor U44496 (N_44496,N_44077,N_44017);
and U44497 (N_44497,N_44148,N_44077);
and U44498 (N_44498,N_44170,N_44198);
nand U44499 (N_44499,N_44034,N_44027);
nor U44500 (N_44500,N_44274,N_44457);
xnor U44501 (N_44501,N_44277,N_44458);
or U44502 (N_44502,N_44388,N_44473);
and U44503 (N_44503,N_44396,N_44304);
nor U44504 (N_44504,N_44346,N_44355);
nand U44505 (N_44505,N_44393,N_44257);
xnor U44506 (N_44506,N_44439,N_44498);
and U44507 (N_44507,N_44282,N_44333);
nor U44508 (N_44508,N_44496,N_44276);
xor U44509 (N_44509,N_44275,N_44329);
xnor U44510 (N_44510,N_44381,N_44459);
nand U44511 (N_44511,N_44464,N_44418);
nor U44512 (N_44512,N_44387,N_44408);
nor U44513 (N_44513,N_44309,N_44348);
nand U44514 (N_44514,N_44331,N_44443);
nor U44515 (N_44515,N_44343,N_44477);
or U44516 (N_44516,N_44420,N_44310);
and U44517 (N_44517,N_44373,N_44425);
and U44518 (N_44518,N_44287,N_44493);
and U44519 (N_44519,N_44261,N_44266);
or U44520 (N_44520,N_44295,N_44422);
xnor U44521 (N_44521,N_44273,N_44410);
xnor U44522 (N_44522,N_44340,N_44305);
nor U44523 (N_44523,N_44444,N_44474);
xnor U44524 (N_44524,N_44298,N_44369);
nand U44525 (N_44525,N_44398,N_44437);
nor U44526 (N_44526,N_44278,N_44446);
nor U44527 (N_44527,N_44460,N_44478);
and U44528 (N_44528,N_44349,N_44491);
nand U44529 (N_44529,N_44365,N_44389);
or U44530 (N_44530,N_44361,N_44302);
or U44531 (N_44531,N_44301,N_44354);
and U44532 (N_44532,N_44313,N_44484);
nand U44533 (N_44533,N_44258,N_44450);
or U44534 (N_44534,N_44378,N_44417);
or U44535 (N_44535,N_44463,N_44454);
and U44536 (N_44536,N_44337,N_44395);
or U44537 (N_44537,N_44462,N_44488);
xnor U44538 (N_44538,N_44400,N_44392);
xor U44539 (N_44539,N_44341,N_44441);
nor U44540 (N_44540,N_44289,N_44427);
and U44541 (N_44541,N_44359,N_44263);
nand U44542 (N_44542,N_44296,N_44468);
nor U44543 (N_44543,N_44481,N_44499);
and U44544 (N_44544,N_44353,N_44494);
nand U44545 (N_44545,N_44384,N_44428);
nand U44546 (N_44546,N_44344,N_44419);
xnor U44547 (N_44547,N_44345,N_44470);
nor U44548 (N_44548,N_44382,N_44267);
xnor U44549 (N_44549,N_44440,N_44367);
xor U44550 (N_44550,N_44442,N_44467);
or U44551 (N_44551,N_44405,N_44312);
or U44552 (N_44552,N_44351,N_44433);
nor U44553 (N_44553,N_44311,N_44307);
and U44554 (N_44554,N_44268,N_44317);
or U44555 (N_44555,N_44320,N_44436);
nand U44556 (N_44556,N_44448,N_44322);
xor U44557 (N_44557,N_44366,N_44326);
nor U44558 (N_44558,N_44291,N_44456);
nor U44559 (N_44559,N_44449,N_44487);
or U44560 (N_44560,N_44414,N_44330);
or U44561 (N_44561,N_44479,N_44283);
nor U44562 (N_44562,N_44285,N_44374);
or U44563 (N_44563,N_44306,N_44411);
nand U44564 (N_44564,N_44390,N_44380);
xnor U44565 (N_44565,N_44292,N_44471);
nand U44566 (N_44566,N_44371,N_44453);
nand U44567 (N_44567,N_44327,N_44492);
xor U44568 (N_44568,N_44251,N_44476);
nand U44569 (N_44569,N_44451,N_44397);
and U44570 (N_44570,N_44250,N_44391);
nand U44571 (N_44571,N_44497,N_44452);
or U44572 (N_44572,N_44426,N_44415);
xor U44573 (N_44573,N_44352,N_44407);
or U44574 (N_44574,N_44413,N_44315);
nand U44575 (N_44575,N_44466,N_44416);
xnor U44576 (N_44576,N_44447,N_44430);
xor U44577 (N_44577,N_44356,N_44265);
nor U44578 (N_44578,N_44338,N_44280);
nand U44579 (N_44579,N_44435,N_44429);
nor U44580 (N_44580,N_44256,N_44379);
nor U44581 (N_44581,N_44264,N_44303);
nor U44582 (N_44582,N_44421,N_44318);
nand U44583 (N_44583,N_44342,N_44368);
and U44584 (N_44584,N_44288,N_44297);
nand U44585 (N_44585,N_44423,N_44431);
xnor U44586 (N_44586,N_44269,N_44316);
or U44587 (N_44587,N_44461,N_44270);
and U44588 (N_44588,N_44386,N_44486);
xor U44589 (N_44589,N_44299,N_44253);
xnor U44590 (N_44590,N_44455,N_44360);
nand U44591 (N_44591,N_44482,N_44409);
or U44592 (N_44592,N_44321,N_44434);
and U44593 (N_44593,N_44485,N_44377);
or U44594 (N_44594,N_44332,N_44490);
xor U44595 (N_44595,N_44324,N_44293);
or U44596 (N_44596,N_44406,N_44336);
nand U44597 (N_44597,N_44475,N_44254);
xnor U44598 (N_44598,N_44372,N_44364);
or U44599 (N_44599,N_44358,N_44335);
and U44600 (N_44600,N_44383,N_44375);
and U44601 (N_44601,N_44271,N_44480);
nor U44602 (N_44602,N_44357,N_44432);
or U44603 (N_44603,N_44259,N_44403);
or U44604 (N_44604,N_44347,N_44376);
nor U44605 (N_44605,N_44394,N_44339);
nand U44606 (N_44606,N_44472,N_44300);
nand U44607 (N_44607,N_44286,N_44279);
nand U44608 (N_44608,N_44362,N_44363);
or U44609 (N_44609,N_44438,N_44281);
or U44610 (N_44610,N_44319,N_44404);
or U44611 (N_44611,N_44465,N_44350);
nor U44612 (N_44612,N_44424,N_44252);
nand U44613 (N_44613,N_44489,N_44325);
or U44614 (N_44614,N_44334,N_44370);
and U44615 (N_44615,N_44401,N_44469);
xor U44616 (N_44616,N_44260,N_44385);
nor U44617 (N_44617,N_44399,N_44323);
or U44618 (N_44618,N_44308,N_44483);
nand U44619 (N_44619,N_44272,N_44495);
nand U44620 (N_44620,N_44328,N_44262);
xor U44621 (N_44621,N_44255,N_44290);
nand U44622 (N_44622,N_44402,N_44314);
or U44623 (N_44623,N_44445,N_44284);
nand U44624 (N_44624,N_44294,N_44412);
nor U44625 (N_44625,N_44315,N_44370);
or U44626 (N_44626,N_44462,N_44323);
or U44627 (N_44627,N_44427,N_44331);
nand U44628 (N_44628,N_44449,N_44260);
nor U44629 (N_44629,N_44252,N_44440);
and U44630 (N_44630,N_44488,N_44497);
nand U44631 (N_44631,N_44410,N_44433);
and U44632 (N_44632,N_44388,N_44313);
nand U44633 (N_44633,N_44473,N_44256);
or U44634 (N_44634,N_44397,N_44338);
xnor U44635 (N_44635,N_44433,N_44471);
nor U44636 (N_44636,N_44310,N_44410);
and U44637 (N_44637,N_44348,N_44409);
nand U44638 (N_44638,N_44356,N_44407);
nor U44639 (N_44639,N_44307,N_44446);
nand U44640 (N_44640,N_44307,N_44414);
nor U44641 (N_44641,N_44274,N_44470);
nand U44642 (N_44642,N_44262,N_44495);
nand U44643 (N_44643,N_44293,N_44365);
nand U44644 (N_44644,N_44310,N_44274);
or U44645 (N_44645,N_44455,N_44439);
nor U44646 (N_44646,N_44338,N_44439);
nor U44647 (N_44647,N_44487,N_44491);
and U44648 (N_44648,N_44383,N_44386);
xnor U44649 (N_44649,N_44419,N_44408);
xor U44650 (N_44650,N_44405,N_44305);
xnor U44651 (N_44651,N_44392,N_44440);
xor U44652 (N_44652,N_44304,N_44351);
or U44653 (N_44653,N_44458,N_44368);
xor U44654 (N_44654,N_44449,N_44274);
or U44655 (N_44655,N_44457,N_44492);
nand U44656 (N_44656,N_44252,N_44331);
and U44657 (N_44657,N_44410,N_44342);
xor U44658 (N_44658,N_44417,N_44399);
or U44659 (N_44659,N_44363,N_44412);
or U44660 (N_44660,N_44255,N_44344);
nand U44661 (N_44661,N_44337,N_44312);
nand U44662 (N_44662,N_44424,N_44321);
nand U44663 (N_44663,N_44405,N_44383);
nor U44664 (N_44664,N_44292,N_44421);
xnor U44665 (N_44665,N_44284,N_44483);
nand U44666 (N_44666,N_44339,N_44276);
nand U44667 (N_44667,N_44364,N_44392);
xnor U44668 (N_44668,N_44480,N_44352);
and U44669 (N_44669,N_44320,N_44288);
and U44670 (N_44670,N_44356,N_44258);
or U44671 (N_44671,N_44255,N_44279);
or U44672 (N_44672,N_44332,N_44406);
xor U44673 (N_44673,N_44453,N_44279);
nor U44674 (N_44674,N_44413,N_44433);
and U44675 (N_44675,N_44398,N_44390);
xor U44676 (N_44676,N_44424,N_44255);
nand U44677 (N_44677,N_44341,N_44427);
or U44678 (N_44678,N_44415,N_44340);
nor U44679 (N_44679,N_44348,N_44482);
nand U44680 (N_44680,N_44273,N_44260);
xnor U44681 (N_44681,N_44392,N_44264);
and U44682 (N_44682,N_44438,N_44447);
and U44683 (N_44683,N_44295,N_44447);
xnor U44684 (N_44684,N_44250,N_44354);
nand U44685 (N_44685,N_44317,N_44344);
nor U44686 (N_44686,N_44342,N_44313);
nand U44687 (N_44687,N_44356,N_44289);
and U44688 (N_44688,N_44496,N_44410);
and U44689 (N_44689,N_44290,N_44456);
nor U44690 (N_44690,N_44421,N_44305);
nand U44691 (N_44691,N_44370,N_44375);
nor U44692 (N_44692,N_44327,N_44400);
or U44693 (N_44693,N_44358,N_44437);
or U44694 (N_44694,N_44320,N_44428);
and U44695 (N_44695,N_44437,N_44266);
xor U44696 (N_44696,N_44363,N_44409);
nand U44697 (N_44697,N_44480,N_44359);
or U44698 (N_44698,N_44311,N_44407);
nor U44699 (N_44699,N_44271,N_44455);
and U44700 (N_44700,N_44408,N_44497);
xnor U44701 (N_44701,N_44452,N_44253);
nor U44702 (N_44702,N_44491,N_44272);
or U44703 (N_44703,N_44455,N_44365);
xnor U44704 (N_44704,N_44475,N_44387);
nor U44705 (N_44705,N_44254,N_44257);
and U44706 (N_44706,N_44329,N_44450);
nand U44707 (N_44707,N_44427,N_44457);
xnor U44708 (N_44708,N_44430,N_44496);
and U44709 (N_44709,N_44424,N_44352);
or U44710 (N_44710,N_44496,N_44351);
nand U44711 (N_44711,N_44409,N_44424);
nor U44712 (N_44712,N_44421,N_44389);
or U44713 (N_44713,N_44298,N_44302);
nand U44714 (N_44714,N_44338,N_44385);
nor U44715 (N_44715,N_44377,N_44435);
and U44716 (N_44716,N_44475,N_44352);
xnor U44717 (N_44717,N_44472,N_44278);
nor U44718 (N_44718,N_44365,N_44326);
or U44719 (N_44719,N_44368,N_44444);
nand U44720 (N_44720,N_44298,N_44362);
xnor U44721 (N_44721,N_44407,N_44499);
xnor U44722 (N_44722,N_44488,N_44252);
and U44723 (N_44723,N_44395,N_44416);
nand U44724 (N_44724,N_44349,N_44316);
nand U44725 (N_44725,N_44458,N_44325);
or U44726 (N_44726,N_44341,N_44474);
and U44727 (N_44727,N_44400,N_44476);
or U44728 (N_44728,N_44487,N_44460);
nand U44729 (N_44729,N_44406,N_44420);
or U44730 (N_44730,N_44313,N_44399);
nand U44731 (N_44731,N_44467,N_44455);
and U44732 (N_44732,N_44338,N_44389);
nand U44733 (N_44733,N_44465,N_44378);
and U44734 (N_44734,N_44321,N_44480);
xnor U44735 (N_44735,N_44455,N_44282);
xnor U44736 (N_44736,N_44323,N_44276);
and U44737 (N_44737,N_44450,N_44295);
and U44738 (N_44738,N_44439,N_44251);
and U44739 (N_44739,N_44466,N_44293);
xnor U44740 (N_44740,N_44421,N_44368);
nor U44741 (N_44741,N_44479,N_44340);
nand U44742 (N_44742,N_44486,N_44264);
nor U44743 (N_44743,N_44388,N_44307);
or U44744 (N_44744,N_44287,N_44443);
nand U44745 (N_44745,N_44363,N_44498);
xnor U44746 (N_44746,N_44257,N_44455);
and U44747 (N_44747,N_44395,N_44421);
xor U44748 (N_44748,N_44420,N_44376);
nor U44749 (N_44749,N_44392,N_44317);
or U44750 (N_44750,N_44702,N_44568);
or U44751 (N_44751,N_44683,N_44526);
xor U44752 (N_44752,N_44689,N_44728);
nor U44753 (N_44753,N_44679,N_44600);
xnor U44754 (N_44754,N_44532,N_44536);
nand U44755 (N_44755,N_44601,N_44732);
or U44756 (N_44756,N_44572,N_44593);
xnor U44757 (N_44757,N_44517,N_44652);
or U44758 (N_44758,N_44725,N_44576);
or U44759 (N_44759,N_44610,N_44554);
or U44760 (N_44760,N_44705,N_44509);
and U44761 (N_44761,N_44710,N_44715);
or U44762 (N_44762,N_44606,N_44579);
or U44763 (N_44763,N_44604,N_44574);
nand U44764 (N_44764,N_44546,N_44567);
nand U44765 (N_44765,N_44558,N_44621);
or U44766 (N_44766,N_44588,N_44748);
nor U44767 (N_44767,N_44680,N_44739);
and U44768 (N_44768,N_44659,N_44687);
nand U44769 (N_44769,N_44556,N_44584);
and U44770 (N_44770,N_44592,N_44605);
nand U44771 (N_44771,N_44667,N_44632);
or U44772 (N_44772,N_44587,N_44607);
or U44773 (N_44773,N_44562,N_44653);
nor U44774 (N_44774,N_44553,N_44525);
nor U44775 (N_44775,N_44520,N_44696);
nand U44776 (N_44776,N_44531,N_44620);
xor U44777 (N_44777,N_44528,N_44668);
xor U44778 (N_44778,N_44665,N_44586);
nor U44779 (N_44779,N_44743,N_44717);
nand U44780 (N_44780,N_44565,N_44590);
nand U44781 (N_44781,N_44618,N_44640);
and U44782 (N_44782,N_44540,N_44548);
xor U44783 (N_44783,N_44631,N_44662);
xor U44784 (N_44784,N_44542,N_44523);
and U44785 (N_44785,N_44639,N_44619);
nor U44786 (N_44786,N_44514,N_44693);
nor U44787 (N_44787,N_44697,N_44564);
and U44788 (N_44788,N_44711,N_44518);
and U44789 (N_44789,N_44596,N_44660);
or U44790 (N_44790,N_44651,N_44527);
or U44791 (N_44791,N_44718,N_44716);
and U44792 (N_44792,N_44740,N_44714);
or U44793 (N_44793,N_44649,N_44581);
and U44794 (N_44794,N_44585,N_44577);
nand U44795 (N_44795,N_44747,N_44661);
and U44796 (N_44796,N_44583,N_44547);
xor U44797 (N_44797,N_44676,N_44549);
xor U44798 (N_44798,N_44684,N_44641);
nand U44799 (N_44799,N_44603,N_44742);
xnor U44800 (N_44800,N_44686,N_44628);
nand U44801 (N_44801,N_44681,N_44695);
nor U44802 (N_44802,N_44543,N_44623);
nor U44803 (N_44803,N_44597,N_44522);
nor U44804 (N_44804,N_44612,N_44589);
nand U44805 (N_44805,N_44704,N_44736);
nor U44806 (N_44806,N_44741,N_44580);
nor U44807 (N_44807,N_44730,N_44550);
and U44808 (N_44808,N_44537,N_44723);
and U44809 (N_44809,N_44719,N_44595);
xor U44810 (N_44810,N_44529,N_44734);
xnor U44811 (N_44811,N_44638,N_44534);
and U44812 (N_44812,N_44654,N_44677);
nor U44813 (N_44813,N_44643,N_44658);
or U44814 (N_44814,N_44615,N_44663);
xor U44815 (N_44815,N_44608,N_44678);
nand U44816 (N_44816,N_44670,N_44506);
nor U44817 (N_44817,N_44647,N_44512);
and U44818 (N_44818,N_44671,N_44707);
nand U44819 (N_44819,N_44625,N_44648);
nor U44820 (N_44820,N_44629,N_44561);
xor U44821 (N_44821,N_44505,N_44692);
or U44822 (N_44822,N_44613,N_44735);
nor U44823 (N_44823,N_44669,N_44573);
xnor U44824 (N_44824,N_44519,N_44566);
nand U44825 (N_44825,N_44511,N_44733);
nor U44826 (N_44826,N_44570,N_44644);
nor U44827 (N_44827,N_44578,N_44555);
nand U44828 (N_44828,N_44616,N_44657);
and U44829 (N_44829,N_44535,N_44617);
nand U44830 (N_44830,N_44666,N_44501);
nor U44831 (N_44831,N_44557,N_44709);
or U44832 (N_44832,N_44521,N_44571);
or U44833 (N_44833,N_44591,N_44552);
nor U44834 (N_44834,N_44722,N_44599);
nor U44835 (N_44835,N_44515,N_44626);
nor U44836 (N_44836,N_44624,N_44682);
or U44837 (N_44837,N_44611,N_44563);
nand U44838 (N_44838,N_44672,N_44614);
nand U44839 (N_44839,N_44721,N_44706);
or U44840 (N_44840,N_44694,N_44720);
nand U44841 (N_44841,N_44634,N_44630);
nand U44842 (N_44842,N_44701,N_44646);
and U44843 (N_44843,N_44602,N_44575);
nand U44844 (N_44844,N_44691,N_44622);
nor U44845 (N_44845,N_44675,N_44727);
and U44846 (N_44846,N_44745,N_44533);
nand U44847 (N_44847,N_44656,N_44504);
nor U44848 (N_44848,N_44664,N_44636);
and U44849 (N_44849,N_44642,N_44738);
nor U44850 (N_44850,N_44545,N_44541);
nand U44851 (N_44851,N_44516,N_44713);
nand U44852 (N_44852,N_44530,N_44685);
and U44853 (N_44853,N_44544,N_44729);
xor U44854 (N_44854,N_44635,N_44560);
nor U44855 (N_44855,N_44650,N_44724);
nor U44856 (N_44856,N_44712,N_44538);
or U44857 (N_44857,N_44645,N_44627);
xnor U44858 (N_44858,N_44513,N_44569);
nand U44859 (N_44859,N_44539,N_44703);
nand U44860 (N_44860,N_44744,N_44609);
nor U44861 (N_44861,N_44633,N_44690);
and U44862 (N_44862,N_44500,N_44594);
and U44863 (N_44863,N_44746,N_44559);
xnor U44864 (N_44864,N_44698,N_44737);
and U44865 (N_44865,N_44502,N_44551);
nand U44866 (N_44866,N_44524,N_44708);
or U44867 (N_44867,N_44655,N_44688);
and U44868 (N_44868,N_44674,N_44673);
xor U44869 (N_44869,N_44582,N_44749);
nor U44870 (N_44870,N_44598,N_44510);
xor U44871 (N_44871,N_44637,N_44731);
xnor U44872 (N_44872,N_44508,N_44503);
nand U44873 (N_44873,N_44700,N_44699);
or U44874 (N_44874,N_44507,N_44726);
or U44875 (N_44875,N_44589,N_44650);
nand U44876 (N_44876,N_44700,N_44591);
or U44877 (N_44877,N_44595,N_44576);
nand U44878 (N_44878,N_44600,N_44500);
nor U44879 (N_44879,N_44710,N_44507);
nor U44880 (N_44880,N_44558,N_44670);
nand U44881 (N_44881,N_44680,N_44531);
or U44882 (N_44882,N_44557,N_44692);
xnor U44883 (N_44883,N_44543,N_44589);
or U44884 (N_44884,N_44695,N_44722);
nand U44885 (N_44885,N_44712,N_44739);
nand U44886 (N_44886,N_44621,N_44605);
and U44887 (N_44887,N_44737,N_44544);
xor U44888 (N_44888,N_44683,N_44657);
and U44889 (N_44889,N_44619,N_44666);
nor U44890 (N_44890,N_44541,N_44643);
and U44891 (N_44891,N_44722,N_44605);
or U44892 (N_44892,N_44634,N_44576);
or U44893 (N_44893,N_44730,N_44706);
and U44894 (N_44894,N_44735,N_44586);
nand U44895 (N_44895,N_44722,N_44577);
or U44896 (N_44896,N_44708,N_44680);
and U44897 (N_44897,N_44714,N_44718);
nor U44898 (N_44898,N_44638,N_44581);
or U44899 (N_44899,N_44606,N_44709);
xor U44900 (N_44900,N_44544,N_44555);
and U44901 (N_44901,N_44645,N_44702);
nand U44902 (N_44902,N_44588,N_44505);
or U44903 (N_44903,N_44554,N_44616);
or U44904 (N_44904,N_44655,N_44518);
nor U44905 (N_44905,N_44744,N_44707);
and U44906 (N_44906,N_44680,N_44509);
nor U44907 (N_44907,N_44629,N_44746);
nand U44908 (N_44908,N_44536,N_44709);
and U44909 (N_44909,N_44549,N_44743);
nand U44910 (N_44910,N_44695,N_44562);
xnor U44911 (N_44911,N_44512,N_44737);
and U44912 (N_44912,N_44589,N_44637);
nand U44913 (N_44913,N_44723,N_44510);
nor U44914 (N_44914,N_44542,N_44571);
nand U44915 (N_44915,N_44514,N_44599);
nor U44916 (N_44916,N_44734,N_44633);
and U44917 (N_44917,N_44547,N_44619);
or U44918 (N_44918,N_44726,N_44691);
or U44919 (N_44919,N_44674,N_44620);
xor U44920 (N_44920,N_44713,N_44669);
nor U44921 (N_44921,N_44591,N_44587);
and U44922 (N_44922,N_44748,N_44623);
and U44923 (N_44923,N_44709,N_44574);
nand U44924 (N_44924,N_44668,N_44516);
or U44925 (N_44925,N_44542,N_44525);
nand U44926 (N_44926,N_44701,N_44744);
and U44927 (N_44927,N_44647,N_44530);
nand U44928 (N_44928,N_44654,N_44571);
nor U44929 (N_44929,N_44570,N_44663);
or U44930 (N_44930,N_44610,N_44685);
nand U44931 (N_44931,N_44740,N_44629);
and U44932 (N_44932,N_44519,N_44734);
and U44933 (N_44933,N_44574,N_44515);
xnor U44934 (N_44934,N_44728,N_44701);
nand U44935 (N_44935,N_44628,N_44554);
xnor U44936 (N_44936,N_44608,N_44665);
nor U44937 (N_44937,N_44674,N_44529);
or U44938 (N_44938,N_44685,N_44725);
and U44939 (N_44939,N_44651,N_44518);
nand U44940 (N_44940,N_44650,N_44648);
nor U44941 (N_44941,N_44595,N_44744);
xor U44942 (N_44942,N_44576,N_44558);
and U44943 (N_44943,N_44683,N_44682);
or U44944 (N_44944,N_44544,N_44671);
or U44945 (N_44945,N_44634,N_44538);
xor U44946 (N_44946,N_44660,N_44656);
nand U44947 (N_44947,N_44637,N_44560);
xor U44948 (N_44948,N_44510,N_44686);
xnor U44949 (N_44949,N_44716,N_44514);
nand U44950 (N_44950,N_44561,N_44539);
xor U44951 (N_44951,N_44705,N_44565);
nand U44952 (N_44952,N_44635,N_44723);
xor U44953 (N_44953,N_44626,N_44516);
nand U44954 (N_44954,N_44535,N_44722);
nor U44955 (N_44955,N_44525,N_44692);
nand U44956 (N_44956,N_44528,N_44714);
nor U44957 (N_44957,N_44612,N_44619);
nor U44958 (N_44958,N_44657,N_44726);
xor U44959 (N_44959,N_44586,N_44502);
xor U44960 (N_44960,N_44629,N_44708);
nand U44961 (N_44961,N_44645,N_44678);
and U44962 (N_44962,N_44705,N_44503);
nor U44963 (N_44963,N_44649,N_44673);
or U44964 (N_44964,N_44700,N_44728);
or U44965 (N_44965,N_44673,N_44660);
nor U44966 (N_44966,N_44724,N_44631);
or U44967 (N_44967,N_44663,N_44672);
nor U44968 (N_44968,N_44686,N_44673);
or U44969 (N_44969,N_44638,N_44641);
or U44970 (N_44970,N_44627,N_44728);
nand U44971 (N_44971,N_44745,N_44585);
xnor U44972 (N_44972,N_44683,N_44705);
nor U44973 (N_44973,N_44518,N_44576);
or U44974 (N_44974,N_44618,N_44716);
nor U44975 (N_44975,N_44640,N_44728);
and U44976 (N_44976,N_44581,N_44663);
xor U44977 (N_44977,N_44655,N_44683);
or U44978 (N_44978,N_44526,N_44647);
nor U44979 (N_44979,N_44582,N_44524);
nand U44980 (N_44980,N_44619,N_44702);
xor U44981 (N_44981,N_44638,N_44649);
or U44982 (N_44982,N_44515,N_44571);
and U44983 (N_44983,N_44609,N_44671);
nand U44984 (N_44984,N_44682,N_44727);
nor U44985 (N_44985,N_44578,N_44738);
or U44986 (N_44986,N_44658,N_44697);
nor U44987 (N_44987,N_44693,N_44713);
and U44988 (N_44988,N_44739,N_44603);
xnor U44989 (N_44989,N_44550,N_44652);
nand U44990 (N_44990,N_44589,N_44603);
or U44991 (N_44991,N_44737,N_44703);
nor U44992 (N_44992,N_44503,N_44669);
nor U44993 (N_44993,N_44737,N_44669);
nor U44994 (N_44994,N_44652,N_44634);
nand U44995 (N_44995,N_44630,N_44736);
nand U44996 (N_44996,N_44634,N_44715);
xor U44997 (N_44997,N_44545,N_44530);
and U44998 (N_44998,N_44686,N_44551);
or U44999 (N_44999,N_44533,N_44685);
nor U45000 (N_45000,N_44771,N_44956);
or U45001 (N_45001,N_44849,N_44850);
xor U45002 (N_45002,N_44803,N_44962);
xor U45003 (N_45003,N_44780,N_44930);
and U45004 (N_45004,N_44934,N_44901);
nor U45005 (N_45005,N_44801,N_44983);
nor U45006 (N_45006,N_44835,N_44790);
nand U45007 (N_45007,N_44991,N_44958);
nor U45008 (N_45008,N_44856,N_44777);
and U45009 (N_45009,N_44989,N_44758);
or U45010 (N_45010,N_44907,N_44815);
xnor U45011 (N_45011,N_44865,N_44751);
nor U45012 (N_45012,N_44951,N_44939);
xnor U45013 (N_45013,N_44887,N_44757);
and U45014 (N_45014,N_44840,N_44832);
and U45015 (N_45015,N_44903,N_44820);
or U45016 (N_45016,N_44769,N_44954);
and U45017 (N_45017,N_44784,N_44898);
or U45018 (N_45018,N_44935,N_44948);
and U45019 (N_45019,N_44817,N_44911);
xor U45020 (N_45020,N_44816,N_44848);
nand U45021 (N_45021,N_44897,N_44885);
nor U45022 (N_45022,N_44767,N_44896);
and U45023 (N_45023,N_44957,N_44860);
nand U45024 (N_45024,N_44905,N_44988);
or U45025 (N_45025,N_44838,N_44900);
nand U45026 (N_45026,N_44852,N_44833);
or U45027 (N_45027,N_44812,N_44967);
or U45028 (N_45028,N_44764,N_44982);
and U45029 (N_45029,N_44807,N_44936);
nor U45030 (N_45030,N_44760,N_44893);
or U45031 (N_45031,N_44914,N_44974);
xor U45032 (N_45032,N_44789,N_44793);
and U45033 (N_45033,N_44808,N_44968);
nand U45034 (N_45034,N_44920,N_44891);
or U45035 (N_45035,N_44762,N_44965);
nor U45036 (N_45036,N_44794,N_44834);
nor U45037 (N_45037,N_44821,N_44964);
nand U45038 (N_45038,N_44750,N_44972);
and U45039 (N_45039,N_44824,N_44944);
and U45040 (N_45040,N_44785,N_44980);
xnor U45041 (N_45041,N_44947,N_44768);
nand U45042 (N_45042,N_44997,N_44960);
nand U45043 (N_45043,N_44828,N_44846);
nor U45044 (N_45044,N_44858,N_44950);
and U45045 (N_45045,N_44831,N_44880);
nor U45046 (N_45046,N_44921,N_44875);
xnor U45047 (N_45047,N_44864,N_44919);
nor U45048 (N_45048,N_44773,N_44895);
nor U45049 (N_45049,N_44863,N_44753);
or U45050 (N_45050,N_44873,N_44952);
or U45051 (N_45051,N_44841,N_44899);
xor U45052 (N_45052,N_44942,N_44839);
nor U45053 (N_45053,N_44862,N_44995);
xnor U45054 (N_45054,N_44929,N_44867);
nor U45055 (N_45055,N_44906,N_44979);
xor U45056 (N_45056,N_44937,N_44869);
or U45057 (N_45057,N_44940,N_44759);
nor U45058 (N_45058,N_44910,N_44798);
or U45059 (N_45059,N_44998,N_44969);
xor U45060 (N_45060,N_44872,N_44933);
nand U45061 (N_45061,N_44826,N_44804);
or U45062 (N_45062,N_44772,N_44908);
and U45063 (N_45063,N_44992,N_44822);
xnor U45064 (N_45064,N_44763,N_44961);
nor U45065 (N_45065,N_44938,N_44941);
nor U45066 (N_45066,N_44986,N_44836);
nand U45067 (N_45067,N_44859,N_44851);
xor U45068 (N_45068,N_44970,N_44778);
nor U45069 (N_45069,N_44868,N_44829);
nand U45070 (N_45070,N_44978,N_44928);
nor U45071 (N_45071,N_44857,N_44999);
nor U45072 (N_45072,N_44976,N_44915);
nor U45073 (N_45073,N_44966,N_44902);
nor U45074 (N_45074,N_44913,N_44878);
nor U45075 (N_45075,N_44830,N_44809);
nand U45076 (N_45076,N_44977,N_44925);
and U45077 (N_45077,N_44870,N_44783);
and U45078 (N_45078,N_44927,N_44802);
and U45079 (N_45079,N_44877,N_44752);
or U45080 (N_45080,N_44797,N_44883);
and U45081 (N_45081,N_44892,N_44882);
or U45082 (N_45082,N_44909,N_44792);
nand U45083 (N_45083,N_44786,N_44886);
xor U45084 (N_45084,N_44782,N_44827);
nand U45085 (N_45085,N_44781,N_44795);
and U45086 (N_45086,N_44990,N_44926);
or U45087 (N_45087,N_44791,N_44818);
nand U45088 (N_45088,N_44963,N_44814);
xnor U45089 (N_45089,N_44844,N_44973);
and U45090 (N_45090,N_44861,N_44775);
xnor U45091 (N_45091,N_44923,N_44955);
xor U45092 (N_45092,N_44842,N_44922);
nor U45093 (N_45093,N_44853,N_44806);
xnor U45094 (N_45094,N_44805,N_44949);
xnor U45095 (N_45095,N_44774,N_44984);
xnor U45096 (N_45096,N_44912,N_44994);
nor U45097 (N_45097,N_44787,N_44871);
nand U45098 (N_45098,N_44971,N_44766);
xor U45099 (N_45099,N_44981,N_44931);
and U45100 (N_45100,N_44888,N_44917);
and U45101 (N_45101,N_44776,N_44854);
nor U45102 (N_45102,N_44985,N_44975);
and U45103 (N_45103,N_44945,N_44996);
and U45104 (N_45104,N_44845,N_44765);
or U45105 (N_45105,N_44770,N_44924);
nor U45106 (N_45106,N_44987,N_44855);
xnor U45107 (N_45107,N_44953,N_44959);
nand U45108 (N_45108,N_44946,N_44918);
and U45109 (N_45109,N_44819,N_44823);
and U45110 (N_45110,N_44810,N_44788);
and U45111 (N_45111,N_44876,N_44890);
or U45112 (N_45112,N_44943,N_44884);
nand U45113 (N_45113,N_44813,N_44796);
xor U45114 (N_45114,N_44811,N_44866);
nor U45115 (N_45115,N_44800,N_44874);
and U45116 (N_45116,N_44837,N_44889);
nor U45117 (N_45117,N_44761,N_44754);
xor U45118 (N_45118,N_44881,N_44932);
and U45119 (N_45119,N_44799,N_44904);
or U45120 (N_45120,N_44779,N_44847);
and U45121 (N_45121,N_44993,N_44879);
xnor U45122 (N_45122,N_44916,N_44755);
xor U45123 (N_45123,N_44843,N_44894);
xor U45124 (N_45124,N_44825,N_44756);
or U45125 (N_45125,N_44951,N_44959);
nand U45126 (N_45126,N_44895,N_44919);
xnor U45127 (N_45127,N_44867,N_44838);
and U45128 (N_45128,N_44915,N_44823);
nor U45129 (N_45129,N_44833,N_44950);
and U45130 (N_45130,N_44826,N_44786);
xnor U45131 (N_45131,N_44910,N_44912);
nand U45132 (N_45132,N_44868,N_44896);
nor U45133 (N_45133,N_44824,N_44871);
nand U45134 (N_45134,N_44877,N_44946);
or U45135 (N_45135,N_44952,N_44827);
and U45136 (N_45136,N_44756,N_44791);
xnor U45137 (N_45137,N_44955,N_44972);
or U45138 (N_45138,N_44890,N_44790);
nand U45139 (N_45139,N_44844,N_44793);
and U45140 (N_45140,N_44972,N_44894);
xor U45141 (N_45141,N_44796,N_44883);
and U45142 (N_45142,N_44888,N_44839);
or U45143 (N_45143,N_44849,N_44918);
nand U45144 (N_45144,N_44803,N_44888);
and U45145 (N_45145,N_44978,N_44842);
nand U45146 (N_45146,N_44915,N_44975);
xnor U45147 (N_45147,N_44900,N_44876);
and U45148 (N_45148,N_44807,N_44771);
or U45149 (N_45149,N_44800,N_44917);
or U45150 (N_45150,N_44774,N_44822);
xnor U45151 (N_45151,N_44902,N_44818);
nor U45152 (N_45152,N_44934,N_44892);
and U45153 (N_45153,N_44801,N_44871);
or U45154 (N_45154,N_44945,N_44934);
and U45155 (N_45155,N_44989,N_44803);
nor U45156 (N_45156,N_44991,N_44797);
and U45157 (N_45157,N_44990,N_44820);
and U45158 (N_45158,N_44832,N_44910);
nand U45159 (N_45159,N_44910,N_44896);
and U45160 (N_45160,N_44766,N_44864);
xor U45161 (N_45161,N_44891,N_44955);
xnor U45162 (N_45162,N_44816,N_44977);
or U45163 (N_45163,N_44789,N_44970);
or U45164 (N_45164,N_44896,N_44948);
and U45165 (N_45165,N_44939,N_44772);
nand U45166 (N_45166,N_44906,N_44921);
or U45167 (N_45167,N_44788,N_44752);
nor U45168 (N_45168,N_44980,N_44916);
nand U45169 (N_45169,N_44805,N_44819);
nand U45170 (N_45170,N_44884,N_44958);
or U45171 (N_45171,N_44961,N_44835);
nor U45172 (N_45172,N_44974,N_44764);
xor U45173 (N_45173,N_44829,N_44770);
nor U45174 (N_45174,N_44957,N_44804);
nand U45175 (N_45175,N_44884,N_44767);
nor U45176 (N_45176,N_44807,N_44954);
and U45177 (N_45177,N_44969,N_44836);
or U45178 (N_45178,N_44968,N_44810);
xor U45179 (N_45179,N_44873,N_44871);
nand U45180 (N_45180,N_44821,N_44969);
and U45181 (N_45181,N_44886,N_44978);
nor U45182 (N_45182,N_44811,N_44883);
nor U45183 (N_45183,N_44991,N_44796);
nor U45184 (N_45184,N_44800,N_44962);
nor U45185 (N_45185,N_44757,N_44937);
nor U45186 (N_45186,N_44975,N_44779);
xnor U45187 (N_45187,N_44980,N_44838);
nor U45188 (N_45188,N_44877,N_44842);
or U45189 (N_45189,N_44925,N_44910);
xnor U45190 (N_45190,N_44891,N_44778);
xor U45191 (N_45191,N_44937,N_44956);
or U45192 (N_45192,N_44942,N_44751);
and U45193 (N_45193,N_44841,N_44764);
and U45194 (N_45194,N_44910,N_44983);
or U45195 (N_45195,N_44995,N_44940);
and U45196 (N_45196,N_44751,N_44826);
or U45197 (N_45197,N_44760,N_44817);
nand U45198 (N_45198,N_44839,N_44772);
xor U45199 (N_45199,N_44811,N_44886);
and U45200 (N_45200,N_44793,N_44817);
xor U45201 (N_45201,N_44988,N_44834);
nand U45202 (N_45202,N_44782,N_44786);
or U45203 (N_45203,N_44809,N_44934);
nand U45204 (N_45204,N_44995,N_44765);
nand U45205 (N_45205,N_44970,N_44779);
or U45206 (N_45206,N_44924,N_44826);
nor U45207 (N_45207,N_44944,N_44885);
xnor U45208 (N_45208,N_44886,N_44857);
xor U45209 (N_45209,N_44994,N_44806);
or U45210 (N_45210,N_44969,N_44863);
nor U45211 (N_45211,N_44889,N_44982);
and U45212 (N_45212,N_44850,N_44822);
and U45213 (N_45213,N_44779,N_44943);
xor U45214 (N_45214,N_44932,N_44798);
nand U45215 (N_45215,N_44934,N_44974);
and U45216 (N_45216,N_44860,N_44772);
or U45217 (N_45217,N_44969,N_44897);
or U45218 (N_45218,N_44756,N_44905);
nand U45219 (N_45219,N_44818,N_44908);
nand U45220 (N_45220,N_44775,N_44949);
or U45221 (N_45221,N_44794,N_44932);
and U45222 (N_45222,N_44837,N_44897);
or U45223 (N_45223,N_44778,N_44976);
nor U45224 (N_45224,N_44988,N_44895);
nand U45225 (N_45225,N_44921,N_44972);
or U45226 (N_45226,N_44960,N_44814);
xor U45227 (N_45227,N_44913,N_44859);
or U45228 (N_45228,N_44793,N_44883);
nand U45229 (N_45229,N_44974,N_44838);
xnor U45230 (N_45230,N_44854,N_44784);
xor U45231 (N_45231,N_44911,N_44851);
nor U45232 (N_45232,N_44895,N_44917);
and U45233 (N_45233,N_44829,N_44821);
and U45234 (N_45234,N_44928,N_44855);
nor U45235 (N_45235,N_44767,N_44934);
nand U45236 (N_45236,N_44754,N_44830);
nand U45237 (N_45237,N_44853,N_44802);
nor U45238 (N_45238,N_44755,N_44825);
and U45239 (N_45239,N_44890,N_44943);
nor U45240 (N_45240,N_44931,N_44800);
nand U45241 (N_45241,N_44845,N_44853);
xnor U45242 (N_45242,N_44827,N_44786);
or U45243 (N_45243,N_44848,N_44962);
and U45244 (N_45244,N_44857,N_44980);
xor U45245 (N_45245,N_44848,N_44859);
or U45246 (N_45246,N_44773,N_44955);
nor U45247 (N_45247,N_44914,N_44820);
nand U45248 (N_45248,N_44778,N_44800);
nor U45249 (N_45249,N_44825,N_44797);
nand U45250 (N_45250,N_45155,N_45075);
nor U45251 (N_45251,N_45096,N_45182);
and U45252 (N_45252,N_45143,N_45063);
and U45253 (N_45253,N_45059,N_45227);
nand U45254 (N_45254,N_45161,N_45231);
xnor U45255 (N_45255,N_45127,N_45093);
nor U45256 (N_45256,N_45171,N_45049);
nand U45257 (N_45257,N_45176,N_45151);
xor U45258 (N_45258,N_45000,N_45104);
nand U45259 (N_45259,N_45193,N_45056);
and U45260 (N_45260,N_45244,N_45240);
nand U45261 (N_45261,N_45236,N_45062);
xnor U45262 (N_45262,N_45027,N_45140);
nor U45263 (N_45263,N_45030,N_45011);
xnor U45264 (N_45264,N_45195,N_45068);
or U45265 (N_45265,N_45054,N_45088);
nor U45266 (N_45266,N_45098,N_45239);
and U45267 (N_45267,N_45097,N_45095);
and U45268 (N_45268,N_45100,N_45103);
nor U45269 (N_45269,N_45246,N_45142);
nand U45270 (N_45270,N_45058,N_45150);
nand U45271 (N_45271,N_45043,N_45067);
and U45272 (N_45272,N_45038,N_45078);
xnor U45273 (N_45273,N_45119,N_45156);
xor U45274 (N_45274,N_45123,N_45218);
xnor U45275 (N_45275,N_45225,N_45069);
nor U45276 (N_45276,N_45124,N_45133);
and U45277 (N_45277,N_45178,N_45209);
or U45278 (N_45278,N_45114,N_45175);
or U45279 (N_45279,N_45129,N_45180);
or U45280 (N_45280,N_45145,N_45061);
nand U45281 (N_45281,N_45048,N_45020);
or U45282 (N_45282,N_45091,N_45102);
xnor U45283 (N_45283,N_45122,N_45237);
and U45284 (N_45284,N_45118,N_45066);
xor U45285 (N_45285,N_45014,N_45206);
xor U45286 (N_45286,N_45041,N_45031);
nand U45287 (N_45287,N_45163,N_45029);
xor U45288 (N_45288,N_45057,N_45212);
xor U45289 (N_45289,N_45198,N_45099);
xor U45290 (N_45290,N_45016,N_45185);
nand U45291 (N_45291,N_45036,N_45044);
and U45292 (N_45292,N_45089,N_45189);
nor U45293 (N_45293,N_45019,N_45247);
or U45294 (N_45294,N_45033,N_45208);
nand U45295 (N_45295,N_45039,N_45169);
or U45296 (N_45296,N_45073,N_45232);
nand U45297 (N_45297,N_45235,N_45139);
nor U45298 (N_45298,N_45170,N_45224);
and U45299 (N_45299,N_45008,N_45165);
and U45300 (N_45300,N_45147,N_45108);
nor U45301 (N_45301,N_45005,N_45092);
and U45302 (N_45302,N_45221,N_45132);
nor U45303 (N_45303,N_45172,N_45110);
nand U45304 (N_45304,N_45077,N_45112);
and U45305 (N_45305,N_45245,N_45157);
xnor U45306 (N_45306,N_45186,N_45130);
and U45307 (N_45307,N_45074,N_45146);
nor U45308 (N_45308,N_45002,N_45177);
or U45309 (N_45309,N_45148,N_45022);
xor U45310 (N_45310,N_45080,N_45120);
or U45311 (N_45311,N_45040,N_45107);
nor U45312 (N_45312,N_45051,N_45128);
or U45313 (N_45313,N_45179,N_45183);
nor U45314 (N_45314,N_45081,N_45234);
nand U45315 (N_45315,N_45187,N_45013);
nor U45316 (N_45316,N_45135,N_45079);
xnor U45317 (N_45317,N_45228,N_45154);
xor U45318 (N_45318,N_45162,N_45060);
or U45319 (N_45319,N_45160,N_45085);
nor U45320 (N_45320,N_45047,N_45070);
nand U45321 (N_45321,N_45199,N_45113);
or U45322 (N_45322,N_45149,N_45249);
nand U45323 (N_45323,N_45076,N_45217);
nand U45324 (N_45324,N_45190,N_45134);
xor U45325 (N_45325,N_45213,N_45201);
xnor U45326 (N_45326,N_45012,N_45037);
or U45327 (N_45327,N_45086,N_45238);
nor U45328 (N_45328,N_45084,N_45050);
xnor U45329 (N_45329,N_45072,N_45001);
nor U45330 (N_45330,N_45222,N_45215);
xor U45331 (N_45331,N_45010,N_45055);
and U45332 (N_45332,N_45087,N_45025);
xor U45333 (N_45333,N_45211,N_45064);
or U45334 (N_45334,N_45153,N_45184);
nand U45335 (N_45335,N_45106,N_45216);
and U45336 (N_45336,N_45094,N_45115);
and U45337 (N_45337,N_45028,N_45131);
nand U45338 (N_45338,N_45017,N_45023);
and U45339 (N_45339,N_45125,N_45181);
or U45340 (N_45340,N_45109,N_45045);
nor U45341 (N_45341,N_45082,N_45152);
xor U45342 (N_45342,N_45226,N_45210);
and U45343 (N_45343,N_45242,N_45003);
or U45344 (N_45344,N_45083,N_45046);
or U45345 (N_45345,N_45009,N_45053);
nor U45346 (N_45346,N_45144,N_45233);
nand U45347 (N_45347,N_45071,N_45035);
nand U45348 (N_45348,N_45200,N_45243);
nor U45349 (N_45349,N_45241,N_45214);
and U45350 (N_45350,N_45158,N_45204);
or U45351 (N_45351,N_45202,N_45164);
xor U45352 (N_45352,N_45174,N_45101);
and U45353 (N_45353,N_45141,N_45117);
or U45354 (N_45354,N_45126,N_45024);
and U45355 (N_45355,N_45026,N_45137);
nor U45356 (N_45356,N_45229,N_45015);
or U45357 (N_45357,N_45223,N_45166);
nor U45358 (N_45358,N_45052,N_45136);
xnor U45359 (N_45359,N_45220,N_45197);
xor U45360 (N_45360,N_45065,N_45203);
xnor U45361 (N_45361,N_45105,N_45207);
xor U45362 (N_45362,N_45194,N_45196);
or U45363 (N_45363,N_45219,N_45021);
and U45364 (N_45364,N_45192,N_45034);
or U45365 (N_45365,N_45191,N_45188);
nor U45366 (N_45366,N_45032,N_45018);
nand U45367 (N_45367,N_45205,N_45121);
nand U45368 (N_45368,N_45138,N_45173);
and U45369 (N_45369,N_45159,N_45007);
xor U45370 (N_45370,N_45042,N_45116);
or U45371 (N_45371,N_45167,N_45168);
nor U45372 (N_45372,N_45248,N_45004);
nand U45373 (N_45373,N_45230,N_45090);
nor U45374 (N_45374,N_45006,N_45111);
or U45375 (N_45375,N_45168,N_45111);
nor U45376 (N_45376,N_45187,N_45118);
nand U45377 (N_45377,N_45020,N_45149);
nor U45378 (N_45378,N_45220,N_45212);
xor U45379 (N_45379,N_45134,N_45205);
and U45380 (N_45380,N_45190,N_45088);
xnor U45381 (N_45381,N_45188,N_45068);
or U45382 (N_45382,N_45222,N_45060);
nor U45383 (N_45383,N_45090,N_45216);
nor U45384 (N_45384,N_45101,N_45049);
nor U45385 (N_45385,N_45227,N_45022);
xor U45386 (N_45386,N_45067,N_45227);
nor U45387 (N_45387,N_45104,N_45215);
nand U45388 (N_45388,N_45034,N_45031);
nand U45389 (N_45389,N_45056,N_45131);
nand U45390 (N_45390,N_45226,N_45070);
and U45391 (N_45391,N_45046,N_45222);
nand U45392 (N_45392,N_45045,N_45067);
nand U45393 (N_45393,N_45111,N_45157);
and U45394 (N_45394,N_45229,N_45032);
xor U45395 (N_45395,N_45001,N_45130);
or U45396 (N_45396,N_45147,N_45082);
or U45397 (N_45397,N_45169,N_45194);
nand U45398 (N_45398,N_45139,N_45006);
nor U45399 (N_45399,N_45210,N_45201);
nand U45400 (N_45400,N_45242,N_45238);
nor U45401 (N_45401,N_45235,N_45044);
xor U45402 (N_45402,N_45021,N_45064);
or U45403 (N_45403,N_45144,N_45141);
nor U45404 (N_45404,N_45115,N_45236);
or U45405 (N_45405,N_45027,N_45102);
and U45406 (N_45406,N_45186,N_45116);
nor U45407 (N_45407,N_45097,N_45098);
nand U45408 (N_45408,N_45068,N_45205);
or U45409 (N_45409,N_45163,N_45024);
nand U45410 (N_45410,N_45224,N_45064);
nand U45411 (N_45411,N_45153,N_45240);
xor U45412 (N_45412,N_45074,N_45247);
nand U45413 (N_45413,N_45055,N_45077);
xor U45414 (N_45414,N_45240,N_45105);
and U45415 (N_45415,N_45212,N_45062);
and U45416 (N_45416,N_45185,N_45078);
xor U45417 (N_45417,N_45065,N_45148);
nand U45418 (N_45418,N_45212,N_45003);
xnor U45419 (N_45419,N_45127,N_45068);
xnor U45420 (N_45420,N_45018,N_45122);
nor U45421 (N_45421,N_45022,N_45033);
nand U45422 (N_45422,N_45241,N_45168);
nand U45423 (N_45423,N_45178,N_45122);
xor U45424 (N_45424,N_45158,N_45081);
nand U45425 (N_45425,N_45145,N_45241);
or U45426 (N_45426,N_45055,N_45151);
nand U45427 (N_45427,N_45047,N_45187);
or U45428 (N_45428,N_45195,N_45055);
xnor U45429 (N_45429,N_45087,N_45209);
nand U45430 (N_45430,N_45065,N_45242);
and U45431 (N_45431,N_45044,N_45227);
or U45432 (N_45432,N_45059,N_45066);
nor U45433 (N_45433,N_45077,N_45118);
nand U45434 (N_45434,N_45078,N_45207);
or U45435 (N_45435,N_45123,N_45118);
and U45436 (N_45436,N_45212,N_45221);
nand U45437 (N_45437,N_45007,N_45169);
nor U45438 (N_45438,N_45039,N_45179);
and U45439 (N_45439,N_45055,N_45013);
xor U45440 (N_45440,N_45052,N_45121);
xor U45441 (N_45441,N_45163,N_45104);
xnor U45442 (N_45442,N_45074,N_45085);
or U45443 (N_45443,N_45161,N_45103);
or U45444 (N_45444,N_45213,N_45018);
or U45445 (N_45445,N_45241,N_45046);
nor U45446 (N_45446,N_45025,N_45061);
nor U45447 (N_45447,N_45096,N_45017);
xnor U45448 (N_45448,N_45212,N_45069);
or U45449 (N_45449,N_45149,N_45030);
nand U45450 (N_45450,N_45111,N_45047);
and U45451 (N_45451,N_45132,N_45068);
nor U45452 (N_45452,N_45041,N_45070);
or U45453 (N_45453,N_45059,N_45047);
nor U45454 (N_45454,N_45206,N_45162);
nand U45455 (N_45455,N_45143,N_45102);
nand U45456 (N_45456,N_45116,N_45151);
xnor U45457 (N_45457,N_45067,N_45170);
nor U45458 (N_45458,N_45082,N_45158);
or U45459 (N_45459,N_45200,N_45076);
or U45460 (N_45460,N_45190,N_45050);
nand U45461 (N_45461,N_45095,N_45046);
nand U45462 (N_45462,N_45237,N_45057);
and U45463 (N_45463,N_45036,N_45128);
nand U45464 (N_45464,N_45109,N_45190);
or U45465 (N_45465,N_45111,N_45046);
or U45466 (N_45466,N_45174,N_45089);
nor U45467 (N_45467,N_45234,N_45194);
xnor U45468 (N_45468,N_45147,N_45077);
xor U45469 (N_45469,N_45008,N_45078);
nor U45470 (N_45470,N_45182,N_45198);
nor U45471 (N_45471,N_45104,N_45141);
and U45472 (N_45472,N_45063,N_45180);
nor U45473 (N_45473,N_45184,N_45210);
nand U45474 (N_45474,N_45097,N_45118);
or U45475 (N_45475,N_45044,N_45015);
and U45476 (N_45476,N_45140,N_45093);
xor U45477 (N_45477,N_45111,N_45010);
nand U45478 (N_45478,N_45166,N_45178);
or U45479 (N_45479,N_45233,N_45028);
or U45480 (N_45480,N_45193,N_45192);
and U45481 (N_45481,N_45239,N_45086);
nor U45482 (N_45482,N_45198,N_45183);
nor U45483 (N_45483,N_45035,N_45110);
and U45484 (N_45484,N_45174,N_45014);
and U45485 (N_45485,N_45013,N_45212);
nor U45486 (N_45486,N_45134,N_45046);
and U45487 (N_45487,N_45223,N_45077);
nor U45488 (N_45488,N_45085,N_45070);
nor U45489 (N_45489,N_45154,N_45041);
nor U45490 (N_45490,N_45164,N_45206);
xnor U45491 (N_45491,N_45193,N_45068);
or U45492 (N_45492,N_45099,N_45240);
and U45493 (N_45493,N_45218,N_45053);
xor U45494 (N_45494,N_45134,N_45135);
and U45495 (N_45495,N_45204,N_45176);
xor U45496 (N_45496,N_45036,N_45057);
nor U45497 (N_45497,N_45165,N_45162);
or U45498 (N_45498,N_45020,N_45090);
nor U45499 (N_45499,N_45188,N_45058);
xor U45500 (N_45500,N_45423,N_45256);
xor U45501 (N_45501,N_45355,N_45454);
nand U45502 (N_45502,N_45318,N_45384);
nor U45503 (N_45503,N_45349,N_45329);
or U45504 (N_45504,N_45331,N_45417);
xnor U45505 (N_45505,N_45413,N_45484);
and U45506 (N_45506,N_45451,N_45481);
or U45507 (N_45507,N_45492,N_45358);
xnor U45508 (N_45508,N_45493,N_45496);
or U45509 (N_45509,N_45469,N_45411);
or U45510 (N_45510,N_45498,N_45401);
nand U45511 (N_45511,N_45323,N_45332);
xnor U45512 (N_45512,N_45370,N_45379);
or U45513 (N_45513,N_45425,N_45457);
nand U45514 (N_45514,N_45404,N_45347);
nor U45515 (N_45515,N_45278,N_45385);
and U45516 (N_45516,N_45488,N_45475);
or U45517 (N_45517,N_45486,N_45434);
nor U45518 (N_45518,N_45298,N_45452);
nor U45519 (N_45519,N_45325,N_45461);
or U45520 (N_45520,N_45357,N_45302);
or U45521 (N_45521,N_45383,N_45261);
nand U45522 (N_45522,N_45435,N_45443);
or U45523 (N_45523,N_45395,N_45415);
nor U45524 (N_45524,N_45303,N_45499);
and U45525 (N_45525,N_45436,N_45408);
nand U45526 (N_45526,N_45263,N_45269);
nand U45527 (N_45527,N_45271,N_45444);
xnor U45528 (N_45528,N_45262,N_45348);
nand U45529 (N_45529,N_45316,N_45440);
and U45530 (N_45530,N_45466,N_45346);
xnor U45531 (N_45531,N_45448,N_45367);
and U45532 (N_45532,N_45251,N_45343);
or U45533 (N_45533,N_45283,N_45429);
and U45534 (N_45534,N_45468,N_45427);
nor U45535 (N_45535,N_45458,N_45338);
and U45536 (N_45536,N_45313,N_45356);
and U45537 (N_45537,N_45477,N_45396);
xnor U45538 (N_45538,N_45365,N_45490);
nand U45539 (N_45539,N_45467,N_45340);
or U45540 (N_45540,N_45437,N_45254);
and U45541 (N_45541,N_45321,N_45482);
or U45542 (N_45542,N_45288,N_45293);
nand U45543 (N_45543,N_45366,N_45259);
nand U45544 (N_45544,N_45315,N_45300);
and U45545 (N_45545,N_45352,N_45373);
and U45546 (N_45546,N_45497,N_45433);
and U45547 (N_45547,N_45409,N_45460);
xnor U45548 (N_45548,N_45465,N_45334);
and U45549 (N_45549,N_45277,N_45491);
nor U45550 (N_45550,N_45473,N_45445);
nand U45551 (N_45551,N_45374,N_45361);
or U45552 (N_45552,N_45264,N_45418);
nand U45553 (N_45553,N_45431,N_45462);
xor U45554 (N_45554,N_45380,N_45474);
or U45555 (N_45555,N_45324,N_45397);
nand U45556 (N_45556,N_45412,N_45489);
or U45557 (N_45557,N_45399,N_45398);
xor U45558 (N_45558,N_45414,N_45341);
nand U45559 (N_45559,N_45319,N_45459);
xnor U45560 (N_45560,N_45472,N_45387);
or U45561 (N_45561,N_45279,N_45297);
nor U45562 (N_45562,N_45339,N_45270);
xor U45563 (N_45563,N_45394,N_45291);
nand U45564 (N_45564,N_45406,N_45426);
xor U45565 (N_45565,N_45268,N_45280);
or U45566 (N_45566,N_45450,N_45393);
nand U45567 (N_45567,N_45378,N_45281);
or U45568 (N_45568,N_45287,N_45369);
nor U45569 (N_45569,N_45336,N_45307);
and U45570 (N_45570,N_45483,N_45267);
or U45571 (N_45571,N_45308,N_45344);
or U45572 (N_45572,N_45284,N_45351);
and U45573 (N_45573,N_45273,N_45400);
nand U45574 (N_45574,N_45446,N_45416);
nor U45575 (N_45575,N_45363,N_45337);
and U45576 (N_45576,N_45388,N_45449);
and U45577 (N_45577,N_45342,N_45455);
and U45578 (N_45578,N_45391,N_45402);
and U45579 (N_45579,N_45295,N_45276);
and U45580 (N_45580,N_45260,N_45392);
or U45581 (N_45581,N_45381,N_45330);
xnor U45582 (N_45582,N_45403,N_45432);
xor U45583 (N_45583,N_45453,N_45447);
nand U45584 (N_45584,N_45377,N_45422);
nor U45585 (N_45585,N_45290,N_45304);
or U45586 (N_45586,N_45255,N_45258);
xor U45587 (N_45587,N_45311,N_45353);
nand U45588 (N_45588,N_45257,N_45487);
nand U45589 (N_45589,N_45350,N_45345);
or U45590 (N_45590,N_45372,N_45424);
xor U45591 (N_45591,N_45275,N_45296);
nand U45592 (N_45592,N_45428,N_45320);
xor U45593 (N_45593,N_45478,N_45360);
nand U45594 (N_45594,N_45368,N_45252);
and U45595 (N_45595,N_45274,N_45327);
nand U45596 (N_45596,N_45289,N_45407);
or U45597 (N_45597,N_45463,N_45305);
nor U45598 (N_45598,N_45326,N_45476);
nor U45599 (N_45599,N_45285,N_45354);
nand U45600 (N_45600,N_45362,N_45494);
xnor U45601 (N_45601,N_45333,N_45410);
xor U45602 (N_45602,N_45282,N_45470);
xor U45603 (N_45603,N_45438,N_45389);
xor U45604 (N_45604,N_45382,N_45420);
nand U45605 (N_45605,N_45364,N_45421);
and U45606 (N_45606,N_45371,N_45265);
nor U45607 (N_45607,N_45312,N_45292);
xor U45608 (N_45608,N_45294,N_45480);
nor U45609 (N_45609,N_45286,N_45328);
or U45610 (N_45610,N_45314,N_45495);
and U45611 (N_45611,N_45299,N_45439);
nand U45612 (N_45612,N_45266,N_45310);
nand U45613 (N_45613,N_45464,N_45430);
or U45614 (N_45614,N_45456,N_45390);
xnor U45615 (N_45615,N_45376,N_45405);
or U45616 (N_45616,N_45479,N_45253);
or U45617 (N_45617,N_45306,N_45359);
nand U45618 (N_45618,N_45272,N_45250);
xnor U45619 (N_45619,N_45375,N_45471);
xor U45620 (N_45620,N_45485,N_45317);
xnor U45621 (N_45621,N_45442,N_45322);
and U45622 (N_45622,N_45419,N_45309);
nand U45623 (N_45623,N_45441,N_45386);
or U45624 (N_45624,N_45335,N_45301);
or U45625 (N_45625,N_45267,N_45292);
and U45626 (N_45626,N_45485,N_45283);
xor U45627 (N_45627,N_45463,N_45378);
nor U45628 (N_45628,N_45271,N_45257);
nor U45629 (N_45629,N_45333,N_45438);
and U45630 (N_45630,N_45472,N_45486);
nand U45631 (N_45631,N_45408,N_45396);
or U45632 (N_45632,N_45431,N_45281);
and U45633 (N_45633,N_45447,N_45464);
or U45634 (N_45634,N_45284,N_45325);
and U45635 (N_45635,N_45497,N_45371);
xnor U45636 (N_45636,N_45475,N_45445);
nand U45637 (N_45637,N_45320,N_45260);
or U45638 (N_45638,N_45467,N_45300);
and U45639 (N_45639,N_45346,N_45492);
xnor U45640 (N_45640,N_45363,N_45283);
xor U45641 (N_45641,N_45302,N_45468);
or U45642 (N_45642,N_45339,N_45256);
xor U45643 (N_45643,N_45412,N_45392);
or U45644 (N_45644,N_45382,N_45345);
nand U45645 (N_45645,N_45368,N_45339);
nand U45646 (N_45646,N_45293,N_45451);
and U45647 (N_45647,N_45268,N_45306);
nor U45648 (N_45648,N_45424,N_45420);
xnor U45649 (N_45649,N_45284,N_45344);
and U45650 (N_45650,N_45365,N_45452);
nand U45651 (N_45651,N_45415,N_45486);
nor U45652 (N_45652,N_45397,N_45448);
nand U45653 (N_45653,N_45283,N_45372);
or U45654 (N_45654,N_45499,N_45351);
nor U45655 (N_45655,N_45341,N_45409);
and U45656 (N_45656,N_45395,N_45312);
and U45657 (N_45657,N_45263,N_45368);
nand U45658 (N_45658,N_45364,N_45444);
nand U45659 (N_45659,N_45444,N_45399);
xor U45660 (N_45660,N_45279,N_45418);
or U45661 (N_45661,N_45310,N_45436);
xnor U45662 (N_45662,N_45448,N_45471);
nand U45663 (N_45663,N_45323,N_45489);
nor U45664 (N_45664,N_45343,N_45495);
and U45665 (N_45665,N_45477,N_45272);
nor U45666 (N_45666,N_45393,N_45491);
nand U45667 (N_45667,N_45432,N_45329);
and U45668 (N_45668,N_45326,N_45433);
nand U45669 (N_45669,N_45333,N_45403);
nand U45670 (N_45670,N_45465,N_45354);
nand U45671 (N_45671,N_45267,N_45376);
nand U45672 (N_45672,N_45435,N_45342);
xor U45673 (N_45673,N_45493,N_45361);
nand U45674 (N_45674,N_45394,N_45461);
and U45675 (N_45675,N_45420,N_45487);
or U45676 (N_45676,N_45466,N_45323);
xor U45677 (N_45677,N_45309,N_45391);
nand U45678 (N_45678,N_45455,N_45396);
nor U45679 (N_45679,N_45309,N_45422);
and U45680 (N_45680,N_45398,N_45387);
and U45681 (N_45681,N_45251,N_45329);
and U45682 (N_45682,N_45413,N_45328);
xor U45683 (N_45683,N_45342,N_45452);
and U45684 (N_45684,N_45493,N_45403);
xnor U45685 (N_45685,N_45352,N_45285);
nor U45686 (N_45686,N_45295,N_45445);
xnor U45687 (N_45687,N_45432,N_45465);
xor U45688 (N_45688,N_45427,N_45334);
and U45689 (N_45689,N_45453,N_45263);
or U45690 (N_45690,N_45319,N_45300);
xnor U45691 (N_45691,N_45298,N_45472);
and U45692 (N_45692,N_45313,N_45266);
nand U45693 (N_45693,N_45277,N_45494);
nor U45694 (N_45694,N_45464,N_45325);
or U45695 (N_45695,N_45382,N_45323);
xnor U45696 (N_45696,N_45327,N_45419);
nand U45697 (N_45697,N_45288,N_45465);
and U45698 (N_45698,N_45388,N_45408);
nand U45699 (N_45699,N_45282,N_45263);
or U45700 (N_45700,N_45293,N_45253);
nor U45701 (N_45701,N_45489,N_45475);
nor U45702 (N_45702,N_45285,N_45278);
and U45703 (N_45703,N_45377,N_45371);
nand U45704 (N_45704,N_45330,N_45365);
or U45705 (N_45705,N_45455,N_45482);
nand U45706 (N_45706,N_45480,N_45267);
nor U45707 (N_45707,N_45421,N_45307);
and U45708 (N_45708,N_45416,N_45407);
nor U45709 (N_45709,N_45468,N_45309);
and U45710 (N_45710,N_45419,N_45279);
nor U45711 (N_45711,N_45462,N_45387);
and U45712 (N_45712,N_45289,N_45406);
nor U45713 (N_45713,N_45408,N_45447);
nor U45714 (N_45714,N_45354,N_45253);
nand U45715 (N_45715,N_45393,N_45313);
and U45716 (N_45716,N_45357,N_45404);
nor U45717 (N_45717,N_45357,N_45308);
xnor U45718 (N_45718,N_45435,N_45421);
nor U45719 (N_45719,N_45403,N_45328);
nor U45720 (N_45720,N_45342,N_45289);
or U45721 (N_45721,N_45294,N_45418);
nand U45722 (N_45722,N_45323,N_45435);
xnor U45723 (N_45723,N_45468,N_45449);
and U45724 (N_45724,N_45275,N_45316);
or U45725 (N_45725,N_45456,N_45347);
xor U45726 (N_45726,N_45328,N_45468);
nand U45727 (N_45727,N_45497,N_45486);
and U45728 (N_45728,N_45442,N_45479);
nand U45729 (N_45729,N_45428,N_45469);
xnor U45730 (N_45730,N_45328,N_45333);
nor U45731 (N_45731,N_45487,N_45294);
nor U45732 (N_45732,N_45299,N_45397);
nor U45733 (N_45733,N_45293,N_45415);
xor U45734 (N_45734,N_45427,N_45257);
nor U45735 (N_45735,N_45438,N_45422);
nor U45736 (N_45736,N_45433,N_45377);
or U45737 (N_45737,N_45385,N_45454);
and U45738 (N_45738,N_45344,N_45462);
nor U45739 (N_45739,N_45290,N_45298);
and U45740 (N_45740,N_45441,N_45476);
nand U45741 (N_45741,N_45259,N_45378);
nor U45742 (N_45742,N_45429,N_45467);
or U45743 (N_45743,N_45408,N_45283);
xnor U45744 (N_45744,N_45386,N_45336);
nand U45745 (N_45745,N_45491,N_45439);
xor U45746 (N_45746,N_45311,N_45408);
nand U45747 (N_45747,N_45341,N_45433);
and U45748 (N_45748,N_45429,N_45320);
nor U45749 (N_45749,N_45411,N_45278);
and U45750 (N_45750,N_45579,N_45616);
nand U45751 (N_45751,N_45571,N_45522);
or U45752 (N_45752,N_45576,N_45739);
xnor U45753 (N_45753,N_45558,N_45705);
xnor U45754 (N_45754,N_45557,N_45749);
and U45755 (N_45755,N_45517,N_45574);
nand U45756 (N_45756,N_45707,N_45635);
nand U45757 (N_45757,N_45505,N_45511);
and U45758 (N_45758,N_45527,N_45691);
and U45759 (N_45759,N_45649,N_45748);
nor U45760 (N_45760,N_45550,N_45622);
xnor U45761 (N_45761,N_45524,N_45608);
or U45762 (N_45762,N_45658,N_45681);
or U45763 (N_45763,N_45640,N_45662);
nand U45764 (N_45764,N_45518,N_45516);
nor U45765 (N_45765,N_45699,N_45580);
or U45766 (N_45766,N_45500,N_45602);
and U45767 (N_45767,N_45686,N_45521);
nor U45768 (N_45768,N_45718,N_45530);
xnor U45769 (N_45769,N_45634,N_45697);
or U45770 (N_45770,N_45528,N_45721);
nand U45771 (N_45771,N_45565,N_45730);
or U45772 (N_45772,N_45514,N_45740);
and U45773 (N_45773,N_45611,N_45531);
or U45774 (N_45774,N_45694,N_45667);
or U45775 (N_45775,N_45601,N_45570);
nand U45776 (N_45776,N_45727,N_45656);
xor U45777 (N_45777,N_45737,N_45666);
nor U45778 (N_45778,N_45659,N_45591);
nor U45779 (N_45779,N_45606,N_45588);
xnor U45780 (N_45780,N_45501,N_45726);
xor U45781 (N_45781,N_45729,N_45600);
xor U45782 (N_45782,N_45716,N_45504);
nand U45783 (N_45783,N_45675,N_45563);
nand U45784 (N_45784,N_45626,N_45668);
and U45785 (N_45785,N_45643,N_45743);
xnor U45786 (N_45786,N_45566,N_45738);
nand U45787 (N_45787,N_45541,N_45586);
or U45788 (N_45788,N_45556,N_45693);
and U45789 (N_45789,N_45513,N_45545);
and U45790 (N_45790,N_45597,N_45650);
nand U45791 (N_45791,N_45746,N_45619);
nor U45792 (N_45792,N_45663,N_45560);
xor U45793 (N_45793,N_45725,N_45630);
xnor U45794 (N_45794,N_45529,N_45515);
nor U45795 (N_45795,N_45655,N_45645);
and U45796 (N_45796,N_45661,N_45657);
nor U45797 (N_45797,N_45672,N_45583);
nor U45798 (N_45798,N_45701,N_45651);
nand U45799 (N_45799,N_45589,N_45625);
and U45800 (N_45800,N_45555,N_45603);
nor U45801 (N_45801,N_45723,N_45562);
nor U45802 (N_45802,N_45720,N_45722);
nor U45803 (N_45803,N_45536,N_45612);
nand U45804 (N_45804,N_45508,N_45506);
or U45805 (N_45805,N_45741,N_45654);
xor U45806 (N_45806,N_45677,N_45641);
xor U45807 (N_45807,N_45599,N_45680);
nor U45808 (N_45808,N_45559,N_45647);
nand U45809 (N_45809,N_45569,N_45624);
and U45810 (N_45810,N_45582,N_45593);
nor U45811 (N_45811,N_45639,N_45585);
and U45812 (N_45812,N_45548,N_45510);
nand U45813 (N_45813,N_45735,N_45715);
nand U45814 (N_45814,N_45708,N_45638);
and U45815 (N_45815,N_45590,N_45682);
nor U45816 (N_45816,N_45728,N_45532);
xor U45817 (N_45817,N_45538,N_45724);
nand U45818 (N_45818,N_45642,N_45710);
or U45819 (N_45819,N_45575,N_45533);
nand U45820 (N_45820,N_45687,N_45535);
nor U45821 (N_45821,N_45678,N_45676);
nand U45822 (N_45822,N_45564,N_45523);
nor U45823 (N_45823,N_45671,N_45660);
nand U45824 (N_45824,N_45632,N_45711);
or U45825 (N_45825,N_45549,N_45706);
and U45826 (N_45826,N_45685,N_45547);
and U45827 (N_45827,N_45598,N_45542);
nor U45828 (N_45828,N_45712,N_45644);
xor U45829 (N_45829,N_45594,N_45747);
nor U45830 (N_45830,N_45731,N_45546);
or U45831 (N_45831,N_45700,N_45652);
and U45832 (N_45832,N_45552,N_45665);
xor U45833 (N_45833,N_45502,N_45698);
nor U45834 (N_45834,N_45573,N_45709);
or U45835 (N_45835,N_45539,N_45604);
xnor U45836 (N_45836,N_45745,N_45587);
and U45837 (N_45837,N_45683,N_45736);
nor U45838 (N_45838,N_45537,N_45633);
or U45839 (N_45839,N_45631,N_45702);
nand U45840 (N_45840,N_45595,N_45526);
xor U45841 (N_45841,N_45503,N_45567);
and U45842 (N_45842,N_45534,N_45653);
nand U45843 (N_45843,N_45719,N_45629);
nor U45844 (N_45844,N_45674,N_45636);
or U45845 (N_45845,N_45605,N_45554);
nor U45846 (N_45846,N_45615,N_45696);
nand U45847 (N_45847,N_45561,N_45607);
xnor U45848 (N_45848,N_45520,N_45540);
and U45849 (N_45849,N_45692,N_45610);
or U45850 (N_45850,N_45509,N_45614);
nand U45851 (N_45851,N_45673,N_45617);
nand U45852 (N_45852,N_45581,N_45512);
nor U45853 (N_45853,N_45703,N_45670);
xor U45854 (N_45854,N_45507,N_45568);
nand U45855 (N_45855,N_45713,N_45689);
or U45856 (N_45856,N_45577,N_45592);
or U45857 (N_45857,N_45733,N_45646);
or U45858 (N_45858,N_45551,N_45695);
nand U45859 (N_45859,N_45742,N_45543);
xnor U45860 (N_45860,N_45669,N_45623);
and U45861 (N_45861,N_45596,N_45584);
and U45862 (N_45862,N_45704,N_45621);
and U45863 (N_45863,N_45525,N_45578);
xnor U45864 (N_45864,N_45717,N_45744);
and U45865 (N_45865,N_45714,N_45519);
and U45866 (N_45866,N_45684,N_45620);
or U45867 (N_45867,N_45553,N_45609);
or U45868 (N_45868,N_45648,N_45679);
or U45869 (N_45869,N_45664,N_45618);
nand U45870 (N_45870,N_45628,N_45732);
nand U45871 (N_45871,N_45637,N_45688);
and U45872 (N_45872,N_45627,N_45613);
or U45873 (N_45873,N_45734,N_45690);
or U45874 (N_45874,N_45572,N_45544);
nor U45875 (N_45875,N_45639,N_45709);
xnor U45876 (N_45876,N_45536,N_45595);
or U45877 (N_45877,N_45693,N_45617);
or U45878 (N_45878,N_45738,N_45743);
nor U45879 (N_45879,N_45748,N_45615);
nor U45880 (N_45880,N_45687,N_45705);
and U45881 (N_45881,N_45626,N_45612);
or U45882 (N_45882,N_45737,N_45707);
nand U45883 (N_45883,N_45598,N_45744);
nor U45884 (N_45884,N_45534,N_45742);
nand U45885 (N_45885,N_45594,N_45534);
nand U45886 (N_45886,N_45723,N_45739);
or U45887 (N_45887,N_45561,N_45559);
xnor U45888 (N_45888,N_45663,N_45508);
or U45889 (N_45889,N_45593,N_45635);
or U45890 (N_45890,N_45733,N_45517);
nand U45891 (N_45891,N_45577,N_45557);
nor U45892 (N_45892,N_45550,N_45647);
or U45893 (N_45893,N_45634,N_45604);
nor U45894 (N_45894,N_45559,N_45537);
or U45895 (N_45895,N_45695,N_45686);
and U45896 (N_45896,N_45579,N_45705);
nor U45897 (N_45897,N_45678,N_45582);
xnor U45898 (N_45898,N_45642,N_45628);
nand U45899 (N_45899,N_45582,N_45710);
nor U45900 (N_45900,N_45737,N_45554);
and U45901 (N_45901,N_45602,N_45648);
and U45902 (N_45902,N_45503,N_45653);
or U45903 (N_45903,N_45653,N_45728);
xnor U45904 (N_45904,N_45716,N_45725);
nor U45905 (N_45905,N_45679,N_45731);
or U45906 (N_45906,N_45667,N_45655);
or U45907 (N_45907,N_45562,N_45594);
nand U45908 (N_45908,N_45670,N_45676);
nor U45909 (N_45909,N_45645,N_45726);
xor U45910 (N_45910,N_45542,N_45545);
and U45911 (N_45911,N_45684,N_45654);
xnor U45912 (N_45912,N_45693,N_45506);
or U45913 (N_45913,N_45608,N_45593);
and U45914 (N_45914,N_45566,N_45501);
nand U45915 (N_45915,N_45557,N_45538);
and U45916 (N_45916,N_45588,N_45720);
or U45917 (N_45917,N_45642,N_45532);
or U45918 (N_45918,N_45530,N_45680);
or U45919 (N_45919,N_45638,N_45609);
or U45920 (N_45920,N_45626,N_45560);
or U45921 (N_45921,N_45687,N_45518);
nor U45922 (N_45922,N_45595,N_45560);
nand U45923 (N_45923,N_45520,N_45575);
and U45924 (N_45924,N_45739,N_45603);
or U45925 (N_45925,N_45613,N_45725);
nand U45926 (N_45926,N_45727,N_45660);
and U45927 (N_45927,N_45553,N_45500);
nand U45928 (N_45928,N_45592,N_45571);
and U45929 (N_45929,N_45659,N_45513);
or U45930 (N_45930,N_45616,N_45613);
nor U45931 (N_45931,N_45701,N_45501);
nor U45932 (N_45932,N_45654,N_45713);
or U45933 (N_45933,N_45511,N_45723);
xnor U45934 (N_45934,N_45530,N_45584);
xor U45935 (N_45935,N_45705,N_45673);
or U45936 (N_45936,N_45646,N_45650);
xnor U45937 (N_45937,N_45501,N_45658);
nand U45938 (N_45938,N_45715,N_45675);
nor U45939 (N_45939,N_45683,N_45544);
or U45940 (N_45940,N_45684,N_45543);
xnor U45941 (N_45941,N_45621,N_45571);
nor U45942 (N_45942,N_45558,N_45563);
xnor U45943 (N_45943,N_45716,N_45508);
nor U45944 (N_45944,N_45685,N_45671);
or U45945 (N_45945,N_45748,N_45706);
xor U45946 (N_45946,N_45706,N_45722);
or U45947 (N_45947,N_45716,N_45548);
xnor U45948 (N_45948,N_45540,N_45589);
xor U45949 (N_45949,N_45507,N_45647);
nand U45950 (N_45950,N_45562,N_45610);
or U45951 (N_45951,N_45577,N_45567);
xnor U45952 (N_45952,N_45732,N_45538);
nand U45953 (N_45953,N_45555,N_45630);
or U45954 (N_45954,N_45709,N_45538);
nor U45955 (N_45955,N_45717,N_45515);
or U45956 (N_45956,N_45603,N_45504);
or U45957 (N_45957,N_45539,N_45507);
nand U45958 (N_45958,N_45590,N_45683);
and U45959 (N_45959,N_45520,N_45602);
and U45960 (N_45960,N_45631,N_45735);
and U45961 (N_45961,N_45652,N_45726);
nand U45962 (N_45962,N_45677,N_45536);
nor U45963 (N_45963,N_45652,N_45600);
or U45964 (N_45964,N_45549,N_45614);
or U45965 (N_45965,N_45656,N_45624);
and U45966 (N_45966,N_45742,N_45730);
or U45967 (N_45967,N_45522,N_45687);
or U45968 (N_45968,N_45660,N_45661);
and U45969 (N_45969,N_45744,N_45524);
nor U45970 (N_45970,N_45502,N_45534);
xnor U45971 (N_45971,N_45730,N_45713);
nand U45972 (N_45972,N_45683,N_45720);
or U45973 (N_45973,N_45643,N_45576);
xor U45974 (N_45974,N_45502,N_45712);
or U45975 (N_45975,N_45661,N_45725);
nand U45976 (N_45976,N_45579,N_45731);
and U45977 (N_45977,N_45507,N_45573);
nor U45978 (N_45978,N_45583,N_45639);
and U45979 (N_45979,N_45610,N_45661);
xor U45980 (N_45980,N_45538,N_45588);
and U45981 (N_45981,N_45638,N_45550);
and U45982 (N_45982,N_45649,N_45728);
nor U45983 (N_45983,N_45698,N_45561);
nand U45984 (N_45984,N_45699,N_45641);
and U45985 (N_45985,N_45558,N_45643);
nand U45986 (N_45986,N_45567,N_45559);
xnor U45987 (N_45987,N_45675,N_45508);
or U45988 (N_45988,N_45742,N_45557);
or U45989 (N_45989,N_45586,N_45648);
or U45990 (N_45990,N_45713,N_45537);
nor U45991 (N_45991,N_45537,N_45586);
nand U45992 (N_45992,N_45586,N_45571);
nor U45993 (N_45993,N_45533,N_45749);
nand U45994 (N_45994,N_45607,N_45628);
nor U45995 (N_45995,N_45728,N_45668);
nand U45996 (N_45996,N_45630,N_45655);
nand U45997 (N_45997,N_45576,N_45701);
nand U45998 (N_45998,N_45594,N_45619);
or U45999 (N_45999,N_45638,N_45635);
or U46000 (N_46000,N_45994,N_45865);
xnor U46001 (N_46001,N_45971,N_45788);
nand U46002 (N_46002,N_45955,N_45773);
nor U46003 (N_46003,N_45995,N_45886);
nor U46004 (N_46004,N_45912,N_45963);
and U46005 (N_46005,N_45989,N_45943);
xor U46006 (N_46006,N_45841,N_45812);
or U46007 (N_46007,N_45809,N_45801);
nor U46008 (N_46008,N_45802,N_45873);
nor U46009 (N_46009,N_45923,N_45858);
xnor U46010 (N_46010,N_45902,N_45753);
nor U46011 (N_46011,N_45959,N_45849);
nand U46012 (N_46012,N_45933,N_45766);
or U46013 (N_46013,N_45780,N_45875);
nor U46014 (N_46014,N_45961,N_45761);
nor U46015 (N_46015,N_45915,N_45774);
xnor U46016 (N_46016,N_45920,N_45817);
nand U46017 (N_46017,N_45755,N_45895);
or U46018 (N_46018,N_45868,N_45975);
nor U46019 (N_46019,N_45863,N_45756);
or U46020 (N_46020,N_45917,N_45960);
or U46021 (N_46021,N_45785,N_45847);
xor U46022 (N_46022,N_45832,N_45776);
nor U46023 (N_46023,N_45987,N_45979);
or U46024 (N_46024,N_45767,N_45792);
or U46025 (N_46025,N_45811,N_45821);
and U46026 (N_46026,N_45837,N_45947);
xnor U46027 (N_46027,N_45793,N_45938);
and U46028 (N_46028,N_45814,N_45757);
nand U46029 (N_46029,N_45983,N_45940);
or U46030 (N_46030,N_45911,N_45953);
or U46031 (N_46031,N_45877,N_45931);
or U46032 (N_46032,N_45787,N_45999);
nor U46033 (N_46033,N_45908,N_45997);
nand U46034 (N_46034,N_45867,N_45881);
nand U46035 (N_46035,N_45790,N_45857);
xnor U46036 (N_46036,N_45891,N_45796);
nor U46037 (N_46037,N_45779,N_45883);
and U46038 (N_46038,N_45866,N_45916);
nor U46039 (N_46039,N_45884,N_45958);
xor U46040 (N_46040,N_45752,N_45998);
xnor U46041 (N_46041,N_45860,N_45764);
or U46042 (N_46042,N_45977,N_45988);
and U46043 (N_46043,N_45826,N_45909);
xnor U46044 (N_46044,N_45869,N_45944);
xor U46045 (N_46045,N_45799,N_45816);
nor U46046 (N_46046,N_45850,N_45855);
or U46047 (N_46047,N_45922,N_45833);
xnor U46048 (N_46048,N_45771,N_45907);
and U46049 (N_46049,N_45996,N_45784);
and U46050 (N_46050,N_45934,N_45954);
and U46051 (N_46051,N_45951,N_45921);
and U46052 (N_46052,N_45949,N_45897);
nand U46053 (N_46053,N_45758,N_45791);
nor U46054 (N_46054,N_45765,N_45828);
xor U46055 (N_46055,N_45770,N_45992);
and U46056 (N_46056,N_45763,N_45798);
nor U46057 (N_46057,N_45950,N_45901);
xor U46058 (N_46058,N_45819,N_45781);
nor U46059 (N_46059,N_45818,N_45824);
xnor U46060 (N_46060,N_45903,N_45978);
nand U46061 (N_46061,N_45965,N_45990);
xor U46062 (N_46062,N_45854,N_45823);
nor U46063 (N_46063,N_45794,N_45852);
or U46064 (N_46064,N_45892,N_45810);
nand U46065 (N_46065,N_45926,N_45929);
or U46066 (N_46066,N_45825,N_45806);
nand U46067 (N_46067,N_45967,N_45807);
xor U46068 (N_46068,N_45851,N_45972);
nand U46069 (N_46069,N_45772,N_45845);
and U46070 (N_46070,N_45969,N_45910);
xor U46071 (N_46071,N_45946,N_45751);
and U46072 (N_46072,N_45924,N_45803);
and U46073 (N_46073,N_45984,N_45896);
and U46074 (N_46074,N_45843,N_45830);
xnor U46075 (N_46075,N_45804,N_45941);
nor U46076 (N_46076,N_45846,N_45880);
nor U46077 (N_46077,N_45893,N_45905);
and U46078 (N_46078,N_45900,N_45831);
and U46079 (N_46079,N_45864,N_45839);
nor U46080 (N_46080,N_45870,N_45840);
or U46081 (N_46081,N_45957,N_45861);
nor U46082 (N_46082,N_45822,N_45885);
nor U46083 (N_46083,N_45948,N_45750);
or U46084 (N_46084,N_45836,N_45976);
nand U46085 (N_46085,N_45800,N_45942);
and U46086 (N_46086,N_45859,N_45945);
xnor U46087 (N_46087,N_45842,N_45918);
xnor U46088 (N_46088,N_45887,N_45930);
and U46089 (N_46089,N_45936,N_45789);
xor U46090 (N_46090,N_45835,N_45939);
xnor U46091 (N_46091,N_45913,N_45894);
or U46092 (N_46092,N_45925,N_45985);
nand U46093 (N_46093,N_45874,N_45966);
xor U46094 (N_46094,N_45890,N_45759);
or U46095 (N_46095,N_45876,N_45899);
xnor U46096 (N_46096,N_45919,N_45815);
nor U46097 (N_46097,N_45856,N_45993);
or U46098 (N_46098,N_45782,N_45878);
nor U46099 (N_46099,N_45754,N_45805);
xor U46100 (N_46100,N_45968,N_45879);
or U46101 (N_46101,N_45862,N_45872);
or U46102 (N_46102,N_45838,N_45898);
xor U46103 (N_46103,N_45914,N_45760);
xor U46104 (N_46104,N_45829,N_45795);
and U46105 (N_46105,N_45980,N_45991);
and U46106 (N_46106,N_45848,N_45962);
nor U46107 (N_46107,N_45981,N_45889);
xor U46108 (N_46108,N_45882,N_45834);
nand U46109 (N_46109,N_45775,N_45797);
nand U46110 (N_46110,N_45769,N_45964);
nand U46111 (N_46111,N_45970,N_45853);
nor U46112 (N_46112,N_45986,N_45973);
and U46113 (N_46113,N_45820,N_45786);
nand U46114 (N_46114,N_45906,N_45871);
nand U46115 (N_46115,N_45935,N_45904);
and U46116 (N_46116,N_45956,N_45937);
nor U46117 (N_46117,N_45827,N_45982);
or U46118 (N_46118,N_45813,N_45778);
or U46119 (N_46119,N_45927,N_45932);
or U46120 (N_46120,N_45808,N_45928);
or U46121 (N_46121,N_45952,N_45844);
and U46122 (N_46122,N_45777,N_45768);
and U46123 (N_46123,N_45888,N_45762);
or U46124 (N_46124,N_45783,N_45974);
or U46125 (N_46125,N_45901,N_45995);
and U46126 (N_46126,N_45817,N_45827);
nor U46127 (N_46127,N_45853,N_45886);
xnor U46128 (N_46128,N_45961,N_45783);
or U46129 (N_46129,N_45922,N_45861);
nor U46130 (N_46130,N_45757,N_45835);
and U46131 (N_46131,N_45781,N_45887);
nor U46132 (N_46132,N_45963,N_45948);
and U46133 (N_46133,N_45876,N_45814);
nor U46134 (N_46134,N_45799,N_45982);
or U46135 (N_46135,N_45867,N_45821);
or U46136 (N_46136,N_45752,N_45813);
and U46137 (N_46137,N_45814,N_45857);
or U46138 (N_46138,N_45837,N_45867);
or U46139 (N_46139,N_45904,N_45849);
xnor U46140 (N_46140,N_45911,N_45825);
or U46141 (N_46141,N_45834,N_45778);
xor U46142 (N_46142,N_45989,N_45954);
and U46143 (N_46143,N_45981,N_45847);
or U46144 (N_46144,N_45872,N_45828);
nand U46145 (N_46145,N_45818,N_45987);
and U46146 (N_46146,N_45799,N_45935);
and U46147 (N_46147,N_45954,N_45826);
xnor U46148 (N_46148,N_45781,N_45892);
xor U46149 (N_46149,N_45981,N_45871);
nor U46150 (N_46150,N_45778,N_45974);
nor U46151 (N_46151,N_45765,N_45977);
and U46152 (N_46152,N_45779,N_45785);
nor U46153 (N_46153,N_45806,N_45888);
xnor U46154 (N_46154,N_45791,N_45865);
xor U46155 (N_46155,N_45992,N_45817);
or U46156 (N_46156,N_45858,N_45950);
or U46157 (N_46157,N_45962,N_45878);
xnor U46158 (N_46158,N_45768,N_45979);
or U46159 (N_46159,N_45821,N_45859);
or U46160 (N_46160,N_45805,N_45886);
xor U46161 (N_46161,N_45902,N_45810);
and U46162 (N_46162,N_45923,N_45831);
nand U46163 (N_46163,N_45786,N_45939);
xnor U46164 (N_46164,N_45982,N_45909);
or U46165 (N_46165,N_45782,N_45975);
xor U46166 (N_46166,N_45992,N_45877);
nand U46167 (N_46167,N_45878,N_45755);
nand U46168 (N_46168,N_45822,N_45754);
and U46169 (N_46169,N_45884,N_45954);
and U46170 (N_46170,N_45867,N_45882);
nor U46171 (N_46171,N_45931,N_45924);
xnor U46172 (N_46172,N_45983,N_45878);
or U46173 (N_46173,N_45767,N_45950);
xor U46174 (N_46174,N_45935,N_45810);
and U46175 (N_46175,N_45878,N_45934);
nor U46176 (N_46176,N_45761,N_45883);
and U46177 (N_46177,N_45898,N_45787);
and U46178 (N_46178,N_45879,N_45898);
or U46179 (N_46179,N_45915,N_45813);
xnor U46180 (N_46180,N_45906,N_45917);
or U46181 (N_46181,N_45959,N_45962);
nor U46182 (N_46182,N_45915,N_45841);
and U46183 (N_46183,N_45837,N_45930);
nand U46184 (N_46184,N_45795,N_45888);
and U46185 (N_46185,N_45828,N_45937);
xor U46186 (N_46186,N_45913,N_45886);
nand U46187 (N_46187,N_45846,N_45901);
nor U46188 (N_46188,N_45774,N_45763);
and U46189 (N_46189,N_45857,N_45786);
nand U46190 (N_46190,N_45912,N_45802);
nor U46191 (N_46191,N_45843,N_45793);
and U46192 (N_46192,N_45767,N_45972);
nand U46193 (N_46193,N_45763,N_45955);
nand U46194 (N_46194,N_45830,N_45991);
and U46195 (N_46195,N_45859,N_45800);
and U46196 (N_46196,N_45823,N_45889);
nand U46197 (N_46197,N_45911,N_45834);
nand U46198 (N_46198,N_45815,N_45965);
nor U46199 (N_46199,N_45932,N_45755);
and U46200 (N_46200,N_45933,N_45872);
and U46201 (N_46201,N_45958,N_45933);
nand U46202 (N_46202,N_45763,N_45970);
nand U46203 (N_46203,N_45879,N_45759);
nor U46204 (N_46204,N_45953,N_45969);
nor U46205 (N_46205,N_45982,N_45851);
nor U46206 (N_46206,N_45765,N_45941);
or U46207 (N_46207,N_45903,N_45793);
nand U46208 (N_46208,N_45811,N_45752);
or U46209 (N_46209,N_45820,N_45813);
nand U46210 (N_46210,N_45964,N_45823);
nand U46211 (N_46211,N_45900,N_45753);
xor U46212 (N_46212,N_45868,N_45920);
xor U46213 (N_46213,N_45923,N_45915);
nand U46214 (N_46214,N_45960,N_45997);
and U46215 (N_46215,N_45913,N_45924);
nand U46216 (N_46216,N_45922,N_45920);
nor U46217 (N_46217,N_45894,N_45759);
and U46218 (N_46218,N_45961,N_45863);
or U46219 (N_46219,N_45897,N_45858);
or U46220 (N_46220,N_45775,N_45960);
and U46221 (N_46221,N_45913,N_45906);
and U46222 (N_46222,N_45893,N_45898);
or U46223 (N_46223,N_45963,N_45900);
xnor U46224 (N_46224,N_45962,N_45979);
xor U46225 (N_46225,N_45994,N_45793);
and U46226 (N_46226,N_45922,N_45923);
or U46227 (N_46227,N_45993,N_45762);
or U46228 (N_46228,N_45802,N_45895);
nor U46229 (N_46229,N_45948,N_45901);
nor U46230 (N_46230,N_45764,N_45894);
xor U46231 (N_46231,N_45989,N_45894);
and U46232 (N_46232,N_45874,N_45896);
nor U46233 (N_46233,N_45963,N_45981);
or U46234 (N_46234,N_45908,N_45771);
or U46235 (N_46235,N_45923,N_45961);
nand U46236 (N_46236,N_45868,N_45763);
or U46237 (N_46237,N_45767,N_45817);
or U46238 (N_46238,N_45765,N_45884);
xor U46239 (N_46239,N_45794,N_45972);
or U46240 (N_46240,N_45808,N_45781);
and U46241 (N_46241,N_45839,N_45959);
or U46242 (N_46242,N_45870,N_45765);
and U46243 (N_46243,N_45931,N_45857);
nand U46244 (N_46244,N_45810,N_45989);
and U46245 (N_46245,N_45759,N_45932);
nor U46246 (N_46246,N_45877,N_45986);
nor U46247 (N_46247,N_45752,N_45959);
nor U46248 (N_46248,N_45920,N_45993);
nand U46249 (N_46249,N_45851,N_45984);
or U46250 (N_46250,N_46072,N_46107);
or U46251 (N_46251,N_46192,N_46211);
and U46252 (N_46252,N_46184,N_46030);
nor U46253 (N_46253,N_46081,N_46171);
and U46254 (N_46254,N_46153,N_46177);
or U46255 (N_46255,N_46045,N_46005);
xor U46256 (N_46256,N_46068,N_46145);
xnor U46257 (N_46257,N_46006,N_46013);
or U46258 (N_46258,N_46056,N_46008);
or U46259 (N_46259,N_46239,N_46098);
nor U46260 (N_46260,N_46168,N_46039);
xnor U46261 (N_46261,N_46240,N_46135);
nor U46262 (N_46262,N_46009,N_46046);
and U46263 (N_46263,N_46034,N_46036);
nand U46264 (N_46264,N_46178,N_46246);
and U46265 (N_46265,N_46043,N_46132);
nand U46266 (N_46266,N_46076,N_46058);
nand U46267 (N_46267,N_46194,N_46041);
nand U46268 (N_46268,N_46065,N_46084);
and U46269 (N_46269,N_46229,N_46183);
and U46270 (N_46270,N_46237,N_46222);
and U46271 (N_46271,N_46015,N_46071);
nand U46272 (N_46272,N_46025,N_46121);
and U46273 (N_46273,N_46028,N_46219);
nor U46274 (N_46274,N_46108,N_46161);
or U46275 (N_46275,N_46055,N_46129);
and U46276 (N_46276,N_46086,N_46131);
xor U46277 (N_46277,N_46149,N_46180);
and U46278 (N_46278,N_46124,N_46191);
or U46279 (N_46279,N_46249,N_46226);
nand U46280 (N_46280,N_46190,N_46163);
nand U46281 (N_46281,N_46220,N_46140);
xor U46282 (N_46282,N_46127,N_46155);
xnor U46283 (N_46283,N_46148,N_46067);
or U46284 (N_46284,N_46066,N_46095);
or U46285 (N_46285,N_46119,N_46196);
or U46286 (N_46286,N_46130,N_46169);
and U46287 (N_46287,N_46186,N_46099);
nand U46288 (N_46288,N_46032,N_46059);
nor U46289 (N_46289,N_46234,N_46014);
or U46290 (N_46290,N_46231,N_46233);
xor U46291 (N_46291,N_46115,N_46199);
nor U46292 (N_46292,N_46112,N_46089);
nand U46293 (N_46293,N_46210,N_46012);
or U46294 (N_46294,N_46111,N_46128);
xor U46295 (N_46295,N_46026,N_46151);
nand U46296 (N_46296,N_46187,N_46003);
or U46297 (N_46297,N_46212,N_46174);
xnor U46298 (N_46298,N_46203,N_46200);
xor U46299 (N_46299,N_46204,N_46104);
xnor U46300 (N_46300,N_46173,N_46117);
or U46301 (N_46301,N_46054,N_46159);
nand U46302 (N_46302,N_46092,N_46214);
nand U46303 (N_46303,N_46218,N_46053);
nand U46304 (N_46304,N_46074,N_46040);
or U46305 (N_46305,N_46018,N_46181);
and U46306 (N_46306,N_46142,N_46031);
or U46307 (N_46307,N_46134,N_46179);
and U46308 (N_46308,N_46205,N_46238);
and U46309 (N_46309,N_46110,N_46088);
or U46310 (N_46310,N_46101,N_46096);
nand U46311 (N_46311,N_46091,N_46216);
or U46312 (N_46312,N_46133,N_46202);
or U46313 (N_46313,N_46138,N_46002);
xnor U46314 (N_46314,N_46152,N_46077);
and U46315 (N_46315,N_46080,N_46073);
nand U46316 (N_46316,N_46158,N_46165);
nor U46317 (N_46317,N_46209,N_46000);
nor U46318 (N_46318,N_46069,N_46215);
or U46319 (N_46319,N_46198,N_46182);
and U46320 (N_46320,N_46090,N_46075);
nand U46321 (N_46321,N_46156,N_46241);
nand U46322 (N_46322,N_46038,N_46166);
and U46323 (N_46323,N_46035,N_46011);
nand U46324 (N_46324,N_46019,N_46118);
nand U46325 (N_46325,N_46123,N_46172);
and U46326 (N_46326,N_46193,N_46082);
or U46327 (N_46327,N_46247,N_46060);
or U46328 (N_46328,N_46024,N_46010);
xnor U46329 (N_46329,N_46244,N_46230);
and U46330 (N_46330,N_46044,N_46120);
nor U46331 (N_46331,N_46245,N_46016);
or U46332 (N_46332,N_46062,N_46021);
xor U46333 (N_46333,N_46146,N_46052);
xnor U46334 (N_46334,N_46147,N_46162);
nand U46335 (N_46335,N_46243,N_46160);
nor U46336 (N_46336,N_46049,N_46139);
or U46337 (N_46337,N_46126,N_46175);
and U46338 (N_46338,N_46157,N_46232);
xor U46339 (N_46339,N_46235,N_46078);
and U46340 (N_46340,N_46087,N_46213);
or U46341 (N_46341,N_46197,N_46027);
or U46342 (N_46342,N_46201,N_46102);
and U46343 (N_46343,N_46094,N_46063);
xor U46344 (N_46344,N_46051,N_46105);
and U46345 (N_46345,N_46001,N_46122);
nand U46346 (N_46346,N_46224,N_46217);
or U46347 (N_46347,N_46236,N_46114);
nor U46348 (N_46348,N_46042,N_46164);
or U46349 (N_46349,N_46004,N_46103);
and U46350 (N_46350,N_46109,N_46136);
xnor U46351 (N_46351,N_46225,N_46223);
xnor U46352 (N_46352,N_46170,N_46227);
or U46353 (N_46353,N_46029,N_46017);
or U46354 (N_46354,N_46167,N_46022);
and U46355 (N_46355,N_46048,N_46064);
nor U46356 (N_46356,N_46047,N_46050);
or U46357 (N_46357,N_46113,N_46020);
and U46358 (N_46358,N_46125,N_46141);
nand U46359 (N_46359,N_46207,N_46023);
nand U46360 (N_46360,N_46248,N_46185);
and U46361 (N_46361,N_46144,N_46189);
or U46362 (N_46362,N_46221,N_46093);
or U46363 (N_46363,N_46100,N_46057);
and U46364 (N_46364,N_46037,N_46143);
or U46365 (N_46365,N_46083,N_46206);
xnor U46366 (N_46366,N_46228,N_46242);
nor U46367 (N_46367,N_46106,N_46176);
xnor U46368 (N_46368,N_46061,N_46150);
xor U46369 (N_46369,N_46079,N_46188);
xnor U46370 (N_46370,N_46097,N_46070);
nand U46371 (N_46371,N_46116,N_46007);
nor U46372 (N_46372,N_46033,N_46137);
or U46373 (N_46373,N_46195,N_46154);
xor U46374 (N_46374,N_46085,N_46208);
nand U46375 (N_46375,N_46059,N_46114);
xor U46376 (N_46376,N_46204,N_46112);
nand U46377 (N_46377,N_46244,N_46082);
or U46378 (N_46378,N_46223,N_46085);
xnor U46379 (N_46379,N_46068,N_46060);
and U46380 (N_46380,N_46221,N_46157);
and U46381 (N_46381,N_46057,N_46108);
xnor U46382 (N_46382,N_46120,N_46236);
xor U46383 (N_46383,N_46051,N_46113);
or U46384 (N_46384,N_46201,N_46055);
nand U46385 (N_46385,N_46148,N_46075);
and U46386 (N_46386,N_46119,N_46222);
or U46387 (N_46387,N_46053,N_46224);
nor U46388 (N_46388,N_46234,N_46044);
and U46389 (N_46389,N_46103,N_46210);
or U46390 (N_46390,N_46149,N_46092);
nand U46391 (N_46391,N_46109,N_46048);
or U46392 (N_46392,N_46192,N_46028);
and U46393 (N_46393,N_46073,N_46156);
and U46394 (N_46394,N_46129,N_46223);
or U46395 (N_46395,N_46235,N_46184);
and U46396 (N_46396,N_46123,N_46217);
nor U46397 (N_46397,N_46215,N_46093);
nand U46398 (N_46398,N_46136,N_46145);
nor U46399 (N_46399,N_46040,N_46065);
xnor U46400 (N_46400,N_46207,N_46160);
xnor U46401 (N_46401,N_46024,N_46233);
and U46402 (N_46402,N_46213,N_46127);
or U46403 (N_46403,N_46230,N_46075);
and U46404 (N_46404,N_46152,N_46158);
nor U46405 (N_46405,N_46039,N_46104);
nor U46406 (N_46406,N_46247,N_46141);
and U46407 (N_46407,N_46044,N_46206);
nand U46408 (N_46408,N_46150,N_46112);
or U46409 (N_46409,N_46131,N_46184);
nand U46410 (N_46410,N_46009,N_46020);
xor U46411 (N_46411,N_46190,N_46202);
or U46412 (N_46412,N_46168,N_46100);
xnor U46413 (N_46413,N_46065,N_46165);
or U46414 (N_46414,N_46164,N_46044);
nor U46415 (N_46415,N_46144,N_46058);
or U46416 (N_46416,N_46231,N_46234);
or U46417 (N_46417,N_46219,N_46137);
or U46418 (N_46418,N_46059,N_46058);
and U46419 (N_46419,N_46199,N_46145);
xnor U46420 (N_46420,N_46129,N_46202);
xnor U46421 (N_46421,N_46097,N_46176);
nor U46422 (N_46422,N_46231,N_46056);
xnor U46423 (N_46423,N_46015,N_46112);
or U46424 (N_46424,N_46090,N_46231);
xnor U46425 (N_46425,N_46188,N_46182);
or U46426 (N_46426,N_46192,N_46152);
nand U46427 (N_46427,N_46067,N_46160);
and U46428 (N_46428,N_46170,N_46018);
nand U46429 (N_46429,N_46243,N_46085);
nor U46430 (N_46430,N_46149,N_46222);
and U46431 (N_46431,N_46078,N_46146);
nor U46432 (N_46432,N_46038,N_46075);
xnor U46433 (N_46433,N_46161,N_46157);
nand U46434 (N_46434,N_46165,N_46116);
nor U46435 (N_46435,N_46089,N_46029);
and U46436 (N_46436,N_46155,N_46247);
or U46437 (N_46437,N_46141,N_46187);
nand U46438 (N_46438,N_46118,N_46166);
or U46439 (N_46439,N_46085,N_46148);
xor U46440 (N_46440,N_46111,N_46198);
xor U46441 (N_46441,N_46025,N_46081);
xnor U46442 (N_46442,N_46016,N_46147);
and U46443 (N_46443,N_46023,N_46102);
nor U46444 (N_46444,N_46130,N_46154);
nand U46445 (N_46445,N_46046,N_46049);
nor U46446 (N_46446,N_46221,N_46012);
xor U46447 (N_46447,N_46118,N_46039);
xor U46448 (N_46448,N_46038,N_46187);
nor U46449 (N_46449,N_46060,N_46127);
and U46450 (N_46450,N_46142,N_46074);
or U46451 (N_46451,N_46176,N_46191);
and U46452 (N_46452,N_46081,N_46037);
or U46453 (N_46453,N_46244,N_46059);
or U46454 (N_46454,N_46127,N_46180);
or U46455 (N_46455,N_46003,N_46112);
and U46456 (N_46456,N_46032,N_46100);
or U46457 (N_46457,N_46239,N_46136);
nand U46458 (N_46458,N_46058,N_46245);
xor U46459 (N_46459,N_46206,N_46192);
nor U46460 (N_46460,N_46209,N_46194);
xor U46461 (N_46461,N_46236,N_46041);
nor U46462 (N_46462,N_46087,N_46204);
and U46463 (N_46463,N_46226,N_46187);
or U46464 (N_46464,N_46185,N_46159);
and U46465 (N_46465,N_46017,N_46222);
or U46466 (N_46466,N_46148,N_46147);
nor U46467 (N_46467,N_46147,N_46040);
nand U46468 (N_46468,N_46153,N_46038);
or U46469 (N_46469,N_46084,N_46015);
nand U46470 (N_46470,N_46143,N_46133);
or U46471 (N_46471,N_46024,N_46180);
or U46472 (N_46472,N_46148,N_46058);
or U46473 (N_46473,N_46084,N_46049);
and U46474 (N_46474,N_46124,N_46152);
and U46475 (N_46475,N_46071,N_46105);
or U46476 (N_46476,N_46075,N_46165);
xor U46477 (N_46477,N_46179,N_46193);
nand U46478 (N_46478,N_46248,N_46058);
nor U46479 (N_46479,N_46032,N_46114);
and U46480 (N_46480,N_46169,N_46196);
nand U46481 (N_46481,N_46099,N_46112);
or U46482 (N_46482,N_46061,N_46106);
nor U46483 (N_46483,N_46128,N_46190);
and U46484 (N_46484,N_46025,N_46128);
and U46485 (N_46485,N_46063,N_46045);
or U46486 (N_46486,N_46243,N_46128);
nand U46487 (N_46487,N_46185,N_46075);
nand U46488 (N_46488,N_46069,N_46017);
or U46489 (N_46489,N_46208,N_46126);
nand U46490 (N_46490,N_46102,N_46183);
nor U46491 (N_46491,N_46065,N_46100);
and U46492 (N_46492,N_46089,N_46030);
or U46493 (N_46493,N_46239,N_46221);
or U46494 (N_46494,N_46197,N_46144);
and U46495 (N_46495,N_46180,N_46085);
nand U46496 (N_46496,N_46030,N_46205);
nor U46497 (N_46497,N_46202,N_46128);
nor U46498 (N_46498,N_46003,N_46080);
and U46499 (N_46499,N_46219,N_46187);
or U46500 (N_46500,N_46470,N_46261);
or U46501 (N_46501,N_46413,N_46474);
nand U46502 (N_46502,N_46294,N_46485);
nand U46503 (N_46503,N_46357,N_46283);
nand U46504 (N_46504,N_46303,N_46489);
nand U46505 (N_46505,N_46346,N_46458);
nor U46506 (N_46506,N_46439,N_46441);
and U46507 (N_46507,N_46277,N_46463);
nand U46508 (N_46508,N_46311,N_46358);
nor U46509 (N_46509,N_46384,N_46268);
or U46510 (N_46510,N_46396,N_46348);
xor U46511 (N_46511,N_46481,N_46267);
nor U46512 (N_46512,N_46304,N_46265);
or U46513 (N_46513,N_46334,N_46479);
nand U46514 (N_46514,N_46299,N_46289);
nor U46515 (N_46515,N_46271,N_46350);
or U46516 (N_46516,N_46386,N_46445);
nand U46517 (N_46517,N_46250,N_46467);
nand U46518 (N_46518,N_46272,N_46459);
nand U46519 (N_46519,N_46259,N_46438);
or U46520 (N_46520,N_46476,N_46340);
nand U46521 (N_46521,N_46302,N_46468);
and U46522 (N_46522,N_46310,N_46366);
xor U46523 (N_46523,N_46359,N_46351);
nand U46524 (N_46524,N_46446,N_46473);
and U46525 (N_46525,N_46253,N_46430);
nand U46526 (N_46526,N_46332,N_46280);
nor U46527 (N_46527,N_46330,N_46297);
or U46528 (N_46528,N_46404,N_46497);
nand U46529 (N_46529,N_46451,N_46492);
xnor U46530 (N_46530,N_46282,N_46314);
nand U46531 (N_46531,N_46493,N_46490);
xor U46532 (N_46532,N_46354,N_46369);
and U46533 (N_46533,N_46405,N_46312);
nand U46534 (N_46534,N_46365,N_46275);
and U46535 (N_46535,N_46411,N_46427);
and U46536 (N_46536,N_46382,N_46373);
xnor U46537 (N_46537,N_46429,N_46360);
xnor U46538 (N_46538,N_46424,N_46447);
nor U46539 (N_46539,N_46449,N_46252);
xor U46540 (N_46540,N_46442,N_46440);
and U46541 (N_46541,N_46389,N_46431);
xor U46542 (N_46542,N_46378,N_46420);
nand U46543 (N_46543,N_46270,N_46323);
nor U46544 (N_46544,N_46412,N_46408);
nor U46545 (N_46545,N_46327,N_46251);
nor U46546 (N_46546,N_46324,N_46333);
nor U46547 (N_46547,N_46347,N_46495);
or U46548 (N_46548,N_46484,N_46264);
nand U46549 (N_46549,N_46421,N_46279);
xnor U46550 (N_46550,N_46343,N_46452);
nor U46551 (N_46551,N_46383,N_46276);
nand U46552 (N_46552,N_46262,N_46388);
nand U46553 (N_46553,N_46335,N_46472);
nand U46554 (N_46554,N_46336,N_46345);
and U46555 (N_46555,N_46494,N_46273);
xnor U46556 (N_46556,N_46296,N_46301);
nor U46557 (N_46557,N_46255,N_46319);
or U46558 (N_46558,N_46361,N_46368);
nor U46559 (N_46559,N_46318,N_46260);
nor U46560 (N_46560,N_46326,N_46456);
xor U46561 (N_46561,N_46370,N_46480);
xor U46562 (N_46562,N_46414,N_46305);
nor U46563 (N_46563,N_46422,N_46356);
nand U46564 (N_46564,N_46290,N_46407);
xor U46565 (N_46565,N_46313,N_46392);
and U46566 (N_46566,N_46399,N_46258);
nor U46567 (N_46567,N_46433,N_46434);
or U46568 (N_46568,N_46423,N_46342);
nand U46569 (N_46569,N_46465,N_46328);
nor U46570 (N_46570,N_46418,N_46287);
or U46571 (N_46571,N_46362,N_46380);
xor U46572 (N_46572,N_46466,N_46448);
nand U46573 (N_46573,N_46464,N_46352);
xor U46574 (N_46574,N_46391,N_46406);
nand U46575 (N_46575,N_46403,N_46417);
nand U46576 (N_46576,N_46400,N_46371);
xor U46577 (N_46577,N_46372,N_46455);
or U46578 (N_46578,N_46288,N_46321);
nand U46579 (N_46579,N_46322,N_46339);
nor U46580 (N_46580,N_46409,N_46374);
nand U46581 (N_46581,N_46278,N_46376);
xnor U46582 (N_46582,N_46460,N_46266);
nor U46583 (N_46583,N_46401,N_46394);
xnor U46584 (N_46584,N_46315,N_46381);
xnor U46585 (N_46585,N_46415,N_46496);
nor U46586 (N_46586,N_46344,N_46367);
and U46587 (N_46587,N_46457,N_46390);
and U46588 (N_46588,N_46329,N_46478);
xor U46589 (N_46589,N_46471,N_46461);
or U46590 (N_46590,N_46462,N_46307);
nor U46591 (N_46591,N_46385,N_46402);
nor U46592 (N_46592,N_46488,N_46483);
nor U46593 (N_46593,N_46263,N_46274);
and U46594 (N_46594,N_46395,N_46377);
nor U46595 (N_46595,N_46375,N_46353);
nand U46596 (N_46596,N_46317,N_46341);
and U46597 (N_46597,N_46337,N_46428);
nor U46598 (N_46598,N_46499,N_46285);
and U46599 (N_46599,N_46349,N_46487);
or U46600 (N_46600,N_46482,N_46331);
and U46601 (N_46601,N_46325,N_46425);
or U46602 (N_46602,N_46306,N_46269);
nor U46603 (N_46603,N_46469,N_46300);
nand U46604 (N_46604,N_46397,N_46355);
nor U46605 (N_46605,N_46309,N_46432);
xor U46606 (N_46606,N_46491,N_46410);
or U46607 (N_46607,N_46286,N_46293);
or U46608 (N_46608,N_46292,N_46393);
or U46609 (N_46609,N_46387,N_46257);
xnor U46610 (N_46610,N_46320,N_46475);
nor U46611 (N_46611,N_46443,N_46291);
nor U46612 (N_46612,N_46364,N_46398);
xor U46613 (N_46613,N_46316,N_46363);
and U46614 (N_46614,N_46437,N_46416);
and U46615 (N_46615,N_46284,N_46379);
and U46616 (N_46616,N_46254,N_46454);
nor U46617 (N_46617,N_46338,N_46256);
or U46618 (N_46618,N_46477,N_46298);
nor U46619 (N_46619,N_46436,N_46426);
xnor U46620 (N_46620,N_46486,N_46281);
and U46621 (N_46621,N_46444,N_46450);
nand U46622 (N_46622,N_46295,N_46308);
nand U46623 (N_46623,N_46453,N_46498);
nor U46624 (N_46624,N_46435,N_46419);
xnor U46625 (N_46625,N_46439,N_46437);
or U46626 (N_46626,N_46309,N_46433);
nand U46627 (N_46627,N_46317,N_46475);
nor U46628 (N_46628,N_46410,N_46300);
or U46629 (N_46629,N_46300,N_46403);
xor U46630 (N_46630,N_46338,N_46399);
nand U46631 (N_46631,N_46446,N_46351);
nor U46632 (N_46632,N_46490,N_46485);
nor U46633 (N_46633,N_46265,N_46383);
or U46634 (N_46634,N_46340,N_46296);
or U46635 (N_46635,N_46345,N_46312);
xnor U46636 (N_46636,N_46262,N_46306);
xnor U46637 (N_46637,N_46474,N_46301);
or U46638 (N_46638,N_46467,N_46266);
or U46639 (N_46639,N_46387,N_46287);
nor U46640 (N_46640,N_46456,N_46497);
and U46641 (N_46641,N_46451,N_46360);
nand U46642 (N_46642,N_46341,N_46254);
or U46643 (N_46643,N_46393,N_46468);
or U46644 (N_46644,N_46366,N_46380);
xnor U46645 (N_46645,N_46406,N_46314);
xor U46646 (N_46646,N_46337,N_46482);
and U46647 (N_46647,N_46405,N_46291);
and U46648 (N_46648,N_46461,N_46275);
and U46649 (N_46649,N_46341,N_46297);
or U46650 (N_46650,N_46309,N_46266);
nand U46651 (N_46651,N_46256,N_46411);
nor U46652 (N_46652,N_46358,N_46250);
nor U46653 (N_46653,N_46257,N_46468);
and U46654 (N_46654,N_46369,N_46375);
xnor U46655 (N_46655,N_46489,N_46436);
nand U46656 (N_46656,N_46300,N_46396);
nor U46657 (N_46657,N_46432,N_46358);
nor U46658 (N_46658,N_46308,N_46430);
xor U46659 (N_46659,N_46259,N_46443);
and U46660 (N_46660,N_46354,N_46256);
nand U46661 (N_46661,N_46464,N_46330);
or U46662 (N_46662,N_46452,N_46471);
nor U46663 (N_46663,N_46292,N_46336);
and U46664 (N_46664,N_46311,N_46469);
nand U46665 (N_46665,N_46439,N_46352);
nand U46666 (N_46666,N_46455,N_46499);
xnor U46667 (N_46667,N_46256,N_46454);
nand U46668 (N_46668,N_46349,N_46376);
nand U46669 (N_46669,N_46284,N_46319);
nand U46670 (N_46670,N_46360,N_46310);
or U46671 (N_46671,N_46366,N_46356);
or U46672 (N_46672,N_46364,N_46313);
or U46673 (N_46673,N_46444,N_46377);
or U46674 (N_46674,N_46462,N_46393);
nor U46675 (N_46675,N_46387,N_46379);
or U46676 (N_46676,N_46302,N_46339);
or U46677 (N_46677,N_46368,N_46335);
or U46678 (N_46678,N_46355,N_46281);
and U46679 (N_46679,N_46332,N_46327);
xnor U46680 (N_46680,N_46294,N_46342);
nor U46681 (N_46681,N_46482,N_46328);
and U46682 (N_46682,N_46399,N_46392);
nor U46683 (N_46683,N_46411,N_46301);
and U46684 (N_46684,N_46267,N_46399);
or U46685 (N_46685,N_46393,N_46453);
nand U46686 (N_46686,N_46364,N_46459);
and U46687 (N_46687,N_46452,N_46329);
and U46688 (N_46688,N_46422,N_46478);
xnor U46689 (N_46689,N_46253,N_46265);
or U46690 (N_46690,N_46447,N_46271);
nand U46691 (N_46691,N_46426,N_46498);
nor U46692 (N_46692,N_46252,N_46304);
xor U46693 (N_46693,N_46329,N_46356);
and U46694 (N_46694,N_46285,N_46486);
or U46695 (N_46695,N_46283,N_46278);
xnor U46696 (N_46696,N_46477,N_46265);
xor U46697 (N_46697,N_46260,N_46359);
and U46698 (N_46698,N_46269,N_46320);
or U46699 (N_46699,N_46465,N_46347);
xor U46700 (N_46700,N_46396,N_46473);
nor U46701 (N_46701,N_46307,N_46372);
and U46702 (N_46702,N_46488,N_46441);
or U46703 (N_46703,N_46440,N_46302);
or U46704 (N_46704,N_46414,N_46289);
or U46705 (N_46705,N_46322,N_46308);
xor U46706 (N_46706,N_46354,N_46435);
nand U46707 (N_46707,N_46393,N_46348);
or U46708 (N_46708,N_46386,N_46297);
nor U46709 (N_46709,N_46286,N_46360);
nor U46710 (N_46710,N_46372,N_46438);
nor U46711 (N_46711,N_46302,N_46324);
nand U46712 (N_46712,N_46328,N_46488);
or U46713 (N_46713,N_46489,N_46347);
or U46714 (N_46714,N_46253,N_46467);
or U46715 (N_46715,N_46474,N_46314);
nand U46716 (N_46716,N_46316,N_46414);
nand U46717 (N_46717,N_46426,N_46301);
nand U46718 (N_46718,N_46424,N_46463);
xnor U46719 (N_46719,N_46256,N_46439);
nor U46720 (N_46720,N_46281,N_46290);
nand U46721 (N_46721,N_46303,N_46381);
xor U46722 (N_46722,N_46365,N_46409);
xor U46723 (N_46723,N_46449,N_46386);
and U46724 (N_46724,N_46487,N_46459);
xor U46725 (N_46725,N_46268,N_46406);
xor U46726 (N_46726,N_46481,N_46413);
or U46727 (N_46727,N_46397,N_46493);
and U46728 (N_46728,N_46416,N_46320);
xor U46729 (N_46729,N_46411,N_46486);
xor U46730 (N_46730,N_46298,N_46413);
or U46731 (N_46731,N_46352,N_46447);
or U46732 (N_46732,N_46478,N_46310);
nand U46733 (N_46733,N_46405,N_46443);
nand U46734 (N_46734,N_46451,N_46334);
and U46735 (N_46735,N_46258,N_46333);
or U46736 (N_46736,N_46326,N_46373);
or U46737 (N_46737,N_46430,N_46403);
or U46738 (N_46738,N_46263,N_46421);
xor U46739 (N_46739,N_46415,N_46268);
nor U46740 (N_46740,N_46266,N_46444);
nor U46741 (N_46741,N_46340,N_46426);
and U46742 (N_46742,N_46380,N_46441);
and U46743 (N_46743,N_46483,N_46498);
or U46744 (N_46744,N_46327,N_46362);
nand U46745 (N_46745,N_46251,N_46270);
xnor U46746 (N_46746,N_46476,N_46409);
xor U46747 (N_46747,N_46477,N_46428);
nor U46748 (N_46748,N_46366,N_46330);
nand U46749 (N_46749,N_46352,N_46470);
nand U46750 (N_46750,N_46573,N_46562);
or U46751 (N_46751,N_46710,N_46544);
nand U46752 (N_46752,N_46684,N_46654);
nor U46753 (N_46753,N_46570,N_46548);
nand U46754 (N_46754,N_46707,N_46557);
or U46755 (N_46755,N_46723,N_46554);
and U46756 (N_46756,N_46526,N_46641);
nor U46757 (N_46757,N_46728,N_46613);
nand U46758 (N_46758,N_46511,N_46620);
or U46759 (N_46759,N_46740,N_46632);
or U46760 (N_46760,N_46715,N_46651);
nor U46761 (N_46761,N_46605,N_46576);
nand U46762 (N_46762,N_46578,N_46599);
or U46763 (N_46763,N_46595,N_46666);
nand U46764 (N_46764,N_46509,N_46726);
xor U46765 (N_46765,N_46542,N_46628);
nor U46766 (N_46766,N_46579,N_46656);
or U46767 (N_46767,N_46593,N_46518);
nand U46768 (N_46768,N_46541,N_46712);
and U46769 (N_46769,N_46692,N_46618);
nand U46770 (N_46770,N_46742,N_46686);
or U46771 (N_46771,N_46670,N_46673);
nand U46772 (N_46772,N_46659,N_46635);
or U46773 (N_46773,N_46722,N_46743);
nand U46774 (N_46774,N_46683,N_46504);
or U46775 (N_46775,N_46729,N_46727);
or U46776 (N_46776,N_46567,N_46506);
xor U46777 (N_46777,N_46560,N_46581);
or U46778 (N_46778,N_46564,N_46552);
xor U46779 (N_46779,N_46649,N_46633);
nor U46780 (N_46780,N_46720,N_46711);
nand U46781 (N_46781,N_46690,N_46555);
nor U46782 (N_46782,N_46592,N_46547);
nor U46783 (N_46783,N_46736,N_46627);
nor U46784 (N_46784,N_46553,N_46622);
and U46785 (N_46785,N_46596,N_46660);
or U46786 (N_46786,N_46508,N_46536);
or U46787 (N_46787,N_46519,N_46730);
nor U46788 (N_46788,N_46708,N_46677);
xnor U46789 (N_46789,N_46513,N_46588);
and U46790 (N_46790,N_46533,N_46500);
nor U46791 (N_46791,N_46643,N_46693);
nand U46792 (N_46792,N_46540,N_46668);
or U46793 (N_46793,N_46636,N_46574);
nand U46794 (N_46794,N_46631,N_46522);
nor U46795 (N_46795,N_46517,N_46721);
nand U46796 (N_46796,N_46746,N_46674);
nor U46797 (N_46797,N_46646,N_46587);
or U46798 (N_46798,N_46714,N_46697);
nor U46799 (N_46799,N_46741,N_46688);
nand U46800 (N_46800,N_46705,N_46507);
nor U46801 (N_46801,N_46634,N_46655);
xor U46802 (N_46802,N_46629,N_46737);
nand U46803 (N_46803,N_46621,N_46543);
xnor U46804 (N_46804,N_46590,N_46700);
or U46805 (N_46805,N_46589,N_46550);
nor U46806 (N_46806,N_46691,N_46568);
and U46807 (N_46807,N_46725,N_46551);
xor U46808 (N_46808,N_46528,N_46662);
and U46809 (N_46809,N_46665,N_46642);
and U46810 (N_46810,N_46699,N_46682);
or U46811 (N_46811,N_46702,N_46709);
or U46812 (N_46812,N_46565,N_46625);
nor U46813 (N_46813,N_46652,N_46524);
nand U46814 (N_46814,N_46657,N_46604);
xor U46815 (N_46815,N_46719,N_46529);
and U46816 (N_46816,N_46644,N_46745);
and U46817 (N_46817,N_46505,N_46577);
or U46818 (N_46818,N_46521,N_46640);
nor U46819 (N_46819,N_46503,N_46580);
nand U46820 (N_46820,N_46734,N_46600);
nor U46821 (N_46821,N_46516,N_46534);
xnor U46822 (N_46822,N_46537,N_46515);
xnor U46823 (N_46823,N_46523,N_46698);
and U46824 (N_46824,N_46716,N_46585);
nand U46825 (N_46825,N_46538,N_46658);
nand U46826 (N_46826,N_46501,N_46749);
xnor U46827 (N_46827,N_46694,N_46731);
or U46828 (N_46828,N_46663,N_46603);
or U46829 (N_46829,N_46739,N_46539);
nor U46830 (N_46830,N_46681,N_46616);
nor U46831 (N_46831,N_46675,N_46612);
or U46832 (N_46832,N_46591,N_46549);
nand U46833 (N_46833,N_46701,N_46623);
or U46834 (N_46834,N_46678,N_46624);
nor U46835 (N_46835,N_46672,N_46704);
nor U46836 (N_46836,N_46546,N_46676);
and U46837 (N_46837,N_46639,N_46569);
or U46838 (N_46838,N_46615,N_46650);
nand U46839 (N_46839,N_46610,N_46563);
nor U46840 (N_46840,N_46582,N_46748);
xor U46841 (N_46841,N_46607,N_46706);
or U46842 (N_46842,N_46724,N_46661);
nor U46843 (N_46843,N_46695,N_46689);
nor U46844 (N_46844,N_46531,N_46648);
nand U46845 (N_46845,N_46703,N_46594);
nand U46846 (N_46846,N_46514,N_46575);
nor U46847 (N_46847,N_46611,N_46638);
or U46848 (N_46848,N_46597,N_46671);
nor U46849 (N_46849,N_46556,N_46732);
nor U46850 (N_46850,N_46619,N_46617);
and U46851 (N_46851,N_46606,N_46717);
nor U46852 (N_46852,N_46669,N_46510);
nor U46853 (N_46853,N_46502,N_46647);
or U46854 (N_46854,N_46626,N_46713);
nand U46855 (N_46855,N_46679,N_46566);
nand U46856 (N_46856,N_46572,N_46601);
xor U46857 (N_46857,N_46747,N_46680);
xnor U46858 (N_46858,N_46525,N_46667);
or U46859 (N_46859,N_46609,N_46558);
and U46860 (N_46860,N_46696,N_46530);
nand U46861 (N_46861,N_46738,N_46744);
or U46862 (N_46862,N_46735,N_46718);
nand U46863 (N_46863,N_46602,N_46614);
and U46864 (N_46864,N_46586,N_46608);
or U46865 (N_46865,N_46571,N_46630);
xor U46866 (N_46866,N_46584,N_46512);
xor U46867 (N_46867,N_46645,N_46583);
nand U46868 (N_46868,N_46535,N_46520);
nor U46869 (N_46869,N_46561,N_46559);
nor U46870 (N_46870,N_46637,N_46527);
nor U46871 (N_46871,N_46664,N_46687);
xnor U46872 (N_46872,N_46545,N_46685);
or U46873 (N_46873,N_46653,N_46733);
or U46874 (N_46874,N_46532,N_46598);
nor U46875 (N_46875,N_46539,N_46605);
xor U46876 (N_46876,N_46582,N_46646);
and U46877 (N_46877,N_46600,N_46690);
xor U46878 (N_46878,N_46692,N_46577);
or U46879 (N_46879,N_46549,N_46714);
and U46880 (N_46880,N_46736,N_46603);
xor U46881 (N_46881,N_46569,N_46725);
xor U46882 (N_46882,N_46507,N_46720);
and U46883 (N_46883,N_46556,N_46508);
nor U46884 (N_46884,N_46732,N_46719);
and U46885 (N_46885,N_46598,N_46571);
and U46886 (N_46886,N_46657,N_46601);
nor U46887 (N_46887,N_46629,N_46601);
xnor U46888 (N_46888,N_46727,N_46707);
xor U46889 (N_46889,N_46588,N_46537);
xor U46890 (N_46890,N_46660,N_46632);
nand U46891 (N_46891,N_46612,N_46668);
nor U46892 (N_46892,N_46571,N_46723);
and U46893 (N_46893,N_46723,N_46704);
or U46894 (N_46894,N_46536,N_46543);
nand U46895 (N_46895,N_46601,N_46529);
nor U46896 (N_46896,N_46719,N_46601);
or U46897 (N_46897,N_46658,N_46596);
nor U46898 (N_46898,N_46547,N_46719);
nand U46899 (N_46899,N_46513,N_46587);
or U46900 (N_46900,N_46607,N_46617);
nand U46901 (N_46901,N_46519,N_46616);
nand U46902 (N_46902,N_46707,N_46518);
and U46903 (N_46903,N_46520,N_46734);
xor U46904 (N_46904,N_46614,N_46674);
nand U46905 (N_46905,N_46675,N_46638);
and U46906 (N_46906,N_46686,N_46592);
or U46907 (N_46907,N_46509,N_46560);
nand U46908 (N_46908,N_46746,N_46673);
xnor U46909 (N_46909,N_46599,N_46703);
or U46910 (N_46910,N_46704,N_46700);
and U46911 (N_46911,N_46515,N_46603);
or U46912 (N_46912,N_46534,N_46585);
nor U46913 (N_46913,N_46539,N_46578);
nand U46914 (N_46914,N_46657,N_46680);
nor U46915 (N_46915,N_46735,N_46505);
xor U46916 (N_46916,N_46623,N_46603);
and U46917 (N_46917,N_46579,N_46583);
or U46918 (N_46918,N_46564,N_46589);
and U46919 (N_46919,N_46554,N_46560);
xnor U46920 (N_46920,N_46699,N_46593);
nand U46921 (N_46921,N_46544,N_46518);
and U46922 (N_46922,N_46683,N_46727);
or U46923 (N_46923,N_46578,N_46541);
xor U46924 (N_46924,N_46626,N_46618);
or U46925 (N_46925,N_46522,N_46570);
nand U46926 (N_46926,N_46531,N_46668);
and U46927 (N_46927,N_46565,N_46626);
xnor U46928 (N_46928,N_46742,N_46598);
xor U46929 (N_46929,N_46583,N_46673);
nor U46930 (N_46930,N_46703,N_46598);
or U46931 (N_46931,N_46613,N_46554);
xnor U46932 (N_46932,N_46510,N_46603);
nor U46933 (N_46933,N_46662,N_46536);
or U46934 (N_46934,N_46515,N_46503);
nor U46935 (N_46935,N_46515,N_46527);
nand U46936 (N_46936,N_46693,N_46741);
xnor U46937 (N_46937,N_46732,N_46525);
and U46938 (N_46938,N_46722,N_46662);
xor U46939 (N_46939,N_46639,N_46509);
nor U46940 (N_46940,N_46738,N_46587);
nor U46941 (N_46941,N_46656,N_46673);
and U46942 (N_46942,N_46551,N_46732);
or U46943 (N_46943,N_46608,N_46653);
xor U46944 (N_46944,N_46685,N_46679);
nor U46945 (N_46945,N_46614,N_46541);
nor U46946 (N_46946,N_46521,N_46625);
and U46947 (N_46947,N_46644,N_46562);
and U46948 (N_46948,N_46717,N_46647);
nand U46949 (N_46949,N_46648,N_46621);
nand U46950 (N_46950,N_46571,N_46577);
nor U46951 (N_46951,N_46712,N_46738);
and U46952 (N_46952,N_46621,N_46725);
nand U46953 (N_46953,N_46531,N_46522);
and U46954 (N_46954,N_46566,N_46654);
nor U46955 (N_46955,N_46719,N_46550);
xor U46956 (N_46956,N_46690,N_46627);
nor U46957 (N_46957,N_46642,N_46675);
and U46958 (N_46958,N_46503,N_46706);
and U46959 (N_46959,N_46665,N_46743);
xnor U46960 (N_46960,N_46709,N_46658);
nand U46961 (N_46961,N_46562,N_46560);
nand U46962 (N_46962,N_46741,N_46544);
or U46963 (N_46963,N_46620,N_46635);
xnor U46964 (N_46964,N_46541,N_46670);
or U46965 (N_46965,N_46669,N_46715);
nand U46966 (N_46966,N_46743,N_46711);
nand U46967 (N_46967,N_46661,N_46572);
or U46968 (N_46968,N_46711,N_46526);
nand U46969 (N_46969,N_46518,N_46706);
nor U46970 (N_46970,N_46664,N_46545);
xor U46971 (N_46971,N_46532,N_46539);
nor U46972 (N_46972,N_46593,N_46671);
nor U46973 (N_46973,N_46530,N_46686);
nand U46974 (N_46974,N_46708,N_46508);
or U46975 (N_46975,N_46599,N_46564);
and U46976 (N_46976,N_46695,N_46509);
or U46977 (N_46977,N_46682,N_46540);
nor U46978 (N_46978,N_46702,N_46527);
nand U46979 (N_46979,N_46741,N_46636);
nor U46980 (N_46980,N_46590,N_46702);
and U46981 (N_46981,N_46561,N_46531);
xnor U46982 (N_46982,N_46649,N_46674);
nand U46983 (N_46983,N_46659,N_46519);
nand U46984 (N_46984,N_46639,N_46504);
or U46985 (N_46985,N_46557,N_46715);
and U46986 (N_46986,N_46576,N_46509);
or U46987 (N_46987,N_46535,N_46550);
or U46988 (N_46988,N_46524,N_46522);
and U46989 (N_46989,N_46690,N_46529);
and U46990 (N_46990,N_46506,N_46510);
xnor U46991 (N_46991,N_46577,N_46705);
nand U46992 (N_46992,N_46676,N_46605);
and U46993 (N_46993,N_46676,N_46707);
and U46994 (N_46994,N_46576,N_46701);
or U46995 (N_46995,N_46700,N_46516);
and U46996 (N_46996,N_46648,N_46564);
nor U46997 (N_46997,N_46607,N_46576);
nor U46998 (N_46998,N_46500,N_46510);
nor U46999 (N_46999,N_46695,N_46610);
and U47000 (N_47000,N_46873,N_46781);
and U47001 (N_47001,N_46933,N_46851);
xnor U47002 (N_47002,N_46960,N_46845);
nand U47003 (N_47003,N_46903,N_46794);
nand U47004 (N_47004,N_46853,N_46802);
nand U47005 (N_47005,N_46756,N_46917);
and U47006 (N_47006,N_46982,N_46833);
and U47007 (N_47007,N_46754,N_46855);
nor U47008 (N_47008,N_46818,N_46950);
and U47009 (N_47009,N_46866,N_46963);
xnor U47010 (N_47010,N_46916,N_46809);
or U47011 (N_47011,N_46790,N_46772);
nand U47012 (N_47012,N_46951,N_46832);
xnor U47013 (N_47013,N_46762,N_46997);
and U47014 (N_47014,N_46959,N_46806);
nand U47015 (N_47015,N_46848,N_46860);
nand U47016 (N_47016,N_46890,N_46911);
xnor U47017 (N_47017,N_46760,N_46824);
xnor U47018 (N_47018,N_46887,N_46808);
nand U47019 (N_47019,N_46952,N_46977);
nand U47020 (N_47020,N_46953,N_46944);
and U47021 (N_47021,N_46861,N_46787);
xnor U47022 (N_47022,N_46966,N_46888);
nand U47023 (N_47023,N_46918,N_46976);
nand U47024 (N_47024,N_46989,N_46862);
nor U47025 (N_47025,N_46967,N_46858);
nand U47026 (N_47026,N_46948,N_46821);
and U47027 (N_47027,N_46854,N_46786);
nor U47028 (N_47028,N_46978,N_46990);
nor U47029 (N_47029,N_46767,N_46882);
or U47030 (N_47030,N_46949,N_46840);
or U47031 (N_47031,N_46900,N_46946);
xor U47032 (N_47032,N_46773,N_46938);
nand U47033 (N_47033,N_46896,N_46765);
nor U47034 (N_47034,N_46912,N_46969);
nand U47035 (N_47035,N_46807,N_46926);
or U47036 (N_47036,N_46775,N_46774);
xnor U47037 (N_47037,N_46909,N_46995);
nand U47038 (N_47038,N_46906,N_46752);
nand U47039 (N_47039,N_46919,N_46972);
nand U47040 (N_47040,N_46799,N_46834);
or U47041 (N_47041,N_46849,N_46962);
xnor U47042 (N_47042,N_46889,N_46788);
xor U47043 (N_47043,N_46867,N_46979);
and U47044 (N_47044,N_46935,N_46886);
nor U47045 (N_47045,N_46898,N_46954);
or U47046 (N_47046,N_46884,N_46871);
xor U47047 (N_47047,N_46914,N_46863);
xor U47048 (N_47048,N_46936,N_46784);
nand U47049 (N_47049,N_46941,N_46856);
and U47050 (N_47050,N_46757,N_46876);
and U47051 (N_47051,N_46750,N_46835);
xor U47052 (N_47052,N_46846,N_46779);
xor U47053 (N_47053,N_46928,N_46811);
nor U47054 (N_47054,N_46793,N_46920);
and U47055 (N_47055,N_46796,N_46769);
nand U47056 (N_47056,N_46838,N_46828);
or U47057 (N_47057,N_46885,N_46763);
or U47058 (N_47058,N_46829,N_46870);
or U47059 (N_47059,N_46819,N_46910);
or U47060 (N_47060,N_46820,N_46764);
xnor U47061 (N_47061,N_46998,N_46837);
or U47062 (N_47062,N_46991,N_46894);
and U47063 (N_47063,N_46785,N_46907);
and U47064 (N_47064,N_46927,N_46815);
and U47065 (N_47065,N_46899,N_46847);
nor U47066 (N_47066,N_46755,N_46973);
nand U47067 (N_47067,N_46924,N_46999);
and U47068 (N_47068,N_46804,N_46816);
and U47069 (N_47069,N_46922,N_46874);
nand U47070 (N_47070,N_46823,N_46932);
and U47071 (N_47071,N_46805,N_46956);
nand U47072 (N_47072,N_46825,N_46993);
nand U47073 (N_47073,N_46822,N_46942);
or U47074 (N_47074,N_46988,N_46893);
nor U47075 (N_47075,N_46992,N_46766);
nor U47076 (N_47076,N_46843,N_46925);
nand U47077 (N_47077,N_46761,N_46996);
xnor U47078 (N_47078,N_46868,N_46872);
and U47079 (N_47079,N_46880,N_46751);
nand U47080 (N_47080,N_46844,N_46891);
or U47081 (N_47081,N_46957,N_46929);
nor U47082 (N_47082,N_46826,N_46778);
xor U47083 (N_47083,N_46897,N_46810);
nor U47084 (N_47084,N_46883,N_46792);
xnor U47085 (N_47085,N_46813,N_46961);
xnor U47086 (N_47086,N_46994,N_46913);
nor U47087 (N_47087,N_46817,N_46939);
and U47088 (N_47088,N_46943,N_46937);
nand U47089 (N_47089,N_46955,N_46812);
and U47090 (N_47090,N_46798,N_46892);
or U47091 (N_47091,N_46921,N_46859);
nand U47092 (N_47092,N_46789,N_46841);
or U47093 (N_47093,N_46968,N_46881);
nand U47094 (N_47094,N_46852,N_46947);
or U47095 (N_47095,N_46777,N_46970);
nand U47096 (N_47096,N_46895,N_46800);
and U47097 (N_47097,N_46864,N_46902);
nor U47098 (N_47098,N_46770,N_46865);
or U47099 (N_47099,N_46827,N_46836);
xor U47100 (N_47100,N_46964,N_46879);
and U47101 (N_47101,N_46759,N_46877);
xor U47102 (N_47102,N_46975,N_46839);
nor U47103 (N_47103,N_46797,N_46878);
and U47104 (N_47104,N_46830,N_46987);
or U47105 (N_47105,N_46958,N_46753);
nand U47106 (N_47106,N_46930,N_46869);
xor U47107 (N_47107,N_46814,N_46901);
nor U47108 (N_47108,N_46904,N_46842);
nor U47109 (N_47109,N_46965,N_46780);
and U47110 (N_47110,N_46980,N_46908);
or U47111 (N_47111,N_46791,N_46831);
nor U47112 (N_47112,N_46974,N_46984);
xnor U47113 (N_47113,N_46986,N_46801);
and U47114 (N_47114,N_46776,N_46758);
nor U47115 (N_47115,N_46981,N_46923);
xnor U47116 (N_47116,N_46783,N_46905);
nor U47117 (N_47117,N_46985,N_46945);
or U47118 (N_47118,N_46857,N_46971);
nor U47119 (N_47119,N_46803,N_46915);
nor U47120 (N_47120,N_46931,N_46940);
nand U47121 (N_47121,N_46934,N_46768);
nor U47122 (N_47122,N_46771,N_46850);
or U47123 (N_47123,N_46983,N_46875);
xnor U47124 (N_47124,N_46795,N_46782);
or U47125 (N_47125,N_46752,N_46821);
or U47126 (N_47126,N_46971,N_46908);
nor U47127 (N_47127,N_46978,N_46814);
or U47128 (N_47128,N_46813,N_46946);
nor U47129 (N_47129,N_46834,N_46995);
nand U47130 (N_47130,N_46767,N_46964);
and U47131 (N_47131,N_46966,N_46973);
or U47132 (N_47132,N_46912,N_46833);
nor U47133 (N_47133,N_46886,N_46845);
xnor U47134 (N_47134,N_46848,N_46844);
nand U47135 (N_47135,N_46846,N_46767);
xor U47136 (N_47136,N_46790,N_46796);
and U47137 (N_47137,N_46799,N_46879);
or U47138 (N_47138,N_46933,N_46876);
or U47139 (N_47139,N_46829,N_46986);
and U47140 (N_47140,N_46844,N_46853);
and U47141 (N_47141,N_46961,N_46751);
xor U47142 (N_47142,N_46821,N_46964);
or U47143 (N_47143,N_46979,N_46975);
nor U47144 (N_47144,N_46999,N_46876);
nand U47145 (N_47145,N_46962,N_46998);
nor U47146 (N_47146,N_46966,N_46833);
nor U47147 (N_47147,N_46842,N_46987);
nor U47148 (N_47148,N_46855,N_46850);
nand U47149 (N_47149,N_46797,N_46795);
xnor U47150 (N_47150,N_46996,N_46983);
xnor U47151 (N_47151,N_46869,N_46818);
nor U47152 (N_47152,N_46873,N_46852);
nand U47153 (N_47153,N_46871,N_46765);
nand U47154 (N_47154,N_46970,N_46904);
xnor U47155 (N_47155,N_46831,N_46918);
xnor U47156 (N_47156,N_46829,N_46927);
and U47157 (N_47157,N_46796,N_46953);
or U47158 (N_47158,N_46965,N_46812);
and U47159 (N_47159,N_46758,N_46935);
and U47160 (N_47160,N_46852,N_46750);
nand U47161 (N_47161,N_46971,N_46969);
xnor U47162 (N_47162,N_46926,N_46850);
or U47163 (N_47163,N_46823,N_46752);
nand U47164 (N_47164,N_46852,N_46936);
nand U47165 (N_47165,N_46851,N_46958);
and U47166 (N_47166,N_46820,N_46949);
nor U47167 (N_47167,N_46928,N_46861);
nor U47168 (N_47168,N_46763,N_46783);
nand U47169 (N_47169,N_46910,N_46911);
and U47170 (N_47170,N_46879,N_46850);
or U47171 (N_47171,N_46910,N_46817);
and U47172 (N_47172,N_46982,N_46938);
xor U47173 (N_47173,N_46787,N_46978);
nor U47174 (N_47174,N_46853,N_46937);
nor U47175 (N_47175,N_46994,N_46976);
nor U47176 (N_47176,N_46793,N_46997);
nand U47177 (N_47177,N_46837,N_46829);
nand U47178 (N_47178,N_46865,N_46786);
xor U47179 (N_47179,N_46799,N_46838);
xor U47180 (N_47180,N_46906,N_46813);
xnor U47181 (N_47181,N_46774,N_46797);
and U47182 (N_47182,N_46817,N_46820);
or U47183 (N_47183,N_46967,N_46817);
and U47184 (N_47184,N_46836,N_46999);
nor U47185 (N_47185,N_46892,N_46897);
nand U47186 (N_47186,N_46993,N_46954);
nor U47187 (N_47187,N_46829,N_46938);
nand U47188 (N_47188,N_46959,N_46767);
nand U47189 (N_47189,N_46752,N_46859);
and U47190 (N_47190,N_46809,N_46991);
nand U47191 (N_47191,N_46924,N_46952);
nand U47192 (N_47192,N_46861,N_46992);
and U47193 (N_47193,N_46773,N_46855);
or U47194 (N_47194,N_46973,N_46855);
nand U47195 (N_47195,N_46790,N_46935);
nand U47196 (N_47196,N_46949,N_46963);
nand U47197 (N_47197,N_46969,N_46945);
nor U47198 (N_47198,N_46802,N_46883);
xor U47199 (N_47199,N_46899,N_46848);
or U47200 (N_47200,N_46799,N_46950);
xnor U47201 (N_47201,N_46939,N_46974);
nand U47202 (N_47202,N_46868,N_46807);
nor U47203 (N_47203,N_46822,N_46986);
xor U47204 (N_47204,N_46890,N_46938);
nor U47205 (N_47205,N_46926,N_46904);
xor U47206 (N_47206,N_46957,N_46897);
nor U47207 (N_47207,N_46865,N_46853);
nor U47208 (N_47208,N_46858,N_46881);
xor U47209 (N_47209,N_46770,N_46932);
and U47210 (N_47210,N_46764,N_46849);
nor U47211 (N_47211,N_46817,N_46848);
nor U47212 (N_47212,N_46809,N_46846);
or U47213 (N_47213,N_46920,N_46921);
xnor U47214 (N_47214,N_46765,N_46761);
nand U47215 (N_47215,N_46795,N_46853);
nand U47216 (N_47216,N_46937,N_46768);
xnor U47217 (N_47217,N_46783,N_46825);
nor U47218 (N_47218,N_46868,N_46806);
and U47219 (N_47219,N_46866,N_46864);
and U47220 (N_47220,N_46825,N_46798);
xor U47221 (N_47221,N_46857,N_46865);
and U47222 (N_47222,N_46779,N_46781);
nand U47223 (N_47223,N_46870,N_46905);
or U47224 (N_47224,N_46958,N_46825);
xor U47225 (N_47225,N_46950,N_46882);
nand U47226 (N_47226,N_46968,N_46849);
nand U47227 (N_47227,N_46888,N_46946);
and U47228 (N_47228,N_46929,N_46773);
nand U47229 (N_47229,N_46867,N_46957);
or U47230 (N_47230,N_46902,N_46777);
or U47231 (N_47231,N_46815,N_46824);
xor U47232 (N_47232,N_46822,N_46752);
nor U47233 (N_47233,N_46833,N_46778);
or U47234 (N_47234,N_46815,N_46756);
or U47235 (N_47235,N_46898,N_46851);
or U47236 (N_47236,N_46901,N_46799);
and U47237 (N_47237,N_46841,N_46918);
nor U47238 (N_47238,N_46881,N_46922);
and U47239 (N_47239,N_46833,N_46792);
xor U47240 (N_47240,N_46871,N_46908);
nor U47241 (N_47241,N_46875,N_46804);
xor U47242 (N_47242,N_46771,N_46787);
and U47243 (N_47243,N_46783,N_46856);
nand U47244 (N_47244,N_46922,N_46784);
and U47245 (N_47245,N_46851,N_46838);
nand U47246 (N_47246,N_46791,N_46889);
nand U47247 (N_47247,N_46946,N_46894);
xor U47248 (N_47248,N_46847,N_46784);
and U47249 (N_47249,N_46756,N_46880);
and U47250 (N_47250,N_47208,N_47241);
and U47251 (N_47251,N_47151,N_47182);
nor U47252 (N_47252,N_47081,N_47043);
and U47253 (N_47253,N_47195,N_47082);
and U47254 (N_47254,N_47244,N_47114);
nand U47255 (N_47255,N_47227,N_47231);
and U47256 (N_47256,N_47073,N_47130);
nor U47257 (N_47257,N_47197,N_47121);
nor U47258 (N_47258,N_47229,N_47233);
xor U47259 (N_47259,N_47133,N_47041);
or U47260 (N_47260,N_47018,N_47023);
nand U47261 (N_47261,N_47185,N_47000);
or U47262 (N_47262,N_47074,N_47207);
xor U47263 (N_47263,N_47045,N_47052);
xor U47264 (N_47264,N_47174,N_47139);
nor U47265 (N_47265,N_47040,N_47015);
and U47266 (N_47266,N_47021,N_47149);
nand U47267 (N_47267,N_47028,N_47214);
xor U47268 (N_47268,N_47055,N_47078);
xor U47269 (N_47269,N_47030,N_47091);
and U47270 (N_47270,N_47228,N_47221);
or U47271 (N_47271,N_47198,N_47202);
or U47272 (N_47272,N_47215,N_47012);
and U47273 (N_47273,N_47039,N_47058);
nor U47274 (N_47274,N_47193,N_47016);
and U47275 (N_47275,N_47169,N_47076);
and U47276 (N_47276,N_47167,N_47051);
xnor U47277 (N_47277,N_47070,N_47180);
and U47278 (N_47278,N_47205,N_47104);
nand U47279 (N_47279,N_47099,N_47036);
nor U47280 (N_47280,N_47212,N_47173);
xor U47281 (N_47281,N_47145,N_47044);
or U47282 (N_47282,N_47237,N_47171);
or U47283 (N_47283,N_47084,N_47154);
or U47284 (N_47284,N_47129,N_47249);
nor U47285 (N_47285,N_47248,N_47068);
or U47286 (N_47286,N_47179,N_47006);
xnor U47287 (N_47287,N_47013,N_47218);
or U47288 (N_47288,N_47189,N_47005);
nor U47289 (N_47289,N_47163,N_47216);
xor U47290 (N_47290,N_47035,N_47062);
and U47291 (N_47291,N_47206,N_47141);
or U47292 (N_47292,N_47191,N_47155);
nor U47293 (N_47293,N_47079,N_47026);
and U47294 (N_47294,N_47022,N_47106);
nor U47295 (N_47295,N_47111,N_47232);
nor U47296 (N_47296,N_47222,N_47007);
and U47297 (N_47297,N_47042,N_47177);
and U47298 (N_47298,N_47083,N_47108);
and U47299 (N_47299,N_47020,N_47172);
xnor U47300 (N_47300,N_47008,N_47048);
xor U47301 (N_47301,N_47245,N_47032);
nand U47302 (N_47302,N_47019,N_47127);
xnor U47303 (N_47303,N_47029,N_47004);
or U47304 (N_47304,N_47053,N_47132);
nor U47305 (N_47305,N_47238,N_47120);
and U47306 (N_47306,N_47112,N_47162);
and U47307 (N_47307,N_47147,N_47211);
nand U47308 (N_47308,N_47164,N_47159);
or U47309 (N_47309,N_47090,N_47061);
nand U47310 (N_47310,N_47095,N_47085);
or U47311 (N_47311,N_47209,N_47246);
nor U47312 (N_47312,N_47200,N_47247);
and U47313 (N_47313,N_47033,N_47077);
or U47314 (N_47314,N_47158,N_47119);
nand U47315 (N_47315,N_47105,N_47025);
and U47316 (N_47316,N_47086,N_47188);
xnor U47317 (N_47317,N_47037,N_47092);
nor U47318 (N_47318,N_47064,N_47063);
xnor U47319 (N_47319,N_47134,N_47113);
and U47320 (N_47320,N_47181,N_47009);
xor U47321 (N_47321,N_47116,N_47156);
nand U47322 (N_47322,N_47034,N_47187);
nor U47323 (N_47323,N_47102,N_47240);
nand U47324 (N_47324,N_47183,N_47213);
and U47325 (N_47325,N_47176,N_47072);
or U47326 (N_47326,N_47242,N_47136);
nor U47327 (N_47327,N_47060,N_47153);
or U47328 (N_47328,N_47219,N_47002);
xnor U47329 (N_47329,N_47057,N_47087);
xnor U47330 (N_47330,N_47047,N_47031);
nor U47331 (N_47331,N_47075,N_47168);
nand U47332 (N_47332,N_47192,N_47160);
and U47333 (N_47333,N_47148,N_47201);
or U47334 (N_47334,N_47056,N_47103);
xor U47335 (N_47335,N_47146,N_47065);
and U47336 (N_47336,N_47128,N_47170);
nor U47337 (N_47337,N_47050,N_47080);
or U47338 (N_47338,N_47010,N_47093);
nand U47339 (N_47339,N_47003,N_47235);
or U47340 (N_47340,N_47194,N_47143);
and U47341 (N_47341,N_47017,N_47220);
or U47342 (N_47342,N_47117,N_47234);
or U47343 (N_47343,N_47125,N_47210);
or U47344 (N_47344,N_47178,N_47142);
xnor U47345 (N_47345,N_47027,N_47066);
xor U47346 (N_47346,N_47223,N_47165);
nor U47347 (N_47347,N_47049,N_47109);
nor U47348 (N_47348,N_47230,N_47097);
or U47349 (N_47349,N_47059,N_47225);
nor U47350 (N_47350,N_47089,N_47144);
nand U47351 (N_47351,N_47118,N_47126);
xnor U47352 (N_47352,N_47186,N_47152);
and U47353 (N_47353,N_47038,N_47199);
nor U47354 (N_47354,N_47098,N_47131);
xor U47355 (N_47355,N_47166,N_47150);
and U47356 (N_47356,N_47124,N_47140);
nand U47357 (N_47357,N_47024,N_47224);
or U47358 (N_47358,N_47243,N_47236);
nor U47359 (N_47359,N_47115,N_47101);
or U47360 (N_47360,N_47011,N_47123);
or U47361 (N_47361,N_47122,N_47094);
or U47362 (N_47362,N_47175,N_47226);
and U47363 (N_47363,N_47014,N_47107);
and U47364 (N_47364,N_47069,N_47096);
or U47365 (N_47365,N_47184,N_47138);
and U47366 (N_47366,N_47046,N_47137);
nand U47367 (N_47367,N_47217,N_47001);
xor U47368 (N_47368,N_47110,N_47190);
or U47369 (N_47369,N_47161,N_47203);
xor U47370 (N_47370,N_47239,N_47157);
nand U47371 (N_47371,N_47196,N_47100);
nor U47372 (N_47372,N_47067,N_47135);
xor U47373 (N_47373,N_47204,N_47088);
or U47374 (N_47374,N_47054,N_47071);
or U47375 (N_47375,N_47030,N_47113);
nand U47376 (N_47376,N_47231,N_47086);
and U47377 (N_47377,N_47113,N_47106);
nand U47378 (N_47378,N_47134,N_47135);
or U47379 (N_47379,N_47093,N_47214);
nand U47380 (N_47380,N_47211,N_47240);
nor U47381 (N_47381,N_47093,N_47083);
or U47382 (N_47382,N_47144,N_47006);
or U47383 (N_47383,N_47215,N_47168);
nor U47384 (N_47384,N_47237,N_47021);
xor U47385 (N_47385,N_47192,N_47091);
and U47386 (N_47386,N_47217,N_47060);
or U47387 (N_47387,N_47050,N_47235);
nor U47388 (N_47388,N_47130,N_47203);
or U47389 (N_47389,N_47135,N_47199);
xor U47390 (N_47390,N_47138,N_47132);
or U47391 (N_47391,N_47056,N_47151);
nor U47392 (N_47392,N_47040,N_47014);
nor U47393 (N_47393,N_47231,N_47195);
xor U47394 (N_47394,N_47097,N_47126);
nand U47395 (N_47395,N_47056,N_47096);
xor U47396 (N_47396,N_47212,N_47247);
and U47397 (N_47397,N_47213,N_47104);
or U47398 (N_47398,N_47226,N_47027);
nand U47399 (N_47399,N_47133,N_47167);
and U47400 (N_47400,N_47209,N_47142);
xor U47401 (N_47401,N_47103,N_47236);
or U47402 (N_47402,N_47166,N_47067);
nor U47403 (N_47403,N_47104,N_47105);
nor U47404 (N_47404,N_47025,N_47201);
nand U47405 (N_47405,N_47153,N_47233);
or U47406 (N_47406,N_47057,N_47217);
or U47407 (N_47407,N_47055,N_47020);
nand U47408 (N_47408,N_47158,N_47022);
nand U47409 (N_47409,N_47217,N_47069);
xnor U47410 (N_47410,N_47084,N_47246);
and U47411 (N_47411,N_47154,N_47156);
and U47412 (N_47412,N_47101,N_47107);
or U47413 (N_47413,N_47247,N_47183);
nor U47414 (N_47414,N_47244,N_47193);
nand U47415 (N_47415,N_47182,N_47174);
xor U47416 (N_47416,N_47232,N_47058);
nand U47417 (N_47417,N_47056,N_47057);
nand U47418 (N_47418,N_47110,N_47101);
and U47419 (N_47419,N_47244,N_47177);
or U47420 (N_47420,N_47068,N_47008);
and U47421 (N_47421,N_47073,N_47071);
and U47422 (N_47422,N_47040,N_47185);
and U47423 (N_47423,N_47058,N_47028);
nor U47424 (N_47424,N_47141,N_47009);
xor U47425 (N_47425,N_47128,N_47008);
or U47426 (N_47426,N_47186,N_47208);
nand U47427 (N_47427,N_47075,N_47087);
nor U47428 (N_47428,N_47248,N_47203);
or U47429 (N_47429,N_47190,N_47213);
xnor U47430 (N_47430,N_47042,N_47138);
xor U47431 (N_47431,N_47003,N_47008);
nor U47432 (N_47432,N_47002,N_47091);
xor U47433 (N_47433,N_47225,N_47072);
xnor U47434 (N_47434,N_47168,N_47219);
xor U47435 (N_47435,N_47109,N_47032);
nor U47436 (N_47436,N_47213,N_47090);
nand U47437 (N_47437,N_47024,N_47217);
xor U47438 (N_47438,N_47220,N_47154);
nand U47439 (N_47439,N_47099,N_47086);
or U47440 (N_47440,N_47125,N_47248);
or U47441 (N_47441,N_47050,N_47243);
nand U47442 (N_47442,N_47228,N_47163);
or U47443 (N_47443,N_47131,N_47021);
and U47444 (N_47444,N_47216,N_47211);
and U47445 (N_47445,N_47147,N_47087);
and U47446 (N_47446,N_47071,N_47077);
xor U47447 (N_47447,N_47001,N_47153);
nand U47448 (N_47448,N_47222,N_47002);
nand U47449 (N_47449,N_47177,N_47205);
nor U47450 (N_47450,N_47184,N_47200);
nand U47451 (N_47451,N_47235,N_47180);
nand U47452 (N_47452,N_47150,N_47146);
or U47453 (N_47453,N_47102,N_47029);
and U47454 (N_47454,N_47062,N_47090);
xnor U47455 (N_47455,N_47035,N_47005);
nor U47456 (N_47456,N_47147,N_47141);
or U47457 (N_47457,N_47113,N_47055);
nor U47458 (N_47458,N_47208,N_47203);
nor U47459 (N_47459,N_47213,N_47020);
xor U47460 (N_47460,N_47094,N_47017);
or U47461 (N_47461,N_47162,N_47128);
nor U47462 (N_47462,N_47240,N_47241);
nand U47463 (N_47463,N_47195,N_47128);
and U47464 (N_47464,N_47158,N_47129);
or U47465 (N_47465,N_47004,N_47116);
and U47466 (N_47466,N_47119,N_47193);
xor U47467 (N_47467,N_47060,N_47049);
nor U47468 (N_47468,N_47163,N_47101);
or U47469 (N_47469,N_47146,N_47018);
and U47470 (N_47470,N_47074,N_47015);
and U47471 (N_47471,N_47031,N_47011);
xnor U47472 (N_47472,N_47012,N_47162);
xnor U47473 (N_47473,N_47202,N_47201);
xnor U47474 (N_47474,N_47207,N_47166);
and U47475 (N_47475,N_47025,N_47078);
nand U47476 (N_47476,N_47044,N_47027);
and U47477 (N_47477,N_47042,N_47182);
nor U47478 (N_47478,N_47163,N_47121);
or U47479 (N_47479,N_47023,N_47138);
xnor U47480 (N_47480,N_47154,N_47038);
nand U47481 (N_47481,N_47063,N_47226);
xnor U47482 (N_47482,N_47166,N_47168);
xnor U47483 (N_47483,N_47116,N_47228);
or U47484 (N_47484,N_47077,N_47056);
and U47485 (N_47485,N_47022,N_47011);
nand U47486 (N_47486,N_47110,N_47167);
nand U47487 (N_47487,N_47203,N_47018);
nor U47488 (N_47488,N_47247,N_47079);
nand U47489 (N_47489,N_47111,N_47083);
or U47490 (N_47490,N_47078,N_47073);
nor U47491 (N_47491,N_47184,N_47146);
or U47492 (N_47492,N_47199,N_47063);
nor U47493 (N_47493,N_47042,N_47111);
xnor U47494 (N_47494,N_47080,N_47207);
nand U47495 (N_47495,N_47158,N_47192);
nor U47496 (N_47496,N_47152,N_47121);
xnor U47497 (N_47497,N_47182,N_47186);
nand U47498 (N_47498,N_47095,N_47055);
xor U47499 (N_47499,N_47148,N_47184);
or U47500 (N_47500,N_47455,N_47291);
nand U47501 (N_47501,N_47437,N_47279);
xor U47502 (N_47502,N_47469,N_47419);
or U47503 (N_47503,N_47485,N_47302);
nor U47504 (N_47504,N_47400,N_47314);
and U47505 (N_47505,N_47289,N_47316);
or U47506 (N_47506,N_47357,N_47466);
nand U47507 (N_47507,N_47348,N_47405);
nand U47508 (N_47508,N_47395,N_47346);
and U47509 (N_47509,N_47392,N_47262);
or U47510 (N_47510,N_47402,N_47491);
nand U47511 (N_47511,N_47382,N_47411);
nor U47512 (N_47512,N_47454,N_47322);
and U47513 (N_47513,N_47443,N_47494);
and U47514 (N_47514,N_47296,N_47353);
or U47515 (N_47515,N_47492,N_47299);
nor U47516 (N_47516,N_47452,N_47385);
and U47517 (N_47517,N_47301,N_47380);
or U47518 (N_47518,N_47265,N_47424);
nand U47519 (N_47519,N_47420,N_47343);
xor U47520 (N_47520,N_47376,N_47495);
nand U47521 (N_47521,N_47393,N_47375);
xor U47522 (N_47522,N_47497,N_47383);
xor U47523 (N_47523,N_47297,N_47363);
and U47524 (N_47524,N_47406,N_47251);
or U47525 (N_47525,N_47269,N_47445);
nor U47526 (N_47526,N_47471,N_47473);
or U47527 (N_47527,N_47447,N_47386);
nor U47528 (N_47528,N_47467,N_47446);
xor U47529 (N_47529,N_47464,N_47461);
nand U47530 (N_47530,N_47309,N_47440);
xnor U47531 (N_47531,N_47431,N_47428);
and U47532 (N_47532,N_47490,N_47426);
nor U47533 (N_47533,N_47499,N_47449);
and U47534 (N_47534,N_47336,N_47324);
nor U47535 (N_47535,N_47368,N_47276);
xnor U47536 (N_47536,N_47326,N_47480);
and U47537 (N_47537,N_47366,N_47468);
xor U47538 (N_47538,N_47481,N_47321);
xor U47539 (N_47539,N_47422,N_47441);
nand U47540 (N_47540,N_47329,N_47423);
and U47541 (N_47541,N_47408,N_47378);
and U47542 (N_47542,N_47381,N_47260);
nor U47543 (N_47543,N_47303,N_47401);
nand U47544 (N_47544,N_47493,N_47338);
nand U47545 (N_47545,N_47414,N_47367);
nand U47546 (N_47546,N_47475,N_47288);
and U47547 (N_47547,N_47365,N_47352);
xor U47548 (N_47548,N_47325,N_47281);
nor U47549 (N_47549,N_47263,N_47486);
nand U47550 (N_47550,N_47310,N_47427);
xor U47551 (N_47551,N_47472,N_47394);
and U47552 (N_47552,N_47295,N_47489);
xnor U47553 (N_47553,N_47470,N_47293);
nor U47554 (N_47554,N_47323,N_47388);
or U47555 (N_47555,N_47305,N_47369);
and U47556 (N_47556,N_47498,N_47258);
nand U47557 (N_47557,N_47341,N_47488);
nand U47558 (N_47558,N_47317,N_47355);
and U47559 (N_47559,N_47476,N_47404);
and U47560 (N_47560,N_47273,N_47478);
nor U47561 (N_47561,N_47290,N_47390);
and U47562 (N_47562,N_47415,N_47334);
nand U47563 (N_47563,N_47298,N_47274);
and U47564 (N_47564,N_47287,N_47278);
and U47565 (N_47565,N_47487,N_47474);
nand U47566 (N_47566,N_47407,N_47271);
nand U47567 (N_47567,N_47308,N_47362);
xor U47568 (N_47568,N_47379,N_47372);
nor U47569 (N_47569,N_47272,N_47425);
and U47570 (N_47570,N_47444,N_47284);
nor U47571 (N_47571,N_47280,N_47306);
and U47572 (N_47572,N_47257,N_47304);
nand U47573 (N_47573,N_47311,N_47389);
and U47574 (N_47574,N_47307,N_47433);
xnor U47575 (N_47575,N_47451,N_47384);
nand U47576 (N_47576,N_47370,N_47377);
or U47577 (N_47577,N_47320,N_47361);
and U47578 (N_47578,N_47403,N_47465);
nor U47579 (N_47579,N_47429,N_47391);
xor U47580 (N_47580,N_47268,N_47371);
xor U47581 (N_47581,N_47277,N_47267);
nor U47582 (N_47582,N_47459,N_47318);
and U47583 (N_47583,N_47270,N_47436);
nand U47584 (N_47584,N_47409,N_47477);
nor U47585 (N_47585,N_47337,N_47350);
or U47586 (N_47586,N_47250,N_47332);
nor U47587 (N_47587,N_47458,N_47315);
nand U47588 (N_47588,N_47434,N_47418);
and U47589 (N_47589,N_47416,N_47253);
xnor U47590 (N_47590,N_47432,N_47286);
nand U47591 (N_47591,N_47359,N_47300);
or U47592 (N_47592,N_47460,N_47259);
or U47593 (N_47593,N_47349,N_47364);
and U47594 (N_47594,N_47285,N_47435);
nor U47595 (N_47595,N_47342,N_47254);
xor U47596 (N_47596,N_47313,N_47453);
nand U47597 (N_47597,N_47327,N_47430);
nor U47598 (N_47598,N_47328,N_47331);
xnor U47599 (N_47599,N_47399,N_47484);
nor U47600 (N_47600,N_47312,N_47360);
xnor U47601 (N_47601,N_47374,N_47256);
nor U47602 (N_47602,N_47330,N_47261);
or U47603 (N_47603,N_47457,N_47417);
nor U47604 (N_47604,N_47396,N_47292);
nand U47605 (N_47605,N_47439,N_47345);
and U47606 (N_47606,N_47335,N_47387);
nand U47607 (N_47607,N_47339,N_47319);
and U47608 (N_47608,N_47354,N_47483);
nor U47609 (N_47609,N_47479,N_47294);
xor U47610 (N_47610,N_47410,N_47456);
xnor U47611 (N_47611,N_47442,N_47333);
and U47612 (N_47612,N_47496,N_47282);
nor U47613 (N_47613,N_47463,N_47340);
or U47614 (N_47614,N_47264,N_47421);
nand U47615 (N_47615,N_47373,N_47462);
or U47616 (N_47616,N_47438,N_47358);
nand U47617 (N_47617,N_47450,N_47255);
xnor U47618 (N_47618,N_47413,N_47351);
nand U47619 (N_47619,N_47482,N_47275);
or U47620 (N_47620,N_47266,N_47252);
nor U47621 (N_47621,N_47398,N_47344);
and U47622 (N_47622,N_47397,N_47412);
or U47623 (N_47623,N_47448,N_47347);
nor U47624 (N_47624,N_47283,N_47356);
nor U47625 (N_47625,N_47392,N_47489);
nand U47626 (N_47626,N_47340,N_47372);
xnor U47627 (N_47627,N_47433,N_47287);
or U47628 (N_47628,N_47400,N_47427);
or U47629 (N_47629,N_47254,N_47445);
or U47630 (N_47630,N_47254,N_47375);
or U47631 (N_47631,N_47344,N_47328);
and U47632 (N_47632,N_47364,N_47432);
nand U47633 (N_47633,N_47288,N_47483);
or U47634 (N_47634,N_47259,N_47481);
xnor U47635 (N_47635,N_47354,N_47267);
nor U47636 (N_47636,N_47428,N_47284);
and U47637 (N_47637,N_47328,N_47358);
nor U47638 (N_47638,N_47386,N_47311);
nor U47639 (N_47639,N_47342,N_47335);
nand U47640 (N_47640,N_47441,N_47285);
nand U47641 (N_47641,N_47422,N_47252);
or U47642 (N_47642,N_47449,N_47456);
or U47643 (N_47643,N_47320,N_47414);
xor U47644 (N_47644,N_47328,N_47313);
nand U47645 (N_47645,N_47483,N_47256);
and U47646 (N_47646,N_47415,N_47366);
or U47647 (N_47647,N_47422,N_47420);
nand U47648 (N_47648,N_47468,N_47309);
xnor U47649 (N_47649,N_47343,N_47291);
xor U47650 (N_47650,N_47323,N_47396);
xnor U47651 (N_47651,N_47325,N_47397);
nand U47652 (N_47652,N_47386,N_47266);
and U47653 (N_47653,N_47388,N_47274);
and U47654 (N_47654,N_47433,N_47372);
and U47655 (N_47655,N_47381,N_47436);
nand U47656 (N_47656,N_47270,N_47252);
nand U47657 (N_47657,N_47447,N_47266);
nor U47658 (N_47658,N_47499,N_47363);
nor U47659 (N_47659,N_47487,N_47351);
nand U47660 (N_47660,N_47306,N_47272);
or U47661 (N_47661,N_47321,N_47295);
or U47662 (N_47662,N_47425,N_47334);
or U47663 (N_47663,N_47401,N_47407);
or U47664 (N_47664,N_47250,N_47428);
or U47665 (N_47665,N_47331,N_47388);
nand U47666 (N_47666,N_47335,N_47369);
nand U47667 (N_47667,N_47498,N_47450);
and U47668 (N_47668,N_47374,N_47288);
and U47669 (N_47669,N_47438,N_47467);
or U47670 (N_47670,N_47379,N_47375);
xor U47671 (N_47671,N_47275,N_47423);
nand U47672 (N_47672,N_47296,N_47496);
nand U47673 (N_47673,N_47381,N_47469);
or U47674 (N_47674,N_47323,N_47478);
nor U47675 (N_47675,N_47404,N_47337);
nor U47676 (N_47676,N_47462,N_47364);
and U47677 (N_47677,N_47464,N_47336);
or U47678 (N_47678,N_47407,N_47481);
nand U47679 (N_47679,N_47410,N_47354);
or U47680 (N_47680,N_47380,N_47324);
and U47681 (N_47681,N_47343,N_47359);
nor U47682 (N_47682,N_47456,N_47294);
and U47683 (N_47683,N_47436,N_47398);
and U47684 (N_47684,N_47490,N_47304);
or U47685 (N_47685,N_47332,N_47267);
nand U47686 (N_47686,N_47347,N_47334);
nor U47687 (N_47687,N_47278,N_47279);
nand U47688 (N_47688,N_47396,N_47438);
nor U47689 (N_47689,N_47369,N_47468);
xnor U47690 (N_47690,N_47462,N_47298);
and U47691 (N_47691,N_47349,N_47469);
xnor U47692 (N_47692,N_47421,N_47364);
nand U47693 (N_47693,N_47339,N_47272);
or U47694 (N_47694,N_47465,N_47424);
nor U47695 (N_47695,N_47373,N_47260);
nor U47696 (N_47696,N_47457,N_47472);
or U47697 (N_47697,N_47442,N_47427);
or U47698 (N_47698,N_47326,N_47351);
xnor U47699 (N_47699,N_47281,N_47443);
nor U47700 (N_47700,N_47494,N_47276);
or U47701 (N_47701,N_47436,N_47422);
and U47702 (N_47702,N_47470,N_47490);
xor U47703 (N_47703,N_47254,N_47393);
or U47704 (N_47704,N_47325,N_47376);
and U47705 (N_47705,N_47443,N_47462);
nor U47706 (N_47706,N_47457,N_47306);
nand U47707 (N_47707,N_47426,N_47380);
nand U47708 (N_47708,N_47297,N_47393);
nor U47709 (N_47709,N_47483,N_47379);
nand U47710 (N_47710,N_47482,N_47477);
or U47711 (N_47711,N_47455,N_47330);
or U47712 (N_47712,N_47479,N_47484);
xor U47713 (N_47713,N_47337,N_47313);
or U47714 (N_47714,N_47433,N_47427);
or U47715 (N_47715,N_47426,N_47488);
nor U47716 (N_47716,N_47356,N_47306);
nor U47717 (N_47717,N_47430,N_47455);
or U47718 (N_47718,N_47303,N_47389);
xnor U47719 (N_47719,N_47384,N_47473);
nor U47720 (N_47720,N_47265,N_47404);
or U47721 (N_47721,N_47424,N_47371);
xnor U47722 (N_47722,N_47318,N_47361);
xnor U47723 (N_47723,N_47475,N_47267);
or U47724 (N_47724,N_47385,N_47456);
or U47725 (N_47725,N_47396,N_47378);
nand U47726 (N_47726,N_47363,N_47446);
nor U47727 (N_47727,N_47416,N_47492);
nor U47728 (N_47728,N_47350,N_47315);
nand U47729 (N_47729,N_47350,N_47347);
and U47730 (N_47730,N_47493,N_47324);
nor U47731 (N_47731,N_47250,N_47403);
or U47732 (N_47732,N_47274,N_47355);
xnor U47733 (N_47733,N_47345,N_47467);
nor U47734 (N_47734,N_47319,N_47268);
xor U47735 (N_47735,N_47485,N_47336);
nor U47736 (N_47736,N_47338,N_47326);
nor U47737 (N_47737,N_47422,N_47470);
nor U47738 (N_47738,N_47360,N_47361);
or U47739 (N_47739,N_47463,N_47305);
and U47740 (N_47740,N_47351,N_47386);
nand U47741 (N_47741,N_47450,N_47287);
nor U47742 (N_47742,N_47492,N_47334);
and U47743 (N_47743,N_47343,N_47269);
nor U47744 (N_47744,N_47495,N_47373);
xor U47745 (N_47745,N_47392,N_47251);
nand U47746 (N_47746,N_47282,N_47338);
or U47747 (N_47747,N_47364,N_47297);
and U47748 (N_47748,N_47345,N_47479);
nand U47749 (N_47749,N_47253,N_47427);
and U47750 (N_47750,N_47703,N_47552);
nand U47751 (N_47751,N_47673,N_47643);
nor U47752 (N_47752,N_47695,N_47551);
nor U47753 (N_47753,N_47610,N_47504);
and U47754 (N_47754,N_47585,N_47502);
nand U47755 (N_47755,N_47635,N_47580);
and U47756 (N_47756,N_47664,N_47640);
xor U47757 (N_47757,N_47656,N_47590);
nand U47758 (N_47758,N_47676,N_47633);
xnor U47759 (N_47759,N_47538,N_47732);
or U47760 (N_47760,N_47661,N_47639);
nor U47761 (N_47761,N_47745,N_47668);
or U47762 (N_47762,N_47748,N_47607);
nor U47763 (N_47763,N_47726,N_47540);
xor U47764 (N_47764,N_47677,N_47577);
nand U47765 (N_47765,N_47730,N_47563);
xor U47766 (N_47766,N_47518,N_47562);
nand U47767 (N_47767,N_47615,N_47687);
and U47768 (N_47768,N_47506,N_47729);
nor U47769 (N_47769,N_47605,N_47725);
nor U47770 (N_47770,N_47702,N_47681);
and U47771 (N_47771,N_47628,N_47644);
nand U47772 (N_47772,N_47549,N_47523);
or U47773 (N_47773,N_47537,N_47625);
xor U47774 (N_47774,N_47527,N_47684);
nand U47775 (N_47775,N_47561,N_47631);
nand U47776 (N_47776,N_47743,N_47682);
xor U47777 (N_47777,N_47581,N_47651);
nor U47778 (N_47778,N_47595,N_47742);
or U47779 (N_47779,N_47629,N_47622);
or U47780 (N_47780,N_47544,N_47569);
and U47781 (N_47781,N_47733,N_47530);
xor U47782 (N_47782,N_47621,N_47711);
or U47783 (N_47783,N_47637,N_47672);
and U47784 (N_47784,N_47571,N_47653);
or U47785 (N_47785,N_47611,N_47529);
xnor U47786 (N_47786,N_47578,N_47620);
or U47787 (N_47787,N_47604,N_47536);
and U47788 (N_47788,N_47565,N_47632);
nor U47789 (N_47789,N_47545,N_47626);
nand U47790 (N_47790,N_47613,N_47746);
nand U47791 (N_47791,N_47698,N_47624);
or U47792 (N_47792,N_47718,N_47557);
nand U47793 (N_47793,N_47704,N_47650);
or U47794 (N_47794,N_47596,N_47548);
or U47795 (N_47795,N_47511,N_47706);
nand U47796 (N_47796,N_47539,N_47696);
nand U47797 (N_47797,N_47707,N_47522);
nand U47798 (N_47798,N_47587,N_47679);
xnor U47799 (N_47799,N_47671,N_47597);
and U47800 (N_47800,N_47603,N_47659);
nor U47801 (N_47801,N_47609,N_47608);
xor U47802 (N_47802,N_47598,N_47560);
nor U47803 (N_47803,N_47734,N_47646);
nor U47804 (N_47804,N_47505,N_47737);
and U47805 (N_47805,N_47602,N_47614);
nor U47806 (N_47806,N_47749,N_47642);
nand U47807 (N_47807,N_47619,N_47573);
and U47808 (N_47808,N_47735,N_47747);
or U47809 (N_47809,N_47574,N_47520);
xor U47810 (N_47810,N_47701,N_47727);
nor U47811 (N_47811,N_47678,N_47591);
nor U47812 (N_47812,N_47712,N_47645);
nor U47813 (N_47813,N_47720,N_47666);
or U47814 (N_47814,N_47630,N_47547);
xnor U47815 (N_47815,N_47594,N_47713);
nor U47816 (N_47816,N_47508,N_47567);
xnor U47817 (N_47817,N_47623,N_47516);
nand U47818 (N_47818,N_47691,N_47510);
nor U47819 (N_47819,N_47665,N_47572);
or U47820 (N_47820,N_47667,N_47692);
nor U47821 (N_47821,N_47689,N_47709);
xnor U47822 (N_47822,N_47579,N_47641);
nand U47823 (N_47823,N_47513,N_47674);
and U47824 (N_47824,N_47638,N_47660);
or U47825 (N_47825,N_47584,N_47558);
xnor U47826 (N_47826,N_47546,N_47738);
or U47827 (N_47827,N_47503,N_47708);
nor U47828 (N_47828,N_47532,N_47501);
and U47829 (N_47829,N_47535,N_47583);
nand U47830 (N_47830,N_47740,N_47627);
nor U47831 (N_47831,N_47741,N_47568);
and U47832 (N_47832,N_47710,N_47570);
xor U47833 (N_47833,N_47582,N_47721);
or U47834 (N_47834,N_47699,N_47517);
nor U47835 (N_47835,N_47618,N_47533);
or U47836 (N_47836,N_47715,N_47512);
or U47837 (N_47837,N_47648,N_47556);
and U47838 (N_47838,N_47521,N_47575);
or U47839 (N_47839,N_47514,N_47680);
or U47840 (N_47840,N_47601,N_47550);
and U47841 (N_47841,N_47693,N_47526);
nand U47842 (N_47842,N_47599,N_47576);
or U47843 (N_47843,N_47600,N_47588);
or U47844 (N_47844,N_47524,N_47553);
or U47845 (N_47845,N_47700,N_47647);
xor U47846 (N_47846,N_47649,N_47688);
xnor U47847 (N_47847,N_47652,N_47714);
and U47848 (N_47848,N_47531,N_47606);
xor U47849 (N_47849,N_47685,N_47555);
and U47850 (N_47850,N_47564,N_47592);
nand U47851 (N_47851,N_47655,N_47654);
xnor U47852 (N_47852,N_47683,N_47705);
nor U47853 (N_47853,N_47543,N_47612);
nor U47854 (N_47854,N_47541,N_47559);
xnor U47855 (N_47855,N_47617,N_47719);
and U47856 (N_47856,N_47589,N_47739);
or U47857 (N_47857,N_47525,N_47593);
xor U47858 (N_47858,N_47686,N_47728);
or U47859 (N_47859,N_47519,N_47542);
nor U47860 (N_47860,N_47697,N_47669);
nand U47861 (N_47861,N_47586,N_47663);
nand U47862 (N_47862,N_47634,N_47736);
or U47863 (N_47863,N_47723,N_47509);
nand U47864 (N_47864,N_47507,N_47717);
nor U47865 (N_47865,N_47566,N_47636);
nor U47866 (N_47866,N_47515,N_47724);
nand U47867 (N_47867,N_47716,N_47731);
and U47868 (N_47868,N_47657,N_47616);
or U47869 (N_47869,N_47528,N_47500);
nand U47870 (N_47870,N_47694,N_47662);
xor U47871 (N_47871,N_47675,N_47744);
nand U47872 (N_47872,N_47670,N_47658);
xor U47873 (N_47873,N_47722,N_47534);
and U47874 (N_47874,N_47690,N_47554);
or U47875 (N_47875,N_47725,N_47666);
and U47876 (N_47876,N_47692,N_47594);
nor U47877 (N_47877,N_47521,N_47630);
xor U47878 (N_47878,N_47725,N_47742);
or U47879 (N_47879,N_47515,N_47608);
nand U47880 (N_47880,N_47582,N_47516);
or U47881 (N_47881,N_47507,N_47555);
nor U47882 (N_47882,N_47600,N_47745);
or U47883 (N_47883,N_47525,N_47568);
nor U47884 (N_47884,N_47535,N_47616);
or U47885 (N_47885,N_47537,N_47596);
nand U47886 (N_47886,N_47650,N_47509);
nand U47887 (N_47887,N_47602,N_47542);
and U47888 (N_47888,N_47585,N_47568);
nand U47889 (N_47889,N_47614,N_47716);
nand U47890 (N_47890,N_47591,N_47574);
nand U47891 (N_47891,N_47615,N_47658);
or U47892 (N_47892,N_47530,N_47721);
or U47893 (N_47893,N_47586,N_47745);
nor U47894 (N_47894,N_47609,N_47567);
or U47895 (N_47895,N_47748,N_47731);
nand U47896 (N_47896,N_47580,N_47646);
xnor U47897 (N_47897,N_47647,N_47654);
or U47898 (N_47898,N_47554,N_47534);
and U47899 (N_47899,N_47672,N_47650);
nor U47900 (N_47900,N_47510,N_47712);
xor U47901 (N_47901,N_47604,N_47694);
or U47902 (N_47902,N_47645,N_47626);
nor U47903 (N_47903,N_47515,N_47561);
or U47904 (N_47904,N_47577,N_47734);
nand U47905 (N_47905,N_47531,N_47735);
xnor U47906 (N_47906,N_47506,N_47726);
or U47907 (N_47907,N_47688,N_47653);
xnor U47908 (N_47908,N_47681,N_47614);
nor U47909 (N_47909,N_47639,N_47609);
nand U47910 (N_47910,N_47539,N_47700);
or U47911 (N_47911,N_47621,N_47678);
nand U47912 (N_47912,N_47559,N_47585);
and U47913 (N_47913,N_47649,N_47557);
and U47914 (N_47914,N_47691,N_47613);
or U47915 (N_47915,N_47637,N_47682);
xor U47916 (N_47916,N_47607,N_47717);
nor U47917 (N_47917,N_47684,N_47634);
nor U47918 (N_47918,N_47539,N_47603);
nand U47919 (N_47919,N_47642,N_47689);
and U47920 (N_47920,N_47622,N_47597);
nand U47921 (N_47921,N_47561,N_47624);
nor U47922 (N_47922,N_47533,N_47673);
nor U47923 (N_47923,N_47543,N_47572);
nor U47924 (N_47924,N_47702,N_47523);
xor U47925 (N_47925,N_47613,N_47589);
and U47926 (N_47926,N_47620,N_47628);
and U47927 (N_47927,N_47709,N_47539);
nand U47928 (N_47928,N_47733,N_47671);
and U47929 (N_47929,N_47741,N_47703);
nor U47930 (N_47930,N_47509,N_47517);
and U47931 (N_47931,N_47557,N_47519);
xnor U47932 (N_47932,N_47548,N_47512);
nand U47933 (N_47933,N_47527,N_47740);
xor U47934 (N_47934,N_47729,N_47626);
nand U47935 (N_47935,N_47533,N_47654);
xor U47936 (N_47936,N_47679,N_47536);
nor U47937 (N_47937,N_47569,N_47703);
xor U47938 (N_47938,N_47740,N_47678);
and U47939 (N_47939,N_47689,N_47576);
nor U47940 (N_47940,N_47745,N_47596);
nor U47941 (N_47941,N_47630,N_47574);
and U47942 (N_47942,N_47566,N_47538);
or U47943 (N_47943,N_47665,N_47560);
nand U47944 (N_47944,N_47558,N_47635);
nand U47945 (N_47945,N_47649,N_47589);
and U47946 (N_47946,N_47600,N_47743);
nor U47947 (N_47947,N_47529,N_47682);
xor U47948 (N_47948,N_47544,N_47718);
xor U47949 (N_47949,N_47625,N_47599);
or U47950 (N_47950,N_47737,N_47663);
nand U47951 (N_47951,N_47555,N_47502);
nand U47952 (N_47952,N_47630,N_47672);
nand U47953 (N_47953,N_47548,N_47672);
or U47954 (N_47954,N_47664,N_47533);
nand U47955 (N_47955,N_47703,N_47665);
nand U47956 (N_47956,N_47517,N_47528);
nand U47957 (N_47957,N_47710,N_47734);
or U47958 (N_47958,N_47556,N_47670);
xor U47959 (N_47959,N_47606,N_47626);
xor U47960 (N_47960,N_47668,N_47565);
or U47961 (N_47961,N_47525,N_47621);
and U47962 (N_47962,N_47640,N_47632);
nor U47963 (N_47963,N_47642,N_47522);
and U47964 (N_47964,N_47639,N_47548);
or U47965 (N_47965,N_47524,N_47549);
nor U47966 (N_47966,N_47530,N_47520);
or U47967 (N_47967,N_47599,N_47700);
nand U47968 (N_47968,N_47517,N_47690);
nand U47969 (N_47969,N_47529,N_47532);
nand U47970 (N_47970,N_47589,N_47721);
or U47971 (N_47971,N_47594,N_47513);
and U47972 (N_47972,N_47506,N_47643);
and U47973 (N_47973,N_47550,N_47534);
xnor U47974 (N_47974,N_47563,N_47547);
and U47975 (N_47975,N_47715,N_47508);
xnor U47976 (N_47976,N_47720,N_47596);
or U47977 (N_47977,N_47557,N_47558);
xnor U47978 (N_47978,N_47620,N_47509);
nand U47979 (N_47979,N_47683,N_47513);
and U47980 (N_47980,N_47747,N_47510);
or U47981 (N_47981,N_47577,N_47567);
nor U47982 (N_47982,N_47636,N_47650);
nand U47983 (N_47983,N_47631,N_47657);
xnor U47984 (N_47984,N_47556,N_47614);
and U47985 (N_47985,N_47686,N_47687);
xor U47986 (N_47986,N_47545,N_47649);
and U47987 (N_47987,N_47555,N_47548);
or U47988 (N_47988,N_47656,N_47647);
xnor U47989 (N_47989,N_47556,N_47532);
and U47990 (N_47990,N_47519,N_47582);
and U47991 (N_47991,N_47527,N_47516);
nand U47992 (N_47992,N_47647,N_47713);
nor U47993 (N_47993,N_47523,N_47628);
or U47994 (N_47994,N_47513,N_47536);
xor U47995 (N_47995,N_47650,N_47544);
nor U47996 (N_47996,N_47515,N_47595);
or U47997 (N_47997,N_47589,N_47741);
nor U47998 (N_47998,N_47743,N_47675);
nor U47999 (N_47999,N_47700,N_47584);
xor U48000 (N_48000,N_47817,N_47804);
and U48001 (N_48001,N_47768,N_47770);
nor U48002 (N_48002,N_47913,N_47823);
nand U48003 (N_48003,N_47959,N_47896);
or U48004 (N_48004,N_47938,N_47761);
or U48005 (N_48005,N_47919,N_47840);
nand U48006 (N_48006,N_47951,N_47971);
nand U48007 (N_48007,N_47925,N_47926);
xor U48008 (N_48008,N_47810,N_47859);
nor U48009 (N_48009,N_47750,N_47844);
nand U48010 (N_48010,N_47862,N_47942);
xnor U48011 (N_48011,N_47880,N_47993);
xnor U48012 (N_48012,N_47955,N_47991);
nor U48013 (N_48013,N_47910,N_47776);
and U48014 (N_48014,N_47820,N_47899);
nor U48015 (N_48015,N_47866,N_47774);
and U48016 (N_48016,N_47863,N_47924);
or U48017 (N_48017,N_47754,N_47867);
or U48018 (N_48018,N_47992,N_47763);
or U48019 (N_48019,N_47996,N_47802);
or U48020 (N_48020,N_47818,N_47846);
xnor U48021 (N_48021,N_47922,N_47794);
and U48022 (N_48022,N_47855,N_47758);
xor U48023 (N_48023,N_47895,N_47787);
xor U48024 (N_48024,N_47871,N_47915);
nand U48025 (N_48025,N_47962,N_47885);
nor U48026 (N_48026,N_47970,N_47829);
nand U48027 (N_48027,N_47958,N_47981);
and U48028 (N_48028,N_47904,N_47872);
xnor U48029 (N_48029,N_47850,N_47982);
xnor U48030 (N_48030,N_47916,N_47785);
and U48031 (N_48031,N_47997,N_47941);
nand U48032 (N_48032,N_47824,N_47886);
nand U48033 (N_48033,N_47994,N_47847);
nand U48034 (N_48034,N_47861,N_47799);
or U48035 (N_48035,N_47759,N_47827);
nor U48036 (N_48036,N_47778,N_47845);
or U48037 (N_48037,N_47858,N_47833);
nor U48038 (N_48038,N_47983,N_47979);
or U48039 (N_48039,N_47835,N_47821);
nor U48040 (N_48040,N_47936,N_47877);
xnor U48041 (N_48041,N_47832,N_47752);
xor U48042 (N_48042,N_47853,N_47826);
and U48043 (N_48043,N_47812,N_47813);
or U48044 (N_48044,N_47881,N_47811);
nor U48045 (N_48045,N_47753,N_47838);
nand U48046 (N_48046,N_47900,N_47920);
or U48047 (N_48047,N_47793,N_47999);
nor U48048 (N_48048,N_47909,N_47831);
and U48049 (N_48049,N_47894,N_47775);
nand U48050 (N_48050,N_47978,N_47888);
or U48051 (N_48051,N_47756,N_47966);
xnor U48052 (N_48052,N_47876,N_47998);
xor U48053 (N_48053,N_47932,N_47929);
nand U48054 (N_48054,N_47782,N_47908);
or U48055 (N_48055,N_47828,N_47977);
nor U48056 (N_48056,N_47949,N_47792);
nor U48057 (N_48057,N_47773,N_47819);
xor U48058 (N_48058,N_47825,N_47973);
nor U48059 (N_48059,N_47934,N_47954);
or U48060 (N_48060,N_47766,N_47907);
xor U48061 (N_48061,N_47995,N_47755);
nand U48062 (N_48062,N_47928,N_47972);
nand U48063 (N_48063,N_47807,N_47901);
xor U48064 (N_48064,N_47964,N_47976);
nand U48065 (N_48065,N_47987,N_47795);
nor U48066 (N_48066,N_47956,N_47854);
and U48067 (N_48067,N_47918,N_47751);
nand U48068 (N_48068,N_47891,N_47953);
nor U48069 (N_48069,N_47931,N_47937);
xnor U48070 (N_48070,N_47975,N_47914);
nor U48071 (N_48071,N_47765,N_47893);
xnor U48072 (N_48072,N_47961,N_47944);
and U48073 (N_48073,N_47767,N_47805);
xnor U48074 (N_48074,N_47798,N_47852);
nor U48075 (N_48075,N_47963,N_47809);
nand U48076 (N_48076,N_47988,N_47803);
or U48077 (N_48077,N_47797,N_47796);
nor U48078 (N_48078,N_47860,N_47839);
or U48079 (N_48079,N_47906,N_47801);
or U48080 (N_48080,N_47948,N_47874);
nand U48081 (N_48081,N_47757,N_47952);
nor U48082 (N_48082,N_47878,N_47923);
or U48083 (N_48083,N_47791,N_47869);
and U48084 (N_48084,N_47806,N_47887);
and U48085 (N_48085,N_47921,N_47892);
xnor U48086 (N_48086,N_47837,N_47902);
nand U48087 (N_48087,N_47815,N_47967);
and U48088 (N_48088,N_47890,N_47762);
nand U48089 (N_48089,N_47889,N_47764);
and U48090 (N_48090,N_47968,N_47879);
xor U48091 (N_48091,N_47911,N_47980);
or U48092 (N_48092,N_47769,N_47842);
xor U48093 (N_48093,N_47884,N_47781);
nor U48094 (N_48094,N_47865,N_47816);
xor U48095 (N_48095,N_47989,N_47783);
xnor U48096 (N_48096,N_47772,N_47822);
and U48097 (N_48097,N_47903,N_47974);
or U48098 (N_48098,N_47986,N_47830);
nand U48099 (N_48099,N_47912,N_47873);
and U48100 (N_48100,N_47950,N_47939);
nand U48101 (N_48101,N_47870,N_47933);
xor U48102 (N_48102,N_47905,N_47943);
nand U48103 (N_48103,N_47857,N_47848);
or U48104 (N_48104,N_47843,N_47984);
and U48105 (N_48105,N_47786,N_47882);
nand U48106 (N_48106,N_47836,N_47834);
xnor U48107 (N_48107,N_47969,N_47875);
xnor U48108 (N_48108,N_47841,N_47780);
or U48109 (N_48109,N_47897,N_47985);
or U48110 (N_48110,N_47849,N_47898);
and U48111 (N_48111,N_47779,N_47864);
nand U48112 (N_48112,N_47777,N_47760);
or U48113 (N_48113,N_47771,N_47784);
or U48114 (N_48114,N_47917,N_47930);
nand U48115 (N_48115,N_47957,N_47788);
or U48116 (N_48116,N_47856,N_47790);
and U48117 (N_48117,N_47960,N_47965);
nand U48118 (N_48118,N_47789,N_47851);
nor U48119 (N_48119,N_47800,N_47940);
nand U48120 (N_48120,N_47947,N_47883);
xnor U48121 (N_48121,N_47935,N_47868);
nor U48122 (N_48122,N_47808,N_47946);
xnor U48123 (N_48123,N_47927,N_47814);
nand U48124 (N_48124,N_47990,N_47945);
and U48125 (N_48125,N_47897,N_47941);
or U48126 (N_48126,N_47766,N_47833);
and U48127 (N_48127,N_47786,N_47862);
or U48128 (N_48128,N_47967,N_47776);
nor U48129 (N_48129,N_47761,N_47956);
nand U48130 (N_48130,N_47973,N_47814);
and U48131 (N_48131,N_47927,N_47774);
and U48132 (N_48132,N_47760,N_47790);
and U48133 (N_48133,N_47861,N_47946);
nand U48134 (N_48134,N_47761,N_47800);
nor U48135 (N_48135,N_47891,N_47796);
xnor U48136 (N_48136,N_47866,N_47876);
nand U48137 (N_48137,N_47965,N_47970);
nor U48138 (N_48138,N_47938,N_47931);
nand U48139 (N_48139,N_47772,N_47970);
or U48140 (N_48140,N_47975,N_47866);
xor U48141 (N_48141,N_47822,N_47776);
and U48142 (N_48142,N_47837,N_47967);
xor U48143 (N_48143,N_47864,N_47815);
and U48144 (N_48144,N_47836,N_47789);
or U48145 (N_48145,N_47825,N_47822);
nand U48146 (N_48146,N_47793,N_47908);
nand U48147 (N_48147,N_47804,N_47886);
nor U48148 (N_48148,N_47934,N_47966);
or U48149 (N_48149,N_47983,N_47961);
or U48150 (N_48150,N_47766,N_47882);
nand U48151 (N_48151,N_47946,N_47772);
xnor U48152 (N_48152,N_47987,N_47775);
nand U48153 (N_48153,N_47822,N_47828);
or U48154 (N_48154,N_47953,N_47930);
or U48155 (N_48155,N_47783,N_47778);
xor U48156 (N_48156,N_47990,N_47800);
nor U48157 (N_48157,N_47829,N_47893);
and U48158 (N_48158,N_47787,N_47816);
xor U48159 (N_48159,N_47932,N_47993);
nor U48160 (N_48160,N_47964,N_47884);
nor U48161 (N_48161,N_47980,N_47851);
xnor U48162 (N_48162,N_47898,N_47956);
and U48163 (N_48163,N_47842,N_47838);
nand U48164 (N_48164,N_47888,N_47849);
and U48165 (N_48165,N_47917,N_47761);
nor U48166 (N_48166,N_47813,N_47944);
xnor U48167 (N_48167,N_47792,N_47796);
or U48168 (N_48168,N_47789,N_47937);
and U48169 (N_48169,N_47885,N_47827);
nor U48170 (N_48170,N_47928,N_47920);
xor U48171 (N_48171,N_47942,N_47838);
nor U48172 (N_48172,N_47944,N_47873);
nor U48173 (N_48173,N_47787,N_47855);
nand U48174 (N_48174,N_47848,N_47893);
or U48175 (N_48175,N_47931,N_47979);
and U48176 (N_48176,N_47794,N_47998);
nor U48177 (N_48177,N_47940,N_47792);
or U48178 (N_48178,N_47919,N_47793);
or U48179 (N_48179,N_47956,N_47936);
or U48180 (N_48180,N_47848,N_47853);
and U48181 (N_48181,N_47992,N_47972);
and U48182 (N_48182,N_47959,N_47771);
nand U48183 (N_48183,N_47871,N_47793);
and U48184 (N_48184,N_47933,N_47830);
or U48185 (N_48185,N_47901,N_47955);
nor U48186 (N_48186,N_47830,N_47997);
and U48187 (N_48187,N_47791,N_47783);
and U48188 (N_48188,N_47829,N_47934);
nand U48189 (N_48189,N_47969,N_47850);
xnor U48190 (N_48190,N_47890,N_47879);
xor U48191 (N_48191,N_47786,N_47758);
or U48192 (N_48192,N_47869,N_47954);
and U48193 (N_48193,N_47959,N_47929);
xnor U48194 (N_48194,N_47814,N_47896);
xor U48195 (N_48195,N_47848,N_47995);
or U48196 (N_48196,N_47856,N_47829);
xor U48197 (N_48197,N_47875,N_47834);
nand U48198 (N_48198,N_47886,N_47887);
xnor U48199 (N_48199,N_47864,N_47936);
nor U48200 (N_48200,N_47759,N_47791);
and U48201 (N_48201,N_47844,N_47772);
nand U48202 (N_48202,N_47847,N_47849);
xor U48203 (N_48203,N_47764,N_47905);
nor U48204 (N_48204,N_47845,N_47952);
xor U48205 (N_48205,N_47994,N_47815);
xnor U48206 (N_48206,N_47770,N_47895);
nand U48207 (N_48207,N_47761,N_47826);
xor U48208 (N_48208,N_47991,N_47902);
nor U48209 (N_48209,N_47983,N_47965);
nor U48210 (N_48210,N_47902,N_47951);
nand U48211 (N_48211,N_47785,N_47990);
nand U48212 (N_48212,N_47905,N_47967);
nor U48213 (N_48213,N_47809,N_47758);
and U48214 (N_48214,N_47766,N_47782);
and U48215 (N_48215,N_47906,N_47928);
xor U48216 (N_48216,N_47914,N_47819);
nand U48217 (N_48217,N_47986,N_47918);
and U48218 (N_48218,N_47996,N_47984);
or U48219 (N_48219,N_47857,N_47832);
and U48220 (N_48220,N_47946,N_47900);
nand U48221 (N_48221,N_47849,N_47790);
and U48222 (N_48222,N_47991,N_47972);
xor U48223 (N_48223,N_47784,N_47899);
xnor U48224 (N_48224,N_47909,N_47849);
nor U48225 (N_48225,N_47812,N_47928);
or U48226 (N_48226,N_47896,N_47917);
nor U48227 (N_48227,N_47993,N_47897);
nand U48228 (N_48228,N_47764,N_47869);
nor U48229 (N_48229,N_47944,N_47900);
nand U48230 (N_48230,N_47911,N_47790);
or U48231 (N_48231,N_47865,N_47986);
xnor U48232 (N_48232,N_47802,N_47861);
nand U48233 (N_48233,N_47965,N_47923);
or U48234 (N_48234,N_47774,N_47896);
xor U48235 (N_48235,N_47753,N_47916);
and U48236 (N_48236,N_47818,N_47847);
nand U48237 (N_48237,N_47945,N_47852);
nor U48238 (N_48238,N_47873,N_47934);
and U48239 (N_48239,N_47809,N_47915);
and U48240 (N_48240,N_47819,N_47893);
nor U48241 (N_48241,N_47924,N_47959);
nor U48242 (N_48242,N_47873,N_47916);
xnor U48243 (N_48243,N_47861,N_47962);
or U48244 (N_48244,N_47900,N_47908);
nor U48245 (N_48245,N_47845,N_47859);
and U48246 (N_48246,N_47959,N_47759);
and U48247 (N_48247,N_47870,N_47993);
and U48248 (N_48248,N_47753,N_47872);
xor U48249 (N_48249,N_47984,N_47787);
nor U48250 (N_48250,N_48234,N_48105);
and U48251 (N_48251,N_48111,N_48049);
nand U48252 (N_48252,N_48216,N_48108);
nor U48253 (N_48253,N_48047,N_48177);
nand U48254 (N_48254,N_48221,N_48244);
or U48255 (N_48255,N_48018,N_48107);
xor U48256 (N_48256,N_48238,N_48205);
xnor U48257 (N_48257,N_48134,N_48008);
or U48258 (N_48258,N_48161,N_48157);
nand U48259 (N_48259,N_48182,N_48003);
and U48260 (N_48260,N_48053,N_48191);
nor U48261 (N_48261,N_48071,N_48204);
and U48262 (N_48262,N_48084,N_48214);
xor U48263 (N_48263,N_48009,N_48183);
or U48264 (N_48264,N_48167,N_48020);
and U48265 (N_48265,N_48110,N_48227);
and U48266 (N_48266,N_48101,N_48125);
nor U48267 (N_48267,N_48207,N_48029);
or U48268 (N_48268,N_48173,N_48141);
or U48269 (N_48269,N_48092,N_48233);
xor U48270 (N_48270,N_48129,N_48096);
nand U48271 (N_48271,N_48219,N_48210);
and U48272 (N_48272,N_48079,N_48147);
nand U48273 (N_48273,N_48225,N_48198);
or U48274 (N_48274,N_48061,N_48231);
nand U48275 (N_48275,N_48081,N_48247);
or U48276 (N_48276,N_48099,N_48013);
xnor U48277 (N_48277,N_48104,N_48056);
nand U48278 (N_48278,N_48067,N_48217);
nor U48279 (N_48279,N_48162,N_48033);
or U48280 (N_48280,N_48241,N_48039);
or U48281 (N_48281,N_48022,N_48041);
and U48282 (N_48282,N_48196,N_48048);
and U48283 (N_48283,N_48072,N_48117);
nor U48284 (N_48284,N_48232,N_48154);
and U48285 (N_48285,N_48121,N_48119);
nor U48286 (N_48286,N_48181,N_48188);
or U48287 (N_48287,N_48034,N_48103);
nand U48288 (N_48288,N_48069,N_48211);
nor U48289 (N_48289,N_48091,N_48059);
or U48290 (N_48290,N_48073,N_48058);
nor U48291 (N_48291,N_48136,N_48001);
xor U48292 (N_48292,N_48109,N_48124);
nor U48293 (N_48293,N_48040,N_48249);
nand U48294 (N_48294,N_48209,N_48195);
nand U48295 (N_48295,N_48206,N_48193);
and U48296 (N_48296,N_48045,N_48032);
nor U48297 (N_48297,N_48150,N_48128);
or U48298 (N_48298,N_48226,N_48122);
xor U48299 (N_48299,N_48131,N_48095);
or U48300 (N_48300,N_48021,N_48246);
and U48301 (N_48301,N_48007,N_48203);
or U48302 (N_48302,N_48153,N_48170);
or U48303 (N_48303,N_48126,N_48160);
nand U48304 (N_48304,N_48120,N_48236);
nand U48305 (N_48305,N_48215,N_48037);
nand U48306 (N_48306,N_48123,N_48023);
xnor U48307 (N_48307,N_48189,N_48164);
and U48308 (N_48308,N_48240,N_48118);
xnor U48309 (N_48309,N_48149,N_48218);
or U48310 (N_48310,N_48026,N_48074);
xnor U48311 (N_48311,N_48057,N_48075);
and U48312 (N_48312,N_48086,N_48012);
xnor U48313 (N_48313,N_48082,N_48165);
nand U48314 (N_48314,N_48184,N_48144);
and U48315 (N_48315,N_48024,N_48199);
xor U48316 (N_48316,N_48077,N_48201);
and U48317 (N_48317,N_48006,N_48200);
or U48318 (N_48318,N_48004,N_48017);
or U48319 (N_48319,N_48031,N_48087);
nand U48320 (N_48320,N_48163,N_48133);
xor U48321 (N_48321,N_48186,N_48098);
or U48322 (N_48322,N_48005,N_48043);
nand U48323 (N_48323,N_48171,N_48235);
xor U48324 (N_48324,N_48097,N_48187);
or U48325 (N_48325,N_48116,N_48155);
and U48326 (N_48326,N_48194,N_48025);
nand U48327 (N_48327,N_48089,N_48054);
nor U48328 (N_48328,N_48027,N_48080);
nand U48329 (N_48329,N_48093,N_48036);
and U48330 (N_48330,N_48142,N_48132);
or U48331 (N_48331,N_48028,N_48062);
and U48332 (N_48332,N_48148,N_48145);
nand U48333 (N_48333,N_48090,N_48063);
nand U48334 (N_48334,N_48202,N_48172);
or U48335 (N_48335,N_48002,N_48168);
or U48336 (N_48336,N_48228,N_48010);
nand U48337 (N_48337,N_48190,N_48180);
nand U48338 (N_48338,N_48175,N_48248);
or U48339 (N_48339,N_48220,N_48152);
xor U48340 (N_48340,N_48014,N_48078);
and U48341 (N_48341,N_48208,N_48035);
or U48342 (N_48342,N_48055,N_48178);
nand U48343 (N_48343,N_48222,N_48016);
nand U48344 (N_48344,N_48019,N_48011);
or U48345 (N_48345,N_48242,N_48066);
xor U48346 (N_48346,N_48051,N_48237);
or U48347 (N_48347,N_48223,N_48185);
or U48348 (N_48348,N_48243,N_48130);
nand U48349 (N_48349,N_48156,N_48070);
and U48350 (N_48350,N_48076,N_48224);
and U48351 (N_48351,N_48176,N_48113);
nor U48352 (N_48352,N_48197,N_48137);
xor U48353 (N_48353,N_48038,N_48138);
or U48354 (N_48354,N_48169,N_48046);
nand U48355 (N_48355,N_48192,N_48245);
xnor U48356 (N_48356,N_48015,N_48127);
nor U48357 (N_48357,N_48151,N_48112);
and U48358 (N_48358,N_48139,N_48083);
xor U48359 (N_48359,N_48146,N_48064);
and U48360 (N_48360,N_48174,N_48158);
xor U48361 (N_48361,N_48088,N_48050);
nor U48362 (N_48362,N_48159,N_48229);
or U48363 (N_48363,N_48179,N_48135);
nor U48364 (N_48364,N_48212,N_48140);
xor U48365 (N_48365,N_48030,N_48094);
xnor U48366 (N_48366,N_48106,N_48052);
nor U48367 (N_48367,N_48102,N_48060);
xnor U48368 (N_48368,N_48114,N_48143);
or U48369 (N_48369,N_48115,N_48100);
and U48370 (N_48370,N_48166,N_48085);
nor U48371 (N_48371,N_48230,N_48239);
and U48372 (N_48372,N_48044,N_48000);
nand U48373 (N_48373,N_48065,N_48068);
xor U48374 (N_48374,N_48213,N_48042);
nand U48375 (N_48375,N_48150,N_48064);
nand U48376 (N_48376,N_48160,N_48221);
nor U48377 (N_48377,N_48100,N_48244);
nor U48378 (N_48378,N_48039,N_48131);
nor U48379 (N_48379,N_48113,N_48249);
nand U48380 (N_48380,N_48073,N_48063);
xor U48381 (N_48381,N_48167,N_48087);
xor U48382 (N_48382,N_48205,N_48136);
nor U48383 (N_48383,N_48001,N_48211);
nor U48384 (N_48384,N_48018,N_48092);
nor U48385 (N_48385,N_48177,N_48028);
and U48386 (N_48386,N_48003,N_48031);
xor U48387 (N_48387,N_48197,N_48033);
or U48388 (N_48388,N_48008,N_48171);
and U48389 (N_48389,N_48206,N_48213);
nand U48390 (N_48390,N_48178,N_48118);
nor U48391 (N_48391,N_48050,N_48221);
or U48392 (N_48392,N_48023,N_48091);
nand U48393 (N_48393,N_48110,N_48233);
or U48394 (N_48394,N_48226,N_48165);
xor U48395 (N_48395,N_48091,N_48173);
or U48396 (N_48396,N_48099,N_48210);
or U48397 (N_48397,N_48163,N_48041);
nor U48398 (N_48398,N_48227,N_48059);
xnor U48399 (N_48399,N_48222,N_48145);
or U48400 (N_48400,N_48165,N_48212);
nand U48401 (N_48401,N_48136,N_48244);
xor U48402 (N_48402,N_48106,N_48157);
and U48403 (N_48403,N_48213,N_48138);
nor U48404 (N_48404,N_48126,N_48199);
and U48405 (N_48405,N_48232,N_48166);
and U48406 (N_48406,N_48071,N_48224);
and U48407 (N_48407,N_48071,N_48020);
nand U48408 (N_48408,N_48162,N_48062);
and U48409 (N_48409,N_48069,N_48063);
and U48410 (N_48410,N_48090,N_48243);
or U48411 (N_48411,N_48194,N_48152);
nand U48412 (N_48412,N_48004,N_48032);
xor U48413 (N_48413,N_48034,N_48156);
or U48414 (N_48414,N_48231,N_48221);
nand U48415 (N_48415,N_48008,N_48179);
xnor U48416 (N_48416,N_48202,N_48080);
or U48417 (N_48417,N_48037,N_48141);
and U48418 (N_48418,N_48149,N_48071);
nand U48419 (N_48419,N_48047,N_48145);
nand U48420 (N_48420,N_48035,N_48229);
or U48421 (N_48421,N_48109,N_48242);
xor U48422 (N_48422,N_48175,N_48161);
nor U48423 (N_48423,N_48090,N_48165);
or U48424 (N_48424,N_48235,N_48187);
or U48425 (N_48425,N_48140,N_48081);
or U48426 (N_48426,N_48119,N_48064);
and U48427 (N_48427,N_48138,N_48026);
xnor U48428 (N_48428,N_48144,N_48065);
nand U48429 (N_48429,N_48234,N_48120);
xor U48430 (N_48430,N_48030,N_48198);
nor U48431 (N_48431,N_48169,N_48153);
and U48432 (N_48432,N_48058,N_48187);
nand U48433 (N_48433,N_48097,N_48152);
nand U48434 (N_48434,N_48049,N_48136);
nand U48435 (N_48435,N_48179,N_48232);
xnor U48436 (N_48436,N_48123,N_48105);
xnor U48437 (N_48437,N_48056,N_48132);
nand U48438 (N_48438,N_48001,N_48120);
nor U48439 (N_48439,N_48241,N_48016);
or U48440 (N_48440,N_48154,N_48042);
nand U48441 (N_48441,N_48150,N_48060);
xnor U48442 (N_48442,N_48129,N_48186);
and U48443 (N_48443,N_48236,N_48042);
xnor U48444 (N_48444,N_48206,N_48212);
or U48445 (N_48445,N_48191,N_48160);
and U48446 (N_48446,N_48084,N_48132);
nand U48447 (N_48447,N_48055,N_48079);
and U48448 (N_48448,N_48237,N_48017);
and U48449 (N_48449,N_48051,N_48190);
or U48450 (N_48450,N_48101,N_48109);
xnor U48451 (N_48451,N_48227,N_48069);
nand U48452 (N_48452,N_48076,N_48236);
or U48453 (N_48453,N_48228,N_48198);
or U48454 (N_48454,N_48086,N_48016);
and U48455 (N_48455,N_48188,N_48120);
nor U48456 (N_48456,N_48100,N_48206);
and U48457 (N_48457,N_48041,N_48222);
nand U48458 (N_48458,N_48195,N_48182);
nand U48459 (N_48459,N_48146,N_48246);
xnor U48460 (N_48460,N_48086,N_48020);
and U48461 (N_48461,N_48072,N_48027);
xnor U48462 (N_48462,N_48047,N_48084);
xor U48463 (N_48463,N_48122,N_48151);
nor U48464 (N_48464,N_48183,N_48239);
nand U48465 (N_48465,N_48040,N_48031);
xor U48466 (N_48466,N_48142,N_48168);
nor U48467 (N_48467,N_48150,N_48124);
xnor U48468 (N_48468,N_48135,N_48111);
nor U48469 (N_48469,N_48181,N_48152);
and U48470 (N_48470,N_48093,N_48030);
nand U48471 (N_48471,N_48216,N_48014);
xor U48472 (N_48472,N_48030,N_48155);
xor U48473 (N_48473,N_48172,N_48230);
nor U48474 (N_48474,N_48242,N_48146);
xnor U48475 (N_48475,N_48178,N_48222);
nand U48476 (N_48476,N_48107,N_48176);
and U48477 (N_48477,N_48094,N_48189);
nand U48478 (N_48478,N_48062,N_48097);
nand U48479 (N_48479,N_48098,N_48012);
or U48480 (N_48480,N_48137,N_48100);
or U48481 (N_48481,N_48235,N_48051);
xor U48482 (N_48482,N_48243,N_48221);
and U48483 (N_48483,N_48171,N_48242);
and U48484 (N_48484,N_48209,N_48034);
nor U48485 (N_48485,N_48145,N_48186);
xnor U48486 (N_48486,N_48137,N_48201);
nand U48487 (N_48487,N_48111,N_48175);
and U48488 (N_48488,N_48095,N_48052);
nor U48489 (N_48489,N_48092,N_48095);
and U48490 (N_48490,N_48220,N_48161);
and U48491 (N_48491,N_48165,N_48005);
xor U48492 (N_48492,N_48125,N_48175);
nand U48493 (N_48493,N_48247,N_48127);
xor U48494 (N_48494,N_48219,N_48040);
nor U48495 (N_48495,N_48151,N_48065);
nand U48496 (N_48496,N_48008,N_48219);
nor U48497 (N_48497,N_48084,N_48107);
or U48498 (N_48498,N_48007,N_48178);
or U48499 (N_48499,N_48094,N_48190);
and U48500 (N_48500,N_48494,N_48274);
nand U48501 (N_48501,N_48465,N_48359);
nand U48502 (N_48502,N_48317,N_48369);
xor U48503 (N_48503,N_48483,N_48295);
xor U48504 (N_48504,N_48496,N_48443);
or U48505 (N_48505,N_48441,N_48415);
nor U48506 (N_48506,N_48458,N_48285);
nand U48507 (N_48507,N_48300,N_48347);
or U48508 (N_48508,N_48325,N_48457);
nand U48509 (N_48509,N_48391,N_48345);
or U48510 (N_48510,N_48375,N_48297);
nand U48511 (N_48511,N_48272,N_48394);
and U48512 (N_48512,N_48407,N_48451);
nor U48513 (N_48513,N_48251,N_48376);
or U48514 (N_48514,N_48477,N_48481);
or U48515 (N_48515,N_48401,N_48257);
xor U48516 (N_48516,N_48308,N_48473);
xnor U48517 (N_48517,N_48396,N_48342);
or U48518 (N_48518,N_48373,N_48314);
or U48519 (N_48519,N_48408,N_48392);
or U48520 (N_48520,N_48493,N_48269);
and U48521 (N_48521,N_48474,N_48307);
nand U48522 (N_48522,N_48312,N_48447);
nand U48523 (N_48523,N_48405,N_48476);
xnor U48524 (N_48524,N_48350,N_48420);
nand U48525 (N_48525,N_48260,N_48414);
nand U48526 (N_48526,N_48337,N_48482);
nand U48527 (N_48527,N_48360,N_48331);
nand U48528 (N_48528,N_48398,N_48271);
and U48529 (N_48529,N_48416,N_48436);
or U48530 (N_48530,N_48366,N_48438);
nand U48531 (N_48531,N_48378,N_48439);
nand U48532 (N_48532,N_48385,N_48426);
nor U48533 (N_48533,N_48397,N_48454);
or U48534 (N_48534,N_48425,N_48365);
nor U48535 (N_48535,N_48291,N_48298);
nor U48536 (N_48536,N_48252,N_48403);
nor U48537 (N_48537,N_48363,N_48364);
or U48538 (N_48538,N_48448,N_48402);
nor U48539 (N_48539,N_48288,N_48404);
nor U48540 (N_48540,N_48282,N_48362);
nand U48541 (N_48541,N_48491,N_48498);
or U48542 (N_48542,N_48351,N_48313);
nor U48543 (N_48543,N_48464,N_48333);
nand U48544 (N_48544,N_48380,N_48480);
xnor U48545 (N_48545,N_48290,N_48283);
nor U48546 (N_48546,N_48265,N_48440);
or U48547 (N_48547,N_48344,N_48395);
or U48548 (N_48548,N_48338,N_48446);
nand U48549 (N_48549,N_48349,N_48497);
and U48550 (N_48550,N_48450,N_48302);
or U48551 (N_48551,N_48423,N_48456);
xnor U48552 (N_48552,N_48460,N_48270);
and U48553 (N_48553,N_48368,N_48422);
xor U48554 (N_48554,N_48452,N_48304);
xor U48555 (N_48555,N_48462,N_48389);
nand U48556 (N_48556,N_48455,N_48284);
xnor U48557 (N_48557,N_48318,N_48387);
or U48558 (N_48558,N_48281,N_48268);
or U48559 (N_48559,N_48437,N_48264);
and U48560 (N_48560,N_48335,N_48419);
or U48561 (N_48561,N_48386,N_48254);
and U48562 (N_48562,N_48445,N_48316);
and U48563 (N_48563,N_48383,N_48323);
nor U48564 (N_48564,N_48390,N_48329);
xnor U48565 (N_48565,N_48348,N_48399);
or U48566 (N_48566,N_48336,N_48276);
xnor U48567 (N_48567,N_48469,N_48301);
xor U48568 (N_48568,N_48352,N_48296);
nand U48569 (N_48569,N_48412,N_48332);
nor U48570 (N_48570,N_48490,N_48478);
nand U48571 (N_48571,N_48287,N_48303);
or U48572 (N_48572,N_48255,N_48495);
or U48573 (N_48573,N_48358,N_48261);
or U48574 (N_48574,N_48311,N_48306);
xnor U48575 (N_48575,N_48411,N_48367);
and U48576 (N_48576,N_48413,N_48353);
nor U48577 (N_48577,N_48292,N_48294);
xnor U48578 (N_48578,N_48467,N_48315);
xor U48579 (N_48579,N_48355,N_48289);
or U48580 (N_48580,N_48424,N_48371);
nor U48581 (N_48581,N_48499,N_48434);
or U48582 (N_48582,N_48322,N_48479);
and U48583 (N_48583,N_48463,N_48339);
xor U48584 (N_48584,N_48453,N_48319);
nand U48585 (N_48585,N_48370,N_48262);
nor U48586 (N_48586,N_48267,N_48418);
xnor U48587 (N_48587,N_48277,N_48340);
nand U48588 (N_48588,N_48273,N_48382);
or U48589 (N_48589,N_48472,N_48361);
and U48590 (N_48590,N_48321,N_48393);
nand U48591 (N_48591,N_48357,N_48466);
nor U48592 (N_48592,N_48410,N_48259);
xnor U48593 (N_48593,N_48280,N_48379);
nor U48594 (N_48594,N_48489,N_48459);
nor U48595 (N_48595,N_48492,N_48305);
nor U48596 (N_48596,N_48330,N_48384);
xor U48597 (N_48597,N_48309,N_48324);
xnor U48598 (N_48598,N_48320,N_48488);
xor U48599 (N_48599,N_48471,N_48409);
nor U48600 (N_48600,N_48343,N_48432);
or U48601 (N_48601,N_48326,N_48356);
nand U48602 (N_48602,N_48279,N_48374);
or U48603 (N_48603,N_48381,N_48470);
and U48604 (N_48604,N_48468,N_48310);
xor U48605 (N_48605,N_48433,N_48263);
nand U48606 (N_48606,N_48372,N_48442);
xnor U48607 (N_48607,N_48354,N_48253);
nor U48608 (N_48608,N_48334,N_48417);
nand U48609 (N_48609,N_48377,N_48435);
or U48610 (N_48610,N_48461,N_48256);
and U48611 (N_48611,N_48299,N_48266);
or U48612 (N_48612,N_48275,N_48449);
xnor U48613 (N_48613,N_48341,N_48388);
nand U48614 (N_48614,N_48346,N_48485);
nor U48615 (N_48615,N_48258,N_48428);
and U48616 (N_48616,N_48431,N_48286);
xor U48617 (N_48617,N_48400,N_48427);
and U48618 (N_48618,N_48430,N_48429);
and U48619 (N_48619,N_48475,N_48406);
xor U48620 (N_48620,N_48484,N_48328);
xnor U48621 (N_48621,N_48486,N_48278);
nand U48622 (N_48622,N_48250,N_48293);
or U48623 (N_48623,N_48421,N_48444);
or U48624 (N_48624,N_48327,N_48487);
or U48625 (N_48625,N_48263,N_48278);
and U48626 (N_48626,N_48359,N_48301);
xnor U48627 (N_48627,N_48263,N_48476);
and U48628 (N_48628,N_48474,N_48266);
or U48629 (N_48629,N_48394,N_48438);
xor U48630 (N_48630,N_48449,N_48314);
and U48631 (N_48631,N_48452,N_48409);
or U48632 (N_48632,N_48455,N_48341);
xor U48633 (N_48633,N_48431,N_48398);
or U48634 (N_48634,N_48344,N_48374);
nand U48635 (N_48635,N_48491,N_48455);
nand U48636 (N_48636,N_48421,N_48382);
and U48637 (N_48637,N_48299,N_48392);
nand U48638 (N_48638,N_48352,N_48461);
or U48639 (N_48639,N_48347,N_48467);
nand U48640 (N_48640,N_48276,N_48398);
and U48641 (N_48641,N_48394,N_48294);
xnor U48642 (N_48642,N_48329,N_48375);
nor U48643 (N_48643,N_48324,N_48494);
and U48644 (N_48644,N_48279,N_48252);
or U48645 (N_48645,N_48358,N_48335);
xor U48646 (N_48646,N_48420,N_48476);
nor U48647 (N_48647,N_48340,N_48331);
nand U48648 (N_48648,N_48348,N_48371);
nor U48649 (N_48649,N_48381,N_48266);
and U48650 (N_48650,N_48437,N_48458);
and U48651 (N_48651,N_48273,N_48453);
xor U48652 (N_48652,N_48469,N_48311);
and U48653 (N_48653,N_48499,N_48259);
xnor U48654 (N_48654,N_48345,N_48362);
or U48655 (N_48655,N_48273,N_48475);
nand U48656 (N_48656,N_48482,N_48423);
and U48657 (N_48657,N_48265,N_48418);
nor U48658 (N_48658,N_48331,N_48396);
and U48659 (N_48659,N_48377,N_48346);
xor U48660 (N_48660,N_48257,N_48486);
nor U48661 (N_48661,N_48261,N_48487);
and U48662 (N_48662,N_48395,N_48324);
or U48663 (N_48663,N_48384,N_48425);
and U48664 (N_48664,N_48255,N_48491);
and U48665 (N_48665,N_48480,N_48343);
nand U48666 (N_48666,N_48385,N_48404);
and U48667 (N_48667,N_48405,N_48455);
xor U48668 (N_48668,N_48478,N_48270);
xor U48669 (N_48669,N_48296,N_48262);
xnor U48670 (N_48670,N_48338,N_48255);
and U48671 (N_48671,N_48403,N_48372);
and U48672 (N_48672,N_48451,N_48261);
and U48673 (N_48673,N_48306,N_48256);
nand U48674 (N_48674,N_48434,N_48257);
and U48675 (N_48675,N_48351,N_48438);
nor U48676 (N_48676,N_48367,N_48382);
and U48677 (N_48677,N_48377,N_48417);
xor U48678 (N_48678,N_48251,N_48333);
xor U48679 (N_48679,N_48328,N_48296);
nor U48680 (N_48680,N_48373,N_48360);
nor U48681 (N_48681,N_48359,N_48326);
nand U48682 (N_48682,N_48358,N_48481);
nor U48683 (N_48683,N_48448,N_48284);
xor U48684 (N_48684,N_48386,N_48477);
nor U48685 (N_48685,N_48288,N_48385);
xor U48686 (N_48686,N_48272,N_48340);
nor U48687 (N_48687,N_48285,N_48306);
nor U48688 (N_48688,N_48485,N_48441);
xor U48689 (N_48689,N_48465,N_48324);
and U48690 (N_48690,N_48292,N_48277);
xor U48691 (N_48691,N_48378,N_48255);
or U48692 (N_48692,N_48480,N_48296);
or U48693 (N_48693,N_48254,N_48452);
or U48694 (N_48694,N_48311,N_48387);
xnor U48695 (N_48695,N_48417,N_48367);
and U48696 (N_48696,N_48278,N_48411);
nand U48697 (N_48697,N_48471,N_48401);
or U48698 (N_48698,N_48354,N_48496);
or U48699 (N_48699,N_48270,N_48321);
xnor U48700 (N_48700,N_48460,N_48429);
nand U48701 (N_48701,N_48396,N_48283);
nor U48702 (N_48702,N_48289,N_48325);
and U48703 (N_48703,N_48443,N_48494);
nor U48704 (N_48704,N_48252,N_48379);
nor U48705 (N_48705,N_48318,N_48472);
nor U48706 (N_48706,N_48298,N_48277);
xor U48707 (N_48707,N_48453,N_48419);
nor U48708 (N_48708,N_48316,N_48288);
and U48709 (N_48709,N_48477,N_48254);
nor U48710 (N_48710,N_48434,N_48255);
or U48711 (N_48711,N_48476,N_48460);
and U48712 (N_48712,N_48321,N_48256);
and U48713 (N_48713,N_48487,N_48270);
or U48714 (N_48714,N_48375,N_48492);
or U48715 (N_48715,N_48345,N_48405);
and U48716 (N_48716,N_48499,N_48446);
nand U48717 (N_48717,N_48396,N_48291);
nor U48718 (N_48718,N_48415,N_48472);
or U48719 (N_48719,N_48290,N_48307);
or U48720 (N_48720,N_48306,N_48291);
and U48721 (N_48721,N_48354,N_48256);
xnor U48722 (N_48722,N_48370,N_48283);
and U48723 (N_48723,N_48286,N_48455);
nor U48724 (N_48724,N_48346,N_48392);
and U48725 (N_48725,N_48326,N_48393);
xnor U48726 (N_48726,N_48323,N_48356);
or U48727 (N_48727,N_48482,N_48463);
nor U48728 (N_48728,N_48378,N_48254);
nand U48729 (N_48729,N_48464,N_48306);
xnor U48730 (N_48730,N_48252,N_48499);
xor U48731 (N_48731,N_48435,N_48279);
and U48732 (N_48732,N_48483,N_48255);
nand U48733 (N_48733,N_48313,N_48462);
nand U48734 (N_48734,N_48300,N_48433);
or U48735 (N_48735,N_48441,N_48289);
xnor U48736 (N_48736,N_48258,N_48429);
nand U48737 (N_48737,N_48478,N_48402);
nor U48738 (N_48738,N_48412,N_48478);
xor U48739 (N_48739,N_48271,N_48418);
nor U48740 (N_48740,N_48375,N_48252);
and U48741 (N_48741,N_48498,N_48309);
or U48742 (N_48742,N_48367,N_48341);
nor U48743 (N_48743,N_48355,N_48419);
or U48744 (N_48744,N_48372,N_48371);
or U48745 (N_48745,N_48476,N_48497);
or U48746 (N_48746,N_48478,N_48331);
nand U48747 (N_48747,N_48495,N_48364);
xor U48748 (N_48748,N_48253,N_48280);
nand U48749 (N_48749,N_48426,N_48271);
nor U48750 (N_48750,N_48664,N_48597);
nor U48751 (N_48751,N_48513,N_48579);
nand U48752 (N_48752,N_48660,N_48507);
or U48753 (N_48753,N_48606,N_48748);
nand U48754 (N_48754,N_48652,N_48742);
xnor U48755 (N_48755,N_48633,N_48612);
and U48756 (N_48756,N_48725,N_48509);
and U48757 (N_48757,N_48678,N_48666);
xor U48758 (N_48758,N_48663,N_48711);
or U48759 (N_48759,N_48685,N_48578);
nand U48760 (N_48760,N_48592,N_48686);
xnor U48761 (N_48761,N_48604,N_48532);
xor U48762 (N_48762,N_48676,N_48733);
nand U48763 (N_48763,N_48671,N_48672);
xor U48764 (N_48764,N_48608,N_48627);
or U48765 (N_48765,N_48646,N_48587);
nand U48766 (N_48766,N_48525,N_48719);
and U48767 (N_48767,N_48591,N_48538);
xnor U48768 (N_48768,N_48503,N_48500);
and U48769 (N_48769,N_48512,N_48514);
and U48770 (N_48770,N_48595,N_48736);
nor U48771 (N_48771,N_48528,N_48710);
or U48772 (N_48772,N_48524,N_48644);
nor U48773 (N_48773,N_48623,N_48529);
nor U48774 (N_48774,N_48674,N_48728);
nor U48775 (N_48775,N_48629,N_48694);
or U48776 (N_48776,N_48647,N_48642);
nor U48777 (N_48777,N_48508,N_48635);
nor U48778 (N_48778,N_48583,N_48703);
nor U48779 (N_48779,N_48562,N_48723);
or U48780 (N_48780,N_48568,N_48746);
xnor U48781 (N_48781,N_48540,N_48731);
nor U48782 (N_48782,N_48721,N_48610);
nand U48783 (N_48783,N_48621,N_48543);
nor U48784 (N_48784,N_48636,N_48639);
nor U48785 (N_48785,N_48716,N_48522);
and U48786 (N_48786,N_48670,N_48744);
or U48787 (N_48787,N_48563,N_48519);
or U48788 (N_48788,N_48580,N_48501);
and U48789 (N_48789,N_48677,N_48707);
nor U48790 (N_48790,N_48545,N_48649);
xor U48791 (N_48791,N_48617,N_48510);
nand U48792 (N_48792,N_48593,N_48502);
nand U48793 (N_48793,N_48523,N_48586);
or U48794 (N_48794,N_48506,N_48609);
and U48795 (N_48795,N_48556,N_48620);
nor U48796 (N_48796,N_48605,N_48565);
nand U48797 (N_48797,N_48738,N_48706);
xnor U48798 (N_48798,N_48526,N_48521);
or U48799 (N_48799,N_48640,N_48741);
xnor U48800 (N_48800,N_48722,N_48541);
xor U48801 (N_48801,N_48717,N_48714);
or U48802 (N_48802,N_48618,N_48504);
nand U48803 (N_48803,N_48691,N_48675);
and U48804 (N_48804,N_48570,N_48684);
nand U48805 (N_48805,N_48724,N_48622);
nand U48806 (N_48806,N_48625,N_48534);
xor U48807 (N_48807,N_48705,N_48704);
nand U48808 (N_48808,N_48602,N_48628);
or U48809 (N_48809,N_48700,N_48564);
and U48810 (N_48810,N_48661,N_48645);
xnor U48811 (N_48811,N_48600,N_48544);
and U48812 (N_48812,N_48619,N_48702);
nand U48813 (N_48813,N_48690,N_48582);
nand U48814 (N_48814,N_48547,N_48734);
and U48815 (N_48815,N_48624,N_48553);
nand U48816 (N_48816,N_48740,N_48511);
or U48817 (N_48817,N_48658,N_48551);
nor U48818 (N_48818,N_48546,N_48552);
or U48819 (N_48819,N_48662,N_48516);
nand U48820 (N_48820,N_48683,N_48571);
xor U48821 (N_48821,N_48550,N_48613);
xor U48822 (N_48822,N_48577,N_48693);
and U48823 (N_48823,N_48695,N_48650);
nand U48824 (N_48824,N_48667,N_48549);
xor U48825 (N_48825,N_48708,N_48615);
nand U48826 (N_48826,N_48648,N_48626);
nand U48827 (N_48827,N_48729,N_48634);
and U48828 (N_48828,N_48669,N_48699);
or U48829 (N_48829,N_48697,N_48701);
or U48830 (N_48830,N_48656,N_48745);
and U48831 (N_48831,N_48726,N_48637);
and U48832 (N_48832,N_48611,N_48680);
and U48833 (N_48833,N_48631,N_48659);
nand U48834 (N_48834,N_48668,N_48588);
xor U48835 (N_48835,N_48689,N_48590);
and U48836 (N_48836,N_48589,N_48585);
or U48837 (N_48837,N_48696,N_48687);
nand U48838 (N_48838,N_48692,N_48632);
or U48839 (N_48839,N_48520,N_48630);
and U48840 (N_48840,N_48530,N_48720);
or U48841 (N_48841,N_48575,N_48581);
nor U48842 (N_48842,N_48688,N_48735);
xnor U48843 (N_48843,N_48555,N_48584);
nor U48844 (N_48844,N_48657,N_48572);
or U48845 (N_48845,N_48535,N_48557);
and U48846 (N_48846,N_48569,N_48709);
xnor U48847 (N_48847,N_48749,N_48505);
and U48848 (N_48848,N_48517,N_48601);
nand U48849 (N_48849,N_48641,N_48643);
nand U48850 (N_48850,N_48537,N_48638);
xor U48851 (N_48851,N_48682,N_48713);
xor U48852 (N_48852,N_48743,N_48559);
or U48853 (N_48853,N_48739,N_48727);
nor U48854 (N_48854,N_48558,N_48566);
xnor U48855 (N_48855,N_48596,N_48536);
or U48856 (N_48856,N_48576,N_48653);
or U48857 (N_48857,N_48598,N_48747);
nand U48858 (N_48858,N_48616,N_48718);
nor U48859 (N_48859,N_48567,N_48654);
nand U48860 (N_48860,N_48548,N_48603);
xor U48861 (N_48861,N_48539,N_48651);
and U48862 (N_48862,N_48574,N_48531);
xnor U48863 (N_48863,N_48607,N_48730);
and U48864 (N_48864,N_48679,N_48737);
or U48865 (N_48865,N_48542,N_48712);
xor U48866 (N_48866,N_48594,N_48673);
nor U48867 (N_48867,N_48732,N_48518);
or U48868 (N_48868,N_48560,N_48681);
xnor U48869 (N_48869,N_48715,N_48533);
or U48870 (N_48870,N_48599,N_48554);
or U48871 (N_48871,N_48665,N_48573);
or U48872 (N_48872,N_48698,N_48561);
nor U48873 (N_48873,N_48614,N_48515);
nand U48874 (N_48874,N_48655,N_48527);
or U48875 (N_48875,N_48590,N_48746);
nand U48876 (N_48876,N_48683,N_48660);
or U48877 (N_48877,N_48524,N_48578);
or U48878 (N_48878,N_48609,N_48692);
nor U48879 (N_48879,N_48593,N_48667);
nand U48880 (N_48880,N_48653,N_48633);
and U48881 (N_48881,N_48559,N_48515);
nor U48882 (N_48882,N_48566,N_48518);
and U48883 (N_48883,N_48675,N_48717);
and U48884 (N_48884,N_48709,N_48714);
or U48885 (N_48885,N_48722,N_48669);
and U48886 (N_48886,N_48611,N_48647);
and U48887 (N_48887,N_48738,N_48657);
or U48888 (N_48888,N_48701,N_48528);
xnor U48889 (N_48889,N_48641,N_48728);
xnor U48890 (N_48890,N_48654,N_48557);
or U48891 (N_48891,N_48573,N_48617);
xor U48892 (N_48892,N_48596,N_48610);
nor U48893 (N_48893,N_48663,N_48554);
xnor U48894 (N_48894,N_48580,N_48547);
or U48895 (N_48895,N_48523,N_48688);
and U48896 (N_48896,N_48621,N_48514);
nand U48897 (N_48897,N_48512,N_48549);
nor U48898 (N_48898,N_48615,N_48582);
and U48899 (N_48899,N_48582,N_48530);
nor U48900 (N_48900,N_48618,N_48511);
or U48901 (N_48901,N_48603,N_48723);
nand U48902 (N_48902,N_48531,N_48658);
and U48903 (N_48903,N_48525,N_48606);
or U48904 (N_48904,N_48714,N_48625);
nand U48905 (N_48905,N_48657,N_48723);
and U48906 (N_48906,N_48697,N_48724);
or U48907 (N_48907,N_48624,N_48548);
xor U48908 (N_48908,N_48731,N_48647);
nor U48909 (N_48909,N_48547,N_48729);
and U48910 (N_48910,N_48560,N_48600);
xnor U48911 (N_48911,N_48648,N_48519);
nor U48912 (N_48912,N_48703,N_48532);
nand U48913 (N_48913,N_48584,N_48626);
xor U48914 (N_48914,N_48681,N_48593);
nor U48915 (N_48915,N_48691,N_48657);
nand U48916 (N_48916,N_48614,N_48640);
and U48917 (N_48917,N_48731,N_48553);
xor U48918 (N_48918,N_48748,N_48734);
nand U48919 (N_48919,N_48529,N_48504);
xor U48920 (N_48920,N_48531,N_48654);
xnor U48921 (N_48921,N_48742,N_48704);
or U48922 (N_48922,N_48720,N_48723);
xnor U48923 (N_48923,N_48518,N_48547);
xnor U48924 (N_48924,N_48699,N_48609);
or U48925 (N_48925,N_48730,N_48676);
nor U48926 (N_48926,N_48638,N_48738);
xor U48927 (N_48927,N_48581,N_48542);
xnor U48928 (N_48928,N_48674,N_48530);
xnor U48929 (N_48929,N_48697,N_48710);
xor U48930 (N_48930,N_48695,N_48687);
xnor U48931 (N_48931,N_48580,N_48579);
and U48932 (N_48932,N_48689,N_48503);
nor U48933 (N_48933,N_48603,N_48690);
xnor U48934 (N_48934,N_48597,N_48552);
nor U48935 (N_48935,N_48596,N_48589);
and U48936 (N_48936,N_48577,N_48616);
nand U48937 (N_48937,N_48514,N_48672);
nor U48938 (N_48938,N_48571,N_48720);
xor U48939 (N_48939,N_48705,N_48659);
and U48940 (N_48940,N_48692,N_48671);
or U48941 (N_48941,N_48746,N_48565);
nor U48942 (N_48942,N_48661,N_48515);
xor U48943 (N_48943,N_48674,N_48631);
or U48944 (N_48944,N_48644,N_48625);
and U48945 (N_48945,N_48645,N_48650);
and U48946 (N_48946,N_48594,N_48644);
or U48947 (N_48947,N_48721,N_48647);
xnor U48948 (N_48948,N_48693,N_48672);
nand U48949 (N_48949,N_48557,N_48634);
xnor U48950 (N_48950,N_48617,N_48511);
and U48951 (N_48951,N_48696,N_48698);
or U48952 (N_48952,N_48542,N_48687);
xor U48953 (N_48953,N_48705,N_48565);
and U48954 (N_48954,N_48686,N_48724);
nand U48955 (N_48955,N_48516,N_48550);
and U48956 (N_48956,N_48586,N_48583);
or U48957 (N_48957,N_48636,N_48679);
or U48958 (N_48958,N_48723,N_48505);
nor U48959 (N_48959,N_48674,N_48696);
xnor U48960 (N_48960,N_48576,N_48665);
xor U48961 (N_48961,N_48713,N_48689);
nor U48962 (N_48962,N_48529,N_48727);
and U48963 (N_48963,N_48570,N_48614);
and U48964 (N_48964,N_48602,N_48672);
nand U48965 (N_48965,N_48710,N_48726);
xnor U48966 (N_48966,N_48616,N_48633);
and U48967 (N_48967,N_48633,N_48555);
xor U48968 (N_48968,N_48635,N_48708);
or U48969 (N_48969,N_48719,N_48662);
and U48970 (N_48970,N_48609,N_48611);
nor U48971 (N_48971,N_48574,N_48528);
and U48972 (N_48972,N_48642,N_48515);
nor U48973 (N_48973,N_48544,N_48562);
nor U48974 (N_48974,N_48694,N_48731);
nand U48975 (N_48975,N_48606,N_48716);
and U48976 (N_48976,N_48711,N_48547);
xnor U48977 (N_48977,N_48718,N_48500);
nor U48978 (N_48978,N_48634,N_48593);
xnor U48979 (N_48979,N_48602,N_48627);
or U48980 (N_48980,N_48559,N_48685);
or U48981 (N_48981,N_48738,N_48533);
xor U48982 (N_48982,N_48695,N_48742);
nand U48983 (N_48983,N_48653,N_48694);
or U48984 (N_48984,N_48741,N_48727);
and U48985 (N_48985,N_48664,N_48583);
or U48986 (N_48986,N_48533,N_48670);
or U48987 (N_48987,N_48633,N_48512);
and U48988 (N_48988,N_48508,N_48540);
or U48989 (N_48989,N_48540,N_48680);
or U48990 (N_48990,N_48694,N_48633);
nor U48991 (N_48991,N_48696,N_48742);
and U48992 (N_48992,N_48703,N_48709);
and U48993 (N_48993,N_48583,N_48612);
or U48994 (N_48994,N_48560,N_48574);
nor U48995 (N_48995,N_48695,N_48704);
xnor U48996 (N_48996,N_48655,N_48593);
nor U48997 (N_48997,N_48572,N_48733);
xor U48998 (N_48998,N_48639,N_48587);
nand U48999 (N_48999,N_48539,N_48663);
or U49000 (N_49000,N_48796,N_48889);
and U49001 (N_49001,N_48888,N_48978);
and U49002 (N_49002,N_48852,N_48854);
xnor U49003 (N_49003,N_48877,N_48938);
nor U49004 (N_49004,N_48947,N_48935);
and U49005 (N_49005,N_48945,N_48855);
xnor U49006 (N_49006,N_48863,N_48974);
nand U49007 (N_49007,N_48962,N_48750);
xor U49008 (N_49008,N_48794,N_48925);
and U49009 (N_49009,N_48799,N_48891);
nor U49010 (N_49010,N_48783,N_48982);
nand U49011 (N_49011,N_48956,N_48987);
xor U49012 (N_49012,N_48981,N_48814);
nor U49013 (N_49013,N_48934,N_48932);
or U49014 (N_49014,N_48904,N_48804);
xnor U49015 (N_49015,N_48807,N_48884);
and U49016 (N_49016,N_48805,N_48984);
nand U49017 (N_49017,N_48753,N_48998);
and U49018 (N_49018,N_48903,N_48908);
nand U49019 (N_49019,N_48853,N_48819);
or U49020 (N_49020,N_48955,N_48882);
nor U49021 (N_49021,N_48772,N_48911);
and U49022 (N_49022,N_48788,N_48972);
or U49023 (N_49023,N_48951,N_48913);
nand U49024 (N_49024,N_48936,N_48810);
and U49025 (N_49025,N_48970,N_48781);
and U49026 (N_49026,N_48880,N_48848);
xnor U49027 (N_49027,N_48886,N_48774);
nor U49028 (N_49028,N_48791,N_48988);
or U49029 (N_49029,N_48968,N_48948);
nand U49030 (N_49030,N_48875,N_48887);
or U49031 (N_49031,N_48818,N_48760);
or U49032 (N_49032,N_48761,N_48907);
nand U49033 (N_49033,N_48975,N_48926);
and U49034 (N_49034,N_48865,N_48801);
and U49035 (N_49035,N_48993,N_48942);
or U49036 (N_49036,N_48780,N_48901);
or U49037 (N_49037,N_48830,N_48851);
xor U49038 (N_49038,N_48892,N_48828);
nand U49039 (N_49039,N_48792,N_48953);
nand U49040 (N_49040,N_48829,N_48977);
or U49041 (N_49041,N_48834,N_48841);
or U49042 (N_49042,N_48806,N_48831);
nor U49043 (N_49043,N_48812,N_48835);
xor U49044 (N_49044,N_48895,N_48837);
and U49045 (N_49045,N_48905,N_48967);
xor U49046 (N_49046,N_48966,N_48943);
nand U49047 (N_49047,N_48960,N_48906);
or U49048 (N_49048,N_48986,N_48756);
nor U49049 (N_49049,N_48857,N_48881);
nand U49050 (N_49050,N_48929,N_48838);
nand U49051 (N_49051,N_48850,N_48847);
nand U49052 (N_49052,N_48826,N_48817);
nand U49053 (N_49053,N_48918,N_48859);
or U49054 (N_49054,N_48840,N_48973);
or U49055 (N_49055,N_48846,N_48985);
xnor U49056 (N_49056,N_48861,N_48959);
nor U49057 (N_49057,N_48897,N_48964);
nand U49058 (N_49058,N_48969,N_48786);
xnor U49059 (N_49059,N_48765,N_48770);
xnor U49060 (N_49060,N_48946,N_48940);
or U49061 (N_49061,N_48950,N_48784);
and U49062 (N_49062,N_48954,N_48894);
nand U49063 (N_49063,N_48979,N_48755);
and U49064 (N_49064,N_48787,N_48839);
nand U49065 (N_49065,N_48776,N_48927);
and U49066 (N_49066,N_48937,N_48758);
xor U49067 (N_49067,N_48797,N_48757);
nand U49068 (N_49068,N_48991,N_48754);
nor U49069 (N_49069,N_48873,N_48782);
and U49070 (N_49070,N_48871,N_48976);
or U49071 (N_49071,N_48914,N_48775);
nor U49072 (N_49072,N_48763,N_48823);
xor U49073 (N_49073,N_48767,N_48922);
xor U49074 (N_49074,N_48921,N_48836);
xnor U49075 (N_49075,N_48872,N_48971);
nand U49076 (N_49076,N_48762,N_48996);
or U49077 (N_49077,N_48923,N_48919);
nand U49078 (N_49078,N_48764,N_48856);
and U49079 (N_49079,N_48866,N_48999);
nor U49080 (N_49080,N_48957,N_48825);
or U49081 (N_49081,N_48909,N_48990);
or U49082 (N_49082,N_48883,N_48924);
and U49083 (N_49083,N_48902,N_48885);
nor U49084 (N_49084,N_48751,N_48773);
xnor U49085 (N_49085,N_48821,N_48789);
nor U49086 (N_49086,N_48952,N_48832);
xor U49087 (N_49087,N_48790,N_48980);
nor U49088 (N_49088,N_48898,N_48778);
nand U49089 (N_49089,N_48768,N_48766);
nor U49090 (N_49090,N_48879,N_48900);
or U49091 (N_49091,N_48822,N_48933);
or U49092 (N_49092,N_48916,N_48949);
nand U49093 (N_49093,N_48800,N_48798);
xnor U49094 (N_49094,N_48878,N_48824);
or U49095 (N_49095,N_48845,N_48869);
or U49096 (N_49096,N_48896,N_48862);
or U49097 (N_49097,N_48793,N_48820);
or U49098 (N_49098,N_48803,N_48868);
nand U49099 (N_49099,N_48870,N_48983);
xnor U49100 (N_49100,N_48997,N_48802);
or U49101 (N_49101,N_48842,N_48963);
nand U49102 (N_49102,N_48910,N_48769);
and U49103 (N_49103,N_48771,N_48915);
and U49104 (N_49104,N_48874,N_48912);
or U49105 (N_49105,N_48994,N_48899);
nor U49106 (N_49106,N_48941,N_48867);
nor U49107 (N_49107,N_48864,N_48928);
or U49108 (N_49108,N_48920,N_48759);
or U49109 (N_49109,N_48860,N_48795);
and U49110 (N_49110,N_48958,N_48811);
and U49111 (N_49111,N_48989,N_48849);
nor U49112 (N_49112,N_48777,N_48992);
xor U49113 (N_49113,N_48815,N_48833);
nor U49114 (N_49114,N_48965,N_48939);
nor U49115 (N_49115,N_48995,N_48785);
or U49116 (N_49116,N_48890,N_48779);
nand U49117 (N_49117,N_48931,N_48858);
nand U49118 (N_49118,N_48752,N_48808);
or U49119 (N_49119,N_48917,N_48844);
xnor U49120 (N_49120,N_48816,N_48944);
and U49121 (N_49121,N_48876,N_48813);
and U49122 (N_49122,N_48827,N_48893);
nand U49123 (N_49123,N_48809,N_48961);
nor U49124 (N_49124,N_48930,N_48843);
nand U49125 (N_49125,N_48789,N_48949);
nand U49126 (N_49126,N_48851,N_48991);
or U49127 (N_49127,N_48912,N_48997);
nor U49128 (N_49128,N_48970,N_48892);
and U49129 (N_49129,N_48873,N_48885);
nand U49130 (N_49130,N_48773,N_48869);
or U49131 (N_49131,N_48917,N_48979);
xnor U49132 (N_49132,N_48833,N_48862);
nand U49133 (N_49133,N_48908,N_48917);
xor U49134 (N_49134,N_48976,N_48805);
xor U49135 (N_49135,N_48811,N_48995);
and U49136 (N_49136,N_48903,N_48855);
nor U49137 (N_49137,N_48844,N_48981);
nand U49138 (N_49138,N_48838,N_48776);
xor U49139 (N_49139,N_48971,N_48914);
and U49140 (N_49140,N_48778,N_48981);
nand U49141 (N_49141,N_48951,N_48826);
nand U49142 (N_49142,N_48934,N_48870);
xor U49143 (N_49143,N_48765,N_48982);
nand U49144 (N_49144,N_48853,N_48995);
nand U49145 (N_49145,N_48975,N_48993);
nand U49146 (N_49146,N_48819,N_48956);
and U49147 (N_49147,N_48832,N_48838);
xor U49148 (N_49148,N_48870,N_48754);
nand U49149 (N_49149,N_48848,N_48782);
nor U49150 (N_49150,N_48751,N_48855);
and U49151 (N_49151,N_48842,N_48871);
nor U49152 (N_49152,N_48812,N_48801);
xnor U49153 (N_49153,N_48979,N_48805);
and U49154 (N_49154,N_48883,N_48988);
xor U49155 (N_49155,N_48874,N_48891);
nand U49156 (N_49156,N_48925,N_48775);
nor U49157 (N_49157,N_48981,N_48802);
nor U49158 (N_49158,N_48954,N_48843);
xnor U49159 (N_49159,N_48836,N_48963);
and U49160 (N_49160,N_48922,N_48843);
nand U49161 (N_49161,N_48781,N_48907);
xnor U49162 (N_49162,N_48892,N_48818);
and U49163 (N_49163,N_48753,N_48929);
or U49164 (N_49164,N_48857,N_48783);
xnor U49165 (N_49165,N_48884,N_48813);
and U49166 (N_49166,N_48903,N_48971);
nand U49167 (N_49167,N_48904,N_48823);
nand U49168 (N_49168,N_48757,N_48939);
nand U49169 (N_49169,N_48753,N_48905);
nor U49170 (N_49170,N_48935,N_48940);
nor U49171 (N_49171,N_48932,N_48900);
and U49172 (N_49172,N_48960,N_48778);
nand U49173 (N_49173,N_48904,N_48854);
nor U49174 (N_49174,N_48782,N_48964);
and U49175 (N_49175,N_48980,N_48829);
nand U49176 (N_49176,N_48906,N_48920);
xnor U49177 (N_49177,N_48974,N_48963);
or U49178 (N_49178,N_48851,N_48884);
nand U49179 (N_49179,N_48969,N_48826);
or U49180 (N_49180,N_48878,N_48875);
and U49181 (N_49181,N_48836,N_48896);
or U49182 (N_49182,N_48825,N_48762);
nor U49183 (N_49183,N_48812,N_48870);
or U49184 (N_49184,N_48847,N_48853);
nand U49185 (N_49185,N_48852,N_48914);
nor U49186 (N_49186,N_48944,N_48900);
or U49187 (N_49187,N_48817,N_48887);
xnor U49188 (N_49188,N_48848,N_48938);
and U49189 (N_49189,N_48884,N_48763);
nand U49190 (N_49190,N_48771,N_48833);
xor U49191 (N_49191,N_48901,N_48847);
or U49192 (N_49192,N_48983,N_48833);
nand U49193 (N_49193,N_48887,N_48879);
nor U49194 (N_49194,N_48926,N_48928);
nor U49195 (N_49195,N_48789,N_48903);
or U49196 (N_49196,N_48969,N_48825);
nand U49197 (N_49197,N_48806,N_48779);
xor U49198 (N_49198,N_48962,N_48836);
nand U49199 (N_49199,N_48846,N_48841);
and U49200 (N_49200,N_48780,N_48789);
nor U49201 (N_49201,N_48968,N_48964);
and U49202 (N_49202,N_48853,N_48803);
nor U49203 (N_49203,N_48801,N_48936);
xor U49204 (N_49204,N_48865,N_48823);
nor U49205 (N_49205,N_48878,N_48961);
nor U49206 (N_49206,N_48971,N_48885);
nor U49207 (N_49207,N_48778,N_48823);
nand U49208 (N_49208,N_48939,N_48934);
xor U49209 (N_49209,N_48829,N_48967);
or U49210 (N_49210,N_48784,N_48791);
nand U49211 (N_49211,N_48874,N_48776);
or U49212 (N_49212,N_48842,N_48989);
xor U49213 (N_49213,N_48919,N_48825);
nor U49214 (N_49214,N_48933,N_48873);
or U49215 (N_49215,N_48823,N_48815);
nor U49216 (N_49216,N_48953,N_48982);
nor U49217 (N_49217,N_48927,N_48891);
nand U49218 (N_49218,N_48790,N_48822);
nand U49219 (N_49219,N_48975,N_48957);
nand U49220 (N_49220,N_48874,N_48959);
nand U49221 (N_49221,N_48948,N_48751);
or U49222 (N_49222,N_48966,N_48970);
xnor U49223 (N_49223,N_48778,N_48943);
and U49224 (N_49224,N_48759,N_48778);
and U49225 (N_49225,N_48811,N_48970);
nor U49226 (N_49226,N_48984,N_48759);
or U49227 (N_49227,N_48943,N_48772);
and U49228 (N_49228,N_48759,N_48981);
and U49229 (N_49229,N_48982,N_48850);
or U49230 (N_49230,N_48791,N_48978);
nand U49231 (N_49231,N_48983,N_48801);
and U49232 (N_49232,N_48782,N_48972);
xor U49233 (N_49233,N_48933,N_48953);
xnor U49234 (N_49234,N_48907,N_48941);
xnor U49235 (N_49235,N_48986,N_48882);
nand U49236 (N_49236,N_48996,N_48960);
or U49237 (N_49237,N_48993,N_48785);
and U49238 (N_49238,N_48806,N_48795);
nand U49239 (N_49239,N_48879,N_48877);
nand U49240 (N_49240,N_48763,N_48963);
and U49241 (N_49241,N_48985,N_48822);
nor U49242 (N_49242,N_48925,N_48813);
and U49243 (N_49243,N_48910,N_48899);
or U49244 (N_49244,N_48869,N_48873);
and U49245 (N_49245,N_48942,N_48854);
nor U49246 (N_49246,N_48960,N_48939);
nand U49247 (N_49247,N_48766,N_48951);
or U49248 (N_49248,N_48971,N_48944);
xor U49249 (N_49249,N_48951,N_48832);
nor U49250 (N_49250,N_49061,N_49238);
xor U49251 (N_49251,N_49080,N_49024);
or U49252 (N_49252,N_49130,N_49164);
nor U49253 (N_49253,N_49030,N_49202);
and U49254 (N_49254,N_49100,N_49028);
nand U49255 (N_49255,N_49219,N_49146);
nor U49256 (N_49256,N_49009,N_49233);
nand U49257 (N_49257,N_49026,N_49208);
and U49258 (N_49258,N_49195,N_49232);
nor U49259 (N_49259,N_49122,N_49016);
and U49260 (N_49260,N_49018,N_49211);
xnor U49261 (N_49261,N_49156,N_49025);
nor U49262 (N_49262,N_49085,N_49147);
or U49263 (N_49263,N_49227,N_49082);
and U49264 (N_49264,N_49029,N_49043);
nor U49265 (N_49265,N_49126,N_49128);
nand U49266 (N_49266,N_49201,N_49078);
nand U49267 (N_49267,N_49022,N_49042);
and U49268 (N_49268,N_49239,N_49039);
xnor U49269 (N_49269,N_49160,N_49065);
nor U49270 (N_49270,N_49194,N_49235);
and U49271 (N_49271,N_49151,N_49037);
and U49272 (N_49272,N_49124,N_49175);
nand U49273 (N_49273,N_49129,N_49079);
xor U49274 (N_49274,N_49209,N_49084);
nor U49275 (N_49275,N_49047,N_49172);
or U49276 (N_49276,N_49125,N_49188);
xor U49277 (N_49277,N_49155,N_49000);
or U49278 (N_49278,N_49107,N_49032);
xnor U49279 (N_49279,N_49117,N_49200);
nand U49280 (N_49280,N_49051,N_49105);
xor U49281 (N_49281,N_49135,N_49249);
and U49282 (N_49282,N_49119,N_49215);
and U49283 (N_49283,N_49169,N_49138);
and U49284 (N_49284,N_49098,N_49236);
and U49285 (N_49285,N_49132,N_49040);
xor U49286 (N_49286,N_49052,N_49162);
or U49287 (N_49287,N_49001,N_49190);
or U49288 (N_49288,N_49068,N_49027);
or U49289 (N_49289,N_49224,N_49178);
or U49290 (N_49290,N_49181,N_49210);
and U49291 (N_49291,N_49187,N_49139);
and U49292 (N_49292,N_49007,N_49110);
xor U49293 (N_49293,N_49091,N_49087);
or U49294 (N_49294,N_49168,N_49141);
nor U49295 (N_49295,N_49222,N_49218);
and U49296 (N_49296,N_49193,N_49205);
and U49297 (N_49297,N_49152,N_49101);
nor U49298 (N_49298,N_49161,N_49011);
or U49299 (N_49299,N_49242,N_49230);
nor U49300 (N_49300,N_49140,N_49183);
xor U49301 (N_49301,N_49213,N_49012);
nor U49302 (N_49302,N_49176,N_49246);
nand U49303 (N_49303,N_49153,N_49165);
xor U49304 (N_49304,N_49111,N_49173);
and U49305 (N_49305,N_49217,N_49099);
xnor U49306 (N_49306,N_49064,N_49220);
and U49307 (N_49307,N_49020,N_49229);
and U49308 (N_49308,N_49106,N_49159);
nor U49309 (N_49309,N_49184,N_49131);
or U49310 (N_49310,N_49189,N_49203);
or U49311 (N_49311,N_49243,N_49148);
xor U49312 (N_49312,N_49017,N_49121);
or U49313 (N_49313,N_49060,N_49036);
and U49314 (N_49314,N_49077,N_49045);
or U49315 (N_49315,N_49102,N_49248);
nor U49316 (N_49316,N_49163,N_49134);
or U49317 (N_49317,N_49096,N_49145);
and U49318 (N_49318,N_49247,N_49180);
nor U49319 (N_49319,N_49245,N_49035);
nand U49320 (N_49320,N_49171,N_49179);
nand U49321 (N_49321,N_49204,N_49056);
nor U49322 (N_49322,N_49109,N_49231);
or U49323 (N_49323,N_49240,N_49090);
and U49324 (N_49324,N_49019,N_49041);
nor U49325 (N_49325,N_49226,N_49113);
and U49326 (N_49326,N_49021,N_49166);
nand U49327 (N_49327,N_49023,N_49136);
and U49328 (N_49328,N_49144,N_49075);
and U49329 (N_49329,N_49057,N_49088);
nor U49330 (N_49330,N_49066,N_49014);
nand U49331 (N_49331,N_49225,N_49103);
or U49332 (N_49332,N_49033,N_49055);
xor U49333 (N_49333,N_49133,N_49071);
nand U49334 (N_49334,N_49069,N_49063);
nor U49335 (N_49335,N_49223,N_49089);
xnor U49336 (N_49336,N_49093,N_49054);
xor U49337 (N_49337,N_49237,N_49207);
nand U49338 (N_49338,N_49120,N_49182);
or U49339 (N_49339,N_49157,N_49008);
nand U49340 (N_49340,N_49038,N_49199);
nand U49341 (N_49341,N_49074,N_49058);
or U49342 (N_49342,N_49228,N_49196);
xor U49343 (N_49343,N_49059,N_49095);
or U49344 (N_49344,N_49150,N_49062);
and U49345 (N_49345,N_49216,N_49115);
or U49346 (N_49346,N_49073,N_49143);
or U49347 (N_49347,N_49244,N_49170);
or U49348 (N_49348,N_49154,N_49198);
nor U49349 (N_49349,N_49212,N_49006);
nand U49350 (N_49350,N_49005,N_49081);
and U49351 (N_49351,N_49049,N_49108);
nor U49352 (N_49352,N_49142,N_49083);
or U49353 (N_49353,N_49097,N_49053);
nand U49354 (N_49354,N_49137,N_49092);
nor U49355 (N_49355,N_49048,N_49076);
nor U49356 (N_49356,N_49034,N_49191);
xnor U49357 (N_49357,N_49185,N_49174);
nor U49358 (N_49358,N_49072,N_49031);
nor U49359 (N_49359,N_49197,N_49116);
nand U49360 (N_49360,N_49167,N_49241);
nand U49361 (N_49361,N_49112,N_49046);
and U49362 (N_49362,N_49067,N_49004);
or U49363 (N_49363,N_49186,N_49118);
or U49364 (N_49364,N_49123,N_49044);
nor U49365 (N_49365,N_49002,N_49015);
xor U49366 (N_49366,N_49192,N_49010);
and U49367 (N_49367,N_49221,N_49114);
nor U49368 (N_49368,N_49086,N_49094);
and U49369 (N_49369,N_49149,N_49013);
and U49370 (N_49370,N_49127,N_49070);
nand U49371 (N_49371,N_49177,N_49206);
or U49372 (N_49372,N_49214,N_49104);
or U49373 (N_49373,N_49158,N_49003);
nand U49374 (N_49374,N_49050,N_49234);
xor U49375 (N_49375,N_49042,N_49181);
or U49376 (N_49376,N_49021,N_49217);
and U49377 (N_49377,N_49037,N_49168);
nand U49378 (N_49378,N_49085,N_49184);
nand U49379 (N_49379,N_49009,N_49220);
and U49380 (N_49380,N_49203,N_49011);
or U49381 (N_49381,N_49121,N_49089);
or U49382 (N_49382,N_49230,N_49036);
and U49383 (N_49383,N_49153,N_49034);
nand U49384 (N_49384,N_49036,N_49059);
or U49385 (N_49385,N_49073,N_49120);
nand U49386 (N_49386,N_49085,N_49189);
nor U49387 (N_49387,N_49092,N_49220);
or U49388 (N_49388,N_49046,N_49237);
and U49389 (N_49389,N_49157,N_49197);
xnor U49390 (N_49390,N_49019,N_49039);
xnor U49391 (N_49391,N_49111,N_49094);
xor U49392 (N_49392,N_49135,N_49073);
nor U49393 (N_49393,N_49221,N_49030);
nand U49394 (N_49394,N_49033,N_49112);
xnor U49395 (N_49395,N_49104,N_49097);
or U49396 (N_49396,N_49220,N_49095);
or U49397 (N_49397,N_49240,N_49104);
and U49398 (N_49398,N_49167,N_49082);
nor U49399 (N_49399,N_49137,N_49169);
nor U49400 (N_49400,N_49096,N_49185);
or U49401 (N_49401,N_49228,N_49110);
nor U49402 (N_49402,N_49069,N_49199);
and U49403 (N_49403,N_49062,N_49063);
nand U49404 (N_49404,N_49174,N_49225);
nand U49405 (N_49405,N_49188,N_49032);
and U49406 (N_49406,N_49078,N_49198);
nand U49407 (N_49407,N_49030,N_49035);
xor U49408 (N_49408,N_49239,N_49116);
and U49409 (N_49409,N_49003,N_49088);
or U49410 (N_49410,N_49223,N_49026);
or U49411 (N_49411,N_49047,N_49072);
nand U49412 (N_49412,N_49093,N_49118);
nand U49413 (N_49413,N_49078,N_49152);
nor U49414 (N_49414,N_49116,N_49098);
xor U49415 (N_49415,N_49027,N_49111);
or U49416 (N_49416,N_49064,N_49242);
nand U49417 (N_49417,N_49205,N_49234);
nand U49418 (N_49418,N_49180,N_49170);
xnor U49419 (N_49419,N_49072,N_49142);
xnor U49420 (N_49420,N_49184,N_49177);
xor U49421 (N_49421,N_49067,N_49027);
or U49422 (N_49422,N_49205,N_49030);
xor U49423 (N_49423,N_49101,N_49109);
and U49424 (N_49424,N_49182,N_49044);
or U49425 (N_49425,N_49056,N_49157);
nand U49426 (N_49426,N_49218,N_49244);
xnor U49427 (N_49427,N_49003,N_49201);
nor U49428 (N_49428,N_49033,N_49012);
nand U49429 (N_49429,N_49200,N_49131);
and U49430 (N_49430,N_49176,N_49059);
nor U49431 (N_49431,N_49120,N_49067);
xnor U49432 (N_49432,N_49019,N_49078);
xor U49433 (N_49433,N_49067,N_49249);
and U49434 (N_49434,N_49144,N_49127);
and U49435 (N_49435,N_49055,N_49067);
nor U49436 (N_49436,N_49222,N_49141);
or U49437 (N_49437,N_49215,N_49165);
or U49438 (N_49438,N_49152,N_49035);
nand U49439 (N_49439,N_49171,N_49198);
nand U49440 (N_49440,N_49190,N_49145);
nor U49441 (N_49441,N_49181,N_49082);
and U49442 (N_49442,N_49012,N_49066);
or U49443 (N_49443,N_49134,N_49216);
or U49444 (N_49444,N_49019,N_49097);
or U49445 (N_49445,N_49079,N_49056);
or U49446 (N_49446,N_49041,N_49140);
nor U49447 (N_49447,N_49201,N_49061);
nor U49448 (N_49448,N_49060,N_49090);
xor U49449 (N_49449,N_49100,N_49031);
or U49450 (N_49450,N_49086,N_49044);
or U49451 (N_49451,N_49126,N_49083);
xnor U49452 (N_49452,N_49046,N_49241);
or U49453 (N_49453,N_49240,N_49213);
xor U49454 (N_49454,N_49226,N_49150);
xnor U49455 (N_49455,N_49058,N_49025);
or U49456 (N_49456,N_49216,N_49190);
and U49457 (N_49457,N_49244,N_49044);
and U49458 (N_49458,N_49103,N_49067);
nor U49459 (N_49459,N_49079,N_49015);
nand U49460 (N_49460,N_49075,N_49147);
xnor U49461 (N_49461,N_49227,N_49118);
or U49462 (N_49462,N_49072,N_49010);
xor U49463 (N_49463,N_49035,N_49130);
nand U49464 (N_49464,N_49023,N_49167);
xnor U49465 (N_49465,N_49000,N_49018);
nand U49466 (N_49466,N_49046,N_49239);
xor U49467 (N_49467,N_49164,N_49162);
or U49468 (N_49468,N_49055,N_49143);
nor U49469 (N_49469,N_49204,N_49060);
or U49470 (N_49470,N_49172,N_49231);
and U49471 (N_49471,N_49199,N_49125);
nand U49472 (N_49472,N_49130,N_49042);
and U49473 (N_49473,N_49211,N_49134);
nand U49474 (N_49474,N_49174,N_49067);
nor U49475 (N_49475,N_49246,N_49235);
and U49476 (N_49476,N_49185,N_49097);
or U49477 (N_49477,N_49060,N_49201);
xnor U49478 (N_49478,N_49048,N_49172);
and U49479 (N_49479,N_49157,N_49174);
or U49480 (N_49480,N_49082,N_49096);
xnor U49481 (N_49481,N_49140,N_49021);
or U49482 (N_49482,N_49193,N_49025);
or U49483 (N_49483,N_49074,N_49218);
xor U49484 (N_49484,N_49138,N_49053);
or U49485 (N_49485,N_49018,N_49231);
xnor U49486 (N_49486,N_49193,N_49018);
nand U49487 (N_49487,N_49120,N_49061);
nand U49488 (N_49488,N_49197,N_49172);
nand U49489 (N_49489,N_49052,N_49080);
or U49490 (N_49490,N_49043,N_49044);
nor U49491 (N_49491,N_49236,N_49176);
nand U49492 (N_49492,N_49169,N_49044);
or U49493 (N_49493,N_49198,N_49227);
nand U49494 (N_49494,N_49149,N_49151);
xor U49495 (N_49495,N_49160,N_49221);
nand U49496 (N_49496,N_49236,N_49198);
and U49497 (N_49497,N_49078,N_49069);
and U49498 (N_49498,N_49059,N_49077);
or U49499 (N_49499,N_49248,N_49035);
xnor U49500 (N_49500,N_49270,N_49384);
and U49501 (N_49501,N_49407,N_49309);
and U49502 (N_49502,N_49261,N_49341);
or U49503 (N_49503,N_49347,N_49281);
and U49504 (N_49504,N_49367,N_49269);
and U49505 (N_49505,N_49414,N_49410);
xnor U49506 (N_49506,N_49396,N_49420);
nand U49507 (N_49507,N_49417,N_49320);
xor U49508 (N_49508,N_49278,N_49326);
xor U49509 (N_49509,N_49291,N_49302);
nand U49510 (N_49510,N_49333,N_49354);
nor U49511 (N_49511,N_49352,N_49475);
xor U49512 (N_49512,N_49332,N_49345);
xnor U49513 (N_49513,N_49426,N_49455);
xor U49514 (N_49514,N_49469,N_49301);
nand U49515 (N_49515,N_49280,N_49365);
nand U49516 (N_49516,N_49342,N_49299);
nor U49517 (N_49517,N_49316,N_49292);
and U49518 (N_49518,N_49441,N_49380);
or U49519 (N_49519,N_49275,N_49449);
xnor U49520 (N_49520,N_49386,N_49321);
nor U49521 (N_49521,N_49256,N_49425);
nor U49522 (N_49522,N_49266,N_49436);
or U49523 (N_49523,N_49461,N_49418);
or U49524 (N_49524,N_49494,N_49412);
nor U49525 (N_49525,N_49390,N_49351);
xor U49526 (N_49526,N_49404,N_49328);
and U49527 (N_49527,N_49471,N_49374);
and U49528 (N_49528,N_49307,N_49327);
xnor U49529 (N_49529,N_49489,N_49388);
and U49530 (N_49530,N_49424,N_49429);
or U49531 (N_49531,N_49257,N_49498);
nor U49532 (N_49532,N_49479,N_49303);
xnor U49533 (N_49533,N_49437,N_49411);
or U49534 (N_49534,N_49274,N_49336);
xnor U49535 (N_49535,N_49346,N_49376);
and U49536 (N_49536,N_49446,N_49428);
xor U49537 (N_49537,N_49311,N_49491);
and U49538 (N_49538,N_49268,N_49381);
and U49539 (N_49539,N_49325,N_49285);
nor U49540 (N_49540,N_49392,N_49402);
or U49541 (N_49541,N_49403,N_49416);
nand U49542 (N_49542,N_49393,N_49370);
and U49543 (N_49543,N_49443,N_49298);
xor U49544 (N_49544,N_49377,N_49276);
and U49545 (N_49545,N_49456,N_49331);
or U49546 (N_49546,N_49375,N_49366);
nand U49547 (N_49547,N_49277,N_49383);
xor U49548 (N_49548,N_49305,N_49379);
and U49549 (N_49549,N_49259,N_49310);
xor U49550 (N_49550,N_49427,N_49460);
or U49551 (N_49551,N_49435,N_49415);
or U49552 (N_49552,N_49401,N_49398);
or U49553 (N_49553,N_49265,N_49294);
or U49554 (N_49554,N_49260,N_49431);
nor U49555 (N_49555,N_49438,N_49329);
nand U49556 (N_49556,N_49286,N_49391);
nor U49557 (N_49557,N_49434,N_49335);
xnor U49558 (N_49558,N_49338,N_49382);
nor U49559 (N_49559,N_49421,N_49451);
or U49560 (N_49560,N_49452,N_49394);
xnor U49561 (N_49561,N_49348,N_49314);
nand U49562 (N_49562,N_49323,N_49355);
xor U49563 (N_49563,N_49363,N_49293);
or U49564 (N_49564,N_49272,N_49462);
and U49565 (N_49565,N_49319,N_49350);
nor U49566 (N_49566,N_49330,N_49306);
xnor U49567 (N_49567,N_49444,N_49251);
nand U49568 (N_49568,N_49495,N_49397);
xnor U49569 (N_49569,N_49254,N_49487);
nand U49570 (N_49570,N_49480,N_49468);
and U49571 (N_49571,N_49344,N_49334);
and U49572 (N_49572,N_49357,N_49486);
nor U49573 (N_49573,N_49463,N_49317);
or U49574 (N_49574,N_49283,N_49490);
and U49575 (N_49575,N_49454,N_49297);
nor U49576 (N_49576,N_49282,N_49408);
and U49577 (N_49577,N_49478,N_49253);
or U49578 (N_49578,N_49409,N_49296);
xor U49579 (N_49579,N_49358,N_49343);
xor U49580 (N_49580,N_49440,N_49324);
or U49581 (N_49581,N_49493,N_49442);
or U49582 (N_49582,N_49273,N_49385);
or U49583 (N_49583,N_49279,N_49477);
and U49584 (N_49584,N_49371,N_49264);
and U49585 (N_49585,N_49322,N_49483);
nor U49586 (N_49586,N_49308,N_49387);
or U49587 (N_49587,N_49473,N_49476);
xor U49588 (N_49588,N_49423,N_49439);
nand U49589 (N_49589,N_49482,N_49422);
xnor U49590 (N_49590,N_49368,N_49406);
and U49591 (N_49591,N_49481,N_49389);
xnor U49592 (N_49592,N_49399,N_49361);
nor U49593 (N_49593,N_49252,N_49372);
nor U49594 (N_49594,N_49450,N_49405);
xor U49595 (N_49595,N_49413,N_49267);
and U49596 (N_49596,N_49432,N_49378);
and U49597 (N_49597,N_49349,N_49304);
and U49598 (N_49598,N_49395,N_49464);
nor U49599 (N_49599,N_49289,N_49430);
xor U49600 (N_49600,N_49499,N_49359);
nand U49601 (N_49601,N_49445,N_49467);
nand U49602 (N_49602,N_49356,N_49447);
or U49603 (N_49603,N_49258,N_49492);
or U49604 (N_49604,N_49474,N_49496);
xor U49605 (N_49605,N_49488,N_49312);
or U49606 (N_49606,N_49340,N_49470);
and U49607 (N_49607,N_49458,N_49448);
or U49608 (N_49608,N_49369,N_49262);
xor U49609 (N_49609,N_49315,N_49295);
xnor U49610 (N_49610,N_49484,N_49290);
xor U49611 (N_49611,N_49300,N_49453);
and U49612 (N_49612,N_49419,N_49339);
and U49613 (N_49613,N_49313,N_49263);
xnor U49614 (N_49614,N_49485,N_49360);
xor U49615 (N_49615,N_49255,N_49459);
nor U49616 (N_49616,N_49364,N_49465);
or U49617 (N_49617,N_49373,N_49433);
and U49618 (N_49618,N_49472,N_49457);
nor U49619 (N_49619,N_49284,N_49400);
nand U49620 (N_49620,N_49337,N_49318);
and U49621 (N_49621,N_49271,N_49250);
nor U49622 (N_49622,N_49353,N_49287);
or U49623 (N_49623,N_49362,N_49497);
xor U49624 (N_49624,N_49466,N_49288);
nor U49625 (N_49625,N_49348,N_49355);
nor U49626 (N_49626,N_49377,N_49473);
nand U49627 (N_49627,N_49354,N_49360);
and U49628 (N_49628,N_49354,N_49400);
and U49629 (N_49629,N_49254,N_49300);
nand U49630 (N_49630,N_49397,N_49385);
nor U49631 (N_49631,N_49363,N_49375);
xnor U49632 (N_49632,N_49250,N_49461);
and U49633 (N_49633,N_49250,N_49251);
nor U49634 (N_49634,N_49253,N_49379);
or U49635 (N_49635,N_49328,N_49443);
xnor U49636 (N_49636,N_49423,N_49369);
and U49637 (N_49637,N_49257,N_49264);
or U49638 (N_49638,N_49376,N_49317);
or U49639 (N_49639,N_49288,N_49451);
nor U49640 (N_49640,N_49336,N_49466);
and U49641 (N_49641,N_49261,N_49443);
and U49642 (N_49642,N_49444,N_49254);
nor U49643 (N_49643,N_49478,N_49272);
or U49644 (N_49644,N_49383,N_49293);
or U49645 (N_49645,N_49414,N_49304);
nor U49646 (N_49646,N_49387,N_49292);
nor U49647 (N_49647,N_49309,N_49300);
nor U49648 (N_49648,N_49445,N_49327);
and U49649 (N_49649,N_49374,N_49393);
nand U49650 (N_49650,N_49283,N_49292);
nor U49651 (N_49651,N_49478,N_49340);
or U49652 (N_49652,N_49432,N_49416);
xnor U49653 (N_49653,N_49454,N_49408);
nor U49654 (N_49654,N_49331,N_49409);
or U49655 (N_49655,N_49434,N_49393);
nand U49656 (N_49656,N_49495,N_49479);
or U49657 (N_49657,N_49401,N_49353);
and U49658 (N_49658,N_49494,N_49253);
and U49659 (N_49659,N_49437,N_49266);
nor U49660 (N_49660,N_49398,N_49460);
xnor U49661 (N_49661,N_49377,N_49302);
or U49662 (N_49662,N_49305,N_49355);
nor U49663 (N_49663,N_49308,N_49384);
nor U49664 (N_49664,N_49417,N_49419);
or U49665 (N_49665,N_49331,N_49376);
xor U49666 (N_49666,N_49288,N_49254);
nor U49667 (N_49667,N_49416,N_49327);
and U49668 (N_49668,N_49261,N_49296);
nor U49669 (N_49669,N_49367,N_49471);
nand U49670 (N_49670,N_49340,N_49450);
nor U49671 (N_49671,N_49397,N_49250);
nor U49672 (N_49672,N_49297,N_49307);
or U49673 (N_49673,N_49418,N_49252);
xor U49674 (N_49674,N_49408,N_49446);
and U49675 (N_49675,N_49487,N_49493);
or U49676 (N_49676,N_49481,N_49257);
or U49677 (N_49677,N_49294,N_49498);
and U49678 (N_49678,N_49376,N_49480);
nor U49679 (N_49679,N_49497,N_49477);
and U49680 (N_49680,N_49257,N_49275);
nand U49681 (N_49681,N_49321,N_49270);
and U49682 (N_49682,N_49255,N_49351);
nor U49683 (N_49683,N_49311,N_49376);
and U49684 (N_49684,N_49396,N_49474);
nand U49685 (N_49685,N_49420,N_49252);
nand U49686 (N_49686,N_49379,N_49327);
nand U49687 (N_49687,N_49356,N_49340);
or U49688 (N_49688,N_49274,N_49258);
nor U49689 (N_49689,N_49480,N_49319);
nor U49690 (N_49690,N_49422,N_49321);
and U49691 (N_49691,N_49456,N_49408);
or U49692 (N_49692,N_49495,N_49296);
nand U49693 (N_49693,N_49252,N_49317);
and U49694 (N_49694,N_49272,N_49460);
nand U49695 (N_49695,N_49358,N_49315);
xnor U49696 (N_49696,N_49438,N_49275);
and U49697 (N_49697,N_49323,N_49421);
and U49698 (N_49698,N_49363,N_49351);
or U49699 (N_49699,N_49352,N_49351);
xnor U49700 (N_49700,N_49360,N_49405);
and U49701 (N_49701,N_49371,N_49451);
or U49702 (N_49702,N_49443,N_49485);
and U49703 (N_49703,N_49454,N_49271);
nand U49704 (N_49704,N_49260,N_49314);
nor U49705 (N_49705,N_49370,N_49318);
nand U49706 (N_49706,N_49482,N_49471);
nor U49707 (N_49707,N_49442,N_49282);
or U49708 (N_49708,N_49438,N_49373);
and U49709 (N_49709,N_49434,N_49345);
and U49710 (N_49710,N_49341,N_49325);
nor U49711 (N_49711,N_49461,N_49339);
xnor U49712 (N_49712,N_49499,N_49343);
nor U49713 (N_49713,N_49338,N_49440);
nand U49714 (N_49714,N_49263,N_49279);
xor U49715 (N_49715,N_49458,N_49271);
nand U49716 (N_49716,N_49420,N_49416);
nor U49717 (N_49717,N_49344,N_49363);
nand U49718 (N_49718,N_49459,N_49447);
and U49719 (N_49719,N_49391,N_49389);
and U49720 (N_49720,N_49281,N_49415);
nor U49721 (N_49721,N_49425,N_49447);
xnor U49722 (N_49722,N_49474,N_49472);
nor U49723 (N_49723,N_49425,N_49294);
nand U49724 (N_49724,N_49259,N_49337);
xnor U49725 (N_49725,N_49287,N_49493);
nor U49726 (N_49726,N_49339,N_49483);
xnor U49727 (N_49727,N_49419,N_49402);
nand U49728 (N_49728,N_49494,N_49405);
or U49729 (N_49729,N_49343,N_49303);
nor U49730 (N_49730,N_49267,N_49404);
and U49731 (N_49731,N_49427,N_49413);
or U49732 (N_49732,N_49417,N_49300);
xnor U49733 (N_49733,N_49471,N_49255);
nand U49734 (N_49734,N_49443,N_49255);
nor U49735 (N_49735,N_49362,N_49425);
and U49736 (N_49736,N_49495,N_49422);
or U49737 (N_49737,N_49372,N_49344);
nor U49738 (N_49738,N_49482,N_49295);
nor U49739 (N_49739,N_49460,N_49334);
nor U49740 (N_49740,N_49382,N_49455);
nor U49741 (N_49741,N_49493,N_49267);
nor U49742 (N_49742,N_49421,N_49284);
or U49743 (N_49743,N_49264,N_49263);
or U49744 (N_49744,N_49316,N_49423);
nand U49745 (N_49745,N_49377,N_49419);
and U49746 (N_49746,N_49358,N_49296);
xor U49747 (N_49747,N_49419,N_49426);
or U49748 (N_49748,N_49404,N_49311);
nand U49749 (N_49749,N_49422,N_49309);
nor U49750 (N_49750,N_49702,N_49685);
nand U49751 (N_49751,N_49543,N_49654);
nor U49752 (N_49752,N_49738,N_49650);
xnor U49753 (N_49753,N_49540,N_49668);
and U49754 (N_49754,N_49512,N_49730);
and U49755 (N_49755,N_49719,N_49595);
nor U49756 (N_49756,N_49708,N_49601);
or U49757 (N_49757,N_49693,N_49676);
nand U49758 (N_49758,N_49602,N_49529);
xnor U49759 (N_49759,N_49617,N_49591);
xnor U49760 (N_49760,N_49694,N_49735);
nor U49761 (N_49761,N_49727,N_49532);
nor U49762 (N_49762,N_49633,N_49689);
and U49763 (N_49763,N_49516,N_49651);
or U49764 (N_49764,N_49639,N_49579);
xnor U49765 (N_49765,N_49523,N_49544);
nor U49766 (N_49766,N_49627,N_49582);
xnor U49767 (N_49767,N_49570,N_49691);
or U49768 (N_49768,N_49722,N_49636);
or U49769 (N_49769,N_49548,N_49649);
and U49770 (N_49770,N_49584,N_49632);
xnor U49771 (N_49771,N_49561,N_49553);
and U49772 (N_49772,N_49747,N_49521);
nand U49773 (N_49773,N_49531,N_49625);
or U49774 (N_49774,N_49736,N_49733);
or U49775 (N_49775,N_49509,N_49552);
xnor U49776 (N_49776,N_49661,N_49678);
nand U49777 (N_49777,N_49669,N_49593);
xnor U49778 (N_49778,N_49729,N_49506);
xor U49779 (N_49779,N_49671,N_49630);
nand U49780 (N_49780,N_49674,N_49711);
or U49781 (N_49781,N_49684,N_49728);
nand U49782 (N_49782,N_49605,N_49610);
and U49783 (N_49783,N_49742,N_49511);
nand U49784 (N_49784,N_49551,N_49594);
nor U49785 (N_49785,N_49657,N_49589);
or U49786 (N_49786,N_49637,N_49745);
nand U49787 (N_49787,N_49624,N_49581);
xor U49788 (N_49788,N_49635,N_49629);
xnor U49789 (N_49789,N_49740,N_49749);
and U49790 (N_49790,N_49704,N_49718);
nand U49791 (N_49791,N_49717,N_49574);
or U49792 (N_49792,N_49500,N_49638);
nor U49793 (N_49793,N_49703,N_49746);
nand U49794 (N_49794,N_49670,N_49712);
or U49795 (N_49795,N_49731,N_49588);
xnor U49796 (N_49796,N_49677,N_49664);
nor U49797 (N_49797,N_49599,N_49628);
and U49798 (N_49798,N_49675,N_49501);
nand U49799 (N_49799,N_49520,N_49707);
xnor U49800 (N_49800,N_49616,N_49504);
and U49801 (N_49801,N_49518,N_49695);
nand U49802 (N_49802,N_49573,N_49541);
and U49803 (N_49803,N_49600,N_49580);
and U49804 (N_49804,N_49748,N_49549);
or U49805 (N_49805,N_49560,N_49534);
nand U49806 (N_49806,N_49732,N_49655);
nand U49807 (N_49807,N_49725,N_49585);
and U49808 (N_49808,N_49696,N_49699);
or U49809 (N_49809,N_49612,N_49620);
nor U49810 (N_49810,N_49556,N_49557);
or U49811 (N_49811,N_49713,N_49503);
and U49812 (N_49812,N_49744,N_49608);
or U49813 (N_49813,N_49537,N_49538);
nor U49814 (N_49814,N_49653,N_49575);
xor U49815 (N_49815,N_49568,N_49542);
nand U49816 (N_49816,N_49586,N_49663);
and U49817 (N_49817,N_49646,N_49641);
nor U49818 (N_49818,N_49592,N_49618);
or U49819 (N_49819,N_49614,N_49715);
and U49820 (N_49820,N_49527,N_49507);
or U49821 (N_49821,N_49720,N_49710);
or U49822 (N_49822,N_49564,N_49621);
nand U49823 (N_49823,N_49539,N_49578);
and U49824 (N_49824,N_49697,N_49567);
xor U49825 (N_49825,N_49554,N_49606);
xor U49826 (N_49826,N_49563,N_49645);
xor U49827 (N_49827,N_49739,N_49598);
and U49828 (N_49828,N_49626,N_49513);
or U49829 (N_49829,N_49743,N_49686);
or U49830 (N_49830,N_49660,N_49546);
nand U49831 (N_49831,N_49596,N_49615);
or U49832 (N_49832,N_49652,N_49700);
nor U49833 (N_49833,N_49648,N_49672);
or U49834 (N_49834,N_49536,N_49545);
and U49835 (N_49835,N_49643,N_49514);
xor U49836 (N_49836,N_49692,N_49709);
or U49837 (N_49837,N_49623,N_49622);
nand U49838 (N_49838,N_49666,N_49665);
nand U49839 (N_49839,N_49519,N_49611);
xnor U49840 (N_49840,N_49688,N_49690);
xor U49841 (N_49841,N_49714,N_49662);
nor U49842 (N_49842,N_49634,N_49656);
nand U49843 (N_49843,N_49547,N_49644);
or U49844 (N_49844,N_49555,N_49642);
nand U49845 (N_49845,N_49682,N_49524);
nor U49846 (N_49846,N_49515,N_49525);
nand U49847 (N_49847,N_49680,N_49631);
nor U49848 (N_49848,N_49530,N_49522);
xor U49849 (N_49849,N_49679,N_49597);
and U49850 (N_49850,N_49559,N_49706);
nor U49851 (N_49851,N_49683,N_49647);
or U49852 (N_49852,N_49619,N_49659);
nor U49853 (N_49853,N_49658,N_49566);
nand U49854 (N_49854,N_49741,N_49528);
nand U49855 (N_49855,N_49673,N_49577);
and U49856 (N_49856,N_49737,N_49572);
or U49857 (N_49857,N_49510,N_49604);
nand U49858 (N_49858,N_49550,N_49502);
nand U49859 (N_49859,N_49590,N_49734);
nand U49860 (N_49860,N_49716,N_49558);
or U49861 (N_49861,N_49569,N_49640);
and U49862 (N_49862,N_49565,N_49533);
nand U49863 (N_49863,N_49607,N_49517);
xor U49864 (N_49864,N_49508,N_49721);
and U49865 (N_49865,N_49613,N_49705);
and U49866 (N_49866,N_49609,N_49667);
xor U49867 (N_49867,N_49576,N_49583);
and U49868 (N_49868,N_49571,N_49723);
xnor U49869 (N_49869,N_49535,N_49603);
and U49870 (N_49870,N_49698,N_49526);
nand U49871 (N_49871,N_49724,N_49505);
nand U49872 (N_49872,N_49681,N_49687);
nand U49873 (N_49873,N_49701,N_49587);
and U49874 (N_49874,N_49726,N_49562);
nor U49875 (N_49875,N_49652,N_49695);
and U49876 (N_49876,N_49655,N_49694);
or U49877 (N_49877,N_49736,N_49740);
and U49878 (N_49878,N_49626,N_49569);
xor U49879 (N_49879,N_49720,N_49695);
xor U49880 (N_49880,N_49562,N_49591);
xnor U49881 (N_49881,N_49641,N_49703);
and U49882 (N_49882,N_49738,N_49565);
and U49883 (N_49883,N_49738,N_49633);
and U49884 (N_49884,N_49747,N_49738);
or U49885 (N_49885,N_49601,N_49615);
nor U49886 (N_49886,N_49534,N_49716);
or U49887 (N_49887,N_49578,N_49597);
nand U49888 (N_49888,N_49532,N_49521);
or U49889 (N_49889,N_49728,N_49749);
and U49890 (N_49890,N_49555,N_49684);
xor U49891 (N_49891,N_49699,N_49520);
or U49892 (N_49892,N_49676,N_49569);
xnor U49893 (N_49893,N_49671,N_49560);
xnor U49894 (N_49894,N_49628,N_49506);
nor U49895 (N_49895,N_49658,N_49746);
or U49896 (N_49896,N_49610,N_49526);
nand U49897 (N_49897,N_49617,N_49717);
nor U49898 (N_49898,N_49744,N_49661);
nor U49899 (N_49899,N_49632,N_49540);
xnor U49900 (N_49900,N_49683,N_49574);
nor U49901 (N_49901,N_49659,N_49687);
xor U49902 (N_49902,N_49504,N_49617);
nor U49903 (N_49903,N_49618,N_49666);
or U49904 (N_49904,N_49510,N_49624);
nor U49905 (N_49905,N_49538,N_49611);
and U49906 (N_49906,N_49748,N_49650);
and U49907 (N_49907,N_49525,N_49638);
and U49908 (N_49908,N_49587,N_49644);
nor U49909 (N_49909,N_49620,N_49696);
nand U49910 (N_49910,N_49539,N_49536);
or U49911 (N_49911,N_49583,N_49637);
nand U49912 (N_49912,N_49557,N_49552);
nor U49913 (N_49913,N_49519,N_49710);
and U49914 (N_49914,N_49569,N_49673);
xor U49915 (N_49915,N_49598,N_49714);
or U49916 (N_49916,N_49685,N_49649);
and U49917 (N_49917,N_49531,N_49548);
and U49918 (N_49918,N_49504,N_49615);
or U49919 (N_49919,N_49689,N_49703);
or U49920 (N_49920,N_49503,N_49614);
and U49921 (N_49921,N_49587,N_49744);
nand U49922 (N_49922,N_49719,N_49567);
or U49923 (N_49923,N_49717,N_49516);
or U49924 (N_49924,N_49684,N_49517);
and U49925 (N_49925,N_49733,N_49681);
nand U49926 (N_49926,N_49502,N_49666);
xor U49927 (N_49927,N_49530,N_49502);
nand U49928 (N_49928,N_49622,N_49684);
and U49929 (N_49929,N_49623,N_49597);
xnor U49930 (N_49930,N_49583,N_49704);
nand U49931 (N_49931,N_49624,N_49674);
nor U49932 (N_49932,N_49662,N_49674);
nor U49933 (N_49933,N_49618,N_49531);
nand U49934 (N_49934,N_49626,N_49724);
and U49935 (N_49935,N_49500,N_49600);
nor U49936 (N_49936,N_49620,N_49590);
nand U49937 (N_49937,N_49511,N_49719);
xnor U49938 (N_49938,N_49566,N_49623);
and U49939 (N_49939,N_49731,N_49535);
xor U49940 (N_49940,N_49729,N_49657);
and U49941 (N_49941,N_49726,N_49579);
nor U49942 (N_49942,N_49514,N_49552);
nand U49943 (N_49943,N_49614,N_49561);
and U49944 (N_49944,N_49749,N_49585);
xor U49945 (N_49945,N_49689,N_49600);
nor U49946 (N_49946,N_49606,N_49743);
nand U49947 (N_49947,N_49548,N_49674);
and U49948 (N_49948,N_49546,N_49733);
and U49949 (N_49949,N_49561,N_49740);
nor U49950 (N_49950,N_49607,N_49673);
nand U49951 (N_49951,N_49531,N_49717);
and U49952 (N_49952,N_49560,N_49565);
nor U49953 (N_49953,N_49631,N_49660);
xor U49954 (N_49954,N_49715,N_49703);
and U49955 (N_49955,N_49593,N_49531);
xnor U49956 (N_49956,N_49727,N_49520);
nand U49957 (N_49957,N_49707,N_49690);
nand U49958 (N_49958,N_49575,N_49536);
xor U49959 (N_49959,N_49500,N_49699);
or U49960 (N_49960,N_49522,N_49567);
and U49961 (N_49961,N_49506,N_49605);
nor U49962 (N_49962,N_49699,N_49518);
or U49963 (N_49963,N_49500,N_49621);
nor U49964 (N_49964,N_49656,N_49708);
xor U49965 (N_49965,N_49682,N_49665);
or U49966 (N_49966,N_49616,N_49678);
nand U49967 (N_49967,N_49703,N_49533);
or U49968 (N_49968,N_49613,N_49647);
nand U49969 (N_49969,N_49704,N_49501);
or U49970 (N_49970,N_49625,N_49732);
nand U49971 (N_49971,N_49730,N_49667);
nor U49972 (N_49972,N_49743,N_49734);
xor U49973 (N_49973,N_49540,N_49687);
nor U49974 (N_49974,N_49540,N_49562);
nand U49975 (N_49975,N_49543,N_49708);
or U49976 (N_49976,N_49628,N_49564);
nand U49977 (N_49977,N_49698,N_49684);
and U49978 (N_49978,N_49645,N_49622);
nor U49979 (N_49979,N_49709,N_49565);
nand U49980 (N_49980,N_49517,N_49626);
or U49981 (N_49981,N_49629,N_49706);
and U49982 (N_49982,N_49543,N_49566);
and U49983 (N_49983,N_49589,N_49708);
and U49984 (N_49984,N_49638,N_49563);
xor U49985 (N_49985,N_49501,N_49693);
nand U49986 (N_49986,N_49595,N_49557);
nand U49987 (N_49987,N_49716,N_49693);
xor U49988 (N_49988,N_49553,N_49728);
nand U49989 (N_49989,N_49598,N_49552);
and U49990 (N_49990,N_49701,N_49731);
or U49991 (N_49991,N_49597,N_49504);
nor U49992 (N_49992,N_49605,N_49572);
xnor U49993 (N_49993,N_49722,N_49547);
nor U49994 (N_49994,N_49530,N_49599);
nand U49995 (N_49995,N_49621,N_49525);
xor U49996 (N_49996,N_49703,N_49530);
or U49997 (N_49997,N_49639,N_49719);
xor U49998 (N_49998,N_49649,N_49619);
or U49999 (N_49999,N_49658,N_49535);
or UO_0 (O_0,N_49944,N_49757);
nand UO_1 (O_1,N_49963,N_49943);
or UO_2 (O_2,N_49873,N_49761);
or UO_3 (O_3,N_49758,N_49980);
nor UO_4 (O_4,N_49966,N_49784);
and UO_5 (O_5,N_49998,N_49799);
nand UO_6 (O_6,N_49831,N_49989);
nand UO_7 (O_7,N_49935,N_49789);
or UO_8 (O_8,N_49820,N_49934);
nor UO_9 (O_9,N_49952,N_49882);
or UO_10 (O_10,N_49792,N_49876);
and UO_11 (O_11,N_49996,N_49920);
xnor UO_12 (O_12,N_49833,N_49970);
xnor UO_13 (O_13,N_49986,N_49909);
and UO_14 (O_14,N_49810,N_49767);
nand UO_15 (O_15,N_49990,N_49959);
and UO_16 (O_16,N_49913,N_49903);
nand UO_17 (O_17,N_49933,N_49777);
nand UO_18 (O_18,N_49973,N_49778);
and UO_19 (O_19,N_49886,N_49848);
and UO_20 (O_20,N_49866,N_49826);
xnor UO_21 (O_21,N_49864,N_49994);
and UO_22 (O_22,N_49905,N_49861);
nand UO_23 (O_23,N_49960,N_49962);
xor UO_24 (O_24,N_49993,N_49982);
nor UO_25 (O_25,N_49830,N_49981);
nand UO_26 (O_26,N_49971,N_49768);
or UO_27 (O_27,N_49954,N_49921);
nor UO_28 (O_28,N_49991,N_49754);
xor UO_29 (O_29,N_49797,N_49992);
nand UO_30 (O_30,N_49819,N_49798);
nor UO_31 (O_31,N_49849,N_49919);
nor UO_32 (O_32,N_49813,N_49822);
or UO_33 (O_33,N_49958,N_49891);
or UO_34 (O_34,N_49785,N_49773);
nand UO_35 (O_35,N_49832,N_49979);
or UO_36 (O_36,N_49926,N_49805);
and UO_37 (O_37,N_49786,N_49915);
xor UO_38 (O_38,N_49867,N_49751);
xnor UO_39 (O_39,N_49840,N_49829);
xnor UO_40 (O_40,N_49923,N_49776);
or UO_41 (O_41,N_49818,N_49899);
xor UO_42 (O_42,N_49850,N_49951);
nor UO_43 (O_43,N_49756,N_49955);
or UO_44 (O_44,N_49922,N_49760);
or UO_45 (O_45,N_49846,N_49937);
nor UO_46 (O_46,N_49801,N_49869);
or UO_47 (O_47,N_49878,N_49775);
xor UO_48 (O_48,N_49800,N_49811);
or UO_49 (O_49,N_49824,N_49835);
nor UO_50 (O_50,N_49875,N_49770);
xnor UO_51 (O_51,N_49780,N_49918);
or UO_52 (O_52,N_49950,N_49807);
and UO_53 (O_53,N_49839,N_49927);
xor UO_54 (O_54,N_49852,N_49974);
nand UO_55 (O_55,N_49942,N_49774);
xnor UO_56 (O_56,N_49984,N_49803);
xor UO_57 (O_57,N_49881,N_49834);
or UO_58 (O_58,N_49844,N_49809);
nor UO_59 (O_59,N_49936,N_49940);
or UO_60 (O_60,N_49985,N_49945);
or UO_61 (O_61,N_49977,N_49892);
nor UO_62 (O_62,N_49925,N_49860);
or UO_63 (O_63,N_49791,N_49859);
nand UO_64 (O_64,N_49978,N_49872);
and UO_65 (O_65,N_49788,N_49947);
xnor UO_66 (O_66,N_49825,N_49908);
xor UO_67 (O_67,N_49928,N_49750);
nor UO_68 (O_68,N_49972,N_49888);
nand UO_69 (O_69,N_49781,N_49783);
nor UO_70 (O_70,N_49790,N_49865);
nor UO_71 (O_71,N_49896,N_49828);
xnor UO_72 (O_72,N_49912,N_49975);
nand UO_73 (O_73,N_49956,N_49893);
nor UO_74 (O_74,N_49999,N_49890);
or UO_75 (O_75,N_49874,N_49957);
nor UO_76 (O_76,N_49794,N_49766);
nor UO_77 (O_77,N_49900,N_49763);
xnor UO_78 (O_78,N_49983,N_49806);
and UO_79 (O_79,N_49887,N_49988);
xor UO_80 (O_80,N_49939,N_49862);
or UO_81 (O_81,N_49858,N_49845);
and UO_82 (O_82,N_49949,N_49787);
and UO_83 (O_83,N_49817,N_49910);
xor UO_84 (O_84,N_49965,N_49837);
nand UO_85 (O_85,N_49968,N_49827);
nor UO_86 (O_86,N_49863,N_49821);
nand UO_87 (O_87,N_49895,N_49883);
and UO_88 (O_88,N_49847,N_49841);
xnor UO_89 (O_89,N_49857,N_49901);
or UO_90 (O_90,N_49953,N_49853);
and UO_91 (O_91,N_49843,N_49997);
or UO_92 (O_92,N_49964,N_49894);
or UO_93 (O_93,N_49884,N_49836);
nand UO_94 (O_94,N_49976,N_49880);
nand UO_95 (O_95,N_49995,N_49842);
nor UO_96 (O_96,N_49816,N_49904);
xnor UO_97 (O_97,N_49948,N_49795);
xnor UO_98 (O_98,N_49987,N_49897);
nor UO_99 (O_99,N_49856,N_49782);
xor UO_100 (O_100,N_49779,N_49932);
nor UO_101 (O_101,N_49814,N_49914);
or UO_102 (O_102,N_49885,N_49838);
xnor UO_103 (O_103,N_49815,N_49796);
nor UO_104 (O_104,N_49911,N_49772);
or UO_105 (O_105,N_49906,N_49946);
nand UO_106 (O_106,N_49855,N_49967);
and UO_107 (O_107,N_49931,N_49907);
nor UO_108 (O_108,N_49879,N_49793);
nor UO_109 (O_109,N_49812,N_49930);
or UO_110 (O_110,N_49802,N_49969);
xnor UO_111 (O_111,N_49941,N_49769);
nand UO_112 (O_112,N_49808,N_49771);
nand UO_113 (O_113,N_49902,N_49961);
or UO_114 (O_114,N_49917,N_49898);
or UO_115 (O_115,N_49755,N_49854);
xnor UO_116 (O_116,N_49938,N_49765);
nor UO_117 (O_117,N_49823,N_49924);
xor UO_118 (O_118,N_49804,N_49762);
xnor UO_119 (O_119,N_49870,N_49752);
nand UO_120 (O_120,N_49753,N_49871);
nor UO_121 (O_121,N_49877,N_49868);
nor UO_122 (O_122,N_49764,N_49759);
nand UO_123 (O_123,N_49929,N_49851);
nand UO_124 (O_124,N_49916,N_49889);
and UO_125 (O_125,N_49961,N_49976);
nor UO_126 (O_126,N_49956,N_49799);
nand UO_127 (O_127,N_49945,N_49900);
and UO_128 (O_128,N_49873,N_49890);
and UO_129 (O_129,N_49969,N_49890);
nand UO_130 (O_130,N_49943,N_49925);
or UO_131 (O_131,N_49840,N_49751);
xor UO_132 (O_132,N_49890,N_49966);
xnor UO_133 (O_133,N_49862,N_49971);
nand UO_134 (O_134,N_49830,N_49870);
nor UO_135 (O_135,N_49840,N_49834);
xnor UO_136 (O_136,N_49784,N_49997);
nand UO_137 (O_137,N_49794,N_49863);
nor UO_138 (O_138,N_49792,N_49963);
and UO_139 (O_139,N_49755,N_49935);
or UO_140 (O_140,N_49777,N_49904);
and UO_141 (O_141,N_49905,N_49758);
or UO_142 (O_142,N_49750,N_49904);
or UO_143 (O_143,N_49849,N_49997);
or UO_144 (O_144,N_49770,N_49888);
nor UO_145 (O_145,N_49852,N_49927);
nand UO_146 (O_146,N_49833,N_49926);
and UO_147 (O_147,N_49912,N_49982);
and UO_148 (O_148,N_49835,N_49892);
or UO_149 (O_149,N_49915,N_49798);
xnor UO_150 (O_150,N_49858,N_49902);
or UO_151 (O_151,N_49814,N_49888);
nand UO_152 (O_152,N_49757,N_49776);
and UO_153 (O_153,N_49930,N_49938);
xor UO_154 (O_154,N_49915,N_49783);
or UO_155 (O_155,N_49978,N_49907);
xor UO_156 (O_156,N_49851,N_49817);
xnor UO_157 (O_157,N_49750,N_49826);
nor UO_158 (O_158,N_49907,N_49996);
or UO_159 (O_159,N_49897,N_49836);
or UO_160 (O_160,N_49994,N_49946);
and UO_161 (O_161,N_49775,N_49965);
or UO_162 (O_162,N_49788,N_49962);
nor UO_163 (O_163,N_49754,N_49837);
nand UO_164 (O_164,N_49863,N_49828);
or UO_165 (O_165,N_49862,N_49970);
nor UO_166 (O_166,N_49973,N_49861);
nand UO_167 (O_167,N_49996,N_49835);
nand UO_168 (O_168,N_49793,N_49813);
and UO_169 (O_169,N_49793,N_49847);
and UO_170 (O_170,N_49944,N_49808);
and UO_171 (O_171,N_49881,N_49763);
and UO_172 (O_172,N_49801,N_49813);
nor UO_173 (O_173,N_49832,N_49960);
xor UO_174 (O_174,N_49750,N_49982);
and UO_175 (O_175,N_49874,N_49953);
nor UO_176 (O_176,N_49916,N_49899);
xor UO_177 (O_177,N_49928,N_49950);
xor UO_178 (O_178,N_49916,N_49984);
or UO_179 (O_179,N_49854,N_49909);
xnor UO_180 (O_180,N_49902,N_49799);
and UO_181 (O_181,N_49878,N_49923);
nor UO_182 (O_182,N_49837,N_49850);
nand UO_183 (O_183,N_49921,N_49876);
nor UO_184 (O_184,N_49835,N_49843);
xor UO_185 (O_185,N_49811,N_49780);
and UO_186 (O_186,N_49834,N_49933);
and UO_187 (O_187,N_49896,N_49836);
xor UO_188 (O_188,N_49751,N_49918);
nor UO_189 (O_189,N_49880,N_49968);
or UO_190 (O_190,N_49801,N_49930);
nor UO_191 (O_191,N_49982,N_49987);
xor UO_192 (O_192,N_49935,N_49763);
and UO_193 (O_193,N_49970,N_49853);
xor UO_194 (O_194,N_49977,N_49981);
nand UO_195 (O_195,N_49788,N_49988);
nor UO_196 (O_196,N_49880,N_49825);
or UO_197 (O_197,N_49919,N_49841);
or UO_198 (O_198,N_49835,N_49906);
and UO_199 (O_199,N_49971,N_49882);
or UO_200 (O_200,N_49771,N_49957);
nor UO_201 (O_201,N_49871,N_49771);
xor UO_202 (O_202,N_49986,N_49951);
nor UO_203 (O_203,N_49760,N_49814);
nand UO_204 (O_204,N_49877,N_49904);
nand UO_205 (O_205,N_49934,N_49802);
nand UO_206 (O_206,N_49993,N_49923);
nor UO_207 (O_207,N_49941,N_49953);
and UO_208 (O_208,N_49930,N_49811);
xor UO_209 (O_209,N_49815,N_49851);
and UO_210 (O_210,N_49800,N_49927);
or UO_211 (O_211,N_49877,N_49796);
or UO_212 (O_212,N_49762,N_49866);
or UO_213 (O_213,N_49894,N_49789);
and UO_214 (O_214,N_49945,N_49915);
or UO_215 (O_215,N_49769,N_49795);
and UO_216 (O_216,N_49946,N_49764);
nor UO_217 (O_217,N_49770,N_49788);
nor UO_218 (O_218,N_49937,N_49953);
and UO_219 (O_219,N_49831,N_49822);
and UO_220 (O_220,N_49808,N_49799);
and UO_221 (O_221,N_49996,N_49778);
nor UO_222 (O_222,N_49885,N_49823);
xnor UO_223 (O_223,N_49936,N_49835);
xor UO_224 (O_224,N_49970,N_49790);
and UO_225 (O_225,N_49789,N_49929);
and UO_226 (O_226,N_49786,N_49832);
xnor UO_227 (O_227,N_49958,N_49928);
nand UO_228 (O_228,N_49937,N_49917);
xor UO_229 (O_229,N_49883,N_49850);
nand UO_230 (O_230,N_49928,N_49874);
xnor UO_231 (O_231,N_49756,N_49957);
or UO_232 (O_232,N_49755,N_49821);
or UO_233 (O_233,N_49951,N_49861);
nor UO_234 (O_234,N_49776,N_49838);
xnor UO_235 (O_235,N_49963,N_49802);
or UO_236 (O_236,N_49764,N_49799);
or UO_237 (O_237,N_49872,N_49772);
and UO_238 (O_238,N_49898,N_49888);
and UO_239 (O_239,N_49903,N_49754);
nor UO_240 (O_240,N_49919,N_49975);
and UO_241 (O_241,N_49865,N_49806);
nor UO_242 (O_242,N_49760,N_49875);
xnor UO_243 (O_243,N_49758,N_49885);
nor UO_244 (O_244,N_49770,N_49750);
nand UO_245 (O_245,N_49986,N_49803);
nand UO_246 (O_246,N_49913,N_49862);
and UO_247 (O_247,N_49932,N_49965);
nor UO_248 (O_248,N_49842,N_49770);
and UO_249 (O_249,N_49950,N_49803);
nor UO_250 (O_250,N_49802,N_49977);
or UO_251 (O_251,N_49881,N_49895);
nand UO_252 (O_252,N_49809,N_49801);
nand UO_253 (O_253,N_49756,N_49797);
and UO_254 (O_254,N_49786,N_49804);
xnor UO_255 (O_255,N_49901,N_49973);
and UO_256 (O_256,N_49862,N_49877);
xnor UO_257 (O_257,N_49797,N_49870);
xor UO_258 (O_258,N_49795,N_49811);
nand UO_259 (O_259,N_49898,N_49983);
xor UO_260 (O_260,N_49890,N_49769);
or UO_261 (O_261,N_49756,N_49851);
or UO_262 (O_262,N_49913,N_49864);
or UO_263 (O_263,N_49894,N_49980);
xor UO_264 (O_264,N_49785,N_49969);
nand UO_265 (O_265,N_49819,N_49852);
xor UO_266 (O_266,N_49890,N_49841);
xor UO_267 (O_267,N_49995,N_49870);
or UO_268 (O_268,N_49829,N_49760);
and UO_269 (O_269,N_49895,N_49924);
or UO_270 (O_270,N_49931,N_49946);
nor UO_271 (O_271,N_49878,N_49965);
nand UO_272 (O_272,N_49963,N_49789);
and UO_273 (O_273,N_49856,N_49863);
nand UO_274 (O_274,N_49889,N_49766);
nor UO_275 (O_275,N_49858,N_49844);
or UO_276 (O_276,N_49850,N_49953);
or UO_277 (O_277,N_49803,N_49775);
nand UO_278 (O_278,N_49900,N_49887);
and UO_279 (O_279,N_49814,N_49883);
and UO_280 (O_280,N_49895,N_49979);
xnor UO_281 (O_281,N_49919,N_49933);
xor UO_282 (O_282,N_49928,N_49931);
or UO_283 (O_283,N_49759,N_49990);
or UO_284 (O_284,N_49964,N_49927);
xnor UO_285 (O_285,N_49935,N_49993);
nand UO_286 (O_286,N_49893,N_49813);
or UO_287 (O_287,N_49778,N_49799);
xnor UO_288 (O_288,N_49896,N_49867);
or UO_289 (O_289,N_49907,N_49846);
xor UO_290 (O_290,N_49993,N_49851);
nor UO_291 (O_291,N_49772,N_49775);
nand UO_292 (O_292,N_49888,N_49763);
nand UO_293 (O_293,N_49939,N_49891);
nor UO_294 (O_294,N_49766,N_49780);
nor UO_295 (O_295,N_49855,N_49830);
xnor UO_296 (O_296,N_49875,N_49779);
or UO_297 (O_297,N_49967,N_49807);
nor UO_298 (O_298,N_49979,N_49828);
xnor UO_299 (O_299,N_49840,N_49997);
nor UO_300 (O_300,N_49854,N_49837);
nor UO_301 (O_301,N_49982,N_49975);
xor UO_302 (O_302,N_49769,N_49976);
xor UO_303 (O_303,N_49757,N_49935);
or UO_304 (O_304,N_49816,N_49793);
and UO_305 (O_305,N_49870,N_49937);
xor UO_306 (O_306,N_49862,N_49972);
xor UO_307 (O_307,N_49903,N_49923);
and UO_308 (O_308,N_49751,N_49825);
or UO_309 (O_309,N_49872,N_49775);
nand UO_310 (O_310,N_49975,N_49786);
or UO_311 (O_311,N_49882,N_49941);
nor UO_312 (O_312,N_49793,N_49784);
nand UO_313 (O_313,N_49914,N_49974);
nor UO_314 (O_314,N_49764,N_49758);
nand UO_315 (O_315,N_49853,N_49929);
or UO_316 (O_316,N_49786,N_49867);
xor UO_317 (O_317,N_49894,N_49970);
or UO_318 (O_318,N_49783,N_49992);
nor UO_319 (O_319,N_49879,N_49954);
or UO_320 (O_320,N_49819,N_49751);
xor UO_321 (O_321,N_49780,N_49956);
nor UO_322 (O_322,N_49992,N_49836);
or UO_323 (O_323,N_49950,N_49764);
xnor UO_324 (O_324,N_49818,N_49936);
or UO_325 (O_325,N_49997,N_49770);
or UO_326 (O_326,N_49958,N_49975);
and UO_327 (O_327,N_49926,N_49953);
nand UO_328 (O_328,N_49913,N_49797);
and UO_329 (O_329,N_49989,N_49754);
nand UO_330 (O_330,N_49809,N_49920);
xor UO_331 (O_331,N_49801,N_49885);
xor UO_332 (O_332,N_49789,N_49881);
nand UO_333 (O_333,N_49763,N_49981);
or UO_334 (O_334,N_49932,N_49924);
nand UO_335 (O_335,N_49871,N_49960);
xor UO_336 (O_336,N_49843,N_49896);
or UO_337 (O_337,N_49775,N_49966);
nor UO_338 (O_338,N_49763,N_49953);
nor UO_339 (O_339,N_49934,N_49775);
or UO_340 (O_340,N_49819,N_49982);
nand UO_341 (O_341,N_49839,N_49910);
and UO_342 (O_342,N_49795,N_49958);
nor UO_343 (O_343,N_49947,N_49853);
nand UO_344 (O_344,N_49979,N_49921);
and UO_345 (O_345,N_49855,N_49937);
or UO_346 (O_346,N_49918,N_49942);
nor UO_347 (O_347,N_49871,N_49989);
and UO_348 (O_348,N_49989,N_49903);
nor UO_349 (O_349,N_49930,N_49899);
and UO_350 (O_350,N_49945,N_49950);
nand UO_351 (O_351,N_49775,N_49819);
and UO_352 (O_352,N_49995,N_49922);
or UO_353 (O_353,N_49994,N_49859);
xnor UO_354 (O_354,N_49794,N_49994);
and UO_355 (O_355,N_49831,N_49758);
nand UO_356 (O_356,N_49958,N_49919);
and UO_357 (O_357,N_49949,N_49920);
and UO_358 (O_358,N_49917,N_49909);
nor UO_359 (O_359,N_49983,N_49824);
nor UO_360 (O_360,N_49895,N_49874);
nor UO_361 (O_361,N_49988,N_49910);
and UO_362 (O_362,N_49939,N_49876);
nor UO_363 (O_363,N_49991,N_49756);
xor UO_364 (O_364,N_49801,N_49880);
or UO_365 (O_365,N_49986,N_49926);
or UO_366 (O_366,N_49881,N_49850);
nor UO_367 (O_367,N_49898,N_49877);
or UO_368 (O_368,N_49925,N_49831);
nand UO_369 (O_369,N_49827,N_49880);
nor UO_370 (O_370,N_49947,N_49804);
or UO_371 (O_371,N_49805,N_49820);
nor UO_372 (O_372,N_49798,N_49752);
and UO_373 (O_373,N_49859,N_49828);
nor UO_374 (O_374,N_49838,N_49906);
or UO_375 (O_375,N_49833,N_49962);
nand UO_376 (O_376,N_49965,N_49779);
nand UO_377 (O_377,N_49842,N_49909);
xor UO_378 (O_378,N_49970,N_49887);
nor UO_379 (O_379,N_49821,N_49815);
or UO_380 (O_380,N_49831,N_49935);
or UO_381 (O_381,N_49866,N_49951);
nor UO_382 (O_382,N_49957,N_49791);
and UO_383 (O_383,N_49782,N_49794);
and UO_384 (O_384,N_49961,N_49932);
nand UO_385 (O_385,N_49900,N_49877);
and UO_386 (O_386,N_49783,N_49920);
nand UO_387 (O_387,N_49893,N_49824);
or UO_388 (O_388,N_49860,N_49929);
nor UO_389 (O_389,N_49932,N_49989);
xor UO_390 (O_390,N_49934,N_49996);
and UO_391 (O_391,N_49949,N_49945);
nor UO_392 (O_392,N_49887,N_49863);
xnor UO_393 (O_393,N_49896,N_49816);
xnor UO_394 (O_394,N_49831,N_49791);
and UO_395 (O_395,N_49816,N_49760);
and UO_396 (O_396,N_49924,N_49879);
and UO_397 (O_397,N_49796,N_49790);
xor UO_398 (O_398,N_49955,N_49778);
nor UO_399 (O_399,N_49918,N_49832);
and UO_400 (O_400,N_49759,N_49769);
or UO_401 (O_401,N_49918,N_49888);
nand UO_402 (O_402,N_49762,N_49872);
nand UO_403 (O_403,N_49989,N_49941);
xor UO_404 (O_404,N_49892,N_49921);
xnor UO_405 (O_405,N_49860,N_49872);
and UO_406 (O_406,N_49875,N_49833);
or UO_407 (O_407,N_49981,N_49838);
and UO_408 (O_408,N_49779,N_49836);
xor UO_409 (O_409,N_49946,N_49923);
or UO_410 (O_410,N_49900,N_49917);
nor UO_411 (O_411,N_49917,N_49842);
or UO_412 (O_412,N_49803,N_49981);
or UO_413 (O_413,N_49784,N_49940);
nor UO_414 (O_414,N_49777,N_49937);
nand UO_415 (O_415,N_49882,N_49914);
and UO_416 (O_416,N_49807,N_49767);
or UO_417 (O_417,N_49987,N_49848);
or UO_418 (O_418,N_49936,N_49886);
or UO_419 (O_419,N_49904,N_49832);
nor UO_420 (O_420,N_49958,N_49790);
nor UO_421 (O_421,N_49768,N_49785);
nand UO_422 (O_422,N_49937,N_49795);
xor UO_423 (O_423,N_49981,N_49976);
and UO_424 (O_424,N_49820,N_49986);
xnor UO_425 (O_425,N_49997,N_49999);
or UO_426 (O_426,N_49819,N_49883);
nand UO_427 (O_427,N_49809,N_49909);
and UO_428 (O_428,N_49794,N_49751);
and UO_429 (O_429,N_49762,N_49975);
and UO_430 (O_430,N_49822,N_49826);
nor UO_431 (O_431,N_49777,N_49836);
and UO_432 (O_432,N_49855,N_49758);
nand UO_433 (O_433,N_49964,N_49948);
and UO_434 (O_434,N_49977,N_49989);
nand UO_435 (O_435,N_49971,N_49801);
nor UO_436 (O_436,N_49904,N_49861);
and UO_437 (O_437,N_49986,N_49874);
xnor UO_438 (O_438,N_49766,N_49868);
nand UO_439 (O_439,N_49765,N_49947);
or UO_440 (O_440,N_49901,N_49783);
nor UO_441 (O_441,N_49772,N_49855);
or UO_442 (O_442,N_49973,N_49862);
nor UO_443 (O_443,N_49861,N_49930);
and UO_444 (O_444,N_49943,N_49917);
and UO_445 (O_445,N_49981,N_49972);
nand UO_446 (O_446,N_49798,N_49992);
xor UO_447 (O_447,N_49784,N_49777);
and UO_448 (O_448,N_49792,N_49954);
and UO_449 (O_449,N_49945,N_49857);
nand UO_450 (O_450,N_49918,N_49987);
nor UO_451 (O_451,N_49832,N_49817);
or UO_452 (O_452,N_49955,N_49800);
xnor UO_453 (O_453,N_49982,N_49949);
nand UO_454 (O_454,N_49757,N_49872);
nor UO_455 (O_455,N_49808,N_49931);
nor UO_456 (O_456,N_49818,N_49916);
or UO_457 (O_457,N_49755,N_49751);
nor UO_458 (O_458,N_49893,N_49784);
nand UO_459 (O_459,N_49785,N_49860);
and UO_460 (O_460,N_49854,N_49874);
or UO_461 (O_461,N_49827,N_49873);
nand UO_462 (O_462,N_49860,N_49758);
nor UO_463 (O_463,N_49899,N_49761);
or UO_464 (O_464,N_49845,N_49892);
nand UO_465 (O_465,N_49844,N_49760);
and UO_466 (O_466,N_49912,N_49893);
and UO_467 (O_467,N_49900,N_49752);
nand UO_468 (O_468,N_49863,N_49790);
and UO_469 (O_469,N_49837,N_49916);
and UO_470 (O_470,N_49869,N_49867);
and UO_471 (O_471,N_49767,N_49756);
nand UO_472 (O_472,N_49867,N_49989);
and UO_473 (O_473,N_49914,N_49801);
nand UO_474 (O_474,N_49999,N_49756);
nor UO_475 (O_475,N_49937,N_49871);
or UO_476 (O_476,N_49780,N_49908);
or UO_477 (O_477,N_49814,N_49834);
nor UO_478 (O_478,N_49878,N_49810);
and UO_479 (O_479,N_49944,N_49827);
xor UO_480 (O_480,N_49987,N_49776);
nand UO_481 (O_481,N_49979,N_49865);
nor UO_482 (O_482,N_49976,N_49876);
nand UO_483 (O_483,N_49843,N_49930);
nor UO_484 (O_484,N_49905,N_49759);
and UO_485 (O_485,N_49983,N_49952);
xor UO_486 (O_486,N_49988,N_49814);
xnor UO_487 (O_487,N_49966,N_49924);
or UO_488 (O_488,N_49844,N_49987);
nor UO_489 (O_489,N_49878,N_49777);
xor UO_490 (O_490,N_49847,N_49935);
or UO_491 (O_491,N_49831,N_49795);
nand UO_492 (O_492,N_49859,N_49840);
or UO_493 (O_493,N_49905,N_49845);
xnor UO_494 (O_494,N_49804,N_49816);
xnor UO_495 (O_495,N_49755,N_49764);
xnor UO_496 (O_496,N_49841,N_49949);
or UO_497 (O_497,N_49968,N_49834);
nor UO_498 (O_498,N_49988,N_49842);
xnor UO_499 (O_499,N_49835,N_49942);
nor UO_500 (O_500,N_49873,N_49769);
and UO_501 (O_501,N_49791,N_49841);
nand UO_502 (O_502,N_49817,N_49988);
nor UO_503 (O_503,N_49985,N_49887);
or UO_504 (O_504,N_49834,N_49803);
and UO_505 (O_505,N_49755,N_49963);
or UO_506 (O_506,N_49839,N_49896);
nor UO_507 (O_507,N_49968,N_49928);
nand UO_508 (O_508,N_49855,N_49933);
nor UO_509 (O_509,N_49862,N_49897);
nor UO_510 (O_510,N_49971,N_49907);
nand UO_511 (O_511,N_49813,N_49967);
or UO_512 (O_512,N_49880,N_49814);
xnor UO_513 (O_513,N_49911,N_49985);
or UO_514 (O_514,N_49911,N_49926);
nor UO_515 (O_515,N_49888,N_49788);
or UO_516 (O_516,N_49885,N_49798);
xnor UO_517 (O_517,N_49956,N_49944);
or UO_518 (O_518,N_49795,N_49908);
xnor UO_519 (O_519,N_49752,N_49971);
or UO_520 (O_520,N_49845,N_49859);
nand UO_521 (O_521,N_49845,N_49984);
nor UO_522 (O_522,N_49788,N_49758);
or UO_523 (O_523,N_49901,N_49840);
or UO_524 (O_524,N_49876,N_49795);
and UO_525 (O_525,N_49946,N_49834);
xnor UO_526 (O_526,N_49959,N_49893);
nand UO_527 (O_527,N_49888,N_49912);
or UO_528 (O_528,N_49769,N_49799);
nor UO_529 (O_529,N_49838,N_49912);
nand UO_530 (O_530,N_49952,N_49771);
and UO_531 (O_531,N_49895,N_49996);
and UO_532 (O_532,N_49968,N_49906);
xnor UO_533 (O_533,N_49976,N_49823);
nor UO_534 (O_534,N_49948,N_49920);
nand UO_535 (O_535,N_49842,N_49875);
or UO_536 (O_536,N_49856,N_49852);
or UO_537 (O_537,N_49754,N_49938);
and UO_538 (O_538,N_49836,N_49959);
nor UO_539 (O_539,N_49777,N_49865);
or UO_540 (O_540,N_49765,N_49979);
xor UO_541 (O_541,N_49945,N_49855);
xor UO_542 (O_542,N_49955,N_49773);
and UO_543 (O_543,N_49982,N_49915);
xnor UO_544 (O_544,N_49986,N_49898);
xor UO_545 (O_545,N_49805,N_49953);
nor UO_546 (O_546,N_49799,N_49921);
nor UO_547 (O_547,N_49783,N_49770);
nor UO_548 (O_548,N_49821,N_49971);
and UO_549 (O_549,N_49949,N_49830);
nand UO_550 (O_550,N_49939,N_49894);
or UO_551 (O_551,N_49798,N_49952);
xnor UO_552 (O_552,N_49946,N_49832);
nor UO_553 (O_553,N_49949,N_49848);
nor UO_554 (O_554,N_49950,N_49918);
and UO_555 (O_555,N_49825,N_49904);
and UO_556 (O_556,N_49843,N_49956);
xnor UO_557 (O_557,N_49957,N_49865);
nand UO_558 (O_558,N_49952,N_49902);
xor UO_559 (O_559,N_49849,N_49989);
and UO_560 (O_560,N_49860,N_49918);
nor UO_561 (O_561,N_49977,N_49983);
xnor UO_562 (O_562,N_49916,N_49761);
nor UO_563 (O_563,N_49860,N_49951);
xnor UO_564 (O_564,N_49810,N_49850);
xor UO_565 (O_565,N_49937,N_49827);
nand UO_566 (O_566,N_49904,N_49796);
and UO_567 (O_567,N_49894,N_49794);
and UO_568 (O_568,N_49753,N_49776);
xor UO_569 (O_569,N_49929,N_49968);
or UO_570 (O_570,N_49977,N_49841);
xor UO_571 (O_571,N_49938,N_49928);
or UO_572 (O_572,N_49895,N_49819);
xnor UO_573 (O_573,N_49899,N_49842);
nand UO_574 (O_574,N_49893,N_49974);
or UO_575 (O_575,N_49850,N_49967);
xor UO_576 (O_576,N_49886,N_49867);
or UO_577 (O_577,N_49983,N_49825);
nor UO_578 (O_578,N_49912,N_49851);
and UO_579 (O_579,N_49888,N_49886);
xor UO_580 (O_580,N_49898,N_49914);
and UO_581 (O_581,N_49791,N_49856);
nand UO_582 (O_582,N_49826,N_49841);
nor UO_583 (O_583,N_49858,N_49814);
nor UO_584 (O_584,N_49779,N_49950);
xnor UO_585 (O_585,N_49932,N_49962);
or UO_586 (O_586,N_49909,N_49812);
nor UO_587 (O_587,N_49851,N_49821);
nor UO_588 (O_588,N_49859,N_49777);
nor UO_589 (O_589,N_49866,N_49920);
and UO_590 (O_590,N_49979,N_49776);
nand UO_591 (O_591,N_49860,N_49791);
and UO_592 (O_592,N_49928,N_49821);
and UO_593 (O_593,N_49911,N_49798);
xor UO_594 (O_594,N_49971,N_49776);
or UO_595 (O_595,N_49877,N_49971);
nand UO_596 (O_596,N_49786,N_49972);
xor UO_597 (O_597,N_49860,N_49934);
xnor UO_598 (O_598,N_49751,N_49980);
nor UO_599 (O_599,N_49975,N_49806);
nor UO_600 (O_600,N_49929,N_49827);
nor UO_601 (O_601,N_49982,N_49820);
and UO_602 (O_602,N_49946,N_49966);
xor UO_603 (O_603,N_49888,N_49943);
nand UO_604 (O_604,N_49982,N_49921);
xor UO_605 (O_605,N_49814,N_49974);
xnor UO_606 (O_606,N_49954,N_49828);
and UO_607 (O_607,N_49767,N_49860);
nor UO_608 (O_608,N_49847,N_49788);
and UO_609 (O_609,N_49969,N_49888);
and UO_610 (O_610,N_49755,N_49849);
nor UO_611 (O_611,N_49866,N_49789);
nor UO_612 (O_612,N_49915,N_49754);
or UO_613 (O_613,N_49943,N_49786);
nor UO_614 (O_614,N_49992,N_49841);
or UO_615 (O_615,N_49986,N_49943);
nand UO_616 (O_616,N_49933,N_49790);
nand UO_617 (O_617,N_49850,N_49806);
nand UO_618 (O_618,N_49878,N_49754);
xnor UO_619 (O_619,N_49874,N_49897);
nand UO_620 (O_620,N_49988,N_49981);
nor UO_621 (O_621,N_49886,N_49971);
xnor UO_622 (O_622,N_49767,N_49774);
nor UO_623 (O_623,N_49753,N_49836);
nand UO_624 (O_624,N_49979,N_49769);
nand UO_625 (O_625,N_49855,N_49910);
or UO_626 (O_626,N_49985,N_49952);
or UO_627 (O_627,N_49848,N_49854);
nor UO_628 (O_628,N_49975,N_49916);
nor UO_629 (O_629,N_49980,N_49793);
xor UO_630 (O_630,N_49773,N_49954);
or UO_631 (O_631,N_49871,N_49997);
and UO_632 (O_632,N_49816,N_49861);
and UO_633 (O_633,N_49772,N_49802);
or UO_634 (O_634,N_49854,N_49804);
nand UO_635 (O_635,N_49853,N_49801);
and UO_636 (O_636,N_49810,N_49830);
or UO_637 (O_637,N_49900,N_49834);
nor UO_638 (O_638,N_49855,N_49971);
and UO_639 (O_639,N_49951,N_49811);
or UO_640 (O_640,N_49902,N_49762);
nand UO_641 (O_641,N_49789,N_49900);
xor UO_642 (O_642,N_49771,N_49931);
xor UO_643 (O_643,N_49928,N_49981);
nor UO_644 (O_644,N_49889,N_49954);
nand UO_645 (O_645,N_49931,N_49836);
or UO_646 (O_646,N_49972,N_49971);
nand UO_647 (O_647,N_49950,N_49937);
xor UO_648 (O_648,N_49874,N_49954);
nand UO_649 (O_649,N_49847,N_49764);
and UO_650 (O_650,N_49900,N_49813);
nand UO_651 (O_651,N_49996,N_49891);
nand UO_652 (O_652,N_49758,N_49999);
or UO_653 (O_653,N_49855,N_49778);
and UO_654 (O_654,N_49965,N_49951);
and UO_655 (O_655,N_49931,N_49775);
nor UO_656 (O_656,N_49867,N_49774);
xnor UO_657 (O_657,N_49755,N_49844);
and UO_658 (O_658,N_49924,N_49878);
nor UO_659 (O_659,N_49875,N_49781);
or UO_660 (O_660,N_49769,N_49782);
or UO_661 (O_661,N_49945,N_49921);
nor UO_662 (O_662,N_49823,N_49967);
and UO_663 (O_663,N_49996,N_49765);
nand UO_664 (O_664,N_49818,N_49952);
nand UO_665 (O_665,N_49765,N_49942);
and UO_666 (O_666,N_49852,N_49861);
and UO_667 (O_667,N_49955,N_49766);
and UO_668 (O_668,N_49761,N_49839);
nor UO_669 (O_669,N_49907,N_49810);
xor UO_670 (O_670,N_49981,N_49758);
or UO_671 (O_671,N_49798,N_49777);
or UO_672 (O_672,N_49985,N_49895);
and UO_673 (O_673,N_49987,N_49771);
or UO_674 (O_674,N_49805,N_49767);
and UO_675 (O_675,N_49932,N_49796);
nand UO_676 (O_676,N_49855,N_49991);
and UO_677 (O_677,N_49911,N_49877);
xnor UO_678 (O_678,N_49865,N_49873);
nand UO_679 (O_679,N_49822,N_49789);
or UO_680 (O_680,N_49886,N_49943);
nand UO_681 (O_681,N_49932,N_49851);
and UO_682 (O_682,N_49846,N_49909);
or UO_683 (O_683,N_49806,N_49869);
nand UO_684 (O_684,N_49915,N_49909);
or UO_685 (O_685,N_49969,N_49896);
nand UO_686 (O_686,N_49797,N_49817);
or UO_687 (O_687,N_49774,N_49911);
or UO_688 (O_688,N_49958,N_49797);
or UO_689 (O_689,N_49778,N_49972);
nand UO_690 (O_690,N_49925,N_49930);
nor UO_691 (O_691,N_49876,N_49822);
or UO_692 (O_692,N_49832,N_49896);
nor UO_693 (O_693,N_49771,N_49917);
xnor UO_694 (O_694,N_49959,N_49857);
nand UO_695 (O_695,N_49756,N_49985);
and UO_696 (O_696,N_49944,N_49873);
and UO_697 (O_697,N_49767,N_49968);
nand UO_698 (O_698,N_49928,N_49952);
nor UO_699 (O_699,N_49807,N_49834);
nand UO_700 (O_700,N_49913,N_49960);
xor UO_701 (O_701,N_49902,N_49820);
nor UO_702 (O_702,N_49984,N_49964);
nor UO_703 (O_703,N_49835,N_49995);
nor UO_704 (O_704,N_49849,N_49917);
nor UO_705 (O_705,N_49965,N_49804);
xnor UO_706 (O_706,N_49867,N_49828);
or UO_707 (O_707,N_49923,N_49763);
or UO_708 (O_708,N_49938,N_49870);
and UO_709 (O_709,N_49858,N_49888);
nor UO_710 (O_710,N_49761,N_49966);
or UO_711 (O_711,N_49825,N_49830);
nand UO_712 (O_712,N_49879,N_49893);
xnor UO_713 (O_713,N_49871,N_49841);
or UO_714 (O_714,N_49950,N_49978);
and UO_715 (O_715,N_49805,N_49868);
xor UO_716 (O_716,N_49895,N_49997);
or UO_717 (O_717,N_49862,N_49984);
nand UO_718 (O_718,N_49753,N_49811);
nand UO_719 (O_719,N_49827,N_49804);
xnor UO_720 (O_720,N_49853,N_49831);
xor UO_721 (O_721,N_49755,N_49991);
nand UO_722 (O_722,N_49750,N_49811);
xor UO_723 (O_723,N_49961,N_49995);
nor UO_724 (O_724,N_49783,N_49790);
and UO_725 (O_725,N_49942,N_49842);
nand UO_726 (O_726,N_49783,N_49912);
and UO_727 (O_727,N_49773,N_49799);
nand UO_728 (O_728,N_49923,N_49920);
and UO_729 (O_729,N_49951,N_49979);
xnor UO_730 (O_730,N_49794,N_49901);
xnor UO_731 (O_731,N_49892,N_49818);
nor UO_732 (O_732,N_49889,N_49883);
and UO_733 (O_733,N_49812,N_49938);
xor UO_734 (O_734,N_49932,N_49983);
nand UO_735 (O_735,N_49870,N_49916);
nand UO_736 (O_736,N_49786,N_49770);
nor UO_737 (O_737,N_49963,N_49974);
or UO_738 (O_738,N_49985,N_49928);
nand UO_739 (O_739,N_49947,N_49771);
or UO_740 (O_740,N_49784,N_49832);
and UO_741 (O_741,N_49753,N_49825);
and UO_742 (O_742,N_49892,N_49900);
xor UO_743 (O_743,N_49880,N_49993);
xor UO_744 (O_744,N_49936,N_49856);
and UO_745 (O_745,N_49961,N_49830);
xor UO_746 (O_746,N_49850,N_49815);
xor UO_747 (O_747,N_49908,N_49970);
and UO_748 (O_748,N_49920,N_49970);
or UO_749 (O_749,N_49784,N_49802);
or UO_750 (O_750,N_49889,N_49921);
nor UO_751 (O_751,N_49919,N_49896);
nor UO_752 (O_752,N_49901,N_49827);
or UO_753 (O_753,N_49837,N_49901);
xor UO_754 (O_754,N_49798,N_49868);
nor UO_755 (O_755,N_49945,N_49880);
nor UO_756 (O_756,N_49895,N_49757);
xor UO_757 (O_757,N_49949,N_49875);
nor UO_758 (O_758,N_49926,N_49780);
nor UO_759 (O_759,N_49890,N_49812);
or UO_760 (O_760,N_49823,N_49865);
xor UO_761 (O_761,N_49759,N_49832);
xor UO_762 (O_762,N_49906,N_49788);
and UO_763 (O_763,N_49915,N_49817);
and UO_764 (O_764,N_49999,N_49896);
nand UO_765 (O_765,N_49966,N_49753);
and UO_766 (O_766,N_49853,N_49896);
or UO_767 (O_767,N_49974,N_49826);
or UO_768 (O_768,N_49818,N_49944);
nor UO_769 (O_769,N_49824,N_49827);
nor UO_770 (O_770,N_49832,N_49801);
nor UO_771 (O_771,N_49951,N_49908);
and UO_772 (O_772,N_49963,N_49999);
xnor UO_773 (O_773,N_49879,N_49982);
nor UO_774 (O_774,N_49820,N_49949);
nand UO_775 (O_775,N_49987,N_49857);
nand UO_776 (O_776,N_49946,N_49890);
and UO_777 (O_777,N_49998,N_49901);
nor UO_778 (O_778,N_49831,N_49834);
xnor UO_779 (O_779,N_49982,N_49940);
xnor UO_780 (O_780,N_49846,N_49764);
or UO_781 (O_781,N_49948,N_49808);
and UO_782 (O_782,N_49968,N_49829);
nor UO_783 (O_783,N_49822,N_49982);
xnor UO_784 (O_784,N_49891,N_49908);
nor UO_785 (O_785,N_49965,N_49985);
and UO_786 (O_786,N_49860,N_49777);
or UO_787 (O_787,N_49931,N_49823);
and UO_788 (O_788,N_49907,N_49838);
and UO_789 (O_789,N_49879,N_49813);
or UO_790 (O_790,N_49759,N_49992);
nor UO_791 (O_791,N_49994,N_49873);
nor UO_792 (O_792,N_49755,N_49763);
and UO_793 (O_793,N_49758,N_49817);
and UO_794 (O_794,N_49791,N_49986);
and UO_795 (O_795,N_49911,N_49890);
xnor UO_796 (O_796,N_49886,N_49952);
nand UO_797 (O_797,N_49823,N_49872);
nand UO_798 (O_798,N_49765,N_49928);
or UO_799 (O_799,N_49931,N_49839);
nor UO_800 (O_800,N_49857,N_49819);
and UO_801 (O_801,N_49757,N_49773);
and UO_802 (O_802,N_49811,N_49948);
nand UO_803 (O_803,N_49754,N_49769);
xnor UO_804 (O_804,N_49991,N_49913);
or UO_805 (O_805,N_49887,N_49936);
and UO_806 (O_806,N_49837,N_49872);
or UO_807 (O_807,N_49904,N_49995);
xnor UO_808 (O_808,N_49770,N_49785);
and UO_809 (O_809,N_49792,N_49822);
and UO_810 (O_810,N_49765,N_49935);
xor UO_811 (O_811,N_49999,N_49903);
nor UO_812 (O_812,N_49833,N_49848);
or UO_813 (O_813,N_49774,N_49765);
nor UO_814 (O_814,N_49810,N_49759);
xor UO_815 (O_815,N_49810,N_49936);
nor UO_816 (O_816,N_49811,N_49812);
or UO_817 (O_817,N_49941,N_49943);
xnor UO_818 (O_818,N_49899,N_49939);
or UO_819 (O_819,N_49826,N_49917);
nand UO_820 (O_820,N_49979,N_49919);
nor UO_821 (O_821,N_49829,N_49962);
xor UO_822 (O_822,N_49768,N_49826);
xor UO_823 (O_823,N_49985,N_49862);
or UO_824 (O_824,N_49922,N_49777);
or UO_825 (O_825,N_49940,N_49873);
or UO_826 (O_826,N_49985,N_49960);
xor UO_827 (O_827,N_49823,N_49832);
nand UO_828 (O_828,N_49950,N_49781);
nand UO_829 (O_829,N_49836,N_49801);
or UO_830 (O_830,N_49985,N_49864);
or UO_831 (O_831,N_49998,N_49916);
and UO_832 (O_832,N_49814,N_49825);
nand UO_833 (O_833,N_49759,N_49825);
nand UO_834 (O_834,N_49910,N_49786);
xnor UO_835 (O_835,N_49967,N_49952);
xor UO_836 (O_836,N_49901,N_49957);
xor UO_837 (O_837,N_49857,N_49790);
and UO_838 (O_838,N_49782,N_49889);
or UO_839 (O_839,N_49917,N_49887);
xor UO_840 (O_840,N_49948,N_49861);
nand UO_841 (O_841,N_49754,N_49950);
xnor UO_842 (O_842,N_49867,N_49999);
or UO_843 (O_843,N_49881,N_49892);
nor UO_844 (O_844,N_49766,N_49975);
nand UO_845 (O_845,N_49882,N_49844);
xor UO_846 (O_846,N_49890,N_49916);
xor UO_847 (O_847,N_49946,N_49952);
or UO_848 (O_848,N_49877,N_49856);
xnor UO_849 (O_849,N_49954,N_49933);
nor UO_850 (O_850,N_49824,N_49840);
nand UO_851 (O_851,N_49931,N_49826);
or UO_852 (O_852,N_49818,N_49799);
nand UO_853 (O_853,N_49926,N_49979);
or UO_854 (O_854,N_49798,N_49815);
xor UO_855 (O_855,N_49946,N_49915);
and UO_856 (O_856,N_49976,N_49808);
nand UO_857 (O_857,N_49833,N_49759);
or UO_858 (O_858,N_49887,N_49785);
or UO_859 (O_859,N_49987,N_49975);
nor UO_860 (O_860,N_49859,N_49957);
xor UO_861 (O_861,N_49811,N_49808);
nand UO_862 (O_862,N_49806,N_49961);
and UO_863 (O_863,N_49877,N_49876);
or UO_864 (O_864,N_49816,N_49966);
xnor UO_865 (O_865,N_49884,N_49909);
nand UO_866 (O_866,N_49945,N_49834);
nor UO_867 (O_867,N_49756,N_49990);
or UO_868 (O_868,N_49767,N_49804);
and UO_869 (O_869,N_49779,N_49831);
nand UO_870 (O_870,N_49914,N_49932);
and UO_871 (O_871,N_49988,N_49885);
nand UO_872 (O_872,N_49800,N_49958);
and UO_873 (O_873,N_49814,N_49756);
nor UO_874 (O_874,N_49858,N_49949);
and UO_875 (O_875,N_49914,N_49873);
or UO_876 (O_876,N_49904,N_49953);
nand UO_877 (O_877,N_49815,N_49948);
nand UO_878 (O_878,N_49875,N_49754);
or UO_879 (O_879,N_49854,N_49931);
or UO_880 (O_880,N_49807,N_49830);
xor UO_881 (O_881,N_49825,N_49750);
or UO_882 (O_882,N_49874,N_49801);
and UO_883 (O_883,N_49825,N_49967);
nor UO_884 (O_884,N_49833,N_49859);
and UO_885 (O_885,N_49863,N_49899);
or UO_886 (O_886,N_49846,N_49833);
xnor UO_887 (O_887,N_49808,N_49982);
or UO_888 (O_888,N_49823,N_49760);
or UO_889 (O_889,N_49754,N_49986);
and UO_890 (O_890,N_49959,N_49938);
and UO_891 (O_891,N_49868,N_49942);
xnor UO_892 (O_892,N_49930,N_49890);
nor UO_893 (O_893,N_49861,N_49854);
nand UO_894 (O_894,N_49863,N_49905);
nand UO_895 (O_895,N_49870,N_49889);
xnor UO_896 (O_896,N_49811,N_49761);
and UO_897 (O_897,N_49827,N_49956);
nand UO_898 (O_898,N_49997,N_49964);
and UO_899 (O_899,N_49876,N_49919);
nand UO_900 (O_900,N_49992,N_49772);
xor UO_901 (O_901,N_49952,N_49941);
nor UO_902 (O_902,N_49894,N_49889);
nor UO_903 (O_903,N_49986,N_49952);
nand UO_904 (O_904,N_49951,N_49851);
and UO_905 (O_905,N_49950,N_49793);
or UO_906 (O_906,N_49852,N_49871);
and UO_907 (O_907,N_49833,N_49807);
nand UO_908 (O_908,N_49815,N_49845);
nand UO_909 (O_909,N_49876,N_49967);
and UO_910 (O_910,N_49819,N_49877);
xor UO_911 (O_911,N_49850,N_49931);
xnor UO_912 (O_912,N_49990,N_49903);
xor UO_913 (O_913,N_49805,N_49943);
nand UO_914 (O_914,N_49768,N_49990);
nand UO_915 (O_915,N_49820,N_49930);
nor UO_916 (O_916,N_49923,N_49853);
and UO_917 (O_917,N_49882,N_49996);
or UO_918 (O_918,N_49837,N_49911);
and UO_919 (O_919,N_49760,N_49872);
and UO_920 (O_920,N_49756,N_49914);
xor UO_921 (O_921,N_49936,N_49864);
nor UO_922 (O_922,N_49862,N_49986);
and UO_923 (O_923,N_49817,N_49913);
nor UO_924 (O_924,N_49811,N_49833);
or UO_925 (O_925,N_49943,N_49818);
or UO_926 (O_926,N_49994,N_49838);
or UO_927 (O_927,N_49939,N_49834);
nand UO_928 (O_928,N_49818,N_49917);
nor UO_929 (O_929,N_49864,N_49901);
and UO_930 (O_930,N_49960,N_49945);
nor UO_931 (O_931,N_49858,N_49778);
xnor UO_932 (O_932,N_49819,N_49755);
and UO_933 (O_933,N_49751,N_49848);
or UO_934 (O_934,N_49911,N_49874);
and UO_935 (O_935,N_49976,N_49877);
nor UO_936 (O_936,N_49898,N_49948);
xor UO_937 (O_937,N_49846,N_49883);
and UO_938 (O_938,N_49854,N_49869);
xor UO_939 (O_939,N_49827,N_49890);
and UO_940 (O_940,N_49973,N_49896);
and UO_941 (O_941,N_49967,N_49884);
or UO_942 (O_942,N_49845,N_49991);
nand UO_943 (O_943,N_49815,N_49917);
nand UO_944 (O_944,N_49781,N_49753);
and UO_945 (O_945,N_49998,N_49807);
nor UO_946 (O_946,N_49953,N_49892);
or UO_947 (O_947,N_49829,N_49753);
xnor UO_948 (O_948,N_49847,N_49941);
and UO_949 (O_949,N_49832,N_49902);
nor UO_950 (O_950,N_49898,N_49922);
xor UO_951 (O_951,N_49965,N_49976);
nand UO_952 (O_952,N_49835,N_49869);
nor UO_953 (O_953,N_49905,N_49880);
and UO_954 (O_954,N_49866,N_49942);
or UO_955 (O_955,N_49996,N_49989);
and UO_956 (O_956,N_49971,N_49795);
nand UO_957 (O_957,N_49804,N_49985);
xor UO_958 (O_958,N_49878,N_49999);
or UO_959 (O_959,N_49837,N_49789);
and UO_960 (O_960,N_49757,N_49986);
nand UO_961 (O_961,N_49952,N_49989);
and UO_962 (O_962,N_49841,N_49779);
and UO_963 (O_963,N_49978,N_49985);
xor UO_964 (O_964,N_49801,N_49843);
nor UO_965 (O_965,N_49991,N_49771);
and UO_966 (O_966,N_49781,N_49834);
nand UO_967 (O_967,N_49805,N_49814);
xor UO_968 (O_968,N_49984,N_49981);
and UO_969 (O_969,N_49789,N_49760);
and UO_970 (O_970,N_49778,N_49790);
or UO_971 (O_971,N_49977,N_49771);
or UO_972 (O_972,N_49861,N_49870);
or UO_973 (O_973,N_49830,N_49782);
nor UO_974 (O_974,N_49873,N_49850);
nand UO_975 (O_975,N_49763,N_49972);
or UO_976 (O_976,N_49857,N_49876);
nand UO_977 (O_977,N_49792,N_49843);
and UO_978 (O_978,N_49969,N_49901);
nand UO_979 (O_979,N_49755,N_49951);
or UO_980 (O_980,N_49995,N_49958);
nor UO_981 (O_981,N_49864,N_49949);
nand UO_982 (O_982,N_49798,N_49849);
nand UO_983 (O_983,N_49945,N_49810);
nor UO_984 (O_984,N_49925,N_49963);
xor UO_985 (O_985,N_49961,N_49753);
or UO_986 (O_986,N_49967,N_49913);
and UO_987 (O_987,N_49990,N_49875);
nand UO_988 (O_988,N_49925,N_49759);
nand UO_989 (O_989,N_49770,N_49752);
nand UO_990 (O_990,N_49751,N_49875);
nor UO_991 (O_991,N_49962,N_49775);
or UO_992 (O_992,N_49886,N_49973);
and UO_993 (O_993,N_49814,N_49911);
and UO_994 (O_994,N_49974,N_49947);
and UO_995 (O_995,N_49760,N_49801);
nand UO_996 (O_996,N_49791,N_49995);
nand UO_997 (O_997,N_49936,N_49770);
nor UO_998 (O_998,N_49917,N_49964);
nand UO_999 (O_999,N_49795,N_49885);
nor UO_1000 (O_1000,N_49994,N_49829);
nand UO_1001 (O_1001,N_49991,N_49762);
and UO_1002 (O_1002,N_49904,N_49967);
nand UO_1003 (O_1003,N_49954,N_49953);
nor UO_1004 (O_1004,N_49911,N_49941);
nand UO_1005 (O_1005,N_49879,N_49899);
nand UO_1006 (O_1006,N_49771,N_49839);
nand UO_1007 (O_1007,N_49934,N_49867);
nor UO_1008 (O_1008,N_49981,N_49805);
xor UO_1009 (O_1009,N_49963,N_49870);
or UO_1010 (O_1010,N_49897,N_49969);
xor UO_1011 (O_1011,N_49845,N_49939);
xnor UO_1012 (O_1012,N_49892,N_49860);
or UO_1013 (O_1013,N_49986,N_49821);
nor UO_1014 (O_1014,N_49879,N_49754);
and UO_1015 (O_1015,N_49954,N_49806);
or UO_1016 (O_1016,N_49756,N_49951);
xnor UO_1017 (O_1017,N_49826,N_49776);
xnor UO_1018 (O_1018,N_49869,N_49845);
nand UO_1019 (O_1019,N_49864,N_49890);
or UO_1020 (O_1020,N_49886,N_49920);
xnor UO_1021 (O_1021,N_49932,N_49927);
xnor UO_1022 (O_1022,N_49997,N_49767);
nand UO_1023 (O_1023,N_49954,N_49947);
or UO_1024 (O_1024,N_49989,N_49906);
or UO_1025 (O_1025,N_49990,N_49978);
nor UO_1026 (O_1026,N_49777,N_49997);
nand UO_1027 (O_1027,N_49984,N_49789);
nor UO_1028 (O_1028,N_49845,N_49782);
nor UO_1029 (O_1029,N_49852,N_49837);
or UO_1030 (O_1030,N_49933,N_49899);
and UO_1031 (O_1031,N_49839,N_49810);
or UO_1032 (O_1032,N_49931,N_49991);
and UO_1033 (O_1033,N_49947,N_49884);
or UO_1034 (O_1034,N_49805,N_49756);
xor UO_1035 (O_1035,N_49895,N_49910);
and UO_1036 (O_1036,N_49765,N_49908);
xor UO_1037 (O_1037,N_49861,N_49968);
or UO_1038 (O_1038,N_49753,N_49998);
xnor UO_1039 (O_1039,N_49968,N_49787);
xor UO_1040 (O_1040,N_49793,N_49908);
or UO_1041 (O_1041,N_49992,N_49880);
xor UO_1042 (O_1042,N_49753,N_49895);
or UO_1043 (O_1043,N_49969,N_49780);
xnor UO_1044 (O_1044,N_49937,N_49820);
nor UO_1045 (O_1045,N_49994,N_49768);
or UO_1046 (O_1046,N_49966,N_49991);
or UO_1047 (O_1047,N_49871,N_49750);
nand UO_1048 (O_1048,N_49798,N_49847);
nor UO_1049 (O_1049,N_49918,N_49993);
or UO_1050 (O_1050,N_49882,N_49988);
nor UO_1051 (O_1051,N_49834,N_49855);
or UO_1052 (O_1052,N_49979,N_49846);
xnor UO_1053 (O_1053,N_49848,N_49919);
nand UO_1054 (O_1054,N_49842,N_49934);
or UO_1055 (O_1055,N_49885,N_49814);
and UO_1056 (O_1056,N_49792,N_49983);
xor UO_1057 (O_1057,N_49856,N_49805);
nand UO_1058 (O_1058,N_49822,N_49867);
nand UO_1059 (O_1059,N_49896,N_49796);
or UO_1060 (O_1060,N_49963,N_49763);
nand UO_1061 (O_1061,N_49943,N_49821);
nand UO_1062 (O_1062,N_49934,N_49801);
xor UO_1063 (O_1063,N_49754,N_49810);
nand UO_1064 (O_1064,N_49885,N_49919);
xnor UO_1065 (O_1065,N_49969,N_49861);
and UO_1066 (O_1066,N_49797,N_49981);
and UO_1067 (O_1067,N_49826,N_49785);
nand UO_1068 (O_1068,N_49839,N_49792);
nand UO_1069 (O_1069,N_49948,N_49872);
and UO_1070 (O_1070,N_49947,N_49887);
and UO_1071 (O_1071,N_49985,N_49816);
nand UO_1072 (O_1072,N_49843,N_49882);
nor UO_1073 (O_1073,N_49938,N_49996);
and UO_1074 (O_1074,N_49912,N_49827);
and UO_1075 (O_1075,N_49967,N_49985);
xnor UO_1076 (O_1076,N_49965,N_49841);
or UO_1077 (O_1077,N_49942,N_49890);
and UO_1078 (O_1078,N_49966,N_49882);
nand UO_1079 (O_1079,N_49782,N_49777);
nand UO_1080 (O_1080,N_49790,N_49832);
or UO_1081 (O_1081,N_49807,N_49763);
nand UO_1082 (O_1082,N_49847,N_49971);
nor UO_1083 (O_1083,N_49926,N_49821);
xnor UO_1084 (O_1084,N_49944,N_49926);
nand UO_1085 (O_1085,N_49858,N_49953);
xor UO_1086 (O_1086,N_49894,N_49961);
xnor UO_1087 (O_1087,N_49866,N_49896);
and UO_1088 (O_1088,N_49809,N_49967);
xnor UO_1089 (O_1089,N_49871,N_49847);
nand UO_1090 (O_1090,N_49773,N_49892);
or UO_1091 (O_1091,N_49854,N_49983);
nor UO_1092 (O_1092,N_49775,N_49906);
nand UO_1093 (O_1093,N_49841,N_49830);
or UO_1094 (O_1094,N_49816,N_49939);
and UO_1095 (O_1095,N_49801,N_49795);
or UO_1096 (O_1096,N_49941,N_49948);
nand UO_1097 (O_1097,N_49803,N_49990);
xor UO_1098 (O_1098,N_49986,N_49776);
xor UO_1099 (O_1099,N_49815,N_49753);
xnor UO_1100 (O_1100,N_49855,N_49890);
and UO_1101 (O_1101,N_49844,N_49968);
nor UO_1102 (O_1102,N_49885,N_49773);
nor UO_1103 (O_1103,N_49979,N_49958);
xnor UO_1104 (O_1104,N_49975,N_49951);
xnor UO_1105 (O_1105,N_49866,N_49755);
and UO_1106 (O_1106,N_49832,N_49752);
and UO_1107 (O_1107,N_49903,N_49956);
nand UO_1108 (O_1108,N_49999,N_49938);
nor UO_1109 (O_1109,N_49850,N_49855);
nand UO_1110 (O_1110,N_49874,N_49991);
nand UO_1111 (O_1111,N_49855,N_49818);
nor UO_1112 (O_1112,N_49872,N_49843);
nor UO_1113 (O_1113,N_49800,N_49828);
or UO_1114 (O_1114,N_49908,N_49986);
and UO_1115 (O_1115,N_49995,N_49948);
nor UO_1116 (O_1116,N_49960,N_49815);
xor UO_1117 (O_1117,N_49901,N_49939);
xnor UO_1118 (O_1118,N_49797,N_49811);
and UO_1119 (O_1119,N_49785,N_49893);
xor UO_1120 (O_1120,N_49849,N_49954);
nand UO_1121 (O_1121,N_49946,N_49857);
nor UO_1122 (O_1122,N_49793,N_49806);
or UO_1123 (O_1123,N_49944,N_49964);
nand UO_1124 (O_1124,N_49868,N_49862);
nand UO_1125 (O_1125,N_49762,N_49971);
nand UO_1126 (O_1126,N_49869,N_49945);
xor UO_1127 (O_1127,N_49809,N_49959);
nand UO_1128 (O_1128,N_49880,N_49799);
xor UO_1129 (O_1129,N_49901,N_49759);
and UO_1130 (O_1130,N_49846,N_49752);
nor UO_1131 (O_1131,N_49750,N_49880);
nor UO_1132 (O_1132,N_49819,N_49886);
or UO_1133 (O_1133,N_49829,N_49886);
or UO_1134 (O_1134,N_49912,N_49808);
and UO_1135 (O_1135,N_49974,N_49902);
nor UO_1136 (O_1136,N_49801,N_49864);
nand UO_1137 (O_1137,N_49961,N_49756);
nand UO_1138 (O_1138,N_49992,N_49820);
nand UO_1139 (O_1139,N_49912,N_49786);
nor UO_1140 (O_1140,N_49975,N_49873);
xnor UO_1141 (O_1141,N_49786,N_49956);
and UO_1142 (O_1142,N_49908,N_49853);
xnor UO_1143 (O_1143,N_49750,N_49991);
and UO_1144 (O_1144,N_49807,N_49916);
or UO_1145 (O_1145,N_49899,N_49759);
xor UO_1146 (O_1146,N_49971,N_49783);
and UO_1147 (O_1147,N_49800,N_49949);
xnor UO_1148 (O_1148,N_49766,N_49895);
and UO_1149 (O_1149,N_49927,N_49844);
nand UO_1150 (O_1150,N_49787,N_49935);
nand UO_1151 (O_1151,N_49902,N_49949);
nor UO_1152 (O_1152,N_49772,N_49991);
xnor UO_1153 (O_1153,N_49791,N_49938);
nor UO_1154 (O_1154,N_49815,N_49968);
xor UO_1155 (O_1155,N_49793,N_49966);
and UO_1156 (O_1156,N_49837,N_49937);
and UO_1157 (O_1157,N_49952,N_49760);
nor UO_1158 (O_1158,N_49989,N_49803);
xor UO_1159 (O_1159,N_49965,N_49894);
or UO_1160 (O_1160,N_49851,N_49766);
nand UO_1161 (O_1161,N_49803,N_49959);
nor UO_1162 (O_1162,N_49769,N_49929);
or UO_1163 (O_1163,N_49987,N_49894);
xor UO_1164 (O_1164,N_49795,N_49753);
nor UO_1165 (O_1165,N_49834,N_49884);
xnor UO_1166 (O_1166,N_49911,N_49853);
nor UO_1167 (O_1167,N_49804,N_49848);
or UO_1168 (O_1168,N_49751,N_49869);
xor UO_1169 (O_1169,N_49931,N_49971);
xor UO_1170 (O_1170,N_49976,N_49778);
or UO_1171 (O_1171,N_49815,N_49944);
nor UO_1172 (O_1172,N_49785,N_49922);
nor UO_1173 (O_1173,N_49849,N_49766);
or UO_1174 (O_1174,N_49821,N_49871);
or UO_1175 (O_1175,N_49995,N_49822);
or UO_1176 (O_1176,N_49797,N_49764);
nor UO_1177 (O_1177,N_49971,N_49925);
and UO_1178 (O_1178,N_49778,N_49863);
nor UO_1179 (O_1179,N_49765,N_49815);
nand UO_1180 (O_1180,N_49902,N_49816);
and UO_1181 (O_1181,N_49995,N_49801);
or UO_1182 (O_1182,N_49999,N_49875);
nand UO_1183 (O_1183,N_49881,N_49917);
nand UO_1184 (O_1184,N_49957,N_49928);
and UO_1185 (O_1185,N_49818,N_49891);
and UO_1186 (O_1186,N_49815,N_49807);
and UO_1187 (O_1187,N_49840,N_49962);
nand UO_1188 (O_1188,N_49787,N_49896);
or UO_1189 (O_1189,N_49951,N_49750);
xor UO_1190 (O_1190,N_49988,N_49881);
or UO_1191 (O_1191,N_49808,N_49756);
nor UO_1192 (O_1192,N_49898,N_49864);
and UO_1193 (O_1193,N_49868,N_49763);
nand UO_1194 (O_1194,N_49882,N_49875);
nor UO_1195 (O_1195,N_49762,N_49915);
or UO_1196 (O_1196,N_49774,N_49957);
nor UO_1197 (O_1197,N_49802,N_49781);
or UO_1198 (O_1198,N_49884,N_49958);
nor UO_1199 (O_1199,N_49789,N_49928);
xnor UO_1200 (O_1200,N_49839,N_49770);
nand UO_1201 (O_1201,N_49815,N_49950);
and UO_1202 (O_1202,N_49884,N_49811);
or UO_1203 (O_1203,N_49841,N_49788);
and UO_1204 (O_1204,N_49998,N_49759);
and UO_1205 (O_1205,N_49790,N_49794);
nand UO_1206 (O_1206,N_49758,N_49770);
nand UO_1207 (O_1207,N_49871,N_49756);
nor UO_1208 (O_1208,N_49896,N_49886);
or UO_1209 (O_1209,N_49894,N_49923);
nand UO_1210 (O_1210,N_49803,N_49976);
or UO_1211 (O_1211,N_49942,N_49818);
nor UO_1212 (O_1212,N_49841,N_49799);
xnor UO_1213 (O_1213,N_49927,N_49808);
nor UO_1214 (O_1214,N_49848,N_49766);
xnor UO_1215 (O_1215,N_49941,N_49908);
nor UO_1216 (O_1216,N_49836,N_49803);
or UO_1217 (O_1217,N_49792,N_49860);
xnor UO_1218 (O_1218,N_49814,N_49824);
or UO_1219 (O_1219,N_49891,N_49782);
xor UO_1220 (O_1220,N_49779,N_49894);
or UO_1221 (O_1221,N_49864,N_49802);
nor UO_1222 (O_1222,N_49870,N_49909);
nor UO_1223 (O_1223,N_49793,N_49826);
and UO_1224 (O_1224,N_49773,N_49818);
and UO_1225 (O_1225,N_49883,N_49822);
nor UO_1226 (O_1226,N_49762,N_49752);
nor UO_1227 (O_1227,N_49929,N_49783);
nand UO_1228 (O_1228,N_49925,N_49797);
xor UO_1229 (O_1229,N_49920,N_49841);
nand UO_1230 (O_1230,N_49809,N_49972);
xor UO_1231 (O_1231,N_49850,N_49926);
xor UO_1232 (O_1232,N_49968,N_49893);
nand UO_1233 (O_1233,N_49975,N_49805);
or UO_1234 (O_1234,N_49765,N_49758);
nor UO_1235 (O_1235,N_49912,N_49750);
or UO_1236 (O_1236,N_49785,N_49866);
and UO_1237 (O_1237,N_49892,N_49814);
and UO_1238 (O_1238,N_49971,N_49913);
and UO_1239 (O_1239,N_49955,N_49868);
or UO_1240 (O_1240,N_49967,N_49976);
and UO_1241 (O_1241,N_49892,N_49771);
or UO_1242 (O_1242,N_49827,N_49759);
xnor UO_1243 (O_1243,N_49811,N_49777);
and UO_1244 (O_1244,N_49969,N_49970);
xnor UO_1245 (O_1245,N_49909,N_49811);
or UO_1246 (O_1246,N_49960,N_49899);
xnor UO_1247 (O_1247,N_49876,N_49812);
or UO_1248 (O_1248,N_49828,N_49909);
xnor UO_1249 (O_1249,N_49864,N_49803);
nand UO_1250 (O_1250,N_49937,N_49766);
and UO_1251 (O_1251,N_49953,N_49798);
xnor UO_1252 (O_1252,N_49856,N_49923);
or UO_1253 (O_1253,N_49940,N_49760);
and UO_1254 (O_1254,N_49796,N_49894);
xor UO_1255 (O_1255,N_49772,N_49833);
nand UO_1256 (O_1256,N_49961,N_49941);
xnor UO_1257 (O_1257,N_49952,N_49906);
and UO_1258 (O_1258,N_49967,N_49773);
or UO_1259 (O_1259,N_49892,N_49919);
and UO_1260 (O_1260,N_49965,N_49962);
xnor UO_1261 (O_1261,N_49981,N_49902);
or UO_1262 (O_1262,N_49887,N_49855);
and UO_1263 (O_1263,N_49893,N_49850);
nand UO_1264 (O_1264,N_49897,N_49844);
nor UO_1265 (O_1265,N_49834,N_49955);
or UO_1266 (O_1266,N_49904,N_49838);
or UO_1267 (O_1267,N_49785,N_49952);
or UO_1268 (O_1268,N_49789,N_49869);
nor UO_1269 (O_1269,N_49792,N_49977);
nand UO_1270 (O_1270,N_49791,N_49976);
or UO_1271 (O_1271,N_49934,N_49800);
nand UO_1272 (O_1272,N_49967,N_49790);
nor UO_1273 (O_1273,N_49830,N_49996);
nor UO_1274 (O_1274,N_49937,N_49908);
xnor UO_1275 (O_1275,N_49841,N_49892);
xnor UO_1276 (O_1276,N_49914,N_49867);
xor UO_1277 (O_1277,N_49771,N_49973);
nand UO_1278 (O_1278,N_49990,N_49828);
xnor UO_1279 (O_1279,N_49819,N_49969);
nand UO_1280 (O_1280,N_49907,N_49911);
nand UO_1281 (O_1281,N_49823,N_49783);
or UO_1282 (O_1282,N_49764,N_49750);
or UO_1283 (O_1283,N_49751,N_49828);
nand UO_1284 (O_1284,N_49779,N_49929);
nor UO_1285 (O_1285,N_49784,N_49896);
nor UO_1286 (O_1286,N_49874,N_49889);
nand UO_1287 (O_1287,N_49859,N_49996);
nand UO_1288 (O_1288,N_49813,N_49803);
nand UO_1289 (O_1289,N_49888,N_49817);
nor UO_1290 (O_1290,N_49807,N_49972);
and UO_1291 (O_1291,N_49861,N_49889);
and UO_1292 (O_1292,N_49869,N_49898);
xor UO_1293 (O_1293,N_49914,N_49842);
nor UO_1294 (O_1294,N_49776,N_49813);
or UO_1295 (O_1295,N_49863,N_49833);
and UO_1296 (O_1296,N_49883,N_49997);
nand UO_1297 (O_1297,N_49793,N_49939);
or UO_1298 (O_1298,N_49925,N_49776);
or UO_1299 (O_1299,N_49925,N_49886);
or UO_1300 (O_1300,N_49960,N_49932);
and UO_1301 (O_1301,N_49922,N_49899);
nand UO_1302 (O_1302,N_49845,N_49970);
and UO_1303 (O_1303,N_49985,N_49818);
nand UO_1304 (O_1304,N_49853,N_49763);
or UO_1305 (O_1305,N_49950,N_49829);
or UO_1306 (O_1306,N_49752,N_49795);
or UO_1307 (O_1307,N_49765,N_49759);
and UO_1308 (O_1308,N_49792,N_49770);
and UO_1309 (O_1309,N_49849,N_49870);
xor UO_1310 (O_1310,N_49812,N_49900);
xnor UO_1311 (O_1311,N_49811,N_49822);
xnor UO_1312 (O_1312,N_49987,N_49850);
xor UO_1313 (O_1313,N_49932,N_49826);
or UO_1314 (O_1314,N_49879,N_49952);
and UO_1315 (O_1315,N_49910,N_49815);
xnor UO_1316 (O_1316,N_49878,N_49938);
xnor UO_1317 (O_1317,N_49895,N_49926);
xor UO_1318 (O_1318,N_49954,N_49976);
nor UO_1319 (O_1319,N_49795,N_49962);
nand UO_1320 (O_1320,N_49971,N_49980);
or UO_1321 (O_1321,N_49970,N_49936);
and UO_1322 (O_1322,N_49939,N_49948);
nor UO_1323 (O_1323,N_49869,N_49922);
or UO_1324 (O_1324,N_49953,N_49987);
and UO_1325 (O_1325,N_49958,N_49806);
and UO_1326 (O_1326,N_49798,N_49811);
nand UO_1327 (O_1327,N_49903,N_49870);
nor UO_1328 (O_1328,N_49949,N_49844);
and UO_1329 (O_1329,N_49904,N_49998);
or UO_1330 (O_1330,N_49831,N_49959);
nand UO_1331 (O_1331,N_49768,N_49835);
nor UO_1332 (O_1332,N_49996,N_49914);
nand UO_1333 (O_1333,N_49776,N_49954);
nand UO_1334 (O_1334,N_49919,N_49996);
nor UO_1335 (O_1335,N_49856,N_49772);
and UO_1336 (O_1336,N_49939,N_49782);
nand UO_1337 (O_1337,N_49954,N_49916);
xnor UO_1338 (O_1338,N_49786,N_49905);
or UO_1339 (O_1339,N_49925,N_49861);
nor UO_1340 (O_1340,N_49920,N_49763);
nand UO_1341 (O_1341,N_49753,N_49917);
or UO_1342 (O_1342,N_49952,N_49910);
nor UO_1343 (O_1343,N_49806,N_49962);
and UO_1344 (O_1344,N_49954,N_49939);
nor UO_1345 (O_1345,N_49942,N_49776);
nand UO_1346 (O_1346,N_49992,N_49999);
or UO_1347 (O_1347,N_49921,N_49969);
and UO_1348 (O_1348,N_49782,N_49841);
or UO_1349 (O_1349,N_49751,N_49984);
xor UO_1350 (O_1350,N_49880,N_49979);
or UO_1351 (O_1351,N_49892,N_49992);
and UO_1352 (O_1352,N_49770,N_49778);
nor UO_1353 (O_1353,N_49806,N_49960);
or UO_1354 (O_1354,N_49843,N_49935);
nand UO_1355 (O_1355,N_49912,N_49970);
and UO_1356 (O_1356,N_49993,N_49871);
nand UO_1357 (O_1357,N_49786,N_49860);
nor UO_1358 (O_1358,N_49837,N_49759);
nor UO_1359 (O_1359,N_49999,N_49810);
and UO_1360 (O_1360,N_49937,N_49825);
and UO_1361 (O_1361,N_49912,N_49755);
nand UO_1362 (O_1362,N_49784,N_49876);
nor UO_1363 (O_1363,N_49868,N_49867);
and UO_1364 (O_1364,N_49912,N_49952);
xor UO_1365 (O_1365,N_49928,N_49803);
and UO_1366 (O_1366,N_49754,N_49952);
nor UO_1367 (O_1367,N_49870,N_49912);
or UO_1368 (O_1368,N_49811,N_49993);
nor UO_1369 (O_1369,N_49780,N_49851);
or UO_1370 (O_1370,N_49850,N_49789);
nand UO_1371 (O_1371,N_49883,N_49768);
and UO_1372 (O_1372,N_49968,N_49853);
nor UO_1373 (O_1373,N_49937,N_49800);
xnor UO_1374 (O_1374,N_49828,N_49837);
nor UO_1375 (O_1375,N_49831,N_49846);
nand UO_1376 (O_1376,N_49966,N_49917);
xnor UO_1377 (O_1377,N_49848,N_49986);
and UO_1378 (O_1378,N_49890,N_49814);
or UO_1379 (O_1379,N_49951,N_49805);
nand UO_1380 (O_1380,N_49813,N_49891);
or UO_1381 (O_1381,N_49920,N_49755);
nand UO_1382 (O_1382,N_49952,N_49759);
nand UO_1383 (O_1383,N_49961,N_49923);
xor UO_1384 (O_1384,N_49837,N_49791);
or UO_1385 (O_1385,N_49798,N_49844);
nor UO_1386 (O_1386,N_49971,N_49812);
nor UO_1387 (O_1387,N_49976,N_49910);
and UO_1388 (O_1388,N_49913,N_49892);
xor UO_1389 (O_1389,N_49798,N_49957);
nor UO_1390 (O_1390,N_49892,N_49989);
xor UO_1391 (O_1391,N_49874,N_49779);
and UO_1392 (O_1392,N_49761,N_49864);
and UO_1393 (O_1393,N_49775,N_49810);
or UO_1394 (O_1394,N_49843,N_49809);
or UO_1395 (O_1395,N_49825,N_49847);
nand UO_1396 (O_1396,N_49790,N_49795);
and UO_1397 (O_1397,N_49838,N_49789);
nor UO_1398 (O_1398,N_49933,N_49935);
nor UO_1399 (O_1399,N_49770,N_49912);
or UO_1400 (O_1400,N_49815,N_49928);
nor UO_1401 (O_1401,N_49804,N_49932);
and UO_1402 (O_1402,N_49756,N_49983);
xnor UO_1403 (O_1403,N_49899,N_49823);
nand UO_1404 (O_1404,N_49925,N_49933);
xnor UO_1405 (O_1405,N_49878,N_49792);
and UO_1406 (O_1406,N_49985,N_49814);
nor UO_1407 (O_1407,N_49786,N_49856);
and UO_1408 (O_1408,N_49965,N_49810);
nand UO_1409 (O_1409,N_49822,N_49899);
and UO_1410 (O_1410,N_49843,N_49837);
and UO_1411 (O_1411,N_49878,N_49964);
nand UO_1412 (O_1412,N_49978,N_49894);
and UO_1413 (O_1413,N_49886,N_49987);
xor UO_1414 (O_1414,N_49832,N_49808);
and UO_1415 (O_1415,N_49846,N_49897);
xor UO_1416 (O_1416,N_49886,N_49816);
xor UO_1417 (O_1417,N_49974,N_49883);
nand UO_1418 (O_1418,N_49775,N_49900);
or UO_1419 (O_1419,N_49767,N_49898);
nand UO_1420 (O_1420,N_49959,N_49801);
nand UO_1421 (O_1421,N_49880,N_49850);
nor UO_1422 (O_1422,N_49753,N_49875);
nor UO_1423 (O_1423,N_49816,N_49940);
xor UO_1424 (O_1424,N_49906,N_49993);
xor UO_1425 (O_1425,N_49778,N_49847);
and UO_1426 (O_1426,N_49897,N_49769);
and UO_1427 (O_1427,N_49812,N_49752);
or UO_1428 (O_1428,N_49895,N_49971);
nand UO_1429 (O_1429,N_49977,N_49756);
and UO_1430 (O_1430,N_49904,N_49965);
xor UO_1431 (O_1431,N_49884,N_49829);
nor UO_1432 (O_1432,N_49853,N_49803);
nand UO_1433 (O_1433,N_49943,N_49839);
or UO_1434 (O_1434,N_49849,N_49828);
nor UO_1435 (O_1435,N_49989,N_49979);
nor UO_1436 (O_1436,N_49863,N_49941);
nand UO_1437 (O_1437,N_49917,N_49942);
nand UO_1438 (O_1438,N_49977,N_49866);
nand UO_1439 (O_1439,N_49814,N_49769);
nand UO_1440 (O_1440,N_49779,N_49960);
nand UO_1441 (O_1441,N_49792,N_49903);
or UO_1442 (O_1442,N_49989,N_49790);
nor UO_1443 (O_1443,N_49953,N_49794);
nand UO_1444 (O_1444,N_49967,N_49844);
nor UO_1445 (O_1445,N_49897,N_49858);
or UO_1446 (O_1446,N_49784,N_49972);
xnor UO_1447 (O_1447,N_49784,N_49754);
nand UO_1448 (O_1448,N_49907,N_49942);
nand UO_1449 (O_1449,N_49835,N_49821);
xor UO_1450 (O_1450,N_49952,N_49963);
or UO_1451 (O_1451,N_49830,N_49797);
xor UO_1452 (O_1452,N_49785,N_49958);
nand UO_1453 (O_1453,N_49954,N_49970);
and UO_1454 (O_1454,N_49836,N_49881);
or UO_1455 (O_1455,N_49815,N_49794);
nand UO_1456 (O_1456,N_49813,N_49970);
or UO_1457 (O_1457,N_49910,N_49838);
xor UO_1458 (O_1458,N_49888,N_49945);
nand UO_1459 (O_1459,N_49924,N_49962);
and UO_1460 (O_1460,N_49992,N_49840);
nor UO_1461 (O_1461,N_49788,N_49959);
xor UO_1462 (O_1462,N_49985,N_49871);
nand UO_1463 (O_1463,N_49796,N_49893);
and UO_1464 (O_1464,N_49950,N_49864);
and UO_1465 (O_1465,N_49865,N_49911);
and UO_1466 (O_1466,N_49764,N_49952);
nand UO_1467 (O_1467,N_49778,N_49964);
nor UO_1468 (O_1468,N_49922,N_49902);
xor UO_1469 (O_1469,N_49941,N_49899);
or UO_1470 (O_1470,N_49777,N_49763);
nand UO_1471 (O_1471,N_49948,N_49839);
xor UO_1472 (O_1472,N_49774,N_49975);
nor UO_1473 (O_1473,N_49880,N_49813);
nor UO_1474 (O_1474,N_49974,N_49989);
and UO_1475 (O_1475,N_49938,N_49941);
xnor UO_1476 (O_1476,N_49811,N_49893);
or UO_1477 (O_1477,N_49803,N_49947);
nand UO_1478 (O_1478,N_49891,N_49964);
xor UO_1479 (O_1479,N_49825,N_49909);
nand UO_1480 (O_1480,N_49996,N_49890);
or UO_1481 (O_1481,N_49980,N_49911);
nor UO_1482 (O_1482,N_49815,N_49966);
nor UO_1483 (O_1483,N_49817,N_49954);
or UO_1484 (O_1484,N_49789,N_49893);
or UO_1485 (O_1485,N_49813,N_49975);
nand UO_1486 (O_1486,N_49948,N_49950);
or UO_1487 (O_1487,N_49950,N_49757);
or UO_1488 (O_1488,N_49981,N_49878);
or UO_1489 (O_1489,N_49778,N_49832);
nand UO_1490 (O_1490,N_49912,N_49866);
and UO_1491 (O_1491,N_49947,N_49852);
and UO_1492 (O_1492,N_49800,N_49812);
nor UO_1493 (O_1493,N_49862,N_49960);
xor UO_1494 (O_1494,N_49822,N_49940);
and UO_1495 (O_1495,N_49947,N_49916);
nor UO_1496 (O_1496,N_49810,N_49922);
and UO_1497 (O_1497,N_49909,N_49830);
xor UO_1498 (O_1498,N_49886,N_49856);
or UO_1499 (O_1499,N_49876,N_49845);
nand UO_1500 (O_1500,N_49759,N_49959);
xor UO_1501 (O_1501,N_49808,N_49919);
or UO_1502 (O_1502,N_49752,N_49826);
nand UO_1503 (O_1503,N_49996,N_49948);
or UO_1504 (O_1504,N_49929,N_49758);
or UO_1505 (O_1505,N_49897,N_49790);
or UO_1506 (O_1506,N_49914,N_49800);
nor UO_1507 (O_1507,N_49811,N_49991);
xor UO_1508 (O_1508,N_49757,N_49962);
or UO_1509 (O_1509,N_49862,N_49759);
nand UO_1510 (O_1510,N_49877,N_49842);
nand UO_1511 (O_1511,N_49982,N_49974);
nand UO_1512 (O_1512,N_49957,N_49750);
nor UO_1513 (O_1513,N_49871,N_49805);
nand UO_1514 (O_1514,N_49983,N_49880);
and UO_1515 (O_1515,N_49843,N_49813);
nand UO_1516 (O_1516,N_49954,N_49917);
xnor UO_1517 (O_1517,N_49890,N_49994);
nor UO_1518 (O_1518,N_49760,N_49766);
nand UO_1519 (O_1519,N_49777,N_49805);
nor UO_1520 (O_1520,N_49794,N_49909);
nand UO_1521 (O_1521,N_49811,N_49784);
nor UO_1522 (O_1522,N_49778,N_49817);
or UO_1523 (O_1523,N_49892,N_49961);
xor UO_1524 (O_1524,N_49960,N_49997);
or UO_1525 (O_1525,N_49847,N_49779);
xor UO_1526 (O_1526,N_49768,N_49763);
nand UO_1527 (O_1527,N_49987,N_49966);
nand UO_1528 (O_1528,N_49795,N_49990);
and UO_1529 (O_1529,N_49870,N_49842);
xor UO_1530 (O_1530,N_49873,N_49980);
nor UO_1531 (O_1531,N_49819,N_49768);
xnor UO_1532 (O_1532,N_49857,N_49863);
nor UO_1533 (O_1533,N_49754,N_49867);
or UO_1534 (O_1534,N_49839,N_49821);
or UO_1535 (O_1535,N_49865,N_49759);
nand UO_1536 (O_1536,N_49827,N_49931);
nor UO_1537 (O_1537,N_49994,N_49978);
and UO_1538 (O_1538,N_49761,N_49845);
nand UO_1539 (O_1539,N_49985,N_49843);
nand UO_1540 (O_1540,N_49815,N_49963);
and UO_1541 (O_1541,N_49778,N_49898);
and UO_1542 (O_1542,N_49964,N_49954);
nor UO_1543 (O_1543,N_49974,N_49925);
nor UO_1544 (O_1544,N_49753,N_49918);
nand UO_1545 (O_1545,N_49914,N_49871);
or UO_1546 (O_1546,N_49797,N_49824);
xor UO_1547 (O_1547,N_49821,N_49931);
nor UO_1548 (O_1548,N_49839,N_49888);
or UO_1549 (O_1549,N_49961,N_49821);
nand UO_1550 (O_1550,N_49766,N_49756);
and UO_1551 (O_1551,N_49750,N_49907);
and UO_1552 (O_1552,N_49872,N_49974);
xnor UO_1553 (O_1553,N_49764,N_49901);
xor UO_1554 (O_1554,N_49980,N_49947);
and UO_1555 (O_1555,N_49846,N_49919);
or UO_1556 (O_1556,N_49821,N_49847);
or UO_1557 (O_1557,N_49984,N_49796);
and UO_1558 (O_1558,N_49808,N_49942);
nor UO_1559 (O_1559,N_49865,N_49784);
or UO_1560 (O_1560,N_49856,N_49794);
nand UO_1561 (O_1561,N_49974,N_49891);
nor UO_1562 (O_1562,N_49932,N_49912);
nand UO_1563 (O_1563,N_49937,N_49957);
xnor UO_1564 (O_1564,N_49961,N_49766);
nand UO_1565 (O_1565,N_49919,N_49987);
or UO_1566 (O_1566,N_49895,N_49770);
or UO_1567 (O_1567,N_49811,N_49755);
xnor UO_1568 (O_1568,N_49991,N_49814);
nand UO_1569 (O_1569,N_49902,N_49800);
and UO_1570 (O_1570,N_49862,N_49840);
nand UO_1571 (O_1571,N_49909,N_49912);
nand UO_1572 (O_1572,N_49784,N_49835);
xnor UO_1573 (O_1573,N_49799,N_49783);
or UO_1574 (O_1574,N_49810,N_49888);
nor UO_1575 (O_1575,N_49819,N_49832);
nor UO_1576 (O_1576,N_49819,N_49985);
nand UO_1577 (O_1577,N_49800,N_49861);
nor UO_1578 (O_1578,N_49925,N_49864);
nor UO_1579 (O_1579,N_49898,N_49913);
or UO_1580 (O_1580,N_49866,N_49952);
and UO_1581 (O_1581,N_49842,N_49814);
xnor UO_1582 (O_1582,N_49975,N_49902);
nand UO_1583 (O_1583,N_49767,N_49834);
xor UO_1584 (O_1584,N_49984,N_49996);
and UO_1585 (O_1585,N_49973,N_49905);
and UO_1586 (O_1586,N_49822,N_49770);
and UO_1587 (O_1587,N_49904,N_49826);
and UO_1588 (O_1588,N_49756,N_49821);
nand UO_1589 (O_1589,N_49816,N_49882);
nor UO_1590 (O_1590,N_49970,N_49891);
xor UO_1591 (O_1591,N_49775,N_49849);
nand UO_1592 (O_1592,N_49776,N_49886);
and UO_1593 (O_1593,N_49935,N_49888);
or UO_1594 (O_1594,N_49802,N_49765);
xnor UO_1595 (O_1595,N_49985,N_49969);
nor UO_1596 (O_1596,N_49800,N_49978);
or UO_1597 (O_1597,N_49981,N_49959);
and UO_1598 (O_1598,N_49957,N_49960);
xor UO_1599 (O_1599,N_49867,N_49964);
nand UO_1600 (O_1600,N_49918,N_49797);
and UO_1601 (O_1601,N_49955,N_49752);
nand UO_1602 (O_1602,N_49917,N_49976);
and UO_1603 (O_1603,N_49924,N_49920);
nor UO_1604 (O_1604,N_49854,N_49991);
xnor UO_1605 (O_1605,N_49910,N_49812);
nor UO_1606 (O_1606,N_49811,N_49792);
nand UO_1607 (O_1607,N_49924,N_49946);
nand UO_1608 (O_1608,N_49926,N_49750);
or UO_1609 (O_1609,N_49939,N_49846);
nor UO_1610 (O_1610,N_49841,N_49929);
nand UO_1611 (O_1611,N_49964,N_49916);
nor UO_1612 (O_1612,N_49999,N_49781);
and UO_1613 (O_1613,N_49972,N_49903);
xnor UO_1614 (O_1614,N_49976,N_49875);
and UO_1615 (O_1615,N_49973,N_49853);
xnor UO_1616 (O_1616,N_49968,N_49965);
nand UO_1617 (O_1617,N_49803,N_49857);
and UO_1618 (O_1618,N_49908,N_49945);
or UO_1619 (O_1619,N_49836,N_49989);
and UO_1620 (O_1620,N_49924,N_49794);
or UO_1621 (O_1621,N_49833,N_49793);
xor UO_1622 (O_1622,N_49960,N_49879);
nand UO_1623 (O_1623,N_49843,N_49757);
or UO_1624 (O_1624,N_49816,N_49910);
xnor UO_1625 (O_1625,N_49916,N_49872);
and UO_1626 (O_1626,N_49893,N_49829);
or UO_1627 (O_1627,N_49976,N_49817);
and UO_1628 (O_1628,N_49968,N_49912);
or UO_1629 (O_1629,N_49883,N_49758);
xnor UO_1630 (O_1630,N_49766,N_49929);
nand UO_1631 (O_1631,N_49761,N_49838);
nand UO_1632 (O_1632,N_49755,N_49770);
xnor UO_1633 (O_1633,N_49853,N_49989);
or UO_1634 (O_1634,N_49798,N_49896);
xnor UO_1635 (O_1635,N_49954,N_49856);
nand UO_1636 (O_1636,N_49938,N_49882);
nor UO_1637 (O_1637,N_49786,N_49957);
and UO_1638 (O_1638,N_49964,N_49992);
nor UO_1639 (O_1639,N_49984,N_49828);
or UO_1640 (O_1640,N_49771,N_49773);
nand UO_1641 (O_1641,N_49830,N_49832);
and UO_1642 (O_1642,N_49853,N_49868);
xnor UO_1643 (O_1643,N_49797,N_49786);
nand UO_1644 (O_1644,N_49826,N_49761);
and UO_1645 (O_1645,N_49763,N_49955);
and UO_1646 (O_1646,N_49918,N_49774);
nand UO_1647 (O_1647,N_49828,N_49945);
nand UO_1648 (O_1648,N_49794,N_49768);
and UO_1649 (O_1649,N_49760,N_49995);
xor UO_1650 (O_1650,N_49750,N_49805);
xor UO_1651 (O_1651,N_49911,N_49864);
nor UO_1652 (O_1652,N_49807,N_49776);
or UO_1653 (O_1653,N_49879,N_49876);
nor UO_1654 (O_1654,N_49854,N_49771);
nor UO_1655 (O_1655,N_49798,N_49826);
xor UO_1656 (O_1656,N_49912,N_49973);
nand UO_1657 (O_1657,N_49930,N_49860);
xor UO_1658 (O_1658,N_49758,N_49984);
or UO_1659 (O_1659,N_49790,N_49874);
nor UO_1660 (O_1660,N_49992,N_49854);
nand UO_1661 (O_1661,N_49948,N_49893);
nand UO_1662 (O_1662,N_49903,N_49839);
xnor UO_1663 (O_1663,N_49837,N_49836);
and UO_1664 (O_1664,N_49860,N_49945);
and UO_1665 (O_1665,N_49982,N_49882);
nand UO_1666 (O_1666,N_49760,N_49915);
xnor UO_1667 (O_1667,N_49799,N_49882);
or UO_1668 (O_1668,N_49899,N_49836);
nor UO_1669 (O_1669,N_49901,N_49868);
or UO_1670 (O_1670,N_49963,N_49865);
and UO_1671 (O_1671,N_49931,N_49929);
xor UO_1672 (O_1672,N_49809,N_49942);
nand UO_1673 (O_1673,N_49856,N_49768);
nand UO_1674 (O_1674,N_49849,N_49853);
and UO_1675 (O_1675,N_49804,N_49857);
nor UO_1676 (O_1676,N_49988,N_49816);
nor UO_1677 (O_1677,N_49869,N_49775);
and UO_1678 (O_1678,N_49820,N_49984);
and UO_1679 (O_1679,N_49837,N_49770);
nand UO_1680 (O_1680,N_49827,N_49883);
xor UO_1681 (O_1681,N_49758,N_49898);
nand UO_1682 (O_1682,N_49991,N_49908);
and UO_1683 (O_1683,N_49822,N_49984);
nor UO_1684 (O_1684,N_49913,N_49760);
and UO_1685 (O_1685,N_49902,N_49854);
or UO_1686 (O_1686,N_49804,N_49806);
and UO_1687 (O_1687,N_49811,N_49916);
nand UO_1688 (O_1688,N_49780,N_49921);
and UO_1689 (O_1689,N_49893,N_49777);
nand UO_1690 (O_1690,N_49904,N_49811);
nand UO_1691 (O_1691,N_49971,N_49797);
or UO_1692 (O_1692,N_49810,N_49909);
nor UO_1693 (O_1693,N_49770,N_49915);
and UO_1694 (O_1694,N_49874,N_49808);
xnor UO_1695 (O_1695,N_49920,N_49936);
and UO_1696 (O_1696,N_49766,N_49870);
xnor UO_1697 (O_1697,N_49849,N_49948);
or UO_1698 (O_1698,N_49965,N_49997);
xor UO_1699 (O_1699,N_49981,N_49983);
xor UO_1700 (O_1700,N_49859,N_49973);
or UO_1701 (O_1701,N_49854,N_49904);
nand UO_1702 (O_1702,N_49948,N_49852);
nor UO_1703 (O_1703,N_49915,N_49880);
xor UO_1704 (O_1704,N_49764,N_49785);
xnor UO_1705 (O_1705,N_49839,N_49797);
nor UO_1706 (O_1706,N_49978,N_49827);
nor UO_1707 (O_1707,N_49862,N_49872);
and UO_1708 (O_1708,N_49898,N_49802);
or UO_1709 (O_1709,N_49986,N_49916);
xor UO_1710 (O_1710,N_49811,N_49851);
nand UO_1711 (O_1711,N_49809,N_49977);
and UO_1712 (O_1712,N_49766,N_49927);
and UO_1713 (O_1713,N_49956,N_49995);
or UO_1714 (O_1714,N_49833,N_49972);
or UO_1715 (O_1715,N_49852,N_49934);
nand UO_1716 (O_1716,N_49884,N_49824);
and UO_1717 (O_1717,N_49947,N_49996);
or UO_1718 (O_1718,N_49925,N_49900);
nand UO_1719 (O_1719,N_49802,N_49869);
or UO_1720 (O_1720,N_49990,N_49753);
and UO_1721 (O_1721,N_49865,N_49971);
and UO_1722 (O_1722,N_49788,N_49870);
or UO_1723 (O_1723,N_49801,N_49996);
nor UO_1724 (O_1724,N_49760,N_49885);
nand UO_1725 (O_1725,N_49888,N_49904);
xor UO_1726 (O_1726,N_49818,N_49814);
nor UO_1727 (O_1727,N_49798,N_49856);
and UO_1728 (O_1728,N_49899,N_49837);
or UO_1729 (O_1729,N_49751,N_49897);
nand UO_1730 (O_1730,N_49800,N_49756);
nand UO_1731 (O_1731,N_49870,N_49795);
xnor UO_1732 (O_1732,N_49938,N_49916);
or UO_1733 (O_1733,N_49966,N_49803);
nand UO_1734 (O_1734,N_49927,N_49942);
nand UO_1735 (O_1735,N_49787,N_49930);
or UO_1736 (O_1736,N_49757,N_49857);
or UO_1737 (O_1737,N_49954,N_49779);
nor UO_1738 (O_1738,N_49959,N_49807);
nor UO_1739 (O_1739,N_49920,N_49776);
xor UO_1740 (O_1740,N_49866,N_49891);
nand UO_1741 (O_1741,N_49890,N_49750);
and UO_1742 (O_1742,N_49868,N_49835);
and UO_1743 (O_1743,N_49931,N_49785);
or UO_1744 (O_1744,N_49848,N_49845);
and UO_1745 (O_1745,N_49883,N_49916);
nand UO_1746 (O_1746,N_49992,N_49988);
xor UO_1747 (O_1747,N_49904,N_49813);
nor UO_1748 (O_1748,N_49784,N_49929);
xor UO_1749 (O_1749,N_49895,N_49778);
nand UO_1750 (O_1750,N_49999,N_49989);
or UO_1751 (O_1751,N_49834,N_49995);
nor UO_1752 (O_1752,N_49954,N_49996);
or UO_1753 (O_1753,N_49845,N_49954);
or UO_1754 (O_1754,N_49838,N_49755);
nor UO_1755 (O_1755,N_49843,N_49797);
or UO_1756 (O_1756,N_49840,N_49993);
and UO_1757 (O_1757,N_49764,N_49790);
xnor UO_1758 (O_1758,N_49802,N_49970);
and UO_1759 (O_1759,N_49755,N_49921);
xnor UO_1760 (O_1760,N_49854,N_49994);
and UO_1761 (O_1761,N_49848,N_49900);
and UO_1762 (O_1762,N_49981,N_49868);
xor UO_1763 (O_1763,N_49959,N_49770);
or UO_1764 (O_1764,N_49779,N_49984);
nor UO_1765 (O_1765,N_49943,N_49804);
nand UO_1766 (O_1766,N_49832,N_49833);
and UO_1767 (O_1767,N_49902,N_49763);
xnor UO_1768 (O_1768,N_49898,N_49964);
and UO_1769 (O_1769,N_49903,N_49890);
or UO_1770 (O_1770,N_49956,N_49797);
nor UO_1771 (O_1771,N_49974,N_49878);
or UO_1772 (O_1772,N_49804,N_49945);
xor UO_1773 (O_1773,N_49811,N_49818);
nor UO_1774 (O_1774,N_49824,N_49772);
nor UO_1775 (O_1775,N_49843,N_49804);
or UO_1776 (O_1776,N_49979,N_49824);
or UO_1777 (O_1777,N_49922,N_49759);
xor UO_1778 (O_1778,N_49963,N_49923);
nand UO_1779 (O_1779,N_49751,N_49839);
nand UO_1780 (O_1780,N_49769,N_49778);
nor UO_1781 (O_1781,N_49858,N_49988);
nor UO_1782 (O_1782,N_49750,N_49840);
or UO_1783 (O_1783,N_49943,N_49935);
or UO_1784 (O_1784,N_49783,N_49875);
or UO_1785 (O_1785,N_49927,N_49792);
xor UO_1786 (O_1786,N_49770,N_49795);
nand UO_1787 (O_1787,N_49759,N_49956);
xor UO_1788 (O_1788,N_49887,N_49784);
xor UO_1789 (O_1789,N_49911,N_49893);
nand UO_1790 (O_1790,N_49925,N_49942);
nor UO_1791 (O_1791,N_49846,N_49941);
nor UO_1792 (O_1792,N_49886,N_49855);
xor UO_1793 (O_1793,N_49990,N_49930);
nor UO_1794 (O_1794,N_49894,N_49932);
nand UO_1795 (O_1795,N_49869,N_49999);
and UO_1796 (O_1796,N_49779,N_49840);
nor UO_1797 (O_1797,N_49759,N_49818);
xnor UO_1798 (O_1798,N_49821,N_49937);
or UO_1799 (O_1799,N_49971,N_49813);
or UO_1800 (O_1800,N_49865,N_49775);
nand UO_1801 (O_1801,N_49830,N_49883);
nor UO_1802 (O_1802,N_49792,N_49926);
and UO_1803 (O_1803,N_49843,N_49866);
or UO_1804 (O_1804,N_49753,N_49859);
nor UO_1805 (O_1805,N_49805,N_49807);
or UO_1806 (O_1806,N_49780,N_49837);
nor UO_1807 (O_1807,N_49862,N_49921);
nand UO_1808 (O_1808,N_49962,N_49994);
and UO_1809 (O_1809,N_49871,N_49802);
nand UO_1810 (O_1810,N_49904,N_49948);
and UO_1811 (O_1811,N_49846,N_49974);
or UO_1812 (O_1812,N_49926,N_49899);
and UO_1813 (O_1813,N_49825,N_49853);
xor UO_1814 (O_1814,N_49908,N_49956);
nand UO_1815 (O_1815,N_49845,N_49945);
and UO_1816 (O_1816,N_49826,N_49928);
xor UO_1817 (O_1817,N_49969,N_49877);
or UO_1818 (O_1818,N_49772,N_49963);
or UO_1819 (O_1819,N_49934,N_49925);
xnor UO_1820 (O_1820,N_49897,N_49905);
or UO_1821 (O_1821,N_49881,N_49956);
and UO_1822 (O_1822,N_49996,N_49950);
xnor UO_1823 (O_1823,N_49932,N_49823);
or UO_1824 (O_1824,N_49764,N_49923);
xnor UO_1825 (O_1825,N_49968,N_49915);
nor UO_1826 (O_1826,N_49966,N_49985);
nand UO_1827 (O_1827,N_49785,N_49942);
nor UO_1828 (O_1828,N_49884,N_49767);
xor UO_1829 (O_1829,N_49757,N_49998);
nor UO_1830 (O_1830,N_49803,N_49992);
xnor UO_1831 (O_1831,N_49870,N_49908);
and UO_1832 (O_1832,N_49888,N_49777);
nand UO_1833 (O_1833,N_49985,N_49815);
xnor UO_1834 (O_1834,N_49986,N_49793);
nor UO_1835 (O_1835,N_49990,N_49791);
or UO_1836 (O_1836,N_49982,N_49837);
nand UO_1837 (O_1837,N_49988,N_49832);
and UO_1838 (O_1838,N_49763,N_49826);
nand UO_1839 (O_1839,N_49880,N_49883);
xor UO_1840 (O_1840,N_49960,N_49949);
and UO_1841 (O_1841,N_49932,N_49974);
and UO_1842 (O_1842,N_49779,N_49835);
xor UO_1843 (O_1843,N_49987,N_49908);
nor UO_1844 (O_1844,N_49951,N_49877);
xnor UO_1845 (O_1845,N_49898,N_49962);
nand UO_1846 (O_1846,N_49757,N_49817);
and UO_1847 (O_1847,N_49996,N_49845);
nand UO_1848 (O_1848,N_49909,N_49832);
and UO_1849 (O_1849,N_49898,N_49885);
or UO_1850 (O_1850,N_49976,N_49771);
and UO_1851 (O_1851,N_49969,N_49904);
nor UO_1852 (O_1852,N_49824,N_49768);
nand UO_1853 (O_1853,N_49814,N_49754);
and UO_1854 (O_1854,N_49795,N_49757);
and UO_1855 (O_1855,N_49961,N_49888);
nand UO_1856 (O_1856,N_49998,N_49751);
nor UO_1857 (O_1857,N_49796,N_49910);
and UO_1858 (O_1858,N_49822,N_49851);
nor UO_1859 (O_1859,N_49782,N_49988);
nor UO_1860 (O_1860,N_49940,N_49841);
or UO_1861 (O_1861,N_49911,N_49754);
nor UO_1862 (O_1862,N_49752,N_49791);
xor UO_1863 (O_1863,N_49891,N_49918);
nand UO_1864 (O_1864,N_49827,N_49916);
nor UO_1865 (O_1865,N_49843,N_49869);
and UO_1866 (O_1866,N_49769,N_49982);
and UO_1867 (O_1867,N_49840,N_49998);
xor UO_1868 (O_1868,N_49789,N_49980);
nor UO_1869 (O_1869,N_49829,N_49841);
or UO_1870 (O_1870,N_49931,N_49756);
and UO_1871 (O_1871,N_49751,N_49978);
and UO_1872 (O_1872,N_49803,N_49758);
or UO_1873 (O_1873,N_49899,N_49906);
or UO_1874 (O_1874,N_49757,N_49845);
and UO_1875 (O_1875,N_49946,N_49987);
nand UO_1876 (O_1876,N_49930,N_49917);
nand UO_1877 (O_1877,N_49806,N_49826);
and UO_1878 (O_1878,N_49923,N_49939);
nor UO_1879 (O_1879,N_49973,N_49801);
or UO_1880 (O_1880,N_49928,N_49941);
or UO_1881 (O_1881,N_49950,N_49897);
and UO_1882 (O_1882,N_49912,N_49935);
or UO_1883 (O_1883,N_49961,N_49936);
nor UO_1884 (O_1884,N_49938,N_49837);
nand UO_1885 (O_1885,N_49990,N_49991);
and UO_1886 (O_1886,N_49926,N_49936);
and UO_1887 (O_1887,N_49866,N_49927);
or UO_1888 (O_1888,N_49927,N_49916);
or UO_1889 (O_1889,N_49768,N_49956);
and UO_1890 (O_1890,N_49934,N_49757);
nor UO_1891 (O_1891,N_49933,N_49889);
and UO_1892 (O_1892,N_49823,N_49804);
nor UO_1893 (O_1893,N_49786,N_49830);
nand UO_1894 (O_1894,N_49810,N_49804);
or UO_1895 (O_1895,N_49989,N_49881);
or UO_1896 (O_1896,N_49930,N_49797);
nor UO_1897 (O_1897,N_49934,N_49989);
and UO_1898 (O_1898,N_49778,N_49824);
xor UO_1899 (O_1899,N_49861,N_49811);
nor UO_1900 (O_1900,N_49798,N_49932);
and UO_1901 (O_1901,N_49877,N_49809);
nor UO_1902 (O_1902,N_49813,N_49810);
and UO_1903 (O_1903,N_49951,N_49871);
and UO_1904 (O_1904,N_49837,N_49926);
xnor UO_1905 (O_1905,N_49827,N_49869);
xor UO_1906 (O_1906,N_49907,N_49826);
xor UO_1907 (O_1907,N_49820,N_49912);
xnor UO_1908 (O_1908,N_49982,N_49840);
and UO_1909 (O_1909,N_49806,N_49797);
nand UO_1910 (O_1910,N_49920,N_49855);
or UO_1911 (O_1911,N_49891,N_49863);
and UO_1912 (O_1912,N_49804,N_49852);
or UO_1913 (O_1913,N_49950,N_49938);
nand UO_1914 (O_1914,N_49916,N_49908);
xor UO_1915 (O_1915,N_49836,N_49980);
nand UO_1916 (O_1916,N_49838,N_49867);
nand UO_1917 (O_1917,N_49836,N_49901);
xnor UO_1918 (O_1918,N_49931,N_49949);
xor UO_1919 (O_1919,N_49855,N_49988);
nand UO_1920 (O_1920,N_49766,N_49984);
nor UO_1921 (O_1921,N_49774,N_49773);
nor UO_1922 (O_1922,N_49882,N_49855);
nor UO_1923 (O_1923,N_49820,N_49891);
and UO_1924 (O_1924,N_49923,N_49852);
xor UO_1925 (O_1925,N_49973,N_49819);
nor UO_1926 (O_1926,N_49797,N_49935);
nand UO_1927 (O_1927,N_49790,N_49854);
and UO_1928 (O_1928,N_49936,N_49832);
xor UO_1929 (O_1929,N_49843,N_49943);
nand UO_1930 (O_1930,N_49866,N_49943);
and UO_1931 (O_1931,N_49826,N_49895);
xor UO_1932 (O_1932,N_49920,N_49914);
or UO_1933 (O_1933,N_49750,N_49837);
and UO_1934 (O_1934,N_49978,N_49996);
nand UO_1935 (O_1935,N_49801,N_49788);
and UO_1936 (O_1936,N_49800,N_49783);
and UO_1937 (O_1937,N_49987,N_49805);
nand UO_1938 (O_1938,N_49788,N_49796);
xnor UO_1939 (O_1939,N_49886,N_49753);
or UO_1940 (O_1940,N_49922,N_49762);
nand UO_1941 (O_1941,N_49811,N_49912);
and UO_1942 (O_1942,N_49902,N_49805);
nand UO_1943 (O_1943,N_49874,N_49891);
xnor UO_1944 (O_1944,N_49856,N_49946);
nor UO_1945 (O_1945,N_49939,N_49766);
nor UO_1946 (O_1946,N_49931,N_49753);
and UO_1947 (O_1947,N_49891,N_49808);
or UO_1948 (O_1948,N_49916,N_49937);
nand UO_1949 (O_1949,N_49840,N_49886);
xor UO_1950 (O_1950,N_49856,N_49921);
xnor UO_1951 (O_1951,N_49783,N_49949);
or UO_1952 (O_1952,N_49788,N_49912);
and UO_1953 (O_1953,N_49795,N_49987);
nand UO_1954 (O_1954,N_49880,N_49897);
nor UO_1955 (O_1955,N_49920,N_49822);
nor UO_1956 (O_1956,N_49796,N_49763);
or UO_1957 (O_1957,N_49884,N_49986);
or UO_1958 (O_1958,N_49806,N_49817);
nand UO_1959 (O_1959,N_49900,N_49797);
and UO_1960 (O_1960,N_49793,N_49887);
nor UO_1961 (O_1961,N_49935,N_49817);
nor UO_1962 (O_1962,N_49779,N_49867);
nand UO_1963 (O_1963,N_49831,N_49771);
nor UO_1964 (O_1964,N_49908,N_49971);
nand UO_1965 (O_1965,N_49805,N_49904);
nand UO_1966 (O_1966,N_49796,N_49898);
and UO_1967 (O_1967,N_49973,N_49828);
or UO_1968 (O_1968,N_49925,N_49788);
and UO_1969 (O_1969,N_49753,N_49869);
xnor UO_1970 (O_1970,N_49769,N_49828);
nand UO_1971 (O_1971,N_49900,N_49915);
or UO_1972 (O_1972,N_49771,N_49966);
xnor UO_1973 (O_1973,N_49900,N_49780);
or UO_1974 (O_1974,N_49758,N_49968);
and UO_1975 (O_1975,N_49992,N_49969);
nor UO_1976 (O_1976,N_49956,N_49803);
nor UO_1977 (O_1977,N_49892,N_49827);
xor UO_1978 (O_1978,N_49940,N_49973);
nor UO_1979 (O_1979,N_49944,N_49913);
and UO_1980 (O_1980,N_49967,N_49802);
and UO_1981 (O_1981,N_49986,N_49945);
nand UO_1982 (O_1982,N_49916,N_49929);
nor UO_1983 (O_1983,N_49963,N_49779);
or UO_1984 (O_1984,N_49885,N_49800);
nand UO_1985 (O_1985,N_49931,N_49796);
and UO_1986 (O_1986,N_49967,N_49830);
xnor UO_1987 (O_1987,N_49837,N_49820);
or UO_1988 (O_1988,N_49920,N_49972);
or UO_1989 (O_1989,N_49908,N_49886);
nand UO_1990 (O_1990,N_49890,N_49882);
or UO_1991 (O_1991,N_49763,N_49992);
nor UO_1992 (O_1992,N_49930,N_49783);
nand UO_1993 (O_1993,N_49942,N_49974);
or UO_1994 (O_1994,N_49812,N_49865);
and UO_1995 (O_1995,N_49960,N_49896);
nor UO_1996 (O_1996,N_49800,N_49841);
nor UO_1997 (O_1997,N_49954,N_49946);
or UO_1998 (O_1998,N_49922,N_49804);
nor UO_1999 (O_1999,N_49966,N_49978);
nand UO_2000 (O_2000,N_49895,N_49815);
nand UO_2001 (O_2001,N_49969,N_49773);
or UO_2002 (O_2002,N_49995,N_49759);
or UO_2003 (O_2003,N_49829,N_49989);
nand UO_2004 (O_2004,N_49860,N_49927);
xnor UO_2005 (O_2005,N_49950,N_49840);
xor UO_2006 (O_2006,N_49867,N_49952);
xnor UO_2007 (O_2007,N_49903,N_49911);
nand UO_2008 (O_2008,N_49803,N_49954);
xor UO_2009 (O_2009,N_49953,N_49789);
or UO_2010 (O_2010,N_49999,N_49759);
xnor UO_2011 (O_2011,N_49847,N_49942);
and UO_2012 (O_2012,N_49840,N_49954);
and UO_2013 (O_2013,N_49952,N_49827);
and UO_2014 (O_2014,N_49833,N_49902);
and UO_2015 (O_2015,N_49896,N_49883);
nand UO_2016 (O_2016,N_49864,N_49991);
or UO_2017 (O_2017,N_49959,N_49886);
nor UO_2018 (O_2018,N_49775,N_49913);
and UO_2019 (O_2019,N_49841,N_49866);
and UO_2020 (O_2020,N_49869,N_49873);
nand UO_2021 (O_2021,N_49885,N_49813);
or UO_2022 (O_2022,N_49860,N_49820);
nand UO_2023 (O_2023,N_49751,N_49922);
xnor UO_2024 (O_2024,N_49960,N_49986);
xor UO_2025 (O_2025,N_49826,N_49947);
nor UO_2026 (O_2026,N_49808,N_49943);
nor UO_2027 (O_2027,N_49889,N_49828);
nor UO_2028 (O_2028,N_49955,N_49956);
nand UO_2029 (O_2029,N_49753,N_49754);
nand UO_2030 (O_2030,N_49995,N_49936);
nor UO_2031 (O_2031,N_49993,N_49822);
xnor UO_2032 (O_2032,N_49756,N_49930);
or UO_2033 (O_2033,N_49897,N_49797);
or UO_2034 (O_2034,N_49943,N_49949);
and UO_2035 (O_2035,N_49865,N_49848);
or UO_2036 (O_2036,N_49930,N_49937);
and UO_2037 (O_2037,N_49903,N_49892);
nor UO_2038 (O_2038,N_49794,N_49911);
and UO_2039 (O_2039,N_49809,N_49992);
nand UO_2040 (O_2040,N_49773,N_49979);
nand UO_2041 (O_2041,N_49943,N_49861);
or UO_2042 (O_2042,N_49951,N_49954);
and UO_2043 (O_2043,N_49834,N_49911);
xor UO_2044 (O_2044,N_49889,N_49982);
or UO_2045 (O_2045,N_49940,N_49829);
nand UO_2046 (O_2046,N_49800,N_49803);
nor UO_2047 (O_2047,N_49750,N_49970);
or UO_2048 (O_2048,N_49870,N_49799);
or UO_2049 (O_2049,N_49757,N_49896);
and UO_2050 (O_2050,N_49855,N_49947);
and UO_2051 (O_2051,N_49809,N_49817);
nand UO_2052 (O_2052,N_49989,N_49960);
or UO_2053 (O_2053,N_49750,N_49858);
nand UO_2054 (O_2054,N_49858,N_49921);
nand UO_2055 (O_2055,N_49849,N_49987);
or UO_2056 (O_2056,N_49810,N_49789);
nor UO_2057 (O_2057,N_49930,N_49788);
xor UO_2058 (O_2058,N_49805,N_49830);
nor UO_2059 (O_2059,N_49808,N_49838);
xor UO_2060 (O_2060,N_49933,N_49912);
nor UO_2061 (O_2061,N_49996,N_49941);
nor UO_2062 (O_2062,N_49808,N_49800);
and UO_2063 (O_2063,N_49782,N_49946);
nor UO_2064 (O_2064,N_49929,N_49863);
nand UO_2065 (O_2065,N_49852,N_49797);
nand UO_2066 (O_2066,N_49917,N_49936);
xor UO_2067 (O_2067,N_49991,N_49899);
nand UO_2068 (O_2068,N_49957,N_49873);
nand UO_2069 (O_2069,N_49982,N_49861);
or UO_2070 (O_2070,N_49878,N_49907);
and UO_2071 (O_2071,N_49794,N_49961);
nand UO_2072 (O_2072,N_49915,N_49898);
nand UO_2073 (O_2073,N_49983,N_49829);
nand UO_2074 (O_2074,N_49904,N_49853);
or UO_2075 (O_2075,N_49867,N_49962);
and UO_2076 (O_2076,N_49962,N_49802);
and UO_2077 (O_2077,N_49767,N_49964);
or UO_2078 (O_2078,N_49946,N_49774);
xnor UO_2079 (O_2079,N_49951,N_49853);
nand UO_2080 (O_2080,N_49949,N_49881);
or UO_2081 (O_2081,N_49973,N_49902);
or UO_2082 (O_2082,N_49854,N_49893);
nor UO_2083 (O_2083,N_49905,N_49762);
or UO_2084 (O_2084,N_49786,N_49782);
and UO_2085 (O_2085,N_49869,N_49979);
nand UO_2086 (O_2086,N_49873,N_49961);
nand UO_2087 (O_2087,N_49918,N_49953);
nand UO_2088 (O_2088,N_49909,N_49788);
and UO_2089 (O_2089,N_49773,N_49907);
and UO_2090 (O_2090,N_49774,N_49951);
or UO_2091 (O_2091,N_49945,N_49783);
xor UO_2092 (O_2092,N_49982,N_49957);
xnor UO_2093 (O_2093,N_49837,N_49873);
xnor UO_2094 (O_2094,N_49889,N_49958);
or UO_2095 (O_2095,N_49776,N_49775);
xor UO_2096 (O_2096,N_49845,N_49770);
nor UO_2097 (O_2097,N_49950,N_49968);
or UO_2098 (O_2098,N_49980,N_49782);
nand UO_2099 (O_2099,N_49913,N_49997);
nor UO_2100 (O_2100,N_49896,N_49852);
and UO_2101 (O_2101,N_49774,N_49849);
nor UO_2102 (O_2102,N_49788,N_49956);
or UO_2103 (O_2103,N_49915,N_49935);
nand UO_2104 (O_2104,N_49784,N_49957);
or UO_2105 (O_2105,N_49932,N_49874);
nand UO_2106 (O_2106,N_49902,N_49986);
nor UO_2107 (O_2107,N_49769,N_49884);
nor UO_2108 (O_2108,N_49987,N_49925);
and UO_2109 (O_2109,N_49913,N_49838);
or UO_2110 (O_2110,N_49768,N_49860);
and UO_2111 (O_2111,N_49825,N_49867);
nor UO_2112 (O_2112,N_49797,N_49959);
and UO_2113 (O_2113,N_49957,N_49985);
xor UO_2114 (O_2114,N_49772,N_49818);
nor UO_2115 (O_2115,N_49937,N_49792);
nor UO_2116 (O_2116,N_49895,N_49962);
xor UO_2117 (O_2117,N_49960,N_49943);
xnor UO_2118 (O_2118,N_49835,N_49845);
nor UO_2119 (O_2119,N_49899,N_49903);
and UO_2120 (O_2120,N_49772,N_49896);
nor UO_2121 (O_2121,N_49797,N_49964);
nand UO_2122 (O_2122,N_49889,N_49946);
or UO_2123 (O_2123,N_49952,N_49801);
nor UO_2124 (O_2124,N_49826,N_49865);
xnor UO_2125 (O_2125,N_49778,N_49933);
nand UO_2126 (O_2126,N_49919,N_49863);
xnor UO_2127 (O_2127,N_49862,N_49777);
xnor UO_2128 (O_2128,N_49764,N_49961);
nand UO_2129 (O_2129,N_49838,N_49882);
and UO_2130 (O_2130,N_49754,N_49831);
and UO_2131 (O_2131,N_49759,N_49933);
xnor UO_2132 (O_2132,N_49881,N_49921);
nor UO_2133 (O_2133,N_49779,N_49888);
or UO_2134 (O_2134,N_49763,N_49779);
nor UO_2135 (O_2135,N_49949,N_49922);
nand UO_2136 (O_2136,N_49953,N_49951);
xor UO_2137 (O_2137,N_49871,N_49862);
or UO_2138 (O_2138,N_49887,N_49892);
nor UO_2139 (O_2139,N_49972,N_49820);
nor UO_2140 (O_2140,N_49986,N_49755);
and UO_2141 (O_2141,N_49815,N_49839);
or UO_2142 (O_2142,N_49977,N_49888);
and UO_2143 (O_2143,N_49764,N_49777);
nand UO_2144 (O_2144,N_49860,N_49986);
and UO_2145 (O_2145,N_49776,N_49962);
or UO_2146 (O_2146,N_49922,N_49955);
or UO_2147 (O_2147,N_49866,N_49797);
xor UO_2148 (O_2148,N_49968,N_49888);
and UO_2149 (O_2149,N_49929,N_49891);
or UO_2150 (O_2150,N_49763,N_49877);
nor UO_2151 (O_2151,N_49763,N_49825);
or UO_2152 (O_2152,N_49956,N_49816);
xnor UO_2153 (O_2153,N_49925,N_49786);
nor UO_2154 (O_2154,N_49983,N_49933);
or UO_2155 (O_2155,N_49805,N_49799);
or UO_2156 (O_2156,N_49898,N_49875);
xor UO_2157 (O_2157,N_49913,N_49778);
xnor UO_2158 (O_2158,N_49977,N_49779);
nor UO_2159 (O_2159,N_49885,N_49819);
and UO_2160 (O_2160,N_49983,N_49871);
nand UO_2161 (O_2161,N_49894,N_49912);
nor UO_2162 (O_2162,N_49900,N_49971);
and UO_2163 (O_2163,N_49912,N_49954);
or UO_2164 (O_2164,N_49838,N_49797);
nand UO_2165 (O_2165,N_49814,N_49826);
nand UO_2166 (O_2166,N_49847,N_49827);
and UO_2167 (O_2167,N_49796,N_49752);
nand UO_2168 (O_2168,N_49757,N_49798);
and UO_2169 (O_2169,N_49843,N_49756);
nand UO_2170 (O_2170,N_49866,N_49832);
xor UO_2171 (O_2171,N_49759,N_49883);
xnor UO_2172 (O_2172,N_49756,N_49769);
xnor UO_2173 (O_2173,N_49855,N_49759);
or UO_2174 (O_2174,N_49764,N_49884);
nor UO_2175 (O_2175,N_49815,N_49958);
nand UO_2176 (O_2176,N_49839,N_49863);
or UO_2177 (O_2177,N_49789,N_49927);
xor UO_2178 (O_2178,N_49980,N_49826);
xnor UO_2179 (O_2179,N_49761,N_49939);
xor UO_2180 (O_2180,N_49799,N_49754);
and UO_2181 (O_2181,N_49800,N_49954);
xnor UO_2182 (O_2182,N_49820,N_49996);
nor UO_2183 (O_2183,N_49875,N_49888);
or UO_2184 (O_2184,N_49777,N_49840);
or UO_2185 (O_2185,N_49930,N_49926);
nor UO_2186 (O_2186,N_49837,N_49778);
xor UO_2187 (O_2187,N_49874,N_49821);
nand UO_2188 (O_2188,N_49864,N_49779);
xnor UO_2189 (O_2189,N_49793,N_49982);
nor UO_2190 (O_2190,N_49848,N_49907);
nand UO_2191 (O_2191,N_49985,N_49764);
and UO_2192 (O_2192,N_49892,N_49915);
nor UO_2193 (O_2193,N_49807,N_49869);
and UO_2194 (O_2194,N_49967,N_49866);
xnor UO_2195 (O_2195,N_49787,N_49872);
and UO_2196 (O_2196,N_49765,N_49834);
or UO_2197 (O_2197,N_49972,N_49875);
and UO_2198 (O_2198,N_49753,N_49988);
nor UO_2199 (O_2199,N_49935,N_49890);
and UO_2200 (O_2200,N_49942,N_49932);
and UO_2201 (O_2201,N_49880,N_49888);
and UO_2202 (O_2202,N_49753,N_49853);
and UO_2203 (O_2203,N_49782,N_49886);
or UO_2204 (O_2204,N_49936,N_49857);
nor UO_2205 (O_2205,N_49986,N_49806);
nand UO_2206 (O_2206,N_49917,N_49757);
and UO_2207 (O_2207,N_49773,N_49790);
and UO_2208 (O_2208,N_49768,N_49916);
and UO_2209 (O_2209,N_49767,N_49779);
nor UO_2210 (O_2210,N_49788,N_49781);
nor UO_2211 (O_2211,N_49781,N_49754);
nor UO_2212 (O_2212,N_49791,N_49946);
nor UO_2213 (O_2213,N_49799,N_49989);
xor UO_2214 (O_2214,N_49993,N_49939);
and UO_2215 (O_2215,N_49890,N_49785);
nor UO_2216 (O_2216,N_49991,N_49969);
or UO_2217 (O_2217,N_49917,N_49780);
nor UO_2218 (O_2218,N_49992,N_49831);
xnor UO_2219 (O_2219,N_49968,N_49958);
xnor UO_2220 (O_2220,N_49970,N_49995);
and UO_2221 (O_2221,N_49940,N_49918);
or UO_2222 (O_2222,N_49961,N_49928);
xor UO_2223 (O_2223,N_49987,N_49882);
or UO_2224 (O_2224,N_49956,N_49811);
and UO_2225 (O_2225,N_49794,N_49907);
nor UO_2226 (O_2226,N_49917,N_49989);
or UO_2227 (O_2227,N_49825,N_49762);
nand UO_2228 (O_2228,N_49975,N_49931);
nor UO_2229 (O_2229,N_49868,N_49898);
and UO_2230 (O_2230,N_49839,N_49986);
and UO_2231 (O_2231,N_49954,N_49862);
xnor UO_2232 (O_2232,N_49881,N_49773);
xnor UO_2233 (O_2233,N_49878,N_49846);
nor UO_2234 (O_2234,N_49913,N_49925);
xor UO_2235 (O_2235,N_49859,N_49843);
and UO_2236 (O_2236,N_49911,N_49778);
xor UO_2237 (O_2237,N_49949,N_49887);
and UO_2238 (O_2238,N_49859,N_49902);
and UO_2239 (O_2239,N_49913,N_49781);
nand UO_2240 (O_2240,N_49934,N_49985);
xor UO_2241 (O_2241,N_49880,N_49777);
xor UO_2242 (O_2242,N_49875,N_49923);
xor UO_2243 (O_2243,N_49983,N_49972);
xor UO_2244 (O_2244,N_49965,N_49760);
or UO_2245 (O_2245,N_49926,N_49752);
nand UO_2246 (O_2246,N_49968,N_49842);
or UO_2247 (O_2247,N_49871,N_49833);
nand UO_2248 (O_2248,N_49834,N_49887);
nor UO_2249 (O_2249,N_49814,N_49752);
nor UO_2250 (O_2250,N_49852,N_49855);
nand UO_2251 (O_2251,N_49750,N_49841);
or UO_2252 (O_2252,N_49971,N_49901);
xnor UO_2253 (O_2253,N_49751,N_49799);
nor UO_2254 (O_2254,N_49840,N_49951);
xor UO_2255 (O_2255,N_49945,N_49771);
and UO_2256 (O_2256,N_49846,N_49948);
and UO_2257 (O_2257,N_49759,N_49839);
nand UO_2258 (O_2258,N_49969,N_49984);
and UO_2259 (O_2259,N_49792,N_49932);
or UO_2260 (O_2260,N_49914,N_49846);
or UO_2261 (O_2261,N_49909,N_49877);
or UO_2262 (O_2262,N_49908,N_49936);
or UO_2263 (O_2263,N_49918,N_49877);
and UO_2264 (O_2264,N_49841,N_49945);
nor UO_2265 (O_2265,N_49791,N_49853);
nand UO_2266 (O_2266,N_49857,N_49860);
and UO_2267 (O_2267,N_49850,N_49938);
or UO_2268 (O_2268,N_49777,N_49999);
and UO_2269 (O_2269,N_49895,N_49845);
xor UO_2270 (O_2270,N_49914,N_49849);
or UO_2271 (O_2271,N_49975,N_49753);
nor UO_2272 (O_2272,N_49967,N_49788);
nand UO_2273 (O_2273,N_49909,N_49953);
or UO_2274 (O_2274,N_49870,N_49818);
nor UO_2275 (O_2275,N_49883,N_49984);
and UO_2276 (O_2276,N_49976,N_49939);
or UO_2277 (O_2277,N_49845,N_49943);
nor UO_2278 (O_2278,N_49991,N_49829);
xnor UO_2279 (O_2279,N_49849,N_49793);
nand UO_2280 (O_2280,N_49911,N_49782);
or UO_2281 (O_2281,N_49891,N_49768);
nor UO_2282 (O_2282,N_49894,N_49956);
or UO_2283 (O_2283,N_49755,N_49765);
nand UO_2284 (O_2284,N_49882,N_49962);
or UO_2285 (O_2285,N_49809,N_49768);
nor UO_2286 (O_2286,N_49972,N_49917);
nor UO_2287 (O_2287,N_49805,N_49968);
nand UO_2288 (O_2288,N_49840,N_49921);
and UO_2289 (O_2289,N_49999,N_49757);
and UO_2290 (O_2290,N_49795,N_49760);
nand UO_2291 (O_2291,N_49855,N_49796);
and UO_2292 (O_2292,N_49939,N_49790);
or UO_2293 (O_2293,N_49792,N_49914);
and UO_2294 (O_2294,N_49890,N_49940);
and UO_2295 (O_2295,N_49835,N_49785);
and UO_2296 (O_2296,N_49927,N_49832);
nor UO_2297 (O_2297,N_49764,N_49768);
or UO_2298 (O_2298,N_49775,N_49811);
xnor UO_2299 (O_2299,N_49843,N_49909);
or UO_2300 (O_2300,N_49937,N_49878);
nand UO_2301 (O_2301,N_49816,N_49899);
nand UO_2302 (O_2302,N_49781,N_49998);
nand UO_2303 (O_2303,N_49976,N_49872);
and UO_2304 (O_2304,N_49995,N_49823);
nand UO_2305 (O_2305,N_49959,N_49824);
nand UO_2306 (O_2306,N_49988,N_49991);
xnor UO_2307 (O_2307,N_49936,N_49881);
and UO_2308 (O_2308,N_49850,N_49805);
or UO_2309 (O_2309,N_49845,N_49873);
and UO_2310 (O_2310,N_49906,N_49918);
nand UO_2311 (O_2311,N_49934,N_49909);
and UO_2312 (O_2312,N_49779,N_49806);
nor UO_2313 (O_2313,N_49917,N_49928);
xnor UO_2314 (O_2314,N_49829,N_49807);
or UO_2315 (O_2315,N_49949,N_49971);
xnor UO_2316 (O_2316,N_49928,N_49786);
and UO_2317 (O_2317,N_49864,N_49763);
or UO_2318 (O_2318,N_49856,N_49985);
or UO_2319 (O_2319,N_49750,N_49809);
xor UO_2320 (O_2320,N_49871,N_49998);
and UO_2321 (O_2321,N_49852,N_49846);
nor UO_2322 (O_2322,N_49861,N_49977);
and UO_2323 (O_2323,N_49934,N_49825);
or UO_2324 (O_2324,N_49763,N_49837);
xnor UO_2325 (O_2325,N_49808,N_49791);
or UO_2326 (O_2326,N_49886,N_49934);
or UO_2327 (O_2327,N_49765,N_49784);
or UO_2328 (O_2328,N_49992,N_49766);
or UO_2329 (O_2329,N_49850,N_49841);
xnor UO_2330 (O_2330,N_49862,N_49806);
and UO_2331 (O_2331,N_49760,N_49882);
and UO_2332 (O_2332,N_49966,N_49956);
xnor UO_2333 (O_2333,N_49986,N_49834);
nor UO_2334 (O_2334,N_49973,N_49787);
and UO_2335 (O_2335,N_49963,N_49903);
and UO_2336 (O_2336,N_49897,N_49893);
nor UO_2337 (O_2337,N_49991,N_49951);
xnor UO_2338 (O_2338,N_49985,N_49989);
nand UO_2339 (O_2339,N_49975,N_49807);
or UO_2340 (O_2340,N_49894,N_49753);
or UO_2341 (O_2341,N_49913,N_49928);
and UO_2342 (O_2342,N_49859,N_49784);
and UO_2343 (O_2343,N_49986,N_49807);
nand UO_2344 (O_2344,N_49842,N_49921);
or UO_2345 (O_2345,N_49779,N_49760);
nand UO_2346 (O_2346,N_49897,N_49818);
nor UO_2347 (O_2347,N_49769,N_49818);
and UO_2348 (O_2348,N_49859,N_49974);
and UO_2349 (O_2349,N_49935,N_49842);
or UO_2350 (O_2350,N_49972,N_49831);
xor UO_2351 (O_2351,N_49812,N_49814);
and UO_2352 (O_2352,N_49833,N_49830);
and UO_2353 (O_2353,N_49873,N_49872);
nor UO_2354 (O_2354,N_49946,N_49798);
or UO_2355 (O_2355,N_49919,N_49968);
xnor UO_2356 (O_2356,N_49898,N_49809);
nor UO_2357 (O_2357,N_49839,N_49862);
or UO_2358 (O_2358,N_49898,N_49786);
nand UO_2359 (O_2359,N_49992,N_49811);
nand UO_2360 (O_2360,N_49766,N_49900);
xor UO_2361 (O_2361,N_49902,N_49823);
nor UO_2362 (O_2362,N_49779,N_49944);
nand UO_2363 (O_2363,N_49855,N_49857);
xor UO_2364 (O_2364,N_49834,N_49973);
or UO_2365 (O_2365,N_49952,N_49751);
and UO_2366 (O_2366,N_49781,N_49918);
nor UO_2367 (O_2367,N_49902,N_49970);
and UO_2368 (O_2368,N_49937,N_49942);
xor UO_2369 (O_2369,N_49895,N_49785);
nor UO_2370 (O_2370,N_49798,N_49755);
nand UO_2371 (O_2371,N_49868,N_49989);
or UO_2372 (O_2372,N_49933,N_49794);
xor UO_2373 (O_2373,N_49995,N_49772);
xor UO_2374 (O_2374,N_49770,N_49796);
nor UO_2375 (O_2375,N_49918,N_49978);
or UO_2376 (O_2376,N_49863,N_49993);
and UO_2377 (O_2377,N_49836,N_49872);
or UO_2378 (O_2378,N_49815,N_49939);
and UO_2379 (O_2379,N_49863,N_49804);
or UO_2380 (O_2380,N_49863,N_49755);
nor UO_2381 (O_2381,N_49991,N_49815);
xor UO_2382 (O_2382,N_49816,N_49891);
nand UO_2383 (O_2383,N_49796,N_49869);
nand UO_2384 (O_2384,N_49975,N_49894);
and UO_2385 (O_2385,N_49907,N_49755);
nand UO_2386 (O_2386,N_49976,N_49811);
nor UO_2387 (O_2387,N_49931,N_49780);
xor UO_2388 (O_2388,N_49768,N_49814);
and UO_2389 (O_2389,N_49979,N_49945);
or UO_2390 (O_2390,N_49806,N_49955);
or UO_2391 (O_2391,N_49822,N_49886);
nand UO_2392 (O_2392,N_49878,N_49884);
xnor UO_2393 (O_2393,N_49993,N_49841);
and UO_2394 (O_2394,N_49937,N_49999);
and UO_2395 (O_2395,N_49750,N_49985);
nor UO_2396 (O_2396,N_49940,N_49844);
or UO_2397 (O_2397,N_49989,N_49762);
and UO_2398 (O_2398,N_49840,N_49966);
nand UO_2399 (O_2399,N_49833,N_49784);
xor UO_2400 (O_2400,N_49803,N_49865);
xor UO_2401 (O_2401,N_49961,N_49935);
xnor UO_2402 (O_2402,N_49780,N_49790);
nor UO_2403 (O_2403,N_49833,N_49795);
nor UO_2404 (O_2404,N_49767,N_49878);
xor UO_2405 (O_2405,N_49987,N_49984);
nor UO_2406 (O_2406,N_49942,N_49896);
nand UO_2407 (O_2407,N_49914,N_49751);
xor UO_2408 (O_2408,N_49809,N_49946);
and UO_2409 (O_2409,N_49799,N_49926);
nor UO_2410 (O_2410,N_49856,N_49774);
nor UO_2411 (O_2411,N_49856,N_49959);
and UO_2412 (O_2412,N_49961,N_49970);
and UO_2413 (O_2413,N_49948,N_49794);
or UO_2414 (O_2414,N_49786,N_49796);
nand UO_2415 (O_2415,N_49985,N_49924);
nand UO_2416 (O_2416,N_49988,N_49894);
nor UO_2417 (O_2417,N_49857,N_49955);
xnor UO_2418 (O_2418,N_49940,N_49777);
and UO_2419 (O_2419,N_49851,N_49781);
nor UO_2420 (O_2420,N_49952,N_49905);
nor UO_2421 (O_2421,N_49870,N_49791);
and UO_2422 (O_2422,N_49923,N_49910);
nand UO_2423 (O_2423,N_49990,N_49928);
and UO_2424 (O_2424,N_49860,N_49962);
nand UO_2425 (O_2425,N_49865,N_49834);
or UO_2426 (O_2426,N_49950,N_49992);
nand UO_2427 (O_2427,N_49852,N_49812);
and UO_2428 (O_2428,N_49933,N_49860);
or UO_2429 (O_2429,N_49770,N_49847);
xnor UO_2430 (O_2430,N_49990,N_49778);
xnor UO_2431 (O_2431,N_49845,N_49769);
xor UO_2432 (O_2432,N_49867,N_49760);
or UO_2433 (O_2433,N_49866,N_49903);
xnor UO_2434 (O_2434,N_49765,N_49756);
nand UO_2435 (O_2435,N_49920,N_49902);
and UO_2436 (O_2436,N_49870,N_49961);
xnor UO_2437 (O_2437,N_49968,N_49981);
nand UO_2438 (O_2438,N_49781,N_49892);
and UO_2439 (O_2439,N_49886,N_49996);
xor UO_2440 (O_2440,N_49937,N_49991);
or UO_2441 (O_2441,N_49873,N_49886);
nor UO_2442 (O_2442,N_49848,N_49959);
nand UO_2443 (O_2443,N_49794,N_49913);
xnor UO_2444 (O_2444,N_49926,N_49834);
and UO_2445 (O_2445,N_49884,N_49906);
or UO_2446 (O_2446,N_49796,N_49795);
nor UO_2447 (O_2447,N_49957,N_49753);
and UO_2448 (O_2448,N_49852,N_49817);
and UO_2449 (O_2449,N_49972,N_49990);
xnor UO_2450 (O_2450,N_49803,N_49763);
xor UO_2451 (O_2451,N_49999,N_49765);
nor UO_2452 (O_2452,N_49802,N_49914);
xor UO_2453 (O_2453,N_49994,N_49851);
xnor UO_2454 (O_2454,N_49951,N_49943);
and UO_2455 (O_2455,N_49800,N_49926);
xor UO_2456 (O_2456,N_49898,N_49765);
nand UO_2457 (O_2457,N_49830,N_49934);
or UO_2458 (O_2458,N_49819,N_49792);
and UO_2459 (O_2459,N_49989,N_49778);
xor UO_2460 (O_2460,N_49937,N_49775);
or UO_2461 (O_2461,N_49934,N_49844);
and UO_2462 (O_2462,N_49956,N_49784);
and UO_2463 (O_2463,N_49918,N_49892);
nand UO_2464 (O_2464,N_49873,N_49918);
nor UO_2465 (O_2465,N_49780,N_49907);
nand UO_2466 (O_2466,N_49867,N_49946);
xor UO_2467 (O_2467,N_49923,N_49881);
and UO_2468 (O_2468,N_49835,N_49752);
nand UO_2469 (O_2469,N_49825,N_49928);
xnor UO_2470 (O_2470,N_49829,N_49816);
nor UO_2471 (O_2471,N_49951,N_49826);
or UO_2472 (O_2472,N_49871,N_49870);
or UO_2473 (O_2473,N_49973,N_49952);
nand UO_2474 (O_2474,N_49995,N_49860);
and UO_2475 (O_2475,N_49932,N_49803);
xnor UO_2476 (O_2476,N_49895,N_49992);
nor UO_2477 (O_2477,N_49930,N_49813);
nor UO_2478 (O_2478,N_49978,N_49809);
nor UO_2479 (O_2479,N_49778,N_49856);
nand UO_2480 (O_2480,N_49973,N_49844);
and UO_2481 (O_2481,N_49986,N_49983);
and UO_2482 (O_2482,N_49957,N_49987);
or UO_2483 (O_2483,N_49888,N_49990);
xnor UO_2484 (O_2484,N_49836,N_49771);
or UO_2485 (O_2485,N_49785,N_49921);
and UO_2486 (O_2486,N_49878,N_49967);
or UO_2487 (O_2487,N_49963,N_49832);
and UO_2488 (O_2488,N_49783,N_49985);
or UO_2489 (O_2489,N_49820,N_49925);
or UO_2490 (O_2490,N_49888,N_49753);
nor UO_2491 (O_2491,N_49883,N_49953);
xnor UO_2492 (O_2492,N_49964,N_49782);
and UO_2493 (O_2493,N_49917,N_49991);
nor UO_2494 (O_2494,N_49803,N_49940);
and UO_2495 (O_2495,N_49927,N_49977);
nand UO_2496 (O_2496,N_49784,N_49998);
xor UO_2497 (O_2497,N_49889,N_49792);
or UO_2498 (O_2498,N_49862,N_49791);
or UO_2499 (O_2499,N_49995,N_49933);
nor UO_2500 (O_2500,N_49784,N_49796);
and UO_2501 (O_2501,N_49853,N_49860);
nor UO_2502 (O_2502,N_49973,N_49823);
or UO_2503 (O_2503,N_49966,N_49979);
xor UO_2504 (O_2504,N_49791,N_49913);
xor UO_2505 (O_2505,N_49962,N_49995);
or UO_2506 (O_2506,N_49880,N_49798);
xnor UO_2507 (O_2507,N_49958,N_49804);
xnor UO_2508 (O_2508,N_49750,N_49772);
and UO_2509 (O_2509,N_49968,N_49776);
nand UO_2510 (O_2510,N_49983,N_49861);
and UO_2511 (O_2511,N_49875,N_49931);
nand UO_2512 (O_2512,N_49826,N_49854);
or UO_2513 (O_2513,N_49838,N_49769);
or UO_2514 (O_2514,N_49991,N_49958);
nand UO_2515 (O_2515,N_49763,N_49790);
or UO_2516 (O_2516,N_49969,N_49947);
or UO_2517 (O_2517,N_49759,N_49819);
xnor UO_2518 (O_2518,N_49793,N_49756);
nor UO_2519 (O_2519,N_49904,N_49952);
and UO_2520 (O_2520,N_49783,N_49789);
nand UO_2521 (O_2521,N_49957,N_49851);
xnor UO_2522 (O_2522,N_49840,N_49916);
nand UO_2523 (O_2523,N_49862,N_49794);
or UO_2524 (O_2524,N_49877,N_49890);
and UO_2525 (O_2525,N_49821,N_49823);
nor UO_2526 (O_2526,N_49968,N_49895);
nand UO_2527 (O_2527,N_49949,N_49798);
nor UO_2528 (O_2528,N_49788,N_49828);
or UO_2529 (O_2529,N_49967,N_49834);
nand UO_2530 (O_2530,N_49824,N_49751);
nor UO_2531 (O_2531,N_49975,N_49769);
xor UO_2532 (O_2532,N_49854,N_49953);
or UO_2533 (O_2533,N_49991,N_49858);
or UO_2534 (O_2534,N_49992,N_49915);
nand UO_2535 (O_2535,N_49996,N_49962);
or UO_2536 (O_2536,N_49982,N_49909);
nor UO_2537 (O_2537,N_49753,N_49902);
and UO_2538 (O_2538,N_49870,N_49860);
or UO_2539 (O_2539,N_49893,N_49835);
and UO_2540 (O_2540,N_49905,N_49957);
and UO_2541 (O_2541,N_49806,N_49861);
xnor UO_2542 (O_2542,N_49847,N_49839);
nand UO_2543 (O_2543,N_49946,N_49912);
and UO_2544 (O_2544,N_49756,N_49833);
and UO_2545 (O_2545,N_49884,N_49990);
or UO_2546 (O_2546,N_49954,N_49895);
or UO_2547 (O_2547,N_49846,N_49913);
xor UO_2548 (O_2548,N_49856,N_49835);
nor UO_2549 (O_2549,N_49782,N_49816);
nand UO_2550 (O_2550,N_49789,N_49961);
nor UO_2551 (O_2551,N_49755,N_49868);
xnor UO_2552 (O_2552,N_49840,N_49965);
nand UO_2553 (O_2553,N_49750,N_49932);
xor UO_2554 (O_2554,N_49960,N_49763);
or UO_2555 (O_2555,N_49762,N_49933);
or UO_2556 (O_2556,N_49821,N_49777);
nor UO_2557 (O_2557,N_49898,N_49950);
xor UO_2558 (O_2558,N_49955,N_49885);
nor UO_2559 (O_2559,N_49897,N_49798);
or UO_2560 (O_2560,N_49863,N_49837);
nor UO_2561 (O_2561,N_49906,N_49988);
nand UO_2562 (O_2562,N_49839,N_49959);
or UO_2563 (O_2563,N_49784,N_49911);
nand UO_2564 (O_2564,N_49895,N_49955);
nor UO_2565 (O_2565,N_49894,N_49846);
or UO_2566 (O_2566,N_49981,N_49937);
and UO_2567 (O_2567,N_49767,N_49816);
nand UO_2568 (O_2568,N_49937,N_49986);
nor UO_2569 (O_2569,N_49925,N_49982);
nand UO_2570 (O_2570,N_49980,N_49813);
nand UO_2571 (O_2571,N_49868,N_49994);
or UO_2572 (O_2572,N_49863,N_49881);
and UO_2573 (O_2573,N_49879,N_49921);
nand UO_2574 (O_2574,N_49762,N_49924);
xor UO_2575 (O_2575,N_49854,N_49885);
nand UO_2576 (O_2576,N_49807,N_49791);
and UO_2577 (O_2577,N_49893,N_49996);
and UO_2578 (O_2578,N_49828,N_49795);
nor UO_2579 (O_2579,N_49815,N_49954);
or UO_2580 (O_2580,N_49906,N_49787);
nor UO_2581 (O_2581,N_49806,N_49924);
and UO_2582 (O_2582,N_49928,N_49779);
xnor UO_2583 (O_2583,N_49756,N_49878);
and UO_2584 (O_2584,N_49907,N_49954);
xnor UO_2585 (O_2585,N_49978,N_49895);
xnor UO_2586 (O_2586,N_49969,N_49810);
nand UO_2587 (O_2587,N_49897,N_49995);
or UO_2588 (O_2588,N_49995,N_49928);
nor UO_2589 (O_2589,N_49864,N_49824);
nand UO_2590 (O_2590,N_49969,N_49895);
xor UO_2591 (O_2591,N_49861,N_49826);
nor UO_2592 (O_2592,N_49797,N_49850);
or UO_2593 (O_2593,N_49973,N_49989);
xnor UO_2594 (O_2594,N_49893,N_49775);
or UO_2595 (O_2595,N_49987,N_49816);
nand UO_2596 (O_2596,N_49896,N_49902);
and UO_2597 (O_2597,N_49869,N_49913);
and UO_2598 (O_2598,N_49970,N_49998);
or UO_2599 (O_2599,N_49879,N_49915);
xor UO_2600 (O_2600,N_49790,N_49883);
and UO_2601 (O_2601,N_49952,N_49993);
or UO_2602 (O_2602,N_49813,N_49943);
nand UO_2603 (O_2603,N_49914,N_49997);
and UO_2604 (O_2604,N_49777,N_49919);
nor UO_2605 (O_2605,N_49985,N_49860);
nor UO_2606 (O_2606,N_49975,N_49883);
nand UO_2607 (O_2607,N_49777,N_49794);
and UO_2608 (O_2608,N_49840,N_49845);
and UO_2609 (O_2609,N_49987,N_49783);
nand UO_2610 (O_2610,N_49752,N_49893);
nand UO_2611 (O_2611,N_49877,N_49839);
and UO_2612 (O_2612,N_49827,N_49982);
and UO_2613 (O_2613,N_49780,N_49924);
nor UO_2614 (O_2614,N_49867,N_49936);
nand UO_2615 (O_2615,N_49869,N_49929);
or UO_2616 (O_2616,N_49952,N_49838);
or UO_2617 (O_2617,N_49942,N_49941);
or UO_2618 (O_2618,N_49915,N_49761);
nor UO_2619 (O_2619,N_49958,N_49783);
and UO_2620 (O_2620,N_49904,N_49983);
xnor UO_2621 (O_2621,N_49868,N_49859);
xor UO_2622 (O_2622,N_49896,N_49805);
nor UO_2623 (O_2623,N_49868,N_49996);
nor UO_2624 (O_2624,N_49984,N_49885);
nor UO_2625 (O_2625,N_49955,N_49954);
and UO_2626 (O_2626,N_49789,N_49910);
xor UO_2627 (O_2627,N_49783,N_49865);
xnor UO_2628 (O_2628,N_49985,N_49977);
nor UO_2629 (O_2629,N_49963,N_49783);
nor UO_2630 (O_2630,N_49967,N_49756);
xor UO_2631 (O_2631,N_49913,N_49786);
nor UO_2632 (O_2632,N_49827,N_49871);
nand UO_2633 (O_2633,N_49871,N_49963);
nor UO_2634 (O_2634,N_49795,N_49765);
nand UO_2635 (O_2635,N_49859,N_49856);
nor UO_2636 (O_2636,N_49892,N_49914);
nand UO_2637 (O_2637,N_49967,N_49910);
xor UO_2638 (O_2638,N_49780,N_49750);
xor UO_2639 (O_2639,N_49786,N_49815);
xnor UO_2640 (O_2640,N_49801,N_49943);
nand UO_2641 (O_2641,N_49826,N_49888);
nand UO_2642 (O_2642,N_49839,N_49752);
nor UO_2643 (O_2643,N_49815,N_49876);
xor UO_2644 (O_2644,N_49945,N_49854);
nand UO_2645 (O_2645,N_49883,N_49832);
nor UO_2646 (O_2646,N_49788,N_49834);
nor UO_2647 (O_2647,N_49797,N_49928);
and UO_2648 (O_2648,N_49833,N_49824);
nand UO_2649 (O_2649,N_49885,N_49948);
nor UO_2650 (O_2650,N_49942,N_49966);
nand UO_2651 (O_2651,N_49913,N_49999);
nand UO_2652 (O_2652,N_49800,N_49996);
nor UO_2653 (O_2653,N_49978,N_49774);
or UO_2654 (O_2654,N_49999,N_49961);
or UO_2655 (O_2655,N_49804,N_49908);
nor UO_2656 (O_2656,N_49909,N_49836);
nor UO_2657 (O_2657,N_49850,N_49836);
nand UO_2658 (O_2658,N_49860,N_49921);
nor UO_2659 (O_2659,N_49992,N_49819);
or UO_2660 (O_2660,N_49933,N_49826);
nor UO_2661 (O_2661,N_49879,N_49971);
and UO_2662 (O_2662,N_49982,N_49802);
xnor UO_2663 (O_2663,N_49842,N_49901);
and UO_2664 (O_2664,N_49923,N_49800);
nand UO_2665 (O_2665,N_49906,N_49848);
and UO_2666 (O_2666,N_49911,N_49758);
nand UO_2667 (O_2667,N_49831,N_49919);
nand UO_2668 (O_2668,N_49803,N_49999);
or UO_2669 (O_2669,N_49910,N_49776);
or UO_2670 (O_2670,N_49820,N_49761);
nand UO_2671 (O_2671,N_49878,N_49998);
nand UO_2672 (O_2672,N_49969,N_49836);
and UO_2673 (O_2673,N_49846,N_49756);
or UO_2674 (O_2674,N_49970,N_49765);
or UO_2675 (O_2675,N_49829,N_49952);
nand UO_2676 (O_2676,N_49997,N_49823);
or UO_2677 (O_2677,N_49788,N_49995);
or UO_2678 (O_2678,N_49801,N_49807);
nand UO_2679 (O_2679,N_49858,N_49832);
xor UO_2680 (O_2680,N_49855,N_49928);
xor UO_2681 (O_2681,N_49778,N_49970);
xor UO_2682 (O_2682,N_49758,N_49856);
or UO_2683 (O_2683,N_49840,N_49876);
xor UO_2684 (O_2684,N_49958,N_49763);
and UO_2685 (O_2685,N_49909,N_49901);
nand UO_2686 (O_2686,N_49879,N_49922);
and UO_2687 (O_2687,N_49865,N_49847);
and UO_2688 (O_2688,N_49948,N_49966);
and UO_2689 (O_2689,N_49830,N_49836);
nor UO_2690 (O_2690,N_49802,N_49930);
nor UO_2691 (O_2691,N_49986,N_49843);
and UO_2692 (O_2692,N_49895,N_49975);
and UO_2693 (O_2693,N_49960,N_49958);
and UO_2694 (O_2694,N_49934,N_49868);
nand UO_2695 (O_2695,N_49972,N_49764);
xnor UO_2696 (O_2696,N_49880,N_49800);
nor UO_2697 (O_2697,N_49755,N_49968);
or UO_2698 (O_2698,N_49793,N_49900);
xnor UO_2699 (O_2699,N_49965,N_49870);
xnor UO_2700 (O_2700,N_49875,N_49816);
and UO_2701 (O_2701,N_49801,N_49776);
or UO_2702 (O_2702,N_49930,N_49968);
nand UO_2703 (O_2703,N_49909,N_49921);
xnor UO_2704 (O_2704,N_49976,N_49926);
xor UO_2705 (O_2705,N_49933,N_49924);
nor UO_2706 (O_2706,N_49921,N_49837);
xor UO_2707 (O_2707,N_49927,N_49855);
nor UO_2708 (O_2708,N_49988,N_49921);
and UO_2709 (O_2709,N_49769,N_49750);
and UO_2710 (O_2710,N_49959,N_49813);
nand UO_2711 (O_2711,N_49794,N_49798);
and UO_2712 (O_2712,N_49847,N_49866);
xor UO_2713 (O_2713,N_49912,N_49798);
nor UO_2714 (O_2714,N_49799,N_49795);
xor UO_2715 (O_2715,N_49901,N_49792);
nand UO_2716 (O_2716,N_49831,N_49878);
xnor UO_2717 (O_2717,N_49968,N_49821);
nor UO_2718 (O_2718,N_49795,N_49910);
nand UO_2719 (O_2719,N_49941,N_49806);
or UO_2720 (O_2720,N_49816,N_49995);
nand UO_2721 (O_2721,N_49935,N_49804);
and UO_2722 (O_2722,N_49891,N_49827);
xor UO_2723 (O_2723,N_49918,N_49871);
xor UO_2724 (O_2724,N_49975,N_49911);
or UO_2725 (O_2725,N_49959,N_49782);
or UO_2726 (O_2726,N_49754,N_49777);
and UO_2727 (O_2727,N_49970,N_49844);
xor UO_2728 (O_2728,N_49999,N_49889);
and UO_2729 (O_2729,N_49910,N_49840);
xor UO_2730 (O_2730,N_49963,N_49756);
nand UO_2731 (O_2731,N_49894,N_49971);
nor UO_2732 (O_2732,N_49877,N_49885);
nor UO_2733 (O_2733,N_49990,N_49804);
or UO_2734 (O_2734,N_49799,N_49829);
nor UO_2735 (O_2735,N_49778,N_49974);
nor UO_2736 (O_2736,N_49963,N_49861);
nand UO_2737 (O_2737,N_49775,N_49935);
xnor UO_2738 (O_2738,N_49936,N_49938);
or UO_2739 (O_2739,N_49825,N_49949);
or UO_2740 (O_2740,N_49865,N_49753);
or UO_2741 (O_2741,N_49753,N_49956);
nor UO_2742 (O_2742,N_49838,N_49865);
nor UO_2743 (O_2743,N_49924,N_49859);
or UO_2744 (O_2744,N_49958,N_49893);
and UO_2745 (O_2745,N_49816,N_49846);
xnor UO_2746 (O_2746,N_49984,N_49832);
or UO_2747 (O_2747,N_49880,N_49917);
or UO_2748 (O_2748,N_49836,N_49766);
or UO_2749 (O_2749,N_49861,N_49894);
xnor UO_2750 (O_2750,N_49920,N_49759);
or UO_2751 (O_2751,N_49850,N_49940);
nor UO_2752 (O_2752,N_49948,N_49972);
and UO_2753 (O_2753,N_49802,N_49770);
xor UO_2754 (O_2754,N_49852,N_49932);
xor UO_2755 (O_2755,N_49977,N_49788);
nand UO_2756 (O_2756,N_49885,N_49797);
nand UO_2757 (O_2757,N_49779,N_49859);
and UO_2758 (O_2758,N_49783,N_49808);
or UO_2759 (O_2759,N_49994,N_49943);
nand UO_2760 (O_2760,N_49817,N_49881);
nor UO_2761 (O_2761,N_49882,N_49972);
nor UO_2762 (O_2762,N_49854,N_49968);
nand UO_2763 (O_2763,N_49975,N_49884);
nor UO_2764 (O_2764,N_49934,N_49803);
nor UO_2765 (O_2765,N_49833,N_49835);
xor UO_2766 (O_2766,N_49784,N_49834);
nand UO_2767 (O_2767,N_49866,N_49933);
or UO_2768 (O_2768,N_49991,N_49822);
nand UO_2769 (O_2769,N_49805,N_49908);
and UO_2770 (O_2770,N_49892,N_49880);
and UO_2771 (O_2771,N_49831,N_49990);
nand UO_2772 (O_2772,N_49955,N_49984);
nand UO_2773 (O_2773,N_49860,N_49972);
and UO_2774 (O_2774,N_49987,N_49976);
nand UO_2775 (O_2775,N_49892,N_49934);
and UO_2776 (O_2776,N_49901,N_49917);
nor UO_2777 (O_2777,N_49919,N_49984);
nand UO_2778 (O_2778,N_49951,N_49809);
or UO_2779 (O_2779,N_49787,N_49776);
nor UO_2780 (O_2780,N_49806,N_49919);
nor UO_2781 (O_2781,N_49999,N_49947);
nor UO_2782 (O_2782,N_49755,N_49985);
xor UO_2783 (O_2783,N_49765,N_49863);
and UO_2784 (O_2784,N_49993,N_49798);
or UO_2785 (O_2785,N_49850,N_49918);
or UO_2786 (O_2786,N_49967,N_49808);
and UO_2787 (O_2787,N_49924,N_49955);
and UO_2788 (O_2788,N_49993,N_49870);
nor UO_2789 (O_2789,N_49970,N_49996);
xor UO_2790 (O_2790,N_49914,N_49770);
and UO_2791 (O_2791,N_49765,N_49817);
xor UO_2792 (O_2792,N_49804,N_49865);
xor UO_2793 (O_2793,N_49823,N_49814);
nand UO_2794 (O_2794,N_49769,N_49770);
xnor UO_2795 (O_2795,N_49922,N_49934);
or UO_2796 (O_2796,N_49945,N_49813);
nor UO_2797 (O_2797,N_49824,N_49932);
xnor UO_2798 (O_2798,N_49994,N_49896);
or UO_2799 (O_2799,N_49825,N_49984);
nor UO_2800 (O_2800,N_49823,N_49948);
nor UO_2801 (O_2801,N_49773,N_49975);
nand UO_2802 (O_2802,N_49976,N_49955);
and UO_2803 (O_2803,N_49985,N_49873);
and UO_2804 (O_2804,N_49897,N_49920);
xnor UO_2805 (O_2805,N_49970,N_49882);
and UO_2806 (O_2806,N_49827,N_49856);
or UO_2807 (O_2807,N_49828,N_49928);
and UO_2808 (O_2808,N_49915,N_49773);
or UO_2809 (O_2809,N_49841,N_49867);
xnor UO_2810 (O_2810,N_49975,N_49984);
nor UO_2811 (O_2811,N_49885,N_49881);
or UO_2812 (O_2812,N_49947,N_49844);
or UO_2813 (O_2813,N_49960,N_49999);
or UO_2814 (O_2814,N_49960,N_49764);
or UO_2815 (O_2815,N_49868,N_49987);
nand UO_2816 (O_2816,N_49931,N_49997);
and UO_2817 (O_2817,N_49759,N_49887);
nand UO_2818 (O_2818,N_49984,N_49874);
or UO_2819 (O_2819,N_49869,N_49820);
nor UO_2820 (O_2820,N_49957,N_49946);
or UO_2821 (O_2821,N_49810,N_49905);
xor UO_2822 (O_2822,N_49863,N_49851);
xor UO_2823 (O_2823,N_49852,N_49824);
nand UO_2824 (O_2824,N_49909,N_49831);
xnor UO_2825 (O_2825,N_49918,N_49843);
or UO_2826 (O_2826,N_49804,N_49836);
or UO_2827 (O_2827,N_49888,N_49952);
nand UO_2828 (O_2828,N_49785,N_49787);
xor UO_2829 (O_2829,N_49856,N_49928);
nor UO_2830 (O_2830,N_49981,N_49771);
or UO_2831 (O_2831,N_49884,N_49845);
nand UO_2832 (O_2832,N_49987,N_49870);
nor UO_2833 (O_2833,N_49929,N_49917);
nor UO_2834 (O_2834,N_49770,N_49919);
nand UO_2835 (O_2835,N_49890,N_49983);
xor UO_2836 (O_2836,N_49755,N_49997);
and UO_2837 (O_2837,N_49993,N_49905);
or UO_2838 (O_2838,N_49956,N_49885);
and UO_2839 (O_2839,N_49798,N_49788);
nand UO_2840 (O_2840,N_49978,N_49987);
nor UO_2841 (O_2841,N_49918,N_49759);
or UO_2842 (O_2842,N_49758,N_49810);
nand UO_2843 (O_2843,N_49998,N_49989);
xor UO_2844 (O_2844,N_49847,N_49750);
and UO_2845 (O_2845,N_49924,N_49853);
or UO_2846 (O_2846,N_49998,N_49965);
xor UO_2847 (O_2847,N_49827,N_49798);
xor UO_2848 (O_2848,N_49816,N_49831);
nand UO_2849 (O_2849,N_49773,N_49947);
nor UO_2850 (O_2850,N_49945,N_49876);
xnor UO_2851 (O_2851,N_49793,N_49995);
nor UO_2852 (O_2852,N_49880,N_49881);
nand UO_2853 (O_2853,N_49858,N_49923);
nor UO_2854 (O_2854,N_49852,N_49971);
nor UO_2855 (O_2855,N_49920,N_49901);
or UO_2856 (O_2856,N_49952,N_49922);
xor UO_2857 (O_2857,N_49763,N_49811);
xnor UO_2858 (O_2858,N_49752,N_49875);
or UO_2859 (O_2859,N_49763,N_49766);
nor UO_2860 (O_2860,N_49773,N_49899);
xnor UO_2861 (O_2861,N_49820,N_49785);
and UO_2862 (O_2862,N_49864,N_49764);
and UO_2863 (O_2863,N_49987,N_49808);
nor UO_2864 (O_2864,N_49977,N_49878);
nor UO_2865 (O_2865,N_49766,N_49842);
and UO_2866 (O_2866,N_49894,N_49895);
or UO_2867 (O_2867,N_49869,N_49924);
and UO_2868 (O_2868,N_49955,N_49859);
nand UO_2869 (O_2869,N_49982,N_49886);
or UO_2870 (O_2870,N_49910,N_49940);
or UO_2871 (O_2871,N_49891,N_49893);
or UO_2872 (O_2872,N_49842,N_49810);
xnor UO_2873 (O_2873,N_49983,N_49923);
and UO_2874 (O_2874,N_49885,N_49880);
nor UO_2875 (O_2875,N_49972,N_49980);
nand UO_2876 (O_2876,N_49900,N_49760);
and UO_2877 (O_2877,N_49750,N_49868);
nand UO_2878 (O_2878,N_49830,N_49997);
nand UO_2879 (O_2879,N_49969,N_49811);
nor UO_2880 (O_2880,N_49814,N_49907);
or UO_2881 (O_2881,N_49750,N_49836);
nand UO_2882 (O_2882,N_49750,N_49885);
nor UO_2883 (O_2883,N_49866,N_49751);
or UO_2884 (O_2884,N_49826,N_49813);
xnor UO_2885 (O_2885,N_49945,N_49987);
and UO_2886 (O_2886,N_49899,N_49895);
xor UO_2887 (O_2887,N_49803,N_49872);
and UO_2888 (O_2888,N_49877,N_49832);
or UO_2889 (O_2889,N_49936,N_49947);
nor UO_2890 (O_2890,N_49934,N_49959);
nor UO_2891 (O_2891,N_49978,N_49973);
nand UO_2892 (O_2892,N_49858,N_49813);
or UO_2893 (O_2893,N_49972,N_49977);
or UO_2894 (O_2894,N_49800,N_49770);
nand UO_2895 (O_2895,N_49871,N_49834);
nor UO_2896 (O_2896,N_49924,N_49760);
or UO_2897 (O_2897,N_49903,N_49779);
nor UO_2898 (O_2898,N_49782,N_49914);
nand UO_2899 (O_2899,N_49857,N_49889);
nor UO_2900 (O_2900,N_49768,N_49950);
nand UO_2901 (O_2901,N_49807,N_49753);
nor UO_2902 (O_2902,N_49817,N_49962);
and UO_2903 (O_2903,N_49767,N_49937);
nand UO_2904 (O_2904,N_49923,N_49960);
and UO_2905 (O_2905,N_49923,N_49806);
nand UO_2906 (O_2906,N_49934,N_49967);
nor UO_2907 (O_2907,N_49785,N_49751);
xor UO_2908 (O_2908,N_49997,N_49983);
and UO_2909 (O_2909,N_49873,N_49993);
xnor UO_2910 (O_2910,N_49990,N_49909);
and UO_2911 (O_2911,N_49860,N_49988);
nor UO_2912 (O_2912,N_49950,N_49834);
and UO_2913 (O_2913,N_49863,N_49831);
or UO_2914 (O_2914,N_49998,N_49898);
nand UO_2915 (O_2915,N_49865,N_49819);
and UO_2916 (O_2916,N_49979,N_49779);
or UO_2917 (O_2917,N_49807,N_49757);
nor UO_2918 (O_2918,N_49762,N_49761);
nor UO_2919 (O_2919,N_49944,N_49988);
nand UO_2920 (O_2920,N_49808,N_49819);
and UO_2921 (O_2921,N_49993,N_49914);
and UO_2922 (O_2922,N_49997,N_49833);
and UO_2923 (O_2923,N_49977,N_49986);
nor UO_2924 (O_2924,N_49954,N_49971);
nand UO_2925 (O_2925,N_49972,N_49798);
nand UO_2926 (O_2926,N_49777,N_49781);
nand UO_2927 (O_2927,N_49766,N_49981);
or UO_2928 (O_2928,N_49999,N_49948);
xor UO_2929 (O_2929,N_49879,N_49894);
and UO_2930 (O_2930,N_49873,N_49978);
xor UO_2931 (O_2931,N_49958,N_49925);
nor UO_2932 (O_2932,N_49823,N_49888);
nand UO_2933 (O_2933,N_49829,N_49883);
nand UO_2934 (O_2934,N_49790,N_49912);
or UO_2935 (O_2935,N_49864,N_49794);
xnor UO_2936 (O_2936,N_49984,N_49994);
nand UO_2937 (O_2937,N_49755,N_49864);
and UO_2938 (O_2938,N_49876,N_49894);
nand UO_2939 (O_2939,N_49960,N_49787);
and UO_2940 (O_2940,N_49884,N_49920);
or UO_2941 (O_2941,N_49898,N_49988);
and UO_2942 (O_2942,N_49996,N_49775);
nand UO_2943 (O_2943,N_49990,N_49975);
and UO_2944 (O_2944,N_49968,N_49890);
nor UO_2945 (O_2945,N_49837,N_49959);
nor UO_2946 (O_2946,N_49892,N_49787);
or UO_2947 (O_2947,N_49877,N_49953);
xnor UO_2948 (O_2948,N_49844,N_49771);
nor UO_2949 (O_2949,N_49974,N_49793);
and UO_2950 (O_2950,N_49994,N_49887);
nor UO_2951 (O_2951,N_49940,N_49775);
nor UO_2952 (O_2952,N_49990,N_49993);
nand UO_2953 (O_2953,N_49952,N_49885);
or UO_2954 (O_2954,N_49820,N_49799);
nor UO_2955 (O_2955,N_49991,N_49850);
nand UO_2956 (O_2956,N_49880,N_49770);
and UO_2957 (O_2957,N_49838,N_49811);
or UO_2958 (O_2958,N_49916,N_49887);
xnor UO_2959 (O_2959,N_49808,N_49920);
nand UO_2960 (O_2960,N_49813,N_49973);
and UO_2961 (O_2961,N_49830,N_49924);
and UO_2962 (O_2962,N_49958,N_49758);
nor UO_2963 (O_2963,N_49970,N_49897);
nor UO_2964 (O_2964,N_49966,N_49936);
xor UO_2965 (O_2965,N_49862,N_49935);
nor UO_2966 (O_2966,N_49775,N_49836);
or UO_2967 (O_2967,N_49930,N_49804);
and UO_2968 (O_2968,N_49806,N_49829);
and UO_2969 (O_2969,N_49785,N_49984);
nor UO_2970 (O_2970,N_49839,N_49817);
nor UO_2971 (O_2971,N_49810,N_49851);
xor UO_2972 (O_2972,N_49942,N_49864);
xnor UO_2973 (O_2973,N_49758,N_49947);
or UO_2974 (O_2974,N_49936,N_49999);
or UO_2975 (O_2975,N_49890,N_49897);
xor UO_2976 (O_2976,N_49980,N_49938);
nand UO_2977 (O_2977,N_49916,N_49752);
xor UO_2978 (O_2978,N_49843,N_49898);
nor UO_2979 (O_2979,N_49907,N_49779);
xnor UO_2980 (O_2980,N_49826,N_49945);
or UO_2981 (O_2981,N_49997,N_49763);
nand UO_2982 (O_2982,N_49977,N_49992);
nor UO_2983 (O_2983,N_49806,N_49906);
or UO_2984 (O_2984,N_49999,N_49771);
xor UO_2985 (O_2985,N_49814,N_49784);
nor UO_2986 (O_2986,N_49775,N_49953);
and UO_2987 (O_2987,N_49838,N_49963);
or UO_2988 (O_2988,N_49859,N_49892);
or UO_2989 (O_2989,N_49972,N_49781);
or UO_2990 (O_2990,N_49943,N_49921);
nor UO_2991 (O_2991,N_49950,N_49853);
and UO_2992 (O_2992,N_49949,N_49849);
or UO_2993 (O_2993,N_49924,N_49989);
and UO_2994 (O_2994,N_49902,N_49906);
nand UO_2995 (O_2995,N_49825,N_49808);
nor UO_2996 (O_2996,N_49985,N_49876);
or UO_2997 (O_2997,N_49831,N_49963);
or UO_2998 (O_2998,N_49827,N_49963);
xor UO_2999 (O_2999,N_49809,N_49802);
and UO_3000 (O_3000,N_49798,N_49899);
xor UO_3001 (O_3001,N_49925,N_49965);
xor UO_3002 (O_3002,N_49918,N_49957);
nand UO_3003 (O_3003,N_49853,N_49750);
xnor UO_3004 (O_3004,N_49908,N_49935);
nand UO_3005 (O_3005,N_49820,N_49823);
nand UO_3006 (O_3006,N_49775,N_49847);
and UO_3007 (O_3007,N_49828,N_49856);
nor UO_3008 (O_3008,N_49929,N_49848);
or UO_3009 (O_3009,N_49939,N_49890);
xor UO_3010 (O_3010,N_49896,N_49949);
nand UO_3011 (O_3011,N_49887,N_49977);
nand UO_3012 (O_3012,N_49814,N_49762);
nor UO_3013 (O_3013,N_49992,N_49753);
nand UO_3014 (O_3014,N_49913,N_49949);
xnor UO_3015 (O_3015,N_49880,N_49898);
or UO_3016 (O_3016,N_49840,N_49925);
nor UO_3017 (O_3017,N_49869,N_49859);
nor UO_3018 (O_3018,N_49773,N_49787);
or UO_3019 (O_3019,N_49996,N_49759);
nand UO_3020 (O_3020,N_49845,N_49813);
nor UO_3021 (O_3021,N_49971,N_49840);
nor UO_3022 (O_3022,N_49817,N_49847);
nand UO_3023 (O_3023,N_49974,N_49819);
or UO_3024 (O_3024,N_49937,N_49754);
nand UO_3025 (O_3025,N_49957,N_49917);
xor UO_3026 (O_3026,N_49813,N_49933);
xor UO_3027 (O_3027,N_49940,N_49780);
and UO_3028 (O_3028,N_49855,N_49924);
and UO_3029 (O_3029,N_49982,N_49910);
or UO_3030 (O_3030,N_49827,N_49756);
and UO_3031 (O_3031,N_49921,N_49877);
nor UO_3032 (O_3032,N_49926,N_49969);
nor UO_3033 (O_3033,N_49820,N_49924);
xnor UO_3034 (O_3034,N_49796,N_49939);
xor UO_3035 (O_3035,N_49794,N_49811);
nor UO_3036 (O_3036,N_49974,N_49795);
xor UO_3037 (O_3037,N_49908,N_49959);
and UO_3038 (O_3038,N_49869,N_49916);
xor UO_3039 (O_3039,N_49843,N_49853);
and UO_3040 (O_3040,N_49966,N_49960);
and UO_3041 (O_3041,N_49843,N_49897);
nor UO_3042 (O_3042,N_49814,N_49886);
xnor UO_3043 (O_3043,N_49970,N_49898);
nand UO_3044 (O_3044,N_49874,N_49944);
and UO_3045 (O_3045,N_49881,N_49901);
nand UO_3046 (O_3046,N_49931,N_49798);
or UO_3047 (O_3047,N_49859,N_49796);
nand UO_3048 (O_3048,N_49789,N_49854);
nand UO_3049 (O_3049,N_49770,N_49929);
xor UO_3050 (O_3050,N_49960,N_49869);
nand UO_3051 (O_3051,N_49928,N_49887);
xnor UO_3052 (O_3052,N_49941,N_49816);
and UO_3053 (O_3053,N_49769,N_49821);
or UO_3054 (O_3054,N_49855,N_49961);
nand UO_3055 (O_3055,N_49859,N_49911);
xnor UO_3056 (O_3056,N_49948,N_49933);
and UO_3057 (O_3057,N_49758,N_49916);
or UO_3058 (O_3058,N_49828,N_49854);
or UO_3059 (O_3059,N_49888,N_49861);
nand UO_3060 (O_3060,N_49892,N_49988);
or UO_3061 (O_3061,N_49962,N_49976);
nand UO_3062 (O_3062,N_49908,N_49965);
nor UO_3063 (O_3063,N_49878,N_49989);
nor UO_3064 (O_3064,N_49850,N_49812);
and UO_3065 (O_3065,N_49990,N_49781);
and UO_3066 (O_3066,N_49990,N_49833);
nor UO_3067 (O_3067,N_49860,N_49822);
nor UO_3068 (O_3068,N_49956,N_49982);
nand UO_3069 (O_3069,N_49898,N_49770);
nor UO_3070 (O_3070,N_49786,N_49799);
nand UO_3071 (O_3071,N_49875,N_49872);
or UO_3072 (O_3072,N_49830,N_49817);
and UO_3073 (O_3073,N_49913,N_49773);
or UO_3074 (O_3074,N_49761,N_49859);
or UO_3075 (O_3075,N_49869,N_49959);
and UO_3076 (O_3076,N_49879,N_49869);
or UO_3077 (O_3077,N_49912,N_49955);
nor UO_3078 (O_3078,N_49821,N_49890);
nor UO_3079 (O_3079,N_49779,N_49791);
or UO_3080 (O_3080,N_49988,N_49973);
or UO_3081 (O_3081,N_49987,N_49863);
and UO_3082 (O_3082,N_49819,N_49872);
and UO_3083 (O_3083,N_49857,N_49899);
nand UO_3084 (O_3084,N_49869,N_49857);
or UO_3085 (O_3085,N_49840,N_49932);
xnor UO_3086 (O_3086,N_49958,N_49856);
or UO_3087 (O_3087,N_49977,N_49883);
nor UO_3088 (O_3088,N_49804,N_49797);
nand UO_3089 (O_3089,N_49922,N_49877);
nand UO_3090 (O_3090,N_49850,N_49946);
nor UO_3091 (O_3091,N_49792,N_49898);
nor UO_3092 (O_3092,N_49858,N_49964);
and UO_3093 (O_3093,N_49932,N_49819);
and UO_3094 (O_3094,N_49843,N_49967);
xor UO_3095 (O_3095,N_49793,N_49942);
nand UO_3096 (O_3096,N_49900,N_49876);
nor UO_3097 (O_3097,N_49959,N_49865);
nor UO_3098 (O_3098,N_49796,N_49854);
or UO_3099 (O_3099,N_49953,N_49770);
and UO_3100 (O_3100,N_49910,N_49788);
and UO_3101 (O_3101,N_49944,N_49979);
nor UO_3102 (O_3102,N_49817,N_49907);
and UO_3103 (O_3103,N_49959,N_49754);
and UO_3104 (O_3104,N_49986,N_49967);
nand UO_3105 (O_3105,N_49861,N_49842);
nand UO_3106 (O_3106,N_49991,N_49939);
and UO_3107 (O_3107,N_49855,N_49956);
xor UO_3108 (O_3108,N_49966,N_49934);
and UO_3109 (O_3109,N_49959,N_49946);
xnor UO_3110 (O_3110,N_49869,N_49926);
nand UO_3111 (O_3111,N_49870,N_49865);
or UO_3112 (O_3112,N_49961,N_49881);
xnor UO_3113 (O_3113,N_49975,N_49794);
nand UO_3114 (O_3114,N_49906,N_49904);
and UO_3115 (O_3115,N_49971,N_49887);
or UO_3116 (O_3116,N_49914,N_49780);
nand UO_3117 (O_3117,N_49795,N_49904);
nor UO_3118 (O_3118,N_49826,N_49978);
or UO_3119 (O_3119,N_49866,N_49793);
and UO_3120 (O_3120,N_49856,N_49997);
and UO_3121 (O_3121,N_49762,N_49834);
xnor UO_3122 (O_3122,N_49939,N_49887);
nand UO_3123 (O_3123,N_49823,N_49974);
nor UO_3124 (O_3124,N_49811,N_49874);
nand UO_3125 (O_3125,N_49845,N_49827);
nand UO_3126 (O_3126,N_49972,N_49791);
nand UO_3127 (O_3127,N_49751,N_49884);
or UO_3128 (O_3128,N_49981,N_49990);
or UO_3129 (O_3129,N_49956,N_49963);
xnor UO_3130 (O_3130,N_49761,N_49920);
nand UO_3131 (O_3131,N_49817,N_49949);
nand UO_3132 (O_3132,N_49791,N_49761);
nand UO_3133 (O_3133,N_49773,N_49909);
or UO_3134 (O_3134,N_49873,N_49755);
nand UO_3135 (O_3135,N_49872,N_49883);
and UO_3136 (O_3136,N_49831,N_49794);
nor UO_3137 (O_3137,N_49808,N_49869);
and UO_3138 (O_3138,N_49995,N_49943);
nand UO_3139 (O_3139,N_49937,N_49890);
or UO_3140 (O_3140,N_49931,N_49809);
nand UO_3141 (O_3141,N_49871,N_49928);
or UO_3142 (O_3142,N_49870,N_49769);
and UO_3143 (O_3143,N_49793,N_49771);
nor UO_3144 (O_3144,N_49835,N_49925);
nand UO_3145 (O_3145,N_49803,N_49776);
xnor UO_3146 (O_3146,N_49846,N_49876);
xor UO_3147 (O_3147,N_49993,N_49821);
or UO_3148 (O_3148,N_49999,N_49788);
and UO_3149 (O_3149,N_49971,N_49830);
nand UO_3150 (O_3150,N_49950,N_49855);
nor UO_3151 (O_3151,N_49801,N_49884);
and UO_3152 (O_3152,N_49763,N_49776);
nor UO_3153 (O_3153,N_49767,N_49955);
nand UO_3154 (O_3154,N_49760,N_49887);
or UO_3155 (O_3155,N_49847,N_49911);
xor UO_3156 (O_3156,N_49897,N_49768);
nand UO_3157 (O_3157,N_49984,N_49910);
or UO_3158 (O_3158,N_49998,N_49811);
and UO_3159 (O_3159,N_49836,N_49962);
nand UO_3160 (O_3160,N_49845,N_49947);
nor UO_3161 (O_3161,N_49773,N_49910);
xnor UO_3162 (O_3162,N_49937,N_49796);
xor UO_3163 (O_3163,N_49957,N_49903);
xor UO_3164 (O_3164,N_49861,N_49770);
nor UO_3165 (O_3165,N_49769,N_49846);
nor UO_3166 (O_3166,N_49959,N_49798);
and UO_3167 (O_3167,N_49791,N_49969);
nand UO_3168 (O_3168,N_49942,N_49781);
nor UO_3169 (O_3169,N_49926,N_49787);
nor UO_3170 (O_3170,N_49993,N_49780);
nor UO_3171 (O_3171,N_49886,N_49924);
nand UO_3172 (O_3172,N_49961,N_49895);
and UO_3173 (O_3173,N_49971,N_49946);
nor UO_3174 (O_3174,N_49981,N_49899);
or UO_3175 (O_3175,N_49844,N_49983);
nand UO_3176 (O_3176,N_49933,N_49934);
and UO_3177 (O_3177,N_49782,N_49860);
nand UO_3178 (O_3178,N_49938,N_49880);
nor UO_3179 (O_3179,N_49969,N_49799);
nand UO_3180 (O_3180,N_49876,N_49756);
nand UO_3181 (O_3181,N_49831,N_49804);
nor UO_3182 (O_3182,N_49905,N_49875);
and UO_3183 (O_3183,N_49981,N_49897);
xor UO_3184 (O_3184,N_49868,N_49794);
nand UO_3185 (O_3185,N_49798,N_49813);
xor UO_3186 (O_3186,N_49840,N_49906);
xor UO_3187 (O_3187,N_49795,N_49978);
xnor UO_3188 (O_3188,N_49974,N_49937);
or UO_3189 (O_3189,N_49862,N_49883);
or UO_3190 (O_3190,N_49795,N_49864);
xor UO_3191 (O_3191,N_49967,N_49797);
and UO_3192 (O_3192,N_49868,N_49910);
xnor UO_3193 (O_3193,N_49885,N_49981);
nand UO_3194 (O_3194,N_49919,N_49986);
nand UO_3195 (O_3195,N_49947,N_49982);
and UO_3196 (O_3196,N_49963,N_49990);
and UO_3197 (O_3197,N_49871,N_49801);
nand UO_3198 (O_3198,N_49907,N_49811);
and UO_3199 (O_3199,N_49768,N_49996);
and UO_3200 (O_3200,N_49963,N_49860);
nand UO_3201 (O_3201,N_49938,N_49854);
nor UO_3202 (O_3202,N_49962,N_49845);
xor UO_3203 (O_3203,N_49836,N_49855);
or UO_3204 (O_3204,N_49868,N_49887);
nor UO_3205 (O_3205,N_49776,N_49767);
and UO_3206 (O_3206,N_49842,N_49831);
nand UO_3207 (O_3207,N_49926,N_49795);
and UO_3208 (O_3208,N_49961,N_49901);
or UO_3209 (O_3209,N_49797,N_49978);
or UO_3210 (O_3210,N_49879,N_49771);
xnor UO_3211 (O_3211,N_49833,N_49949);
nor UO_3212 (O_3212,N_49857,N_49792);
nor UO_3213 (O_3213,N_49928,N_49850);
nand UO_3214 (O_3214,N_49898,N_49976);
nand UO_3215 (O_3215,N_49797,N_49831);
and UO_3216 (O_3216,N_49958,N_49802);
xor UO_3217 (O_3217,N_49832,N_49859);
nand UO_3218 (O_3218,N_49854,N_49949);
xnor UO_3219 (O_3219,N_49806,N_49971);
nor UO_3220 (O_3220,N_49803,N_49786);
xnor UO_3221 (O_3221,N_49957,N_49767);
or UO_3222 (O_3222,N_49973,N_49839);
and UO_3223 (O_3223,N_49910,N_49825);
or UO_3224 (O_3224,N_49865,N_49895);
nand UO_3225 (O_3225,N_49824,N_49982);
xnor UO_3226 (O_3226,N_49799,N_49757);
nand UO_3227 (O_3227,N_49909,N_49822);
nor UO_3228 (O_3228,N_49922,N_49970);
and UO_3229 (O_3229,N_49827,N_49849);
or UO_3230 (O_3230,N_49986,N_49917);
nand UO_3231 (O_3231,N_49766,N_49866);
or UO_3232 (O_3232,N_49969,N_49997);
xnor UO_3233 (O_3233,N_49965,N_49769);
xor UO_3234 (O_3234,N_49880,N_49805);
or UO_3235 (O_3235,N_49980,N_49869);
nor UO_3236 (O_3236,N_49898,N_49854);
nor UO_3237 (O_3237,N_49859,N_49831);
or UO_3238 (O_3238,N_49801,N_49907);
nand UO_3239 (O_3239,N_49878,N_49844);
or UO_3240 (O_3240,N_49958,N_49777);
nand UO_3241 (O_3241,N_49841,N_49963);
or UO_3242 (O_3242,N_49812,N_49949);
and UO_3243 (O_3243,N_49834,N_49935);
or UO_3244 (O_3244,N_49787,N_49992);
or UO_3245 (O_3245,N_49900,N_49840);
xnor UO_3246 (O_3246,N_49903,N_49884);
xor UO_3247 (O_3247,N_49980,N_49763);
and UO_3248 (O_3248,N_49879,N_49860);
or UO_3249 (O_3249,N_49956,N_49828);
and UO_3250 (O_3250,N_49960,N_49858);
nor UO_3251 (O_3251,N_49753,N_49803);
nor UO_3252 (O_3252,N_49921,N_49905);
nor UO_3253 (O_3253,N_49863,N_49760);
nand UO_3254 (O_3254,N_49867,N_49898);
nand UO_3255 (O_3255,N_49798,N_49861);
nor UO_3256 (O_3256,N_49817,N_49931);
nor UO_3257 (O_3257,N_49855,N_49905);
and UO_3258 (O_3258,N_49988,N_49890);
nand UO_3259 (O_3259,N_49814,N_49875);
and UO_3260 (O_3260,N_49858,N_49819);
nor UO_3261 (O_3261,N_49754,N_49790);
nor UO_3262 (O_3262,N_49835,N_49941);
nand UO_3263 (O_3263,N_49940,N_49944);
xor UO_3264 (O_3264,N_49752,N_49960);
xor UO_3265 (O_3265,N_49942,N_49912);
xnor UO_3266 (O_3266,N_49944,N_49751);
nor UO_3267 (O_3267,N_49882,N_49839);
xor UO_3268 (O_3268,N_49828,N_49762);
xor UO_3269 (O_3269,N_49973,N_49976);
or UO_3270 (O_3270,N_49765,N_49924);
and UO_3271 (O_3271,N_49934,N_49889);
nor UO_3272 (O_3272,N_49801,N_49989);
nor UO_3273 (O_3273,N_49796,N_49867);
or UO_3274 (O_3274,N_49863,N_49945);
nand UO_3275 (O_3275,N_49856,N_49879);
and UO_3276 (O_3276,N_49897,N_49777);
nor UO_3277 (O_3277,N_49923,N_49843);
or UO_3278 (O_3278,N_49760,N_49774);
or UO_3279 (O_3279,N_49946,N_49849);
xor UO_3280 (O_3280,N_49949,N_49880);
and UO_3281 (O_3281,N_49896,N_49880);
or UO_3282 (O_3282,N_49828,N_49923);
xor UO_3283 (O_3283,N_49911,N_49801);
and UO_3284 (O_3284,N_49878,N_49790);
nor UO_3285 (O_3285,N_49821,N_49891);
or UO_3286 (O_3286,N_49988,N_49819);
nor UO_3287 (O_3287,N_49792,N_49790);
nor UO_3288 (O_3288,N_49996,N_49946);
nand UO_3289 (O_3289,N_49846,N_49808);
or UO_3290 (O_3290,N_49882,N_49756);
and UO_3291 (O_3291,N_49932,N_49884);
nand UO_3292 (O_3292,N_49856,N_49830);
nor UO_3293 (O_3293,N_49886,N_49824);
nand UO_3294 (O_3294,N_49837,N_49983);
and UO_3295 (O_3295,N_49957,N_49879);
nor UO_3296 (O_3296,N_49887,N_49756);
nor UO_3297 (O_3297,N_49796,N_49853);
or UO_3298 (O_3298,N_49760,N_49937);
nand UO_3299 (O_3299,N_49888,N_49801);
or UO_3300 (O_3300,N_49961,N_49808);
or UO_3301 (O_3301,N_49768,N_49825);
and UO_3302 (O_3302,N_49847,N_49981);
xnor UO_3303 (O_3303,N_49999,N_49837);
or UO_3304 (O_3304,N_49750,N_49937);
nor UO_3305 (O_3305,N_49817,N_49908);
and UO_3306 (O_3306,N_49873,N_49803);
xor UO_3307 (O_3307,N_49757,N_49806);
or UO_3308 (O_3308,N_49869,N_49830);
xor UO_3309 (O_3309,N_49767,N_49829);
nor UO_3310 (O_3310,N_49783,N_49873);
and UO_3311 (O_3311,N_49791,N_49864);
and UO_3312 (O_3312,N_49825,N_49979);
or UO_3313 (O_3313,N_49987,N_49887);
nand UO_3314 (O_3314,N_49768,N_49894);
or UO_3315 (O_3315,N_49884,N_49957);
xnor UO_3316 (O_3316,N_49883,N_49968);
nand UO_3317 (O_3317,N_49801,N_49956);
xor UO_3318 (O_3318,N_49963,N_49882);
xnor UO_3319 (O_3319,N_49905,N_49807);
or UO_3320 (O_3320,N_49786,N_49902);
nor UO_3321 (O_3321,N_49981,N_49979);
xnor UO_3322 (O_3322,N_49845,N_49976);
or UO_3323 (O_3323,N_49785,N_49947);
xor UO_3324 (O_3324,N_49752,N_49953);
nor UO_3325 (O_3325,N_49800,N_49984);
xor UO_3326 (O_3326,N_49909,N_49902);
and UO_3327 (O_3327,N_49848,N_49915);
xnor UO_3328 (O_3328,N_49983,N_49891);
xor UO_3329 (O_3329,N_49956,N_49927);
and UO_3330 (O_3330,N_49791,N_49899);
and UO_3331 (O_3331,N_49960,N_49972);
and UO_3332 (O_3332,N_49909,N_49943);
or UO_3333 (O_3333,N_49904,N_49900);
or UO_3334 (O_3334,N_49826,N_49916);
or UO_3335 (O_3335,N_49918,N_49909);
or UO_3336 (O_3336,N_49881,N_49929);
nand UO_3337 (O_3337,N_49890,N_49985);
nand UO_3338 (O_3338,N_49884,N_49961);
and UO_3339 (O_3339,N_49873,N_49931);
and UO_3340 (O_3340,N_49911,N_49845);
nor UO_3341 (O_3341,N_49860,N_49967);
xnor UO_3342 (O_3342,N_49849,N_49759);
or UO_3343 (O_3343,N_49878,N_49789);
nand UO_3344 (O_3344,N_49866,N_49889);
or UO_3345 (O_3345,N_49811,N_49813);
nand UO_3346 (O_3346,N_49801,N_49753);
nand UO_3347 (O_3347,N_49778,N_49788);
or UO_3348 (O_3348,N_49832,N_49996);
and UO_3349 (O_3349,N_49871,N_49861);
nand UO_3350 (O_3350,N_49929,N_49790);
nand UO_3351 (O_3351,N_49816,N_49754);
or UO_3352 (O_3352,N_49800,N_49892);
and UO_3353 (O_3353,N_49883,N_49778);
nor UO_3354 (O_3354,N_49977,N_49870);
nand UO_3355 (O_3355,N_49923,N_49981);
nand UO_3356 (O_3356,N_49777,N_49846);
nand UO_3357 (O_3357,N_49933,N_49858);
and UO_3358 (O_3358,N_49766,N_49786);
xnor UO_3359 (O_3359,N_49939,N_49942);
or UO_3360 (O_3360,N_49946,N_49933);
and UO_3361 (O_3361,N_49813,N_49775);
or UO_3362 (O_3362,N_49814,N_49915);
xor UO_3363 (O_3363,N_49886,N_49884);
and UO_3364 (O_3364,N_49893,N_49806);
xor UO_3365 (O_3365,N_49821,N_49998);
xor UO_3366 (O_3366,N_49796,N_49832);
or UO_3367 (O_3367,N_49876,N_49841);
and UO_3368 (O_3368,N_49860,N_49868);
nand UO_3369 (O_3369,N_49790,N_49842);
nand UO_3370 (O_3370,N_49774,N_49836);
xor UO_3371 (O_3371,N_49979,N_49843);
or UO_3372 (O_3372,N_49861,N_49967);
or UO_3373 (O_3373,N_49941,N_49780);
xor UO_3374 (O_3374,N_49853,N_49897);
and UO_3375 (O_3375,N_49905,N_49821);
or UO_3376 (O_3376,N_49948,N_49835);
nand UO_3377 (O_3377,N_49908,N_49988);
xnor UO_3378 (O_3378,N_49955,N_49983);
and UO_3379 (O_3379,N_49985,N_49919);
xor UO_3380 (O_3380,N_49936,N_49955);
nor UO_3381 (O_3381,N_49848,N_49989);
xor UO_3382 (O_3382,N_49819,N_49990);
nand UO_3383 (O_3383,N_49871,N_49929);
nand UO_3384 (O_3384,N_49779,N_49812);
xor UO_3385 (O_3385,N_49891,N_49935);
xor UO_3386 (O_3386,N_49857,N_49835);
xor UO_3387 (O_3387,N_49991,N_49794);
xnor UO_3388 (O_3388,N_49955,N_49950);
nand UO_3389 (O_3389,N_49985,N_49996);
and UO_3390 (O_3390,N_49826,N_49782);
and UO_3391 (O_3391,N_49825,N_49790);
nor UO_3392 (O_3392,N_49952,N_49774);
or UO_3393 (O_3393,N_49978,N_49773);
nor UO_3394 (O_3394,N_49844,N_49928);
nand UO_3395 (O_3395,N_49919,N_49796);
and UO_3396 (O_3396,N_49934,N_49977);
and UO_3397 (O_3397,N_49965,N_49941);
nor UO_3398 (O_3398,N_49836,N_49933);
nor UO_3399 (O_3399,N_49831,N_49944);
xnor UO_3400 (O_3400,N_49844,N_49971);
nand UO_3401 (O_3401,N_49762,N_49794);
nand UO_3402 (O_3402,N_49908,N_49940);
xor UO_3403 (O_3403,N_49993,N_49917);
nand UO_3404 (O_3404,N_49819,N_49947);
nand UO_3405 (O_3405,N_49907,N_49896);
nand UO_3406 (O_3406,N_49940,N_49935);
nand UO_3407 (O_3407,N_49821,N_49766);
nand UO_3408 (O_3408,N_49956,N_49931);
or UO_3409 (O_3409,N_49967,N_49965);
xnor UO_3410 (O_3410,N_49980,N_49912);
and UO_3411 (O_3411,N_49919,N_49792);
or UO_3412 (O_3412,N_49842,N_49758);
or UO_3413 (O_3413,N_49986,N_49785);
xnor UO_3414 (O_3414,N_49889,N_49772);
nand UO_3415 (O_3415,N_49858,N_49810);
or UO_3416 (O_3416,N_49812,N_49981);
or UO_3417 (O_3417,N_49993,N_49865);
nor UO_3418 (O_3418,N_49869,N_49989);
and UO_3419 (O_3419,N_49928,N_49816);
nor UO_3420 (O_3420,N_49808,N_49866);
nor UO_3421 (O_3421,N_49870,N_49855);
nand UO_3422 (O_3422,N_49854,N_49852);
or UO_3423 (O_3423,N_49888,N_49841);
nand UO_3424 (O_3424,N_49888,N_49908);
xor UO_3425 (O_3425,N_49878,N_49921);
nand UO_3426 (O_3426,N_49876,N_49797);
xor UO_3427 (O_3427,N_49751,N_49852);
nand UO_3428 (O_3428,N_49952,N_49957);
or UO_3429 (O_3429,N_49855,N_49769);
and UO_3430 (O_3430,N_49768,N_49914);
nor UO_3431 (O_3431,N_49751,N_49942);
and UO_3432 (O_3432,N_49980,N_49878);
nor UO_3433 (O_3433,N_49887,N_49969);
nor UO_3434 (O_3434,N_49981,N_49889);
nand UO_3435 (O_3435,N_49901,N_49773);
and UO_3436 (O_3436,N_49780,N_49772);
nand UO_3437 (O_3437,N_49789,N_49957);
or UO_3438 (O_3438,N_49803,N_49764);
and UO_3439 (O_3439,N_49753,N_49993);
nand UO_3440 (O_3440,N_49857,N_49898);
nor UO_3441 (O_3441,N_49876,N_49831);
or UO_3442 (O_3442,N_49956,N_49775);
or UO_3443 (O_3443,N_49950,N_49767);
xor UO_3444 (O_3444,N_49972,N_49925);
nand UO_3445 (O_3445,N_49755,N_49983);
nor UO_3446 (O_3446,N_49999,N_49994);
or UO_3447 (O_3447,N_49831,N_49913);
or UO_3448 (O_3448,N_49884,N_49890);
nor UO_3449 (O_3449,N_49828,N_49917);
nand UO_3450 (O_3450,N_49758,N_49861);
nand UO_3451 (O_3451,N_49993,N_49791);
nand UO_3452 (O_3452,N_49853,N_49883);
nor UO_3453 (O_3453,N_49797,N_49864);
or UO_3454 (O_3454,N_49870,N_49943);
nand UO_3455 (O_3455,N_49775,N_49876);
xnor UO_3456 (O_3456,N_49994,N_49894);
nor UO_3457 (O_3457,N_49757,N_49803);
and UO_3458 (O_3458,N_49897,N_49918);
or UO_3459 (O_3459,N_49818,N_49813);
or UO_3460 (O_3460,N_49877,N_49854);
nor UO_3461 (O_3461,N_49880,N_49824);
or UO_3462 (O_3462,N_49957,N_49906);
xnor UO_3463 (O_3463,N_49751,N_49787);
nor UO_3464 (O_3464,N_49929,N_49901);
nor UO_3465 (O_3465,N_49752,N_49764);
xnor UO_3466 (O_3466,N_49766,N_49831);
or UO_3467 (O_3467,N_49769,N_49836);
and UO_3468 (O_3468,N_49873,N_49851);
nand UO_3469 (O_3469,N_49780,N_49803);
xor UO_3470 (O_3470,N_49862,N_49885);
nor UO_3471 (O_3471,N_49774,N_49872);
or UO_3472 (O_3472,N_49980,N_49872);
nand UO_3473 (O_3473,N_49762,N_49847);
nor UO_3474 (O_3474,N_49854,N_49797);
or UO_3475 (O_3475,N_49819,N_49960);
nor UO_3476 (O_3476,N_49803,N_49929);
nand UO_3477 (O_3477,N_49918,N_49859);
nor UO_3478 (O_3478,N_49875,N_49884);
nor UO_3479 (O_3479,N_49842,N_49858);
or UO_3480 (O_3480,N_49757,N_49824);
or UO_3481 (O_3481,N_49923,N_49805);
nor UO_3482 (O_3482,N_49766,N_49860);
or UO_3483 (O_3483,N_49994,N_49911);
xor UO_3484 (O_3484,N_49855,N_49793);
and UO_3485 (O_3485,N_49983,N_49974);
and UO_3486 (O_3486,N_49889,N_49972);
or UO_3487 (O_3487,N_49822,N_49948);
nand UO_3488 (O_3488,N_49822,N_49897);
xnor UO_3489 (O_3489,N_49861,N_49958);
nand UO_3490 (O_3490,N_49975,N_49791);
nor UO_3491 (O_3491,N_49910,N_49900);
nor UO_3492 (O_3492,N_49772,N_49789);
or UO_3493 (O_3493,N_49827,N_49837);
and UO_3494 (O_3494,N_49965,N_49876);
and UO_3495 (O_3495,N_49956,N_49818);
or UO_3496 (O_3496,N_49949,N_49859);
xnor UO_3497 (O_3497,N_49888,N_49966);
nor UO_3498 (O_3498,N_49792,N_49825);
and UO_3499 (O_3499,N_49948,N_49843);
xnor UO_3500 (O_3500,N_49770,N_49954);
nand UO_3501 (O_3501,N_49884,N_49996);
nand UO_3502 (O_3502,N_49975,N_49974);
or UO_3503 (O_3503,N_49889,N_49991);
and UO_3504 (O_3504,N_49813,N_49916);
and UO_3505 (O_3505,N_49916,N_49897);
xnor UO_3506 (O_3506,N_49875,N_49934);
or UO_3507 (O_3507,N_49937,N_49918);
nor UO_3508 (O_3508,N_49814,N_49882);
or UO_3509 (O_3509,N_49885,N_49973);
nor UO_3510 (O_3510,N_49890,N_49879);
and UO_3511 (O_3511,N_49762,N_49903);
or UO_3512 (O_3512,N_49890,N_49801);
and UO_3513 (O_3513,N_49979,N_49804);
xnor UO_3514 (O_3514,N_49924,N_49860);
and UO_3515 (O_3515,N_49769,N_49896);
xor UO_3516 (O_3516,N_49926,N_49882);
or UO_3517 (O_3517,N_49784,N_49927);
and UO_3518 (O_3518,N_49868,N_49849);
nand UO_3519 (O_3519,N_49981,N_49933);
xor UO_3520 (O_3520,N_49998,N_49834);
nor UO_3521 (O_3521,N_49995,N_49872);
xor UO_3522 (O_3522,N_49977,N_49926);
and UO_3523 (O_3523,N_49767,N_49824);
nand UO_3524 (O_3524,N_49956,N_49946);
nor UO_3525 (O_3525,N_49952,N_49893);
nand UO_3526 (O_3526,N_49993,N_49837);
nand UO_3527 (O_3527,N_49994,N_49761);
xor UO_3528 (O_3528,N_49953,N_49769);
and UO_3529 (O_3529,N_49824,N_49976);
or UO_3530 (O_3530,N_49808,N_49887);
or UO_3531 (O_3531,N_49850,N_49857);
and UO_3532 (O_3532,N_49827,N_49813);
and UO_3533 (O_3533,N_49755,N_49784);
or UO_3534 (O_3534,N_49930,N_49775);
xnor UO_3535 (O_3535,N_49968,N_49818);
nor UO_3536 (O_3536,N_49829,N_49792);
nand UO_3537 (O_3537,N_49964,N_49900);
nor UO_3538 (O_3538,N_49943,N_49881);
nor UO_3539 (O_3539,N_49871,N_49791);
and UO_3540 (O_3540,N_49871,N_49940);
xnor UO_3541 (O_3541,N_49788,N_49833);
and UO_3542 (O_3542,N_49772,N_49791);
nor UO_3543 (O_3543,N_49795,N_49884);
xnor UO_3544 (O_3544,N_49752,N_49803);
xnor UO_3545 (O_3545,N_49941,N_49906);
nand UO_3546 (O_3546,N_49865,N_49772);
nand UO_3547 (O_3547,N_49900,N_49898);
nor UO_3548 (O_3548,N_49789,N_49986);
nor UO_3549 (O_3549,N_49903,N_49761);
nand UO_3550 (O_3550,N_49778,N_49762);
xor UO_3551 (O_3551,N_49813,N_49785);
and UO_3552 (O_3552,N_49901,N_49946);
xnor UO_3553 (O_3553,N_49975,N_49833);
xnor UO_3554 (O_3554,N_49799,N_49999);
and UO_3555 (O_3555,N_49969,N_49857);
nand UO_3556 (O_3556,N_49871,N_49958);
nand UO_3557 (O_3557,N_49929,N_49800);
and UO_3558 (O_3558,N_49945,N_49988);
xnor UO_3559 (O_3559,N_49904,N_49988);
or UO_3560 (O_3560,N_49980,N_49934);
or UO_3561 (O_3561,N_49805,N_49974);
nor UO_3562 (O_3562,N_49895,N_49767);
nor UO_3563 (O_3563,N_49863,N_49779);
or UO_3564 (O_3564,N_49801,N_49879);
xnor UO_3565 (O_3565,N_49793,N_49993);
nor UO_3566 (O_3566,N_49943,N_49908);
and UO_3567 (O_3567,N_49808,N_49889);
xor UO_3568 (O_3568,N_49909,N_49995);
and UO_3569 (O_3569,N_49881,N_49828);
xor UO_3570 (O_3570,N_49865,N_49927);
and UO_3571 (O_3571,N_49999,N_49863);
and UO_3572 (O_3572,N_49776,N_49978);
or UO_3573 (O_3573,N_49808,N_49892);
nor UO_3574 (O_3574,N_49860,N_49814);
or UO_3575 (O_3575,N_49921,N_49958);
and UO_3576 (O_3576,N_49774,N_49757);
nor UO_3577 (O_3577,N_49969,N_49752);
xor UO_3578 (O_3578,N_49921,N_49961);
nand UO_3579 (O_3579,N_49780,N_49920);
xor UO_3580 (O_3580,N_49890,N_49823);
and UO_3581 (O_3581,N_49848,N_49883);
and UO_3582 (O_3582,N_49876,N_49978);
or UO_3583 (O_3583,N_49829,N_49904);
nor UO_3584 (O_3584,N_49775,N_49894);
nand UO_3585 (O_3585,N_49962,N_49851);
nand UO_3586 (O_3586,N_49767,N_49758);
nand UO_3587 (O_3587,N_49973,N_49765);
nor UO_3588 (O_3588,N_49831,N_49957);
or UO_3589 (O_3589,N_49854,N_49760);
nor UO_3590 (O_3590,N_49773,N_49982);
and UO_3591 (O_3591,N_49988,N_49755);
nor UO_3592 (O_3592,N_49948,N_49956);
nand UO_3593 (O_3593,N_49838,N_49754);
nand UO_3594 (O_3594,N_49807,N_49813);
and UO_3595 (O_3595,N_49851,N_49783);
nand UO_3596 (O_3596,N_49830,N_49757);
or UO_3597 (O_3597,N_49957,N_49838);
or UO_3598 (O_3598,N_49974,N_49752);
and UO_3599 (O_3599,N_49955,N_49920);
nor UO_3600 (O_3600,N_49843,N_49848);
and UO_3601 (O_3601,N_49956,N_49848);
or UO_3602 (O_3602,N_49844,N_49754);
or UO_3603 (O_3603,N_49957,N_49835);
nor UO_3604 (O_3604,N_49921,N_49955);
nor UO_3605 (O_3605,N_49916,N_49874);
nand UO_3606 (O_3606,N_49783,N_49766);
or UO_3607 (O_3607,N_49984,N_49929);
xor UO_3608 (O_3608,N_49957,N_49967);
nor UO_3609 (O_3609,N_49924,N_49873);
xor UO_3610 (O_3610,N_49875,N_49813);
or UO_3611 (O_3611,N_49830,N_49838);
nand UO_3612 (O_3612,N_49901,N_49933);
nor UO_3613 (O_3613,N_49897,N_49840);
xnor UO_3614 (O_3614,N_49757,N_49923);
or UO_3615 (O_3615,N_49862,N_49782);
nor UO_3616 (O_3616,N_49837,N_49877);
and UO_3617 (O_3617,N_49778,N_49991);
and UO_3618 (O_3618,N_49752,N_49951);
and UO_3619 (O_3619,N_49758,N_49813);
nor UO_3620 (O_3620,N_49970,N_49947);
nand UO_3621 (O_3621,N_49993,N_49858);
and UO_3622 (O_3622,N_49774,N_49937);
and UO_3623 (O_3623,N_49994,N_49970);
or UO_3624 (O_3624,N_49979,N_49808);
nand UO_3625 (O_3625,N_49987,N_49874);
xor UO_3626 (O_3626,N_49905,N_49896);
xnor UO_3627 (O_3627,N_49781,N_49874);
nor UO_3628 (O_3628,N_49764,N_49789);
xor UO_3629 (O_3629,N_49843,N_49938);
and UO_3630 (O_3630,N_49885,N_49825);
nor UO_3631 (O_3631,N_49777,N_49980);
nor UO_3632 (O_3632,N_49976,N_49868);
xnor UO_3633 (O_3633,N_49979,N_49910);
nor UO_3634 (O_3634,N_49955,N_49931);
nor UO_3635 (O_3635,N_49812,N_49912);
nand UO_3636 (O_3636,N_49937,N_49929);
and UO_3637 (O_3637,N_49752,N_49768);
xor UO_3638 (O_3638,N_49987,N_49778);
nor UO_3639 (O_3639,N_49868,N_49935);
nor UO_3640 (O_3640,N_49977,N_49751);
xor UO_3641 (O_3641,N_49763,N_49753);
nor UO_3642 (O_3642,N_49962,N_49837);
nor UO_3643 (O_3643,N_49970,N_49837);
or UO_3644 (O_3644,N_49921,N_49781);
or UO_3645 (O_3645,N_49931,N_49807);
nand UO_3646 (O_3646,N_49753,N_49809);
nand UO_3647 (O_3647,N_49988,N_49996);
nand UO_3648 (O_3648,N_49753,N_49857);
xor UO_3649 (O_3649,N_49758,N_49778);
nor UO_3650 (O_3650,N_49755,N_49783);
and UO_3651 (O_3651,N_49795,N_49812);
nand UO_3652 (O_3652,N_49999,N_49924);
nand UO_3653 (O_3653,N_49913,N_49829);
xnor UO_3654 (O_3654,N_49968,N_49941);
nor UO_3655 (O_3655,N_49920,N_49795);
nor UO_3656 (O_3656,N_49832,N_49917);
and UO_3657 (O_3657,N_49945,N_49861);
nand UO_3658 (O_3658,N_49823,N_49806);
and UO_3659 (O_3659,N_49794,N_49876);
nand UO_3660 (O_3660,N_49931,N_49815);
nor UO_3661 (O_3661,N_49983,N_49886);
nand UO_3662 (O_3662,N_49904,N_49945);
nor UO_3663 (O_3663,N_49793,N_49818);
and UO_3664 (O_3664,N_49927,N_49806);
and UO_3665 (O_3665,N_49900,N_49885);
nor UO_3666 (O_3666,N_49802,N_49999);
nand UO_3667 (O_3667,N_49843,N_49950);
nor UO_3668 (O_3668,N_49879,N_49806);
or UO_3669 (O_3669,N_49813,N_49901);
nor UO_3670 (O_3670,N_49969,N_49816);
nand UO_3671 (O_3671,N_49835,N_49951);
or UO_3672 (O_3672,N_49992,N_49941);
xnor UO_3673 (O_3673,N_49760,N_49986);
xnor UO_3674 (O_3674,N_49797,N_49803);
nor UO_3675 (O_3675,N_49937,N_49889);
or UO_3676 (O_3676,N_49880,N_49757);
nor UO_3677 (O_3677,N_49908,N_49969);
xor UO_3678 (O_3678,N_49940,N_49887);
nor UO_3679 (O_3679,N_49929,N_49993);
nand UO_3680 (O_3680,N_49848,N_49840);
nand UO_3681 (O_3681,N_49874,N_49753);
and UO_3682 (O_3682,N_49948,N_49907);
nand UO_3683 (O_3683,N_49809,N_49860);
nor UO_3684 (O_3684,N_49771,N_49959);
xor UO_3685 (O_3685,N_49779,N_49799);
nor UO_3686 (O_3686,N_49988,N_49966);
nand UO_3687 (O_3687,N_49836,N_49979);
nand UO_3688 (O_3688,N_49776,N_49909);
nor UO_3689 (O_3689,N_49881,N_49757);
nor UO_3690 (O_3690,N_49883,N_49954);
nand UO_3691 (O_3691,N_49921,N_49971);
or UO_3692 (O_3692,N_49830,N_49781);
and UO_3693 (O_3693,N_49987,N_49879);
nand UO_3694 (O_3694,N_49909,N_49999);
xnor UO_3695 (O_3695,N_49851,N_49791);
or UO_3696 (O_3696,N_49976,N_49846);
xor UO_3697 (O_3697,N_49995,N_49974);
nor UO_3698 (O_3698,N_49827,N_49760);
xnor UO_3699 (O_3699,N_49774,N_49846);
and UO_3700 (O_3700,N_49929,N_49947);
and UO_3701 (O_3701,N_49809,N_49933);
xnor UO_3702 (O_3702,N_49776,N_49993);
nor UO_3703 (O_3703,N_49974,N_49798);
xnor UO_3704 (O_3704,N_49851,N_49999);
nor UO_3705 (O_3705,N_49934,N_49763);
or UO_3706 (O_3706,N_49896,N_49975);
nor UO_3707 (O_3707,N_49868,N_49846);
nand UO_3708 (O_3708,N_49773,N_49841);
and UO_3709 (O_3709,N_49771,N_49989);
xnor UO_3710 (O_3710,N_49812,N_49946);
or UO_3711 (O_3711,N_49936,N_49952);
nor UO_3712 (O_3712,N_49811,N_49855);
and UO_3713 (O_3713,N_49769,N_49903);
and UO_3714 (O_3714,N_49858,N_49963);
nand UO_3715 (O_3715,N_49777,N_49775);
xor UO_3716 (O_3716,N_49981,N_49900);
and UO_3717 (O_3717,N_49930,N_49984);
nand UO_3718 (O_3718,N_49913,N_49814);
nand UO_3719 (O_3719,N_49797,N_49853);
nand UO_3720 (O_3720,N_49923,N_49798);
nor UO_3721 (O_3721,N_49782,N_49765);
and UO_3722 (O_3722,N_49891,N_49920);
nor UO_3723 (O_3723,N_49810,N_49884);
nand UO_3724 (O_3724,N_49779,N_49772);
and UO_3725 (O_3725,N_49756,N_49928);
nand UO_3726 (O_3726,N_49842,N_49819);
nor UO_3727 (O_3727,N_49857,N_49941);
nor UO_3728 (O_3728,N_49840,N_49894);
nor UO_3729 (O_3729,N_49899,N_49772);
nand UO_3730 (O_3730,N_49955,N_49992);
xnor UO_3731 (O_3731,N_49968,N_49848);
xor UO_3732 (O_3732,N_49774,N_49981);
xor UO_3733 (O_3733,N_49790,N_49807);
xnor UO_3734 (O_3734,N_49915,N_49933);
nand UO_3735 (O_3735,N_49864,N_49928);
nand UO_3736 (O_3736,N_49836,N_49977);
xnor UO_3737 (O_3737,N_49961,N_49765);
and UO_3738 (O_3738,N_49928,N_49910);
nand UO_3739 (O_3739,N_49920,N_49843);
nand UO_3740 (O_3740,N_49976,N_49858);
nor UO_3741 (O_3741,N_49912,N_49864);
nand UO_3742 (O_3742,N_49971,N_49942);
or UO_3743 (O_3743,N_49792,N_49905);
nor UO_3744 (O_3744,N_49900,N_49990);
xnor UO_3745 (O_3745,N_49953,N_49857);
nand UO_3746 (O_3746,N_49934,N_49874);
xor UO_3747 (O_3747,N_49917,N_49915);
nor UO_3748 (O_3748,N_49808,N_49809);
and UO_3749 (O_3749,N_49854,N_49925);
and UO_3750 (O_3750,N_49758,N_49926);
xor UO_3751 (O_3751,N_49761,N_49780);
or UO_3752 (O_3752,N_49883,N_49924);
xor UO_3753 (O_3753,N_49936,N_49838);
xnor UO_3754 (O_3754,N_49850,N_49861);
or UO_3755 (O_3755,N_49941,N_49778);
or UO_3756 (O_3756,N_49984,N_49912);
nor UO_3757 (O_3757,N_49895,N_49917);
xnor UO_3758 (O_3758,N_49993,N_49946);
and UO_3759 (O_3759,N_49815,N_49766);
xor UO_3760 (O_3760,N_49859,N_49806);
xnor UO_3761 (O_3761,N_49811,N_49938);
or UO_3762 (O_3762,N_49893,N_49906);
or UO_3763 (O_3763,N_49764,N_49922);
nor UO_3764 (O_3764,N_49753,N_49813);
xor UO_3765 (O_3765,N_49776,N_49985);
nor UO_3766 (O_3766,N_49868,N_49864);
or UO_3767 (O_3767,N_49774,N_49916);
nand UO_3768 (O_3768,N_49928,N_49781);
nor UO_3769 (O_3769,N_49927,N_49759);
xor UO_3770 (O_3770,N_49839,N_49768);
nand UO_3771 (O_3771,N_49808,N_49775);
nor UO_3772 (O_3772,N_49755,N_49845);
or UO_3773 (O_3773,N_49794,N_49819);
and UO_3774 (O_3774,N_49804,N_49879);
nor UO_3775 (O_3775,N_49803,N_49862);
xnor UO_3776 (O_3776,N_49919,N_49994);
xnor UO_3777 (O_3777,N_49786,N_49889);
or UO_3778 (O_3778,N_49913,N_49933);
xor UO_3779 (O_3779,N_49773,N_49904);
nand UO_3780 (O_3780,N_49999,N_49826);
nor UO_3781 (O_3781,N_49867,N_49966);
nor UO_3782 (O_3782,N_49993,N_49799);
xnor UO_3783 (O_3783,N_49841,N_49980);
and UO_3784 (O_3784,N_49967,N_49925);
or UO_3785 (O_3785,N_49914,N_49833);
or UO_3786 (O_3786,N_49798,N_49927);
or UO_3787 (O_3787,N_49824,N_49964);
xor UO_3788 (O_3788,N_49872,N_49779);
and UO_3789 (O_3789,N_49751,N_49963);
nor UO_3790 (O_3790,N_49911,N_49989);
xor UO_3791 (O_3791,N_49939,N_49935);
and UO_3792 (O_3792,N_49813,N_49859);
and UO_3793 (O_3793,N_49974,N_49903);
and UO_3794 (O_3794,N_49994,N_49950);
nor UO_3795 (O_3795,N_49889,N_49832);
nor UO_3796 (O_3796,N_49794,N_49779);
and UO_3797 (O_3797,N_49930,N_49989);
nor UO_3798 (O_3798,N_49976,N_49988);
nand UO_3799 (O_3799,N_49760,N_49906);
or UO_3800 (O_3800,N_49823,N_49942);
and UO_3801 (O_3801,N_49832,N_49827);
or UO_3802 (O_3802,N_49915,N_49829);
and UO_3803 (O_3803,N_49949,N_49907);
or UO_3804 (O_3804,N_49839,N_49875);
xor UO_3805 (O_3805,N_49919,N_49787);
and UO_3806 (O_3806,N_49944,N_49840);
xnor UO_3807 (O_3807,N_49818,N_49989);
xor UO_3808 (O_3808,N_49849,N_49898);
and UO_3809 (O_3809,N_49953,N_49792);
and UO_3810 (O_3810,N_49992,N_49997);
nor UO_3811 (O_3811,N_49870,N_49935);
nor UO_3812 (O_3812,N_49866,N_49895);
xnor UO_3813 (O_3813,N_49938,N_49981);
nor UO_3814 (O_3814,N_49975,N_49952);
xor UO_3815 (O_3815,N_49993,N_49902);
and UO_3816 (O_3816,N_49978,N_49842);
and UO_3817 (O_3817,N_49950,N_49839);
and UO_3818 (O_3818,N_49875,N_49977);
and UO_3819 (O_3819,N_49889,N_49978);
nand UO_3820 (O_3820,N_49869,N_49809);
and UO_3821 (O_3821,N_49777,N_49990);
xnor UO_3822 (O_3822,N_49824,N_49861);
and UO_3823 (O_3823,N_49792,N_49799);
nand UO_3824 (O_3824,N_49792,N_49789);
and UO_3825 (O_3825,N_49941,N_49825);
nor UO_3826 (O_3826,N_49853,N_49909);
xor UO_3827 (O_3827,N_49839,N_49968);
nand UO_3828 (O_3828,N_49775,N_49971);
or UO_3829 (O_3829,N_49986,N_49931);
or UO_3830 (O_3830,N_49810,N_49966);
nor UO_3831 (O_3831,N_49999,N_49832);
xor UO_3832 (O_3832,N_49775,N_49952);
nor UO_3833 (O_3833,N_49896,N_49922);
xor UO_3834 (O_3834,N_49846,N_49751);
nor UO_3835 (O_3835,N_49984,N_49873);
xor UO_3836 (O_3836,N_49786,N_49878);
and UO_3837 (O_3837,N_49896,N_49877);
nand UO_3838 (O_3838,N_49829,N_49998);
and UO_3839 (O_3839,N_49806,N_49912);
nor UO_3840 (O_3840,N_49888,N_49919);
and UO_3841 (O_3841,N_49997,N_49878);
and UO_3842 (O_3842,N_49882,N_49790);
nor UO_3843 (O_3843,N_49899,N_49974);
or UO_3844 (O_3844,N_49993,N_49806);
nor UO_3845 (O_3845,N_49985,N_49823);
or UO_3846 (O_3846,N_49979,N_49862);
or UO_3847 (O_3847,N_49843,N_49815);
xor UO_3848 (O_3848,N_49903,N_49917);
nor UO_3849 (O_3849,N_49805,N_49810);
and UO_3850 (O_3850,N_49847,N_49912);
nand UO_3851 (O_3851,N_49974,N_49854);
nand UO_3852 (O_3852,N_49835,N_49840);
xnor UO_3853 (O_3853,N_49818,N_49863);
nand UO_3854 (O_3854,N_49959,N_49969);
and UO_3855 (O_3855,N_49900,N_49976);
nor UO_3856 (O_3856,N_49990,N_49920);
and UO_3857 (O_3857,N_49808,N_49785);
or UO_3858 (O_3858,N_49933,N_49804);
xnor UO_3859 (O_3859,N_49778,N_49825);
nor UO_3860 (O_3860,N_49907,N_49958);
nand UO_3861 (O_3861,N_49946,N_49806);
and UO_3862 (O_3862,N_49818,N_49868);
nand UO_3863 (O_3863,N_49854,N_49928);
nor UO_3864 (O_3864,N_49906,N_49810);
nor UO_3865 (O_3865,N_49927,N_49931);
nand UO_3866 (O_3866,N_49787,N_49835);
or UO_3867 (O_3867,N_49995,N_49849);
xor UO_3868 (O_3868,N_49841,N_49930);
nor UO_3869 (O_3869,N_49866,N_49984);
or UO_3870 (O_3870,N_49795,N_49960);
or UO_3871 (O_3871,N_49857,N_49805);
nand UO_3872 (O_3872,N_49981,N_49777);
nand UO_3873 (O_3873,N_49764,N_49906);
or UO_3874 (O_3874,N_49979,N_49807);
and UO_3875 (O_3875,N_49898,N_49938);
or UO_3876 (O_3876,N_49952,N_49924);
and UO_3877 (O_3877,N_49885,N_49890);
or UO_3878 (O_3878,N_49910,N_49862);
and UO_3879 (O_3879,N_49850,N_49932);
and UO_3880 (O_3880,N_49802,N_49978);
and UO_3881 (O_3881,N_49766,N_49936);
nand UO_3882 (O_3882,N_49919,N_49845);
nand UO_3883 (O_3883,N_49985,N_49875);
nand UO_3884 (O_3884,N_49973,N_49890);
or UO_3885 (O_3885,N_49939,N_49827);
nand UO_3886 (O_3886,N_49793,N_49851);
nor UO_3887 (O_3887,N_49932,N_49944);
and UO_3888 (O_3888,N_49807,N_49923);
or UO_3889 (O_3889,N_49990,N_49927);
or UO_3890 (O_3890,N_49840,N_49907);
nand UO_3891 (O_3891,N_49907,N_49854);
and UO_3892 (O_3892,N_49855,N_49889);
and UO_3893 (O_3893,N_49940,N_49812);
nor UO_3894 (O_3894,N_49931,N_49869);
nand UO_3895 (O_3895,N_49920,N_49998);
nand UO_3896 (O_3896,N_49908,N_49912);
nor UO_3897 (O_3897,N_49809,N_49828);
nor UO_3898 (O_3898,N_49994,N_49836);
and UO_3899 (O_3899,N_49771,N_49875);
or UO_3900 (O_3900,N_49949,N_49911);
nor UO_3901 (O_3901,N_49753,N_49837);
nand UO_3902 (O_3902,N_49905,N_49753);
nor UO_3903 (O_3903,N_49919,N_49929);
nand UO_3904 (O_3904,N_49762,N_49984);
xnor UO_3905 (O_3905,N_49848,N_49927);
xor UO_3906 (O_3906,N_49831,N_49960);
xnor UO_3907 (O_3907,N_49957,N_49864);
nor UO_3908 (O_3908,N_49825,N_49856);
xnor UO_3909 (O_3909,N_49817,N_49933);
xnor UO_3910 (O_3910,N_49774,N_49877);
nand UO_3911 (O_3911,N_49784,N_49858);
and UO_3912 (O_3912,N_49770,N_49774);
nor UO_3913 (O_3913,N_49887,N_49997);
or UO_3914 (O_3914,N_49796,N_49912);
or UO_3915 (O_3915,N_49897,N_49847);
nor UO_3916 (O_3916,N_49861,N_49909);
or UO_3917 (O_3917,N_49912,N_49782);
nor UO_3918 (O_3918,N_49754,N_49842);
xnor UO_3919 (O_3919,N_49979,N_49754);
or UO_3920 (O_3920,N_49793,N_49902);
or UO_3921 (O_3921,N_49892,N_49890);
nand UO_3922 (O_3922,N_49940,N_49856);
nand UO_3923 (O_3923,N_49894,N_49887);
or UO_3924 (O_3924,N_49955,N_49926);
nand UO_3925 (O_3925,N_49981,N_49793);
xnor UO_3926 (O_3926,N_49808,N_49936);
or UO_3927 (O_3927,N_49779,N_49759);
and UO_3928 (O_3928,N_49907,N_49877);
nor UO_3929 (O_3929,N_49802,N_49858);
nand UO_3930 (O_3930,N_49861,N_49868);
xnor UO_3931 (O_3931,N_49782,N_49815);
xor UO_3932 (O_3932,N_49862,N_49892);
or UO_3933 (O_3933,N_49918,N_49866);
nor UO_3934 (O_3934,N_49783,N_49997);
xnor UO_3935 (O_3935,N_49992,N_49791);
nor UO_3936 (O_3936,N_49831,N_49799);
nor UO_3937 (O_3937,N_49819,N_49897);
or UO_3938 (O_3938,N_49989,N_49883);
nand UO_3939 (O_3939,N_49854,N_49903);
nand UO_3940 (O_3940,N_49859,N_49926);
xor UO_3941 (O_3941,N_49756,N_49820);
and UO_3942 (O_3942,N_49927,N_49958);
or UO_3943 (O_3943,N_49933,N_49968);
or UO_3944 (O_3944,N_49909,N_49897);
xor UO_3945 (O_3945,N_49856,N_49951);
and UO_3946 (O_3946,N_49896,N_49780);
and UO_3947 (O_3947,N_49813,N_49789);
xnor UO_3948 (O_3948,N_49813,N_49866);
nor UO_3949 (O_3949,N_49952,N_49830);
xnor UO_3950 (O_3950,N_49770,N_49757);
nor UO_3951 (O_3951,N_49902,N_49931);
or UO_3952 (O_3952,N_49897,N_49771);
nand UO_3953 (O_3953,N_49974,N_49791);
or UO_3954 (O_3954,N_49971,N_49787);
nor UO_3955 (O_3955,N_49861,N_49972);
nand UO_3956 (O_3956,N_49914,N_49937);
xor UO_3957 (O_3957,N_49817,N_49828);
and UO_3958 (O_3958,N_49842,N_49827);
or UO_3959 (O_3959,N_49752,N_49983);
nor UO_3960 (O_3960,N_49842,N_49982);
nand UO_3961 (O_3961,N_49853,N_49886);
and UO_3962 (O_3962,N_49825,N_49922);
and UO_3963 (O_3963,N_49846,N_49884);
xnor UO_3964 (O_3964,N_49780,N_49755);
nand UO_3965 (O_3965,N_49863,N_49838);
xnor UO_3966 (O_3966,N_49856,N_49933);
xnor UO_3967 (O_3967,N_49949,N_49816);
or UO_3968 (O_3968,N_49932,N_49766);
and UO_3969 (O_3969,N_49960,N_49965);
and UO_3970 (O_3970,N_49985,N_49772);
or UO_3971 (O_3971,N_49933,N_49950);
and UO_3972 (O_3972,N_49947,N_49750);
nand UO_3973 (O_3973,N_49916,N_49888);
xnor UO_3974 (O_3974,N_49867,N_49866);
nor UO_3975 (O_3975,N_49888,N_49834);
nand UO_3976 (O_3976,N_49757,N_49976);
nand UO_3977 (O_3977,N_49799,N_49813);
and UO_3978 (O_3978,N_49914,N_49915);
nand UO_3979 (O_3979,N_49796,N_49858);
nor UO_3980 (O_3980,N_49886,N_49818);
or UO_3981 (O_3981,N_49966,N_49886);
or UO_3982 (O_3982,N_49777,N_49856);
or UO_3983 (O_3983,N_49976,N_49765);
or UO_3984 (O_3984,N_49898,N_49826);
and UO_3985 (O_3985,N_49998,N_49816);
nor UO_3986 (O_3986,N_49956,N_49972);
xnor UO_3987 (O_3987,N_49791,N_49873);
nor UO_3988 (O_3988,N_49770,N_49828);
xor UO_3989 (O_3989,N_49982,N_49759);
xnor UO_3990 (O_3990,N_49821,N_49892);
and UO_3991 (O_3991,N_49869,N_49994);
or UO_3992 (O_3992,N_49918,N_49905);
xor UO_3993 (O_3993,N_49970,N_49927);
or UO_3994 (O_3994,N_49906,N_49857);
nand UO_3995 (O_3995,N_49788,N_49821);
nand UO_3996 (O_3996,N_49828,N_49937);
nor UO_3997 (O_3997,N_49903,N_49959);
xnor UO_3998 (O_3998,N_49925,N_49993);
or UO_3999 (O_3999,N_49987,N_49862);
nor UO_4000 (O_4000,N_49944,N_49870);
and UO_4001 (O_4001,N_49956,N_49781);
or UO_4002 (O_4002,N_49776,N_49755);
nand UO_4003 (O_4003,N_49864,N_49972);
or UO_4004 (O_4004,N_49814,N_49965);
xnor UO_4005 (O_4005,N_49983,N_49998);
xnor UO_4006 (O_4006,N_49912,N_49815);
or UO_4007 (O_4007,N_49810,N_49791);
and UO_4008 (O_4008,N_49881,N_49965);
and UO_4009 (O_4009,N_49836,N_49926);
xor UO_4010 (O_4010,N_49799,N_49873);
xor UO_4011 (O_4011,N_49846,N_49819);
nor UO_4012 (O_4012,N_49817,N_49759);
or UO_4013 (O_4013,N_49951,N_49834);
nor UO_4014 (O_4014,N_49966,N_49848);
or UO_4015 (O_4015,N_49923,N_49916);
xnor UO_4016 (O_4016,N_49785,N_49907);
or UO_4017 (O_4017,N_49805,N_49853);
xor UO_4018 (O_4018,N_49955,N_49760);
xnor UO_4019 (O_4019,N_49799,N_49869);
or UO_4020 (O_4020,N_49801,N_49944);
or UO_4021 (O_4021,N_49833,N_49899);
nand UO_4022 (O_4022,N_49761,N_49890);
and UO_4023 (O_4023,N_49855,N_49984);
nor UO_4024 (O_4024,N_49891,N_49832);
and UO_4025 (O_4025,N_49750,N_49848);
nor UO_4026 (O_4026,N_49869,N_49780);
xor UO_4027 (O_4027,N_49862,N_49874);
or UO_4028 (O_4028,N_49795,N_49875);
or UO_4029 (O_4029,N_49756,N_49875);
nand UO_4030 (O_4030,N_49977,N_49890);
nand UO_4031 (O_4031,N_49801,N_49860);
xor UO_4032 (O_4032,N_49767,N_49965);
nor UO_4033 (O_4033,N_49947,N_49769);
or UO_4034 (O_4034,N_49835,N_49908);
nand UO_4035 (O_4035,N_49823,N_49926);
and UO_4036 (O_4036,N_49789,N_49885);
xor UO_4037 (O_4037,N_49769,N_49800);
or UO_4038 (O_4038,N_49824,N_49984);
and UO_4039 (O_4039,N_49904,N_49920);
nand UO_4040 (O_4040,N_49975,N_49840);
and UO_4041 (O_4041,N_49954,N_49887);
or UO_4042 (O_4042,N_49994,N_49770);
xnor UO_4043 (O_4043,N_49802,N_49839);
or UO_4044 (O_4044,N_49939,N_49962);
xnor UO_4045 (O_4045,N_49969,N_49786);
and UO_4046 (O_4046,N_49847,N_49978);
nand UO_4047 (O_4047,N_49978,N_49989);
or UO_4048 (O_4048,N_49838,N_49794);
and UO_4049 (O_4049,N_49989,N_49856);
nor UO_4050 (O_4050,N_49990,N_49767);
or UO_4051 (O_4051,N_49840,N_49866);
or UO_4052 (O_4052,N_49911,N_49751);
nor UO_4053 (O_4053,N_49802,N_49759);
xnor UO_4054 (O_4054,N_49817,N_49947);
and UO_4055 (O_4055,N_49908,N_49858);
nand UO_4056 (O_4056,N_49872,N_49892);
and UO_4057 (O_4057,N_49942,N_49964);
nor UO_4058 (O_4058,N_49777,N_49841);
and UO_4059 (O_4059,N_49823,N_49982);
nand UO_4060 (O_4060,N_49911,N_49861);
or UO_4061 (O_4061,N_49982,N_49881);
or UO_4062 (O_4062,N_49997,N_49897);
nand UO_4063 (O_4063,N_49898,N_49961);
nor UO_4064 (O_4064,N_49821,N_49866);
nand UO_4065 (O_4065,N_49978,N_49848);
nor UO_4066 (O_4066,N_49935,N_49788);
xnor UO_4067 (O_4067,N_49967,N_49921);
nor UO_4068 (O_4068,N_49859,N_49817);
xor UO_4069 (O_4069,N_49920,N_49975);
nand UO_4070 (O_4070,N_49900,N_49985);
nand UO_4071 (O_4071,N_49857,N_49963);
xor UO_4072 (O_4072,N_49806,N_49989);
xnor UO_4073 (O_4073,N_49909,N_49980);
nand UO_4074 (O_4074,N_49786,N_49811);
nor UO_4075 (O_4075,N_49832,N_49881);
and UO_4076 (O_4076,N_49937,N_49912);
and UO_4077 (O_4077,N_49824,N_49908);
or UO_4078 (O_4078,N_49782,N_49802);
xnor UO_4079 (O_4079,N_49830,N_49819);
or UO_4080 (O_4080,N_49780,N_49961);
nand UO_4081 (O_4081,N_49959,N_49844);
and UO_4082 (O_4082,N_49924,N_49854);
nand UO_4083 (O_4083,N_49927,N_49775);
xor UO_4084 (O_4084,N_49895,N_49846);
or UO_4085 (O_4085,N_49791,N_49798);
and UO_4086 (O_4086,N_49798,N_49784);
nand UO_4087 (O_4087,N_49912,N_49830);
and UO_4088 (O_4088,N_49861,N_49817);
and UO_4089 (O_4089,N_49832,N_49920);
or UO_4090 (O_4090,N_49946,N_49872);
nand UO_4091 (O_4091,N_49756,N_49859);
nor UO_4092 (O_4092,N_49820,N_49887);
nand UO_4093 (O_4093,N_49879,N_49805);
and UO_4094 (O_4094,N_49992,N_49994);
xnor UO_4095 (O_4095,N_49888,N_49893);
nor UO_4096 (O_4096,N_49975,N_49784);
and UO_4097 (O_4097,N_49864,N_49869);
nor UO_4098 (O_4098,N_49866,N_49931);
xnor UO_4099 (O_4099,N_49941,N_49862);
and UO_4100 (O_4100,N_49757,N_49898);
nor UO_4101 (O_4101,N_49788,N_49915);
nor UO_4102 (O_4102,N_49840,N_49836);
or UO_4103 (O_4103,N_49783,N_49999);
nand UO_4104 (O_4104,N_49879,N_49796);
xnor UO_4105 (O_4105,N_49892,N_49901);
and UO_4106 (O_4106,N_49934,N_49944);
xnor UO_4107 (O_4107,N_49970,N_49794);
or UO_4108 (O_4108,N_49959,N_49795);
and UO_4109 (O_4109,N_49789,N_49973);
nand UO_4110 (O_4110,N_49834,N_49938);
and UO_4111 (O_4111,N_49824,N_49822);
or UO_4112 (O_4112,N_49998,N_49793);
or UO_4113 (O_4113,N_49755,N_49888);
nor UO_4114 (O_4114,N_49835,N_49950);
or UO_4115 (O_4115,N_49854,N_49880);
nor UO_4116 (O_4116,N_49809,N_49966);
and UO_4117 (O_4117,N_49798,N_49850);
and UO_4118 (O_4118,N_49923,N_49812);
and UO_4119 (O_4119,N_49938,N_49807);
nand UO_4120 (O_4120,N_49924,N_49772);
nand UO_4121 (O_4121,N_49780,N_49861);
or UO_4122 (O_4122,N_49827,N_49975);
nor UO_4123 (O_4123,N_49819,N_49910);
xor UO_4124 (O_4124,N_49998,N_49980);
or UO_4125 (O_4125,N_49809,N_49960);
or UO_4126 (O_4126,N_49836,N_49831);
nand UO_4127 (O_4127,N_49860,N_49862);
nand UO_4128 (O_4128,N_49929,N_49940);
nor UO_4129 (O_4129,N_49948,N_49781);
or UO_4130 (O_4130,N_49778,N_49889);
or UO_4131 (O_4131,N_49956,N_49857);
xnor UO_4132 (O_4132,N_49855,N_49946);
nand UO_4133 (O_4133,N_49931,N_49903);
xor UO_4134 (O_4134,N_49809,N_49873);
xnor UO_4135 (O_4135,N_49859,N_49794);
nor UO_4136 (O_4136,N_49752,N_49842);
xnor UO_4137 (O_4137,N_49857,N_49950);
nand UO_4138 (O_4138,N_49772,N_49948);
or UO_4139 (O_4139,N_49829,N_49764);
or UO_4140 (O_4140,N_49796,N_49830);
nor UO_4141 (O_4141,N_49965,N_49906);
nand UO_4142 (O_4142,N_49838,N_49949);
or UO_4143 (O_4143,N_49941,N_49811);
nand UO_4144 (O_4144,N_49811,N_49877);
nand UO_4145 (O_4145,N_49974,N_49869);
or UO_4146 (O_4146,N_49943,N_49860);
nor UO_4147 (O_4147,N_49929,N_49922);
nor UO_4148 (O_4148,N_49882,N_49999);
or UO_4149 (O_4149,N_49780,N_49776);
or UO_4150 (O_4150,N_49993,N_49854);
or UO_4151 (O_4151,N_49916,N_49893);
or UO_4152 (O_4152,N_49956,N_49939);
and UO_4153 (O_4153,N_49985,N_49980);
nor UO_4154 (O_4154,N_49900,N_49788);
nor UO_4155 (O_4155,N_49965,N_49754);
nand UO_4156 (O_4156,N_49796,N_49772);
nor UO_4157 (O_4157,N_49967,N_49761);
nand UO_4158 (O_4158,N_49921,N_49828);
nand UO_4159 (O_4159,N_49989,N_49994);
and UO_4160 (O_4160,N_49996,N_49840);
nand UO_4161 (O_4161,N_49930,N_49777);
and UO_4162 (O_4162,N_49808,N_49964);
nand UO_4163 (O_4163,N_49958,N_49965);
nor UO_4164 (O_4164,N_49938,N_49833);
and UO_4165 (O_4165,N_49932,N_49908);
xor UO_4166 (O_4166,N_49902,N_49913);
or UO_4167 (O_4167,N_49837,N_49819);
and UO_4168 (O_4168,N_49896,N_49874);
nor UO_4169 (O_4169,N_49894,N_49799);
or UO_4170 (O_4170,N_49841,N_49973);
nor UO_4171 (O_4171,N_49871,N_49845);
and UO_4172 (O_4172,N_49906,N_49770);
and UO_4173 (O_4173,N_49839,N_49835);
xnor UO_4174 (O_4174,N_49887,N_49902);
nand UO_4175 (O_4175,N_49998,N_49820);
nand UO_4176 (O_4176,N_49850,N_49775);
nand UO_4177 (O_4177,N_49920,N_49760);
or UO_4178 (O_4178,N_49870,N_49751);
and UO_4179 (O_4179,N_49854,N_49985);
and UO_4180 (O_4180,N_49975,N_49785);
nand UO_4181 (O_4181,N_49836,N_49865);
nand UO_4182 (O_4182,N_49881,N_49818);
xnor UO_4183 (O_4183,N_49768,N_49862);
or UO_4184 (O_4184,N_49932,N_49761);
xor UO_4185 (O_4185,N_49848,N_49979);
xnor UO_4186 (O_4186,N_49814,N_49811);
nand UO_4187 (O_4187,N_49757,N_49870);
xor UO_4188 (O_4188,N_49799,N_49905);
xor UO_4189 (O_4189,N_49946,N_49935);
and UO_4190 (O_4190,N_49828,N_49879);
nand UO_4191 (O_4191,N_49927,N_49801);
nor UO_4192 (O_4192,N_49980,N_49823);
nand UO_4193 (O_4193,N_49821,N_49995);
nand UO_4194 (O_4194,N_49930,N_49944);
xor UO_4195 (O_4195,N_49805,N_49914);
nand UO_4196 (O_4196,N_49814,N_49970);
and UO_4197 (O_4197,N_49783,N_49922);
xnor UO_4198 (O_4198,N_49940,N_49853);
nor UO_4199 (O_4199,N_49796,N_49810);
nor UO_4200 (O_4200,N_49881,N_49888);
and UO_4201 (O_4201,N_49876,N_49799);
xor UO_4202 (O_4202,N_49921,N_49994);
or UO_4203 (O_4203,N_49754,N_49776);
and UO_4204 (O_4204,N_49974,N_49868);
xor UO_4205 (O_4205,N_49994,N_49926);
xor UO_4206 (O_4206,N_49835,N_49773);
nand UO_4207 (O_4207,N_49850,N_49895);
and UO_4208 (O_4208,N_49902,N_49921);
or UO_4209 (O_4209,N_49846,N_49806);
nand UO_4210 (O_4210,N_49756,N_49858);
and UO_4211 (O_4211,N_49793,N_49882);
xnor UO_4212 (O_4212,N_49841,N_49819);
or UO_4213 (O_4213,N_49897,N_49929);
or UO_4214 (O_4214,N_49849,N_49877);
nor UO_4215 (O_4215,N_49922,N_49779);
nand UO_4216 (O_4216,N_49963,N_49790);
nor UO_4217 (O_4217,N_49856,N_49955);
and UO_4218 (O_4218,N_49817,N_49816);
nand UO_4219 (O_4219,N_49921,N_49830);
nor UO_4220 (O_4220,N_49816,N_49826);
xnor UO_4221 (O_4221,N_49834,N_49772);
nand UO_4222 (O_4222,N_49829,N_49919);
xor UO_4223 (O_4223,N_49888,N_49950);
xnor UO_4224 (O_4224,N_49876,N_49791);
and UO_4225 (O_4225,N_49809,N_49806);
nor UO_4226 (O_4226,N_49829,N_49768);
nand UO_4227 (O_4227,N_49967,N_49907);
xor UO_4228 (O_4228,N_49779,N_49985);
and UO_4229 (O_4229,N_49750,N_49787);
nor UO_4230 (O_4230,N_49810,N_49914);
xnor UO_4231 (O_4231,N_49940,N_49972);
and UO_4232 (O_4232,N_49994,N_49965);
nand UO_4233 (O_4233,N_49944,N_49916);
and UO_4234 (O_4234,N_49752,N_49797);
or UO_4235 (O_4235,N_49878,N_49807);
and UO_4236 (O_4236,N_49936,N_49871);
nand UO_4237 (O_4237,N_49874,N_49828);
or UO_4238 (O_4238,N_49870,N_49928);
or UO_4239 (O_4239,N_49765,N_49794);
and UO_4240 (O_4240,N_49833,N_49771);
nor UO_4241 (O_4241,N_49966,N_49997);
xnor UO_4242 (O_4242,N_49858,N_49952);
nand UO_4243 (O_4243,N_49902,N_49844);
xnor UO_4244 (O_4244,N_49931,N_49844);
nor UO_4245 (O_4245,N_49896,N_49818);
xnor UO_4246 (O_4246,N_49798,N_49970);
xor UO_4247 (O_4247,N_49814,N_49981);
nor UO_4248 (O_4248,N_49821,N_49974);
xor UO_4249 (O_4249,N_49871,N_49795);
and UO_4250 (O_4250,N_49857,N_49840);
nand UO_4251 (O_4251,N_49761,N_49894);
nor UO_4252 (O_4252,N_49966,N_49975);
xor UO_4253 (O_4253,N_49783,N_49877);
nand UO_4254 (O_4254,N_49875,N_49797);
nor UO_4255 (O_4255,N_49943,N_49802);
xor UO_4256 (O_4256,N_49871,N_49855);
nand UO_4257 (O_4257,N_49913,N_49783);
xor UO_4258 (O_4258,N_49835,N_49755);
nor UO_4259 (O_4259,N_49772,N_49752);
nor UO_4260 (O_4260,N_49978,N_49945);
nand UO_4261 (O_4261,N_49890,N_49809);
and UO_4262 (O_4262,N_49959,N_49841);
nand UO_4263 (O_4263,N_49780,N_49767);
and UO_4264 (O_4264,N_49993,N_49889);
or UO_4265 (O_4265,N_49760,N_49782);
and UO_4266 (O_4266,N_49968,N_49911);
nand UO_4267 (O_4267,N_49754,N_49861);
xnor UO_4268 (O_4268,N_49841,N_49924);
xnor UO_4269 (O_4269,N_49836,N_49758);
xnor UO_4270 (O_4270,N_49906,N_49819);
nor UO_4271 (O_4271,N_49966,N_49974);
nand UO_4272 (O_4272,N_49755,N_49790);
xnor UO_4273 (O_4273,N_49958,N_49903);
nor UO_4274 (O_4274,N_49976,N_49840);
or UO_4275 (O_4275,N_49927,N_49973);
nor UO_4276 (O_4276,N_49801,N_49974);
and UO_4277 (O_4277,N_49764,N_49938);
or UO_4278 (O_4278,N_49888,N_49905);
xor UO_4279 (O_4279,N_49872,N_49791);
xnor UO_4280 (O_4280,N_49864,N_49826);
nand UO_4281 (O_4281,N_49820,N_49797);
nor UO_4282 (O_4282,N_49934,N_49900);
or UO_4283 (O_4283,N_49945,N_49897);
or UO_4284 (O_4284,N_49920,N_49805);
nor UO_4285 (O_4285,N_49917,N_49850);
nand UO_4286 (O_4286,N_49828,N_49850);
nor UO_4287 (O_4287,N_49863,N_49858);
or UO_4288 (O_4288,N_49828,N_49805);
and UO_4289 (O_4289,N_49798,N_49975);
nor UO_4290 (O_4290,N_49880,N_49780);
nand UO_4291 (O_4291,N_49902,N_49861);
nand UO_4292 (O_4292,N_49804,N_49820);
or UO_4293 (O_4293,N_49968,N_49990);
nor UO_4294 (O_4294,N_49919,N_49993);
nor UO_4295 (O_4295,N_49814,N_49806);
and UO_4296 (O_4296,N_49880,N_49782);
xor UO_4297 (O_4297,N_49947,N_49777);
nand UO_4298 (O_4298,N_49974,N_49978);
xor UO_4299 (O_4299,N_49846,N_49854);
and UO_4300 (O_4300,N_49930,N_49980);
nand UO_4301 (O_4301,N_49802,N_49937);
xor UO_4302 (O_4302,N_49863,N_49957);
nor UO_4303 (O_4303,N_49834,N_49949);
nand UO_4304 (O_4304,N_49852,N_49938);
nor UO_4305 (O_4305,N_49881,N_49872);
nand UO_4306 (O_4306,N_49801,N_49894);
nand UO_4307 (O_4307,N_49865,N_49926);
nand UO_4308 (O_4308,N_49930,N_49975);
nand UO_4309 (O_4309,N_49808,N_49978);
or UO_4310 (O_4310,N_49753,N_49923);
and UO_4311 (O_4311,N_49986,N_49751);
and UO_4312 (O_4312,N_49995,N_49852);
or UO_4313 (O_4313,N_49868,N_49803);
or UO_4314 (O_4314,N_49968,N_49988);
nand UO_4315 (O_4315,N_49775,N_49828);
or UO_4316 (O_4316,N_49842,N_49974);
xnor UO_4317 (O_4317,N_49859,N_49969);
nor UO_4318 (O_4318,N_49981,N_49946);
nor UO_4319 (O_4319,N_49847,N_49814);
and UO_4320 (O_4320,N_49976,N_49779);
nand UO_4321 (O_4321,N_49834,N_49800);
xnor UO_4322 (O_4322,N_49779,N_49798);
xor UO_4323 (O_4323,N_49921,N_49999);
or UO_4324 (O_4324,N_49767,N_49945);
xor UO_4325 (O_4325,N_49991,N_49943);
nand UO_4326 (O_4326,N_49929,N_49943);
nor UO_4327 (O_4327,N_49917,N_49871);
nand UO_4328 (O_4328,N_49873,N_49816);
or UO_4329 (O_4329,N_49896,N_49812);
nand UO_4330 (O_4330,N_49956,N_49859);
and UO_4331 (O_4331,N_49922,N_49854);
or UO_4332 (O_4332,N_49924,N_49822);
nand UO_4333 (O_4333,N_49835,N_49865);
or UO_4334 (O_4334,N_49761,N_49901);
xor UO_4335 (O_4335,N_49988,N_49800);
nor UO_4336 (O_4336,N_49926,N_49857);
and UO_4337 (O_4337,N_49875,N_49870);
nor UO_4338 (O_4338,N_49849,N_49864);
nand UO_4339 (O_4339,N_49780,N_49828);
nand UO_4340 (O_4340,N_49801,N_49948);
nor UO_4341 (O_4341,N_49910,N_49800);
or UO_4342 (O_4342,N_49870,N_49952);
or UO_4343 (O_4343,N_49874,N_49941);
and UO_4344 (O_4344,N_49991,N_49930);
nor UO_4345 (O_4345,N_49783,N_49988);
or UO_4346 (O_4346,N_49824,N_49867);
and UO_4347 (O_4347,N_49887,N_49937);
and UO_4348 (O_4348,N_49789,N_49853);
xor UO_4349 (O_4349,N_49841,N_49911);
xnor UO_4350 (O_4350,N_49800,N_49898);
nand UO_4351 (O_4351,N_49782,N_49925);
nor UO_4352 (O_4352,N_49774,N_49998);
xnor UO_4353 (O_4353,N_49984,N_49922);
nor UO_4354 (O_4354,N_49997,N_49963);
nand UO_4355 (O_4355,N_49767,N_49823);
xor UO_4356 (O_4356,N_49941,N_49962);
nand UO_4357 (O_4357,N_49850,N_49860);
and UO_4358 (O_4358,N_49984,N_49760);
nand UO_4359 (O_4359,N_49868,N_49831);
nand UO_4360 (O_4360,N_49966,N_49880);
nor UO_4361 (O_4361,N_49814,N_49931);
or UO_4362 (O_4362,N_49933,N_49987);
nor UO_4363 (O_4363,N_49964,N_49785);
or UO_4364 (O_4364,N_49777,N_49896);
nand UO_4365 (O_4365,N_49932,N_49899);
xnor UO_4366 (O_4366,N_49762,N_49841);
nor UO_4367 (O_4367,N_49964,N_49911);
nor UO_4368 (O_4368,N_49787,N_49964);
nand UO_4369 (O_4369,N_49885,N_49903);
xor UO_4370 (O_4370,N_49873,N_49794);
and UO_4371 (O_4371,N_49918,N_49800);
or UO_4372 (O_4372,N_49942,N_49979);
or UO_4373 (O_4373,N_49884,N_49842);
and UO_4374 (O_4374,N_49754,N_49763);
nor UO_4375 (O_4375,N_49912,N_49949);
nand UO_4376 (O_4376,N_49834,N_49849);
and UO_4377 (O_4377,N_49837,N_49842);
xnor UO_4378 (O_4378,N_49923,N_49931);
xor UO_4379 (O_4379,N_49917,N_49764);
xnor UO_4380 (O_4380,N_49836,N_49904);
and UO_4381 (O_4381,N_49962,N_49876);
and UO_4382 (O_4382,N_49945,N_49890);
xnor UO_4383 (O_4383,N_49864,N_49944);
xor UO_4384 (O_4384,N_49828,N_49768);
nor UO_4385 (O_4385,N_49928,N_49988);
or UO_4386 (O_4386,N_49808,N_49855);
and UO_4387 (O_4387,N_49873,N_49925);
nor UO_4388 (O_4388,N_49853,N_49846);
nand UO_4389 (O_4389,N_49888,N_49882);
nor UO_4390 (O_4390,N_49879,N_49818);
or UO_4391 (O_4391,N_49789,N_49814);
or UO_4392 (O_4392,N_49871,N_49776);
and UO_4393 (O_4393,N_49838,N_49848);
nand UO_4394 (O_4394,N_49851,N_49859);
nand UO_4395 (O_4395,N_49776,N_49988);
nand UO_4396 (O_4396,N_49925,N_49986);
xnor UO_4397 (O_4397,N_49845,N_49885);
and UO_4398 (O_4398,N_49779,N_49957);
nor UO_4399 (O_4399,N_49892,N_49750);
nor UO_4400 (O_4400,N_49966,N_49908);
xnor UO_4401 (O_4401,N_49970,N_49777);
and UO_4402 (O_4402,N_49767,N_49752);
xnor UO_4403 (O_4403,N_49823,N_49911);
and UO_4404 (O_4404,N_49761,N_49858);
nand UO_4405 (O_4405,N_49868,N_49900);
or UO_4406 (O_4406,N_49857,N_49791);
and UO_4407 (O_4407,N_49975,N_49888);
xor UO_4408 (O_4408,N_49880,N_49955);
nor UO_4409 (O_4409,N_49903,N_49920);
and UO_4410 (O_4410,N_49862,N_49989);
or UO_4411 (O_4411,N_49840,N_49967);
nor UO_4412 (O_4412,N_49861,N_49937);
nand UO_4413 (O_4413,N_49842,N_49882);
nand UO_4414 (O_4414,N_49824,N_49860);
and UO_4415 (O_4415,N_49879,N_49819);
nand UO_4416 (O_4416,N_49923,N_49985);
or UO_4417 (O_4417,N_49937,N_49818);
nor UO_4418 (O_4418,N_49952,N_49947);
nor UO_4419 (O_4419,N_49789,N_49913);
or UO_4420 (O_4420,N_49782,N_49982);
and UO_4421 (O_4421,N_49766,N_49873);
nand UO_4422 (O_4422,N_49879,N_49944);
xnor UO_4423 (O_4423,N_49878,N_49959);
xor UO_4424 (O_4424,N_49970,N_49830);
nand UO_4425 (O_4425,N_49895,N_49802);
or UO_4426 (O_4426,N_49884,N_49883);
xor UO_4427 (O_4427,N_49912,N_49958);
or UO_4428 (O_4428,N_49808,N_49996);
nand UO_4429 (O_4429,N_49803,N_49854);
and UO_4430 (O_4430,N_49922,N_49812);
nor UO_4431 (O_4431,N_49803,N_49808);
xor UO_4432 (O_4432,N_49776,N_49756);
xor UO_4433 (O_4433,N_49877,N_49999);
nor UO_4434 (O_4434,N_49948,N_49770);
nor UO_4435 (O_4435,N_49904,N_49869);
nor UO_4436 (O_4436,N_49940,N_49967);
nand UO_4437 (O_4437,N_49764,N_49839);
or UO_4438 (O_4438,N_49861,N_49954);
xor UO_4439 (O_4439,N_49874,N_49784);
nand UO_4440 (O_4440,N_49800,N_49922);
nand UO_4441 (O_4441,N_49870,N_49926);
nor UO_4442 (O_4442,N_49817,N_49944);
and UO_4443 (O_4443,N_49978,N_49905);
and UO_4444 (O_4444,N_49920,N_49799);
and UO_4445 (O_4445,N_49919,N_49856);
nor UO_4446 (O_4446,N_49931,N_49852);
xor UO_4447 (O_4447,N_49842,N_49946);
xor UO_4448 (O_4448,N_49885,N_49925);
xor UO_4449 (O_4449,N_49903,N_49914);
or UO_4450 (O_4450,N_49864,N_49861);
nor UO_4451 (O_4451,N_49815,N_49888);
or UO_4452 (O_4452,N_49995,N_49931);
nor UO_4453 (O_4453,N_49935,N_49792);
xnor UO_4454 (O_4454,N_49956,N_49986);
or UO_4455 (O_4455,N_49919,N_49949);
and UO_4456 (O_4456,N_49805,N_49762);
xnor UO_4457 (O_4457,N_49802,N_49847);
and UO_4458 (O_4458,N_49980,N_49799);
nor UO_4459 (O_4459,N_49923,N_49895);
nor UO_4460 (O_4460,N_49959,N_49978);
nor UO_4461 (O_4461,N_49935,N_49949);
nand UO_4462 (O_4462,N_49891,N_49797);
nand UO_4463 (O_4463,N_49816,N_49825);
or UO_4464 (O_4464,N_49934,N_49813);
nor UO_4465 (O_4465,N_49761,N_49757);
nor UO_4466 (O_4466,N_49896,N_49940);
or UO_4467 (O_4467,N_49935,N_49836);
nand UO_4468 (O_4468,N_49962,N_49979);
and UO_4469 (O_4469,N_49858,N_49914);
and UO_4470 (O_4470,N_49906,N_49808);
and UO_4471 (O_4471,N_49829,N_49944);
xor UO_4472 (O_4472,N_49837,N_49974);
nand UO_4473 (O_4473,N_49978,N_49806);
or UO_4474 (O_4474,N_49916,N_49962);
nor UO_4475 (O_4475,N_49943,N_49766);
xor UO_4476 (O_4476,N_49802,N_49860);
nor UO_4477 (O_4477,N_49913,N_49900);
nand UO_4478 (O_4478,N_49952,N_49836);
xnor UO_4479 (O_4479,N_49926,N_49831);
or UO_4480 (O_4480,N_49846,N_49840);
nand UO_4481 (O_4481,N_49957,N_49759);
and UO_4482 (O_4482,N_49780,N_49782);
and UO_4483 (O_4483,N_49752,N_49816);
and UO_4484 (O_4484,N_49913,N_49850);
or UO_4485 (O_4485,N_49808,N_49773);
xor UO_4486 (O_4486,N_49840,N_49994);
nor UO_4487 (O_4487,N_49778,N_49777);
and UO_4488 (O_4488,N_49829,N_49895);
or UO_4489 (O_4489,N_49885,N_49927);
and UO_4490 (O_4490,N_49871,N_49911);
nand UO_4491 (O_4491,N_49937,N_49817);
or UO_4492 (O_4492,N_49973,N_49760);
nand UO_4493 (O_4493,N_49752,N_49978);
or UO_4494 (O_4494,N_49844,N_49768);
nor UO_4495 (O_4495,N_49850,N_49956);
nor UO_4496 (O_4496,N_49908,N_49928);
or UO_4497 (O_4497,N_49981,N_49973);
or UO_4498 (O_4498,N_49924,N_49956);
nand UO_4499 (O_4499,N_49844,N_49821);
and UO_4500 (O_4500,N_49945,N_49943);
nand UO_4501 (O_4501,N_49985,N_49763);
and UO_4502 (O_4502,N_49901,N_49790);
or UO_4503 (O_4503,N_49896,N_49970);
nor UO_4504 (O_4504,N_49928,N_49758);
nand UO_4505 (O_4505,N_49970,N_49775);
nor UO_4506 (O_4506,N_49871,N_49858);
and UO_4507 (O_4507,N_49973,N_49779);
nand UO_4508 (O_4508,N_49852,N_49936);
and UO_4509 (O_4509,N_49950,N_49828);
xor UO_4510 (O_4510,N_49947,N_49893);
or UO_4511 (O_4511,N_49907,N_49763);
or UO_4512 (O_4512,N_49931,N_49959);
or UO_4513 (O_4513,N_49762,N_49951);
xor UO_4514 (O_4514,N_49891,N_49806);
or UO_4515 (O_4515,N_49813,N_49777);
and UO_4516 (O_4516,N_49958,N_49865);
nor UO_4517 (O_4517,N_49845,N_49824);
nor UO_4518 (O_4518,N_49873,N_49773);
nor UO_4519 (O_4519,N_49857,N_49905);
or UO_4520 (O_4520,N_49837,N_49998);
nand UO_4521 (O_4521,N_49979,N_49936);
or UO_4522 (O_4522,N_49896,N_49858);
nand UO_4523 (O_4523,N_49950,N_49962);
nand UO_4524 (O_4524,N_49997,N_49937);
xnor UO_4525 (O_4525,N_49862,N_49821);
nor UO_4526 (O_4526,N_49994,N_49883);
nor UO_4527 (O_4527,N_49807,N_49822);
nand UO_4528 (O_4528,N_49877,N_49906);
nor UO_4529 (O_4529,N_49922,N_49859);
nor UO_4530 (O_4530,N_49949,N_49785);
xor UO_4531 (O_4531,N_49895,N_49859);
nor UO_4532 (O_4532,N_49917,N_49762);
and UO_4533 (O_4533,N_49905,N_49907);
nand UO_4534 (O_4534,N_49895,N_49981);
and UO_4535 (O_4535,N_49903,N_49986);
and UO_4536 (O_4536,N_49873,N_49860);
or UO_4537 (O_4537,N_49754,N_49971);
or UO_4538 (O_4538,N_49967,N_49818);
nand UO_4539 (O_4539,N_49849,N_49894);
and UO_4540 (O_4540,N_49823,N_49875);
or UO_4541 (O_4541,N_49928,N_49754);
or UO_4542 (O_4542,N_49762,N_49977);
nand UO_4543 (O_4543,N_49949,N_49996);
nand UO_4544 (O_4544,N_49786,N_49995);
and UO_4545 (O_4545,N_49754,N_49976);
xnor UO_4546 (O_4546,N_49832,N_49993);
nor UO_4547 (O_4547,N_49881,N_49861);
nor UO_4548 (O_4548,N_49945,N_49914);
nand UO_4549 (O_4549,N_49782,N_49759);
xor UO_4550 (O_4550,N_49934,N_49928);
xor UO_4551 (O_4551,N_49971,N_49769);
nand UO_4552 (O_4552,N_49954,N_49772);
nor UO_4553 (O_4553,N_49983,N_49884);
and UO_4554 (O_4554,N_49846,N_49892);
nand UO_4555 (O_4555,N_49753,N_49983);
and UO_4556 (O_4556,N_49805,N_49881);
and UO_4557 (O_4557,N_49897,N_49765);
xnor UO_4558 (O_4558,N_49794,N_49887);
and UO_4559 (O_4559,N_49973,N_49906);
and UO_4560 (O_4560,N_49980,N_49865);
xor UO_4561 (O_4561,N_49999,N_49933);
xor UO_4562 (O_4562,N_49830,N_49846);
nand UO_4563 (O_4563,N_49885,N_49842);
nand UO_4564 (O_4564,N_49897,N_49814);
nand UO_4565 (O_4565,N_49937,N_49822);
nand UO_4566 (O_4566,N_49951,N_49847);
xnor UO_4567 (O_4567,N_49986,N_49955);
or UO_4568 (O_4568,N_49786,N_49781);
nand UO_4569 (O_4569,N_49792,N_49923);
nor UO_4570 (O_4570,N_49915,N_49908);
or UO_4571 (O_4571,N_49799,N_49967);
xnor UO_4572 (O_4572,N_49962,N_49844);
and UO_4573 (O_4573,N_49840,N_49785);
xor UO_4574 (O_4574,N_49785,N_49959);
nor UO_4575 (O_4575,N_49898,N_49910);
nor UO_4576 (O_4576,N_49800,N_49965);
or UO_4577 (O_4577,N_49931,N_49988);
and UO_4578 (O_4578,N_49914,N_49798);
nand UO_4579 (O_4579,N_49765,N_49807);
xnor UO_4580 (O_4580,N_49845,N_49870);
xnor UO_4581 (O_4581,N_49940,N_49975);
xnor UO_4582 (O_4582,N_49994,N_49821);
nor UO_4583 (O_4583,N_49829,N_49863);
xor UO_4584 (O_4584,N_49818,N_49840);
or UO_4585 (O_4585,N_49966,N_49804);
xor UO_4586 (O_4586,N_49994,N_49990);
or UO_4587 (O_4587,N_49815,N_49988);
nand UO_4588 (O_4588,N_49782,N_49872);
or UO_4589 (O_4589,N_49778,N_49875);
nand UO_4590 (O_4590,N_49889,N_49788);
or UO_4591 (O_4591,N_49789,N_49906);
nand UO_4592 (O_4592,N_49859,N_49896);
or UO_4593 (O_4593,N_49981,N_49862);
or UO_4594 (O_4594,N_49781,N_49839);
nand UO_4595 (O_4595,N_49910,N_49860);
or UO_4596 (O_4596,N_49908,N_49827);
nor UO_4597 (O_4597,N_49913,N_49965);
nand UO_4598 (O_4598,N_49851,N_49879);
and UO_4599 (O_4599,N_49752,N_49838);
nor UO_4600 (O_4600,N_49852,N_49806);
xor UO_4601 (O_4601,N_49986,N_49997);
xor UO_4602 (O_4602,N_49788,N_49800);
nor UO_4603 (O_4603,N_49832,N_49874);
or UO_4604 (O_4604,N_49839,N_49876);
nor UO_4605 (O_4605,N_49951,N_49949);
nand UO_4606 (O_4606,N_49772,N_49983);
and UO_4607 (O_4607,N_49787,N_49844);
xnor UO_4608 (O_4608,N_49785,N_49989);
xnor UO_4609 (O_4609,N_49797,N_49921);
nand UO_4610 (O_4610,N_49825,N_49940);
nor UO_4611 (O_4611,N_49939,N_49973);
or UO_4612 (O_4612,N_49923,N_49933);
nor UO_4613 (O_4613,N_49950,N_49800);
xor UO_4614 (O_4614,N_49924,N_49928);
nor UO_4615 (O_4615,N_49969,N_49979);
nand UO_4616 (O_4616,N_49963,N_49928);
or UO_4617 (O_4617,N_49963,N_49794);
xor UO_4618 (O_4618,N_49970,N_49766);
nor UO_4619 (O_4619,N_49836,N_49888);
nand UO_4620 (O_4620,N_49899,N_49871);
xor UO_4621 (O_4621,N_49878,N_49894);
nand UO_4622 (O_4622,N_49908,N_49927);
nor UO_4623 (O_4623,N_49869,N_49782);
or UO_4624 (O_4624,N_49941,N_49886);
nand UO_4625 (O_4625,N_49963,N_49803);
and UO_4626 (O_4626,N_49822,N_49887);
xnor UO_4627 (O_4627,N_49982,N_49796);
nand UO_4628 (O_4628,N_49758,N_49760);
nor UO_4629 (O_4629,N_49973,N_49900);
nor UO_4630 (O_4630,N_49977,N_49921);
xnor UO_4631 (O_4631,N_49843,N_49870);
or UO_4632 (O_4632,N_49901,N_49793);
and UO_4633 (O_4633,N_49881,N_49755);
nand UO_4634 (O_4634,N_49798,N_49893);
and UO_4635 (O_4635,N_49795,N_49992);
xor UO_4636 (O_4636,N_49782,N_49756);
and UO_4637 (O_4637,N_49894,N_49989);
nor UO_4638 (O_4638,N_49998,N_49881);
xor UO_4639 (O_4639,N_49764,N_49898);
or UO_4640 (O_4640,N_49844,N_49823);
nand UO_4641 (O_4641,N_49946,N_49797);
nor UO_4642 (O_4642,N_49978,N_49871);
xnor UO_4643 (O_4643,N_49994,N_49827);
or UO_4644 (O_4644,N_49894,N_49824);
and UO_4645 (O_4645,N_49830,N_49944);
or UO_4646 (O_4646,N_49840,N_49850);
or UO_4647 (O_4647,N_49769,N_49999);
nor UO_4648 (O_4648,N_49931,N_49841);
xnor UO_4649 (O_4649,N_49829,N_49912);
nand UO_4650 (O_4650,N_49846,N_49975);
xnor UO_4651 (O_4651,N_49868,N_49991);
or UO_4652 (O_4652,N_49787,N_49815);
and UO_4653 (O_4653,N_49925,N_49918);
nand UO_4654 (O_4654,N_49799,N_49777);
and UO_4655 (O_4655,N_49982,N_49996);
or UO_4656 (O_4656,N_49776,N_49891);
xnor UO_4657 (O_4657,N_49865,N_49814);
nand UO_4658 (O_4658,N_49837,N_49803);
or UO_4659 (O_4659,N_49865,N_49802);
nor UO_4660 (O_4660,N_49925,N_49842);
xor UO_4661 (O_4661,N_49963,N_49979);
nand UO_4662 (O_4662,N_49810,N_49867);
nor UO_4663 (O_4663,N_49970,N_49921);
nor UO_4664 (O_4664,N_49792,N_49755);
nand UO_4665 (O_4665,N_49976,N_49847);
nand UO_4666 (O_4666,N_49954,N_49846);
and UO_4667 (O_4667,N_49955,N_49908);
or UO_4668 (O_4668,N_49924,N_49983);
or UO_4669 (O_4669,N_49820,N_49830);
or UO_4670 (O_4670,N_49975,N_49963);
or UO_4671 (O_4671,N_49931,N_49838);
xnor UO_4672 (O_4672,N_49882,N_49822);
nor UO_4673 (O_4673,N_49936,N_49795);
xor UO_4674 (O_4674,N_49974,N_49873);
xnor UO_4675 (O_4675,N_49820,N_49755);
nor UO_4676 (O_4676,N_49824,N_49769);
nand UO_4677 (O_4677,N_49988,N_49769);
nor UO_4678 (O_4678,N_49825,N_49851);
nor UO_4679 (O_4679,N_49784,N_49870);
nand UO_4680 (O_4680,N_49951,N_49758);
nand UO_4681 (O_4681,N_49806,N_49980);
or UO_4682 (O_4682,N_49772,N_49827);
xnor UO_4683 (O_4683,N_49874,N_49776);
or UO_4684 (O_4684,N_49976,N_49760);
or UO_4685 (O_4685,N_49890,N_49998);
xnor UO_4686 (O_4686,N_49968,N_49802);
nor UO_4687 (O_4687,N_49815,N_49926);
or UO_4688 (O_4688,N_49911,N_49809);
and UO_4689 (O_4689,N_49789,N_49925);
xor UO_4690 (O_4690,N_49877,N_49843);
xnor UO_4691 (O_4691,N_49930,N_49898);
xor UO_4692 (O_4692,N_49889,N_49812);
xor UO_4693 (O_4693,N_49956,N_49869);
or UO_4694 (O_4694,N_49848,N_49875);
or UO_4695 (O_4695,N_49878,N_49874);
nand UO_4696 (O_4696,N_49907,N_49856);
xnor UO_4697 (O_4697,N_49881,N_49862);
and UO_4698 (O_4698,N_49876,N_49912);
or UO_4699 (O_4699,N_49980,N_49902);
or UO_4700 (O_4700,N_49901,N_49899);
xnor UO_4701 (O_4701,N_49867,N_49816);
or UO_4702 (O_4702,N_49778,N_49903);
or UO_4703 (O_4703,N_49782,N_49835);
or UO_4704 (O_4704,N_49923,N_49830);
nand UO_4705 (O_4705,N_49802,N_49945);
xor UO_4706 (O_4706,N_49787,N_49768);
xor UO_4707 (O_4707,N_49932,N_49760);
nand UO_4708 (O_4708,N_49944,N_49881);
or UO_4709 (O_4709,N_49788,N_49895);
nor UO_4710 (O_4710,N_49962,N_49910);
and UO_4711 (O_4711,N_49854,N_49976);
and UO_4712 (O_4712,N_49786,N_49828);
xnor UO_4713 (O_4713,N_49787,N_49761);
xnor UO_4714 (O_4714,N_49767,N_49925);
or UO_4715 (O_4715,N_49825,N_49836);
nor UO_4716 (O_4716,N_49962,N_49792);
and UO_4717 (O_4717,N_49973,N_49891);
xnor UO_4718 (O_4718,N_49884,N_49843);
nand UO_4719 (O_4719,N_49920,N_49953);
or UO_4720 (O_4720,N_49884,N_49756);
nor UO_4721 (O_4721,N_49975,N_49972);
and UO_4722 (O_4722,N_49805,N_49865);
xnor UO_4723 (O_4723,N_49964,N_49779);
and UO_4724 (O_4724,N_49827,N_49877);
xnor UO_4725 (O_4725,N_49825,N_49818);
and UO_4726 (O_4726,N_49752,N_49984);
nand UO_4727 (O_4727,N_49989,N_49811);
nor UO_4728 (O_4728,N_49787,N_49839);
nor UO_4729 (O_4729,N_49943,N_49836);
nand UO_4730 (O_4730,N_49992,N_49981);
nor UO_4731 (O_4731,N_49751,N_49936);
nand UO_4732 (O_4732,N_49892,N_49995);
nor UO_4733 (O_4733,N_49857,N_49780);
or UO_4734 (O_4734,N_49769,N_49918);
xnor UO_4735 (O_4735,N_49979,N_49867);
nand UO_4736 (O_4736,N_49760,N_49781);
nand UO_4737 (O_4737,N_49822,N_49830);
xnor UO_4738 (O_4738,N_49860,N_49931);
or UO_4739 (O_4739,N_49937,N_49869);
nand UO_4740 (O_4740,N_49887,N_49862);
and UO_4741 (O_4741,N_49936,N_49912);
or UO_4742 (O_4742,N_49946,N_49920);
nand UO_4743 (O_4743,N_49953,N_49944);
nand UO_4744 (O_4744,N_49979,N_49822);
nor UO_4745 (O_4745,N_49773,N_49839);
nand UO_4746 (O_4746,N_49996,N_49945);
nand UO_4747 (O_4747,N_49904,N_49938);
or UO_4748 (O_4748,N_49790,N_49781);
and UO_4749 (O_4749,N_49873,N_49820);
xnor UO_4750 (O_4750,N_49818,N_49752);
xor UO_4751 (O_4751,N_49755,N_49752);
nand UO_4752 (O_4752,N_49770,N_49843);
xor UO_4753 (O_4753,N_49987,N_49807);
xor UO_4754 (O_4754,N_49839,N_49859);
nor UO_4755 (O_4755,N_49956,N_49878);
or UO_4756 (O_4756,N_49894,N_49866);
xor UO_4757 (O_4757,N_49836,N_49975);
and UO_4758 (O_4758,N_49861,N_49936);
or UO_4759 (O_4759,N_49756,N_49989);
nand UO_4760 (O_4760,N_49963,N_49835);
xor UO_4761 (O_4761,N_49954,N_49974);
and UO_4762 (O_4762,N_49954,N_49978);
or UO_4763 (O_4763,N_49976,N_49935);
or UO_4764 (O_4764,N_49896,N_49854);
or UO_4765 (O_4765,N_49798,N_49999);
nand UO_4766 (O_4766,N_49999,N_49944);
nand UO_4767 (O_4767,N_49804,N_49976);
xnor UO_4768 (O_4768,N_49784,N_49952);
and UO_4769 (O_4769,N_49897,N_49848);
nor UO_4770 (O_4770,N_49817,N_49819);
nand UO_4771 (O_4771,N_49960,N_49760);
xor UO_4772 (O_4772,N_49758,N_49846);
and UO_4773 (O_4773,N_49979,N_49790);
nand UO_4774 (O_4774,N_49983,N_49851);
or UO_4775 (O_4775,N_49940,N_49768);
nand UO_4776 (O_4776,N_49919,N_49772);
nand UO_4777 (O_4777,N_49908,N_49834);
xor UO_4778 (O_4778,N_49823,N_49763);
nor UO_4779 (O_4779,N_49959,N_49958);
and UO_4780 (O_4780,N_49848,N_49998);
nor UO_4781 (O_4781,N_49992,N_49750);
xor UO_4782 (O_4782,N_49877,N_49895);
or UO_4783 (O_4783,N_49794,N_49993);
nand UO_4784 (O_4784,N_49866,N_49817);
xnor UO_4785 (O_4785,N_49774,N_49810);
and UO_4786 (O_4786,N_49800,N_49772);
nor UO_4787 (O_4787,N_49971,N_49805);
nor UO_4788 (O_4788,N_49772,N_49880);
or UO_4789 (O_4789,N_49931,N_49848);
or UO_4790 (O_4790,N_49921,N_49904);
or UO_4791 (O_4791,N_49852,N_49950);
nor UO_4792 (O_4792,N_49885,N_49840);
or UO_4793 (O_4793,N_49984,N_49966);
xnor UO_4794 (O_4794,N_49847,N_49831);
xor UO_4795 (O_4795,N_49931,N_49774);
or UO_4796 (O_4796,N_49977,N_49770);
nor UO_4797 (O_4797,N_49988,N_49793);
nand UO_4798 (O_4798,N_49880,N_49916);
or UO_4799 (O_4799,N_49894,N_49955);
xor UO_4800 (O_4800,N_49925,N_49818);
nand UO_4801 (O_4801,N_49801,N_49833);
or UO_4802 (O_4802,N_49883,N_49752);
and UO_4803 (O_4803,N_49802,N_49836);
and UO_4804 (O_4804,N_49853,N_49866);
and UO_4805 (O_4805,N_49948,N_49983);
nand UO_4806 (O_4806,N_49949,N_49827);
nand UO_4807 (O_4807,N_49752,N_49991);
and UO_4808 (O_4808,N_49790,N_49808);
or UO_4809 (O_4809,N_49982,N_49825);
nand UO_4810 (O_4810,N_49899,N_49783);
xnor UO_4811 (O_4811,N_49779,N_49753);
or UO_4812 (O_4812,N_49981,N_49941);
nand UO_4813 (O_4813,N_49759,N_49943);
and UO_4814 (O_4814,N_49762,N_49930);
nand UO_4815 (O_4815,N_49975,N_49992);
nor UO_4816 (O_4816,N_49888,N_49939);
nor UO_4817 (O_4817,N_49758,N_49822);
nand UO_4818 (O_4818,N_49866,N_49908);
xnor UO_4819 (O_4819,N_49933,N_49828);
xor UO_4820 (O_4820,N_49977,N_49832);
and UO_4821 (O_4821,N_49878,N_49897);
nor UO_4822 (O_4822,N_49990,N_49776);
and UO_4823 (O_4823,N_49878,N_49832);
and UO_4824 (O_4824,N_49780,N_49997);
or UO_4825 (O_4825,N_49839,N_49793);
and UO_4826 (O_4826,N_49876,N_49856);
nor UO_4827 (O_4827,N_49784,N_49822);
or UO_4828 (O_4828,N_49905,N_49765);
and UO_4829 (O_4829,N_49872,N_49812);
nor UO_4830 (O_4830,N_49916,N_49996);
nor UO_4831 (O_4831,N_49760,N_49979);
or UO_4832 (O_4832,N_49783,N_49753);
and UO_4833 (O_4833,N_49843,N_49962);
and UO_4834 (O_4834,N_49885,N_49853);
or UO_4835 (O_4835,N_49935,N_49807);
and UO_4836 (O_4836,N_49772,N_49854);
or UO_4837 (O_4837,N_49984,N_49988);
and UO_4838 (O_4838,N_49981,N_49945);
and UO_4839 (O_4839,N_49789,N_49892);
xor UO_4840 (O_4840,N_49939,N_49817);
or UO_4841 (O_4841,N_49758,N_49967);
nor UO_4842 (O_4842,N_49819,N_49824);
nand UO_4843 (O_4843,N_49844,N_49834);
nand UO_4844 (O_4844,N_49902,N_49985);
nand UO_4845 (O_4845,N_49948,N_49818);
xor UO_4846 (O_4846,N_49931,N_49784);
or UO_4847 (O_4847,N_49974,N_49788);
and UO_4848 (O_4848,N_49976,N_49866);
and UO_4849 (O_4849,N_49915,N_49835);
or UO_4850 (O_4850,N_49891,N_49790);
xnor UO_4851 (O_4851,N_49904,N_49760);
or UO_4852 (O_4852,N_49869,N_49793);
or UO_4853 (O_4853,N_49959,N_49899);
xor UO_4854 (O_4854,N_49754,N_49819);
nand UO_4855 (O_4855,N_49822,N_49763);
nor UO_4856 (O_4856,N_49964,N_49872);
nand UO_4857 (O_4857,N_49980,N_49927);
nand UO_4858 (O_4858,N_49809,N_49800);
xor UO_4859 (O_4859,N_49792,N_49897);
nand UO_4860 (O_4860,N_49930,N_49871);
xor UO_4861 (O_4861,N_49861,N_49856);
and UO_4862 (O_4862,N_49781,N_49794);
and UO_4863 (O_4863,N_49781,N_49939);
and UO_4864 (O_4864,N_49865,N_49791);
xnor UO_4865 (O_4865,N_49910,N_49835);
and UO_4866 (O_4866,N_49803,N_49879);
nor UO_4867 (O_4867,N_49754,N_49901);
nor UO_4868 (O_4868,N_49836,N_49976);
or UO_4869 (O_4869,N_49794,N_49954);
xnor UO_4870 (O_4870,N_49808,N_49890);
nand UO_4871 (O_4871,N_49791,N_49877);
nor UO_4872 (O_4872,N_49831,N_49998);
or UO_4873 (O_4873,N_49860,N_49895);
or UO_4874 (O_4874,N_49990,N_49852);
nand UO_4875 (O_4875,N_49997,N_49934);
or UO_4876 (O_4876,N_49891,N_49868);
xor UO_4877 (O_4877,N_49758,N_49987);
nand UO_4878 (O_4878,N_49835,N_49750);
or UO_4879 (O_4879,N_49964,N_49874);
xor UO_4880 (O_4880,N_49814,N_49918);
nand UO_4881 (O_4881,N_49883,N_49919);
nor UO_4882 (O_4882,N_49758,N_49776);
or UO_4883 (O_4883,N_49775,N_49848);
xnor UO_4884 (O_4884,N_49929,N_49876);
nor UO_4885 (O_4885,N_49754,N_49988);
nand UO_4886 (O_4886,N_49782,N_49866);
xor UO_4887 (O_4887,N_49894,N_49800);
nand UO_4888 (O_4888,N_49766,N_49923);
and UO_4889 (O_4889,N_49863,N_49827);
nand UO_4890 (O_4890,N_49947,N_49759);
xor UO_4891 (O_4891,N_49866,N_49906);
xor UO_4892 (O_4892,N_49755,N_49945);
nor UO_4893 (O_4893,N_49927,N_49777);
nand UO_4894 (O_4894,N_49944,N_49992);
or UO_4895 (O_4895,N_49847,N_49797);
nand UO_4896 (O_4896,N_49796,N_49953);
and UO_4897 (O_4897,N_49779,N_49773);
or UO_4898 (O_4898,N_49902,N_49915);
xor UO_4899 (O_4899,N_49976,N_49927);
nor UO_4900 (O_4900,N_49979,N_49955);
nor UO_4901 (O_4901,N_49750,N_49865);
nor UO_4902 (O_4902,N_49806,N_49988);
nor UO_4903 (O_4903,N_49943,N_49760);
nand UO_4904 (O_4904,N_49765,N_49804);
nand UO_4905 (O_4905,N_49794,N_49893);
nor UO_4906 (O_4906,N_49978,N_49887);
and UO_4907 (O_4907,N_49911,N_49792);
or UO_4908 (O_4908,N_49844,N_49831);
and UO_4909 (O_4909,N_49758,N_49865);
and UO_4910 (O_4910,N_49897,N_49839);
nand UO_4911 (O_4911,N_49898,N_49896);
nand UO_4912 (O_4912,N_49930,N_49771);
nand UO_4913 (O_4913,N_49977,N_49860);
nor UO_4914 (O_4914,N_49961,N_49915);
and UO_4915 (O_4915,N_49783,N_49878);
nor UO_4916 (O_4916,N_49908,N_49849);
xnor UO_4917 (O_4917,N_49849,N_49901);
or UO_4918 (O_4918,N_49829,N_49898);
xor UO_4919 (O_4919,N_49888,N_49852);
nand UO_4920 (O_4920,N_49959,N_49951);
nor UO_4921 (O_4921,N_49859,N_49877);
or UO_4922 (O_4922,N_49779,N_49849);
xnor UO_4923 (O_4923,N_49988,N_49862);
and UO_4924 (O_4924,N_49841,N_49784);
nor UO_4925 (O_4925,N_49845,N_49857);
or UO_4926 (O_4926,N_49920,N_49784);
or UO_4927 (O_4927,N_49978,N_49864);
nor UO_4928 (O_4928,N_49766,N_49867);
xor UO_4929 (O_4929,N_49973,N_49753);
xnor UO_4930 (O_4930,N_49916,N_49850);
and UO_4931 (O_4931,N_49772,N_49753);
nand UO_4932 (O_4932,N_49947,N_49881);
nor UO_4933 (O_4933,N_49930,N_49826);
and UO_4934 (O_4934,N_49896,N_49806);
or UO_4935 (O_4935,N_49853,N_49813);
and UO_4936 (O_4936,N_49932,N_49809);
nor UO_4937 (O_4937,N_49800,N_49766);
nand UO_4938 (O_4938,N_49954,N_49936);
xor UO_4939 (O_4939,N_49932,N_49921);
nor UO_4940 (O_4940,N_49764,N_49927);
xnor UO_4941 (O_4941,N_49797,N_49815);
nor UO_4942 (O_4942,N_49985,N_49784);
nand UO_4943 (O_4943,N_49838,N_49822);
or UO_4944 (O_4944,N_49924,N_49926);
nand UO_4945 (O_4945,N_49872,N_49816);
or UO_4946 (O_4946,N_49940,N_49762);
nand UO_4947 (O_4947,N_49774,N_49873);
or UO_4948 (O_4948,N_49791,N_49886);
xnor UO_4949 (O_4949,N_49893,N_49859);
nand UO_4950 (O_4950,N_49888,N_49804);
nor UO_4951 (O_4951,N_49750,N_49854);
or UO_4952 (O_4952,N_49761,N_49840);
nand UO_4953 (O_4953,N_49754,N_49958);
nor UO_4954 (O_4954,N_49919,N_49785);
xnor UO_4955 (O_4955,N_49926,N_49987);
and UO_4956 (O_4956,N_49777,N_49964);
or UO_4957 (O_4957,N_49798,N_49852);
nor UO_4958 (O_4958,N_49873,N_49781);
xor UO_4959 (O_4959,N_49812,N_49979);
xnor UO_4960 (O_4960,N_49983,N_49832);
nand UO_4961 (O_4961,N_49755,N_49754);
or UO_4962 (O_4962,N_49806,N_49950);
nor UO_4963 (O_4963,N_49840,N_49796);
xor UO_4964 (O_4964,N_49810,N_49985);
xor UO_4965 (O_4965,N_49902,N_49785);
nor UO_4966 (O_4966,N_49813,N_49841);
xor UO_4967 (O_4967,N_49965,N_49860);
nand UO_4968 (O_4968,N_49761,N_49925);
nor UO_4969 (O_4969,N_49907,N_49872);
or UO_4970 (O_4970,N_49952,N_49984);
nand UO_4971 (O_4971,N_49817,N_49853);
xor UO_4972 (O_4972,N_49789,N_49865);
nand UO_4973 (O_4973,N_49919,N_49769);
or UO_4974 (O_4974,N_49959,N_49757);
xnor UO_4975 (O_4975,N_49834,N_49958);
xnor UO_4976 (O_4976,N_49847,N_49845);
nor UO_4977 (O_4977,N_49876,N_49954);
nor UO_4978 (O_4978,N_49786,N_49919);
nand UO_4979 (O_4979,N_49826,N_49975);
nand UO_4980 (O_4980,N_49854,N_49765);
xnor UO_4981 (O_4981,N_49896,N_49794);
and UO_4982 (O_4982,N_49950,N_49851);
and UO_4983 (O_4983,N_49955,N_49914);
xnor UO_4984 (O_4984,N_49958,N_49985);
xnor UO_4985 (O_4985,N_49799,N_49793);
nand UO_4986 (O_4986,N_49995,N_49833);
nand UO_4987 (O_4987,N_49778,N_49785);
and UO_4988 (O_4988,N_49880,N_49870);
nor UO_4989 (O_4989,N_49759,N_49793);
and UO_4990 (O_4990,N_49933,N_49814);
nand UO_4991 (O_4991,N_49833,N_49837);
or UO_4992 (O_4992,N_49771,N_49804);
or UO_4993 (O_4993,N_49897,N_49871);
or UO_4994 (O_4994,N_49962,N_49875);
nand UO_4995 (O_4995,N_49961,N_49836);
and UO_4996 (O_4996,N_49871,N_49888);
xor UO_4997 (O_4997,N_49903,N_49770);
and UO_4998 (O_4998,N_49917,N_49786);
or UO_4999 (O_4999,N_49943,N_49998);
endmodule