module basic_500_3000_500_40_levels_10xor_3(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
nand U0 (N_0,In_47,In_388);
nand U1 (N_1,In_373,In_144);
nor U2 (N_2,In_495,In_42);
nand U3 (N_3,In_151,In_405);
and U4 (N_4,In_398,In_272);
nor U5 (N_5,In_204,In_174);
and U6 (N_6,In_317,In_63);
nor U7 (N_7,In_239,In_200);
or U8 (N_8,In_143,In_43);
and U9 (N_9,In_376,In_220);
nor U10 (N_10,In_154,In_358);
nor U11 (N_11,In_392,In_491);
or U12 (N_12,In_326,In_494);
nand U13 (N_13,In_360,In_250);
or U14 (N_14,In_449,In_319);
or U15 (N_15,In_104,In_114);
nor U16 (N_16,In_247,In_390);
nor U17 (N_17,In_485,In_196);
and U18 (N_18,In_311,In_141);
and U19 (N_19,In_178,In_455);
xnor U20 (N_20,In_87,In_347);
and U21 (N_21,In_349,In_70);
nor U22 (N_22,In_264,In_411);
nand U23 (N_23,In_425,In_75);
and U24 (N_24,In_300,In_28);
and U25 (N_25,In_412,In_5);
nor U26 (N_26,In_361,In_402);
xnor U27 (N_27,In_150,In_122);
xor U28 (N_28,In_216,In_7);
nor U29 (N_29,In_110,In_436);
and U30 (N_30,In_96,In_127);
xnor U31 (N_31,In_18,In_108);
nor U32 (N_32,In_474,In_266);
xnor U33 (N_33,In_168,In_153);
xor U34 (N_34,In_223,In_354);
or U35 (N_35,In_331,In_164);
and U36 (N_36,In_327,In_499);
nor U37 (N_37,In_130,In_212);
or U38 (N_38,In_3,In_440);
or U39 (N_39,In_125,In_83);
nand U40 (N_40,In_41,In_242);
nor U41 (N_41,In_386,In_383);
or U42 (N_42,In_337,In_246);
xor U43 (N_43,In_427,In_470);
nand U44 (N_44,In_410,In_255);
or U45 (N_45,In_172,In_393);
nor U46 (N_46,In_456,In_58);
or U47 (N_47,In_226,In_123);
xor U48 (N_48,In_240,In_290);
xor U49 (N_49,In_184,In_36);
nand U50 (N_50,In_461,In_355);
and U51 (N_51,In_126,In_419);
and U52 (N_52,In_161,In_147);
and U53 (N_53,In_418,In_316);
nor U54 (N_54,In_353,In_265);
nor U55 (N_55,In_9,In_351);
xor U56 (N_56,In_356,In_400);
xnor U57 (N_57,In_284,In_345);
nand U58 (N_58,In_341,In_421);
and U59 (N_59,In_352,In_384);
or U60 (N_60,In_89,In_14);
or U61 (N_61,In_0,In_391);
nand U62 (N_62,In_447,In_237);
nand U63 (N_63,In_112,In_468);
or U64 (N_64,In_395,In_165);
nand U65 (N_65,In_396,In_403);
xor U66 (N_66,In_236,In_78);
xnor U67 (N_67,In_51,In_397);
xnor U68 (N_68,In_282,In_180);
xor U69 (N_69,In_378,In_322);
xor U70 (N_70,In_285,In_404);
xor U71 (N_71,In_364,In_118);
and U72 (N_72,In_206,In_314);
and U73 (N_73,In_371,In_339);
nor U74 (N_74,In_4,In_334);
xnor U75 (N_75,In_202,In_105);
nor U76 (N_76,N_9,In_399);
nor U77 (N_77,In_72,In_203);
nor U78 (N_78,In_234,In_38);
xnor U79 (N_79,N_2,In_169);
and U80 (N_80,N_43,In_444);
nor U81 (N_81,In_305,In_1);
nor U82 (N_82,In_273,N_41);
and U83 (N_83,In_170,In_465);
and U84 (N_84,In_17,In_407);
or U85 (N_85,N_55,In_79);
nand U86 (N_86,In_340,N_53);
nor U87 (N_87,In_61,In_363);
xor U88 (N_88,In_77,In_294);
or U89 (N_89,N_71,In_37);
nand U90 (N_90,In_477,In_16);
and U91 (N_91,N_61,N_29);
nor U92 (N_92,In_156,In_472);
xnor U93 (N_93,In_310,In_35);
and U94 (N_94,In_424,In_454);
or U95 (N_95,In_128,In_306);
and U96 (N_96,In_119,In_475);
xnor U97 (N_97,In_6,In_298);
nor U98 (N_98,In_34,In_365);
nand U99 (N_99,N_12,N_63);
xnor U100 (N_100,In_227,In_244);
and U101 (N_101,In_158,N_50);
or U102 (N_102,N_18,In_377);
nand U103 (N_103,In_445,In_233);
nand U104 (N_104,In_320,N_16);
xnor U105 (N_105,In_323,In_409);
and U106 (N_106,In_488,In_496);
or U107 (N_107,In_271,In_73);
nand U108 (N_108,N_31,In_232);
or U109 (N_109,N_45,N_1);
or U110 (N_110,In_80,In_243);
nand U111 (N_111,In_288,In_394);
or U112 (N_112,In_101,In_277);
or U113 (N_113,In_338,In_434);
nand U114 (N_114,In_189,In_133);
or U115 (N_115,In_201,In_480);
and U116 (N_116,In_177,In_498);
and U117 (N_117,In_92,In_374);
and U118 (N_118,In_65,N_6);
and U119 (N_119,In_56,In_160);
nand U120 (N_120,In_219,N_36);
and U121 (N_121,In_329,In_120);
and U122 (N_122,In_45,In_90);
or U123 (N_123,In_259,In_413);
nor U124 (N_124,N_10,In_224);
or U125 (N_125,N_8,In_218);
nand U126 (N_126,In_382,In_489);
or U127 (N_127,In_457,In_414);
nand U128 (N_128,In_406,In_245);
or U129 (N_129,In_109,N_0);
nand U130 (N_130,In_192,In_380);
or U131 (N_131,In_381,In_46);
or U132 (N_132,In_346,In_486);
and U133 (N_133,In_117,In_71);
xnor U134 (N_134,In_31,N_21);
nor U135 (N_135,In_60,In_401);
or U136 (N_136,In_389,In_370);
xor U137 (N_137,In_208,In_278);
xnor U138 (N_138,In_286,In_32);
xor U139 (N_139,N_27,In_48);
and U140 (N_140,In_124,In_283);
nand U141 (N_141,In_131,N_5);
nor U142 (N_142,In_439,In_52);
and U143 (N_143,In_162,In_94);
or U144 (N_144,In_387,In_299);
or U145 (N_145,N_26,In_121);
xnor U146 (N_146,In_179,In_258);
nor U147 (N_147,In_30,In_279);
nand U148 (N_148,N_19,N_20);
and U149 (N_149,In_59,In_205);
or U150 (N_150,N_104,In_307);
or U151 (N_151,In_438,In_10);
or U152 (N_152,In_187,In_13);
nor U153 (N_153,N_49,N_114);
or U154 (N_154,N_137,In_228);
nor U155 (N_155,In_93,In_473);
nand U156 (N_156,In_487,In_254);
nand U157 (N_157,In_12,In_420);
and U158 (N_158,In_263,N_40);
nor U159 (N_159,In_483,In_238);
xnor U160 (N_160,N_109,In_280);
or U161 (N_161,In_111,In_188);
or U162 (N_162,N_51,N_149);
xor U163 (N_163,N_143,In_183);
xnor U164 (N_164,N_128,N_44);
xor U165 (N_165,N_87,In_350);
or U166 (N_166,N_3,In_462);
nor U167 (N_167,In_357,N_94);
nand U168 (N_168,N_102,In_336);
and U169 (N_169,N_81,In_136);
or U170 (N_170,In_152,In_163);
xor U171 (N_171,In_281,N_115);
and U172 (N_172,In_186,In_146);
xnor U173 (N_173,In_251,In_292);
nor U174 (N_174,In_301,In_287);
xnor U175 (N_175,In_29,In_481);
and U176 (N_176,In_441,In_459);
and U177 (N_177,N_48,In_484);
and U178 (N_178,In_215,In_262);
xnor U179 (N_179,In_21,N_85);
or U180 (N_180,In_466,In_478);
xor U181 (N_181,In_318,In_325);
nand U182 (N_182,N_54,N_126);
nor U183 (N_183,In_39,In_214);
or U184 (N_184,In_241,In_157);
xor U185 (N_185,N_37,In_197);
nor U186 (N_186,In_88,In_23);
nand U187 (N_187,In_417,In_20);
and U188 (N_188,N_56,In_84);
nand U189 (N_189,N_141,In_275);
nand U190 (N_190,In_74,In_348);
xor U191 (N_191,N_64,N_136);
and U192 (N_192,In_268,In_432);
and U193 (N_193,N_70,In_359);
or U194 (N_194,In_295,In_385);
nor U195 (N_195,In_82,N_17);
nand U196 (N_196,In_230,N_25);
nor U197 (N_197,In_100,In_362);
and U198 (N_198,N_146,N_123);
xor U199 (N_199,In_463,In_57);
xnor U200 (N_200,In_257,In_423);
or U201 (N_201,In_293,In_443);
and U202 (N_202,In_54,In_67);
nor U203 (N_203,In_139,In_81);
xnor U204 (N_204,In_191,N_116);
or U205 (N_205,N_148,N_91);
or U206 (N_206,N_147,In_68);
xnor U207 (N_207,In_332,N_105);
and U208 (N_208,In_95,N_58);
or U209 (N_209,In_222,In_452);
nand U210 (N_210,N_57,In_98);
nor U211 (N_211,In_426,N_7);
xnor U212 (N_212,In_235,N_84);
xor U213 (N_213,N_113,N_122);
xnor U214 (N_214,N_127,N_46);
xor U215 (N_215,In_366,In_367);
and U216 (N_216,In_155,In_167);
nand U217 (N_217,In_11,In_106);
nand U218 (N_218,In_431,In_166);
nor U219 (N_219,In_40,In_476);
nor U220 (N_220,N_125,N_22);
and U221 (N_221,In_248,N_106);
and U222 (N_222,N_52,In_76);
nor U223 (N_223,N_88,In_437);
nor U224 (N_224,In_173,N_11);
or U225 (N_225,N_224,In_24);
nand U226 (N_226,N_152,N_15);
or U227 (N_227,N_176,N_167);
or U228 (N_228,N_67,N_221);
and U229 (N_229,In_135,N_142);
nand U230 (N_230,In_269,In_26);
or U231 (N_231,N_206,N_180);
or U232 (N_232,N_145,N_150);
nand U233 (N_233,N_194,N_187);
and U234 (N_234,N_74,N_97);
or U235 (N_235,In_217,N_89);
nor U236 (N_236,In_225,N_220);
or U237 (N_237,In_193,N_65);
nand U238 (N_238,N_42,N_66);
and U239 (N_239,N_14,In_195);
nand U240 (N_240,N_35,In_116);
or U241 (N_241,In_140,In_446);
and U242 (N_242,N_98,N_163);
nor U243 (N_243,In_185,In_422);
or U244 (N_244,In_408,In_450);
or U245 (N_245,In_260,In_213);
nand U246 (N_246,N_169,In_416);
nor U247 (N_247,N_95,N_189);
nand U248 (N_248,N_129,N_208);
nand U249 (N_249,N_80,In_321);
nor U250 (N_250,N_193,N_139);
nor U251 (N_251,N_200,N_130);
nand U252 (N_252,In_207,N_201);
and U253 (N_253,In_330,N_170);
nor U254 (N_254,N_218,N_172);
and U255 (N_255,N_151,N_204);
nor U256 (N_256,In_375,N_174);
xnor U257 (N_257,In_453,N_131);
nand U258 (N_258,In_137,N_183);
and U259 (N_259,In_209,N_112);
or U260 (N_260,In_308,In_303);
xnor U261 (N_261,In_451,In_231);
or U262 (N_262,In_433,In_369);
nand U263 (N_263,In_27,In_53);
or U264 (N_264,N_203,In_50);
nor U265 (N_265,N_86,N_219);
nand U266 (N_266,In_138,In_103);
nand U267 (N_267,In_99,N_23);
and U268 (N_268,N_164,In_296);
and U269 (N_269,N_24,N_178);
or U270 (N_270,In_33,In_458);
and U271 (N_271,In_132,N_184);
xnor U272 (N_272,N_188,In_276);
nand U273 (N_273,In_171,In_467);
nand U274 (N_274,In_312,N_83);
or U275 (N_275,In_210,In_460);
or U276 (N_276,In_49,N_117);
and U277 (N_277,In_115,N_110);
nand U278 (N_278,In_289,N_39);
or U279 (N_279,In_91,N_68);
nand U280 (N_280,N_119,N_157);
or U281 (N_281,In_148,In_309);
and U282 (N_282,N_198,N_107);
xnor U283 (N_283,In_335,N_73);
nor U284 (N_284,In_8,In_199);
xnor U285 (N_285,In_2,N_134);
or U286 (N_286,In_175,N_213);
xnor U287 (N_287,In_86,N_62);
nand U288 (N_288,In_229,In_145);
nor U289 (N_289,In_181,In_379);
xor U290 (N_290,N_182,In_62);
xnor U291 (N_291,N_33,N_196);
xnor U292 (N_292,In_252,In_15);
nor U293 (N_293,N_34,N_179);
nand U294 (N_294,N_13,N_171);
xor U295 (N_295,N_212,In_430);
xnor U296 (N_296,N_28,In_107);
nand U297 (N_297,In_270,N_100);
xor U298 (N_298,N_195,N_132);
and U299 (N_299,In_464,In_302);
or U300 (N_300,N_59,N_78);
nand U301 (N_301,N_283,N_228);
nor U302 (N_302,In_159,In_297);
or U303 (N_303,In_249,N_177);
xnor U304 (N_304,N_234,In_44);
and U305 (N_305,N_226,In_448);
or U306 (N_306,In_442,N_181);
and U307 (N_307,N_215,N_216);
xor U308 (N_308,N_254,In_313);
nor U309 (N_309,N_287,In_469);
nand U310 (N_310,N_199,N_173);
xor U311 (N_311,In_261,N_252);
and U312 (N_312,In_490,N_270);
xor U313 (N_313,N_120,N_133);
and U314 (N_314,N_293,N_144);
and U315 (N_315,In_102,N_76);
nand U316 (N_316,N_79,In_415);
xor U317 (N_317,In_493,N_295);
nand U318 (N_318,N_262,N_241);
nand U319 (N_319,N_75,N_246);
nand U320 (N_320,N_261,N_249);
and U321 (N_321,In_176,N_265);
and U322 (N_322,In_315,In_129);
xor U323 (N_323,In_19,N_258);
nand U324 (N_324,N_251,N_168);
nand U325 (N_325,N_291,N_211);
xnor U326 (N_326,In_492,In_428);
or U327 (N_327,N_286,In_198);
and U328 (N_328,N_255,N_96);
nor U329 (N_329,N_90,N_263);
nor U330 (N_330,N_230,N_297);
xor U331 (N_331,N_207,N_209);
and U332 (N_332,In_85,In_435);
or U333 (N_333,N_118,N_244);
or U334 (N_334,In_97,In_343);
or U335 (N_335,In_291,N_243);
or U336 (N_336,N_253,N_257);
or U337 (N_337,N_225,N_229);
nor U338 (N_338,N_101,N_274);
or U339 (N_339,In_368,N_205);
nand U340 (N_340,In_482,In_304);
nor U341 (N_341,In_253,In_479);
and U342 (N_342,N_269,N_288);
or U343 (N_343,N_140,N_240);
nand U344 (N_344,N_69,N_290);
xor U345 (N_345,N_239,In_497);
nor U346 (N_346,In_211,In_134);
or U347 (N_347,N_217,N_165);
or U348 (N_348,In_182,N_202);
xnor U349 (N_349,N_278,In_113);
nor U350 (N_350,In_190,N_299);
and U351 (N_351,In_344,N_159);
and U352 (N_352,In_64,N_191);
or U353 (N_353,N_162,N_158);
or U354 (N_354,N_277,N_99);
and U355 (N_355,N_285,N_296);
nor U356 (N_356,N_289,N_227);
or U357 (N_357,N_248,In_274);
xor U358 (N_358,N_236,N_235);
or U359 (N_359,N_280,N_121);
nor U360 (N_360,In_194,In_324);
nor U361 (N_361,In_372,N_276);
or U362 (N_362,N_292,In_69);
and U363 (N_363,N_214,N_282);
nand U364 (N_364,N_238,N_271);
nor U365 (N_365,N_190,N_294);
or U366 (N_366,N_232,N_242);
nor U367 (N_367,N_166,N_192);
or U368 (N_368,N_30,N_60);
and U369 (N_369,In_333,N_135);
and U370 (N_370,In_25,N_32);
nand U371 (N_371,N_284,N_38);
nand U372 (N_372,N_231,N_103);
and U373 (N_373,In_66,N_175);
or U374 (N_374,N_250,N_155);
or U375 (N_375,N_361,In_256);
xor U376 (N_376,N_124,N_368);
nor U377 (N_377,N_185,N_360);
nor U378 (N_378,N_354,N_332);
nor U379 (N_379,N_223,N_322);
nand U380 (N_380,N_267,N_245);
or U381 (N_381,N_320,N_313);
or U382 (N_382,N_344,In_221);
or U383 (N_383,N_339,N_348);
xor U384 (N_384,N_323,N_334);
nand U385 (N_385,N_247,N_77);
nor U386 (N_386,N_268,N_342);
or U387 (N_387,N_161,N_340);
xnor U388 (N_388,N_303,N_233);
nor U389 (N_389,N_305,N_331);
or U390 (N_390,N_364,N_371);
or U391 (N_391,N_259,N_325);
or U392 (N_392,N_186,N_353);
nor U393 (N_393,In_22,N_92);
xnor U394 (N_394,N_315,N_275);
nor U395 (N_395,N_314,N_365);
nand U396 (N_396,N_260,N_279);
and U397 (N_397,N_336,N_343);
nand U398 (N_398,N_237,N_256);
or U399 (N_399,N_326,N_366);
or U400 (N_400,N_355,In_267);
nand U401 (N_401,N_337,N_72);
nor U402 (N_402,N_373,N_272);
nand U403 (N_403,N_306,N_304);
xor U404 (N_404,N_222,N_311);
xnor U405 (N_405,N_374,N_266);
nand U406 (N_406,N_358,N_281);
nor U407 (N_407,N_367,N_329);
and U408 (N_408,N_298,N_317);
and U409 (N_409,N_362,N_47);
nor U410 (N_410,N_328,In_471);
nor U411 (N_411,N_210,N_357);
nor U412 (N_412,N_300,N_338);
and U413 (N_413,N_345,N_264);
or U414 (N_414,N_308,N_93);
nand U415 (N_415,In_328,N_302);
nor U416 (N_416,N_319,N_154);
and U417 (N_417,N_301,In_142);
nor U418 (N_418,N_138,N_108);
nor U419 (N_419,N_310,N_318);
nor U420 (N_420,N_349,N_307);
nand U421 (N_421,N_346,In_55);
nor U422 (N_422,N_327,N_324);
and U423 (N_423,N_273,N_156);
nand U424 (N_424,N_321,N_370);
xnor U425 (N_425,N_347,N_350);
xnor U426 (N_426,In_149,N_359);
or U427 (N_427,N_351,In_429);
and U428 (N_428,N_197,N_330);
or U429 (N_429,N_153,N_309);
nand U430 (N_430,N_363,N_352);
nor U431 (N_431,N_316,In_342);
nand U432 (N_432,N_312,N_372);
xnor U433 (N_433,N_111,N_335);
or U434 (N_434,N_341,N_160);
nand U435 (N_435,N_369,N_356);
nand U436 (N_436,N_82,N_333);
or U437 (N_437,N_4,N_330);
xnor U438 (N_438,N_185,N_348);
and U439 (N_439,N_331,N_335);
xnor U440 (N_440,N_108,N_306);
and U441 (N_441,N_264,N_310);
nor U442 (N_442,N_359,N_368);
nand U443 (N_443,In_22,N_356);
or U444 (N_444,N_72,N_160);
nor U445 (N_445,N_124,N_307);
nor U446 (N_446,N_326,N_92);
nand U447 (N_447,N_47,N_349);
nor U448 (N_448,In_429,N_197);
xnor U449 (N_449,N_358,N_360);
or U450 (N_450,N_423,N_432);
and U451 (N_451,N_375,N_411);
nand U452 (N_452,N_448,N_417);
nor U453 (N_453,N_422,N_376);
nor U454 (N_454,N_379,N_391);
nor U455 (N_455,N_389,N_394);
nor U456 (N_456,N_441,N_418);
nand U457 (N_457,N_434,N_415);
and U458 (N_458,N_414,N_438);
nand U459 (N_459,N_384,N_429);
or U460 (N_460,N_408,N_405);
nand U461 (N_461,N_407,N_388);
nand U462 (N_462,N_380,N_400);
xor U463 (N_463,N_419,N_398);
and U464 (N_464,N_399,N_444);
xnor U465 (N_465,N_377,N_410);
nor U466 (N_466,N_436,N_383);
nand U467 (N_467,N_381,N_403);
or U468 (N_468,N_386,N_406);
and U469 (N_469,N_433,N_428);
xnor U470 (N_470,N_401,N_420);
and U471 (N_471,N_443,N_382);
or U472 (N_472,N_392,N_413);
nand U473 (N_473,N_435,N_446);
or U474 (N_474,N_430,N_449);
and U475 (N_475,N_445,N_447);
or U476 (N_476,N_409,N_378);
and U477 (N_477,N_390,N_385);
xor U478 (N_478,N_425,N_421);
and U479 (N_479,N_440,N_442);
nand U480 (N_480,N_437,N_439);
xnor U481 (N_481,N_427,N_431);
and U482 (N_482,N_395,N_412);
and U483 (N_483,N_387,N_424);
and U484 (N_484,N_396,N_393);
and U485 (N_485,N_426,N_402);
nand U486 (N_486,N_416,N_404);
nor U487 (N_487,N_397,N_430);
nor U488 (N_488,N_413,N_438);
nand U489 (N_489,N_413,N_436);
nor U490 (N_490,N_402,N_390);
and U491 (N_491,N_442,N_419);
nand U492 (N_492,N_404,N_424);
nand U493 (N_493,N_431,N_429);
or U494 (N_494,N_399,N_442);
nand U495 (N_495,N_398,N_443);
or U496 (N_496,N_431,N_449);
and U497 (N_497,N_436,N_405);
xnor U498 (N_498,N_428,N_441);
nor U499 (N_499,N_413,N_423);
or U500 (N_500,N_447,N_434);
and U501 (N_501,N_403,N_408);
xor U502 (N_502,N_428,N_415);
nand U503 (N_503,N_420,N_376);
and U504 (N_504,N_405,N_428);
xnor U505 (N_505,N_408,N_437);
nand U506 (N_506,N_414,N_382);
nand U507 (N_507,N_388,N_441);
nor U508 (N_508,N_426,N_444);
xor U509 (N_509,N_433,N_440);
xor U510 (N_510,N_424,N_446);
or U511 (N_511,N_388,N_418);
and U512 (N_512,N_384,N_427);
xnor U513 (N_513,N_398,N_437);
nor U514 (N_514,N_412,N_376);
nand U515 (N_515,N_437,N_384);
or U516 (N_516,N_439,N_435);
nor U517 (N_517,N_387,N_437);
xnor U518 (N_518,N_410,N_446);
xor U519 (N_519,N_381,N_447);
xnor U520 (N_520,N_405,N_441);
or U521 (N_521,N_444,N_436);
nand U522 (N_522,N_388,N_392);
nand U523 (N_523,N_394,N_401);
xnor U524 (N_524,N_414,N_397);
nor U525 (N_525,N_501,N_465);
or U526 (N_526,N_473,N_504);
nor U527 (N_527,N_478,N_479);
and U528 (N_528,N_467,N_459);
and U529 (N_529,N_469,N_472);
nand U530 (N_530,N_455,N_490);
or U531 (N_531,N_476,N_489);
nor U532 (N_532,N_494,N_520);
or U533 (N_533,N_497,N_477);
nor U534 (N_534,N_456,N_492);
or U535 (N_535,N_452,N_460);
xor U536 (N_536,N_499,N_485);
and U537 (N_537,N_481,N_518);
and U538 (N_538,N_510,N_521);
and U539 (N_539,N_487,N_524);
or U540 (N_540,N_515,N_451);
nand U541 (N_541,N_500,N_522);
and U542 (N_542,N_471,N_511);
nor U543 (N_543,N_450,N_486);
and U544 (N_544,N_505,N_506);
and U545 (N_545,N_475,N_502);
xnor U546 (N_546,N_466,N_516);
nor U547 (N_547,N_474,N_458);
xnor U548 (N_548,N_517,N_493);
nor U549 (N_549,N_464,N_488);
and U550 (N_550,N_496,N_509);
and U551 (N_551,N_503,N_514);
and U552 (N_552,N_454,N_480);
nand U553 (N_553,N_513,N_461);
or U554 (N_554,N_484,N_482);
nor U555 (N_555,N_507,N_495);
nor U556 (N_556,N_491,N_462);
nand U557 (N_557,N_512,N_468);
xor U558 (N_558,N_508,N_453);
xnor U559 (N_559,N_519,N_470);
nand U560 (N_560,N_523,N_498);
and U561 (N_561,N_457,N_463);
nor U562 (N_562,N_483,N_512);
nor U563 (N_563,N_453,N_515);
nand U564 (N_564,N_516,N_511);
and U565 (N_565,N_504,N_503);
nor U566 (N_566,N_500,N_495);
xnor U567 (N_567,N_490,N_520);
nand U568 (N_568,N_492,N_453);
nor U569 (N_569,N_506,N_520);
and U570 (N_570,N_469,N_455);
or U571 (N_571,N_483,N_521);
xnor U572 (N_572,N_480,N_488);
nand U573 (N_573,N_506,N_490);
nor U574 (N_574,N_484,N_508);
or U575 (N_575,N_476,N_513);
or U576 (N_576,N_507,N_461);
and U577 (N_577,N_507,N_484);
and U578 (N_578,N_517,N_510);
or U579 (N_579,N_514,N_473);
xor U580 (N_580,N_488,N_504);
and U581 (N_581,N_523,N_524);
nand U582 (N_582,N_465,N_450);
and U583 (N_583,N_454,N_516);
or U584 (N_584,N_453,N_460);
or U585 (N_585,N_456,N_510);
xor U586 (N_586,N_495,N_486);
xnor U587 (N_587,N_501,N_474);
or U588 (N_588,N_459,N_454);
or U589 (N_589,N_524,N_522);
nand U590 (N_590,N_466,N_508);
xor U591 (N_591,N_505,N_516);
and U592 (N_592,N_497,N_509);
nand U593 (N_593,N_520,N_524);
or U594 (N_594,N_471,N_502);
or U595 (N_595,N_490,N_470);
and U596 (N_596,N_524,N_518);
nor U597 (N_597,N_519,N_459);
xor U598 (N_598,N_491,N_472);
or U599 (N_599,N_513,N_517);
xnor U600 (N_600,N_574,N_589);
or U601 (N_601,N_546,N_588);
nor U602 (N_602,N_598,N_558);
nor U603 (N_603,N_567,N_544);
nor U604 (N_604,N_529,N_580);
xor U605 (N_605,N_592,N_555);
nor U606 (N_606,N_547,N_542);
nand U607 (N_607,N_571,N_532);
or U608 (N_608,N_590,N_579);
nand U609 (N_609,N_569,N_565);
or U610 (N_610,N_554,N_534);
nand U611 (N_611,N_556,N_573);
and U612 (N_612,N_575,N_564);
xnor U613 (N_613,N_597,N_583);
nand U614 (N_614,N_533,N_538);
nand U615 (N_615,N_543,N_537);
or U616 (N_616,N_528,N_562);
and U617 (N_617,N_587,N_550);
xnor U618 (N_618,N_527,N_561);
nor U619 (N_619,N_595,N_535);
nor U620 (N_620,N_582,N_560);
nand U621 (N_621,N_539,N_576);
or U622 (N_622,N_566,N_563);
xor U623 (N_623,N_596,N_545);
xor U624 (N_624,N_530,N_572);
xnor U625 (N_625,N_599,N_526);
nand U626 (N_626,N_581,N_578);
nor U627 (N_627,N_594,N_568);
xnor U628 (N_628,N_549,N_553);
nor U629 (N_629,N_577,N_551);
and U630 (N_630,N_584,N_552);
or U631 (N_631,N_536,N_586);
nand U632 (N_632,N_541,N_591);
nor U633 (N_633,N_557,N_593);
xor U634 (N_634,N_570,N_559);
xnor U635 (N_635,N_540,N_531);
nor U636 (N_636,N_585,N_548);
xnor U637 (N_637,N_525,N_570);
and U638 (N_638,N_563,N_540);
and U639 (N_639,N_588,N_593);
nand U640 (N_640,N_555,N_565);
xnor U641 (N_641,N_588,N_556);
or U642 (N_642,N_540,N_565);
nand U643 (N_643,N_567,N_545);
or U644 (N_644,N_588,N_589);
and U645 (N_645,N_565,N_596);
nor U646 (N_646,N_573,N_590);
nor U647 (N_647,N_556,N_542);
nand U648 (N_648,N_599,N_566);
nand U649 (N_649,N_573,N_593);
or U650 (N_650,N_536,N_543);
nor U651 (N_651,N_529,N_587);
nand U652 (N_652,N_552,N_556);
and U653 (N_653,N_569,N_529);
or U654 (N_654,N_568,N_538);
nor U655 (N_655,N_596,N_564);
or U656 (N_656,N_555,N_545);
nor U657 (N_657,N_574,N_538);
or U658 (N_658,N_548,N_574);
or U659 (N_659,N_563,N_594);
nand U660 (N_660,N_536,N_546);
xnor U661 (N_661,N_542,N_574);
nor U662 (N_662,N_547,N_533);
xnor U663 (N_663,N_558,N_586);
and U664 (N_664,N_588,N_532);
xnor U665 (N_665,N_525,N_544);
and U666 (N_666,N_579,N_534);
or U667 (N_667,N_557,N_589);
or U668 (N_668,N_570,N_557);
nor U669 (N_669,N_538,N_565);
xor U670 (N_670,N_543,N_587);
nand U671 (N_671,N_576,N_595);
and U672 (N_672,N_544,N_574);
nand U673 (N_673,N_533,N_544);
nand U674 (N_674,N_589,N_556);
nand U675 (N_675,N_628,N_631);
nand U676 (N_676,N_633,N_617);
or U677 (N_677,N_635,N_671);
nand U678 (N_678,N_603,N_613);
nor U679 (N_679,N_621,N_615);
nand U680 (N_680,N_604,N_611);
or U681 (N_681,N_602,N_636);
and U682 (N_682,N_649,N_622);
nand U683 (N_683,N_663,N_645);
and U684 (N_684,N_659,N_664);
or U685 (N_685,N_643,N_638);
and U686 (N_686,N_670,N_640);
or U687 (N_687,N_655,N_653);
or U688 (N_688,N_648,N_629);
nor U689 (N_689,N_656,N_652);
nor U690 (N_690,N_637,N_641);
nor U691 (N_691,N_660,N_662);
nand U692 (N_692,N_639,N_610);
or U693 (N_693,N_618,N_608);
and U694 (N_694,N_672,N_666);
or U695 (N_695,N_650,N_651);
or U696 (N_696,N_658,N_620);
nand U697 (N_697,N_627,N_612);
and U698 (N_698,N_646,N_634);
and U699 (N_699,N_619,N_625);
or U700 (N_700,N_605,N_674);
or U701 (N_701,N_647,N_632);
and U702 (N_702,N_606,N_673);
nand U703 (N_703,N_623,N_642);
nand U704 (N_704,N_614,N_661);
or U705 (N_705,N_609,N_626);
nand U706 (N_706,N_668,N_657);
and U707 (N_707,N_644,N_624);
and U708 (N_708,N_607,N_654);
and U709 (N_709,N_669,N_601);
or U710 (N_710,N_616,N_630);
nor U711 (N_711,N_667,N_600);
or U712 (N_712,N_665,N_667);
or U713 (N_713,N_627,N_632);
or U714 (N_714,N_660,N_618);
and U715 (N_715,N_648,N_646);
and U716 (N_716,N_614,N_640);
xor U717 (N_717,N_655,N_623);
nor U718 (N_718,N_633,N_673);
nor U719 (N_719,N_665,N_634);
nor U720 (N_720,N_619,N_616);
xnor U721 (N_721,N_636,N_653);
xnor U722 (N_722,N_648,N_633);
and U723 (N_723,N_670,N_608);
nor U724 (N_724,N_603,N_627);
nor U725 (N_725,N_634,N_610);
xnor U726 (N_726,N_643,N_627);
xor U727 (N_727,N_625,N_615);
nand U728 (N_728,N_650,N_600);
nor U729 (N_729,N_628,N_615);
xnor U730 (N_730,N_667,N_639);
or U731 (N_731,N_624,N_632);
and U732 (N_732,N_610,N_624);
xnor U733 (N_733,N_607,N_622);
and U734 (N_734,N_617,N_610);
nor U735 (N_735,N_618,N_610);
and U736 (N_736,N_638,N_639);
and U737 (N_737,N_663,N_670);
xnor U738 (N_738,N_664,N_645);
and U739 (N_739,N_656,N_637);
and U740 (N_740,N_656,N_632);
nor U741 (N_741,N_619,N_614);
nand U742 (N_742,N_630,N_627);
nor U743 (N_743,N_673,N_646);
xor U744 (N_744,N_610,N_623);
or U745 (N_745,N_646,N_602);
and U746 (N_746,N_605,N_658);
nand U747 (N_747,N_600,N_630);
xor U748 (N_748,N_663,N_659);
or U749 (N_749,N_637,N_666);
and U750 (N_750,N_714,N_745);
nor U751 (N_751,N_726,N_704);
nand U752 (N_752,N_741,N_694);
nor U753 (N_753,N_748,N_676);
and U754 (N_754,N_678,N_702);
nor U755 (N_755,N_701,N_730);
xnor U756 (N_756,N_698,N_736);
or U757 (N_757,N_744,N_699);
or U758 (N_758,N_682,N_731);
nor U759 (N_759,N_707,N_717);
or U760 (N_760,N_724,N_738);
and U761 (N_761,N_705,N_715);
or U762 (N_762,N_684,N_719);
xnor U763 (N_763,N_742,N_727);
xnor U764 (N_764,N_746,N_700);
and U765 (N_765,N_675,N_747);
xnor U766 (N_766,N_693,N_743);
or U767 (N_767,N_690,N_729);
nand U768 (N_768,N_734,N_691);
nor U769 (N_769,N_688,N_732);
nand U770 (N_770,N_733,N_728);
nor U771 (N_771,N_680,N_739);
nand U772 (N_772,N_681,N_723);
and U773 (N_773,N_735,N_713);
xor U774 (N_774,N_711,N_708);
xor U775 (N_775,N_696,N_712);
nand U776 (N_776,N_677,N_697);
xnor U777 (N_777,N_689,N_703);
and U778 (N_778,N_740,N_716);
or U779 (N_779,N_706,N_687);
or U780 (N_780,N_695,N_692);
xnor U781 (N_781,N_679,N_749);
or U782 (N_782,N_721,N_720);
nor U783 (N_783,N_722,N_709);
or U784 (N_784,N_686,N_718);
or U785 (N_785,N_685,N_737);
nand U786 (N_786,N_683,N_725);
xor U787 (N_787,N_710,N_696);
xnor U788 (N_788,N_741,N_688);
nand U789 (N_789,N_688,N_681);
nor U790 (N_790,N_681,N_735);
or U791 (N_791,N_740,N_739);
and U792 (N_792,N_723,N_747);
and U793 (N_793,N_679,N_736);
nor U794 (N_794,N_721,N_686);
or U795 (N_795,N_735,N_739);
xor U796 (N_796,N_705,N_676);
or U797 (N_797,N_724,N_740);
or U798 (N_798,N_683,N_744);
nor U799 (N_799,N_709,N_725);
nor U800 (N_800,N_738,N_708);
nor U801 (N_801,N_693,N_696);
and U802 (N_802,N_708,N_687);
xor U803 (N_803,N_747,N_741);
xor U804 (N_804,N_722,N_746);
and U805 (N_805,N_735,N_689);
nor U806 (N_806,N_732,N_705);
and U807 (N_807,N_696,N_682);
nand U808 (N_808,N_694,N_724);
xor U809 (N_809,N_686,N_711);
xnor U810 (N_810,N_725,N_690);
nor U811 (N_811,N_683,N_700);
and U812 (N_812,N_703,N_748);
or U813 (N_813,N_733,N_749);
nor U814 (N_814,N_722,N_700);
nand U815 (N_815,N_739,N_743);
nor U816 (N_816,N_715,N_678);
xor U817 (N_817,N_711,N_739);
nand U818 (N_818,N_745,N_715);
nor U819 (N_819,N_721,N_717);
nand U820 (N_820,N_731,N_701);
nor U821 (N_821,N_737,N_689);
and U822 (N_822,N_681,N_714);
nor U823 (N_823,N_689,N_718);
nor U824 (N_824,N_731,N_746);
or U825 (N_825,N_752,N_823);
nand U826 (N_826,N_761,N_816);
or U827 (N_827,N_798,N_810);
or U828 (N_828,N_780,N_786);
xnor U829 (N_829,N_754,N_772);
and U830 (N_830,N_756,N_760);
xnor U831 (N_831,N_811,N_753);
nor U832 (N_832,N_764,N_778);
or U833 (N_833,N_769,N_815);
nor U834 (N_834,N_757,N_819);
nand U835 (N_835,N_808,N_812);
nand U836 (N_836,N_765,N_791);
and U837 (N_837,N_785,N_751);
nand U838 (N_838,N_795,N_794);
nand U839 (N_839,N_777,N_771);
and U840 (N_840,N_758,N_818);
nor U841 (N_841,N_792,N_762);
or U842 (N_842,N_759,N_804);
nand U843 (N_843,N_805,N_789);
and U844 (N_844,N_793,N_784);
nor U845 (N_845,N_774,N_807);
or U846 (N_846,N_755,N_814);
xor U847 (N_847,N_787,N_783);
xor U848 (N_848,N_813,N_782);
nor U849 (N_849,N_768,N_800);
nor U850 (N_850,N_779,N_797);
nor U851 (N_851,N_770,N_781);
xnor U852 (N_852,N_790,N_817);
or U853 (N_853,N_801,N_803);
nor U854 (N_854,N_799,N_763);
and U855 (N_855,N_773,N_750);
nor U856 (N_856,N_802,N_806);
and U857 (N_857,N_766,N_776);
xor U858 (N_858,N_796,N_824);
or U859 (N_859,N_820,N_775);
nor U860 (N_860,N_788,N_767);
or U861 (N_861,N_821,N_809);
or U862 (N_862,N_822,N_807);
or U863 (N_863,N_807,N_768);
nor U864 (N_864,N_768,N_761);
or U865 (N_865,N_812,N_761);
nor U866 (N_866,N_791,N_760);
nand U867 (N_867,N_796,N_762);
and U868 (N_868,N_767,N_816);
nor U869 (N_869,N_823,N_790);
and U870 (N_870,N_784,N_758);
nor U871 (N_871,N_799,N_784);
nand U872 (N_872,N_761,N_822);
xnor U873 (N_873,N_810,N_780);
and U874 (N_874,N_809,N_819);
and U875 (N_875,N_768,N_776);
nand U876 (N_876,N_778,N_777);
nand U877 (N_877,N_819,N_769);
or U878 (N_878,N_762,N_822);
and U879 (N_879,N_811,N_823);
or U880 (N_880,N_822,N_784);
nor U881 (N_881,N_777,N_776);
or U882 (N_882,N_817,N_770);
and U883 (N_883,N_823,N_809);
nand U884 (N_884,N_793,N_810);
xor U885 (N_885,N_818,N_752);
xnor U886 (N_886,N_750,N_814);
nand U887 (N_887,N_755,N_815);
nand U888 (N_888,N_803,N_753);
nand U889 (N_889,N_808,N_798);
xor U890 (N_890,N_750,N_824);
nor U891 (N_891,N_760,N_770);
nor U892 (N_892,N_751,N_762);
nand U893 (N_893,N_791,N_754);
nand U894 (N_894,N_805,N_752);
and U895 (N_895,N_774,N_758);
nand U896 (N_896,N_764,N_763);
and U897 (N_897,N_824,N_812);
and U898 (N_898,N_779,N_805);
or U899 (N_899,N_795,N_767);
xor U900 (N_900,N_831,N_859);
xor U901 (N_901,N_860,N_856);
nor U902 (N_902,N_846,N_864);
nor U903 (N_903,N_862,N_880);
or U904 (N_904,N_885,N_850);
and U905 (N_905,N_871,N_827);
nand U906 (N_906,N_865,N_845);
nand U907 (N_907,N_854,N_832);
xor U908 (N_908,N_866,N_887);
nand U909 (N_909,N_868,N_839);
nand U910 (N_910,N_840,N_881);
and U911 (N_911,N_836,N_828);
nand U912 (N_912,N_842,N_834);
nor U913 (N_913,N_889,N_884);
and U914 (N_914,N_863,N_851);
or U915 (N_915,N_882,N_844);
xnor U916 (N_916,N_876,N_892);
nor U917 (N_917,N_874,N_886);
and U918 (N_918,N_875,N_826);
or U919 (N_919,N_848,N_883);
xor U920 (N_920,N_837,N_847);
nor U921 (N_921,N_849,N_870);
and U922 (N_922,N_898,N_852);
or U923 (N_923,N_841,N_855);
or U924 (N_924,N_877,N_873);
xnor U925 (N_925,N_879,N_833);
nand U926 (N_926,N_830,N_894);
nor U927 (N_927,N_838,N_890);
or U928 (N_928,N_843,N_835);
nand U929 (N_929,N_888,N_895);
nor U930 (N_930,N_853,N_869);
nand U931 (N_931,N_893,N_861);
or U932 (N_932,N_825,N_897);
nor U933 (N_933,N_896,N_891);
nor U934 (N_934,N_829,N_872);
xnor U935 (N_935,N_899,N_857);
and U936 (N_936,N_858,N_878);
or U937 (N_937,N_867,N_850);
xor U938 (N_938,N_862,N_831);
xor U939 (N_939,N_838,N_866);
nor U940 (N_940,N_835,N_868);
or U941 (N_941,N_845,N_842);
nand U942 (N_942,N_854,N_899);
and U943 (N_943,N_868,N_883);
xnor U944 (N_944,N_872,N_827);
and U945 (N_945,N_863,N_892);
xnor U946 (N_946,N_853,N_894);
xor U947 (N_947,N_865,N_829);
nand U948 (N_948,N_847,N_865);
xnor U949 (N_949,N_879,N_854);
xor U950 (N_950,N_844,N_898);
or U951 (N_951,N_878,N_873);
or U952 (N_952,N_844,N_854);
nand U953 (N_953,N_888,N_889);
nand U954 (N_954,N_874,N_849);
nor U955 (N_955,N_892,N_897);
xor U956 (N_956,N_860,N_871);
xor U957 (N_957,N_853,N_848);
xor U958 (N_958,N_852,N_864);
and U959 (N_959,N_873,N_832);
or U960 (N_960,N_888,N_828);
and U961 (N_961,N_878,N_863);
and U962 (N_962,N_849,N_885);
nor U963 (N_963,N_835,N_859);
xnor U964 (N_964,N_868,N_825);
nand U965 (N_965,N_830,N_834);
or U966 (N_966,N_844,N_885);
xnor U967 (N_967,N_871,N_849);
nor U968 (N_968,N_871,N_837);
and U969 (N_969,N_884,N_866);
nor U970 (N_970,N_846,N_892);
and U971 (N_971,N_858,N_837);
nor U972 (N_972,N_840,N_830);
or U973 (N_973,N_845,N_856);
or U974 (N_974,N_896,N_886);
and U975 (N_975,N_940,N_904);
nand U976 (N_976,N_936,N_944);
or U977 (N_977,N_954,N_952);
xor U978 (N_978,N_924,N_909);
or U979 (N_979,N_928,N_939);
xnor U980 (N_980,N_902,N_925);
nor U981 (N_981,N_960,N_955);
or U982 (N_982,N_912,N_974);
nor U983 (N_983,N_938,N_958);
nand U984 (N_984,N_935,N_949);
nand U985 (N_985,N_914,N_920);
or U986 (N_986,N_971,N_932);
or U987 (N_987,N_908,N_961);
nand U988 (N_988,N_968,N_933);
and U989 (N_989,N_919,N_930);
xnor U990 (N_990,N_934,N_959);
or U991 (N_991,N_946,N_913);
nor U992 (N_992,N_967,N_941);
and U993 (N_993,N_901,N_969);
nand U994 (N_994,N_964,N_910);
xnor U995 (N_995,N_905,N_947);
xnor U996 (N_996,N_927,N_911);
nand U997 (N_997,N_942,N_972);
and U998 (N_998,N_966,N_926);
nor U999 (N_999,N_907,N_970);
nor U1000 (N_1000,N_903,N_943);
nor U1001 (N_1001,N_963,N_937);
or U1002 (N_1002,N_921,N_957);
nor U1003 (N_1003,N_915,N_973);
xor U1004 (N_1004,N_906,N_948);
nand U1005 (N_1005,N_929,N_931);
nand U1006 (N_1006,N_956,N_953);
or U1007 (N_1007,N_918,N_950);
and U1008 (N_1008,N_965,N_916);
and U1009 (N_1009,N_917,N_945);
or U1010 (N_1010,N_962,N_951);
and U1011 (N_1011,N_923,N_922);
xnor U1012 (N_1012,N_900,N_906);
nand U1013 (N_1013,N_948,N_919);
nand U1014 (N_1014,N_929,N_913);
nand U1015 (N_1015,N_970,N_949);
and U1016 (N_1016,N_921,N_944);
or U1017 (N_1017,N_936,N_940);
or U1018 (N_1018,N_927,N_925);
or U1019 (N_1019,N_912,N_903);
and U1020 (N_1020,N_918,N_946);
and U1021 (N_1021,N_904,N_970);
nor U1022 (N_1022,N_936,N_901);
nor U1023 (N_1023,N_926,N_913);
xnor U1024 (N_1024,N_972,N_905);
xor U1025 (N_1025,N_945,N_919);
nor U1026 (N_1026,N_920,N_946);
and U1027 (N_1027,N_952,N_942);
or U1028 (N_1028,N_954,N_961);
nand U1029 (N_1029,N_904,N_939);
or U1030 (N_1030,N_970,N_919);
and U1031 (N_1031,N_914,N_919);
and U1032 (N_1032,N_917,N_924);
or U1033 (N_1033,N_912,N_918);
nor U1034 (N_1034,N_914,N_965);
xor U1035 (N_1035,N_920,N_950);
xnor U1036 (N_1036,N_910,N_959);
or U1037 (N_1037,N_960,N_931);
and U1038 (N_1038,N_914,N_946);
nor U1039 (N_1039,N_950,N_906);
and U1040 (N_1040,N_905,N_955);
nand U1041 (N_1041,N_902,N_935);
and U1042 (N_1042,N_908,N_957);
xor U1043 (N_1043,N_948,N_938);
xor U1044 (N_1044,N_957,N_922);
nor U1045 (N_1045,N_970,N_924);
or U1046 (N_1046,N_965,N_935);
xor U1047 (N_1047,N_914,N_959);
xor U1048 (N_1048,N_930,N_928);
xor U1049 (N_1049,N_947,N_903);
xor U1050 (N_1050,N_988,N_1000);
and U1051 (N_1051,N_979,N_980);
or U1052 (N_1052,N_1032,N_996);
and U1053 (N_1053,N_1004,N_999);
nand U1054 (N_1054,N_1030,N_1025);
nand U1055 (N_1055,N_1046,N_1006);
or U1056 (N_1056,N_1017,N_1001);
and U1057 (N_1057,N_1041,N_1008);
nor U1058 (N_1058,N_1033,N_1034);
or U1059 (N_1059,N_994,N_1023);
xnor U1060 (N_1060,N_1021,N_1020);
or U1061 (N_1061,N_1040,N_1019);
nand U1062 (N_1062,N_1013,N_1045);
or U1063 (N_1063,N_981,N_1014);
nand U1064 (N_1064,N_1022,N_976);
xor U1065 (N_1065,N_1036,N_982);
nand U1066 (N_1066,N_975,N_989);
or U1067 (N_1067,N_1012,N_985);
xor U1068 (N_1068,N_986,N_995);
nand U1069 (N_1069,N_1044,N_997);
and U1070 (N_1070,N_987,N_1002);
or U1071 (N_1071,N_1016,N_1047);
xor U1072 (N_1072,N_1027,N_1035);
or U1073 (N_1073,N_1009,N_1018);
nor U1074 (N_1074,N_1039,N_1048);
or U1075 (N_1075,N_978,N_992);
and U1076 (N_1076,N_1003,N_990);
nor U1077 (N_1077,N_977,N_1043);
nor U1078 (N_1078,N_983,N_1031);
nand U1079 (N_1079,N_1026,N_984);
or U1080 (N_1080,N_1011,N_1015);
xnor U1081 (N_1081,N_1042,N_1038);
nor U1082 (N_1082,N_991,N_1005);
nor U1083 (N_1083,N_1049,N_993);
or U1084 (N_1084,N_1007,N_1028);
nand U1085 (N_1085,N_998,N_1024);
nand U1086 (N_1086,N_1037,N_1029);
or U1087 (N_1087,N_1010,N_982);
or U1088 (N_1088,N_1018,N_1017);
nor U1089 (N_1089,N_1022,N_986);
xor U1090 (N_1090,N_1027,N_986);
and U1091 (N_1091,N_988,N_1040);
nand U1092 (N_1092,N_996,N_999);
nand U1093 (N_1093,N_994,N_1021);
or U1094 (N_1094,N_1000,N_977);
and U1095 (N_1095,N_1037,N_1014);
or U1096 (N_1096,N_985,N_1045);
xor U1097 (N_1097,N_1049,N_987);
nor U1098 (N_1098,N_1041,N_987);
nor U1099 (N_1099,N_985,N_1039);
and U1100 (N_1100,N_1039,N_1047);
nor U1101 (N_1101,N_1022,N_1008);
or U1102 (N_1102,N_1007,N_1021);
and U1103 (N_1103,N_1005,N_1041);
and U1104 (N_1104,N_1010,N_1034);
xor U1105 (N_1105,N_1040,N_1035);
or U1106 (N_1106,N_1037,N_1024);
nand U1107 (N_1107,N_1021,N_1034);
xnor U1108 (N_1108,N_1023,N_1037);
nor U1109 (N_1109,N_1014,N_976);
or U1110 (N_1110,N_1004,N_1029);
and U1111 (N_1111,N_996,N_1020);
and U1112 (N_1112,N_994,N_1024);
and U1113 (N_1113,N_1038,N_1003);
or U1114 (N_1114,N_1026,N_1028);
and U1115 (N_1115,N_1002,N_1006);
nand U1116 (N_1116,N_1034,N_1042);
and U1117 (N_1117,N_1002,N_1043);
nand U1118 (N_1118,N_1049,N_1008);
and U1119 (N_1119,N_979,N_1005);
and U1120 (N_1120,N_997,N_1033);
xor U1121 (N_1121,N_980,N_1014);
and U1122 (N_1122,N_1027,N_981);
nor U1123 (N_1123,N_1021,N_980);
nor U1124 (N_1124,N_1029,N_977);
nor U1125 (N_1125,N_1057,N_1072);
or U1126 (N_1126,N_1061,N_1082);
nand U1127 (N_1127,N_1113,N_1077);
xor U1128 (N_1128,N_1109,N_1100);
nor U1129 (N_1129,N_1104,N_1078);
nor U1130 (N_1130,N_1101,N_1094);
nor U1131 (N_1131,N_1068,N_1116);
nand U1132 (N_1132,N_1105,N_1051);
xnor U1133 (N_1133,N_1050,N_1056);
nand U1134 (N_1134,N_1063,N_1093);
nor U1135 (N_1135,N_1071,N_1066);
and U1136 (N_1136,N_1076,N_1087);
and U1137 (N_1137,N_1070,N_1054);
xnor U1138 (N_1138,N_1086,N_1120);
or U1139 (N_1139,N_1106,N_1081);
or U1140 (N_1140,N_1119,N_1062);
or U1141 (N_1141,N_1080,N_1124);
or U1142 (N_1142,N_1103,N_1114);
or U1143 (N_1143,N_1099,N_1074);
or U1144 (N_1144,N_1073,N_1092);
xor U1145 (N_1145,N_1079,N_1075);
and U1146 (N_1146,N_1102,N_1055);
or U1147 (N_1147,N_1084,N_1052);
nor U1148 (N_1148,N_1065,N_1091);
or U1149 (N_1149,N_1095,N_1108);
xor U1150 (N_1150,N_1118,N_1107);
or U1151 (N_1151,N_1122,N_1089);
and U1152 (N_1152,N_1117,N_1085);
nor U1153 (N_1153,N_1097,N_1053);
nand U1154 (N_1154,N_1064,N_1115);
xor U1155 (N_1155,N_1083,N_1090);
xnor U1156 (N_1156,N_1067,N_1110);
xnor U1157 (N_1157,N_1058,N_1059);
nand U1158 (N_1158,N_1060,N_1098);
nor U1159 (N_1159,N_1111,N_1088);
nor U1160 (N_1160,N_1112,N_1096);
and U1161 (N_1161,N_1069,N_1121);
nand U1162 (N_1162,N_1123,N_1124);
nand U1163 (N_1163,N_1076,N_1068);
nand U1164 (N_1164,N_1112,N_1067);
nor U1165 (N_1165,N_1107,N_1089);
and U1166 (N_1166,N_1101,N_1061);
xnor U1167 (N_1167,N_1097,N_1066);
nor U1168 (N_1168,N_1124,N_1052);
nand U1169 (N_1169,N_1092,N_1117);
xnor U1170 (N_1170,N_1079,N_1122);
or U1171 (N_1171,N_1118,N_1055);
xnor U1172 (N_1172,N_1119,N_1061);
or U1173 (N_1173,N_1107,N_1117);
nand U1174 (N_1174,N_1095,N_1098);
xnor U1175 (N_1175,N_1070,N_1066);
or U1176 (N_1176,N_1050,N_1094);
and U1177 (N_1177,N_1123,N_1054);
or U1178 (N_1178,N_1060,N_1102);
nand U1179 (N_1179,N_1055,N_1076);
or U1180 (N_1180,N_1096,N_1078);
or U1181 (N_1181,N_1051,N_1100);
or U1182 (N_1182,N_1094,N_1086);
or U1183 (N_1183,N_1101,N_1096);
or U1184 (N_1184,N_1120,N_1116);
and U1185 (N_1185,N_1087,N_1080);
xor U1186 (N_1186,N_1110,N_1057);
xnor U1187 (N_1187,N_1113,N_1099);
or U1188 (N_1188,N_1109,N_1089);
or U1189 (N_1189,N_1079,N_1065);
or U1190 (N_1190,N_1056,N_1084);
xnor U1191 (N_1191,N_1113,N_1124);
xor U1192 (N_1192,N_1050,N_1075);
and U1193 (N_1193,N_1079,N_1082);
nor U1194 (N_1194,N_1084,N_1115);
xor U1195 (N_1195,N_1076,N_1102);
xor U1196 (N_1196,N_1113,N_1117);
nor U1197 (N_1197,N_1053,N_1087);
xnor U1198 (N_1198,N_1077,N_1105);
nand U1199 (N_1199,N_1101,N_1112);
or U1200 (N_1200,N_1184,N_1168);
nand U1201 (N_1201,N_1170,N_1127);
nor U1202 (N_1202,N_1189,N_1138);
and U1203 (N_1203,N_1157,N_1146);
nor U1204 (N_1204,N_1181,N_1193);
nand U1205 (N_1205,N_1178,N_1180);
and U1206 (N_1206,N_1143,N_1171);
nor U1207 (N_1207,N_1140,N_1152);
and U1208 (N_1208,N_1162,N_1155);
or U1209 (N_1209,N_1192,N_1172);
or U1210 (N_1210,N_1133,N_1132);
nor U1211 (N_1211,N_1175,N_1130);
nand U1212 (N_1212,N_1190,N_1198);
nor U1213 (N_1213,N_1156,N_1187);
xor U1214 (N_1214,N_1150,N_1185);
nand U1215 (N_1215,N_1176,N_1159);
nor U1216 (N_1216,N_1161,N_1167);
and U1217 (N_1217,N_1154,N_1136);
xor U1218 (N_1218,N_1194,N_1188);
and U1219 (N_1219,N_1158,N_1199);
nand U1220 (N_1220,N_1128,N_1129);
nor U1221 (N_1221,N_1174,N_1182);
nor U1222 (N_1222,N_1135,N_1179);
or U1223 (N_1223,N_1160,N_1186);
nand U1224 (N_1224,N_1142,N_1191);
xnor U1225 (N_1225,N_1149,N_1151);
xor U1226 (N_1226,N_1169,N_1153);
or U1227 (N_1227,N_1134,N_1163);
nand U1228 (N_1228,N_1144,N_1196);
xor U1229 (N_1229,N_1197,N_1137);
nor U1230 (N_1230,N_1139,N_1195);
nand U1231 (N_1231,N_1164,N_1148);
nor U1232 (N_1232,N_1126,N_1131);
nor U1233 (N_1233,N_1177,N_1166);
and U1234 (N_1234,N_1173,N_1125);
xor U1235 (N_1235,N_1141,N_1147);
xor U1236 (N_1236,N_1165,N_1183);
xor U1237 (N_1237,N_1145,N_1147);
nor U1238 (N_1238,N_1147,N_1197);
xor U1239 (N_1239,N_1161,N_1194);
nand U1240 (N_1240,N_1191,N_1129);
or U1241 (N_1241,N_1148,N_1170);
and U1242 (N_1242,N_1177,N_1174);
nand U1243 (N_1243,N_1173,N_1179);
xnor U1244 (N_1244,N_1163,N_1184);
or U1245 (N_1245,N_1146,N_1127);
nor U1246 (N_1246,N_1157,N_1125);
nor U1247 (N_1247,N_1133,N_1136);
nand U1248 (N_1248,N_1137,N_1176);
nor U1249 (N_1249,N_1181,N_1134);
nand U1250 (N_1250,N_1147,N_1174);
or U1251 (N_1251,N_1192,N_1181);
and U1252 (N_1252,N_1173,N_1160);
xnor U1253 (N_1253,N_1166,N_1139);
nand U1254 (N_1254,N_1187,N_1180);
nand U1255 (N_1255,N_1142,N_1141);
and U1256 (N_1256,N_1142,N_1196);
nor U1257 (N_1257,N_1197,N_1138);
nor U1258 (N_1258,N_1179,N_1168);
nor U1259 (N_1259,N_1167,N_1187);
or U1260 (N_1260,N_1176,N_1142);
and U1261 (N_1261,N_1173,N_1143);
nor U1262 (N_1262,N_1136,N_1191);
xor U1263 (N_1263,N_1142,N_1166);
and U1264 (N_1264,N_1136,N_1159);
nor U1265 (N_1265,N_1125,N_1131);
or U1266 (N_1266,N_1149,N_1135);
nor U1267 (N_1267,N_1142,N_1198);
or U1268 (N_1268,N_1184,N_1169);
nand U1269 (N_1269,N_1167,N_1180);
and U1270 (N_1270,N_1180,N_1134);
nor U1271 (N_1271,N_1168,N_1152);
nand U1272 (N_1272,N_1196,N_1195);
nand U1273 (N_1273,N_1142,N_1133);
xor U1274 (N_1274,N_1193,N_1185);
nor U1275 (N_1275,N_1209,N_1226);
xor U1276 (N_1276,N_1253,N_1227);
or U1277 (N_1277,N_1238,N_1216);
or U1278 (N_1278,N_1260,N_1272);
or U1279 (N_1279,N_1265,N_1268);
and U1280 (N_1280,N_1207,N_1222);
nor U1281 (N_1281,N_1240,N_1232);
xor U1282 (N_1282,N_1267,N_1257);
nand U1283 (N_1283,N_1230,N_1245);
nor U1284 (N_1284,N_1270,N_1208);
nor U1285 (N_1285,N_1205,N_1224);
and U1286 (N_1286,N_1254,N_1243);
nor U1287 (N_1287,N_1255,N_1246);
xnor U1288 (N_1288,N_1252,N_1225);
and U1289 (N_1289,N_1237,N_1213);
nand U1290 (N_1290,N_1206,N_1259);
nand U1291 (N_1291,N_1269,N_1212);
or U1292 (N_1292,N_1266,N_1228);
xnor U1293 (N_1293,N_1248,N_1211);
nand U1294 (N_1294,N_1234,N_1210);
or U1295 (N_1295,N_1229,N_1263);
nand U1296 (N_1296,N_1236,N_1215);
nor U1297 (N_1297,N_1264,N_1221);
and U1298 (N_1298,N_1261,N_1256);
or U1299 (N_1299,N_1201,N_1247);
or U1300 (N_1300,N_1223,N_1271);
xnor U1301 (N_1301,N_1217,N_1258);
xnor U1302 (N_1302,N_1250,N_1249);
and U1303 (N_1303,N_1219,N_1203);
nor U1304 (N_1304,N_1220,N_1242);
xnor U1305 (N_1305,N_1241,N_1273);
nor U1306 (N_1306,N_1251,N_1262);
and U1307 (N_1307,N_1231,N_1239);
and U1308 (N_1308,N_1274,N_1235);
and U1309 (N_1309,N_1233,N_1200);
xnor U1310 (N_1310,N_1202,N_1204);
nand U1311 (N_1311,N_1214,N_1244);
nand U1312 (N_1312,N_1218,N_1243);
and U1313 (N_1313,N_1214,N_1232);
nor U1314 (N_1314,N_1256,N_1237);
nor U1315 (N_1315,N_1249,N_1241);
and U1316 (N_1316,N_1257,N_1224);
nand U1317 (N_1317,N_1250,N_1265);
and U1318 (N_1318,N_1246,N_1266);
and U1319 (N_1319,N_1232,N_1223);
or U1320 (N_1320,N_1202,N_1227);
xnor U1321 (N_1321,N_1238,N_1235);
xor U1322 (N_1322,N_1243,N_1256);
xor U1323 (N_1323,N_1247,N_1223);
xor U1324 (N_1324,N_1274,N_1270);
xnor U1325 (N_1325,N_1221,N_1200);
nand U1326 (N_1326,N_1247,N_1272);
nand U1327 (N_1327,N_1251,N_1204);
xor U1328 (N_1328,N_1244,N_1226);
xnor U1329 (N_1329,N_1223,N_1200);
nor U1330 (N_1330,N_1274,N_1250);
and U1331 (N_1331,N_1216,N_1210);
or U1332 (N_1332,N_1202,N_1235);
xnor U1333 (N_1333,N_1248,N_1255);
nand U1334 (N_1334,N_1244,N_1228);
or U1335 (N_1335,N_1200,N_1211);
or U1336 (N_1336,N_1206,N_1242);
nand U1337 (N_1337,N_1209,N_1204);
nand U1338 (N_1338,N_1242,N_1200);
xor U1339 (N_1339,N_1216,N_1226);
xor U1340 (N_1340,N_1226,N_1256);
or U1341 (N_1341,N_1249,N_1218);
nand U1342 (N_1342,N_1266,N_1255);
or U1343 (N_1343,N_1255,N_1254);
or U1344 (N_1344,N_1245,N_1212);
nor U1345 (N_1345,N_1247,N_1237);
and U1346 (N_1346,N_1266,N_1225);
xor U1347 (N_1347,N_1216,N_1222);
or U1348 (N_1348,N_1255,N_1216);
xor U1349 (N_1349,N_1226,N_1223);
nor U1350 (N_1350,N_1344,N_1331);
nand U1351 (N_1351,N_1283,N_1293);
nand U1352 (N_1352,N_1278,N_1321);
nand U1353 (N_1353,N_1334,N_1306);
nor U1354 (N_1354,N_1276,N_1338);
and U1355 (N_1355,N_1335,N_1294);
nand U1356 (N_1356,N_1279,N_1347);
or U1357 (N_1357,N_1312,N_1291);
or U1358 (N_1358,N_1307,N_1319);
and U1359 (N_1359,N_1275,N_1325);
or U1360 (N_1360,N_1277,N_1313);
or U1361 (N_1361,N_1339,N_1349);
nand U1362 (N_1362,N_1343,N_1346);
nand U1363 (N_1363,N_1303,N_1284);
and U1364 (N_1364,N_1345,N_1337);
and U1365 (N_1365,N_1295,N_1288);
and U1366 (N_1366,N_1296,N_1327);
or U1367 (N_1367,N_1336,N_1316);
and U1368 (N_1368,N_1305,N_1333);
nand U1369 (N_1369,N_1300,N_1328);
nor U1370 (N_1370,N_1286,N_1340);
nand U1371 (N_1371,N_1309,N_1311);
xnor U1372 (N_1372,N_1285,N_1323);
and U1373 (N_1373,N_1281,N_1297);
xor U1374 (N_1374,N_1342,N_1280);
or U1375 (N_1375,N_1301,N_1329);
or U1376 (N_1376,N_1304,N_1310);
nand U1377 (N_1377,N_1289,N_1292);
nand U1378 (N_1378,N_1318,N_1290);
xnor U1379 (N_1379,N_1320,N_1308);
nor U1380 (N_1380,N_1287,N_1348);
nor U1381 (N_1381,N_1317,N_1326);
xor U1382 (N_1382,N_1324,N_1299);
and U1383 (N_1383,N_1298,N_1302);
and U1384 (N_1384,N_1282,N_1332);
nor U1385 (N_1385,N_1314,N_1330);
nor U1386 (N_1386,N_1315,N_1322);
xor U1387 (N_1387,N_1341,N_1310);
nand U1388 (N_1388,N_1347,N_1294);
nor U1389 (N_1389,N_1314,N_1349);
nor U1390 (N_1390,N_1278,N_1317);
xnor U1391 (N_1391,N_1309,N_1320);
or U1392 (N_1392,N_1299,N_1344);
nor U1393 (N_1393,N_1335,N_1303);
nor U1394 (N_1394,N_1292,N_1322);
or U1395 (N_1395,N_1311,N_1312);
xnor U1396 (N_1396,N_1329,N_1335);
xor U1397 (N_1397,N_1305,N_1340);
xor U1398 (N_1398,N_1332,N_1349);
nand U1399 (N_1399,N_1299,N_1298);
and U1400 (N_1400,N_1333,N_1286);
or U1401 (N_1401,N_1326,N_1331);
xnor U1402 (N_1402,N_1349,N_1329);
or U1403 (N_1403,N_1328,N_1291);
or U1404 (N_1404,N_1282,N_1305);
xor U1405 (N_1405,N_1306,N_1349);
nor U1406 (N_1406,N_1320,N_1318);
and U1407 (N_1407,N_1330,N_1276);
or U1408 (N_1408,N_1276,N_1284);
nor U1409 (N_1409,N_1314,N_1277);
and U1410 (N_1410,N_1290,N_1279);
or U1411 (N_1411,N_1314,N_1331);
nor U1412 (N_1412,N_1343,N_1334);
nor U1413 (N_1413,N_1347,N_1326);
or U1414 (N_1414,N_1281,N_1325);
and U1415 (N_1415,N_1307,N_1335);
xor U1416 (N_1416,N_1305,N_1337);
and U1417 (N_1417,N_1347,N_1333);
or U1418 (N_1418,N_1302,N_1312);
nand U1419 (N_1419,N_1294,N_1320);
nand U1420 (N_1420,N_1319,N_1280);
xor U1421 (N_1421,N_1316,N_1324);
or U1422 (N_1422,N_1283,N_1326);
nand U1423 (N_1423,N_1331,N_1297);
nand U1424 (N_1424,N_1275,N_1284);
or U1425 (N_1425,N_1417,N_1404);
or U1426 (N_1426,N_1382,N_1391);
and U1427 (N_1427,N_1409,N_1401);
nand U1428 (N_1428,N_1405,N_1396);
or U1429 (N_1429,N_1364,N_1419);
nand U1430 (N_1430,N_1381,N_1420);
nand U1431 (N_1431,N_1403,N_1377);
xnor U1432 (N_1432,N_1378,N_1355);
or U1433 (N_1433,N_1386,N_1353);
nand U1434 (N_1434,N_1422,N_1356);
nand U1435 (N_1435,N_1368,N_1350);
and U1436 (N_1436,N_1384,N_1399);
and U1437 (N_1437,N_1366,N_1395);
nor U1438 (N_1438,N_1371,N_1418);
and U1439 (N_1439,N_1352,N_1361);
nor U1440 (N_1440,N_1365,N_1354);
and U1441 (N_1441,N_1413,N_1374);
xnor U1442 (N_1442,N_1394,N_1370);
or U1443 (N_1443,N_1410,N_1383);
and U1444 (N_1444,N_1414,N_1408);
and U1445 (N_1445,N_1407,N_1369);
nand U1446 (N_1446,N_1390,N_1398);
nor U1447 (N_1447,N_1380,N_1415);
and U1448 (N_1448,N_1387,N_1392);
nor U1449 (N_1449,N_1357,N_1360);
and U1450 (N_1450,N_1412,N_1372);
nor U1451 (N_1451,N_1359,N_1389);
nand U1452 (N_1452,N_1351,N_1423);
nor U1453 (N_1453,N_1400,N_1388);
nor U1454 (N_1454,N_1363,N_1424);
nor U1455 (N_1455,N_1406,N_1416);
xnor U1456 (N_1456,N_1358,N_1393);
xor U1457 (N_1457,N_1367,N_1411);
and U1458 (N_1458,N_1385,N_1362);
or U1459 (N_1459,N_1402,N_1376);
and U1460 (N_1460,N_1397,N_1421);
xor U1461 (N_1461,N_1375,N_1379);
and U1462 (N_1462,N_1373,N_1362);
and U1463 (N_1463,N_1371,N_1353);
or U1464 (N_1464,N_1384,N_1363);
and U1465 (N_1465,N_1397,N_1406);
or U1466 (N_1466,N_1405,N_1404);
or U1467 (N_1467,N_1366,N_1384);
nor U1468 (N_1468,N_1372,N_1357);
and U1469 (N_1469,N_1420,N_1392);
or U1470 (N_1470,N_1354,N_1412);
xnor U1471 (N_1471,N_1393,N_1357);
or U1472 (N_1472,N_1356,N_1368);
xor U1473 (N_1473,N_1361,N_1359);
or U1474 (N_1474,N_1419,N_1421);
nand U1475 (N_1475,N_1409,N_1359);
nor U1476 (N_1476,N_1397,N_1402);
nand U1477 (N_1477,N_1374,N_1417);
and U1478 (N_1478,N_1389,N_1422);
xnor U1479 (N_1479,N_1370,N_1356);
xor U1480 (N_1480,N_1365,N_1408);
nand U1481 (N_1481,N_1356,N_1355);
or U1482 (N_1482,N_1365,N_1386);
nand U1483 (N_1483,N_1409,N_1350);
or U1484 (N_1484,N_1363,N_1392);
nand U1485 (N_1485,N_1374,N_1354);
and U1486 (N_1486,N_1376,N_1405);
xor U1487 (N_1487,N_1420,N_1405);
xnor U1488 (N_1488,N_1351,N_1382);
and U1489 (N_1489,N_1362,N_1387);
xor U1490 (N_1490,N_1382,N_1398);
xnor U1491 (N_1491,N_1368,N_1359);
or U1492 (N_1492,N_1394,N_1395);
nand U1493 (N_1493,N_1362,N_1406);
or U1494 (N_1494,N_1383,N_1382);
nor U1495 (N_1495,N_1350,N_1367);
and U1496 (N_1496,N_1402,N_1420);
xnor U1497 (N_1497,N_1399,N_1388);
xor U1498 (N_1498,N_1404,N_1420);
xnor U1499 (N_1499,N_1356,N_1418);
or U1500 (N_1500,N_1466,N_1455);
and U1501 (N_1501,N_1477,N_1489);
and U1502 (N_1502,N_1428,N_1495);
and U1503 (N_1503,N_1443,N_1450);
xnor U1504 (N_1504,N_1451,N_1458);
xnor U1505 (N_1505,N_1426,N_1459);
or U1506 (N_1506,N_1479,N_1481);
and U1507 (N_1507,N_1438,N_1486);
nor U1508 (N_1508,N_1464,N_1470);
xor U1509 (N_1509,N_1442,N_1425);
or U1510 (N_1510,N_1478,N_1427);
or U1511 (N_1511,N_1499,N_1497);
nand U1512 (N_1512,N_1435,N_1431);
xor U1513 (N_1513,N_1444,N_1430);
xor U1514 (N_1514,N_1490,N_1468);
nor U1515 (N_1515,N_1469,N_1465);
nand U1516 (N_1516,N_1491,N_1482);
nor U1517 (N_1517,N_1429,N_1432);
xnor U1518 (N_1518,N_1496,N_1484);
nor U1519 (N_1519,N_1494,N_1456);
or U1520 (N_1520,N_1471,N_1473);
and U1521 (N_1521,N_1434,N_1492);
nand U1522 (N_1522,N_1452,N_1441);
nor U1523 (N_1523,N_1433,N_1493);
and U1524 (N_1524,N_1445,N_1447);
or U1525 (N_1525,N_1474,N_1463);
nand U1526 (N_1526,N_1440,N_1461);
xnor U1527 (N_1527,N_1488,N_1472);
nor U1528 (N_1528,N_1476,N_1460);
or U1529 (N_1529,N_1437,N_1480);
nand U1530 (N_1530,N_1446,N_1498);
nor U1531 (N_1531,N_1439,N_1457);
nor U1532 (N_1532,N_1467,N_1449);
or U1533 (N_1533,N_1485,N_1487);
nand U1534 (N_1534,N_1462,N_1448);
or U1535 (N_1535,N_1475,N_1454);
nand U1536 (N_1536,N_1436,N_1483);
xnor U1537 (N_1537,N_1453,N_1477);
and U1538 (N_1538,N_1431,N_1488);
nor U1539 (N_1539,N_1479,N_1438);
nor U1540 (N_1540,N_1428,N_1472);
nor U1541 (N_1541,N_1448,N_1472);
xor U1542 (N_1542,N_1484,N_1476);
nor U1543 (N_1543,N_1471,N_1497);
xnor U1544 (N_1544,N_1486,N_1445);
xnor U1545 (N_1545,N_1465,N_1438);
nor U1546 (N_1546,N_1497,N_1429);
or U1547 (N_1547,N_1449,N_1487);
xnor U1548 (N_1548,N_1447,N_1486);
nor U1549 (N_1549,N_1457,N_1440);
or U1550 (N_1550,N_1426,N_1495);
nand U1551 (N_1551,N_1483,N_1425);
or U1552 (N_1552,N_1436,N_1448);
nand U1553 (N_1553,N_1496,N_1480);
xor U1554 (N_1554,N_1474,N_1479);
and U1555 (N_1555,N_1490,N_1485);
nor U1556 (N_1556,N_1469,N_1481);
nor U1557 (N_1557,N_1451,N_1486);
or U1558 (N_1558,N_1485,N_1425);
and U1559 (N_1559,N_1461,N_1446);
nor U1560 (N_1560,N_1456,N_1465);
nor U1561 (N_1561,N_1473,N_1440);
and U1562 (N_1562,N_1482,N_1453);
nand U1563 (N_1563,N_1439,N_1435);
or U1564 (N_1564,N_1494,N_1448);
or U1565 (N_1565,N_1445,N_1429);
xor U1566 (N_1566,N_1498,N_1464);
and U1567 (N_1567,N_1462,N_1480);
xor U1568 (N_1568,N_1485,N_1497);
nand U1569 (N_1569,N_1437,N_1489);
or U1570 (N_1570,N_1483,N_1490);
and U1571 (N_1571,N_1448,N_1498);
nand U1572 (N_1572,N_1465,N_1448);
nand U1573 (N_1573,N_1492,N_1486);
or U1574 (N_1574,N_1436,N_1459);
xnor U1575 (N_1575,N_1547,N_1568);
nor U1576 (N_1576,N_1550,N_1556);
and U1577 (N_1577,N_1517,N_1545);
or U1578 (N_1578,N_1565,N_1564);
or U1579 (N_1579,N_1542,N_1562);
nand U1580 (N_1580,N_1539,N_1522);
or U1581 (N_1581,N_1533,N_1554);
nor U1582 (N_1582,N_1532,N_1555);
nand U1583 (N_1583,N_1538,N_1540);
and U1584 (N_1584,N_1510,N_1544);
nor U1585 (N_1585,N_1525,N_1567);
or U1586 (N_1586,N_1536,N_1535);
xnor U1587 (N_1587,N_1546,N_1528);
nand U1588 (N_1588,N_1551,N_1505);
nor U1589 (N_1589,N_1511,N_1553);
or U1590 (N_1590,N_1543,N_1526);
or U1591 (N_1591,N_1541,N_1512);
and U1592 (N_1592,N_1572,N_1515);
and U1593 (N_1593,N_1563,N_1521);
and U1594 (N_1594,N_1502,N_1529);
xor U1595 (N_1595,N_1508,N_1513);
xnor U1596 (N_1596,N_1534,N_1516);
xor U1597 (N_1597,N_1570,N_1524);
nor U1598 (N_1598,N_1506,N_1519);
nor U1599 (N_1599,N_1514,N_1569);
nand U1600 (N_1600,N_1523,N_1549);
nand U1601 (N_1601,N_1561,N_1530);
nor U1602 (N_1602,N_1558,N_1500);
xnor U1603 (N_1603,N_1520,N_1552);
nor U1604 (N_1604,N_1504,N_1571);
xor U1605 (N_1605,N_1518,N_1531);
nand U1606 (N_1606,N_1574,N_1537);
nand U1607 (N_1607,N_1573,N_1566);
or U1608 (N_1608,N_1507,N_1548);
nor U1609 (N_1609,N_1527,N_1560);
or U1610 (N_1610,N_1509,N_1501);
xor U1611 (N_1611,N_1503,N_1559);
nand U1612 (N_1612,N_1557,N_1540);
and U1613 (N_1613,N_1546,N_1553);
or U1614 (N_1614,N_1547,N_1513);
nor U1615 (N_1615,N_1543,N_1565);
and U1616 (N_1616,N_1546,N_1542);
nand U1617 (N_1617,N_1537,N_1547);
nand U1618 (N_1618,N_1523,N_1520);
nor U1619 (N_1619,N_1542,N_1559);
nor U1620 (N_1620,N_1508,N_1550);
xor U1621 (N_1621,N_1561,N_1546);
nand U1622 (N_1622,N_1551,N_1517);
nand U1623 (N_1623,N_1555,N_1544);
or U1624 (N_1624,N_1533,N_1532);
or U1625 (N_1625,N_1514,N_1513);
or U1626 (N_1626,N_1538,N_1549);
and U1627 (N_1627,N_1503,N_1572);
nor U1628 (N_1628,N_1523,N_1516);
or U1629 (N_1629,N_1543,N_1521);
nand U1630 (N_1630,N_1532,N_1573);
xnor U1631 (N_1631,N_1512,N_1560);
xnor U1632 (N_1632,N_1558,N_1535);
and U1633 (N_1633,N_1574,N_1565);
or U1634 (N_1634,N_1563,N_1526);
and U1635 (N_1635,N_1511,N_1515);
and U1636 (N_1636,N_1526,N_1537);
or U1637 (N_1637,N_1532,N_1544);
xnor U1638 (N_1638,N_1517,N_1534);
xor U1639 (N_1639,N_1571,N_1510);
or U1640 (N_1640,N_1528,N_1541);
nand U1641 (N_1641,N_1536,N_1527);
nor U1642 (N_1642,N_1507,N_1508);
and U1643 (N_1643,N_1518,N_1508);
nor U1644 (N_1644,N_1543,N_1557);
nor U1645 (N_1645,N_1549,N_1546);
nor U1646 (N_1646,N_1521,N_1532);
nand U1647 (N_1647,N_1566,N_1535);
and U1648 (N_1648,N_1521,N_1520);
and U1649 (N_1649,N_1545,N_1541);
nand U1650 (N_1650,N_1608,N_1648);
and U1651 (N_1651,N_1649,N_1628);
xor U1652 (N_1652,N_1637,N_1631);
and U1653 (N_1653,N_1575,N_1630);
nor U1654 (N_1654,N_1636,N_1626);
xor U1655 (N_1655,N_1632,N_1588);
nand U1656 (N_1656,N_1581,N_1615);
nor U1657 (N_1657,N_1589,N_1578);
xor U1658 (N_1658,N_1579,N_1611);
and U1659 (N_1659,N_1600,N_1590);
nor U1660 (N_1660,N_1599,N_1629);
nor U1661 (N_1661,N_1597,N_1621);
and U1662 (N_1662,N_1591,N_1624);
nor U1663 (N_1663,N_1592,N_1576);
and U1664 (N_1664,N_1645,N_1607);
nor U1665 (N_1665,N_1596,N_1598);
and U1666 (N_1666,N_1580,N_1585);
and U1667 (N_1667,N_1620,N_1610);
nor U1668 (N_1668,N_1647,N_1618);
nand U1669 (N_1669,N_1617,N_1634);
xnor U1670 (N_1670,N_1577,N_1601);
or U1671 (N_1671,N_1586,N_1604);
and U1672 (N_1672,N_1644,N_1587);
or U1673 (N_1673,N_1595,N_1582);
or U1674 (N_1674,N_1613,N_1605);
xnor U1675 (N_1675,N_1616,N_1619);
nand U1676 (N_1676,N_1614,N_1602);
or U1677 (N_1677,N_1646,N_1635);
or U1678 (N_1678,N_1606,N_1639);
or U1679 (N_1679,N_1633,N_1623);
and U1680 (N_1680,N_1584,N_1641);
xor U1681 (N_1681,N_1622,N_1638);
nand U1682 (N_1682,N_1612,N_1594);
nand U1683 (N_1683,N_1603,N_1625);
xor U1684 (N_1684,N_1593,N_1642);
nor U1685 (N_1685,N_1643,N_1583);
nand U1686 (N_1686,N_1640,N_1609);
xnor U1687 (N_1687,N_1627,N_1586);
nand U1688 (N_1688,N_1635,N_1644);
or U1689 (N_1689,N_1626,N_1621);
or U1690 (N_1690,N_1635,N_1638);
and U1691 (N_1691,N_1623,N_1605);
nor U1692 (N_1692,N_1608,N_1575);
and U1693 (N_1693,N_1609,N_1610);
nor U1694 (N_1694,N_1611,N_1615);
nand U1695 (N_1695,N_1583,N_1629);
or U1696 (N_1696,N_1616,N_1594);
or U1697 (N_1697,N_1606,N_1594);
and U1698 (N_1698,N_1631,N_1615);
nand U1699 (N_1699,N_1647,N_1621);
and U1700 (N_1700,N_1639,N_1593);
or U1701 (N_1701,N_1594,N_1628);
nand U1702 (N_1702,N_1600,N_1588);
or U1703 (N_1703,N_1592,N_1642);
nor U1704 (N_1704,N_1633,N_1649);
nor U1705 (N_1705,N_1598,N_1640);
or U1706 (N_1706,N_1600,N_1589);
and U1707 (N_1707,N_1599,N_1609);
nand U1708 (N_1708,N_1629,N_1594);
nand U1709 (N_1709,N_1594,N_1593);
and U1710 (N_1710,N_1610,N_1595);
nand U1711 (N_1711,N_1581,N_1610);
nand U1712 (N_1712,N_1642,N_1618);
and U1713 (N_1713,N_1596,N_1635);
nor U1714 (N_1714,N_1587,N_1637);
xor U1715 (N_1715,N_1638,N_1581);
nand U1716 (N_1716,N_1641,N_1593);
or U1717 (N_1717,N_1580,N_1589);
and U1718 (N_1718,N_1629,N_1645);
or U1719 (N_1719,N_1598,N_1601);
xnor U1720 (N_1720,N_1599,N_1619);
nor U1721 (N_1721,N_1601,N_1580);
xor U1722 (N_1722,N_1622,N_1616);
nor U1723 (N_1723,N_1617,N_1610);
or U1724 (N_1724,N_1642,N_1614);
xnor U1725 (N_1725,N_1716,N_1692);
and U1726 (N_1726,N_1655,N_1663);
nor U1727 (N_1727,N_1652,N_1714);
nand U1728 (N_1728,N_1681,N_1688);
or U1729 (N_1729,N_1723,N_1662);
or U1730 (N_1730,N_1683,N_1717);
and U1731 (N_1731,N_1710,N_1677);
nor U1732 (N_1732,N_1709,N_1698);
xor U1733 (N_1733,N_1689,N_1706);
or U1734 (N_1734,N_1721,N_1685);
or U1735 (N_1735,N_1659,N_1653);
nor U1736 (N_1736,N_1668,N_1702);
and U1737 (N_1737,N_1674,N_1720);
nand U1738 (N_1738,N_1711,N_1656);
nand U1739 (N_1739,N_1691,N_1682);
xnor U1740 (N_1740,N_1658,N_1672);
nand U1741 (N_1741,N_1669,N_1678);
nand U1742 (N_1742,N_1700,N_1712);
or U1743 (N_1743,N_1693,N_1675);
nand U1744 (N_1744,N_1679,N_1671);
nand U1745 (N_1745,N_1697,N_1650);
or U1746 (N_1746,N_1666,N_1684);
xor U1747 (N_1747,N_1707,N_1673);
nor U1748 (N_1748,N_1719,N_1722);
or U1749 (N_1749,N_1708,N_1699);
xnor U1750 (N_1750,N_1680,N_1657);
nor U1751 (N_1751,N_1660,N_1664);
nand U1752 (N_1752,N_1704,N_1654);
nor U1753 (N_1753,N_1661,N_1705);
xnor U1754 (N_1754,N_1687,N_1703);
xnor U1755 (N_1755,N_1715,N_1718);
nor U1756 (N_1756,N_1665,N_1695);
or U1757 (N_1757,N_1694,N_1713);
nand U1758 (N_1758,N_1651,N_1701);
nand U1759 (N_1759,N_1676,N_1667);
xor U1760 (N_1760,N_1670,N_1724);
or U1761 (N_1761,N_1686,N_1696);
nand U1762 (N_1762,N_1690,N_1662);
nor U1763 (N_1763,N_1652,N_1710);
nand U1764 (N_1764,N_1652,N_1693);
and U1765 (N_1765,N_1660,N_1693);
or U1766 (N_1766,N_1653,N_1678);
nor U1767 (N_1767,N_1669,N_1654);
nand U1768 (N_1768,N_1695,N_1663);
nor U1769 (N_1769,N_1722,N_1708);
xor U1770 (N_1770,N_1665,N_1662);
and U1771 (N_1771,N_1666,N_1723);
nor U1772 (N_1772,N_1671,N_1724);
and U1773 (N_1773,N_1688,N_1722);
and U1774 (N_1774,N_1701,N_1710);
xor U1775 (N_1775,N_1698,N_1655);
nand U1776 (N_1776,N_1679,N_1684);
nand U1777 (N_1777,N_1697,N_1664);
and U1778 (N_1778,N_1676,N_1688);
xor U1779 (N_1779,N_1720,N_1675);
nand U1780 (N_1780,N_1723,N_1713);
nor U1781 (N_1781,N_1653,N_1685);
xor U1782 (N_1782,N_1689,N_1720);
nor U1783 (N_1783,N_1694,N_1677);
xor U1784 (N_1784,N_1718,N_1700);
or U1785 (N_1785,N_1687,N_1716);
nand U1786 (N_1786,N_1659,N_1671);
xnor U1787 (N_1787,N_1691,N_1663);
xnor U1788 (N_1788,N_1693,N_1690);
nand U1789 (N_1789,N_1652,N_1671);
xnor U1790 (N_1790,N_1652,N_1713);
nand U1791 (N_1791,N_1667,N_1652);
and U1792 (N_1792,N_1688,N_1693);
nand U1793 (N_1793,N_1719,N_1667);
xor U1794 (N_1794,N_1655,N_1685);
or U1795 (N_1795,N_1658,N_1654);
xor U1796 (N_1796,N_1671,N_1675);
nand U1797 (N_1797,N_1724,N_1657);
nor U1798 (N_1798,N_1694,N_1698);
and U1799 (N_1799,N_1689,N_1724);
nor U1800 (N_1800,N_1731,N_1795);
and U1801 (N_1801,N_1792,N_1776);
and U1802 (N_1802,N_1726,N_1799);
and U1803 (N_1803,N_1753,N_1780);
xor U1804 (N_1804,N_1783,N_1736);
nand U1805 (N_1805,N_1790,N_1782);
or U1806 (N_1806,N_1770,N_1727);
nor U1807 (N_1807,N_1744,N_1754);
xor U1808 (N_1808,N_1735,N_1785);
or U1809 (N_1809,N_1756,N_1786);
and U1810 (N_1810,N_1757,N_1750);
and U1811 (N_1811,N_1761,N_1774);
nor U1812 (N_1812,N_1771,N_1747);
nand U1813 (N_1813,N_1739,N_1794);
xnor U1814 (N_1814,N_1737,N_1743);
and U1815 (N_1815,N_1729,N_1796);
nor U1816 (N_1816,N_1777,N_1758);
nor U1817 (N_1817,N_1768,N_1730);
nor U1818 (N_1818,N_1784,N_1775);
or U1819 (N_1819,N_1766,N_1791);
xnor U1820 (N_1820,N_1793,N_1765);
or U1821 (N_1821,N_1773,N_1733);
nand U1822 (N_1822,N_1779,N_1788);
nand U1823 (N_1823,N_1755,N_1728);
xor U1824 (N_1824,N_1746,N_1732);
and U1825 (N_1825,N_1738,N_1767);
nor U1826 (N_1826,N_1762,N_1734);
or U1827 (N_1827,N_1742,N_1752);
xor U1828 (N_1828,N_1759,N_1741);
and U1829 (N_1829,N_1769,N_1797);
nor U1830 (N_1830,N_1725,N_1781);
xor U1831 (N_1831,N_1748,N_1789);
nor U1832 (N_1832,N_1760,N_1764);
nand U1833 (N_1833,N_1772,N_1787);
nand U1834 (N_1834,N_1763,N_1740);
xor U1835 (N_1835,N_1751,N_1778);
nor U1836 (N_1836,N_1749,N_1798);
nand U1837 (N_1837,N_1745,N_1776);
xnor U1838 (N_1838,N_1768,N_1755);
nor U1839 (N_1839,N_1748,N_1750);
nor U1840 (N_1840,N_1742,N_1756);
or U1841 (N_1841,N_1762,N_1732);
and U1842 (N_1842,N_1749,N_1791);
nor U1843 (N_1843,N_1768,N_1791);
or U1844 (N_1844,N_1783,N_1728);
and U1845 (N_1845,N_1752,N_1765);
and U1846 (N_1846,N_1758,N_1735);
nor U1847 (N_1847,N_1756,N_1792);
nand U1848 (N_1848,N_1789,N_1749);
nand U1849 (N_1849,N_1787,N_1785);
xor U1850 (N_1850,N_1745,N_1766);
nand U1851 (N_1851,N_1777,N_1794);
nor U1852 (N_1852,N_1734,N_1769);
nand U1853 (N_1853,N_1730,N_1754);
and U1854 (N_1854,N_1778,N_1734);
and U1855 (N_1855,N_1725,N_1746);
or U1856 (N_1856,N_1730,N_1762);
or U1857 (N_1857,N_1796,N_1726);
and U1858 (N_1858,N_1778,N_1773);
xnor U1859 (N_1859,N_1790,N_1776);
nor U1860 (N_1860,N_1784,N_1747);
or U1861 (N_1861,N_1777,N_1735);
xor U1862 (N_1862,N_1746,N_1771);
nand U1863 (N_1863,N_1796,N_1790);
and U1864 (N_1864,N_1789,N_1747);
and U1865 (N_1865,N_1777,N_1764);
nand U1866 (N_1866,N_1728,N_1797);
nor U1867 (N_1867,N_1799,N_1734);
or U1868 (N_1868,N_1758,N_1796);
or U1869 (N_1869,N_1752,N_1789);
or U1870 (N_1870,N_1774,N_1769);
nand U1871 (N_1871,N_1765,N_1772);
nor U1872 (N_1872,N_1782,N_1796);
nor U1873 (N_1873,N_1732,N_1789);
nand U1874 (N_1874,N_1775,N_1743);
nor U1875 (N_1875,N_1865,N_1850);
or U1876 (N_1876,N_1836,N_1863);
nand U1877 (N_1877,N_1848,N_1822);
nand U1878 (N_1878,N_1845,N_1817);
xnor U1879 (N_1879,N_1846,N_1826);
xnor U1880 (N_1880,N_1800,N_1859);
nand U1881 (N_1881,N_1803,N_1809);
and U1882 (N_1882,N_1819,N_1866);
nor U1883 (N_1883,N_1856,N_1862);
and U1884 (N_1884,N_1840,N_1851);
xnor U1885 (N_1885,N_1823,N_1849);
nor U1886 (N_1886,N_1815,N_1816);
or U1887 (N_1887,N_1870,N_1852);
and U1888 (N_1888,N_1802,N_1820);
nand U1889 (N_1889,N_1842,N_1869);
and U1890 (N_1890,N_1830,N_1847);
xnor U1891 (N_1891,N_1868,N_1806);
xnor U1892 (N_1892,N_1841,N_1864);
and U1893 (N_1893,N_1829,N_1818);
or U1894 (N_1894,N_1812,N_1857);
or U1895 (N_1895,N_1874,N_1814);
xor U1896 (N_1896,N_1839,N_1833);
or U1897 (N_1897,N_1837,N_1838);
or U1898 (N_1898,N_1804,N_1824);
or U1899 (N_1899,N_1855,N_1801);
nor U1900 (N_1900,N_1827,N_1825);
nor U1901 (N_1901,N_1873,N_1853);
xor U1902 (N_1902,N_1813,N_1808);
and U1903 (N_1903,N_1805,N_1831);
nand U1904 (N_1904,N_1810,N_1861);
nor U1905 (N_1905,N_1843,N_1872);
nand U1906 (N_1906,N_1858,N_1854);
xor U1907 (N_1907,N_1828,N_1807);
nor U1908 (N_1908,N_1821,N_1832);
nor U1909 (N_1909,N_1811,N_1835);
and U1910 (N_1910,N_1860,N_1867);
and U1911 (N_1911,N_1844,N_1871);
and U1912 (N_1912,N_1834,N_1859);
nor U1913 (N_1913,N_1809,N_1862);
and U1914 (N_1914,N_1870,N_1860);
nor U1915 (N_1915,N_1813,N_1836);
nor U1916 (N_1916,N_1802,N_1822);
xnor U1917 (N_1917,N_1849,N_1818);
xor U1918 (N_1918,N_1871,N_1800);
and U1919 (N_1919,N_1816,N_1871);
and U1920 (N_1920,N_1836,N_1815);
and U1921 (N_1921,N_1808,N_1824);
and U1922 (N_1922,N_1836,N_1841);
and U1923 (N_1923,N_1865,N_1830);
or U1924 (N_1924,N_1862,N_1803);
nor U1925 (N_1925,N_1814,N_1858);
nand U1926 (N_1926,N_1804,N_1801);
nor U1927 (N_1927,N_1853,N_1864);
nor U1928 (N_1928,N_1849,N_1824);
xnor U1929 (N_1929,N_1822,N_1810);
xnor U1930 (N_1930,N_1843,N_1828);
nor U1931 (N_1931,N_1844,N_1838);
xor U1932 (N_1932,N_1814,N_1837);
or U1933 (N_1933,N_1850,N_1873);
or U1934 (N_1934,N_1810,N_1869);
nor U1935 (N_1935,N_1854,N_1860);
and U1936 (N_1936,N_1861,N_1802);
and U1937 (N_1937,N_1838,N_1873);
nor U1938 (N_1938,N_1807,N_1805);
nand U1939 (N_1939,N_1844,N_1869);
or U1940 (N_1940,N_1804,N_1837);
and U1941 (N_1941,N_1854,N_1802);
and U1942 (N_1942,N_1857,N_1865);
nor U1943 (N_1943,N_1837,N_1844);
and U1944 (N_1944,N_1804,N_1819);
or U1945 (N_1945,N_1840,N_1830);
nand U1946 (N_1946,N_1812,N_1839);
or U1947 (N_1947,N_1822,N_1842);
nand U1948 (N_1948,N_1832,N_1801);
nor U1949 (N_1949,N_1862,N_1832);
and U1950 (N_1950,N_1931,N_1946);
and U1951 (N_1951,N_1898,N_1913);
xor U1952 (N_1952,N_1921,N_1888);
nor U1953 (N_1953,N_1914,N_1887);
nor U1954 (N_1954,N_1909,N_1915);
and U1955 (N_1955,N_1884,N_1935);
and U1956 (N_1956,N_1890,N_1896);
and U1957 (N_1957,N_1947,N_1912);
nand U1958 (N_1958,N_1891,N_1889);
xor U1959 (N_1959,N_1902,N_1934);
nand U1960 (N_1960,N_1918,N_1897);
nand U1961 (N_1961,N_1932,N_1886);
xnor U1962 (N_1962,N_1903,N_1920);
xor U1963 (N_1963,N_1901,N_1938);
or U1964 (N_1964,N_1919,N_1875);
or U1965 (N_1965,N_1905,N_1948);
or U1966 (N_1966,N_1916,N_1944);
nand U1967 (N_1967,N_1892,N_1941);
and U1968 (N_1968,N_1940,N_1895);
or U1969 (N_1969,N_1923,N_1930);
or U1970 (N_1970,N_1917,N_1881);
and U1971 (N_1971,N_1882,N_1911);
xnor U1972 (N_1972,N_1885,N_1937);
nor U1973 (N_1973,N_1943,N_1910);
xor U1974 (N_1974,N_1907,N_1877);
or U1975 (N_1975,N_1883,N_1904);
nand U1976 (N_1976,N_1927,N_1929);
xor U1977 (N_1977,N_1900,N_1933);
or U1978 (N_1978,N_1893,N_1939);
and U1979 (N_1979,N_1928,N_1908);
or U1980 (N_1980,N_1922,N_1906);
nand U1981 (N_1981,N_1945,N_1899);
nor U1982 (N_1982,N_1924,N_1880);
xor U1983 (N_1983,N_1926,N_1925);
nand U1984 (N_1984,N_1879,N_1949);
nand U1985 (N_1985,N_1876,N_1878);
and U1986 (N_1986,N_1894,N_1936);
or U1987 (N_1987,N_1942,N_1913);
nand U1988 (N_1988,N_1884,N_1900);
xor U1989 (N_1989,N_1914,N_1928);
or U1990 (N_1990,N_1885,N_1935);
nand U1991 (N_1991,N_1877,N_1929);
and U1992 (N_1992,N_1940,N_1889);
nand U1993 (N_1993,N_1886,N_1881);
and U1994 (N_1994,N_1938,N_1919);
xnor U1995 (N_1995,N_1939,N_1915);
xor U1996 (N_1996,N_1936,N_1940);
nor U1997 (N_1997,N_1890,N_1947);
or U1998 (N_1998,N_1931,N_1912);
nand U1999 (N_1999,N_1880,N_1891);
nor U2000 (N_2000,N_1944,N_1924);
and U2001 (N_2001,N_1879,N_1893);
and U2002 (N_2002,N_1899,N_1881);
nand U2003 (N_2003,N_1920,N_1915);
nand U2004 (N_2004,N_1943,N_1900);
nand U2005 (N_2005,N_1902,N_1938);
or U2006 (N_2006,N_1948,N_1887);
nor U2007 (N_2007,N_1890,N_1920);
or U2008 (N_2008,N_1932,N_1880);
nand U2009 (N_2009,N_1885,N_1923);
and U2010 (N_2010,N_1938,N_1898);
xor U2011 (N_2011,N_1936,N_1943);
nand U2012 (N_2012,N_1884,N_1897);
or U2013 (N_2013,N_1890,N_1930);
nand U2014 (N_2014,N_1910,N_1946);
xnor U2015 (N_2015,N_1896,N_1881);
or U2016 (N_2016,N_1881,N_1919);
xnor U2017 (N_2017,N_1917,N_1901);
xor U2018 (N_2018,N_1946,N_1890);
and U2019 (N_2019,N_1930,N_1884);
and U2020 (N_2020,N_1945,N_1889);
nor U2021 (N_2021,N_1885,N_1916);
or U2022 (N_2022,N_1926,N_1937);
and U2023 (N_2023,N_1879,N_1908);
xor U2024 (N_2024,N_1896,N_1930);
nand U2025 (N_2025,N_1976,N_2023);
nand U2026 (N_2026,N_1984,N_1971);
and U2027 (N_2027,N_2000,N_1995);
nand U2028 (N_2028,N_1954,N_1990);
nand U2029 (N_2029,N_2022,N_1957);
nor U2030 (N_2030,N_2019,N_2009);
xnor U2031 (N_2031,N_2001,N_2008);
or U2032 (N_2032,N_1999,N_1985);
and U2033 (N_2033,N_1967,N_1956);
nand U2034 (N_2034,N_2013,N_2024);
or U2035 (N_2035,N_2005,N_1950);
xor U2036 (N_2036,N_2016,N_1975);
and U2037 (N_2037,N_1993,N_2010);
nand U2038 (N_2038,N_2015,N_1968);
and U2039 (N_2039,N_1988,N_1964);
nor U2040 (N_2040,N_2007,N_1994);
or U2041 (N_2041,N_1960,N_1963);
nand U2042 (N_2042,N_1998,N_1955);
or U2043 (N_2043,N_1959,N_1974);
nand U2044 (N_2044,N_2014,N_1983);
xnor U2045 (N_2045,N_1972,N_1962);
nand U2046 (N_2046,N_1969,N_1989);
and U2047 (N_2047,N_1986,N_1966);
nor U2048 (N_2048,N_1992,N_2004);
nor U2049 (N_2049,N_2020,N_1952);
xor U2050 (N_2050,N_1965,N_1978);
or U2051 (N_2051,N_1997,N_1953);
and U2052 (N_2052,N_2006,N_1987);
nor U2053 (N_2053,N_2017,N_1996);
nor U2054 (N_2054,N_1977,N_2011);
and U2055 (N_2055,N_1991,N_2021);
nor U2056 (N_2056,N_2018,N_2003);
nor U2057 (N_2057,N_1979,N_2002);
nor U2058 (N_2058,N_1951,N_1981);
and U2059 (N_2059,N_1982,N_1970);
nand U2060 (N_2060,N_1980,N_2012);
or U2061 (N_2061,N_1973,N_1958);
nor U2062 (N_2062,N_1961,N_1980);
xnor U2063 (N_2063,N_2001,N_1991);
or U2064 (N_2064,N_2010,N_1996);
or U2065 (N_2065,N_2021,N_2001);
nand U2066 (N_2066,N_2024,N_1974);
nor U2067 (N_2067,N_1957,N_1965);
nand U2068 (N_2068,N_1964,N_1972);
or U2069 (N_2069,N_1994,N_1963);
or U2070 (N_2070,N_1970,N_1980);
nand U2071 (N_2071,N_1956,N_1999);
nor U2072 (N_2072,N_1975,N_2024);
and U2073 (N_2073,N_1961,N_1952);
nand U2074 (N_2074,N_1977,N_1960);
nand U2075 (N_2075,N_1973,N_2020);
and U2076 (N_2076,N_1978,N_1959);
nor U2077 (N_2077,N_2005,N_1976);
or U2078 (N_2078,N_1962,N_1976);
and U2079 (N_2079,N_1966,N_2004);
nand U2080 (N_2080,N_1962,N_2023);
and U2081 (N_2081,N_2010,N_1975);
xnor U2082 (N_2082,N_2000,N_2005);
nor U2083 (N_2083,N_2012,N_2019);
and U2084 (N_2084,N_1968,N_1967);
nand U2085 (N_2085,N_2018,N_2011);
and U2086 (N_2086,N_2013,N_1997);
or U2087 (N_2087,N_2018,N_1950);
nor U2088 (N_2088,N_1989,N_1963);
nor U2089 (N_2089,N_1975,N_1961);
and U2090 (N_2090,N_1971,N_2022);
or U2091 (N_2091,N_1981,N_2009);
or U2092 (N_2092,N_2015,N_2006);
nand U2093 (N_2093,N_1951,N_2021);
nor U2094 (N_2094,N_2018,N_2001);
or U2095 (N_2095,N_2010,N_2020);
or U2096 (N_2096,N_2013,N_2020);
nor U2097 (N_2097,N_1957,N_1972);
nand U2098 (N_2098,N_1953,N_2017);
nand U2099 (N_2099,N_1955,N_1950);
nor U2100 (N_2100,N_2073,N_2040);
nor U2101 (N_2101,N_2025,N_2061);
nor U2102 (N_2102,N_2029,N_2049);
nor U2103 (N_2103,N_2098,N_2084);
nand U2104 (N_2104,N_2043,N_2069);
and U2105 (N_2105,N_2042,N_2054);
and U2106 (N_2106,N_2027,N_2060);
and U2107 (N_2107,N_2070,N_2089);
and U2108 (N_2108,N_2074,N_2063);
and U2109 (N_2109,N_2062,N_2035);
or U2110 (N_2110,N_2068,N_2026);
xnor U2111 (N_2111,N_2065,N_2097);
and U2112 (N_2112,N_2033,N_2090);
or U2113 (N_2113,N_2076,N_2047);
xor U2114 (N_2114,N_2051,N_2092);
nand U2115 (N_2115,N_2077,N_2080);
xnor U2116 (N_2116,N_2099,N_2048);
and U2117 (N_2117,N_2082,N_2059);
and U2118 (N_2118,N_2066,N_2087);
or U2119 (N_2119,N_2058,N_2088);
and U2120 (N_2120,N_2079,N_2056);
xnor U2121 (N_2121,N_2045,N_2091);
nand U2122 (N_2122,N_2036,N_2034);
and U2123 (N_2123,N_2085,N_2064);
xnor U2124 (N_2124,N_2030,N_2095);
xnor U2125 (N_2125,N_2032,N_2072);
nand U2126 (N_2126,N_2078,N_2057);
nor U2127 (N_2127,N_2046,N_2094);
xnor U2128 (N_2128,N_2067,N_2093);
or U2129 (N_2129,N_2053,N_2081);
xor U2130 (N_2130,N_2083,N_2039);
and U2131 (N_2131,N_2038,N_2050);
nor U2132 (N_2132,N_2031,N_2041);
nand U2133 (N_2133,N_2075,N_2052);
nor U2134 (N_2134,N_2086,N_2055);
or U2135 (N_2135,N_2037,N_2044);
and U2136 (N_2136,N_2071,N_2096);
nor U2137 (N_2137,N_2028,N_2092);
xor U2138 (N_2138,N_2092,N_2057);
and U2139 (N_2139,N_2076,N_2098);
or U2140 (N_2140,N_2090,N_2055);
nand U2141 (N_2141,N_2085,N_2045);
nand U2142 (N_2142,N_2095,N_2026);
or U2143 (N_2143,N_2090,N_2057);
xor U2144 (N_2144,N_2044,N_2048);
nor U2145 (N_2145,N_2088,N_2073);
nand U2146 (N_2146,N_2088,N_2087);
or U2147 (N_2147,N_2067,N_2072);
or U2148 (N_2148,N_2094,N_2055);
nor U2149 (N_2149,N_2084,N_2067);
nand U2150 (N_2150,N_2093,N_2083);
nand U2151 (N_2151,N_2095,N_2050);
nor U2152 (N_2152,N_2047,N_2081);
nand U2153 (N_2153,N_2094,N_2043);
nand U2154 (N_2154,N_2079,N_2042);
xnor U2155 (N_2155,N_2033,N_2044);
or U2156 (N_2156,N_2044,N_2089);
and U2157 (N_2157,N_2094,N_2047);
or U2158 (N_2158,N_2035,N_2061);
xor U2159 (N_2159,N_2099,N_2095);
xnor U2160 (N_2160,N_2073,N_2056);
nor U2161 (N_2161,N_2086,N_2054);
nand U2162 (N_2162,N_2048,N_2064);
nor U2163 (N_2163,N_2068,N_2083);
and U2164 (N_2164,N_2035,N_2052);
nand U2165 (N_2165,N_2043,N_2088);
or U2166 (N_2166,N_2038,N_2041);
nand U2167 (N_2167,N_2041,N_2047);
or U2168 (N_2168,N_2049,N_2031);
or U2169 (N_2169,N_2039,N_2088);
nor U2170 (N_2170,N_2098,N_2062);
nor U2171 (N_2171,N_2026,N_2087);
xor U2172 (N_2172,N_2029,N_2099);
and U2173 (N_2173,N_2074,N_2026);
nand U2174 (N_2174,N_2046,N_2080);
xor U2175 (N_2175,N_2124,N_2115);
nand U2176 (N_2176,N_2134,N_2164);
or U2177 (N_2177,N_2147,N_2165);
xnor U2178 (N_2178,N_2114,N_2159);
or U2179 (N_2179,N_2100,N_2158);
nor U2180 (N_2180,N_2130,N_2135);
nand U2181 (N_2181,N_2138,N_2104);
and U2182 (N_2182,N_2125,N_2121);
nand U2183 (N_2183,N_2108,N_2161);
nor U2184 (N_2184,N_2131,N_2143);
and U2185 (N_2185,N_2122,N_2106);
xnor U2186 (N_2186,N_2169,N_2101);
and U2187 (N_2187,N_2154,N_2155);
xor U2188 (N_2188,N_2146,N_2112);
and U2189 (N_2189,N_2156,N_2126);
or U2190 (N_2190,N_2133,N_2137);
nand U2191 (N_2191,N_2153,N_2149);
xor U2192 (N_2192,N_2113,N_2111);
or U2193 (N_2193,N_2148,N_2118);
nor U2194 (N_2194,N_2116,N_2152);
nor U2195 (N_2195,N_2107,N_2136);
or U2196 (N_2196,N_2110,N_2109);
xnor U2197 (N_2197,N_2162,N_2168);
and U2198 (N_2198,N_2132,N_2170);
or U2199 (N_2199,N_2142,N_2139);
and U2200 (N_2200,N_2117,N_2173);
and U2201 (N_2201,N_2105,N_2119);
nand U2202 (N_2202,N_2127,N_2103);
or U2203 (N_2203,N_2145,N_2129);
xor U2204 (N_2204,N_2157,N_2120);
nand U2205 (N_2205,N_2144,N_2172);
or U2206 (N_2206,N_2151,N_2102);
and U2207 (N_2207,N_2166,N_2128);
and U2208 (N_2208,N_2140,N_2160);
nand U2209 (N_2209,N_2171,N_2141);
or U2210 (N_2210,N_2150,N_2167);
nand U2211 (N_2211,N_2163,N_2123);
and U2212 (N_2212,N_2174,N_2126);
nor U2213 (N_2213,N_2137,N_2125);
xor U2214 (N_2214,N_2124,N_2114);
xnor U2215 (N_2215,N_2134,N_2122);
or U2216 (N_2216,N_2146,N_2137);
nor U2217 (N_2217,N_2134,N_2158);
or U2218 (N_2218,N_2124,N_2159);
nor U2219 (N_2219,N_2102,N_2114);
nand U2220 (N_2220,N_2155,N_2173);
xor U2221 (N_2221,N_2165,N_2122);
or U2222 (N_2222,N_2149,N_2163);
or U2223 (N_2223,N_2102,N_2123);
and U2224 (N_2224,N_2102,N_2141);
or U2225 (N_2225,N_2140,N_2174);
nor U2226 (N_2226,N_2173,N_2118);
and U2227 (N_2227,N_2150,N_2142);
nor U2228 (N_2228,N_2168,N_2166);
and U2229 (N_2229,N_2122,N_2161);
nand U2230 (N_2230,N_2152,N_2160);
and U2231 (N_2231,N_2146,N_2120);
and U2232 (N_2232,N_2112,N_2147);
nor U2233 (N_2233,N_2148,N_2163);
and U2234 (N_2234,N_2144,N_2102);
xor U2235 (N_2235,N_2160,N_2115);
and U2236 (N_2236,N_2101,N_2106);
or U2237 (N_2237,N_2106,N_2126);
nor U2238 (N_2238,N_2159,N_2117);
and U2239 (N_2239,N_2107,N_2158);
or U2240 (N_2240,N_2124,N_2121);
xor U2241 (N_2241,N_2124,N_2112);
or U2242 (N_2242,N_2126,N_2170);
and U2243 (N_2243,N_2119,N_2133);
nand U2244 (N_2244,N_2157,N_2145);
and U2245 (N_2245,N_2123,N_2168);
xor U2246 (N_2246,N_2102,N_2137);
nand U2247 (N_2247,N_2102,N_2111);
or U2248 (N_2248,N_2143,N_2129);
nor U2249 (N_2249,N_2135,N_2147);
or U2250 (N_2250,N_2211,N_2183);
xnor U2251 (N_2251,N_2221,N_2182);
xor U2252 (N_2252,N_2242,N_2247);
xnor U2253 (N_2253,N_2234,N_2217);
and U2254 (N_2254,N_2225,N_2243);
and U2255 (N_2255,N_2226,N_2201);
or U2256 (N_2256,N_2240,N_2185);
and U2257 (N_2257,N_2215,N_2204);
xnor U2258 (N_2258,N_2219,N_2177);
or U2259 (N_2259,N_2244,N_2200);
nor U2260 (N_2260,N_2197,N_2237);
or U2261 (N_2261,N_2212,N_2248);
nor U2262 (N_2262,N_2199,N_2239);
nand U2263 (N_2263,N_2229,N_2224);
xnor U2264 (N_2264,N_2186,N_2246);
or U2265 (N_2265,N_2238,N_2232);
nor U2266 (N_2266,N_2190,N_2202);
or U2267 (N_2267,N_2188,N_2194);
and U2268 (N_2268,N_2210,N_2227);
xor U2269 (N_2269,N_2218,N_2213);
and U2270 (N_2270,N_2245,N_2230);
nand U2271 (N_2271,N_2193,N_2198);
nor U2272 (N_2272,N_2233,N_2175);
nand U2273 (N_2273,N_2206,N_2216);
and U2274 (N_2274,N_2214,N_2180);
nand U2275 (N_2275,N_2220,N_2236);
xor U2276 (N_2276,N_2184,N_2189);
nor U2277 (N_2277,N_2178,N_2187);
and U2278 (N_2278,N_2192,N_2191);
nor U2279 (N_2279,N_2179,N_2223);
or U2280 (N_2280,N_2203,N_2176);
nand U2281 (N_2281,N_2231,N_2241);
or U2282 (N_2282,N_2207,N_2181);
nor U2283 (N_2283,N_2195,N_2208);
and U2284 (N_2284,N_2205,N_2249);
xor U2285 (N_2285,N_2196,N_2228);
or U2286 (N_2286,N_2235,N_2209);
and U2287 (N_2287,N_2222,N_2213);
nand U2288 (N_2288,N_2203,N_2213);
or U2289 (N_2289,N_2196,N_2246);
nor U2290 (N_2290,N_2216,N_2193);
xor U2291 (N_2291,N_2186,N_2195);
or U2292 (N_2292,N_2240,N_2200);
nor U2293 (N_2293,N_2201,N_2229);
nand U2294 (N_2294,N_2242,N_2220);
and U2295 (N_2295,N_2226,N_2231);
nand U2296 (N_2296,N_2246,N_2234);
nand U2297 (N_2297,N_2193,N_2184);
nand U2298 (N_2298,N_2244,N_2231);
xnor U2299 (N_2299,N_2244,N_2195);
nand U2300 (N_2300,N_2205,N_2186);
nand U2301 (N_2301,N_2198,N_2212);
nor U2302 (N_2302,N_2221,N_2199);
or U2303 (N_2303,N_2216,N_2195);
xor U2304 (N_2304,N_2228,N_2216);
and U2305 (N_2305,N_2195,N_2247);
nor U2306 (N_2306,N_2214,N_2201);
or U2307 (N_2307,N_2246,N_2175);
nand U2308 (N_2308,N_2246,N_2233);
nor U2309 (N_2309,N_2192,N_2234);
nand U2310 (N_2310,N_2249,N_2238);
nand U2311 (N_2311,N_2221,N_2187);
nor U2312 (N_2312,N_2191,N_2224);
or U2313 (N_2313,N_2193,N_2188);
nor U2314 (N_2314,N_2176,N_2201);
xnor U2315 (N_2315,N_2211,N_2202);
xnor U2316 (N_2316,N_2188,N_2244);
nor U2317 (N_2317,N_2204,N_2193);
nor U2318 (N_2318,N_2221,N_2227);
nor U2319 (N_2319,N_2178,N_2239);
and U2320 (N_2320,N_2214,N_2213);
and U2321 (N_2321,N_2240,N_2201);
and U2322 (N_2322,N_2207,N_2209);
nor U2323 (N_2323,N_2231,N_2238);
or U2324 (N_2324,N_2223,N_2222);
or U2325 (N_2325,N_2289,N_2277);
nand U2326 (N_2326,N_2262,N_2295);
and U2327 (N_2327,N_2272,N_2282);
or U2328 (N_2328,N_2261,N_2322);
or U2329 (N_2329,N_2302,N_2273);
or U2330 (N_2330,N_2321,N_2290);
and U2331 (N_2331,N_2299,N_2253);
nand U2332 (N_2332,N_2279,N_2259);
nand U2333 (N_2333,N_2264,N_2254);
nand U2334 (N_2334,N_2260,N_2265);
xnor U2335 (N_2335,N_2269,N_2306);
nor U2336 (N_2336,N_2276,N_2263);
and U2337 (N_2337,N_2266,N_2256);
nand U2338 (N_2338,N_2316,N_2257);
and U2339 (N_2339,N_2280,N_2323);
xnor U2340 (N_2340,N_2297,N_2284);
or U2341 (N_2341,N_2281,N_2296);
or U2342 (N_2342,N_2304,N_2294);
or U2343 (N_2343,N_2298,N_2275);
xor U2344 (N_2344,N_2309,N_2317);
xor U2345 (N_2345,N_2301,N_2252);
and U2346 (N_2346,N_2287,N_2324);
nor U2347 (N_2347,N_2314,N_2271);
nor U2348 (N_2348,N_2258,N_2283);
xnor U2349 (N_2349,N_2255,N_2311);
and U2350 (N_2350,N_2315,N_2268);
nor U2351 (N_2351,N_2305,N_2288);
or U2352 (N_2352,N_2320,N_2292);
and U2353 (N_2353,N_2251,N_2274);
nor U2354 (N_2354,N_2285,N_2270);
or U2355 (N_2355,N_2312,N_2267);
and U2356 (N_2356,N_2293,N_2307);
nand U2357 (N_2357,N_2250,N_2308);
nor U2358 (N_2358,N_2300,N_2318);
nand U2359 (N_2359,N_2286,N_2291);
nand U2360 (N_2360,N_2319,N_2278);
xor U2361 (N_2361,N_2303,N_2313);
xnor U2362 (N_2362,N_2310,N_2313);
nand U2363 (N_2363,N_2321,N_2305);
and U2364 (N_2364,N_2256,N_2323);
xnor U2365 (N_2365,N_2319,N_2311);
nor U2366 (N_2366,N_2315,N_2253);
nand U2367 (N_2367,N_2262,N_2303);
and U2368 (N_2368,N_2324,N_2322);
xnor U2369 (N_2369,N_2295,N_2287);
and U2370 (N_2370,N_2312,N_2316);
or U2371 (N_2371,N_2314,N_2261);
xnor U2372 (N_2372,N_2300,N_2290);
nor U2373 (N_2373,N_2297,N_2282);
nand U2374 (N_2374,N_2312,N_2299);
xnor U2375 (N_2375,N_2304,N_2299);
or U2376 (N_2376,N_2320,N_2275);
xor U2377 (N_2377,N_2274,N_2256);
xor U2378 (N_2378,N_2293,N_2292);
and U2379 (N_2379,N_2322,N_2281);
or U2380 (N_2380,N_2300,N_2256);
nand U2381 (N_2381,N_2275,N_2306);
or U2382 (N_2382,N_2303,N_2281);
xor U2383 (N_2383,N_2270,N_2324);
nand U2384 (N_2384,N_2299,N_2317);
xor U2385 (N_2385,N_2306,N_2319);
xor U2386 (N_2386,N_2304,N_2259);
nor U2387 (N_2387,N_2315,N_2321);
and U2388 (N_2388,N_2306,N_2303);
xnor U2389 (N_2389,N_2262,N_2292);
nand U2390 (N_2390,N_2251,N_2275);
xor U2391 (N_2391,N_2306,N_2283);
nand U2392 (N_2392,N_2264,N_2295);
nor U2393 (N_2393,N_2252,N_2280);
xnor U2394 (N_2394,N_2274,N_2262);
nor U2395 (N_2395,N_2291,N_2313);
nand U2396 (N_2396,N_2317,N_2269);
xnor U2397 (N_2397,N_2315,N_2257);
or U2398 (N_2398,N_2296,N_2270);
or U2399 (N_2399,N_2272,N_2292);
xnor U2400 (N_2400,N_2329,N_2398);
and U2401 (N_2401,N_2362,N_2366);
and U2402 (N_2402,N_2392,N_2331);
or U2403 (N_2403,N_2396,N_2381);
xor U2404 (N_2404,N_2387,N_2335);
nor U2405 (N_2405,N_2349,N_2360);
nor U2406 (N_2406,N_2343,N_2374);
or U2407 (N_2407,N_2326,N_2380);
and U2408 (N_2408,N_2399,N_2325);
or U2409 (N_2409,N_2384,N_2375);
and U2410 (N_2410,N_2345,N_2365);
xnor U2411 (N_2411,N_2342,N_2344);
nor U2412 (N_2412,N_2378,N_2334);
and U2413 (N_2413,N_2368,N_2379);
or U2414 (N_2414,N_2397,N_2341);
nand U2415 (N_2415,N_2359,N_2388);
nand U2416 (N_2416,N_2376,N_2393);
nor U2417 (N_2417,N_2337,N_2357);
nor U2418 (N_2418,N_2382,N_2372);
nor U2419 (N_2419,N_2367,N_2356);
xnor U2420 (N_2420,N_2371,N_2373);
nor U2421 (N_2421,N_2354,N_2355);
nor U2422 (N_2422,N_2347,N_2358);
xor U2423 (N_2423,N_2346,N_2377);
nor U2424 (N_2424,N_2351,N_2332);
nor U2425 (N_2425,N_2340,N_2389);
nor U2426 (N_2426,N_2352,N_2395);
nand U2427 (N_2427,N_2330,N_2339);
or U2428 (N_2428,N_2390,N_2394);
nand U2429 (N_2429,N_2369,N_2348);
xor U2430 (N_2430,N_2361,N_2363);
and U2431 (N_2431,N_2364,N_2338);
and U2432 (N_2432,N_2336,N_2350);
and U2433 (N_2433,N_2370,N_2333);
or U2434 (N_2434,N_2328,N_2385);
or U2435 (N_2435,N_2391,N_2353);
nand U2436 (N_2436,N_2386,N_2383);
xnor U2437 (N_2437,N_2327,N_2393);
nor U2438 (N_2438,N_2358,N_2391);
xor U2439 (N_2439,N_2387,N_2343);
or U2440 (N_2440,N_2377,N_2398);
nand U2441 (N_2441,N_2368,N_2348);
and U2442 (N_2442,N_2333,N_2337);
or U2443 (N_2443,N_2371,N_2346);
or U2444 (N_2444,N_2371,N_2331);
or U2445 (N_2445,N_2342,N_2380);
nand U2446 (N_2446,N_2357,N_2333);
nor U2447 (N_2447,N_2387,N_2351);
xnor U2448 (N_2448,N_2385,N_2392);
and U2449 (N_2449,N_2389,N_2331);
and U2450 (N_2450,N_2334,N_2339);
or U2451 (N_2451,N_2353,N_2344);
nand U2452 (N_2452,N_2392,N_2332);
or U2453 (N_2453,N_2339,N_2351);
nor U2454 (N_2454,N_2327,N_2337);
nand U2455 (N_2455,N_2341,N_2378);
nor U2456 (N_2456,N_2374,N_2353);
or U2457 (N_2457,N_2328,N_2371);
nor U2458 (N_2458,N_2328,N_2395);
or U2459 (N_2459,N_2362,N_2367);
nor U2460 (N_2460,N_2376,N_2342);
xor U2461 (N_2461,N_2363,N_2390);
nand U2462 (N_2462,N_2339,N_2344);
or U2463 (N_2463,N_2340,N_2350);
nand U2464 (N_2464,N_2343,N_2354);
xor U2465 (N_2465,N_2360,N_2379);
nand U2466 (N_2466,N_2355,N_2353);
nand U2467 (N_2467,N_2347,N_2386);
or U2468 (N_2468,N_2360,N_2394);
and U2469 (N_2469,N_2348,N_2341);
or U2470 (N_2470,N_2326,N_2333);
xor U2471 (N_2471,N_2349,N_2345);
nand U2472 (N_2472,N_2383,N_2372);
or U2473 (N_2473,N_2347,N_2374);
nor U2474 (N_2474,N_2347,N_2345);
nand U2475 (N_2475,N_2469,N_2458);
nand U2476 (N_2476,N_2416,N_2415);
nor U2477 (N_2477,N_2450,N_2446);
or U2478 (N_2478,N_2465,N_2441);
nand U2479 (N_2479,N_2466,N_2462);
and U2480 (N_2480,N_2431,N_2440);
or U2481 (N_2481,N_2447,N_2412);
nand U2482 (N_2482,N_2470,N_2407);
and U2483 (N_2483,N_2464,N_2402);
or U2484 (N_2484,N_2445,N_2435);
and U2485 (N_2485,N_2472,N_2424);
and U2486 (N_2486,N_2443,N_2461);
xor U2487 (N_2487,N_2409,N_2460);
nor U2488 (N_2488,N_2400,N_2423);
and U2489 (N_2489,N_2429,N_2427);
or U2490 (N_2490,N_2442,N_2434);
nand U2491 (N_2491,N_2422,N_2438);
and U2492 (N_2492,N_2428,N_2404);
or U2493 (N_2493,N_2413,N_2432);
nand U2494 (N_2494,N_2401,N_2454);
xnor U2495 (N_2495,N_2430,N_2439);
nand U2496 (N_2496,N_2456,N_2437);
nor U2497 (N_2497,N_2406,N_2468);
nor U2498 (N_2498,N_2451,N_2463);
nor U2499 (N_2499,N_2449,N_2408);
nor U2500 (N_2500,N_2403,N_2471);
nor U2501 (N_2501,N_2453,N_2420);
and U2502 (N_2502,N_2436,N_2452);
and U2503 (N_2503,N_2459,N_2473);
nand U2504 (N_2504,N_2419,N_2474);
nor U2505 (N_2505,N_2455,N_2444);
and U2506 (N_2506,N_2457,N_2417);
or U2507 (N_2507,N_2411,N_2448);
and U2508 (N_2508,N_2421,N_2425);
or U2509 (N_2509,N_2405,N_2410);
or U2510 (N_2510,N_2467,N_2414);
xnor U2511 (N_2511,N_2433,N_2418);
or U2512 (N_2512,N_2426,N_2470);
and U2513 (N_2513,N_2418,N_2460);
nand U2514 (N_2514,N_2424,N_2404);
nor U2515 (N_2515,N_2448,N_2435);
or U2516 (N_2516,N_2409,N_2463);
or U2517 (N_2517,N_2444,N_2422);
or U2518 (N_2518,N_2456,N_2460);
or U2519 (N_2519,N_2431,N_2409);
and U2520 (N_2520,N_2460,N_2431);
nand U2521 (N_2521,N_2460,N_2438);
or U2522 (N_2522,N_2405,N_2452);
xor U2523 (N_2523,N_2406,N_2410);
xor U2524 (N_2524,N_2408,N_2460);
nand U2525 (N_2525,N_2472,N_2438);
nor U2526 (N_2526,N_2405,N_2407);
nor U2527 (N_2527,N_2412,N_2405);
nor U2528 (N_2528,N_2472,N_2413);
nor U2529 (N_2529,N_2467,N_2465);
nand U2530 (N_2530,N_2448,N_2406);
or U2531 (N_2531,N_2441,N_2433);
and U2532 (N_2532,N_2471,N_2446);
nor U2533 (N_2533,N_2446,N_2465);
xnor U2534 (N_2534,N_2429,N_2446);
xor U2535 (N_2535,N_2446,N_2425);
nand U2536 (N_2536,N_2434,N_2458);
nand U2537 (N_2537,N_2472,N_2403);
nand U2538 (N_2538,N_2468,N_2463);
nor U2539 (N_2539,N_2431,N_2444);
xnor U2540 (N_2540,N_2451,N_2447);
nand U2541 (N_2541,N_2474,N_2450);
xnor U2542 (N_2542,N_2433,N_2454);
and U2543 (N_2543,N_2471,N_2428);
and U2544 (N_2544,N_2400,N_2461);
nand U2545 (N_2545,N_2471,N_2447);
or U2546 (N_2546,N_2413,N_2401);
and U2547 (N_2547,N_2422,N_2455);
nand U2548 (N_2548,N_2458,N_2471);
and U2549 (N_2549,N_2407,N_2458);
nor U2550 (N_2550,N_2496,N_2545);
xnor U2551 (N_2551,N_2521,N_2507);
or U2552 (N_2552,N_2505,N_2548);
nand U2553 (N_2553,N_2504,N_2487);
nand U2554 (N_2554,N_2492,N_2499);
and U2555 (N_2555,N_2485,N_2530);
and U2556 (N_2556,N_2482,N_2518);
or U2557 (N_2557,N_2476,N_2479);
nand U2558 (N_2558,N_2519,N_2490);
xnor U2559 (N_2559,N_2486,N_2533);
nand U2560 (N_2560,N_2495,N_2547);
or U2561 (N_2561,N_2516,N_2475);
or U2562 (N_2562,N_2529,N_2549);
xor U2563 (N_2563,N_2526,N_2524);
and U2564 (N_2564,N_2506,N_2528);
or U2565 (N_2565,N_2512,N_2494);
nor U2566 (N_2566,N_2498,N_2478);
or U2567 (N_2567,N_2546,N_2538);
xnor U2568 (N_2568,N_2509,N_2489);
or U2569 (N_2569,N_2523,N_2532);
xor U2570 (N_2570,N_2511,N_2517);
xor U2571 (N_2571,N_2502,N_2527);
nand U2572 (N_2572,N_2540,N_2542);
or U2573 (N_2573,N_2543,N_2513);
nand U2574 (N_2574,N_2536,N_2493);
nand U2575 (N_2575,N_2484,N_2531);
nand U2576 (N_2576,N_2480,N_2483);
nor U2577 (N_2577,N_2539,N_2501);
and U2578 (N_2578,N_2481,N_2544);
or U2579 (N_2579,N_2522,N_2503);
or U2580 (N_2580,N_2510,N_2508);
and U2581 (N_2581,N_2488,N_2500);
nor U2582 (N_2582,N_2491,N_2514);
nand U2583 (N_2583,N_2534,N_2537);
and U2584 (N_2584,N_2541,N_2477);
nand U2585 (N_2585,N_2497,N_2515);
xnor U2586 (N_2586,N_2535,N_2525);
nor U2587 (N_2587,N_2520,N_2497);
nand U2588 (N_2588,N_2502,N_2506);
or U2589 (N_2589,N_2532,N_2486);
or U2590 (N_2590,N_2526,N_2500);
nor U2591 (N_2591,N_2529,N_2503);
nand U2592 (N_2592,N_2530,N_2529);
nor U2593 (N_2593,N_2501,N_2502);
nor U2594 (N_2594,N_2497,N_2479);
nor U2595 (N_2595,N_2507,N_2539);
and U2596 (N_2596,N_2477,N_2547);
xor U2597 (N_2597,N_2525,N_2489);
and U2598 (N_2598,N_2524,N_2525);
nor U2599 (N_2599,N_2480,N_2508);
or U2600 (N_2600,N_2526,N_2501);
nor U2601 (N_2601,N_2485,N_2515);
xnor U2602 (N_2602,N_2537,N_2505);
nor U2603 (N_2603,N_2549,N_2476);
or U2604 (N_2604,N_2518,N_2535);
or U2605 (N_2605,N_2532,N_2543);
or U2606 (N_2606,N_2537,N_2513);
and U2607 (N_2607,N_2512,N_2534);
and U2608 (N_2608,N_2490,N_2536);
and U2609 (N_2609,N_2528,N_2499);
nand U2610 (N_2610,N_2536,N_2519);
and U2611 (N_2611,N_2477,N_2502);
and U2612 (N_2612,N_2493,N_2498);
or U2613 (N_2613,N_2529,N_2517);
nand U2614 (N_2614,N_2485,N_2540);
and U2615 (N_2615,N_2518,N_2506);
xnor U2616 (N_2616,N_2539,N_2505);
nand U2617 (N_2617,N_2483,N_2512);
nor U2618 (N_2618,N_2476,N_2495);
nor U2619 (N_2619,N_2487,N_2540);
or U2620 (N_2620,N_2498,N_2500);
nand U2621 (N_2621,N_2522,N_2535);
or U2622 (N_2622,N_2485,N_2520);
or U2623 (N_2623,N_2504,N_2538);
xnor U2624 (N_2624,N_2534,N_2487);
xor U2625 (N_2625,N_2618,N_2591);
nor U2626 (N_2626,N_2596,N_2567);
and U2627 (N_2627,N_2572,N_2569);
nand U2628 (N_2628,N_2609,N_2554);
nand U2629 (N_2629,N_2553,N_2555);
or U2630 (N_2630,N_2610,N_2561);
nor U2631 (N_2631,N_2583,N_2563);
or U2632 (N_2632,N_2617,N_2605);
nor U2633 (N_2633,N_2586,N_2623);
nand U2634 (N_2634,N_2620,N_2607);
xor U2635 (N_2635,N_2565,N_2593);
xor U2636 (N_2636,N_2577,N_2589);
and U2637 (N_2637,N_2598,N_2580);
and U2638 (N_2638,N_2611,N_2576);
nor U2639 (N_2639,N_2550,N_2551);
nand U2640 (N_2640,N_2570,N_2579);
nand U2641 (N_2641,N_2571,N_2562);
or U2642 (N_2642,N_2564,N_2574);
nand U2643 (N_2643,N_2614,N_2559);
nor U2644 (N_2644,N_2612,N_2624);
and U2645 (N_2645,N_2557,N_2556);
xor U2646 (N_2646,N_2585,N_2560);
xnor U2647 (N_2647,N_2566,N_2590);
or U2648 (N_2648,N_2599,N_2608);
nor U2649 (N_2649,N_2573,N_2622);
and U2650 (N_2650,N_2584,N_2615);
and U2651 (N_2651,N_2581,N_2594);
nor U2652 (N_2652,N_2582,N_2619);
and U2653 (N_2653,N_2595,N_2616);
nor U2654 (N_2654,N_2597,N_2602);
nand U2655 (N_2655,N_2600,N_2587);
nand U2656 (N_2656,N_2601,N_2603);
nor U2657 (N_2657,N_2568,N_2588);
and U2658 (N_2658,N_2592,N_2606);
nor U2659 (N_2659,N_2604,N_2578);
or U2660 (N_2660,N_2552,N_2621);
or U2661 (N_2661,N_2558,N_2575);
xor U2662 (N_2662,N_2613,N_2609);
or U2663 (N_2663,N_2616,N_2566);
and U2664 (N_2664,N_2605,N_2586);
or U2665 (N_2665,N_2614,N_2578);
nand U2666 (N_2666,N_2552,N_2592);
nand U2667 (N_2667,N_2596,N_2576);
and U2668 (N_2668,N_2578,N_2564);
or U2669 (N_2669,N_2588,N_2620);
or U2670 (N_2670,N_2597,N_2588);
nor U2671 (N_2671,N_2601,N_2590);
nand U2672 (N_2672,N_2580,N_2568);
or U2673 (N_2673,N_2601,N_2552);
nand U2674 (N_2674,N_2560,N_2612);
nor U2675 (N_2675,N_2584,N_2598);
nand U2676 (N_2676,N_2617,N_2567);
xnor U2677 (N_2677,N_2596,N_2571);
nand U2678 (N_2678,N_2624,N_2614);
xnor U2679 (N_2679,N_2568,N_2570);
and U2680 (N_2680,N_2605,N_2589);
or U2681 (N_2681,N_2588,N_2572);
nand U2682 (N_2682,N_2611,N_2582);
nand U2683 (N_2683,N_2575,N_2620);
nand U2684 (N_2684,N_2551,N_2610);
and U2685 (N_2685,N_2611,N_2587);
nand U2686 (N_2686,N_2573,N_2617);
nand U2687 (N_2687,N_2578,N_2569);
or U2688 (N_2688,N_2550,N_2573);
or U2689 (N_2689,N_2565,N_2558);
xor U2690 (N_2690,N_2578,N_2623);
or U2691 (N_2691,N_2567,N_2564);
nor U2692 (N_2692,N_2624,N_2561);
xor U2693 (N_2693,N_2577,N_2553);
and U2694 (N_2694,N_2615,N_2601);
nor U2695 (N_2695,N_2580,N_2595);
and U2696 (N_2696,N_2621,N_2592);
or U2697 (N_2697,N_2594,N_2568);
nand U2698 (N_2698,N_2550,N_2552);
or U2699 (N_2699,N_2559,N_2602);
xor U2700 (N_2700,N_2672,N_2673);
or U2701 (N_2701,N_2671,N_2688);
nand U2702 (N_2702,N_2639,N_2632);
and U2703 (N_2703,N_2656,N_2690);
xor U2704 (N_2704,N_2660,N_2692);
xnor U2705 (N_2705,N_2634,N_2666);
xnor U2706 (N_2706,N_2648,N_2647);
and U2707 (N_2707,N_2662,N_2657);
nor U2708 (N_2708,N_2646,N_2630);
or U2709 (N_2709,N_2637,N_2645);
and U2710 (N_2710,N_2636,N_2653);
and U2711 (N_2711,N_2680,N_2627);
and U2712 (N_2712,N_2644,N_2642);
and U2713 (N_2713,N_2665,N_2663);
xnor U2714 (N_2714,N_2695,N_2674);
nor U2715 (N_2715,N_2628,N_2698);
nand U2716 (N_2716,N_2669,N_2697);
nand U2717 (N_2717,N_2654,N_2689);
nand U2718 (N_2718,N_2641,N_2678);
or U2719 (N_2719,N_2661,N_2691);
nand U2720 (N_2720,N_2635,N_2650);
nand U2721 (N_2721,N_2658,N_2643);
nor U2722 (N_2722,N_2640,N_2686);
nor U2723 (N_2723,N_2676,N_2696);
and U2724 (N_2724,N_2687,N_2699);
nor U2725 (N_2725,N_2693,N_2677);
and U2726 (N_2726,N_2670,N_2649);
and U2727 (N_2727,N_2638,N_2655);
xnor U2728 (N_2728,N_2681,N_2625);
xnor U2729 (N_2729,N_2679,N_2684);
nand U2730 (N_2730,N_2651,N_2659);
nor U2731 (N_2731,N_2631,N_2626);
xnor U2732 (N_2732,N_2682,N_2683);
nand U2733 (N_2733,N_2633,N_2629);
nand U2734 (N_2734,N_2675,N_2664);
nand U2735 (N_2735,N_2685,N_2667);
nor U2736 (N_2736,N_2668,N_2652);
or U2737 (N_2737,N_2694,N_2685);
xnor U2738 (N_2738,N_2658,N_2664);
or U2739 (N_2739,N_2638,N_2660);
and U2740 (N_2740,N_2666,N_2645);
nor U2741 (N_2741,N_2680,N_2660);
nand U2742 (N_2742,N_2684,N_2665);
and U2743 (N_2743,N_2644,N_2662);
xnor U2744 (N_2744,N_2673,N_2643);
and U2745 (N_2745,N_2693,N_2678);
and U2746 (N_2746,N_2637,N_2659);
or U2747 (N_2747,N_2640,N_2641);
nand U2748 (N_2748,N_2628,N_2658);
xor U2749 (N_2749,N_2682,N_2644);
and U2750 (N_2750,N_2665,N_2673);
xnor U2751 (N_2751,N_2655,N_2627);
nand U2752 (N_2752,N_2694,N_2671);
xnor U2753 (N_2753,N_2643,N_2663);
nand U2754 (N_2754,N_2626,N_2647);
nand U2755 (N_2755,N_2656,N_2635);
and U2756 (N_2756,N_2675,N_2649);
xor U2757 (N_2757,N_2685,N_2656);
or U2758 (N_2758,N_2662,N_2625);
and U2759 (N_2759,N_2647,N_2634);
nor U2760 (N_2760,N_2670,N_2656);
nand U2761 (N_2761,N_2672,N_2681);
nand U2762 (N_2762,N_2625,N_2673);
xnor U2763 (N_2763,N_2681,N_2674);
nor U2764 (N_2764,N_2649,N_2644);
xnor U2765 (N_2765,N_2626,N_2637);
or U2766 (N_2766,N_2631,N_2650);
nor U2767 (N_2767,N_2643,N_2692);
xor U2768 (N_2768,N_2689,N_2627);
xnor U2769 (N_2769,N_2693,N_2630);
or U2770 (N_2770,N_2665,N_2626);
nand U2771 (N_2771,N_2629,N_2674);
nand U2772 (N_2772,N_2698,N_2692);
nand U2773 (N_2773,N_2687,N_2659);
nand U2774 (N_2774,N_2636,N_2638);
or U2775 (N_2775,N_2760,N_2751);
nor U2776 (N_2776,N_2723,N_2706);
or U2777 (N_2777,N_2716,N_2737);
or U2778 (N_2778,N_2712,N_2718);
nand U2779 (N_2779,N_2729,N_2709);
or U2780 (N_2780,N_2711,N_2728);
nand U2781 (N_2781,N_2717,N_2774);
or U2782 (N_2782,N_2773,N_2771);
nor U2783 (N_2783,N_2710,N_2741);
or U2784 (N_2784,N_2765,N_2707);
and U2785 (N_2785,N_2713,N_2750);
nand U2786 (N_2786,N_2727,N_2744);
xnor U2787 (N_2787,N_2752,N_2767);
xor U2788 (N_2788,N_2735,N_2768);
nand U2789 (N_2789,N_2734,N_2701);
xor U2790 (N_2790,N_2738,N_2740);
and U2791 (N_2791,N_2721,N_2722);
nand U2792 (N_2792,N_2766,N_2720);
nand U2793 (N_2793,N_2754,N_2748);
and U2794 (N_2794,N_2747,N_2769);
nor U2795 (N_2795,N_2762,N_2733);
nor U2796 (N_2796,N_2763,N_2724);
nand U2797 (N_2797,N_2705,N_2731);
or U2798 (N_2798,N_2753,N_2702);
and U2799 (N_2799,N_2758,N_2755);
nand U2800 (N_2800,N_2719,N_2714);
and U2801 (N_2801,N_2715,N_2730);
nor U2802 (N_2802,N_2742,N_2739);
nor U2803 (N_2803,N_2757,N_2708);
nand U2804 (N_2804,N_2745,N_2759);
xor U2805 (N_2805,N_2736,N_2732);
or U2806 (N_2806,N_2700,N_2761);
xor U2807 (N_2807,N_2772,N_2749);
or U2808 (N_2808,N_2704,N_2726);
xnor U2809 (N_2809,N_2746,N_2756);
or U2810 (N_2810,N_2725,N_2743);
nor U2811 (N_2811,N_2770,N_2764);
nor U2812 (N_2812,N_2703,N_2724);
nand U2813 (N_2813,N_2705,N_2735);
and U2814 (N_2814,N_2763,N_2753);
and U2815 (N_2815,N_2711,N_2720);
xor U2816 (N_2816,N_2727,N_2702);
or U2817 (N_2817,N_2732,N_2752);
or U2818 (N_2818,N_2725,N_2704);
or U2819 (N_2819,N_2708,N_2717);
nand U2820 (N_2820,N_2761,N_2734);
and U2821 (N_2821,N_2721,N_2704);
or U2822 (N_2822,N_2773,N_2769);
xor U2823 (N_2823,N_2704,N_2736);
and U2824 (N_2824,N_2714,N_2726);
nand U2825 (N_2825,N_2766,N_2711);
and U2826 (N_2826,N_2724,N_2755);
and U2827 (N_2827,N_2720,N_2732);
nand U2828 (N_2828,N_2702,N_2741);
nor U2829 (N_2829,N_2722,N_2766);
or U2830 (N_2830,N_2727,N_2724);
nand U2831 (N_2831,N_2727,N_2759);
or U2832 (N_2832,N_2741,N_2719);
and U2833 (N_2833,N_2755,N_2716);
nor U2834 (N_2834,N_2752,N_2736);
xor U2835 (N_2835,N_2700,N_2720);
or U2836 (N_2836,N_2709,N_2724);
nand U2837 (N_2837,N_2707,N_2757);
nand U2838 (N_2838,N_2739,N_2741);
xor U2839 (N_2839,N_2771,N_2746);
nand U2840 (N_2840,N_2768,N_2706);
or U2841 (N_2841,N_2758,N_2761);
nor U2842 (N_2842,N_2739,N_2704);
nand U2843 (N_2843,N_2706,N_2739);
or U2844 (N_2844,N_2738,N_2747);
or U2845 (N_2845,N_2733,N_2757);
nor U2846 (N_2846,N_2725,N_2711);
nand U2847 (N_2847,N_2706,N_2728);
nand U2848 (N_2848,N_2726,N_2709);
or U2849 (N_2849,N_2743,N_2769);
nand U2850 (N_2850,N_2831,N_2799);
nor U2851 (N_2851,N_2829,N_2794);
and U2852 (N_2852,N_2798,N_2779);
or U2853 (N_2853,N_2791,N_2834);
nand U2854 (N_2854,N_2817,N_2807);
nand U2855 (N_2855,N_2827,N_2825);
and U2856 (N_2856,N_2836,N_2804);
and U2857 (N_2857,N_2823,N_2805);
xnor U2858 (N_2858,N_2782,N_2821);
and U2859 (N_2859,N_2810,N_2833);
nor U2860 (N_2860,N_2842,N_2837);
or U2861 (N_2861,N_2838,N_2835);
nand U2862 (N_2862,N_2832,N_2822);
xor U2863 (N_2863,N_2813,N_2806);
or U2864 (N_2864,N_2784,N_2777);
nand U2865 (N_2865,N_2783,N_2819);
nand U2866 (N_2866,N_2796,N_2846);
nor U2867 (N_2867,N_2788,N_2785);
and U2868 (N_2868,N_2786,N_2790);
nand U2869 (N_2869,N_2820,N_2808);
xnor U2870 (N_2870,N_2811,N_2839);
or U2871 (N_2871,N_2775,N_2793);
and U2872 (N_2872,N_2776,N_2795);
nor U2873 (N_2873,N_2841,N_2800);
or U2874 (N_2874,N_2792,N_2789);
or U2875 (N_2875,N_2826,N_2848);
nand U2876 (N_2876,N_2816,N_2840);
or U2877 (N_2877,N_2849,N_2780);
nand U2878 (N_2878,N_2781,N_2802);
and U2879 (N_2879,N_2843,N_2814);
or U2880 (N_2880,N_2830,N_2818);
and U2881 (N_2881,N_2801,N_2845);
or U2882 (N_2882,N_2812,N_2797);
or U2883 (N_2883,N_2824,N_2815);
or U2884 (N_2884,N_2787,N_2844);
and U2885 (N_2885,N_2828,N_2847);
or U2886 (N_2886,N_2778,N_2803);
or U2887 (N_2887,N_2809,N_2780);
or U2888 (N_2888,N_2794,N_2847);
xnor U2889 (N_2889,N_2776,N_2813);
xnor U2890 (N_2890,N_2830,N_2820);
or U2891 (N_2891,N_2842,N_2834);
or U2892 (N_2892,N_2791,N_2845);
nand U2893 (N_2893,N_2829,N_2811);
nand U2894 (N_2894,N_2849,N_2796);
and U2895 (N_2895,N_2825,N_2812);
xor U2896 (N_2896,N_2814,N_2815);
or U2897 (N_2897,N_2796,N_2800);
and U2898 (N_2898,N_2811,N_2815);
xnor U2899 (N_2899,N_2783,N_2789);
xnor U2900 (N_2900,N_2842,N_2824);
xnor U2901 (N_2901,N_2847,N_2800);
xor U2902 (N_2902,N_2830,N_2823);
nand U2903 (N_2903,N_2784,N_2825);
xor U2904 (N_2904,N_2845,N_2784);
nor U2905 (N_2905,N_2848,N_2824);
nor U2906 (N_2906,N_2784,N_2848);
nor U2907 (N_2907,N_2840,N_2785);
xnor U2908 (N_2908,N_2791,N_2795);
nand U2909 (N_2909,N_2823,N_2778);
nand U2910 (N_2910,N_2787,N_2782);
and U2911 (N_2911,N_2818,N_2782);
xor U2912 (N_2912,N_2810,N_2799);
nand U2913 (N_2913,N_2776,N_2843);
nand U2914 (N_2914,N_2811,N_2828);
nor U2915 (N_2915,N_2833,N_2838);
xnor U2916 (N_2916,N_2805,N_2780);
nand U2917 (N_2917,N_2787,N_2812);
nor U2918 (N_2918,N_2809,N_2824);
nand U2919 (N_2919,N_2809,N_2839);
nor U2920 (N_2920,N_2819,N_2844);
xnor U2921 (N_2921,N_2825,N_2778);
nand U2922 (N_2922,N_2803,N_2808);
and U2923 (N_2923,N_2848,N_2841);
and U2924 (N_2924,N_2802,N_2805);
or U2925 (N_2925,N_2884,N_2895);
or U2926 (N_2926,N_2853,N_2909);
nand U2927 (N_2927,N_2887,N_2919);
nand U2928 (N_2928,N_2923,N_2879);
and U2929 (N_2929,N_2903,N_2918);
or U2930 (N_2930,N_2861,N_2898);
xor U2931 (N_2931,N_2872,N_2873);
and U2932 (N_2932,N_2857,N_2920);
xor U2933 (N_2933,N_2875,N_2902);
nor U2934 (N_2934,N_2899,N_2888);
and U2935 (N_2935,N_2868,N_2914);
or U2936 (N_2936,N_2915,N_2892);
nor U2937 (N_2937,N_2878,N_2854);
nor U2938 (N_2938,N_2865,N_2912);
xnor U2939 (N_2939,N_2871,N_2863);
xor U2940 (N_2940,N_2907,N_2864);
and U2941 (N_2941,N_2867,N_2883);
nor U2942 (N_2942,N_2910,N_2881);
xnor U2943 (N_2943,N_2877,N_2901);
nor U2944 (N_2944,N_2869,N_2924);
xor U2945 (N_2945,N_2890,N_2860);
and U2946 (N_2946,N_2855,N_2891);
nand U2947 (N_2947,N_2850,N_2880);
or U2948 (N_2948,N_2852,N_2858);
nor U2949 (N_2949,N_2913,N_2905);
xnor U2950 (N_2950,N_2904,N_2900);
or U2951 (N_2951,N_2876,N_2851);
or U2952 (N_2952,N_2859,N_2911);
nand U2953 (N_2953,N_2896,N_2874);
and U2954 (N_2954,N_2886,N_2897);
nand U2955 (N_2955,N_2870,N_2908);
nand U2956 (N_2956,N_2882,N_2922);
nand U2957 (N_2957,N_2893,N_2866);
xnor U2958 (N_2958,N_2921,N_2894);
xor U2959 (N_2959,N_2906,N_2862);
nor U2960 (N_2960,N_2917,N_2856);
nand U2961 (N_2961,N_2885,N_2916);
and U2962 (N_2962,N_2889,N_2885);
nand U2963 (N_2963,N_2888,N_2920);
nand U2964 (N_2964,N_2903,N_2869);
or U2965 (N_2965,N_2922,N_2902);
xor U2966 (N_2966,N_2883,N_2871);
and U2967 (N_2967,N_2859,N_2885);
xor U2968 (N_2968,N_2863,N_2869);
and U2969 (N_2969,N_2883,N_2856);
xor U2970 (N_2970,N_2908,N_2854);
and U2971 (N_2971,N_2855,N_2921);
xnor U2972 (N_2972,N_2891,N_2861);
or U2973 (N_2973,N_2881,N_2908);
and U2974 (N_2974,N_2883,N_2909);
xnor U2975 (N_2975,N_2894,N_2891);
xnor U2976 (N_2976,N_2895,N_2918);
nor U2977 (N_2977,N_2879,N_2884);
nand U2978 (N_2978,N_2920,N_2872);
nand U2979 (N_2979,N_2898,N_2875);
and U2980 (N_2980,N_2909,N_2857);
or U2981 (N_2981,N_2851,N_2864);
nand U2982 (N_2982,N_2907,N_2885);
nand U2983 (N_2983,N_2882,N_2897);
nor U2984 (N_2984,N_2890,N_2888);
and U2985 (N_2985,N_2883,N_2910);
or U2986 (N_2986,N_2917,N_2915);
and U2987 (N_2987,N_2883,N_2884);
nand U2988 (N_2988,N_2871,N_2924);
and U2989 (N_2989,N_2879,N_2861);
and U2990 (N_2990,N_2883,N_2902);
and U2991 (N_2991,N_2898,N_2892);
or U2992 (N_2992,N_2901,N_2900);
nand U2993 (N_2993,N_2854,N_2890);
nor U2994 (N_2994,N_2891,N_2919);
and U2995 (N_2995,N_2897,N_2893);
nand U2996 (N_2996,N_2921,N_2853);
and U2997 (N_2997,N_2861,N_2866);
xnor U2998 (N_2998,N_2893,N_2917);
xnor U2999 (N_2999,N_2923,N_2854);
xnor UO_0 (O_0,N_2938,N_2953);
nand UO_1 (O_1,N_2925,N_2980);
and UO_2 (O_2,N_2949,N_2967);
nand UO_3 (O_3,N_2935,N_2978);
and UO_4 (O_4,N_2960,N_2997);
or UO_5 (O_5,N_2990,N_2957);
nor UO_6 (O_6,N_2998,N_2955);
nor UO_7 (O_7,N_2965,N_2940);
or UO_8 (O_8,N_2985,N_2977);
nor UO_9 (O_9,N_2968,N_2993);
or UO_10 (O_10,N_2975,N_2976);
nand UO_11 (O_11,N_2926,N_2927);
xnor UO_12 (O_12,N_2928,N_2966);
or UO_13 (O_13,N_2937,N_2987);
nand UO_14 (O_14,N_2972,N_2943);
nor UO_15 (O_15,N_2954,N_2979);
or UO_16 (O_16,N_2946,N_2989);
xnor UO_17 (O_17,N_2931,N_2951);
and UO_18 (O_18,N_2950,N_2983);
xnor UO_19 (O_19,N_2994,N_2934);
nor UO_20 (O_20,N_2974,N_2986);
and UO_21 (O_21,N_2991,N_2947);
or UO_22 (O_22,N_2982,N_2933);
nand UO_23 (O_23,N_2952,N_2996);
xnor UO_24 (O_24,N_2930,N_2948);
xor UO_25 (O_25,N_2973,N_2995);
xnor UO_26 (O_26,N_2988,N_2971);
and UO_27 (O_27,N_2944,N_2939);
nor UO_28 (O_28,N_2964,N_2959);
or UO_29 (O_29,N_2958,N_2969);
nor UO_30 (O_30,N_2932,N_2956);
and UO_31 (O_31,N_2941,N_2942);
nor UO_32 (O_32,N_2962,N_2970);
and UO_33 (O_33,N_2984,N_2992);
nor UO_34 (O_34,N_2961,N_2963);
xnor UO_35 (O_35,N_2981,N_2929);
xnor UO_36 (O_36,N_2945,N_2999);
and UO_37 (O_37,N_2936,N_2927);
or UO_38 (O_38,N_2938,N_2959);
nand UO_39 (O_39,N_2941,N_2979);
and UO_40 (O_40,N_2935,N_2934);
nor UO_41 (O_41,N_2978,N_2993);
xor UO_42 (O_42,N_2993,N_2952);
nand UO_43 (O_43,N_2944,N_2930);
nand UO_44 (O_44,N_2962,N_2965);
nor UO_45 (O_45,N_2979,N_2986);
nand UO_46 (O_46,N_2951,N_2957);
xor UO_47 (O_47,N_2930,N_2929);
nor UO_48 (O_48,N_2992,N_2999);
nor UO_49 (O_49,N_2976,N_2926);
xnor UO_50 (O_50,N_2978,N_2946);
and UO_51 (O_51,N_2958,N_2929);
nand UO_52 (O_52,N_2942,N_2933);
xnor UO_53 (O_53,N_2976,N_2977);
nand UO_54 (O_54,N_2948,N_2958);
xnor UO_55 (O_55,N_2947,N_2989);
and UO_56 (O_56,N_2944,N_2959);
nor UO_57 (O_57,N_2940,N_2959);
nand UO_58 (O_58,N_2972,N_2967);
xor UO_59 (O_59,N_2932,N_2995);
or UO_60 (O_60,N_2983,N_2970);
nor UO_61 (O_61,N_2942,N_2949);
xnor UO_62 (O_62,N_2954,N_2953);
nand UO_63 (O_63,N_2982,N_2948);
nor UO_64 (O_64,N_2987,N_2945);
xor UO_65 (O_65,N_2960,N_2988);
xnor UO_66 (O_66,N_2968,N_2965);
and UO_67 (O_67,N_2937,N_2934);
and UO_68 (O_68,N_2926,N_2989);
or UO_69 (O_69,N_2939,N_2928);
xor UO_70 (O_70,N_2926,N_2936);
nand UO_71 (O_71,N_2949,N_2966);
nand UO_72 (O_72,N_2967,N_2993);
or UO_73 (O_73,N_2955,N_2994);
and UO_74 (O_74,N_2998,N_2975);
and UO_75 (O_75,N_2974,N_2995);
and UO_76 (O_76,N_2957,N_2938);
and UO_77 (O_77,N_2928,N_2935);
and UO_78 (O_78,N_2956,N_2985);
or UO_79 (O_79,N_2976,N_2995);
xor UO_80 (O_80,N_2979,N_2973);
nand UO_81 (O_81,N_2958,N_2960);
nor UO_82 (O_82,N_2947,N_2968);
xnor UO_83 (O_83,N_2999,N_2976);
nand UO_84 (O_84,N_2992,N_2942);
xnor UO_85 (O_85,N_2945,N_2954);
or UO_86 (O_86,N_2949,N_2946);
nor UO_87 (O_87,N_2986,N_2939);
nand UO_88 (O_88,N_2937,N_2941);
xor UO_89 (O_89,N_2980,N_2941);
and UO_90 (O_90,N_2992,N_2966);
xnor UO_91 (O_91,N_2973,N_2992);
or UO_92 (O_92,N_2949,N_2979);
xnor UO_93 (O_93,N_2952,N_2965);
nand UO_94 (O_94,N_2998,N_2963);
xnor UO_95 (O_95,N_2931,N_2964);
and UO_96 (O_96,N_2967,N_2929);
xor UO_97 (O_97,N_2970,N_2999);
nand UO_98 (O_98,N_2936,N_2949);
xnor UO_99 (O_99,N_2948,N_2954);
xor UO_100 (O_100,N_2976,N_2925);
nand UO_101 (O_101,N_2990,N_2931);
nand UO_102 (O_102,N_2990,N_2967);
and UO_103 (O_103,N_2941,N_2932);
nand UO_104 (O_104,N_2999,N_2989);
nand UO_105 (O_105,N_2968,N_2982);
nand UO_106 (O_106,N_2980,N_2959);
or UO_107 (O_107,N_2976,N_2953);
nor UO_108 (O_108,N_2952,N_2942);
nor UO_109 (O_109,N_2951,N_2953);
and UO_110 (O_110,N_2973,N_2942);
nand UO_111 (O_111,N_2958,N_2993);
or UO_112 (O_112,N_2992,N_2944);
nor UO_113 (O_113,N_2998,N_2992);
nand UO_114 (O_114,N_2937,N_2958);
or UO_115 (O_115,N_2931,N_2970);
nand UO_116 (O_116,N_2954,N_2987);
nor UO_117 (O_117,N_2950,N_2963);
or UO_118 (O_118,N_2947,N_2956);
or UO_119 (O_119,N_2952,N_2957);
and UO_120 (O_120,N_2977,N_2936);
or UO_121 (O_121,N_2965,N_2992);
nand UO_122 (O_122,N_2999,N_2955);
nand UO_123 (O_123,N_2925,N_2935);
nand UO_124 (O_124,N_2997,N_2926);
xor UO_125 (O_125,N_2967,N_2994);
and UO_126 (O_126,N_2996,N_2990);
nor UO_127 (O_127,N_2935,N_2937);
nand UO_128 (O_128,N_2999,N_2925);
xor UO_129 (O_129,N_2945,N_2990);
xnor UO_130 (O_130,N_2952,N_2937);
nor UO_131 (O_131,N_2934,N_2986);
nand UO_132 (O_132,N_2964,N_2948);
and UO_133 (O_133,N_2928,N_2948);
and UO_134 (O_134,N_2971,N_2945);
xnor UO_135 (O_135,N_2932,N_2982);
xnor UO_136 (O_136,N_2978,N_2953);
nor UO_137 (O_137,N_2961,N_2935);
and UO_138 (O_138,N_2959,N_2931);
or UO_139 (O_139,N_2946,N_2944);
xor UO_140 (O_140,N_2986,N_2993);
xnor UO_141 (O_141,N_2978,N_2945);
or UO_142 (O_142,N_2949,N_2947);
nand UO_143 (O_143,N_2966,N_2994);
nor UO_144 (O_144,N_2954,N_2968);
and UO_145 (O_145,N_2964,N_2984);
nor UO_146 (O_146,N_2961,N_2959);
or UO_147 (O_147,N_2963,N_2942);
nand UO_148 (O_148,N_2989,N_2984);
nor UO_149 (O_149,N_2927,N_2963);
or UO_150 (O_150,N_2983,N_2949);
nor UO_151 (O_151,N_2948,N_2981);
nor UO_152 (O_152,N_2935,N_2939);
or UO_153 (O_153,N_2950,N_2932);
nor UO_154 (O_154,N_2960,N_2955);
or UO_155 (O_155,N_2947,N_2996);
nor UO_156 (O_156,N_2987,N_2992);
or UO_157 (O_157,N_2930,N_2987);
or UO_158 (O_158,N_2932,N_2955);
or UO_159 (O_159,N_2994,N_2948);
or UO_160 (O_160,N_2984,N_2929);
xor UO_161 (O_161,N_2947,N_2999);
or UO_162 (O_162,N_2927,N_2948);
nand UO_163 (O_163,N_2932,N_2928);
and UO_164 (O_164,N_2960,N_2982);
or UO_165 (O_165,N_2970,N_2975);
xnor UO_166 (O_166,N_2970,N_2950);
or UO_167 (O_167,N_2987,N_2983);
nand UO_168 (O_168,N_2938,N_2961);
or UO_169 (O_169,N_2943,N_2995);
nand UO_170 (O_170,N_2999,N_2938);
xor UO_171 (O_171,N_2966,N_2967);
and UO_172 (O_172,N_2988,N_2997);
or UO_173 (O_173,N_2968,N_2952);
xnor UO_174 (O_174,N_2984,N_2949);
nor UO_175 (O_175,N_2972,N_2999);
nor UO_176 (O_176,N_2968,N_2974);
nand UO_177 (O_177,N_2940,N_2980);
xor UO_178 (O_178,N_2927,N_2994);
nand UO_179 (O_179,N_2964,N_2928);
or UO_180 (O_180,N_2948,N_2952);
and UO_181 (O_181,N_2951,N_2991);
nand UO_182 (O_182,N_2990,N_2972);
and UO_183 (O_183,N_2972,N_2977);
xnor UO_184 (O_184,N_2950,N_2994);
and UO_185 (O_185,N_2995,N_2941);
nand UO_186 (O_186,N_2988,N_2952);
or UO_187 (O_187,N_2967,N_2933);
nor UO_188 (O_188,N_2930,N_2979);
and UO_189 (O_189,N_2937,N_2991);
and UO_190 (O_190,N_2997,N_2928);
or UO_191 (O_191,N_2927,N_2997);
and UO_192 (O_192,N_2956,N_2966);
and UO_193 (O_193,N_2990,N_2981);
and UO_194 (O_194,N_2994,N_2951);
or UO_195 (O_195,N_2962,N_2978);
or UO_196 (O_196,N_2928,N_2944);
and UO_197 (O_197,N_2950,N_2973);
and UO_198 (O_198,N_2933,N_2985);
nor UO_199 (O_199,N_2985,N_2928);
xor UO_200 (O_200,N_2940,N_2956);
nor UO_201 (O_201,N_2968,N_2977);
and UO_202 (O_202,N_2946,N_2977);
nand UO_203 (O_203,N_2999,N_2964);
and UO_204 (O_204,N_2981,N_2955);
xor UO_205 (O_205,N_2998,N_2970);
or UO_206 (O_206,N_2966,N_2981);
xor UO_207 (O_207,N_2992,N_2983);
nand UO_208 (O_208,N_2975,N_2979);
nand UO_209 (O_209,N_2950,N_2941);
and UO_210 (O_210,N_2928,N_2976);
or UO_211 (O_211,N_2994,N_2938);
nand UO_212 (O_212,N_2933,N_2958);
xor UO_213 (O_213,N_2980,N_2989);
or UO_214 (O_214,N_2988,N_2970);
or UO_215 (O_215,N_2977,N_2995);
xnor UO_216 (O_216,N_2940,N_2978);
xor UO_217 (O_217,N_2927,N_2953);
nor UO_218 (O_218,N_2937,N_2972);
xor UO_219 (O_219,N_2933,N_2949);
or UO_220 (O_220,N_2990,N_2936);
and UO_221 (O_221,N_2977,N_2987);
xnor UO_222 (O_222,N_2960,N_2953);
nor UO_223 (O_223,N_2936,N_2995);
or UO_224 (O_224,N_2967,N_2975);
xor UO_225 (O_225,N_2992,N_2935);
and UO_226 (O_226,N_2952,N_2955);
nor UO_227 (O_227,N_2973,N_2983);
and UO_228 (O_228,N_2988,N_2995);
or UO_229 (O_229,N_2941,N_2933);
and UO_230 (O_230,N_2997,N_2983);
nor UO_231 (O_231,N_2972,N_2976);
nor UO_232 (O_232,N_2943,N_2935);
nor UO_233 (O_233,N_2994,N_2969);
and UO_234 (O_234,N_2964,N_2978);
nand UO_235 (O_235,N_2981,N_2935);
or UO_236 (O_236,N_2943,N_2986);
nor UO_237 (O_237,N_2932,N_2946);
nand UO_238 (O_238,N_2933,N_2961);
nand UO_239 (O_239,N_2993,N_2964);
nand UO_240 (O_240,N_2935,N_2964);
or UO_241 (O_241,N_2970,N_2948);
or UO_242 (O_242,N_2962,N_2981);
nor UO_243 (O_243,N_2988,N_2990);
xnor UO_244 (O_244,N_2970,N_2954);
nand UO_245 (O_245,N_2962,N_2960);
or UO_246 (O_246,N_2945,N_2929);
xor UO_247 (O_247,N_2943,N_2953);
and UO_248 (O_248,N_2985,N_2975);
nand UO_249 (O_249,N_2930,N_2958);
xor UO_250 (O_250,N_2975,N_2993);
or UO_251 (O_251,N_2961,N_2988);
nor UO_252 (O_252,N_2940,N_2957);
xnor UO_253 (O_253,N_2932,N_2952);
or UO_254 (O_254,N_2994,N_2932);
nor UO_255 (O_255,N_2932,N_2972);
nand UO_256 (O_256,N_2938,N_2926);
nand UO_257 (O_257,N_2964,N_2953);
xor UO_258 (O_258,N_2963,N_2933);
or UO_259 (O_259,N_2974,N_2984);
nand UO_260 (O_260,N_2975,N_2978);
and UO_261 (O_261,N_2937,N_2940);
nor UO_262 (O_262,N_2930,N_2947);
and UO_263 (O_263,N_2925,N_2993);
or UO_264 (O_264,N_2974,N_2946);
nand UO_265 (O_265,N_2959,N_2953);
xor UO_266 (O_266,N_2931,N_2995);
nor UO_267 (O_267,N_2945,N_2957);
nor UO_268 (O_268,N_2994,N_2928);
nor UO_269 (O_269,N_2991,N_2989);
or UO_270 (O_270,N_2939,N_2977);
nor UO_271 (O_271,N_2972,N_2992);
and UO_272 (O_272,N_2970,N_2951);
or UO_273 (O_273,N_2995,N_2938);
and UO_274 (O_274,N_2936,N_2971);
and UO_275 (O_275,N_2953,N_2961);
nand UO_276 (O_276,N_2984,N_2930);
or UO_277 (O_277,N_2985,N_2941);
and UO_278 (O_278,N_2926,N_2932);
or UO_279 (O_279,N_2993,N_2985);
nand UO_280 (O_280,N_2931,N_2940);
or UO_281 (O_281,N_2962,N_2940);
and UO_282 (O_282,N_2939,N_2955);
nand UO_283 (O_283,N_2948,N_2942);
and UO_284 (O_284,N_2927,N_2988);
or UO_285 (O_285,N_2934,N_2991);
and UO_286 (O_286,N_2958,N_2978);
or UO_287 (O_287,N_2996,N_2975);
nor UO_288 (O_288,N_2935,N_2976);
nand UO_289 (O_289,N_2993,N_2942);
or UO_290 (O_290,N_2967,N_2970);
nand UO_291 (O_291,N_2992,N_2929);
xnor UO_292 (O_292,N_2970,N_2949);
nand UO_293 (O_293,N_2950,N_2933);
and UO_294 (O_294,N_2942,N_2980);
nor UO_295 (O_295,N_2951,N_2984);
xnor UO_296 (O_296,N_2950,N_2961);
nand UO_297 (O_297,N_2984,N_2973);
xor UO_298 (O_298,N_2940,N_2971);
nand UO_299 (O_299,N_2973,N_2998);
nand UO_300 (O_300,N_2998,N_2933);
xor UO_301 (O_301,N_2957,N_2937);
nor UO_302 (O_302,N_2935,N_2971);
nand UO_303 (O_303,N_2977,N_2996);
nand UO_304 (O_304,N_2998,N_2943);
xor UO_305 (O_305,N_2927,N_2969);
nor UO_306 (O_306,N_2973,N_2940);
nor UO_307 (O_307,N_2965,N_2931);
and UO_308 (O_308,N_2963,N_2978);
xor UO_309 (O_309,N_2959,N_2930);
nor UO_310 (O_310,N_2945,N_2996);
nand UO_311 (O_311,N_2931,N_2950);
xor UO_312 (O_312,N_2976,N_2959);
and UO_313 (O_313,N_2930,N_2952);
nand UO_314 (O_314,N_2929,N_2988);
nor UO_315 (O_315,N_2982,N_2941);
or UO_316 (O_316,N_2997,N_2961);
or UO_317 (O_317,N_2983,N_2959);
nand UO_318 (O_318,N_2960,N_2974);
and UO_319 (O_319,N_2940,N_2926);
xnor UO_320 (O_320,N_2962,N_2983);
or UO_321 (O_321,N_2997,N_2929);
and UO_322 (O_322,N_2991,N_2994);
nor UO_323 (O_323,N_2983,N_2934);
nand UO_324 (O_324,N_2964,N_2996);
or UO_325 (O_325,N_2949,N_2943);
nor UO_326 (O_326,N_2956,N_2943);
nand UO_327 (O_327,N_2950,N_2996);
nor UO_328 (O_328,N_2933,N_2953);
or UO_329 (O_329,N_2943,N_2991);
or UO_330 (O_330,N_2942,N_2989);
and UO_331 (O_331,N_2931,N_2979);
xor UO_332 (O_332,N_2949,N_2973);
nor UO_333 (O_333,N_2974,N_2989);
xnor UO_334 (O_334,N_2961,N_2952);
or UO_335 (O_335,N_2998,N_2934);
or UO_336 (O_336,N_2990,N_2994);
and UO_337 (O_337,N_2995,N_2928);
nand UO_338 (O_338,N_2932,N_2951);
and UO_339 (O_339,N_2984,N_2969);
nor UO_340 (O_340,N_2990,N_2987);
nor UO_341 (O_341,N_2960,N_2971);
nor UO_342 (O_342,N_2932,N_2967);
nand UO_343 (O_343,N_2936,N_2960);
nand UO_344 (O_344,N_2962,N_2997);
and UO_345 (O_345,N_2948,N_2940);
xnor UO_346 (O_346,N_2985,N_2995);
or UO_347 (O_347,N_2944,N_2998);
or UO_348 (O_348,N_2997,N_2999);
and UO_349 (O_349,N_2961,N_2965);
nand UO_350 (O_350,N_2943,N_2942);
or UO_351 (O_351,N_2967,N_2969);
or UO_352 (O_352,N_2989,N_2979);
nor UO_353 (O_353,N_2942,N_2931);
nor UO_354 (O_354,N_2970,N_2981);
or UO_355 (O_355,N_2982,N_2936);
and UO_356 (O_356,N_2945,N_2931);
and UO_357 (O_357,N_2991,N_2995);
or UO_358 (O_358,N_2996,N_2959);
or UO_359 (O_359,N_2977,N_2935);
nor UO_360 (O_360,N_2926,N_2977);
or UO_361 (O_361,N_2952,N_2989);
and UO_362 (O_362,N_2935,N_2948);
or UO_363 (O_363,N_2956,N_2964);
nand UO_364 (O_364,N_2937,N_2948);
and UO_365 (O_365,N_2989,N_2957);
nand UO_366 (O_366,N_2930,N_2964);
xor UO_367 (O_367,N_2952,N_2994);
nor UO_368 (O_368,N_2997,N_2976);
or UO_369 (O_369,N_2971,N_2947);
nand UO_370 (O_370,N_2994,N_2972);
or UO_371 (O_371,N_2973,N_2987);
nand UO_372 (O_372,N_2950,N_2945);
xnor UO_373 (O_373,N_2957,N_2996);
xnor UO_374 (O_374,N_2939,N_2965);
xor UO_375 (O_375,N_2954,N_2955);
nand UO_376 (O_376,N_2948,N_2941);
nand UO_377 (O_377,N_2976,N_2978);
nor UO_378 (O_378,N_2975,N_2926);
or UO_379 (O_379,N_2998,N_2939);
nor UO_380 (O_380,N_2987,N_2947);
and UO_381 (O_381,N_2935,N_2959);
nor UO_382 (O_382,N_2964,N_2927);
xnor UO_383 (O_383,N_2971,N_2999);
nand UO_384 (O_384,N_2936,N_2930);
xor UO_385 (O_385,N_2942,N_2979);
or UO_386 (O_386,N_2978,N_2933);
nor UO_387 (O_387,N_2990,N_2929);
nand UO_388 (O_388,N_2989,N_2997);
nor UO_389 (O_389,N_2934,N_2931);
nand UO_390 (O_390,N_2956,N_2953);
xor UO_391 (O_391,N_2988,N_2938);
nand UO_392 (O_392,N_2993,N_2933);
xnor UO_393 (O_393,N_2959,N_2945);
nor UO_394 (O_394,N_2975,N_2952);
nor UO_395 (O_395,N_2997,N_2944);
or UO_396 (O_396,N_2928,N_2992);
nor UO_397 (O_397,N_2931,N_2960);
or UO_398 (O_398,N_2961,N_2991);
nand UO_399 (O_399,N_2986,N_2961);
or UO_400 (O_400,N_2975,N_2950);
and UO_401 (O_401,N_2991,N_2930);
and UO_402 (O_402,N_2995,N_2997);
and UO_403 (O_403,N_2950,N_2955);
xor UO_404 (O_404,N_2973,N_2946);
nor UO_405 (O_405,N_2966,N_2926);
nor UO_406 (O_406,N_2971,N_2980);
nor UO_407 (O_407,N_2952,N_2969);
nor UO_408 (O_408,N_2954,N_2964);
or UO_409 (O_409,N_2937,N_2980);
nor UO_410 (O_410,N_2974,N_2990);
nor UO_411 (O_411,N_2933,N_2931);
nor UO_412 (O_412,N_2959,N_2973);
nand UO_413 (O_413,N_2962,N_2944);
and UO_414 (O_414,N_2974,N_2926);
xor UO_415 (O_415,N_2996,N_2978);
nor UO_416 (O_416,N_2959,N_2971);
nor UO_417 (O_417,N_2943,N_2961);
nor UO_418 (O_418,N_2935,N_2973);
nor UO_419 (O_419,N_2982,N_2980);
or UO_420 (O_420,N_2955,N_2951);
or UO_421 (O_421,N_2940,N_2974);
or UO_422 (O_422,N_2933,N_2946);
xnor UO_423 (O_423,N_2997,N_2963);
and UO_424 (O_424,N_2972,N_2978);
xor UO_425 (O_425,N_2983,N_2969);
nand UO_426 (O_426,N_2971,N_2989);
or UO_427 (O_427,N_2949,N_2972);
nor UO_428 (O_428,N_2927,N_2942);
nor UO_429 (O_429,N_2977,N_2951);
nor UO_430 (O_430,N_2939,N_2970);
xnor UO_431 (O_431,N_2965,N_2985);
or UO_432 (O_432,N_2965,N_2976);
and UO_433 (O_433,N_2996,N_2932);
and UO_434 (O_434,N_2978,N_2970);
and UO_435 (O_435,N_2950,N_2954);
nor UO_436 (O_436,N_2928,N_2945);
xor UO_437 (O_437,N_2966,N_2974);
and UO_438 (O_438,N_2947,N_2927);
and UO_439 (O_439,N_2926,N_2980);
or UO_440 (O_440,N_2964,N_2957);
nand UO_441 (O_441,N_2970,N_2997);
and UO_442 (O_442,N_2926,N_2958);
and UO_443 (O_443,N_2944,N_2974);
and UO_444 (O_444,N_2982,N_2987);
and UO_445 (O_445,N_2990,N_2965);
and UO_446 (O_446,N_2950,N_2935);
or UO_447 (O_447,N_2932,N_2965);
or UO_448 (O_448,N_2972,N_2929);
xnor UO_449 (O_449,N_2991,N_2941);
and UO_450 (O_450,N_2981,N_2994);
and UO_451 (O_451,N_2984,N_2983);
xnor UO_452 (O_452,N_2951,N_2930);
or UO_453 (O_453,N_2971,N_2949);
or UO_454 (O_454,N_2997,N_2933);
nor UO_455 (O_455,N_2943,N_2969);
or UO_456 (O_456,N_2940,N_2967);
nor UO_457 (O_457,N_2927,N_2966);
nand UO_458 (O_458,N_2982,N_2984);
xnor UO_459 (O_459,N_2928,N_2926);
xnor UO_460 (O_460,N_2978,N_2930);
nand UO_461 (O_461,N_2956,N_2988);
or UO_462 (O_462,N_2967,N_2944);
xor UO_463 (O_463,N_2982,N_2986);
or UO_464 (O_464,N_2981,N_2977);
xor UO_465 (O_465,N_2994,N_2986);
nor UO_466 (O_466,N_2956,N_2996);
or UO_467 (O_467,N_2929,N_2991);
xnor UO_468 (O_468,N_2974,N_2953);
nor UO_469 (O_469,N_2933,N_2984);
xnor UO_470 (O_470,N_2962,N_2956);
xor UO_471 (O_471,N_2952,N_2982);
and UO_472 (O_472,N_2971,N_2966);
xnor UO_473 (O_473,N_2989,N_2970);
and UO_474 (O_474,N_2956,N_2984);
xor UO_475 (O_475,N_2951,N_2999);
nor UO_476 (O_476,N_2949,N_2965);
nor UO_477 (O_477,N_2952,N_2987);
or UO_478 (O_478,N_2972,N_2997);
or UO_479 (O_479,N_2939,N_2967);
nor UO_480 (O_480,N_2983,N_2996);
and UO_481 (O_481,N_2930,N_2999);
nor UO_482 (O_482,N_2954,N_2947);
and UO_483 (O_483,N_2942,N_2950);
and UO_484 (O_484,N_2953,N_2942);
xor UO_485 (O_485,N_2990,N_2948);
nor UO_486 (O_486,N_2982,N_2937);
and UO_487 (O_487,N_2939,N_2969);
or UO_488 (O_488,N_2961,N_2984);
and UO_489 (O_489,N_2955,N_2929);
xor UO_490 (O_490,N_2965,N_2999);
and UO_491 (O_491,N_2993,N_2930);
or UO_492 (O_492,N_2938,N_2934);
or UO_493 (O_493,N_2938,N_2945);
xnor UO_494 (O_494,N_2978,N_2928);
or UO_495 (O_495,N_2959,N_2969);
nand UO_496 (O_496,N_2960,N_2964);
or UO_497 (O_497,N_2980,N_2964);
nand UO_498 (O_498,N_2999,N_2932);
or UO_499 (O_499,N_2992,N_2994);
endmodule