module basic_3000_30000_3500_30_levels_10xor_1(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999,N_25000,N_25001,N_25002,N_25003,N_25004,N_25005,N_25006,N_25007,N_25008,N_25009,N_25010,N_25011,N_25012,N_25013,N_25014,N_25015,N_25016,N_25017,N_25018,N_25019,N_25020,N_25021,N_25022,N_25023,N_25024,N_25025,N_25026,N_25027,N_25028,N_25029,N_25030,N_25031,N_25032,N_25033,N_25034,N_25035,N_25036,N_25037,N_25038,N_25039,N_25040,N_25041,N_25042,N_25043,N_25044,N_25045,N_25046,N_25047,N_25048,N_25049,N_25050,N_25051,N_25052,N_25053,N_25054,N_25055,N_25056,N_25057,N_25058,N_25059,N_25060,N_25061,N_25062,N_25063,N_25064,N_25065,N_25066,N_25067,N_25068,N_25069,N_25070,N_25071,N_25072,N_25073,N_25074,N_25075,N_25076,N_25077,N_25078,N_25079,N_25080,N_25081,N_25082,N_25083,N_25084,N_25085,N_25086,N_25087,N_25088,N_25089,N_25090,N_25091,N_25092,N_25093,N_25094,N_25095,N_25096,N_25097,N_25098,N_25099,N_25100,N_25101,N_25102,N_25103,N_25104,N_25105,N_25106,N_25107,N_25108,N_25109,N_25110,N_25111,N_25112,N_25113,N_25114,N_25115,N_25116,N_25117,N_25118,N_25119,N_25120,N_25121,N_25122,N_25123,N_25124,N_25125,N_25126,N_25127,N_25128,N_25129,N_25130,N_25131,N_25132,N_25133,N_25134,N_25135,N_25136,N_25137,N_25138,N_25139,N_25140,N_25141,N_25142,N_25143,N_25144,N_25145,N_25146,N_25147,N_25148,N_25149,N_25150,N_25151,N_25152,N_25153,N_25154,N_25155,N_25156,N_25157,N_25158,N_25159,N_25160,N_25161,N_25162,N_25163,N_25164,N_25165,N_25166,N_25167,N_25168,N_25169,N_25170,N_25171,N_25172,N_25173,N_25174,N_25175,N_25176,N_25177,N_25178,N_25179,N_25180,N_25181,N_25182,N_25183,N_25184,N_25185,N_25186,N_25187,N_25188,N_25189,N_25190,N_25191,N_25192,N_25193,N_25194,N_25195,N_25196,N_25197,N_25198,N_25199,N_25200,N_25201,N_25202,N_25203,N_25204,N_25205,N_25206,N_25207,N_25208,N_25209,N_25210,N_25211,N_25212,N_25213,N_25214,N_25215,N_25216,N_25217,N_25218,N_25219,N_25220,N_25221,N_25222,N_25223,N_25224,N_25225,N_25226,N_25227,N_25228,N_25229,N_25230,N_25231,N_25232,N_25233,N_25234,N_25235,N_25236,N_25237,N_25238,N_25239,N_25240,N_25241,N_25242,N_25243,N_25244,N_25245,N_25246,N_25247,N_25248,N_25249,N_25250,N_25251,N_25252,N_25253,N_25254,N_25255,N_25256,N_25257,N_25258,N_25259,N_25260,N_25261,N_25262,N_25263,N_25264,N_25265,N_25266,N_25267,N_25268,N_25269,N_25270,N_25271,N_25272,N_25273,N_25274,N_25275,N_25276,N_25277,N_25278,N_25279,N_25280,N_25281,N_25282,N_25283,N_25284,N_25285,N_25286,N_25287,N_25288,N_25289,N_25290,N_25291,N_25292,N_25293,N_25294,N_25295,N_25296,N_25297,N_25298,N_25299,N_25300,N_25301,N_25302,N_25303,N_25304,N_25305,N_25306,N_25307,N_25308,N_25309,N_25310,N_25311,N_25312,N_25313,N_25314,N_25315,N_25316,N_25317,N_25318,N_25319,N_25320,N_25321,N_25322,N_25323,N_25324,N_25325,N_25326,N_25327,N_25328,N_25329,N_25330,N_25331,N_25332,N_25333,N_25334,N_25335,N_25336,N_25337,N_25338,N_25339,N_25340,N_25341,N_25342,N_25343,N_25344,N_25345,N_25346,N_25347,N_25348,N_25349,N_25350,N_25351,N_25352,N_25353,N_25354,N_25355,N_25356,N_25357,N_25358,N_25359,N_25360,N_25361,N_25362,N_25363,N_25364,N_25365,N_25366,N_25367,N_25368,N_25369,N_25370,N_25371,N_25372,N_25373,N_25374,N_25375,N_25376,N_25377,N_25378,N_25379,N_25380,N_25381,N_25382,N_25383,N_25384,N_25385,N_25386,N_25387,N_25388,N_25389,N_25390,N_25391,N_25392,N_25393,N_25394,N_25395,N_25396,N_25397,N_25398,N_25399,N_25400,N_25401,N_25402,N_25403,N_25404,N_25405,N_25406,N_25407,N_25408,N_25409,N_25410,N_25411,N_25412,N_25413,N_25414,N_25415,N_25416,N_25417,N_25418,N_25419,N_25420,N_25421,N_25422,N_25423,N_25424,N_25425,N_25426,N_25427,N_25428,N_25429,N_25430,N_25431,N_25432,N_25433,N_25434,N_25435,N_25436,N_25437,N_25438,N_25439,N_25440,N_25441,N_25442,N_25443,N_25444,N_25445,N_25446,N_25447,N_25448,N_25449,N_25450,N_25451,N_25452,N_25453,N_25454,N_25455,N_25456,N_25457,N_25458,N_25459,N_25460,N_25461,N_25462,N_25463,N_25464,N_25465,N_25466,N_25467,N_25468,N_25469,N_25470,N_25471,N_25472,N_25473,N_25474,N_25475,N_25476,N_25477,N_25478,N_25479,N_25480,N_25481,N_25482,N_25483,N_25484,N_25485,N_25486,N_25487,N_25488,N_25489,N_25490,N_25491,N_25492,N_25493,N_25494,N_25495,N_25496,N_25497,N_25498,N_25499,N_25500,N_25501,N_25502,N_25503,N_25504,N_25505,N_25506,N_25507,N_25508,N_25509,N_25510,N_25511,N_25512,N_25513,N_25514,N_25515,N_25516,N_25517,N_25518,N_25519,N_25520,N_25521,N_25522,N_25523,N_25524,N_25525,N_25526,N_25527,N_25528,N_25529,N_25530,N_25531,N_25532,N_25533,N_25534,N_25535,N_25536,N_25537,N_25538,N_25539,N_25540,N_25541,N_25542,N_25543,N_25544,N_25545,N_25546,N_25547,N_25548,N_25549,N_25550,N_25551,N_25552,N_25553,N_25554,N_25555,N_25556,N_25557,N_25558,N_25559,N_25560,N_25561,N_25562,N_25563,N_25564,N_25565,N_25566,N_25567,N_25568,N_25569,N_25570,N_25571,N_25572,N_25573,N_25574,N_25575,N_25576,N_25577,N_25578,N_25579,N_25580,N_25581,N_25582,N_25583,N_25584,N_25585,N_25586,N_25587,N_25588,N_25589,N_25590,N_25591,N_25592,N_25593,N_25594,N_25595,N_25596,N_25597,N_25598,N_25599,N_25600,N_25601,N_25602,N_25603,N_25604,N_25605,N_25606,N_25607,N_25608,N_25609,N_25610,N_25611,N_25612,N_25613,N_25614,N_25615,N_25616,N_25617,N_25618,N_25619,N_25620,N_25621,N_25622,N_25623,N_25624,N_25625,N_25626,N_25627,N_25628,N_25629,N_25630,N_25631,N_25632,N_25633,N_25634,N_25635,N_25636,N_25637,N_25638,N_25639,N_25640,N_25641,N_25642,N_25643,N_25644,N_25645,N_25646,N_25647,N_25648,N_25649,N_25650,N_25651,N_25652,N_25653,N_25654,N_25655,N_25656,N_25657,N_25658,N_25659,N_25660,N_25661,N_25662,N_25663,N_25664,N_25665,N_25666,N_25667,N_25668,N_25669,N_25670,N_25671,N_25672,N_25673,N_25674,N_25675,N_25676,N_25677,N_25678,N_25679,N_25680,N_25681,N_25682,N_25683,N_25684,N_25685,N_25686,N_25687,N_25688,N_25689,N_25690,N_25691,N_25692,N_25693,N_25694,N_25695,N_25696,N_25697,N_25698,N_25699,N_25700,N_25701,N_25702,N_25703,N_25704,N_25705,N_25706,N_25707,N_25708,N_25709,N_25710,N_25711,N_25712,N_25713,N_25714,N_25715,N_25716,N_25717,N_25718,N_25719,N_25720,N_25721,N_25722,N_25723,N_25724,N_25725,N_25726,N_25727,N_25728,N_25729,N_25730,N_25731,N_25732,N_25733,N_25734,N_25735,N_25736,N_25737,N_25738,N_25739,N_25740,N_25741,N_25742,N_25743,N_25744,N_25745,N_25746,N_25747,N_25748,N_25749,N_25750,N_25751,N_25752,N_25753,N_25754,N_25755,N_25756,N_25757,N_25758,N_25759,N_25760,N_25761,N_25762,N_25763,N_25764,N_25765,N_25766,N_25767,N_25768,N_25769,N_25770,N_25771,N_25772,N_25773,N_25774,N_25775,N_25776,N_25777,N_25778,N_25779,N_25780,N_25781,N_25782,N_25783,N_25784,N_25785,N_25786,N_25787,N_25788,N_25789,N_25790,N_25791,N_25792,N_25793,N_25794,N_25795,N_25796,N_25797,N_25798,N_25799,N_25800,N_25801,N_25802,N_25803,N_25804,N_25805,N_25806,N_25807,N_25808,N_25809,N_25810,N_25811,N_25812,N_25813,N_25814,N_25815,N_25816,N_25817,N_25818,N_25819,N_25820,N_25821,N_25822,N_25823,N_25824,N_25825,N_25826,N_25827,N_25828,N_25829,N_25830,N_25831,N_25832,N_25833,N_25834,N_25835,N_25836,N_25837,N_25838,N_25839,N_25840,N_25841,N_25842,N_25843,N_25844,N_25845,N_25846,N_25847,N_25848,N_25849,N_25850,N_25851,N_25852,N_25853,N_25854,N_25855,N_25856,N_25857,N_25858,N_25859,N_25860,N_25861,N_25862,N_25863,N_25864,N_25865,N_25866,N_25867,N_25868,N_25869,N_25870,N_25871,N_25872,N_25873,N_25874,N_25875,N_25876,N_25877,N_25878,N_25879,N_25880,N_25881,N_25882,N_25883,N_25884,N_25885,N_25886,N_25887,N_25888,N_25889,N_25890,N_25891,N_25892,N_25893,N_25894,N_25895,N_25896,N_25897,N_25898,N_25899,N_25900,N_25901,N_25902,N_25903,N_25904,N_25905,N_25906,N_25907,N_25908,N_25909,N_25910,N_25911,N_25912,N_25913,N_25914,N_25915,N_25916,N_25917,N_25918,N_25919,N_25920,N_25921,N_25922,N_25923,N_25924,N_25925,N_25926,N_25927,N_25928,N_25929,N_25930,N_25931,N_25932,N_25933,N_25934,N_25935,N_25936,N_25937,N_25938,N_25939,N_25940,N_25941,N_25942,N_25943,N_25944,N_25945,N_25946,N_25947,N_25948,N_25949,N_25950,N_25951,N_25952,N_25953,N_25954,N_25955,N_25956,N_25957,N_25958,N_25959,N_25960,N_25961,N_25962,N_25963,N_25964,N_25965,N_25966,N_25967,N_25968,N_25969,N_25970,N_25971,N_25972,N_25973,N_25974,N_25975,N_25976,N_25977,N_25978,N_25979,N_25980,N_25981,N_25982,N_25983,N_25984,N_25985,N_25986,N_25987,N_25988,N_25989,N_25990,N_25991,N_25992,N_25993,N_25994,N_25995,N_25996,N_25997,N_25998,N_25999,N_26000,N_26001,N_26002,N_26003,N_26004,N_26005,N_26006,N_26007,N_26008,N_26009,N_26010,N_26011,N_26012,N_26013,N_26014,N_26015,N_26016,N_26017,N_26018,N_26019,N_26020,N_26021,N_26022,N_26023,N_26024,N_26025,N_26026,N_26027,N_26028,N_26029,N_26030,N_26031,N_26032,N_26033,N_26034,N_26035,N_26036,N_26037,N_26038,N_26039,N_26040,N_26041,N_26042,N_26043,N_26044,N_26045,N_26046,N_26047,N_26048,N_26049,N_26050,N_26051,N_26052,N_26053,N_26054,N_26055,N_26056,N_26057,N_26058,N_26059,N_26060,N_26061,N_26062,N_26063,N_26064,N_26065,N_26066,N_26067,N_26068,N_26069,N_26070,N_26071,N_26072,N_26073,N_26074,N_26075,N_26076,N_26077,N_26078,N_26079,N_26080,N_26081,N_26082,N_26083,N_26084,N_26085,N_26086,N_26087,N_26088,N_26089,N_26090,N_26091,N_26092,N_26093,N_26094,N_26095,N_26096,N_26097,N_26098,N_26099,N_26100,N_26101,N_26102,N_26103,N_26104,N_26105,N_26106,N_26107,N_26108,N_26109,N_26110,N_26111,N_26112,N_26113,N_26114,N_26115,N_26116,N_26117,N_26118,N_26119,N_26120,N_26121,N_26122,N_26123,N_26124,N_26125,N_26126,N_26127,N_26128,N_26129,N_26130,N_26131,N_26132,N_26133,N_26134,N_26135,N_26136,N_26137,N_26138,N_26139,N_26140,N_26141,N_26142,N_26143,N_26144,N_26145,N_26146,N_26147,N_26148,N_26149,N_26150,N_26151,N_26152,N_26153,N_26154,N_26155,N_26156,N_26157,N_26158,N_26159,N_26160,N_26161,N_26162,N_26163,N_26164,N_26165,N_26166,N_26167,N_26168,N_26169,N_26170,N_26171,N_26172,N_26173,N_26174,N_26175,N_26176,N_26177,N_26178,N_26179,N_26180,N_26181,N_26182,N_26183,N_26184,N_26185,N_26186,N_26187,N_26188,N_26189,N_26190,N_26191,N_26192,N_26193,N_26194,N_26195,N_26196,N_26197,N_26198,N_26199,N_26200,N_26201,N_26202,N_26203,N_26204,N_26205,N_26206,N_26207,N_26208,N_26209,N_26210,N_26211,N_26212,N_26213,N_26214,N_26215,N_26216,N_26217,N_26218,N_26219,N_26220,N_26221,N_26222,N_26223,N_26224,N_26225,N_26226,N_26227,N_26228,N_26229,N_26230,N_26231,N_26232,N_26233,N_26234,N_26235,N_26236,N_26237,N_26238,N_26239,N_26240,N_26241,N_26242,N_26243,N_26244,N_26245,N_26246,N_26247,N_26248,N_26249,N_26250,N_26251,N_26252,N_26253,N_26254,N_26255,N_26256,N_26257,N_26258,N_26259,N_26260,N_26261,N_26262,N_26263,N_26264,N_26265,N_26266,N_26267,N_26268,N_26269,N_26270,N_26271,N_26272,N_26273,N_26274,N_26275,N_26276,N_26277,N_26278,N_26279,N_26280,N_26281,N_26282,N_26283,N_26284,N_26285,N_26286,N_26287,N_26288,N_26289,N_26290,N_26291,N_26292,N_26293,N_26294,N_26295,N_26296,N_26297,N_26298,N_26299,N_26300,N_26301,N_26302,N_26303,N_26304,N_26305,N_26306,N_26307,N_26308,N_26309,N_26310,N_26311,N_26312,N_26313,N_26314,N_26315,N_26316,N_26317,N_26318,N_26319,N_26320,N_26321,N_26322,N_26323,N_26324,N_26325,N_26326,N_26327,N_26328,N_26329,N_26330,N_26331,N_26332,N_26333,N_26334,N_26335,N_26336,N_26337,N_26338,N_26339,N_26340,N_26341,N_26342,N_26343,N_26344,N_26345,N_26346,N_26347,N_26348,N_26349,N_26350,N_26351,N_26352,N_26353,N_26354,N_26355,N_26356,N_26357,N_26358,N_26359,N_26360,N_26361,N_26362,N_26363,N_26364,N_26365,N_26366,N_26367,N_26368,N_26369,N_26370,N_26371,N_26372,N_26373,N_26374,N_26375,N_26376,N_26377,N_26378,N_26379,N_26380,N_26381,N_26382,N_26383,N_26384,N_26385,N_26386,N_26387,N_26388,N_26389,N_26390,N_26391,N_26392,N_26393,N_26394,N_26395,N_26396,N_26397,N_26398,N_26399,N_26400,N_26401,N_26402,N_26403,N_26404,N_26405,N_26406,N_26407,N_26408,N_26409,N_26410,N_26411,N_26412,N_26413,N_26414,N_26415,N_26416,N_26417,N_26418,N_26419,N_26420,N_26421,N_26422,N_26423,N_26424,N_26425,N_26426,N_26427,N_26428,N_26429,N_26430,N_26431,N_26432,N_26433,N_26434,N_26435,N_26436,N_26437,N_26438,N_26439,N_26440,N_26441,N_26442,N_26443,N_26444,N_26445,N_26446,N_26447,N_26448,N_26449,N_26450,N_26451,N_26452,N_26453,N_26454,N_26455,N_26456,N_26457,N_26458,N_26459,N_26460,N_26461,N_26462,N_26463,N_26464,N_26465,N_26466,N_26467,N_26468,N_26469,N_26470,N_26471,N_26472,N_26473,N_26474,N_26475,N_26476,N_26477,N_26478,N_26479,N_26480,N_26481,N_26482,N_26483,N_26484,N_26485,N_26486,N_26487,N_26488,N_26489,N_26490,N_26491,N_26492,N_26493,N_26494,N_26495,N_26496,N_26497,N_26498,N_26499,N_26500,N_26501,N_26502,N_26503,N_26504,N_26505,N_26506,N_26507,N_26508,N_26509,N_26510,N_26511,N_26512,N_26513,N_26514,N_26515,N_26516,N_26517,N_26518,N_26519,N_26520,N_26521,N_26522,N_26523,N_26524,N_26525,N_26526,N_26527,N_26528,N_26529,N_26530,N_26531,N_26532,N_26533,N_26534,N_26535,N_26536,N_26537,N_26538,N_26539,N_26540,N_26541,N_26542,N_26543,N_26544,N_26545,N_26546,N_26547,N_26548,N_26549,N_26550,N_26551,N_26552,N_26553,N_26554,N_26555,N_26556,N_26557,N_26558,N_26559,N_26560,N_26561,N_26562,N_26563,N_26564,N_26565,N_26566,N_26567,N_26568,N_26569,N_26570,N_26571,N_26572,N_26573,N_26574,N_26575,N_26576,N_26577,N_26578,N_26579,N_26580,N_26581,N_26582,N_26583,N_26584,N_26585,N_26586,N_26587,N_26588,N_26589,N_26590,N_26591,N_26592,N_26593,N_26594,N_26595,N_26596,N_26597,N_26598,N_26599,N_26600,N_26601,N_26602,N_26603,N_26604,N_26605,N_26606,N_26607,N_26608,N_26609,N_26610,N_26611,N_26612,N_26613,N_26614,N_26615,N_26616,N_26617,N_26618,N_26619,N_26620,N_26621,N_26622,N_26623,N_26624,N_26625,N_26626,N_26627,N_26628,N_26629,N_26630,N_26631,N_26632,N_26633,N_26634,N_26635,N_26636,N_26637,N_26638,N_26639,N_26640,N_26641,N_26642,N_26643,N_26644,N_26645,N_26646,N_26647,N_26648,N_26649,N_26650,N_26651,N_26652,N_26653,N_26654,N_26655,N_26656,N_26657,N_26658,N_26659,N_26660,N_26661,N_26662,N_26663,N_26664,N_26665,N_26666,N_26667,N_26668,N_26669,N_26670,N_26671,N_26672,N_26673,N_26674,N_26675,N_26676,N_26677,N_26678,N_26679,N_26680,N_26681,N_26682,N_26683,N_26684,N_26685,N_26686,N_26687,N_26688,N_26689,N_26690,N_26691,N_26692,N_26693,N_26694,N_26695,N_26696,N_26697,N_26698,N_26699,N_26700,N_26701,N_26702,N_26703,N_26704,N_26705,N_26706,N_26707,N_26708,N_26709,N_26710,N_26711,N_26712,N_26713,N_26714,N_26715,N_26716,N_26717,N_26718,N_26719,N_26720,N_26721,N_26722,N_26723,N_26724,N_26725,N_26726,N_26727,N_26728,N_26729,N_26730,N_26731,N_26732,N_26733,N_26734,N_26735,N_26736,N_26737,N_26738,N_26739,N_26740,N_26741,N_26742,N_26743,N_26744,N_26745,N_26746,N_26747,N_26748,N_26749,N_26750,N_26751,N_26752,N_26753,N_26754,N_26755,N_26756,N_26757,N_26758,N_26759,N_26760,N_26761,N_26762,N_26763,N_26764,N_26765,N_26766,N_26767,N_26768,N_26769,N_26770,N_26771,N_26772,N_26773,N_26774,N_26775,N_26776,N_26777,N_26778,N_26779,N_26780,N_26781,N_26782,N_26783,N_26784,N_26785,N_26786,N_26787,N_26788,N_26789,N_26790,N_26791,N_26792,N_26793,N_26794,N_26795,N_26796,N_26797,N_26798,N_26799,N_26800,N_26801,N_26802,N_26803,N_26804,N_26805,N_26806,N_26807,N_26808,N_26809,N_26810,N_26811,N_26812,N_26813,N_26814,N_26815,N_26816,N_26817,N_26818,N_26819,N_26820,N_26821,N_26822,N_26823,N_26824,N_26825,N_26826,N_26827,N_26828,N_26829,N_26830,N_26831,N_26832,N_26833,N_26834,N_26835,N_26836,N_26837,N_26838,N_26839,N_26840,N_26841,N_26842,N_26843,N_26844,N_26845,N_26846,N_26847,N_26848,N_26849,N_26850,N_26851,N_26852,N_26853,N_26854,N_26855,N_26856,N_26857,N_26858,N_26859,N_26860,N_26861,N_26862,N_26863,N_26864,N_26865,N_26866,N_26867,N_26868,N_26869,N_26870,N_26871,N_26872,N_26873,N_26874,N_26875,N_26876,N_26877,N_26878,N_26879,N_26880,N_26881,N_26882,N_26883,N_26884,N_26885,N_26886,N_26887,N_26888,N_26889,N_26890,N_26891,N_26892,N_26893,N_26894,N_26895,N_26896,N_26897,N_26898,N_26899,N_26900,N_26901,N_26902,N_26903,N_26904,N_26905,N_26906,N_26907,N_26908,N_26909,N_26910,N_26911,N_26912,N_26913,N_26914,N_26915,N_26916,N_26917,N_26918,N_26919,N_26920,N_26921,N_26922,N_26923,N_26924,N_26925,N_26926,N_26927,N_26928,N_26929,N_26930,N_26931,N_26932,N_26933,N_26934,N_26935,N_26936,N_26937,N_26938,N_26939,N_26940,N_26941,N_26942,N_26943,N_26944,N_26945,N_26946,N_26947,N_26948,N_26949,N_26950,N_26951,N_26952,N_26953,N_26954,N_26955,N_26956,N_26957,N_26958,N_26959,N_26960,N_26961,N_26962,N_26963,N_26964,N_26965,N_26966,N_26967,N_26968,N_26969,N_26970,N_26971,N_26972,N_26973,N_26974,N_26975,N_26976,N_26977,N_26978,N_26979,N_26980,N_26981,N_26982,N_26983,N_26984,N_26985,N_26986,N_26987,N_26988,N_26989,N_26990,N_26991,N_26992,N_26993,N_26994,N_26995,N_26996,N_26997,N_26998,N_26999,N_27000,N_27001,N_27002,N_27003,N_27004,N_27005,N_27006,N_27007,N_27008,N_27009,N_27010,N_27011,N_27012,N_27013,N_27014,N_27015,N_27016,N_27017,N_27018,N_27019,N_27020,N_27021,N_27022,N_27023,N_27024,N_27025,N_27026,N_27027,N_27028,N_27029,N_27030,N_27031,N_27032,N_27033,N_27034,N_27035,N_27036,N_27037,N_27038,N_27039,N_27040,N_27041,N_27042,N_27043,N_27044,N_27045,N_27046,N_27047,N_27048,N_27049,N_27050,N_27051,N_27052,N_27053,N_27054,N_27055,N_27056,N_27057,N_27058,N_27059,N_27060,N_27061,N_27062,N_27063,N_27064,N_27065,N_27066,N_27067,N_27068,N_27069,N_27070,N_27071,N_27072,N_27073,N_27074,N_27075,N_27076,N_27077,N_27078,N_27079,N_27080,N_27081,N_27082,N_27083,N_27084,N_27085,N_27086,N_27087,N_27088,N_27089,N_27090,N_27091,N_27092,N_27093,N_27094,N_27095,N_27096,N_27097,N_27098,N_27099,N_27100,N_27101,N_27102,N_27103,N_27104,N_27105,N_27106,N_27107,N_27108,N_27109,N_27110,N_27111,N_27112,N_27113,N_27114,N_27115,N_27116,N_27117,N_27118,N_27119,N_27120,N_27121,N_27122,N_27123,N_27124,N_27125,N_27126,N_27127,N_27128,N_27129,N_27130,N_27131,N_27132,N_27133,N_27134,N_27135,N_27136,N_27137,N_27138,N_27139,N_27140,N_27141,N_27142,N_27143,N_27144,N_27145,N_27146,N_27147,N_27148,N_27149,N_27150,N_27151,N_27152,N_27153,N_27154,N_27155,N_27156,N_27157,N_27158,N_27159,N_27160,N_27161,N_27162,N_27163,N_27164,N_27165,N_27166,N_27167,N_27168,N_27169,N_27170,N_27171,N_27172,N_27173,N_27174,N_27175,N_27176,N_27177,N_27178,N_27179,N_27180,N_27181,N_27182,N_27183,N_27184,N_27185,N_27186,N_27187,N_27188,N_27189,N_27190,N_27191,N_27192,N_27193,N_27194,N_27195,N_27196,N_27197,N_27198,N_27199,N_27200,N_27201,N_27202,N_27203,N_27204,N_27205,N_27206,N_27207,N_27208,N_27209,N_27210,N_27211,N_27212,N_27213,N_27214,N_27215,N_27216,N_27217,N_27218,N_27219,N_27220,N_27221,N_27222,N_27223,N_27224,N_27225,N_27226,N_27227,N_27228,N_27229,N_27230,N_27231,N_27232,N_27233,N_27234,N_27235,N_27236,N_27237,N_27238,N_27239,N_27240,N_27241,N_27242,N_27243,N_27244,N_27245,N_27246,N_27247,N_27248,N_27249,N_27250,N_27251,N_27252,N_27253,N_27254,N_27255,N_27256,N_27257,N_27258,N_27259,N_27260,N_27261,N_27262,N_27263,N_27264,N_27265,N_27266,N_27267,N_27268,N_27269,N_27270,N_27271,N_27272,N_27273,N_27274,N_27275,N_27276,N_27277,N_27278,N_27279,N_27280,N_27281,N_27282,N_27283,N_27284,N_27285,N_27286,N_27287,N_27288,N_27289,N_27290,N_27291,N_27292,N_27293,N_27294,N_27295,N_27296,N_27297,N_27298,N_27299,N_27300,N_27301,N_27302,N_27303,N_27304,N_27305,N_27306,N_27307,N_27308,N_27309,N_27310,N_27311,N_27312,N_27313,N_27314,N_27315,N_27316,N_27317,N_27318,N_27319,N_27320,N_27321,N_27322,N_27323,N_27324,N_27325,N_27326,N_27327,N_27328,N_27329,N_27330,N_27331,N_27332,N_27333,N_27334,N_27335,N_27336,N_27337,N_27338,N_27339,N_27340,N_27341,N_27342,N_27343,N_27344,N_27345,N_27346,N_27347,N_27348,N_27349,N_27350,N_27351,N_27352,N_27353,N_27354,N_27355,N_27356,N_27357,N_27358,N_27359,N_27360,N_27361,N_27362,N_27363,N_27364,N_27365,N_27366,N_27367,N_27368,N_27369,N_27370,N_27371,N_27372,N_27373,N_27374,N_27375,N_27376,N_27377,N_27378,N_27379,N_27380,N_27381,N_27382,N_27383,N_27384,N_27385,N_27386,N_27387,N_27388,N_27389,N_27390,N_27391,N_27392,N_27393,N_27394,N_27395,N_27396,N_27397,N_27398,N_27399,N_27400,N_27401,N_27402,N_27403,N_27404,N_27405,N_27406,N_27407,N_27408,N_27409,N_27410,N_27411,N_27412,N_27413,N_27414,N_27415,N_27416,N_27417,N_27418,N_27419,N_27420,N_27421,N_27422,N_27423,N_27424,N_27425,N_27426,N_27427,N_27428,N_27429,N_27430,N_27431,N_27432,N_27433,N_27434,N_27435,N_27436,N_27437,N_27438,N_27439,N_27440,N_27441,N_27442,N_27443,N_27444,N_27445,N_27446,N_27447,N_27448,N_27449,N_27450,N_27451,N_27452,N_27453,N_27454,N_27455,N_27456,N_27457,N_27458,N_27459,N_27460,N_27461,N_27462,N_27463,N_27464,N_27465,N_27466,N_27467,N_27468,N_27469,N_27470,N_27471,N_27472,N_27473,N_27474,N_27475,N_27476,N_27477,N_27478,N_27479,N_27480,N_27481,N_27482,N_27483,N_27484,N_27485,N_27486,N_27487,N_27488,N_27489,N_27490,N_27491,N_27492,N_27493,N_27494,N_27495,N_27496,N_27497,N_27498,N_27499,N_27500,N_27501,N_27502,N_27503,N_27504,N_27505,N_27506,N_27507,N_27508,N_27509,N_27510,N_27511,N_27512,N_27513,N_27514,N_27515,N_27516,N_27517,N_27518,N_27519,N_27520,N_27521,N_27522,N_27523,N_27524,N_27525,N_27526,N_27527,N_27528,N_27529,N_27530,N_27531,N_27532,N_27533,N_27534,N_27535,N_27536,N_27537,N_27538,N_27539,N_27540,N_27541,N_27542,N_27543,N_27544,N_27545,N_27546,N_27547,N_27548,N_27549,N_27550,N_27551,N_27552,N_27553,N_27554,N_27555,N_27556,N_27557,N_27558,N_27559,N_27560,N_27561,N_27562,N_27563,N_27564,N_27565,N_27566,N_27567,N_27568,N_27569,N_27570,N_27571,N_27572,N_27573,N_27574,N_27575,N_27576,N_27577,N_27578,N_27579,N_27580,N_27581,N_27582,N_27583,N_27584,N_27585,N_27586,N_27587,N_27588,N_27589,N_27590,N_27591,N_27592,N_27593,N_27594,N_27595,N_27596,N_27597,N_27598,N_27599,N_27600,N_27601,N_27602,N_27603,N_27604,N_27605,N_27606,N_27607,N_27608,N_27609,N_27610,N_27611,N_27612,N_27613,N_27614,N_27615,N_27616,N_27617,N_27618,N_27619,N_27620,N_27621,N_27622,N_27623,N_27624,N_27625,N_27626,N_27627,N_27628,N_27629,N_27630,N_27631,N_27632,N_27633,N_27634,N_27635,N_27636,N_27637,N_27638,N_27639,N_27640,N_27641,N_27642,N_27643,N_27644,N_27645,N_27646,N_27647,N_27648,N_27649,N_27650,N_27651,N_27652,N_27653,N_27654,N_27655,N_27656,N_27657,N_27658,N_27659,N_27660,N_27661,N_27662,N_27663,N_27664,N_27665,N_27666,N_27667,N_27668,N_27669,N_27670,N_27671,N_27672,N_27673,N_27674,N_27675,N_27676,N_27677,N_27678,N_27679,N_27680,N_27681,N_27682,N_27683,N_27684,N_27685,N_27686,N_27687,N_27688,N_27689,N_27690,N_27691,N_27692,N_27693,N_27694,N_27695,N_27696,N_27697,N_27698,N_27699,N_27700,N_27701,N_27702,N_27703,N_27704,N_27705,N_27706,N_27707,N_27708,N_27709,N_27710,N_27711,N_27712,N_27713,N_27714,N_27715,N_27716,N_27717,N_27718,N_27719,N_27720,N_27721,N_27722,N_27723,N_27724,N_27725,N_27726,N_27727,N_27728,N_27729,N_27730,N_27731,N_27732,N_27733,N_27734,N_27735,N_27736,N_27737,N_27738,N_27739,N_27740,N_27741,N_27742,N_27743,N_27744,N_27745,N_27746,N_27747,N_27748,N_27749,N_27750,N_27751,N_27752,N_27753,N_27754,N_27755,N_27756,N_27757,N_27758,N_27759,N_27760,N_27761,N_27762,N_27763,N_27764,N_27765,N_27766,N_27767,N_27768,N_27769,N_27770,N_27771,N_27772,N_27773,N_27774,N_27775,N_27776,N_27777,N_27778,N_27779,N_27780,N_27781,N_27782,N_27783,N_27784,N_27785,N_27786,N_27787,N_27788,N_27789,N_27790,N_27791,N_27792,N_27793,N_27794,N_27795,N_27796,N_27797,N_27798,N_27799,N_27800,N_27801,N_27802,N_27803,N_27804,N_27805,N_27806,N_27807,N_27808,N_27809,N_27810,N_27811,N_27812,N_27813,N_27814,N_27815,N_27816,N_27817,N_27818,N_27819,N_27820,N_27821,N_27822,N_27823,N_27824,N_27825,N_27826,N_27827,N_27828,N_27829,N_27830,N_27831,N_27832,N_27833,N_27834,N_27835,N_27836,N_27837,N_27838,N_27839,N_27840,N_27841,N_27842,N_27843,N_27844,N_27845,N_27846,N_27847,N_27848,N_27849,N_27850,N_27851,N_27852,N_27853,N_27854,N_27855,N_27856,N_27857,N_27858,N_27859,N_27860,N_27861,N_27862,N_27863,N_27864,N_27865,N_27866,N_27867,N_27868,N_27869,N_27870,N_27871,N_27872,N_27873,N_27874,N_27875,N_27876,N_27877,N_27878,N_27879,N_27880,N_27881,N_27882,N_27883,N_27884,N_27885,N_27886,N_27887,N_27888,N_27889,N_27890,N_27891,N_27892,N_27893,N_27894,N_27895,N_27896,N_27897,N_27898,N_27899,N_27900,N_27901,N_27902,N_27903,N_27904,N_27905,N_27906,N_27907,N_27908,N_27909,N_27910,N_27911,N_27912,N_27913,N_27914,N_27915,N_27916,N_27917,N_27918,N_27919,N_27920,N_27921,N_27922,N_27923,N_27924,N_27925,N_27926,N_27927,N_27928,N_27929,N_27930,N_27931,N_27932,N_27933,N_27934,N_27935,N_27936,N_27937,N_27938,N_27939,N_27940,N_27941,N_27942,N_27943,N_27944,N_27945,N_27946,N_27947,N_27948,N_27949,N_27950,N_27951,N_27952,N_27953,N_27954,N_27955,N_27956,N_27957,N_27958,N_27959,N_27960,N_27961,N_27962,N_27963,N_27964,N_27965,N_27966,N_27967,N_27968,N_27969,N_27970,N_27971,N_27972,N_27973,N_27974,N_27975,N_27976,N_27977,N_27978,N_27979,N_27980,N_27981,N_27982,N_27983,N_27984,N_27985,N_27986,N_27987,N_27988,N_27989,N_27990,N_27991,N_27992,N_27993,N_27994,N_27995,N_27996,N_27997,N_27998,N_27999,N_28000,N_28001,N_28002,N_28003,N_28004,N_28005,N_28006,N_28007,N_28008,N_28009,N_28010,N_28011,N_28012,N_28013,N_28014,N_28015,N_28016,N_28017,N_28018,N_28019,N_28020,N_28021,N_28022,N_28023,N_28024,N_28025,N_28026,N_28027,N_28028,N_28029,N_28030,N_28031,N_28032,N_28033,N_28034,N_28035,N_28036,N_28037,N_28038,N_28039,N_28040,N_28041,N_28042,N_28043,N_28044,N_28045,N_28046,N_28047,N_28048,N_28049,N_28050,N_28051,N_28052,N_28053,N_28054,N_28055,N_28056,N_28057,N_28058,N_28059,N_28060,N_28061,N_28062,N_28063,N_28064,N_28065,N_28066,N_28067,N_28068,N_28069,N_28070,N_28071,N_28072,N_28073,N_28074,N_28075,N_28076,N_28077,N_28078,N_28079,N_28080,N_28081,N_28082,N_28083,N_28084,N_28085,N_28086,N_28087,N_28088,N_28089,N_28090,N_28091,N_28092,N_28093,N_28094,N_28095,N_28096,N_28097,N_28098,N_28099,N_28100,N_28101,N_28102,N_28103,N_28104,N_28105,N_28106,N_28107,N_28108,N_28109,N_28110,N_28111,N_28112,N_28113,N_28114,N_28115,N_28116,N_28117,N_28118,N_28119,N_28120,N_28121,N_28122,N_28123,N_28124,N_28125,N_28126,N_28127,N_28128,N_28129,N_28130,N_28131,N_28132,N_28133,N_28134,N_28135,N_28136,N_28137,N_28138,N_28139,N_28140,N_28141,N_28142,N_28143,N_28144,N_28145,N_28146,N_28147,N_28148,N_28149,N_28150,N_28151,N_28152,N_28153,N_28154,N_28155,N_28156,N_28157,N_28158,N_28159,N_28160,N_28161,N_28162,N_28163,N_28164,N_28165,N_28166,N_28167,N_28168,N_28169,N_28170,N_28171,N_28172,N_28173,N_28174,N_28175,N_28176,N_28177,N_28178,N_28179,N_28180,N_28181,N_28182,N_28183,N_28184,N_28185,N_28186,N_28187,N_28188,N_28189,N_28190,N_28191,N_28192,N_28193,N_28194,N_28195,N_28196,N_28197,N_28198,N_28199,N_28200,N_28201,N_28202,N_28203,N_28204,N_28205,N_28206,N_28207,N_28208,N_28209,N_28210,N_28211,N_28212,N_28213,N_28214,N_28215,N_28216,N_28217,N_28218,N_28219,N_28220,N_28221,N_28222,N_28223,N_28224,N_28225,N_28226,N_28227,N_28228,N_28229,N_28230,N_28231,N_28232,N_28233,N_28234,N_28235,N_28236,N_28237,N_28238,N_28239,N_28240,N_28241,N_28242,N_28243,N_28244,N_28245,N_28246,N_28247,N_28248,N_28249,N_28250,N_28251,N_28252,N_28253,N_28254,N_28255,N_28256,N_28257,N_28258,N_28259,N_28260,N_28261,N_28262,N_28263,N_28264,N_28265,N_28266,N_28267,N_28268,N_28269,N_28270,N_28271,N_28272,N_28273,N_28274,N_28275,N_28276,N_28277,N_28278,N_28279,N_28280,N_28281,N_28282,N_28283,N_28284,N_28285,N_28286,N_28287,N_28288,N_28289,N_28290,N_28291,N_28292,N_28293,N_28294,N_28295,N_28296,N_28297,N_28298,N_28299,N_28300,N_28301,N_28302,N_28303,N_28304,N_28305,N_28306,N_28307,N_28308,N_28309,N_28310,N_28311,N_28312,N_28313,N_28314,N_28315,N_28316,N_28317,N_28318,N_28319,N_28320,N_28321,N_28322,N_28323,N_28324,N_28325,N_28326,N_28327,N_28328,N_28329,N_28330,N_28331,N_28332,N_28333,N_28334,N_28335,N_28336,N_28337,N_28338,N_28339,N_28340,N_28341,N_28342,N_28343,N_28344,N_28345,N_28346,N_28347,N_28348,N_28349,N_28350,N_28351,N_28352,N_28353,N_28354,N_28355,N_28356,N_28357,N_28358,N_28359,N_28360,N_28361,N_28362,N_28363,N_28364,N_28365,N_28366,N_28367,N_28368,N_28369,N_28370,N_28371,N_28372,N_28373,N_28374,N_28375,N_28376,N_28377,N_28378,N_28379,N_28380,N_28381,N_28382,N_28383,N_28384,N_28385,N_28386,N_28387,N_28388,N_28389,N_28390,N_28391,N_28392,N_28393,N_28394,N_28395,N_28396,N_28397,N_28398,N_28399,N_28400,N_28401,N_28402,N_28403,N_28404,N_28405,N_28406,N_28407,N_28408,N_28409,N_28410,N_28411,N_28412,N_28413,N_28414,N_28415,N_28416,N_28417,N_28418,N_28419,N_28420,N_28421,N_28422,N_28423,N_28424,N_28425,N_28426,N_28427,N_28428,N_28429,N_28430,N_28431,N_28432,N_28433,N_28434,N_28435,N_28436,N_28437,N_28438,N_28439,N_28440,N_28441,N_28442,N_28443,N_28444,N_28445,N_28446,N_28447,N_28448,N_28449,N_28450,N_28451,N_28452,N_28453,N_28454,N_28455,N_28456,N_28457,N_28458,N_28459,N_28460,N_28461,N_28462,N_28463,N_28464,N_28465,N_28466,N_28467,N_28468,N_28469,N_28470,N_28471,N_28472,N_28473,N_28474,N_28475,N_28476,N_28477,N_28478,N_28479,N_28480,N_28481,N_28482,N_28483,N_28484,N_28485,N_28486,N_28487,N_28488,N_28489,N_28490,N_28491,N_28492,N_28493,N_28494,N_28495,N_28496,N_28497,N_28498,N_28499,N_28500,N_28501,N_28502,N_28503,N_28504,N_28505,N_28506,N_28507,N_28508,N_28509,N_28510,N_28511,N_28512,N_28513,N_28514,N_28515,N_28516,N_28517,N_28518,N_28519,N_28520,N_28521,N_28522,N_28523,N_28524,N_28525,N_28526,N_28527,N_28528,N_28529,N_28530,N_28531,N_28532,N_28533,N_28534,N_28535,N_28536,N_28537,N_28538,N_28539,N_28540,N_28541,N_28542,N_28543,N_28544,N_28545,N_28546,N_28547,N_28548,N_28549,N_28550,N_28551,N_28552,N_28553,N_28554,N_28555,N_28556,N_28557,N_28558,N_28559,N_28560,N_28561,N_28562,N_28563,N_28564,N_28565,N_28566,N_28567,N_28568,N_28569,N_28570,N_28571,N_28572,N_28573,N_28574,N_28575,N_28576,N_28577,N_28578,N_28579,N_28580,N_28581,N_28582,N_28583,N_28584,N_28585,N_28586,N_28587,N_28588,N_28589,N_28590,N_28591,N_28592,N_28593,N_28594,N_28595,N_28596,N_28597,N_28598,N_28599,N_28600,N_28601,N_28602,N_28603,N_28604,N_28605,N_28606,N_28607,N_28608,N_28609,N_28610,N_28611,N_28612,N_28613,N_28614,N_28615,N_28616,N_28617,N_28618,N_28619,N_28620,N_28621,N_28622,N_28623,N_28624,N_28625,N_28626,N_28627,N_28628,N_28629,N_28630,N_28631,N_28632,N_28633,N_28634,N_28635,N_28636,N_28637,N_28638,N_28639,N_28640,N_28641,N_28642,N_28643,N_28644,N_28645,N_28646,N_28647,N_28648,N_28649,N_28650,N_28651,N_28652,N_28653,N_28654,N_28655,N_28656,N_28657,N_28658,N_28659,N_28660,N_28661,N_28662,N_28663,N_28664,N_28665,N_28666,N_28667,N_28668,N_28669,N_28670,N_28671,N_28672,N_28673,N_28674,N_28675,N_28676,N_28677,N_28678,N_28679,N_28680,N_28681,N_28682,N_28683,N_28684,N_28685,N_28686,N_28687,N_28688,N_28689,N_28690,N_28691,N_28692,N_28693,N_28694,N_28695,N_28696,N_28697,N_28698,N_28699,N_28700,N_28701,N_28702,N_28703,N_28704,N_28705,N_28706,N_28707,N_28708,N_28709,N_28710,N_28711,N_28712,N_28713,N_28714,N_28715,N_28716,N_28717,N_28718,N_28719,N_28720,N_28721,N_28722,N_28723,N_28724,N_28725,N_28726,N_28727,N_28728,N_28729,N_28730,N_28731,N_28732,N_28733,N_28734,N_28735,N_28736,N_28737,N_28738,N_28739,N_28740,N_28741,N_28742,N_28743,N_28744,N_28745,N_28746,N_28747,N_28748,N_28749,N_28750,N_28751,N_28752,N_28753,N_28754,N_28755,N_28756,N_28757,N_28758,N_28759,N_28760,N_28761,N_28762,N_28763,N_28764,N_28765,N_28766,N_28767,N_28768,N_28769,N_28770,N_28771,N_28772,N_28773,N_28774,N_28775,N_28776,N_28777,N_28778,N_28779,N_28780,N_28781,N_28782,N_28783,N_28784,N_28785,N_28786,N_28787,N_28788,N_28789,N_28790,N_28791,N_28792,N_28793,N_28794,N_28795,N_28796,N_28797,N_28798,N_28799,N_28800,N_28801,N_28802,N_28803,N_28804,N_28805,N_28806,N_28807,N_28808,N_28809,N_28810,N_28811,N_28812,N_28813,N_28814,N_28815,N_28816,N_28817,N_28818,N_28819,N_28820,N_28821,N_28822,N_28823,N_28824,N_28825,N_28826,N_28827,N_28828,N_28829,N_28830,N_28831,N_28832,N_28833,N_28834,N_28835,N_28836,N_28837,N_28838,N_28839,N_28840,N_28841,N_28842,N_28843,N_28844,N_28845,N_28846,N_28847,N_28848,N_28849,N_28850,N_28851,N_28852,N_28853,N_28854,N_28855,N_28856,N_28857,N_28858,N_28859,N_28860,N_28861,N_28862,N_28863,N_28864,N_28865,N_28866,N_28867,N_28868,N_28869,N_28870,N_28871,N_28872,N_28873,N_28874,N_28875,N_28876,N_28877,N_28878,N_28879,N_28880,N_28881,N_28882,N_28883,N_28884,N_28885,N_28886,N_28887,N_28888,N_28889,N_28890,N_28891,N_28892,N_28893,N_28894,N_28895,N_28896,N_28897,N_28898,N_28899,N_28900,N_28901,N_28902,N_28903,N_28904,N_28905,N_28906,N_28907,N_28908,N_28909,N_28910,N_28911,N_28912,N_28913,N_28914,N_28915,N_28916,N_28917,N_28918,N_28919,N_28920,N_28921,N_28922,N_28923,N_28924,N_28925,N_28926,N_28927,N_28928,N_28929,N_28930,N_28931,N_28932,N_28933,N_28934,N_28935,N_28936,N_28937,N_28938,N_28939,N_28940,N_28941,N_28942,N_28943,N_28944,N_28945,N_28946,N_28947,N_28948,N_28949,N_28950,N_28951,N_28952,N_28953,N_28954,N_28955,N_28956,N_28957,N_28958,N_28959,N_28960,N_28961,N_28962,N_28963,N_28964,N_28965,N_28966,N_28967,N_28968,N_28969,N_28970,N_28971,N_28972,N_28973,N_28974,N_28975,N_28976,N_28977,N_28978,N_28979,N_28980,N_28981,N_28982,N_28983,N_28984,N_28985,N_28986,N_28987,N_28988,N_28989,N_28990,N_28991,N_28992,N_28993,N_28994,N_28995,N_28996,N_28997,N_28998,N_28999,N_29000,N_29001,N_29002,N_29003,N_29004,N_29005,N_29006,N_29007,N_29008,N_29009,N_29010,N_29011,N_29012,N_29013,N_29014,N_29015,N_29016,N_29017,N_29018,N_29019,N_29020,N_29021,N_29022,N_29023,N_29024,N_29025,N_29026,N_29027,N_29028,N_29029,N_29030,N_29031,N_29032,N_29033,N_29034,N_29035,N_29036,N_29037,N_29038,N_29039,N_29040,N_29041,N_29042,N_29043,N_29044,N_29045,N_29046,N_29047,N_29048,N_29049,N_29050,N_29051,N_29052,N_29053,N_29054,N_29055,N_29056,N_29057,N_29058,N_29059,N_29060,N_29061,N_29062,N_29063,N_29064,N_29065,N_29066,N_29067,N_29068,N_29069,N_29070,N_29071,N_29072,N_29073,N_29074,N_29075,N_29076,N_29077,N_29078,N_29079,N_29080,N_29081,N_29082,N_29083,N_29084,N_29085,N_29086,N_29087,N_29088,N_29089,N_29090,N_29091,N_29092,N_29093,N_29094,N_29095,N_29096,N_29097,N_29098,N_29099,N_29100,N_29101,N_29102,N_29103,N_29104,N_29105,N_29106,N_29107,N_29108,N_29109,N_29110,N_29111,N_29112,N_29113,N_29114,N_29115,N_29116,N_29117,N_29118,N_29119,N_29120,N_29121,N_29122,N_29123,N_29124,N_29125,N_29126,N_29127,N_29128,N_29129,N_29130,N_29131,N_29132,N_29133,N_29134,N_29135,N_29136,N_29137,N_29138,N_29139,N_29140,N_29141,N_29142,N_29143,N_29144,N_29145,N_29146,N_29147,N_29148,N_29149,N_29150,N_29151,N_29152,N_29153,N_29154,N_29155,N_29156,N_29157,N_29158,N_29159,N_29160,N_29161,N_29162,N_29163,N_29164,N_29165,N_29166,N_29167,N_29168,N_29169,N_29170,N_29171,N_29172,N_29173,N_29174,N_29175,N_29176,N_29177,N_29178,N_29179,N_29180,N_29181,N_29182,N_29183,N_29184,N_29185,N_29186,N_29187,N_29188,N_29189,N_29190,N_29191,N_29192,N_29193,N_29194,N_29195,N_29196,N_29197,N_29198,N_29199,N_29200,N_29201,N_29202,N_29203,N_29204,N_29205,N_29206,N_29207,N_29208,N_29209,N_29210,N_29211,N_29212,N_29213,N_29214,N_29215,N_29216,N_29217,N_29218,N_29219,N_29220,N_29221,N_29222,N_29223,N_29224,N_29225,N_29226,N_29227,N_29228,N_29229,N_29230,N_29231,N_29232,N_29233,N_29234,N_29235,N_29236,N_29237,N_29238,N_29239,N_29240,N_29241,N_29242,N_29243,N_29244,N_29245,N_29246,N_29247,N_29248,N_29249,N_29250,N_29251,N_29252,N_29253,N_29254,N_29255,N_29256,N_29257,N_29258,N_29259,N_29260,N_29261,N_29262,N_29263,N_29264,N_29265,N_29266,N_29267,N_29268,N_29269,N_29270,N_29271,N_29272,N_29273,N_29274,N_29275,N_29276,N_29277,N_29278,N_29279,N_29280,N_29281,N_29282,N_29283,N_29284,N_29285,N_29286,N_29287,N_29288,N_29289,N_29290,N_29291,N_29292,N_29293,N_29294,N_29295,N_29296,N_29297,N_29298,N_29299,N_29300,N_29301,N_29302,N_29303,N_29304,N_29305,N_29306,N_29307,N_29308,N_29309,N_29310,N_29311,N_29312,N_29313,N_29314,N_29315,N_29316,N_29317,N_29318,N_29319,N_29320,N_29321,N_29322,N_29323,N_29324,N_29325,N_29326,N_29327,N_29328,N_29329,N_29330,N_29331,N_29332,N_29333,N_29334,N_29335,N_29336,N_29337,N_29338,N_29339,N_29340,N_29341,N_29342,N_29343,N_29344,N_29345,N_29346,N_29347,N_29348,N_29349,N_29350,N_29351,N_29352,N_29353,N_29354,N_29355,N_29356,N_29357,N_29358,N_29359,N_29360,N_29361,N_29362,N_29363,N_29364,N_29365,N_29366,N_29367,N_29368,N_29369,N_29370,N_29371,N_29372,N_29373,N_29374,N_29375,N_29376,N_29377,N_29378,N_29379,N_29380,N_29381,N_29382,N_29383,N_29384,N_29385,N_29386,N_29387,N_29388,N_29389,N_29390,N_29391,N_29392,N_29393,N_29394,N_29395,N_29396,N_29397,N_29398,N_29399,N_29400,N_29401,N_29402,N_29403,N_29404,N_29405,N_29406,N_29407,N_29408,N_29409,N_29410,N_29411,N_29412,N_29413,N_29414,N_29415,N_29416,N_29417,N_29418,N_29419,N_29420,N_29421,N_29422,N_29423,N_29424,N_29425,N_29426,N_29427,N_29428,N_29429,N_29430,N_29431,N_29432,N_29433,N_29434,N_29435,N_29436,N_29437,N_29438,N_29439,N_29440,N_29441,N_29442,N_29443,N_29444,N_29445,N_29446,N_29447,N_29448,N_29449,N_29450,N_29451,N_29452,N_29453,N_29454,N_29455,N_29456,N_29457,N_29458,N_29459,N_29460,N_29461,N_29462,N_29463,N_29464,N_29465,N_29466,N_29467,N_29468,N_29469,N_29470,N_29471,N_29472,N_29473,N_29474,N_29475,N_29476,N_29477,N_29478,N_29479,N_29480,N_29481,N_29482,N_29483,N_29484,N_29485,N_29486,N_29487,N_29488,N_29489,N_29490,N_29491,N_29492,N_29493,N_29494,N_29495,N_29496,N_29497,N_29498,N_29499,N_29500,N_29501,N_29502,N_29503,N_29504,N_29505,N_29506,N_29507,N_29508,N_29509,N_29510,N_29511,N_29512,N_29513,N_29514,N_29515,N_29516,N_29517,N_29518,N_29519,N_29520,N_29521,N_29522,N_29523,N_29524,N_29525,N_29526,N_29527,N_29528,N_29529,N_29530,N_29531,N_29532,N_29533,N_29534,N_29535,N_29536,N_29537,N_29538,N_29539,N_29540,N_29541,N_29542,N_29543,N_29544,N_29545,N_29546,N_29547,N_29548,N_29549,N_29550,N_29551,N_29552,N_29553,N_29554,N_29555,N_29556,N_29557,N_29558,N_29559,N_29560,N_29561,N_29562,N_29563,N_29564,N_29565,N_29566,N_29567,N_29568,N_29569,N_29570,N_29571,N_29572,N_29573,N_29574,N_29575,N_29576,N_29577,N_29578,N_29579,N_29580,N_29581,N_29582,N_29583,N_29584,N_29585,N_29586,N_29587,N_29588,N_29589,N_29590,N_29591,N_29592,N_29593,N_29594,N_29595,N_29596,N_29597,N_29598,N_29599,N_29600,N_29601,N_29602,N_29603,N_29604,N_29605,N_29606,N_29607,N_29608,N_29609,N_29610,N_29611,N_29612,N_29613,N_29614,N_29615,N_29616,N_29617,N_29618,N_29619,N_29620,N_29621,N_29622,N_29623,N_29624,N_29625,N_29626,N_29627,N_29628,N_29629,N_29630,N_29631,N_29632,N_29633,N_29634,N_29635,N_29636,N_29637,N_29638,N_29639,N_29640,N_29641,N_29642,N_29643,N_29644,N_29645,N_29646,N_29647,N_29648,N_29649,N_29650,N_29651,N_29652,N_29653,N_29654,N_29655,N_29656,N_29657,N_29658,N_29659,N_29660,N_29661,N_29662,N_29663,N_29664,N_29665,N_29666,N_29667,N_29668,N_29669,N_29670,N_29671,N_29672,N_29673,N_29674,N_29675,N_29676,N_29677,N_29678,N_29679,N_29680,N_29681,N_29682,N_29683,N_29684,N_29685,N_29686,N_29687,N_29688,N_29689,N_29690,N_29691,N_29692,N_29693,N_29694,N_29695,N_29696,N_29697,N_29698,N_29699,N_29700,N_29701,N_29702,N_29703,N_29704,N_29705,N_29706,N_29707,N_29708,N_29709,N_29710,N_29711,N_29712,N_29713,N_29714,N_29715,N_29716,N_29717,N_29718,N_29719,N_29720,N_29721,N_29722,N_29723,N_29724,N_29725,N_29726,N_29727,N_29728,N_29729,N_29730,N_29731,N_29732,N_29733,N_29734,N_29735,N_29736,N_29737,N_29738,N_29739,N_29740,N_29741,N_29742,N_29743,N_29744,N_29745,N_29746,N_29747,N_29748,N_29749,N_29750,N_29751,N_29752,N_29753,N_29754,N_29755,N_29756,N_29757,N_29758,N_29759,N_29760,N_29761,N_29762,N_29763,N_29764,N_29765,N_29766,N_29767,N_29768,N_29769,N_29770,N_29771,N_29772,N_29773,N_29774,N_29775,N_29776,N_29777,N_29778,N_29779,N_29780,N_29781,N_29782,N_29783,N_29784,N_29785,N_29786,N_29787,N_29788,N_29789,N_29790,N_29791,N_29792,N_29793,N_29794,N_29795,N_29796,N_29797,N_29798,N_29799,N_29800,N_29801,N_29802,N_29803,N_29804,N_29805,N_29806,N_29807,N_29808,N_29809,N_29810,N_29811,N_29812,N_29813,N_29814,N_29815,N_29816,N_29817,N_29818,N_29819,N_29820,N_29821,N_29822,N_29823,N_29824,N_29825,N_29826,N_29827,N_29828,N_29829,N_29830,N_29831,N_29832,N_29833,N_29834,N_29835,N_29836,N_29837,N_29838,N_29839,N_29840,N_29841,N_29842,N_29843,N_29844,N_29845,N_29846,N_29847,N_29848,N_29849,N_29850,N_29851,N_29852,N_29853,N_29854,N_29855,N_29856,N_29857,N_29858,N_29859,N_29860,N_29861,N_29862,N_29863,N_29864,N_29865,N_29866,N_29867,N_29868,N_29869,N_29870,N_29871,N_29872,N_29873,N_29874,N_29875,N_29876,N_29877,N_29878,N_29879,N_29880,N_29881,N_29882,N_29883,N_29884,N_29885,N_29886,N_29887,N_29888,N_29889,N_29890,N_29891,N_29892,N_29893,N_29894,N_29895,N_29896,N_29897,N_29898,N_29899,N_29900,N_29901,N_29902,N_29903,N_29904,N_29905,N_29906,N_29907,N_29908,N_29909,N_29910,N_29911,N_29912,N_29913,N_29914,N_29915,N_29916,N_29917,N_29918,N_29919,N_29920,N_29921,N_29922,N_29923,N_29924,N_29925,N_29926,N_29927,N_29928,N_29929,N_29930,N_29931,N_29932,N_29933,N_29934,N_29935,N_29936,N_29937,N_29938,N_29939,N_29940,N_29941,N_29942,N_29943,N_29944,N_29945,N_29946,N_29947,N_29948,N_29949,N_29950,N_29951,N_29952,N_29953,N_29954,N_29955,N_29956,N_29957,N_29958,N_29959,N_29960,N_29961,N_29962,N_29963,N_29964,N_29965,N_29966,N_29967,N_29968,N_29969,N_29970,N_29971,N_29972,N_29973,N_29974,N_29975,N_29976,N_29977,N_29978,N_29979,N_29980,N_29981,N_29982,N_29983,N_29984,N_29985,N_29986,N_29987,N_29988,N_29989,N_29990,N_29991,N_29992,N_29993,N_29994,N_29995,N_29996,N_29997,N_29998,N_29999;
nand U0 (N_0,In_1063,In_2316);
nor U1 (N_1,In_734,In_344);
nor U2 (N_2,In_175,In_2974);
or U3 (N_3,In_983,In_1148);
and U4 (N_4,In_1214,In_1766);
xor U5 (N_5,In_1136,In_1315);
nor U6 (N_6,In_1706,In_1058);
and U7 (N_7,In_303,In_261);
nand U8 (N_8,In_598,In_913);
xnor U9 (N_9,In_509,In_2467);
or U10 (N_10,In_721,In_1532);
and U11 (N_11,In_2881,In_274);
or U12 (N_12,In_2038,In_1260);
or U13 (N_13,In_1164,In_1209);
or U14 (N_14,In_2817,In_280);
xnor U15 (N_15,In_2325,In_68);
or U16 (N_16,In_2679,In_1756);
and U17 (N_17,In_2207,In_1339);
and U18 (N_18,In_654,In_2146);
nor U19 (N_19,In_2787,In_1720);
and U20 (N_20,In_2491,In_1911);
or U21 (N_21,In_1506,In_2472);
or U22 (N_22,In_882,In_1326);
or U23 (N_23,In_1057,In_1120);
and U24 (N_24,In_1069,In_2105);
and U25 (N_25,In_1351,In_2774);
nor U26 (N_26,In_403,In_2869);
xnor U27 (N_27,In_948,In_2383);
or U28 (N_28,In_2876,In_318);
nand U29 (N_29,In_376,In_2942);
nand U30 (N_30,In_354,In_250);
and U31 (N_31,In_2367,In_239);
xnor U32 (N_32,In_535,In_1549);
xor U33 (N_33,In_2049,In_1806);
or U34 (N_34,In_2500,In_1561);
or U35 (N_35,In_2470,In_1478);
nor U36 (N_36,In_1086,In_883);
xnor U37 (N_37,In_532,In_304);
nor U38 (N_38,In_2537,In_1305);
xnor U39 (N_39,In_778,In_1262);
xnor U40 (N_40,In_1584,In_2543);
nor U41 (N_41,In_1596,In_185);
and U42 (N_42,In_1735,In_398);
nand U43 (N_43,In_169,In_616);
or U44 (N_44,In_1188,In_2311);
xnor U45 (N_45,In_2551,In_1228);
nor U46 (N_46,In_1275,In_789);
or U47 (N_47,In_1744,In_1662);
and U48 (N_48,In_1490,In_162);
nand U49 (N_49,In_377,In_845);
and U50 (N_50,In_462,In_205);
xor U51 (N_51,In_1107,In_1387);
nand U52 (N_52,In_1933,In_2095);
nand U53 (N_53,In_633,In_1129);
nand U54 (N_54,In_2665,In_1978);
or U55 (N_55,In_97,In_1025);
nand U56 (N_56,In_2141,In_2840);
nor U57 (N_57,In_846,In_2647);
nand U58 (N_58,In_1391,In_2969);
xor U59 (N_59,In_2220,In_2976);
or U60 (N_60,In_459,In_1091);
or U61 (N_61,In_2541,In_70);
xnor U62 (N_62,In_2673,In_47);
nor U63 (N_63,In_14,In_1466);
and U64 (N_64,In_2319,In_1151);
nor U65 (N_65,In_1652,In_257);
xor U66 (N_66,In_2520,In_2119);
and U67 (N_67,In_2033,In_66);
nor U68 (N_68,In_1491,In_379);
nand U69 (N_69,In_2608,In_2504);
and U70 (N_70,In_1861,In_2211);
xor U71 (N_71,In_2852,In_309);
or U72 (N_72,In_2687,In_2180);
nand U73 (N_73,In_1500,In_768);
nand U74 (N_74,In_2641,In_368);
or U75 (N_75,In_1464,In_1527);
and U76 (N_76,In_2431,In_1688);
and U77 (N_77,In_498,In_941);
nor U78 (N_78,In_2567,In_2784);
or U79 (N_79,In_744,In_1656);
and U80 (N_80,In_2129,In_517);
or U81 (N_81,In_78,In_2286);
and U82 (N_82,In_2132,In_876);
nand U83 (N_83,In_1150,In_2920);
nor U84 (N_84,In_1049,In_2587);
and U85 (N_85,In_677,In_2492);
nand U86 (N_86,In_329,In_841);
xor U87 (N_87,In_745,In_2973);
xnor U88 (N_88,In_2084,In_2629);
or U89 (N_89,In_1367,In_936);
nor U90 (N_90,In_1795,In_2499);
and U91 (N_91,In_1725,In_699);
xnor U92 (N_92,In_370,In_1711);
or U93 (N_93,In_2360,In_1841);
or U94 (N_94,In_2203,In_2910);
and U95 (N_95,In_1072,In_1447);
nand U96 (N_96,In_953,In_2911);
nand U97 (N_97,In_1190,In_1891);
or U98 (N_98,In_330,In_1421);
nor U99 (N_99,In_640,In_2464);
nand U100 (N_100,In_2337,In_2953);
nand U101 (N_101,In_1272,In_1699);
nand U102 (N_102,In_2285,In_396);
xor U103 (N_103,In_1436,In_2902);
nand U104 (N_104,In_2389,In_1955);
nor U105 (N_105,In_2638,In_51);
nor U106 (N_106,In_2669,In_1237);
nor U107 (N_107,In_1809,In_1541);
nor U108 (N_108,In_2954,In_1404);
or U109 (N_109,In_1383,In_277);
and U110 (N_110,In_945,In_2844);
and U111 (N_111,In_986,In_2009);
or U112 (N_112,In_541,In_1118);
nor U113 (N_113,In_1292,In_942);
nor U114 (N_114,In_2386,In_2210);
nor U115 (N_115,In_1501,In_534);
or U116 (N_116,In_110,In_2232);
or U117 (N_117,In_1369,In_165);
or U118 (N_118,In_1223,In_1818);
or U119 (N_119,In_2826,In_2403);
or U120 (N_120,In_1299,In_2120);
nor U121 (N_121,In_2922,In_2372);
nor U122 (N_122,In_2768,In_907);
nand U123 (N_123,In_988,In_807);
nand U124 (N_124,In_374,In_1590);
or U125 (N_125,In_2864,In_399);
and U126 (N_126,In_2518,In_1226);
xor U127 (N_127,In_1431,In_1771);
nand U128 (N_128,In_1885,In_1511);
nor U129 (N_129,In_95,In_2865);
or U130 (N_130,In_554,In_2975);
nand U131 (N_131,In_890,In_1265);
or U132 (N_132,In_1378,In_1610);
or U133 (N_133,In_1314,In_2018);
nor U134 (N_134,In_24,In_299);
or U135 (N_135,In_1884,In_2233);
xnor U136 (N_136,In_1277,In_638);
xnor U137 (N_137,In_1241,In_1012);
nand U138 (N_138,In_1496,In_1297);
or U139 (N_139,In_946,In_490);
nand U140 (N_140,In_1040,In_158);
xor U141 (N_141,In_588,In_902);
or U142 (N_142,In_88,In_2730);
nand U143 (N_143,In_2596,In_276);
nand U144 (N_144,In_1445,In_606);
or U145 (N_145,In_2221,In_594);
nand U146 (N_146,In_2880,In_64);
xor U147 (N_147,In_1494,In_2845);
xor U148 (N_148,In_1901,In_1635);
nand U149 (N_149,In_2417,In_877);
nand U150 (N_150,In_521,In_2056);
xor U151 (N_151,In_1046,In_1820);
xor U152 (N_152,In_2732,In_1428);
nor U153 (N_153,In_1888,In_247);
xor U154 (N_154,In_1112,In_2167);
or U155 (N_155,In_2086,In_197);
nand U156 (N_156,In_2259,In_2875);
xor U157 (N_157,In_2628,In_189);
and U158 (N_158,In_925,In_825);
or U159 (N_159,In_591,In_834);
or U160 (N_160,In_2956,In_202);
nor U161 (N_161,In_2040,In_319);
and U162 (N_162,In_1186,In_2078);
nor U163 (N_163,In_1044,In_252);
or U164 (N_164,In_2675,In_823);
or U165 (N_165,In_1092,In_2649);
or U166 (N_166,In_411,In_1218);
and U167 (N_167,In_2388,In_2371);
and U168 (N_168,In_2201,In_2468);
and U169 (N_169,In_451,In_1558);
xnor U170 (N_170,In_672,In_2004);
xor U171 (N_171,In_1626,In_796);
nand U172 (N_172,In_1953,In_1497);
or U173 (N_173,In_1559,In_2404);
or U174 (N_174,In_2835,In_1036);
xnor U175 (N_175,In_2109,In_478);
and U176 (N_176,In_1280,In_2216);
or U177 (N_177,In_424,In_2246);
xnor U178 (N_178,In_1109,In_2446);
xor U179 (N_179,In_214,In_748);
nand U180 (N_180,In_790,In_966);
nor U181 (N_181,In_408,In_2517);
or U182 (N_182,In_328,In_653);
nand U183 (N_183,In_469,In_2939);
or U184 (N_184,In_2174,In_472);
nand U185 (N_185,In_1320,In_1357);
or U186 (N_186,In_1894,In_138);
and U187 (N_187,In_23,In_2071);
nand U188 (N_188,In_2481,In_2171);
and U189 (N_189,In_515,In_2026);
xor U190 (N_190,In_1831,In_2946);
xnor U191 (N_191,In_1971,In_1768);
and U192 (N_192,In_2996,In_1442);
or U193 (N_193,In_1227,In_2525);
nor U194 (N_194,In_1104,In_1270);
nor U195 (N_195,In_50,In_414);
or U196 (N_196,In_493,In_1554);
nand U197 (N_197,In_2798,In_146);
or U198 (N_198,In_1889,In_2432);
or U199 (N_199,In_1616,In_2633);
or U200 (N_200,In_2678,In_1144);
or U201 (N_201,In_15,In_2147);
nand U202 (N_202,In_2346,In_2529);
xor U203 (N_203,In_2979,In_767);
or U204 (N_204,In_2117,In_2001);
and U205 (N_205,In_2428,In_1132);
and U206 (N_206,In_2748,In_413);
nand U207 (N_207,In_73,In_1216);
xnor U208 (N_208,In_2085,In_690);
nor U209 (N_209,In_2200,In_1622);
xor U210 (N_210,In_1195,In_2313);
nor U211 (N_211,In_1974,In_288);
nand U212 (N_212,In_1661,In_2879);
nand U213 (N_213,In_2423,In_1191);
nand U214 (N_214,In_242,In_279);
nand U215 (N_215,In_1068,In_1686);
and U216 (N_216,In_660,In_1225);
nor U217 (N_217,In_1805,In_2029);
and U218 (N_218,In_1987,In_1912);
or U219 (N_219,In_2322,In_1585);
xnor U220 (N_220,In_1370,In_2728);
nor U221 (N_221,In_352,In_1028);
xnor U222 (N_222,In_739,In_1870);
nor U223 (N_223,In_2019,In_839);
nor U224 (N_224,In_580,In_2250);
xnor U225 (N_225,In_1542,In_1406);
nor U226 (N_226,In_1878,In_816);
xor U227 (N_227,In_389,In_234);
nand U228 (N_228,In_2381,In_1991);
and U229 (N_229,In_738,In_2590);
xor U230 (N_230,In_974,In_1762);
and U231 (N_231,In_1834,In_1131);
xor U232 (N_232,In_2960,In_2909);
and U233 (N_233,In_2940,In_1269);
nor U234 (N_234,In_1769,In_2637);
or U235 (N_235,In_2471,In_1951);
and U236 (N_236,In_1738,In_160);
and U237 (N_237,In_1531,In_259);
xor U238 (N_238,In_2610,In_1802);
nor U239 (N_239,In_2581,In_2761);
nor U240 (N_240,In_1772,In_1321);
and U241 (N_241,In_2559,In_1116);
nand U242 (N_242,In_121,In_2205);
nand U243 (N_243,In_1565,In_2931);
nor U244 (N_244,In_2726,In_2343);
xnor U245 (N_245,In_1600,In_2682);
or U246 (N_246,In_429,In_1281);
and U247 (N_247,In_1332,In_523);
nand U248 (N_248,In_2883,In_1976);
nand U249 (N_249,In_1928,In_2476);
nor U250 (N_250,In_1819,In_2062);
or U251 (N_251,In_1651,In_1199);
nand U252 (N_252,In_2429,In_696);
nand U253 (N_253,In_180,In_1390);
and U254 (N_254,In_2734,In_148);
nor U255 (N_255,In_2363,In_1755);
nor U256 (N_256,In_1507,In_2459);
nand U257 (N_257,In_1555,In_249);
nor U258 (N_258,In_2722,In_2992);
and U259 (N_259,In_1108,In_1518);
nor U260 (N_260,In_2712,In_793);
or U261 (N_261,In_1207,In_2306);
xnor U262 (N_262,In_1517,In_168);
or U263 (N_263,In_10,In_1366);
and U264 (N_264,In_1776,In_1854);
xnor U265 (N_265,In_1021,In_106);
nand U266 (N_266,In_648,In_992);
and U267 (N_267,In_775,In_2901);
nor U268 (N_268,In_2701,In_1718);
and U269 (N_269,In_1512,In_2827);
nor U270 (N_270,In_2392,In_1790);
nand U271 (N_271,In_2261,In_2776);
nand U272 (N_272,In_1929,In_1476);
or U273 (N_273,In_2842,In_1015);
or U274 (N_274,In_1485,In_1864);
and U275 (N_275,In_1037,In_1405);
xnor U276 (N_276,In_2928,In_2193);
nand U277 (N_277,In_803,In_1601);
and U278 (N_278,In_2605,In_2767);
and U279 (N_279,In_2082,In_2699);
xnor U280 (N_280,In_550,In_641);
or U281 (N_281,In_2899,In_431);
or U282 (N_282,In_1719,In_963);
nand U283 (N_283,In_1373,In_720);
nand U284 (N_284,In_1473,In_1903);
or U285 (N_285,In_72,In_186);
and U286 (N_286,In_1570,In_391);
xnor U287 (N_287,In_642,In_1106);
or U288 (N_288,In_1668,In_2349);
and U289 (N_289,In_2506,In_2290);
xnor U290 (N_290,In_693,In_780);
nand U291 (N_291,In_1372,In_1381);
nor U292 (N_292,In_1073,In_112);
or U293 (N_293,In_76,In_2716);
nand U294 (N_294,In_382,In_2900);
or U295 (N_295,In_2690,In_2568);
nand U296 (N_296,In_2718,In_801);
xor U297 (N_297,In_1973,In_2868);
nand U298 (N_298,In_1710,In_976);
or U299 (N_299,In_1580,In_1060);
or U300 (N_300,In_1777,In_322);
nor U301 (N_301,In_838,In_871);
nand U302 (N_302,In_500,In_1982);
nor U303 (N_303,In_385,In_1403);
nor U304 (N_304,In_2652,In_967);
nor U305 (N_305,In_1014,In_2962);
xor U306 (N_306,In_2195,In_1866);
xnor U307 (N_307,In_1308,In_982);
and U308 (N_308,In_2789,In_1963);
nand U309 (N_309,In_1510,In_2746);
or U310 (N_310,In_2762,In_140);
and U311 (N_311,In_2618,In_784);
or U312 (N_312,In_157,In_1232);
xor U313 (N_313,In_1968,In_474);
nor U314 (N_314,In_114,In_2448);
and U315 (N_315,In_1847,In_2816);
nand U316 (N_316,In_2943,In_624);
and U317 (N_317,In_1171,In_962);
xor U318 (N_318,In_1750,In_19);
nor U319 (N_319,In_2172,In_91);
or U320 (N_320,In_2878,In_390);
or U321 (N_321,In_448,In_903);
and U322 (N_322,In_2870,In_901);
or U323 (N_323,In_2562,In_1443);
xor U324 (N_324,In_1258,In_358);
and U325 (N_325,In_2676,In_2775);
and U326 (N_326,In_2588,In_866);
xnor U327 (N_327,In_446,In_1999);
nor U328 (N_328,In_533,In_2867);
or U329 (N_329,In_199,In_1508);
xor U330 (N_330,In_1293,In_755);
and U331 (N_331,In_2528,In_1222);
and U332 (N_332,In_2489,In_1677);
and U333 (N_333,In_545,In_237);
and U334 (N_334,In_2823,In_2963);
and U335 (N_335,In_269,In_2530);
or U336 (N_336,In_1504,In_881);
nand U337 (N_337,In_2107,In_880);
nor U338 (N_338,In_1594,In_1757);
and U339 (N_339,In_1615,In_501);
nand U340 (N_340,In_814,In_1213);
xor U341 (N_341,In_868,In_2955);
xor U342 (N_342,In_1763,In_1264);
or U343 (N_343,In_2779,In_392);
xor U344 (N_344,In_2563,In_466);
nand U345 (N_345,In_2653,In_644);
and U346 (N_346,In_2917,In_566);
nand U347 (N_347,In_2104,In_294);
or U348 (N_348,In_1001,In_2100);
or U349 (N_349,In_1427,In_1456);
or U350 (N_350,In_1923,In_2044);
or U351 (N_351,In_578,In_235);
and U352 (N_352,In_1915,In_656);
and U353 (N_353,In_2416,In_2438);
nor U354 (N_354,In_286,In_916);
xor U355 (N_355,In_2260,In_2958);
nor U356 (N_356,In_952,In_2137);
and U357 (N_357,In_1238,In_850);
xor U358 (N_358,In_577,In_1880);
or U359 (N_359,In_1306,In_1682);
or U360 (N_360,In_1145,In_464);
and U361 (N_361,In_456,In_2079);
nor U362 (N_362,In_334,In_2197);
and U363 (N_363,In_2967,In_2390);
nor U364 (N_364,In_2045,In_2231);
and U365 (N_365,In_1530,In_774);
nor U366 (N_366,In_2815,In_1231);
nor U367 (N_367,In_21,In_2312);
nand U368 (N_368,In_1630,In_1325);
or U369 (N_369,In_253,In_1817);
and U370 (N_370,In_460,In_912);
or U371 (N_371,In_336,In_1922);
nand U372 (N_372,In_342,In_1965);
or U373 (N_373,In_2185,In_2834);
nor U374 (N_374,In_1417,In_1789);
nand U375 (N_375,In_1949,In_57);
xnor U376 (N_376,In_1563,In_2335);
and U377 (N_377,In_2277,In_461);
or U378 (N_378,In_1128,In_316);
or U379 (N_379,In_1743,In_1051);
and U380 (N_380,In_1869,In_833);
nand U381 (N_381,In_2700,In_2592);
xor U382 (N_382,In_959,In_2188);
xnor U383 (N_383,In_2849,In_2643);
xor U384 (N_384,In_2096,In_2614);
and U385 (N_385,In_1862,In_2198);
or U386 (N_386,In_2184,In_2378);
and U387 (N_387,In_2764,In_958);
nor U388 (N_388,In_2450,In_1647);
xnor U389 (N_389,In_482,In_102);
and U390 (N_390,In_476,In_1583);
and U391 (N_391,In_409,In_206);
nand U392 (N_392,In_2498,In_373);
or U393 (N_393,In_92,In_2664);
nor U394 (N_394,In_2660,In_1451);
xor U395 (N_395,In_2579,In_701);
nor U396 (N_396,In_2304,In_998);
xor U397 (N_397,In_2978,In_607);
nand U398 (N_398,In_593,In_703);
nor U399 (N_399,In_1572,In_1248);
or U400 (N_400,In_1838,In_265);
nand U401 (N_401,In_119,In_1502);
or U402 (N_402,In_1863,In_2624);
nor U403 (N_403,In_2366,In_2175);
xnor U404 (N_404,In_2023,In_512);
or U405 (N_405,In_255,In_2801);
nor U406 (N_406,In_1745,In_1539);
nor U407 (N_407,In_405,In_531);
and U408 (N_408,In_273,In_1059);
and U409 (N_409,In_2075,In_2570);
xor U410 (N_410,In_126,In_233);
and U411 (N_411,In_2797,In_692);
xnor U412 (N_412,In_1544,In_2670);
nand U413 (N_413,In_1048,In_161);
or U414 (N_414,In_989,In_2650);
nor U415 (N_415,In_2756,In_495);
xnor U416 (N_416,In_1620,In_762);
nand U417 (N_417,In_52,In_527);
and U418 (N_418,In_1110,In_2218);
or U419 (N_419,In_950,In_486);
xnor U420 (N_420,In_1545,In_1930);
and U421 (N_421,In_387,In_842);
or U422 (N_422,In_2161,In_2921);
and U423 (N_423,In_2600,In_951);
nor U424 (N_424,In_2727,In_212);
nor U425 (N_425,In_1606,In_179);
xnor U426 (N_426,In_216,In_1007);
and U427 (N_427,In_1200,In_1422);
nand U428 (N_428,In_2703,In_826);
and U429 (N_429,In_182,In_2139);
or U430 (N_430,In_1139,In_568);
or U431 (N_431,In_1039,In_605);
or U432 (N_432,In_1279,In_1934);
and U433 (N_433,In_260,In_1440);
and U434 (N_434,In_1944,In_422);
nand U435 (N_435,In_1437,In_2786);
and U436 (N_436,In_2452,In_2630);
xnor U437 (N_437,In_1017,In_1727);
nand U438 (N_438,In_150,In_196);
and U439 (N_439,In_837,In_1230);
xnor U440 (N_440,In_135,In_2495);
nand U441 (N_441,In_1977,In_315);
or U442 (N_442,In_1618,In_815);
and U443 (N_443,In_2571,In_2987);
or U444 (N_444,In_911,In_940);
xnor U445 (N_445,In_1848,In_2150);
nand U446 (N_446,In_943,In_266);
xor U447 (N_447,In_193,In_1851);
and U448 (N_448,In_1288,In_2951);
nand U449 (N_449,In_1660,In_1240);
or U450 (N_450,In_74,In_442);
xor U451 (N_451,In_87,In_1849);
nand U452 (N_452,In_1206,In_483);
or U453 (N_453,In_2003,In_1474);
or U454 (N_454,In_2811,In_1716);
and U455 (N_455,In_516,In_610);
and U456 (N_456,In_1683,In_2487);
nand U457 (N_457,In_697,In_107);
xor U458 (N_458,In_1815,In_599);
nand U459 (N_459,In_1193,In_449);
nor U460 (N_460,In_1882,In_708);
xor U461 (N_461,In_510,In_1639);
nand U462 (N_462,In_302,In_2);
nor U463 (N_463,In_1992,In_1245);
or U464 (N_464,In_810,In_11);
or U465 (N_465,In_2534,In_1311);
nand U466 (N_466,In_1198,In_1503);
or U467 (N_467,In_2451,In_879);
and U468 (N_468,In_450,In_1407);
and U469 (N_469,In_2245,In_1273);
xor U470 (N_470,In_455,In_2461);
xor U471 (N_471,In_2602,In_2463);
nand U472 (N_472,In_2948,In_975);
nor U473 (N_473,In_2419,In_675);
nand U474 (N_474,In_1548,In_2434);
nor U475 (N_475,In_2279,In_105);
nor U476 (N_476,In_181,In_1868);
and U477 (N_477,In_960,In_2607);
nor U478 (N_478,In_2315,In_2671);
nand U479 (N_479,In_1450,In_108);
nand U480 (N_480,In_2225,In_812);
nand U481 (N_481,In_362,In_34);
nor U482 (N_482,In_1410,In_127);
nand U483 (N_483,In_2620,In_1543);
or U484 (N_484,In_2183,In_932);
nor U485 (N_485,In_740,In_2101);
or U486 (N_486,In_2409,In_1065);
xnor U487 (N_487,In_49,In_520);
nand U488 (N_488,In_2380,In_2138);
xnor U489 (N_489,In_156,In_864);
xnor U490 (N_490,In_93,In_673);
nand U491 (N_491,In_558,In_1394);
nor U492 (N_492,In_792,In_2674);
or U493 (N_493,In_1879,In_592);
nor U494 (N_494,In_2621,In_467);
nand U495 (N_495,In_1364,In_54);
and U496 (N_496,In_2165,In_1631);
or U497 (N_497,In_1823,In_731);
nand U498 (N_498,In_1114,In_629);
xor U499 (N_499,In_1337,In_1778);
nand U500 (N_500,In_104,In_1233);
xor U501 (N_501,In_103,In_1016);
or U502 (N_502,In_1204,In_2970);
or U503 (N_503,In_1788,In_2039);
xnor U504 (N_504,In_1993,In_2333);
nor U505 (N_505,In_928,In_1439);
nor U506 (N_506,In_2267,In_2812);
nor U507 (N_507,In_1876,In_1759);
nand U508 (N_508,In_2024,In_1064);
or U509 (N_509,In_1829,In_529);
nand U510 (N_510,In_659,In_1873);
and U511 (N_511,In_2299,In_458);
nor U512 (N_512,In_321,In_781);
and U513 (N_513,In_1463,In_1538);
or U514 (N_514,In_1843,In_1411);
and U515 (N_515,In_2572,In_477);
or U516 (N_516,In_345,In_711);
xor U517 (N_517,In_918,In_1988);
nor U518 (N_518,In_1493,In_2251);
nand U519 (N_519,In_1197,In_1617);
xnor U520 (N_520,In_1083,In_2426);
xor U521 (N_521,In_122,In_381);
nand U522 (N_522,In_2412,In_923);
nand U523 (N_523,In_1871,In_1737);
and U524 (N_524,In_1027,In_1085);
xor U525 (N_525,In_2187,In_586);
xnor U526 (N_526,In_2391,In_1989);
xor U527 (N_527,In_285,In_1327);
xor U528 (N_528,In_1604,In_2968);
or U529 (N_529,In_2905,In_2912);
nor U530 (N_530,In_45,In_2855);
and U531 (N_531,In_1035,In_1282);
nand U532 (N_532,In_2566,In_1773);
or U533 (N_533,In_1636,In_1966);
nor U534 (N_534,In_899,In_2192);
and U535 (N_535,In_2625,In_832);
and U536 (N_536,In_2918,In_2526);
and U537 (N_537,In_1628,In_650);
xnor U538 (N_538,In_2351,In_678);
nand U539 (N_539,In_2914,In_546);
or U540 (N_540,In_183,In_2007);
or U541 (N_541,In_278,In_990);
and U542 (N_542,In_2757,In_1298);
nand U543 (N_543,In_2418,In_2224);
xor U544 (N_544,In_1938,In_281);
nand U545 (N_545,In_949,In_2384);
or U546 (N_546,In_601,In_84);
nor U547 (N_547,In_904,In_1033);
nor U548 (N_548,In_741,In_195);
nor U549 (N_549,In_2106,In_1576);
xor U550 (N_550,In_2750,In_82);
nand U551 (N_551,In_1892,In_0);
or U552 (N_552,In_2374,In_802);
nand U553 (N_553,In_2656,In_219);
or U554 (N_554,In_83,In_2799);
nor U555 (N_555,In_2689,In_2000);
or U556 (N_556,In_1467,In_134);
and U557 (N_557,In_2846,In_2809);
or U558 (N_558,In_1056,In_427);
nand U559 (N_559,In_1632,In_1430);
nand U560 (N_560,In_2169,In_773);
nor U561 (N_561,In_1157,In_2505);
and U562 (N_562,In_2736,In_898);
or U563 (N_563,In_1368,In_715);
nand U564 (N_564,In_822,In_1452);
or U565 (N_565,In_1874,In_496);
xor U566 (N_566,In_479,In_1495);
xor U567 (N_567,In_1126,In_1123);
nor U568 (N_568,In_1638,In_324);
or U569 (N_569,In_2058,In_2601);
nor U570 (N_570,In_1593,In_263);
xor U571 (N_571,In_1920,In_2108);
nand U572 (N_572,In_2522,In_1498);
nor U573 (N_573,In_2861,In_2832);
and U574 (N_574,In_2222,In_2124);
or U575 (N_575,In_978,In_1424);
nand U576 (N_576,In_1105,In_2773);
nor U577 (N_577,In_2950,In_480);
nand U578 (N_578,In_2615,In_2995);
and U579 (N_579,In_2668,In_1980);
or U580 (N_580,In_538,In_1837);
nor U581 (N_581,In_2408,In_2099);
nor U582 (N_582,In_1627,In_583);
nor U583 (N_583,In_2469,In_349);
or U584 (N_584,In_1811,In_96);
xor U585 (N_585,In_124,In_2145);
or U586 (N_586,In_2329,In_2342);
nand U587 (N_587,In_702,In_808);
xor U588 (N_588,In_1170,In_716);
xor U589 (N_589,In_1154,In_632);
xor U590 (N_590,In_2792,In_1990);
nor U591 (N_591,In_2291,In_2743);
or U592 (N_592,In_2064,In_671);
xnor U593 (N_593,In_441,In_39);
nor U594 (N_594,In_2347,In_2613);
nor U595 (N_595,In_1098,In_2475);
xor U596 (N_596,In_914,In_2751);
and U597 (N_597,In_1916,In_2088);
xnor U598 (N_598,In_1899,In_86);
nor U599 (N_599,In_2176,In_417);
nor U600 (N_600,In_1675,In_2663);
nand U601 (N_601,In_1551,In_2345);
nand U602 (N_602,In_981,In_1746);
or U603 (N_603,In_177,In_2720);
or U604 (N_604,In_1857,In_29);
nor U605 (N_605,In_727,In_1352);
xnor U606 (N_606,In_2655,In_1774);
nand U607 (N_607,In_2723,In_754);
nor U608 (N_608,In_524,In_1972);
xor U609 (N_609,In_2453,In_1441);
nor U610 (N_610,In_2331,In_1330);
or U611 (N_611,In_1896,In_2357);
or U612 (N_612,In_2385,In_753);
xnor U613 (N_613,In_2479,In_2097);
nand U614 (N_614,In_765,In_1887);
and U615 (N_615,In_651,In_2999);
nor U616 (N_616,In_2406,In_835);
xnor U617 (N_617,In_1042,In_282);
nor U618 (N_618,In_1302,In_761);
and U619 (N_619,In_2903,In_1521);
and U620 (N_620,In_1676,In_2893);
xnor U621 (N_621,In_2112,In_2405);
nor U622 (N_622,In_785,In_622);
and U623 (N_623,In_2377,In_2511);
or U624 (N_624,In_730,In_661);
nor U625 (N_625,In_1350,In_468);
nor U626 (N_626,In_1961,In_271);
and U627 (N_627,In_170,In_2254);
nor U628 (N_628,In_2041,In_2046);
nand U629 (N_629,In_631,In_1178);
xor U630 (N_630,In_1099,In_2436);
and U631 (N_631,In_1180,In_2415);
nand U632 (N_632,In_378,In_2081);
nor U633 (N_633,In_2208,In_1655);
and U634 (N_634,In_1687,In_2819);
and U635 (N_635,In_840,In_722);
or U636 (N_636,In_2350,In_1334);
xor U637 (N_637,In_1113,In_862);
nor U638 (N_638,In_669,In_2034);
nand U639 (N_639,In_574,In_2140);
nand U640 (N_640,In_1125,In_2617);
xnor U641 (N_641,In_867,In_312);
or U642 (N_642,In_2164,In_1022);
nand U643 (N_643,In_1026,In_1751);
nand U644 (N_644,In_2072,In_1254);
nor U645 (N_645,In_2810,In_471);
nand U646 (N_646,In_2194,In_2092);
xnor U647 (N_647,In_1850,In_1294);
xor U648 (N_648,In_2407,In_1904);
nor U649 (N_649,In_1426,In_1336);
nand U650 (N_650,In_526,In_2843);
or U651 (N_651,In_1122,In_2556);
and U652 (N_652,In_1183,In_555);
nand U653 (N_653,In_2413,In_2848);
or U654 (N_654,In_1006,In_1797);
nand U655 (N_655,In_2318,In_475);
xnor U656 (N_656,In_445,In_2708);
nor U657 (N_657,In_1019,In_2089);
or U658 (N_658,In_2622,In_1010);
or U659 (N_659,In_668,In_1182);
and U660 (N_660,In_1300,In_2802);
nor U661 (N_661,In_2308,In_724);
or U662 (N_662,In_619,In_2394);
or U663 (N_663,In_1749,In_2509);
and U664 (N_664,In_1986,In_2851);
xnor U665 (N_665,In_1925,In_2593);
nor U666 (N_666,In_2430,In_2991);
or U667 (N_667,In_174,In_1663);
nor U668 (N_668,In_972,In_2281);
and U669 (N_669,In_971,In_2484);
nor U670 (N_670,In_736,In_1697);
nor U671 (N_671,In_1004,In_2118);
nor U672 (N_672,In_709,In_1828);
xnor U673 (N_673,In_149,In_2527);
or U674 (N_674,In_2294,In_2603);
nand U675 (N_675,In_1097,In_691);
xnor U676 (N_676,In_2441,In_797);
nor U677 (N_677,In_1244,In_828);
and U678 (N_678,In_2536,In_2466);
nand U679 (N_679,In_2793,In_844);
or U680 (N_680,In_2264,In_908);
and U681 (N_681,In_1758,In_94);
and U682 (N_682,In_2589,In_848);
xnor U683 (N_683,In_28,In_2070);
and U684 (N_684,In_872,In_2295);
or U685 (N_685,In_20,In_2402);
nor U686 (N_686,In_2936,In_917);
nand U687 (N_687,In_2825,In_2744);
nand U688 (N_688,In_1172,In_2111);
xnor U689 (N_689,In_133,In_1415);
nand U690 (N_690,In_1898,In_1781);
nor U691 (N_691,In_1712,In_836);
or U692 (N_692,In_1935,In_275);
nand U693 (N_693,In_537,In_2783);
nand U694 (N_694,In_2159,In_993);
nand U695 (N_695,In_652,In_1557);
nor U696 (N_696,In_65,In_2008);
xnor U697 (N_697,In_291,In_9);
nor U698 (N_698,In_16,In_970);
xnor U699 (N_699,In_1657,In_2396);
and U700 (N_700,In_886,In_1516);
nor U701 (N_701,In_2606,In_432);
and U702 (N_702,In_926,In_1061);
nand U703 (N_703,In_2609,In_1525);
nand U704 (N_704,In_743,In_2710);
and U705 (N_705,In_2387,In_1475);
or U706 (N_706,In_1534,In_1678);
nor U707 (N_707,In_221,In_1053);
nand U708 (N_708,In_264,In_726);
and U709 (N_709,In_1169,In_357);
nor U710 (N_710,In_2523,In_2257);
and U711 (N_711,In_1247,In_2493);
or U712 (N_712,In_2302,In_2356);
and U713 (N_713,In_2163,In_1645);
nand U714 (N_714,In_646,In_1846);
or U715 (N_715,In_2874,In_1842);
xnor U716 (N_716,In_530,In_2375);
xnor U717 (N_717,In_2740,In_2841);
and U718 (N_718,In_2754,In_1023);
or U719 (N_719,In_2888,In_437);
nor U720 (N_720,In_2646,In_1358);
nand U721 (N_721,In_2204,In_1833);
or U722 (N_722,In_1301,In_782);
and U723 (N_723,In_704,In_1634);
or U724 (N_724,In_1801,In_2866);
nor U725 (N_725,In_2611,In_503);
and U726 (N_726,In_1536,In_2667);
xor U727 (N_727,In_1844,In_2985);
nand U728 (N_728,In_2227,In_2927);
or U729 (N_729,In_1924,In_1361);
nand U730 (N_730,In_340,In_2818);
xnor U731 (N_731,In_1276,In_443);
nor U732 (N_732,In_2065,In_2283);
nor U733 (N_733,In_2573,In_305);
or U734 (N_734,In_1087,In_2830);
and U735 (N_735,In_1783,In_1219);
or U736 (N_736,In_1124,In_1926);
nand U737 (N_737,In_1138,In_1075);
or U738 (N_738,In_2994,In_1767);
nand U739 (N_739,In_536,In_572);
xor U740 (N_740,In_2494,In_2324);
nor U741 (N_741,In_1581,In_217);
xor U742 (N_742,In_2115,In_2437);
nor U743 (N_743,In_705,In_756);
xnor U744 (N_744,In_2980,In_1080);
nand U745 (N_745,In_1942,In_2482);
or U746 (N_746,In_1724,In_2585);
nor U747 (N_747,In_297,In_1459);
and U748 (N_748,In_2275,In_1356);
or U749 (N_749,In_1623,In_1840);
nand U750 (N_750,In_1142,In_53);
or U751 (N_751,In_2552,In_1353);
or U752 (N_752,In_262,In_2486);
and U753 (N_753,In_2270,In_548);
nand U754 (N_754,In_769,In_1155);
nor U755 (N_755,In_1748,In_2560);
nand U756 (N_756,In_895,In_1111);
xnor U757 (N_757,In_805,In_2733);
xnor U758 (N_758,In_1030,In_994);
or U759 (N_759,In_1246,In_2361);
and U760 (N_760,In_1786,In_1723);
and U761 (N_761,In_2713,In_1287);
nor U762 (N_762,In_2747,In_6);
and U763 (N_763,In_2262,In_1796);
xnor U764 (N_764,In_1519,In_1644);
nor U765 (N_765,In_938,In_2131);
and U766 (N_766,In_1076,In_1201);
nor U767 (N_767,In_3,In_999);
nand U768 (N_768,In_2300,In_1734);
nand U769 (N_769,In_2238,In_934);
and U770 (N_770,In_2444,In_395);
nor U771 (N_771,In_2144,In_61);
and U772 (N_772,In_1067,In_980);
nor U773 (N_773,In_270,In_885);
nand U774 (N_774,In_2578,In_245);
nor U775 (N_775,In_2715,In_1483);
xor U776 (N_776,In_1089,In_4);
or U777 (N_777,In_1567,In_2202);
nand U778 (N_778,In_870,In_1444);
xor U779 (N_779,In_1382,In_1696);
or U780 (N_780,In_90,In_1741);
nand U781 (N_781,In_732,In_2457);
nor U782 (N_782,In_300,In_681);
and U783 (N_783,In_2604,In_1189);
xor U784 (N_784,In_436,In_2632);
nand U785 (N_785,In_2162,In_770);
or U786 (N_786,In_1927,In_2640);
nor U787 (N_787,In_1414,In_2938);
nor U788 (N_788,In_2032,In_1344);
xor U789 (N_789,In_98,In_920);
xnor U790 (N_790,In_2237,In_1401);
nor U791 (N_791,In_227,In_597);
and U792 (N_792,In_2020,In_1956);
nand U793 (N_793,In_1454,In_2066);
nor U794 (N_794,In_2691,In_1329);
xnor U795 (N_795,In_204,In_1477);
xor U796 (N_796,In_1520,In_2158);
nand U797 (N_797,In_987,In_1392);
or U798 (N_798,In_2891,In_42);
or U799 (N_799,In_1274,In_636);
nor U800 (N_800,In_1316,In_2997);
nor U801 (N_801,In_2545,In_426);
nor U802 (N_802,In_1453,In_386);
xnor U803 (N_803,In_626,In_1959);
nor U804 (N_804,In_2926,In_338);
or U805 (N_805,In_1692,In_1054);
nand U806 (N_806,In_1304,In_2871);
nor U807 (N_807,In_1236,In_2886);
nor U808 (N_808,In_924,In_2772);
nand U809 (N_809,In_609,In_939);
or U810 (N_810,In_1996,In_1094);
xnor U811 (N_811,In_2447,In_2895);
nand U812 (N_812,In_438,In_688);
nor U813 (N_813,In_404,In_1185);
nor U814 (N_814,In_2885,In_1005);
or U815 (N_815,In_1673,In_1179);
xor U816 (N_816,In_2373,In_2941);
xnor U817 (N_817,In_1156,In_2714);
nand U818 (N_818,In_1785,In_167);
and U819 (N_819,In_1658,In_576);
nor U820 (N_820,In_420,In_184);
xnor U821 (N_821,In_2731,In_1962);
and U822 (N_822,In_2327,In_2341);
xor U823 (N_823,In_821,In_2051);
nand U824 (N_824,In_1793,In_1573);
or U825 (N_825,In_1333,In_1761);
xor U826 (N_826,In_685,In_1814);
and U827 (N_827,In_284,In_713);
nor U828 (N_828,In_518,In_2658);
nor U829 (N_829,In_2364,In_2925);
xor U830 (N_830,In_508,In_410);
nand U831 (N_831,In_1167,In_2239);
nand U832 (N_832,In_1166,In_528);
or U833 (N_833,In_1220,In_2666);
nor U834 (N_834,In_2945,In_1672);
nor U835 (N_835,In_827,In_2685);
or U836 (N_836,In_440,In_718);
or U837 (N_837,In_1434,In_1659);
or U838 (N_838,In_2036,In_2847);
nand U839 (N_839,In_2196,In_2577);
or U840 (N_840,In_2533,In_388);
nand U841 (N_841,In_905,In_552);
nand U842 (N_842,In_1133,In_2707);
nand U843 (N_843,In_1479,In_2554);
and U844 (N_844,In_2397,In_423);
and U845 (N_845,In_359,In_151);
nor U846 (N_846,In_2719,In_2217);
nor U847 (N_847,In_1649,In_612);
and U848 (N_848,In_571,In_2770);
and U849 (N_849,In_847,In_758);
nand U850 (N_850,In_2094,In_1008);
nand U851 (N_851,In_56,In_1695);
nand U852 (N_852,In_930,In_1402);
and U853 (N_853,In_1140,In_1432);
nand U854 (N_854,In_1203,In_2794);
and U855 (N_855,In_806,In_1438);
or U856 (N_856,In_2929,In_1998);
and U857 (N_857,In_2323,In_2272);
or U858 (N_858,In_30,In_2516);
nor U859 (N_859,In_706,In_2133);
or U860 (N_860,In_1130,In_463);
nor U861 (N_861,In_979,In_365);
and U862 (N_862,In_2821,In_412);
or U863 (N_863,In_63,In_2686);
and U864 (N_864,In_1897,In_2873);
or U865 (N_865,In_1782,In_628);
xnor U866 (N_866,In_2644,In_2288);
nor U867 (N_867,In_851,In_2937);
nor U868 (N_868,In_2269,In_2028);
nand U869 (N_869,In_1564,In_2508);
nand U870 (N_870,In_1066,In_1845);
xor U871 (N_871,In_1967,In_751);
nand U872 (N_872,In_1217,In_1587);
or U873 (N_873,In_564,In_491);
xor U874 (N_874,In_1484,In_620);
and U875 (N_875,In_1633,In_1640);
and U876 (N_876,In_906,In_2877);
and U877 (N_877,In_1798,In_2068);
xor U878 (N_878,In_915,In_131);
xnor U879 (N_879,In_1090,In_2753);
nand U880 (N_880,In_788,In_2053);
or U881 (N_881,In_2642,In_707);
nand U882 (N_882,In_1286,In_1794);
nand U883 (N_883,In_858,In_984);
nor U884 (N_884,In_2173,In_137);
and U885 (N_885,In_335,In_350);
xor U886 (N_886,In_2293,In_2755);
or U887 (N_887,In_2704,In_1386);
or U888 (N_888,In_2376,In_2340);
nand U889 (N_889,In_2199,In_2083);
or U890 (N_890,In_854,In_2659);
and U891 (N_891,In_2328,In_2136);
and U892 (N_892,In_2546,In_559);
nand U893 (N_893,In_2694,In_2683);
and U894 (N_894,In_585,In_191);
or U895 (N_895,In_1009,In_320);
or U896 (N_896,In_2368,In_1921);
nor U897 (N_897,In_817,In_549);
nor U898 (N_898,In_1760,In_614);
or U899 (N_899,In_2777,In_337);
nand U900 (N_900,In_771,In_1940);
nor U901 (N_901,In_1586,In_1084);
nor U902 (N_902,In_613,In_2355);
or U903 (N_903,In_2263,In_1446);
xnor U904 (N_904,In_2206,In_1900);
xnor U905 (N_905,In_2025,In_595);
or U906 (N_906,In_236,In_2307);
or U907 (N_907,In_2829,In_779);
nand U908 (N_908,In_1,In_384);
or U909 (N_909,In_366,In_1400);
nor U910 (N_910,In_1611,In_791);
nor U911 (N_911,In_1077,In_1624);
and U912 (N_912,In_447,In_874);
or U913 (N_913,In_117,In_2574);
nor U914 (N_914,In_2977,In_5);
or U915 (N_915,In_2422,In_968);
nor U916 (N_916,In_46,In_1680);
nand U917 (N_917,In_267,In_1803);
nor U918 (N_918,In_2102,In_1176);
or U919 (N_919,In_364,In_215);
nor U920 (N_920,In_60,In_2544);
and U921 (N_921,In_2153,In_857);
xor U922 (N_922,In_153,In_2542);
nand U923 (N_923,In_1713,In_747);
xnor U924 (N_924,In_1621,In_944);
and U925 (N_925,In_166,In_2594);
nand U926 (N_926,In_1465,In_2555);
xnor U927 (N_927,In_211,In_1376);
nor U928 (N_928,In_2090,In_7);
nor U929 (N_929,In_1418,In_1826);
nor U930 (N_930,In_1552,In_1115);
or U931 (N_931,In_1165,In_2828);
xnor U932 (N_932,In_1210,In_2539);
nand U933 (N_933,In_2961,In_1338);
or U934 (N_934,In_2990,In_2330);
nand U935 (N_935,In_228,In_1412);
and U936 (N_936,In_813,In_1654);
xnor U937 (N_937,In_2060,In_1175);
or U938 (N_938,In_1261,In_85);
and U939 (N_939,In_2804,In_218);
nand U940 (N_940,In_2742,In_666);
and U941 (N_941,In_2882,In_1571);
xnor U942 (N_942,In_164,In_58);
or U943 (N_943,In_415,In_1486);
xnor U944 (N_944,In_254,In_1679);
nor U945 (N_945,In_1704,In_1540);
xor U946 (N_946,In_658,In_772);
and U947 (N_947,In_856,In_2709);
or U948 (N_948,In_794,In_2872);
nor U949 (N_949,In_1229,In_1689);
or U950 (N_950,In_2634,In_2395);
nor U951 (N_951,In_565,In_327);
and U952 (N_952,In_2284,In_2182);
xnor U953 (N_953,In_2993,In_596);
nand U954 (N_954,In_289,In_418);
or U955 (N_955,In_208,In_1102);
xnor U956 (N_956,In_1345,In_852);
xnor U957 (N_957,In_602,In_1824);
and U958 (N_958,In_109,In_283);
nor U959 (N_959,In_553,In_2440);
nand U960 (N_960,In_143,In_1560);
nand U961 (N_961,In_2110,In_2549);
or U962 (N_962,In_1174,In_492);
nand U963 (N_963,In_2739,In_798);
xnor U964 (N_964,In_1285,In_2344);
nor U965 (N_965,In_1328,In_1480);
nor U966 (N_966,In_682,In_2091);
nand U967 (N_967,In_2116,In_2935);
nand U968 (N_968,In_1419,In_125);
nor U969 (N_969,In_1290,In_1832);
nand U970 (N_970,In_136,In_2473);
and U971 (N_971,In_1574,In_985);
or U972 (N_972,In_525,In_1941);
nand U973 (N_973,In_1984,In_2688);
and U974 (N_974,In_820,In_2988);
and U975 (N_975,In_194,In_1614);
nor U976 (N_976,In_1162,In_897);
or U977 (N_977,In_670,In_2693);
nor U978 (N_978,In_1257,In_742);
xnor U979 (N_979,In_1855,In_2011);
nor U980 (N_980,In_2309,In_12);
nand U981 (N_981,In_2785,In_2760);
nand U982 (N_982,In_2399,In_1839);
or U983 (N_983,In_2310,In_2897);
or U984 (N_984,In_2265,In_246);
and U985 (N_985,In_2765,In_1469);
and U986 (N_986,In_1095,In_2662);
nand U987 (N_987,In_2780,In_1249);
nand U988 (N_988,In_1018,In_2805);
nand U989 (N_989,In_200,In_1011);
and U990 (N_990,In_2822,In_2488);
and U991 (N_991,In_1578,In_1943);
nor U992 (N_992,In_2352,In_1457);
nand U993 (N_993,In_2547,In_251);
xor U994 (N_994,In_1371,In_400);
xnor U995 (N_995,In_878,In_1255);
xnor U996 (N_996,In_1666,In_665);
and U997 (N_997,In_725,In_737);
nand U998 (N_998,In_100,In_2063);
nor U999 (N_999,In_1733,In_2278);
nor U1000 (N_1000,In_1690,N_641);
nand U1001 (N_1001,N_121,N_450);
and U1002 (N_1002,In_2680,N_271);
and U1003 (N_1003,N_474,In_543);
and U1004 (N_1004,N_940,In_575);
xnor U1005 (N_1005,In_1821,In_2711);
nand U1006 (N_1006,N_930,N_880);
or U1007 (N_1007,N_756,N_511);
nor U1008 (N_1008,In_111,N_156);
nor U1009 (N_1009,In_799,In_2243);
nand U1010 (N_1010,N_19,In_290);
xor U1011 (N_1011,In_1267,N_43);
or U1012 (N_1012,N_825,In_393);
nand U1013 (N_1013,In_2209,N_15);
nor U1014 (N_1014,In_723,In_1860);
xnor U1015 (N_1015,In_973,In_1705);
xnor U1016 (N_1016,In_1078,In_2771);
nand U1017 (N_1017,In_2795,In_957);
xor U1018 (N_1018,In_2896,N_447);
nand U1019 (N_1019,N_349,N_864);
xnor U1020 (N_1020,N_589,N_369);
or U1021 (N_1021,N_766,N_128);
and U1022 (N_1022,In_947,In_617);
xor U1023 (N_1023,In_689,In_1598);
xor U1024 (N_1024,In_2465,In_749);
xnor U1025 (N_1025,In_1134,In_714);
and U1026 (N_1026,In_884,N_431);
and U1027 (N_1027,In_2098,N_329);
xor U1028 (N_1028,N_427,N_300);
xor U1029 (N_1029,N_197,N_762);
or U1030 (N_1030,In_910,In_2122);
or U1031 (N_1031,N_367,N_280);
nand U1032 (N_1032,In_1529,In_369);
nor U1033 (N_1033,In_573,N_21);
xnor U1034 (N_1034,In_2510,N_335);
nor U1035 (N_1035,In_226,In_615);
and U1036 (N_1036,In_2166,In_657);
or U1037 (N_1037,N_304,In_1492);
nor U1038 (N_1038,In_1359,In_1591);
nor U1039 (N_1039,N_494,In_2887);
or U1040 (N_1040,N_807,In_1295);
nor U1041 (N_1041,In_323,In_2439);
or U1042 (N_1042,In_2514,N_153);
nor U1043 (N_1043,N_122,N_316);
xnor U1044 (N_1044,N_261,N_516);
xor U1045 (N_1045,N_902,N_913);
and U1046 (N_1046,N_654,N_536);
nor U1047 (N_1047,N_109,N_859);
and U1048 (N_1048,In_2348,N_24);
and U1049 (N_1049,In_2339,N_174);
nand U1050 (N_1050,In_746,In_891);
and U1051 (N_1051,N_878,In_1082);
nand U1052 (N_1052,In_717,N_527);
nor U1053 (N_1053,N_148,N_343);
nor U1054 (N_1054,In_2503,N_140);
xnor U1055 (N_1055,In_2698,In_2890);
nor U1056 (N_1056,In_1595,In_2057);
nor U1057 (N_1057,N_302,In_733);
nor U1058 (N_1058,In_2321,N_324);
xnor U1059 (N_1059,In_2863,N_77);
nor U1060 (N_1060,In_2702,In_1034);
nand U1061 (N_1061,In_1954,N_10);
and U1062 (N_1062,N_873,In_937);
nor U1063 (N_1063,N_383,N_118);
and U1064 (N_1064,In_1455,In_1858);
xnor U1065 (N_1065,N_308,N_615);
xnor U1066 (N_1066,N_69,In_569);
or U1067 (N_1067,In_1812,N_0);
or U1068 (N_1068,In_1047,N_831);
nand U1069 (N_1069,In_1613,In_1152);
and U1070 (N_1070,N_713,In_2240);
xnor U1071 (N_1071,N_596,In_2460);
nor U1072 (N_1072,N_695,In_2474);
or U1073 (N_1073,In_2548,In_1671);
and U1074 (N_1074,N_740,N_821);
nand U1075 (N_1075,N_939,N_91);
and U1076 (N_1076,In_1685,N_188);
and U1077 (N_1077,N_620,In_203);
nand U1078 (N_1078,In_849,N_269);
nor U1079 (N_1079,N_67,N_292);
and U1080 (N_1080,N_424,N_51);
nor U1081 (N_1081,In_2006,N_818);
xnor U1082 (N_1082,In_1192,In_1458);
and U1083 (N_1083,In_1323,N_531);
xor U1084 (N_1084,N_975,In_1221);
nor U1085 (N_1085,N_433,In_1914);
or U1086 (N_1086,In_1908,In_1556);
nor U1087 (N_1087,In_2565,In_26);
nand U1088 (N_1088,N_346,In_1667);
nor U1089 (N_1089,N_307,In_128);
nand U1090 (N_1090,In_2353,In_2334);
and U1091 (N_1091,N_14,In_1807);
nor U1092 (N_1092,N_960,N_539);
nor U1093 (N_1093,N_764,In_2478);
and U1094 (N_1094,N_26,N_309);
or U1095 (N_1095,N_599,In_859);
xor U1096 (N_1096,N_619,In_1202);
and U1097 (N_1097,N_355,In_637);
nand U1098 (N_1098,N_430,N_636);
and U1099 (N_1099,N_201,N_605);
nand U1100 (N_1100,In_1582,In_1062);
nor U1101 (N_1101,In_101,In_2126);
or U1102 (N_1102,In_1251,N_268);
nand U1103 (N_1103,N_247,N_488);
xor U1104 (N_1104,In_1256,In_1159);
nor U1105 (N_1105,N_915,In_371);
or U1106 (N_1106,In_1983,N_645);
nand U1107 (N_1107,N_769,N_37);
or U1108 (N_1108,In_1958,In_1515);
nor U1109 (N_1109,In_2989,N_951);
nand U1110 (N_1110,N_543,In_560);
or U1111 (N_1111,N_225,N_330);
and U1112 (N_1112,N_138,In_311);
and U1113 (N_1113,N_776,In_1653);
nor U1114 (N_1114,In_2661,N_729);
nor U1115 (N_1115,In_2906,N_87);
nand U1116 (N_1116,In_2157,In_346);
nor U1117 (N_1117,In_1694,N_444);
and U1118 (N_1118,N_783,In_439);
nor U1119 (N_1119,In_1816,In_1703);
and U1120 (N_1120,In_1147,N_390);
xor U1121 (N_1121,N_360,N_560);
nand U1122 (N_1122,In_684,In_40);
and U1123 (N_1123,N_805,In_155);
and U1124 (N_1124,In_1533,N_425);
or U1125 (N_1125,N_443,N_437);
nor U1126 (N_1126,In_1385,In_2241);
nor U1127 (N_1127,N_592,In_402);
or U1128 (N_1128,In_2759,N_706);
and U1129 (N_1129,N_46,N_455);
and U1130 (N_1130,In_32,N_665);
nand U1131 (N_1131,N_312,N_505);
nor U1132 (N_1132,In_31,N_254);
or U1133 (N_1133,In_1939,In_224);
nand U1134 (N_1134,In_889,N_185);
xnor U1135 (N_1135,In_927,In_1528);
nor U1136 (N_1136,In_1603,N_770);
nor U1137 (N_1137,N_139,In_728);
xnor U1138 (N_1138,In_2252,N_249);
xor U1139 (N_1139,In_2933,In_1374);
nand U1140 (N_1140,N_162,In_1253);
nor U1141 (N_1141,N_237,In_383);
xnor U1142 (N_1142,N_794,In_2069);
and U1143 (N_1143,In_2134,In_2186);
and U1144 (N_1144,N_719,In_1081);
or U1145 (N_1145,In_1243,In_2706);
and U1146 (N_1146,In_2502,N_844);
xnor U1147 (N_1147,In_1187,N_632);
and U1148 (N_1148,In_1514,N_876);
or U1149 (N_1149,In_397,In_1312);
and U1150 (N_1150,N_240,In_1168);
nand U1151 (N_1151,N_105,In_172);
nor U1152 (N_1152,N_699,N_896);
xnor U1153 (N_1153,In_1906,N_426);
xor U1154 (N_1154,In_489,N_953);
and U1155 (N_1155,N_751,N_371);
nand U1156 (N_1156,N_119,In_1568);
and U1157 (N_1157,N_374,In_2276);
and U1158 (N_1158,N_63,In_1020);
and U1159 (N_1159,N_838,In_1890);
and U1160 (N_1160,In_1799,In_360);
nand U1161 (N_1161,In_421,In_1399);
nand U1162 (N_1162,N_226,In_481);
and U1163 (N_1163,In_783,N_81);
nand U1164 (N_1164,N_871,In_1707);
and U1165 (N_1165,N_441,In_1945);
or U1166 (N_1166,N_750,In_710);
nor U1167 (N_1167,In_163,N_277);
nor U1168 (N_1168,In_604,N_700);
xor U1169 (N_1169,In_1607,N_31);
or U1170 (N_1170,In_996,N_964);
or U1171 (N_1171,In_2014,N_870);
and U1172 (N_1172,N_976,N_722);
nand U1173 (N_1173,N_354,In_1252);
xnor U1174 (N_1174,In_2932,N_403);
or U1175 (N_1175,In_238,N_743);
xnor U1176 (N_1176,In_1161,In_144);
xor U1177 (N_1177,N_239,N_25);
nor U1178 (N_1178,In_1742,In_130);
nand U1179 (N_1179,In_2580,In_2424);
nand U1180 (N_1180,N_708,N_411);
nand U1181 (N_1181,N_1,In_355);
nor U1182 (N_1182,In_1764,In_2892);
and U1183 (N_1183,N_333,N_581);
nor U1184 (N_1184,N_916,N_887);
and U1185 (N_1185,In_1384,In_579);
or U1186 (N_1186,N_165,N_402);
nor U1187 (N_1187,In_2002,N_550);
nor U1188 (N_1188,In_2540,N_238);
and U1189 (N_1189,N_501,N_855);
and U1190 (N_1190,In_2803,In_2635);
nor U1191 (N_1191,N_52,N_481);
nand U1192 (N_1192,In_1318,N_294);
or U1193 (N_1193,N_670,In_1753);
xnor U1194 (N_1194,N_222,In_1074);
or U1195 (N_1195,In_863,In_2435);
and U1196 (N_1196,N_376,In_1524);
and U1197 (N_1197,N_717,In_372);
xor U1198 (N_1198,N_822,N_339);
or U1199 (N_1199,In_2273,N_946);
or U1200 (N_1200,In_2862,N_515);
nor U1201 (N_1201,In_1792,N_489);
and U1202 (N_1202,In_540,In_241);
or U1203 (N_1203,In_1701,N_907);
nand U1204 (N_1204,N_843,N_208);
or U1205 (N_1205,In_33,N_404);
nor U1206 (N_1206,In_2860,In_1234);
nor U1207 (N_1207,N_845,N_972);
xnor U1208 (N_1208,N_931,In_1349);
nand U1209 (N_1209,In_1702,N_236);
nand U1210 (N_1210,N_204,N_198);
or U1211 (N_1211,N_956,N_624);
xor U1212 (N_1212,N_190,N_123);
nor U1213 (N_1213,In_763,N_246);
xnor U1214 (N_1214,In_209,In_2297);
nand U1215 (N_1215,N_507,In_2127);
xnor U1216 (N_1216,In_1625,In_220);
xor U1217 (N_1217,N_952,N_984);
nand U1218 (N_1218,N_210,N_157);
or U1219 (N_1219,N_469,N_306);
and U1220 (N_1220,In_213,In_1881);
and U1221 (N_1221,N_72,In_2858);
nor U1222 (N_1222,N_38,N_196);
and U1223 (N_1223,In_2048,N_905);
and U1224 (N_1224,In_2485,In_2535);
nand U1225 (N_1225,In_2971,In_457);
or U1226 (N_1226,In_2924,In_1937);
xnor U1227 (N_1227,N_378,In_1602);
xor U1228 (N_1228,In_2215,In_2022);
or U1229 (N_1229,In_2814,In_115);
or U1230 (N_1230,N_385,In_1681);
xnor U1231 (N_1231,In_2684,In_1096);
nor U1232 (N_1232,N_275,In_1700);
xor U1233 (N_1233,In_2061,N_921);
nand U1234 (N_1234,In_1729,N_224);
nand U1235 (N_1235,N_797,In_1468);
xor U1236 (N_1236,N_900,In_1045);
and U1237 (N_1237,N_173,N_804);
or U1238 (N_1238,N_914,N_183);
or U1239 (N_1239,In_2398,N_78);
nand U1240 (N_1240,In_2651,In_1342);
and U1241 (N_1241,In_894,In_2305);
nor U1242 (N_1242,In_679,N_11);
nand U1243 (N_1243,In_1487,N_572);
nand U1244 (N_1244,N_839,N_350);
and U1245 (N_1245,In_1825,In_2477);
or U1246 (N_1246,In_584,In_2490);
nand U1247 (N_1247,In_2151,N_432);
xor U1248 (N_1248,In_2626,N_137);
and U1249 (N_1249,N_212,N_648);
or U1250 (N_1250,N_857,N_809);
nand U1251 (N_1251,N_27,N_777);
nor U1252 (N_1252,N_449,N_672);
nand U1253 (N_1253,In_2143,N_658);
or U1254 (N_1254,N_321,N_60);
nand U1255 (N_1255,N_549,N_879);
and U1256 (N_1256,In_1566,In_965);
nor U1257 (N_1257,N_568,In_1950);
and U1258 (N_1258,In_1271,N_147);
nor U1259 (N_1259,N_142,In_2695);
and U1260 (N_1260,N_647,In_969);
nand U1261 (N_1261,N_755,N_409);
and U1262 (N_1262,N_927,N_435);
and U1263 (N_1263,In_332,N_642);
nor U1264 (N_1264,N_718,N_889);
or U1265 (N_1265,In_2483,N_150);
nor U1266 (N_1266,In_1470,In_843);
nand U1267 (N_1267,In_1284,In_2214);
or U1268 (N_1268,N_396,In_1872);
and U1269 (N_1269,In_380,N_786);
and U1270 (N_1270,In_1041,N_891);
or U1271 (N_1271,In_2177,N_503);
nand U1272 (N_1272,In_1800,N_748);
nor U1273 (N_1273,N_16,In_2113);
nor U1274 (N_1274,In_2957,In_2923);
xnor U1275 (N_1275,In_2135,N_68);
or U1276 (N_1276,In_1779,N_117);
and U1277 (N_1277,N_932,N_657);
xor U1278 (N_1278,In_1088,N_417);
nor U1279 (N_1279,In_2148,In_1946);
nand U1280 (N_1280,N_785,N_169);
xnor U1281 (N_1281,In_1341,N_545);
xnor U1282 (N_1282,In_2796,N_528);
or U1283 (N_1283,N_84,N_479);
nand U1284 (N_1284,N_291,N_577);
xor U1285 (N_1285,N_690,N_135);
nor U1286 (N_1286,In_1461,In_931);
nand U1287 (N_1287,In_1931,N_412);
nand U1288 (N_1288,In_991,N_334);
and U1289 (N_1289,In_1173,In_473);
or U1290 (N_1290,In_2456,In_1331);
or U1291 (N_1291,N_182,N_781);
and U1292 (N_1292,In_1158,In_2538);
and U1293 (N_1293,N_184,In_1296);
or U1294 (N_1294,N_428,N_146);
or U1295 (N_1295,N_293,In_2258);
nor U1296 (N_1296,In_2947,N_968);
nor U1297 (N_1297,N_685,In_2964);
nand U1298 (N_1298,N_365,N_359);
and U1299 (N_1299,In_1913,N_652);
and U1300 (N_1300,N_586,In_1268);
xnor U1301 (N_1301,In_830,In_961);
xnor U1302 (N_1302,In_1810,In_453);
and U1303 (N_1303,N_710,In_2800);
xnor U1304 (N_1304,N_89,N_912);
and U1305 (N_1305,In_935,N_661);
or U1306 (N_1306,N_436,In_2758);
nor U1307 (N_1307,N_116,N_806);
and U1308 (N_1308,In_1117,In_1550);
nand U1309 (N_1309,In_627,In_1208);
and U1310 (N_1310,In_1024,N_943);
xor U1311 (N_1311,In_2983,In_1002);
xor U1312 (N_1312,In_2984,N_676);
nand U1313 (N_1313,N_234,N_908);
nor U1314 (N_1314,N_944,In_2836);
nor U1315 (N_1315,In_1309,N_28);
nor U1316 (N_1316,In_1408,In_860);
nand U1317 (N_1317,N_389,In_634);
nor U1318 (N_1318,In_293,In_2271);
xnor U1319 (N_1319,N_59,In_811);
or U1320 (N_1320,N_74,N_851);
nor U1321 (N_1321,N_570,In_1952);
or U1322 (N_1322,N_7,In_2256);
or U1323 (N_1323,N_442,In_647);
and U1324 (N_1324,N_384,N_653);
nor U1325 (N_1325,In_1003,N_8);
and U1326 (N_1326,N_332,In_141);
nor U1327 (N_1327,N_58,N_850);
and U1328 (N_1328,In_2512,N_500);
or U1329 (N_1329,N_241,In_1395);
xnor U1330 (N_1330,In_1283,In_308);
xnor U1331 (N_1331,In_488,In_2692);
nor U1332 (N_1332,N_714,N_664);
or U1333 (N_1333,N_213,In_1721);
nor U1334 (N_1334,N_22,N_790);
and U1335 (N_1335,In_2645,In_1052);
and U1336 (N_1336,N_361,In_787);
xor U1337 (N_1337,N_858,In_506);
xnor U1338 (N_1338,N_416,In_2042);
xnor U1339 (N_1339,In_2513,N_480);
or U1340 (N_1340,N_50,N_71);
nand U1341 (N_1341,N_98,N_773);
or U1342 (N_1342,N_471,In_2741);
nand U1343 (N_1343,In_700,N_848);
or U1344 (N_1344,N_215,In_1808);
or U1345 (N_1345,N_812,In_1471);
nand U1346 (N_1346,N_363,In_1852);
and U1347 (N_1347,N_338,In_1135);
and U1348 (N_1348,In_1375,In_407);
xor U1349 (N_1349,In_1619,N_440);
nor U1350 (N_1350,In_589,N_659);
nand U1351 (N_1351,In_921,N_235);
or U1352 (N_1352,N_382,N_633);
nand U1353 (N_1353,N_534,N_464);
nor U1354 (N_1354,In_89,N_348);
and U1355 (N_1355,N_888,N_872);
or U1356 (N_1356,In_764,In_2336);
nor U1357 (N_1357,N_410,N_513);
or U1358 (N_1358,In_2103,In_1886);
xnor U1359 (N_1359,In_2820,N_472);
xor U1360 (N_1360,N_506,N_836);
nand U1361 (N_1361,N_780,In_1435);
xnor U1362 (N_1362,In_1709,N_698);
nor U1363 (N_1363,In_1377,In_2908);
nand U1364 (N_1364,In_2575,In_2287);
nor U1365 (N_1365,In_1775,In_2248);
xnor U1366 (N_1366,N_727,N_792);
or U1367 (N_1367,N_823,N_928);
nand U1368 (N_1368,N_454,In_231);
nor U1369 (N_1369,In_1909,In_955);
or U1370 (N_1370,In_2696,N_622);
xnor U1371 (N_1371,In_2959,In_909);
xor U1372 (N_1372,In_454,N_999);
nand U1373 (N_1373,In_2598,N_662);
or U1374 (N_1374,N_761,In_1416);
nand U1375 (N_1375,In_2030,In_2155);
or U1376 (N_1376,In_2519,N_336);
nand U1377 (N_1377,N_232,In_419);
or U1378 (N_1378,N_75,N_612);
or U1379 (N_1379,N_917,N_41);
and U1380 (N_1380,N_906,N_186);
or U1381 (N_1381,In_2631,N_774);
and U1382 (N_1382,N_995,In_2255);
nor U1383 (N_1383,N_650,In_2449);
and U1384 (N_1384,In_1388,In_2005);
nor U1385 (N_1385,N_55,In_470);
nand U1386 (N_1386,N_969,In_229);
and U1387 (N_1387,In_176,In_145);
xor U1388 (N_1388,N_694,In_2123);
nand U1389 (N_1389,In_222,N_919);
nor U1390 (N_1390,In_2745,N_556);
and U1391 (N_1391,In_623,N_646);
and U1392 (N_1392,In_977,In_933);
nor U1393 (N_1393,N_853,N_591);
xnor U1394 (N_1394,N_816,N_967);
or U1395 (N_1395,In_1242,In_36);
xor U1396 (N_1396,N_959,In_1732);
nor U1397 (N_1397,N_97,In_187);
nor U1398 (N_1398,In_363,In_1181);
and U1399 (N_1399,N_893,In_1597);
and U1400 (N_1400,In_1994,In_1266);
nor U1401 (N_1401,N_104,N_211);
or U1402 (N_1402,In_1728,In_2080);
nor U1403 (N_1403,In_2359,In_865);
nand U1404 (N_1404,In_2401,N_911);
or U1405 (N_1405,In_268,N_289);
nor U1406 (N_1406,N_133,In_1684);
nor U1407 (N_1407,N_301,In_1425);
nand U1408 (N_1408,In_1365,N_863);
nand U1409 (N_1409,N_30,In_62);
xnor U1410 (N_1410,N_546,In_1348);
and U1411 (N_1411,N_526,In_2856);
nor U1412 (N_1412,In_1669,N_295);
nor U1413 (N_1413,N_778,N_731);
nand U1414 (N_1414,N_191,In_1481);
nand U1415 (N_1415,N_692,In_347);
and U1416 (N_1416,N_126,N_187);
nor U1417 (N_1417,In_2050,N_90);
or U1418 (N_1418,In_1499,In_2016);
xnor U1419 (N_1419,In_1224,N_265);
xor U1420 (N_1420,N_209,N_895);
xnor U1421 (N_1421,In_430,N_230);
nand U1422 (N_1422,In_1588,In_2919);
xnor U1423 (N_1423,In_22,N_54);
xor U1424 (N_1424,N_419,N_445);
xnor U1425 (N_1425,N_795,N_547);
xnor U1426 (N_1426,In_2497,N_897);
or U1427 (N_1427,N_977,In_1664);
or U1428 (N_1428,In_2584,N_96);
or U1429 (N_1429,N_113,N_758);
nor U1430 (N_1430,N_314,N_493);
nand U1431 (N_1431,N_965,In_2411);
nor U1432 (N_1432,In_434,N_909);
xor U1433 (N_1433,In_643,In_2249);
nor U1434 (N_1434,N_451,N_391);
xnor U1435 (N_1435,N_53,In_2229);
xnor U1436 (N_1436,In_2358,In_2226);
xor U1437 (N_1437,In_2228,In_1429);
nand U1438 (N_1438,In_1736,In_2623);
and U1439 (N_1439,In_600,In_2280);
or U1440 (N_1440,In_954,In_2913);
or U1441 (N_1441,N_723,In_1522);
and U1442 (N_1442,In_2639,N_971);
and U1443 (N_1443,In_1196,In_504);
nand U1444 (N_1444,In_2013,N_651);
nand U1445 (N_1445,In_1997,In_2531);
xor U1446 (N_1446,In_1865,N_108);
nor U1447 (N_1447,In_759,N_910);
nand U1448 (N_1448,In_129,N_167);
nand U1449 (N_1449,In_2952,In_1691);
or U1450 (N_1450,In_243,N_478);
and U1451 (N_1451,N_149,In_2884);
xnor U1452 (N_1452,In_2705,In_2149);
xnor U1453 (N_1453,N_203,N_950);
nor U1454 (N_1454,In_695,N_207);
xnor U1455 (N_1455,N_228,In_210);
and U1456 (N_1456,N_934,N_107);
nand U1457 (N_1457,N_551,In_888);
or U1458 (N_1458,N_45,In_2031);
and U1459 (N_1459,N_144,N_715);
xor U1460 (N_1460,In_99,N_578);
nor U1461 (N_1461,In_2788,N_305);
nor U1462 (N_1462,N_732,In_2236);
and U1463 (N_1463,N_400,N_94);
xnor U1464 (N_1464,N_847,In_118);
xor U1465 (N_1465,In_2087,N_200);
nand U1466 (N_1466,In_1693,In_1100);
and U1467 (N_1467,N_357,N_869);
nand U1468 (N_1468,In_547,In_1747);
nor U1469 (N_1469,In_2160,N_626);
nand U1470 (N_1470,N_678,In_2889);
or U1471 (N_1471,N_625,In_1599);
and U1472 (N_1472,In_1780,In_1346);
xor U1473 (N_1473,In_818,N_533);
xor U1474 (N_1474,In_331,In_75);
xnor U1475 (N_1475,N_571,In_1970);
and U1476 (N_1476,N_554,N_784);
and U1477 (N_1477,N_686,N_155);
xor U1478 (N_1478,N_176,In_2501);
and U1479 (N_1479,In_1324,N_593);
and U1480 (N_1480,N_482,In_2557);
nand U1481 (N_1481,N_904,N_233);
xor U1482 (N_1482,N_553,N_29);
nor U1483 (N_1483,N_803,N_460);
or U1484 (N_1484,N_711,In_343);
xnor U1485 (N_1485,N_492,N_342);
nor U1486 (N_1486,N_925,N_76);
nand U1487 (N_1487,N_635,N_757);
or U1488 (N_1488,N_504,N_453);
xor U1489 (N_1489,In_2986,In_676);
xnor U1490 (N_1490,In_873,N_154);
nand U1491 (N_1491,In_1526,In_48);
xor U1492 (N_1492,N_962,In_1609);
or U1493 (N_1493,N_452,In_2763);
and U1494 (N_1494,In_2998,N_988);
nand U1495 (N_1495,In_1489,In_1038);
and U1496 (N_1496,N_260,N_584);
nand U1497 (N_1497,In_611,In_887);
nor U1498 (N_1498,In_1895,N_600);
nand U1499 (N_1499,N_356,In_2681);
xor U1500 (N_1500,N_106,N_899);
and U1501 (N_1501,N_279,N_555);
xnor U1502 (N_1502,In_786,In_1608);
or U1503 (N_1503,N_978,In_2619);
nor U1504 (N_1504,N_594,In_1642);
and U1505 (N_1505,N_558,In_929);
nor U1506 (N_1506,N_490,In_892);
and U1507 (N_1507,In_2282,In_406);
nand U1508 (N_1508,In_1317,N_216);
and U1509 (N_1509,In_433,In_2179);
xor U1510 (N_1510,N_703,N_865);
or U1511 (N_1511,In_2677,In_190);
nor U1512 (N_1512,N_303,In_1031);
nor U1513 (N_1513,N_512,N_986);
and U1514 (N_1514,N_284,N_407);
and U1515 (N_1515,N_881,In_2833);
xor U1516 (N_1516,In_649,In_8);
and U1517 (N_1517,N_745,N_219);
and U1518 (N_1518,In_2717,In_1013);
nand U1519 (N_1519,N_56,N_47);
and U1520 (N_1520,In_425,N_272);
and U1521 (N_1521,In_1389,In_225);
xor U1522 (N_1522,In_240,N_347);
or U1523 (N_1523,N_151,N_958);
nor U1524 (N_1524,In_139,In_188);
or U1525 (N_1525,N_609,In_2898);
and U1526 (N_1526,In_1708,N_364);
or U1527 (N_1527,In_1340,In_1043);
nand U1528 (N_1528,In_502,In_2838);
and U1529 (N_1529,In_2916,In_2154);
xnor U1530 (N_1530,N_837,N_993);
nor U1531 (N_1531,N_66,N_62);
or U1532 (N_1532,N_875,N_287);
or U1533 (N_1533,N_992,N_521);
and U1534 (N_1534,N_687,N_832);
and U1535 (N_1535,In_1902,N_102);
or U1536 (N_1536,N_476,N_152);
nand U1537 (N_1537,In_292,In_995);
nand U1538 (N_1538,In_2672,N_574);
nand U1539 (N_1539,N_358,In_562);
nor U1540 (N_1540,N_48,In_1093);
and U1541 (N_1541,N_17,In_18);
xnor U1542 (N_1542,N_707,In_1722);
xnor U1543 (N_1543,In_639,In_394);
nor U1544 (N_1544,N_810,In_551);
and U1545 (N_1545,In_375,N_643);
nor U1546 (N_1546,In_587,N_884);
nand U1547 (N_1547,N_381,In_2268);
or U1548 (N_1548,N_573,In_2778);
nand U1549 (N_1549,In_2612,N_112);
nor U1550 (N_1550,N_981,In_2455);
xnor U1551 (N_1551,N_765,N_523);
nor U1552 (N_1552,N_178,In_1177);
nand U1553 (N_1553,N_898,In_2831);
nand U1554 (N_1554,N_752,In_1637);
or U1555 (N_1555,N_569,In_570);
or U1556 (N_1556,N_994,N_989);
and U1557 (N_1557,N_608,N_789);
or U1558 (N_1558,N_736,N_826);
or U1559 (N_1559,N_319,N_901);
or U1560 (N_1560,N_772,In_2289);
nor U1561 (N_1561,In_348,N_206);
nand U1562 (N_1562,N_819,In_452);
nand U1563 (N_1563,N_629,In_729);
xnor U1564 (N_1564,N_70,N_579);
nand U1565 (N_1565,In_494,N_775);
or U1566 (N_1566,N_771,N_175);
or U1567 (N_1567,In_79,N_520);
or U1568 (N_1568,In_201,In_333);
nand U1569 (N_1569,In_511,N_405);
xnor U1570 (N_1570,In_1420,In_120);
nand U1571 (N_1571,In_1650,N_656);
or U1572 (N_1572,In_2915,N_532);
xor U1573 (N_1573,N_487,N_660);
nor U1574 (N_1574,In_2595,N_495);
or U1575 (N_1575,In_557,In_1804);
and U1576 (N_1576,N_386,In_1393);
or U1577 (N_1577,In_2907,In_1379);
or U1578 (N_1578,In_2599,In_561);
nand U1579 (N_1579,In_2369,In_2616);
or U1580 (N_1580,N_65,N_926);
or U1581 (N_1581,In_1589,N_666);
xnor U1582 (N_1582,In_1964,N_296);
and U1583 (N_1583,N_49,In_2296);
nor U1584 (N_1584,N_702,N_483);
or U1585 (N_1585,N_918,N_399);
xor U1586 (N_1586,In_2894,N_408);
and U1587 (N_1587,N_935,In_1835);
xor U1588 (N_1588,In_2442,N_195);
or U1589 (N_1589,In_2454,N_726);
xor U1590 (N_1590,N_885,In_325);
nand U1591 (N_1591,In_1948,In_853);
and U1592 (N_1592,N_575,N_961);
and U1593 (N_1593,N_595,In_1050);
xnor U1594 (N_1594,N_160,In_296);
nor U1595 (N_1595,N_948,In_198);
and U1596 (N_1596,In_1071,In_1905);
xor U1597 (N_1597,N_217,N_580);
xor U1598 (N_1598,In_855,In_2326);
xnor U1599 (N_1599,In_416,N_323);
or U1600 (N_1600,N_617,In_310);
nand U1601 (N_1601,N_255,In_17);
and U1602 (N_1602,In_1960,In_1211);
and U1603 (N_1603,N_630,In_116);
and U1604 (N_1604,N_406,N_738);
nand U1605 (N_1605,N_370,In_444);
or U1606 (N_1606,N_990,In_1488);
xnor U1607 (N_1607,N_677,N_987);
nand U1608 (N_1608,In_1079,In_2266);
nor U1609 (N_1609,In_750,In_1853);
nor U1610 (N_1610,N_563,N_671);
xor U1611 (N_1611,In_608,In_1646);
nand U1612 (N_1612,N_276,N_164);
nor U1613 (N_1613,N_3,In_809);
nand U1614 (N_1614,In_719,N_730);
nand U1615 (N_1615,In_2189,In_1184);
and U1616 (N_1616,N_903,In_667);
or U1617 (N_1617,N_375,In_2338);
xnor U1618 (N_1618,In_207,In_244);
nor U1619 (N_1619,N_125,N_530);
or U1620 (N_1620,In_655,N_963);
or U1621 (N_1621,N_588,In_1449);
nand U1622 (N_1622,In_505,N_418);
nor U1623 (N_1623,N_628,In_1784);
xnor U1624 (N_1624,In_1103,In_1765);
nand U1625 (N_1625,In_2515,N_484);
nand U1626 (N_1626,N_180,In_519);
nand U1627 (N_1627,In_1513,N_674);
nand U1628 (N_1628,In_1141,N_242);
and U1629 (N_1629,In_1562,N_985);
and U1630 (N_1630,N_380,N_486);
and U1631 (N_1631,In_1836,In_2850);
xnor U1632 (N_1632,N_202,In_563);
xnor U1633 (N_1633,N_253,N_701);
xor U1634 (N_1634,In_1995,N_734);
and U1635 (N_1635,N_582,N_742);
or U1636 (N_1636,In_272,N_587);
nor U1637 (N_1637,N_421,In_1754);
and U1638 (N_1638,N_189,In_1919);
nor U1639 (N_1639,N_244,In_2365);
xor U1640 (N_1640,In_1643,In_1859);
nand U1641 (N_1641,In_1698,In_1215);
xnor U1642 (N_1642,In_147,N_79);
or U1643 (N_1643,N_100,In_698);
or U1644 (N_1644,In_2077,In_230);
and U1645 (N_1645,In_2854,In_1822);
xnor U1646 (N_1646,N_439,In_1979);
xnor U1647 (N_1647,N_73,N_327);
or U1648 (N_1648,N_145,N_705);
nand U1649 (N_1649,In_361,N_44);
or U1650 (N_1650,N_639,N_351);
nand U1651 (N_1651,In_178,N_475);
xnor U1652 (N_1652,In_2073,N_9);
xor U1653 (N_1653,In_1509,N_800);
or U1654 (N_1654,In_2806,In_2191);
xnor U1655 (N_1655,N_991,In_1975);
or U1656 (N_1656,In_1355,In_2521);
nor U1657 (N_1657,N_861,In_2303);
xnor U1658 (N_1658,N_20,N_548);
and U1659 (N_1659,N_388,N_457);
nor U1660 (N_1660,N_518,N_136);
nor U1661 (N_1661,In_2561,In_301);
xor U1662 (N_1662,N_627,In_2934);
xor U1663 (N_1663,N_802,N_111);
or U1664 (N_1664,N_741,In_2047);
and U1665 (N_1665,In_645,In_2298);
nand U1666 (N_1666,N_955,In_497);
xnor U1667 (N_1667,N_874,In_1291);
or U1668 (N_1668,In_1715,N_974);
and U1669 (N_1669,N_720,In_77);
xnor U1670 (N_1670,In_625,In_1000);
nor U1671 (N_1671,N_414,In_339);
nor U1672 (N_1672,In_567,In_38);
xnor U1673 (N_1673,N_2,N_936);
or U1674 (N_1674,N_220,N_945);
or U1675 (N_1675,In_635,In_2010);
and U1676 (N_1676,N_697,N_683);
and U1677 (N_1677,In_1347,N_603);
or U1678 (N_1678,N_263,In_674);
nor U1679 (N_1679,N_747,N_709);
nand U1680 (N_1680,N_544,In_2244);
and U1681 (N_1681,In_313,In_2067);
xor U1682 (N_1682,In_353,In_2721);
and U1683 (N_1683,In_1360,In_1674);
nand U1684 (N_1684,In_2379,N_693);
nand U1685 (N_1685,N_285,In_1259);
nor U1686 (N_1686,In_2930,N_82);
or U1687 (N_1687,In_2824,In_1731);
nand U1688 (N_1688,N_669,In_1409);
xor U1689 (N_1689,In_287,N_168);
nor U1690 (N_1690,N_923,N_824);
nand U1691 (N_1691,N_243,N_379);
and U1692 (N_1692,In_1127,N_640);
nand U1693 (N_1693,N_638,N_465);
and U1694 (N_1694,N_218,In_35);
nor U1695 (N_1695,In_542,In_1981);
nor U1696 (N_1696,N_815,In_1239);
and U1697 (N_1697,N_340,N_799);
and U1698 (N_1698,N_458,In_367);
nor U1699 (N_1699,N_733,In_1250);
nor U1700 (N_1700,In_173,N_868);
or U1701 (N_1701,In_513,In_1137);
and U1702 (N_1702,N_115,In_824);
xnor U1703 (N_1703,N_542,In_499);
and U1704 (N_1704,N_331,In_900);
nand U1705 (N_1705,N_231,N_341);
or U1706 (N_1706,In_2156,N_668);
or U1707 (N_1707,N_613,N_817);
or U1708 (N_1708,In_2421,In_1029);
xor U1709 (N_1709,N_368,In_2181);
xor U1710 (N_1710,In_1413,In_603);
and U1711 (N_1711,N_466,N_590);
xnor U1712 (N_1712,In_1149,In_2043);
xnor U1713 (N_1713,In_2168,In_298);
nor U1714 (N_1714,In_630,In_2654);
or U1715 (N_1715,In_2582,N_311);
nand U1716 (N_1716,N_264,In_43);
and U1717 (N_1717,In_2055,In_2213);
nand U1718 (N_1718,N_245,N_177);
nor U1719 (N_1719,In_2725,N_655);
nor U1720 (N_1720,In_2178,In_1163);
xor U1721 (N_1721,In_776,In_2370);
xor U1722 (N_1722,In_69,N_852);
or U1723 (N_1723,In_1278,N_760);
or U1724 (N_1724,In_487,N_663);
or U1725 (N_1725,N_199,N_514);
nor U1726 (N_1726,N_192,N_601);
xnor U1727 (N_1727,N_256,In_256);
nor U1728 (N_1728,N_141,In_248);
nor U1729 (N_1729,N_811,N_798);
xnor U1730 (N_1730,In_2480,In_2219);
or U1731 (N_1731,N_767,In_80);
and U1732 (N_1732,N_924,N_746);
nand U1733 (N_1733,In_2443,In_1947);
and U1734 (N_1734,In_760,N_194);
nand U1735 (N_1735,In_1629,In_2766);
or U1736 (N_1736,N_682,N_675);
nor U1737 (N_1737,N_57,In_1932);
xor U1738 (N_1738,N_882,N_833);
or U1739 (N_1739,In_1160,In_1546);
xnor U1740 (N_1740,N_310,In_2738);
nor U1741 (N_1741,In_1714,N_39);
nand U1742 (N_1742,N_947,N_866);
or U1743 (N_1743,N_814,In_152);
or U1744 (N_1744,N_5,N_813);
and U1745 (N_1745,In_2059,In_1433);
and U1746 (N_1746,In_2724,In_2597);
nand U1747 (N_1747,N_470,N_401);
or U1748 (N_1748,N_721,N_288);
nand U1749 (N_1749,N_938,N_712);
nand U1750 (N_1750,In_1717,In_712);
xor U1751 (N_1751,N_258,N_966);
nor U1752 (N_1752,In_1319,In_2235);
and U1753 (N_1753,N_749,N_725);
and U1754 (N_1754,In_2781,In_507);
or U1755 (N_1755,N_886,In_2410);
nand U1756 (N_1756,In_2813,In_766);
nand U1757 (N_1757,In_1537,In_27);
xnor U1758 (N_1758,N_522,N_362);
and U1759 (N_1759,N_637,N_130);
xor U1760 (N_1760,N_250,In_435);
xnor U1761 (N_1761,In_2121,In_869);
nor U1762 (N_1762,In_81,N_623);
xor U1763 (N_1763,In_132,N_737);
xnor U1764 (N_1764,N_485,N_88);
and U1765 (N_1765,In_1307,In_2253);
and U1766 (N_1766,N_158,N_524);
nand U1767 (N_1767,In_2591,N_286);
or U1768 (N_1768,N_413,N_688);
and U1769 (N_1769,In_306,In_686);
and U1770 (N_1770,In_2170,N_862);
nand U1771 (N_1771,In_544,N_649);
and U1772 (N_1772,In_1462,In_1194);
nand U1773 (N_1773,N_373,In_2190);
and U1774 (N_1774,N_423,In_522);
and U1775 (N_1775,In_1726,N_85);
and U1776 (N_1776,In_1985,N_159);
and U1777 (N_1777,N_259,In_2636);
and U1778 (N_1778,In_581,In_2301);
xor U1779 (N_1779,In_2982,In_964);
or U1780 (N_1780,N_849,In_1791);
nand U1781 (N_1781,N_23,N_13);
or U1782 (N_1782,In_831,N_463);
nand U1783 (N_1783,N_667,N_352);
and U1784 (N_1784,In_1354,N_120);
nor U1785 (N_1785,N_980,In_2017);
nor U1786 (N_1786,N_929,N_537);
or U1787 (N_1787,N_101,N_467);
and U1788 (N_1788,N_86,In_2393);
xor U1789 (N_1789,In_752,N_299);
xor U1790 (N_1790,In_154,N_33);
xnor U1791 (N_1791,In_2564,In_1322);
nand U1792 (N_1792,In_1553,In_1579);
nand U1793 (N_1793,N_438,In_356);
nand U1794 (N_1794,In_1212,N_835);
xor U1795 (N_1795,N_398,In_1289);
nand U1796 (N_1796,In_2037,In_800);
nand U1797 (N_1797,N_267,N_248);
and U1798 (N_1798,In_875,N_892);
and U1799 (N_1799,N_61,N_283);
or U1800 (N_1800,In_539,N_282);
xnor U1801 (N_1801,N_634,In_113);
nand U1802 (N_1802,N_606,N_519);
nand U1803 (N_1803,In_1362,N_320);
nor U1804 (N_1804,In_142,In_2569);
nor U1805 (N_1805,N_477,In_1205);
and U1806 (N_1806,In_2400,N_830);
or U1807 (N_1807,In_2027,N_372);
nand U1808 (N_1808,In_13,N_345);
and U1809 (N_1809,In_2966,In_1143);
and U1810 (N_1810,In_819,In_1665);
nor U1811 (N_1811,In_1612,In_2965);
and U1812 (N_1812,In_2576,N_313);
or U1813 (N_1813,N_942,N_166);
and U1814 (N_1814,In_1893,N_681);
nand U1815 (N_1815,In_757,N_562);
or U1816 (N_1816,In_2524,In_582);
or U1817 (N_1817,In_2648,In_123);
and U1818 (N_1818,N_607,N_12);
nor U1819 (N_1819,N_205,In_1883);
xor U1820 (N_1820,In_171,N_337);
xor U1821 (N_1821,N_883,In_351);
nand U1822 (N_1822,In_2125,N_561);
and U1823 (N_1823,N_462,N_387);
or U1824 (N_1824,In_2586,In_2054);
or U1825 (N_1825,In_2292,N_583);
or U1826 (N_1826,In_44,N_920);
or U1827 (N_1827,N_161,N_124);
xnor U1828 (N_1828,In_680,In_2627);
nor U1829 (N_1829,N_325,In_1740);
nor U1830 (N_1830,N_214,In_401);
nand U1831 (N_1831,In_2857,In_694);
and U1832 (N_1832,In_618,N_179);
or U1833 (N_1833,N_841,N_597);
and U1834 (N_1834,In_2904,N_509);
or U1835 (N_1835,In_1380,N_644);
xnor U1836 (N_1836,N_318,N_827);
nand U1837 (N_1837,In_1472,In_2949);
and U1838 (N_1838,N_274,In_1119);
and U1839 (N_1839,In_2839,N_856);
nand U1840 (N_1840,N_890,In_1830);
nand U1841 (N_1841,In_55,N_497);
nor U1842 (N_1842,In_2769,In_1235);
xnor U1843 (N_1843,In_2737,N_834);
nand U1844 (N_1844,In_556,N_251);
nor U1845 (N_1845,N_604,N_618);
and U1846 (N_1846,N_498,N_680);
nand U1847 (N_1847,In_2382,In_2362);
or U1848 (N_1848,N_468,In_1398);
or U1849 (N_1849,In_861,In_2532);
and U1850 (N_1850,In_1146,N_278);
and U1851 (N_1851,In_2790,N_297);
xnor U1852 (N_1852,N_394,In_1969);
or U1853 (N_1853,N_132,In_2223);
nand U1854 (N_1854,N_735,In_465);
xnor U1855 (N_1855,In_829,N_134);
nor U1856 (N_1856,In_687,In_1343);
nor U1857 (N_1857,N_744,In_1310);
or U1858 (N_1858,In_1752,In_1910);
nor U1859 (N_1859,N_92,N_270);
and U1860 (N_1860,N_114,In_2944);
xnor U1861 (N_1861,In_683,N_877);
xnor U1862 (N_1862,N_456,In_621);
nor U1863 (N_1863,N_353,N_788);
nand U1864 (N_1864,N_80,N_691);
or U1865 (N_1865,In_1505,N_502);
nand U1866 (N_1866,N_724,N_820);
nor U1867 (N_1867,In_2550,N_163);
xor U1868 (N_1868,In_2458,In_922);
nor U1869 (N_1869,In_2212,In_896);
or U1870 (N_1870,In_1813,N_448);
or U1871 (N_1871,N_266,N_415);
nor U1872 (N_1872,N_95,N_842);
xnor U1873 (N_1873,N_508,In_1335);
xor U1874 (N_1874,N_538,In_2247);
and U1875 (N_1875,In_2507,N_728);
nor U1876 (N_1876,In_326,In_1575);
nand U1877 (N_1877,In_1460,N_759);
nor U1878 (N_1878,In_2782,In_2791);
xnor U1879 (N_1879,N_143,N_6);
nand U1880 (N_1880,In_2332,N_611);
nor U1881 (N_1881,N_496,In_2414);
nand U1882 (N_1882,In_2230,In_2496);
and U1883 (N_1883,N_997,N_673);
nor U1884 (N_1884,In_2314,In_1055);
or U1885 (N_1885,N_840,In_1739);
nor U1886 (N_1886,N_631,N_326);
nand U1887 (N_1887,N_979,N_290);
xnor U1888 (N_1888,N_221,In_2052);
nand U1889 (N_1889,In_1877,In_2234);
or U1890 (N_1890,N_377,N_131);
nor U1891 (N_1891,In_2729,In_1263);
xor U1892 (N_1892,In_2128,N_83);
nand U1893 (N_1893,In_37,In_997);
xnor U1894 (N_1894,N_40,N_602);
nand U1895 (N_1895,N_954,N_768);
and U1896 (N_1896,N_229,N_529);
nor U1897 (N_1897,In_1577,N_434);
or U1898 (N_1898,N_557,In_2015);
xnor U1899 (N_1899,In_2427,In_662);
or U1900 (N_1900,N_429,In_2972);
or U1901 (N_1901,N_763,N_252);
or U1902 (N_1902,N_621,N_704);
xor U1903 (N_1903,N_894,In_2553);
nor U1904 (N_1904,N_461,N_397);
and U1905 (N_1905,In_2837,In_893);
nor U1906 (N_1906,In_2445,N_933);
and U1907 (N_1907,N_779,N_34);
and U1908 (N_1908,N_171,N_585);
nand U1909 (N_1909,In_2859,In_2074);
xnor U1910 (N_1910,N_941,In_59);
and U1911 (N_1911,In_2981,N_564);
nor U1912 (N_1912,In_2320,N_782);
nand U1913 (N_1913,N_93,In_1907);
xor U1914 (N_1914,In_1523,N_854);
nand U1915 (N_1915,N_982,N_949);
and U1916 (N_1916,N_420,N_42);
xor U1917 (N_1917,N_793,In_484);
or U1918 (N_1918,In_341,In_1153);
nor U1919 (N_1919,N_996,In_2076);
xnor U1920 (N_1920,N_610,In_258);
xor U1921 (N_1921,N_262,In_1423);
nand U1922 (N_1922,In_1917,In_1121);
nand U1923 (N_1923,N_808,In_2462);
and U1924 (N_1924,N_716,N_739);
or U1925 (N_1925,N_64,In_919);
xor U1926 (N_1926,In_2274,In_2558);
nand U1927 (N_1927,In_1569,In_1397);
or U1928 (N_1928,N_273,N_754);
nand U1929 (N_1929,In_804,N_422);
and U1930 (N_1930,In_1070,N_99);
and U1931 (N_1931,N_525,N_829);
nand U1932 (N_1932,N_684,In_1957);
nor U1933 (N_1933,In_777,In_2021);
or U1934 (N_1934,N_937,N_499);
or U1935 (N_1935,In_1867,In_317);
xnor U1936 (N_1936,N_172,In_2807);
or U1937 (N_1937,In_2354,N_322);
nor U1938 (N_1938,N_517,In_1592);
nor U1939 (N_1939,In_2420,N_957);
nand U1940 (N_1940,In_192,In_232);
and U1941 (N_1941,In_1641,In_2735);
nor U1942 (N_1942,N_181,N_35);
nor U1943 (N_1943,In_795,N_4);
xnor U1944 (N_1944,In_1648,In_223);
and U1945 (N_1945,N_395,N_227);
or U1946 (N_1946,N_170,N_689);
or U1947 (N_1947,N_791,In_2583);
xor U1948 (N_1948,In_1787,N_552);
xnor U1949 (N_1949,N_298,In_1670);
and U1950 (N_1950,In_2093,N_393);
nand U1951 (N_1951,In_71,N_110);
xor U1952 (N_1952,N_223,In_1918);
xor U1953 (N_1953,In_295,In_1936);
nor U1954 (N_1954,N_796,N_540);
nand U1955 (N_1955,In_2697,In_1770);
and U1956 (N_1956,In_2433,In_1313);
or U1957 (N_1957,In_2114,N_535);
and U1958 (N_1958,In_1363,In_1605);
xor U1959 (N_1959,N_344,N_459);
nand U1960 (N_1960,In_2130,N_679);
nor U1961 (N_1961,N_801,N_32);
or U1962 (N_1962,N_970,N_541);
and U1963 (N_1963,N_828,In_428);
nand U1964 (N_1964,In_1101,N_129);
xor U1965 (N_1965,N_565,N_446);
xor U1966 (N_1966,N_193,In_1482);
and U1967 (N_1967,N_867,N_315);
nor U1968 (N_1968,In_1303,In_1547);
nand U1969 (N_1969,N_973,N_696);
xor U1970 (N_1970,In_2808,In_2752);
nor U1971 (N_1971,N_559,In_2425);
and U1972 (N_1972,In_1448,N_567);
or U1973 (N_1973,In_1730,In_41);
and U1974 (N_1974,N_366,In_1535);
xnor U1975 (N_1975,N_616,N_473);
nand U1976 (N_1976,In_2142,N_576);
xor U1977 (N_1977,In_663,In_314);
nor U1978 (N_1978,In_2152,In_25);
xor U1979 (N_1979,In_485,N_317);
and U1980 (N_1980,N_392,N_614);
or U1981 (N_1981,In_956,In_590);
nor U1982 (N_1982,N_328,In_735);
nor U1983 (N_1983,N_598,N_36);
and U1984 (N_1984,N_860,In_159);
nand U1985 (N_1985,In_2012,In_1875);
or U1986 (N_1986,In_1827,N_18);
and U1987 (N_1987,N_787,N_846);
xor U1988 (N_1988,N_566,In_1856);
nor U1989 (N_1989,In_307,In_2853);
and U1990 (N_1990,In_67,In_664);
or U1991 (N_1991,In_2035,N_127);
xor U1992 (N_1992,In_514,N_257);
nand U1993 (N_1993,N_281,N_753);
nand U1994 (N_1994,N_491,In_2749);
and U1995 (N_1995,In_2242,N_103);
nor U1996 (N_1996,In_1032,N_998);
nor U1997 (N_1997,N_510,N_922);
and U1998 (N_1998,In_2657,N_983);
xnor U1999 (N_1999,In_1396,In_2317);
nand U2000 (N_2000,N_1024,N_1184);
nand U2001 (N_2001,N_1565,N_1655);
and U2002 (N_2002,N_1992,N_1075);
xnor U2003 (N_2003,N_1066,N_1708);
and U2004 (N_2004,N_1784,N_1892);
xnor U2005 (N_2005,N_1218,N_1615);
and U2006 (N_2006,N_1225,N_1305);
xnor U2007 (N_2007,N_1256,N_1619);
or U2008 (N_2008,N_1031,N_1377);
xor U2009 (N_2009,N_1012,N_1825);
xnor U2010 (N_2010,N_1984,N_1043);
xor U2011 (N_2011,N_1086,N_1376);
nor U2012 (N_2012,N_1164,N_1903);
xor U2013 (N_2013,N_1966,N_1036);
nand U2014 (N_2014,N_1197,N_1963);
nand U2015 (N_2015,N_1271,N_1872);
and U2016 (N_2016,N_1022,N_1887);
xor U2017 (N_2017,N_1187,N_1250);
and U2018 (N_2018,N_1005,N_1252);
xnor U2019 (N_2019,N_1581,N_1843);
nor U2020 (N_2020,N_1653,N_1120);
or U2021 (N_2021,N_1964,N_1642);
xnor U2022 (N_2022,N_1142,N_1392);
or U2023 (N_2023,N_1794,N_1679);
xor U2024 (N_2024,N_1958,N_1447);
xnor U2025 (N_2025,N_1823,N_1522);
nand U2026 (N_2026,N_1994,N_1782);
nor U2027 (N_2027,N_1322,N_1884);
nor U2028 (N_2028,N_1982,N_1334);
and U2029 (N_2029,N_1803,N_1404);
nor U2030 (N_2030,N_1997,N_1620);
nand U2031 (N_2031,N_1544,N_1241);
and U2032 (N_2032,N_1071,N_1058);
and U2033 (N_2033,N_1283,N_1977);
and U2034 (N_2034,N_1152,N_1870);
and U2035 (N_2035,N_1590,N_1330);
or U2036 (N_2036,N_1659,N_1268);
nor U2037 (N_2037,N_1900,N_1698);
xor U2038 (N_2038,N_1180,N_1924);
or U2039 (N_2039,N_1747,N_1048);
or U2040 (N_2040,N_1101,N_1710);
xor U2041 (N_2041,N_1585,N_1859);
xnor U2042 (N_2042,N_1836,N_1243);
and U2043 (N_2043,N_1213,N_1867);
or U2044 (N_2044,N_1532,N_1652);
xor U2045 (N_2045,N_1403,N_1881);
or U2046 (N_2046,N_1076,N_1743);
and U2047 (N_2047,N_1636,N_1302);
and U2048 (N_2048,N_1774,N_1753);
nand U2049 (N_2049,N_1181,N_1196);
xnor U2050 (N_2050,N_1815,N_1928);
xor U2051 (N_2051,N_1795,N_1761);
nor U2052 (N_2052,N_1441,N_1971);
nor U2053 (N_2053,N_1347,N_1059);
and U2054 (N_2054,N_1510,N_1847);
xnor U2055 (N_2055,N_1809,N_1401);
nand U2056 (N_2056,N_1407,N_1054);
nor U2057 (N_2057,N_1968,N_1814);
and U2058 (N_2058,N_1443,N_1410);
nand U2059 (N_2059,N_1667,N_1008);
or U2060 (N_2060,N_1069,N_1981);
nand U2061 (N_2061,N_1226,N_1912);
nand U2062 (N_2062,N_1039,N_1154);
nand U2063 (N_2063,N_1433,N_1318);
nor U2064 (N_2064,N_1860,N_1098);
nor U2065 (N_2065,N_1995,N_1840);
and U2066 (N_2066,N_1408,N_1808);
and U2067 (N_2067,N_1858,N_1865);
nor U2068 (N_2068,N_1599,N_1432);
xor U2069 (N_2069,N_1260,N_1389);
or U2070 (N_2070,N_1360,N_1844);
or U2071 (N_2071,N_1270,N_1838);
nand U2072 (N_2072,N_1464,N_1788);
xor U2073 (N_2073,N_1215,N_1509);
nor U2074 (N_2074,N_1406,N_1845);
xor U2075 (N_2075,N_1656,N_1733);
nand U2076 (N_2076,N_1987,N_1300);
nand U2077 (N_2077,N_1853,N_1727);
xnor U2078 (N_2078,N_1276,N_1932);
nand U2079 (N_2079,N_1597,N_1923);
or U2080 (N_2080,N_1414,N_1399);
or U2081 (N_2081,N_1337,N_1346);
nand U2082 (N_2082,N_1341,N_1944);
nor U2083 (N_2083,N_1446,N_1244);
and U2084 (N_2084,N_1675,N_1415);
nand U2085 (N_2085,N_1251,N_1961);
and U2086 (N_2086,N_1499,N_1035);
or U2087 (N_2087,N_1933,N_1209);
nand U2088 (N_2088,N_1768,N_1385);
and U2089 (N_2089,N_1044,N_1264);
or U2090 (N_2090,N_1669,N_1574);
nand U2091 (N_2091,N_1624,N_1629);
nand U2092 (N_2092,N_1701,N_1792);
or U2093 (N_2093,N_1426,N_1632);
nand U2094 (N_2094,N_1224,N_1508);
and U2095 (N_2095,N_1553,N_1901);
nand U2096 (N_2096,N_1267,N_1092);
xor U2097 (N_2097,N_1413,N_1592);
xor U2098 (N_2098,N_1458,N_1866);
and U2099 (N_2099,N_1913,N_1748);
or U2100 (N_2100,N_1801,N_1400);
xnor U2101 (N_2101,N_1533,N_1411);
nor U2102 (N_2102,N_1909,N_1373);
or U2103 (N_2103,N_1505,N_1906);
and U2104 (N_2104,N_1545,N_1785);
and U2105 (N_2105,N_1947,N_1674);
nor U2106 (N_2106,N_1393,N_1115);
nor U2107 (N_2107,N_1638,N_1999);
xor U2108 (N_2108,N_1055,N_1145);
or U2109 (N_2109,N_1042,N_1163);
xnor U2110 (N_2110,N_1498,N_1851);
nand U2111 (N_2111,N_1061,N_1731);
nand U2112 (N_2112,N_1095,N_1594);
nor U2113 (N_2113,N_1975,N_1097);
and U2114 (N_2114,N_1375,N_1325);
nor U2115 (N_2115,N_1294,N_1649);
and U2116 (N_2116,N_1333,N_1527);
or U2117 (N_2117,N_1462,N_1626);
xnor U2118 (N_2118,N_1320,N_1538);
xnor U2119 (N_2119,N_1504,N_1986);
nand U2120 (N_2120,N_1328,N_1461);
nand U2121 (N_2121,N_1451,N_1724);
and U2122 (N_2122,N_1770,N_1053);
nor U2123 (N_2123,N_1279,N_1348);
or U2124 (N_2124,N_1262,N_1475);
xor U2125 (N_2125,N_1796,N_1350);
nand U2126 (N_2126,N_1396,N_1526);
and U2127 (N_2127,N_1316,N_1466);
or U2128 (N_2128,N_1745,N_1146);
nor U2129 (N_2129,N_1824,N_1166);
nand U2130 (N_2130,N_1078,N_1848);
and U2131 (N_2131,N_1790,N_1291);
nand U2132 (N_2132,N_1380,N_1394);
nor U2133 (N_2133,N_1205,N_1474);
xor U2134 (N_2134,N_1635,N_1183);
or U2135 (N_2135,N_1106,N_1217);
nand U2136 (N_2136,N_1352,N_1939);
xor U2137 (N_2137,N_1425,N_1686);
and U2138 (N_2138,N_1203,N_1628);
nor U2139 (N_2139,N_1714,N_1861);
nand U2140 (N_2140,N_1662,N_1562);
xor U2141 (N_2141,N_1873,N_1737);
and U2142 (N_2142,N_1816,N_1436);
nor U2143 (N_2143,N_1519,N_1936);
and U2144 (N_2144,N_1927,N_1694);
nor U2145 (N_2145,N_1489,N_1885);
nor U2146 (N_2146,N_1416,N_1613);
nand U2147 (N_2147,N_1969,N_1650);
and U2148 (N_2148,N_1133,N_1530);
and U2149 (N_2149,N_1550,N_1754);
nor U2150 (N_2150,N_1176,N_1729);
xor U2151 (N_2151,N_1678,N_1471);
and U2152 (N_2152,N_1332,N_1494);
nor U2153 (N_2153,N_1324,N_1758);
nand U2154 (N_2154,N_1085,N_1470);
xnor U2155 (N_2155,N_1240,N_1093);
xnor U2156 (N_2156,N_1220,N_1194);
nor U2157 (N_2157,N_1045,N_1552);
nand U2158 (N_2158,N_1204,N_1871);
or U2159 (N_2159,N_1614,N_1455);
xnor U2160 (N_2160,N_1281,N_1088);
or U2161 (N_2161,N_1911,N_1564);
xor U2162 (N_2162,N_1769,N_1070);
and U2163 (N_2163,N_1783,N_1132);
or U2164 (N_2164,N_1517,N_1630);
or U2165 (N_2165,N_1940,N_1955);
or U2166 (N_2166,N_1952,N_1682);
and U2167 (N_2167,N_1431,N_1915);
xnor U2168 (N_2168,N_1398,N_1980);
nand U2169 (N_2169,N_1049,N_1208);
and U2170 (N_2170,N_1547,N_1248);
and U2171 (N_2171,N_1560,N_1864);
nor U2172 (N_2172,N_1643,N_1116);
and U2173 (N_2173,N_1065,N_1503);
xnor U2174 (N_2174,N_1779,N_1402);
or U2175 (N_2175,N_1771,N_1622);
xor U2176 (N_2176,N_1772,N_1569);
nor U2177 (N_2177,N_1200,N_1245);
and U2178 (N_2178,N_1894,N_1368);
nand U2179 (N_2179,N_1391,N_1566);
nor U2180 (N_2180,N_1908,N_1702);
and U2181 (N_2181,N_1949,N_1563);
nor U2182 (N_2182,N_1287,N_1136);
nor U2183 (N_2183,N_1728,N_1606);
and U2184 (N_2184,N_1506,N_1542);
and U2185 (N_2185,N_1645,N_1354);
nand U2186 (N_2186,N_1723,N_1387);
xor U2187 (N_2187,N_1068,N_1237);
or U2188 (N_2188,N_1288,N_1551);
or U2189 (N_2189,N_1732,N_1023);
nand U2190 (N_2190,N_1671,N_1535);
xor U2191 (N_2191,N_1129,N_1979);
nand U2192 (N_2192,N_1060,N_1390);
and U2193 (N_2193,N_1625,N_1442);
or U2194 (N_2194,N_1295,N_1935);
or U2195 (N_2195,N_1378,N_1063);
or U2196 (N_2196,N_1427,N_1018);
xnor U2197 (N_2197,N_1588,N_1835);
nand U2198 (N_2198,N_1718,N_1278);
or U2199 (N_2199,N_1658,N_1104);
or U2200 (N_2200,N_1306,N_1258);
and U2201 (N_2201,N_1050,N_1382);
or U2202 (N_2202,N_1970,N_1962);
or U2203 (N_2203,N_1191,N_1780);
nand U2204 (N_2204,N_1110,N_1673);
or U2205 (N_2205,N_1155,N_1277);
nand U2206 (N_2206,N_1491,N_1323);
nand U2207 (N_2207,N_1990,N_1537);
or U2208 (N_2208,N_1034,N_1459);
and U2209 (N_2209,N_1863,N_1734);
and U2210 (N_2210,N_1046,N_1440);
nand U2211 (N_2211,N_1751,N_1293);
or U2212 (N_2212,N_1381,N_1171);
or U2213 (N_2213,N_1307,N_1107);
or U2214 (N_2214,N_1598,N_1668);
xnor U2215 (N_2215,N_1549,N_1127);
xnor U2216 (N_2216,N_1430,N_1898);
nor U2217 (N_2217,N_1299,N_1880);
xor U2218 (N_2218,N_1239,N_1138);
or U2219 (N_2219,N_1170,N_1317);
nand U2220 (N_2220,N_1819,N_1153);
xnor U2221 (N_2221,N_1789,N_1363);
xor U2222 (N_2222,N_1570,N_1914);
and U2223 (N_2223,N_1917,N_1744);
xnor U2224 (N_2224,N_1822,N_1000);
nor U2225 (N_2225,N_1326,N_1664);
nand U2226 (N_2226,N_1309,N_1760);
xor U2227 (N_2227,N_1931,N_1827);
and U2228 (N_2228,N_1015,N_1072);
nor U2229 (N_2229,N_1140,N_1263);
and U2230 (N_2230,N_1715,N_1134);
and U2231 (N_2231,N_1160,N_1201);
and U2232 (N_2232,N_1879,N_1946);
and U2233 (N_2233,N_1611,N_1223);
nor U2234 (N_2234,N_1806,N_1910);
nor U2235 (N_2235,N_1026,N_1296);
or U2236 (N_2236,N_1988,N_1817);
and U2237 (N_2237,N_1959,N_1482);
nor U2238 (N_2238,N_1998,N_1766);
nor U2239 (N_2239,N_1297,N_1301);
nor U2240 (N_2240,N_1705,N_1595);
nor U2241 (N_2241,N_1463,N_1147);
xnor U2242 (N_2242,N_1228,N_1178);
and U2243 (N_2243,N_1417,N_1591);
or U2244 (N_2244,N_1948,N_1805);
and U2245 (N_2245,N_1736,N_1168);
and U2246 (N_2246,N_1868,N_1521);
and U2247 (N_2247,N_1681,N_1478);
nand U2248 (N_2248,N_1942,N_1916);
and U2249 (N_2249,N_1434,N_1100);
nand U2250 (N_2250,N_1135,N_1090);
xnor U2251 (N_2251,N_1730,N_1144);
nor U2252 (N_2252,N_1830,N_1338);
or U2253 (N_2253,N_1472,N_1460);
xnor U2254 (N_2254,N_1787,N_1339);
and U2255 (N_2255,N_1003,N_1310);
nor U2256 (N_2256,N_1195,N_1738);
or U2257 (N_2257,N_1047,N_1265);
xor U2258 (N_2258,N_1477,N_1212);
nor U2259 (N_2259,N_1584,N_1660);
xor U2260 (N_2260,N_1921,N_1030);
xnor U2261 (N_2261,N_1083,N_1193);
xnor U2262 (N_2262,N_1081,N_1837);
or U2263 (N_2263,N_1541,N_1888);
nor U2264 (N_2264,N_1128,N_1199);
xnor U2265 (N_2265,N_1604,N_1561);
xor U2266 (N_2266,N_1041,N_1109);
nand U2267 (N_2267,N_1148,N_1409);
xor U2268 (N_2268,N_1358,N_1749);
and U2269 (N_2269,N_1716,N_1689);
nand U2270 (N_2270,N_1102,N_1169);
and U2271 (N_2271,N_1516,N_1422);
nand U2272 (N_2272,N_1014,N_1112);
or U2273 (N_2273,N_1143,N_1937);
nor U2274 (N_2274,N_1335,N_1009);
nand U2275 (N_2275,N_1253,N_1395);
or U2276 (N_2276,N_1874,N_1511);
and U2277 (N_2277,N_1465,N_1829);
xor U2278 (N_2278,N_1943,N_1740);
xor U2279 (N_2279,N_1897,N_1839);
or U2280 (N_2280,N_1647,N_1528);
and U2281 (N_2281,N_1087,N_1037);
or U2282 (N_2282,N_1017,N_1807);
and U2283 (N_2283,N_1159,N_1985);
and U2284 (N_2284,N_1567,N_1272);
xor U2285 (N_2285,N_1355,N_1314);
or U2286 (N_2286,N_1878,N_1158);
xor U2287 (N_2287,N_1895,N_1137);
or U2288 (N_2288,N_1211,N_1439);
nor U2289 (N_2289,N_1711,N_1520);
nand U2290 (N_2290,N_1756,N_1820);
or U2291 (N_2291,N_1691,N_1531);
nor U2292 (N_2292,N_1372,N_1596);
nand U2293 (N_2293,N_1618,N_1586);
nand U2294 (N_2294,N_1812,N_1074);
nor U2295 (N_2295,N_1665,N_1122);
or U2296 (N_2296,N_1692,N_1139);
and U2297 (N_2297,N_1362,N_1290);
nor U2298 (N_2298,N_1627,N_1210);
xor U2299 (N_2299,N_1412,N_1367);
nor U2300 (N_2300,N_1266,N_1445);
and U2301 (N_2301,N_1704,N_1573);
or U2302 (N_2302,N_1684,N_1685);
xor U2303 (N_2303,N_1275,N_1548);
nand U2304 (N_2304,N_1468,N_1755);
nand U2305 (N_2305,N_1182,N_1697);
nor U2306 (N_2306,N_1721,N_1846);
xnor U2307 (N_2307,N_1875,N_1831);
nand U2308 (N_2308,N_1905,N_1540);
and U2309 (N_2309,N_1189,N_1007);
xor U2310 (N_2310,N_1001,N_1918);
and U2311 (N_2311,N_1216,N_1173);
or U2312 (N_2312,N_1856,N_1453);
xnor U2313 (N_2313,N_1648,N_1304);
or U2314 (N_2314,N_1119,N_1123);
and U2315 (N_2315,N_1696,N_1719);
or U2316 (N_2316,N_1234,N_1800);
xnor U2317 (N_2317,N_1105,N_1108);
nor U2318 (N_2318,N_1577,N_1423);
or U2319 (N_2319,N_1568,N_1600);
and U2320 (N_2320,N_1991,N_1002);
xnor U2321 (N_2321,N_1725,N_1004);
or U2322 (N_2322,N_1666,N_1616);
nand U2323 (N_2323,N_1424,N_1013);
and U2324 (N_2324,N_1483,N_1557);
and U2325 (N_2325,N_1384,N_1469);
and U2326 (N_2326,N_1500,N_1261);
nand U2327 (N_2327,N_1821,N_1051);
or U2328 (N_2328,N_1623,N_1739);
or U2329 (N_2329,N_1956,N_1292);
or U2330 (N_2330,N_1767,N_1572);
nand U2331 (N_2331,N_1512,N_1490);
nand U2332 (N_2332,N_1811,N_1038);
nand U2333 (N_2333,N_1633,N_1883);
and U2334 (N_2334,N_1765,N_1593);
and U2335 (N_2335,N_1124,N_1327);
nand U2336 (N_2336,N_1534,N_1989);
and U2337 (N_2337,N_1742,N_1951);
nor U2338 (N_2338,N_1269,N_1945);
nor U2339 (N_2339,N_1342,N_1797);
nand U2340 (N_2340,N_1695,N_1331);
xor U2341 (N_2341,N_1383,N_1082);
nand U2342 (N_2342,N_1973,N_1361);
nand U2343 (N_2343,N_1448,N_1161);
nand U2344 (N_2344,N_1273,N_1907);
or U2345 (N_2345,N_1713,N_1198);
or U2346 (N_2346,N_1285,N_1556);
xnor U2347 (N_2347,N_1523,N_1712);
or U2348 (N_2348,N_1693,N_1364);
and U2349 (N_2349,N_1481,N_1663);
and U2350 (N_2350,N_1978,N_1813);
nand U2351 (N_2351,N_1062,N_1850);
nand U2352 (N_2352,N_1099,N_1974);
nand U2353 (N_2353,N_1896,N_1834);
or U2354 (N_2354,N_1759,N_1524);
nand U2355 (N_2355,N_1336,N_1902);
xor U2356 (N_2356,N_1676,N_1492);
or U2357 (N_2357,N_1890,N_1575);
nand U2358 (N_2358,N_1020,N_1476);
or U2359 (N_2359,N_1683,N_1891);
nand U2360 (N_2360,N_1131,N_1379);
nor U2361 (N_2361,N_1941,N_1456);
nand U2362 (N_2362,N_1688,N_1487);
xor U2363 (N_2363,N_1670,N_1227);
xor U2364 (N_2364,N_1365,N_1750);
xnor U2365 (N_2365,N_1162,N_1479);
nand U2366 (N_2366,N_1094,N_1315);
nor U2367 (N_2367,N_1735,N_1202);
or U2368 (N_2368,N_1603,N_1103);
or U2369 (N_2369,N_1558,N_1621);
or U2370 (N_2370,N_1125,N_1993);
xnor U2371 (N_2371,N_1206,N_1904);
and U2372 (N_2372,N_1610,N_1651);
or U2373 (N_2373,N_1920,N_1117);
xor U2374 (N_2374,N_1882,N_1953);
nor U2375 (N_2375,N_1113,N_1777);
nand U2376 (N_2376,N_1057,N_1514);
nand U2377 (N_2377,N_1793,N_1954);
nand U2378 (N_2378,N_1862,N_1033);
nor U2379 (N_2379,N_1231,N_1639);
xnor U2380 (N_2380,N_1156,N_1501);
or U2381 (N_2381,N_1605,N_1799);
or U2382 (N_2382,N_1687,N_1021);
or U2383 (N_2383,N_1452,N_1444);
xor U2384 (N_2384,N_1539,N_1321);
or U2385 (N_2385,N_1717,N_1089);
nor U2386 (N_2386,N_1222,N_1832);
xor U2387 (N_2387,N_1587,N_1852);
or U2388 (N_2388,N_1925,N_1019);
and U2389 (N_2389,N_1221,N_1370);
or U2390 (N_2390,N_1286,N_1157);
xor U2391 (N_2391,N_1421,N_1810);
or U2392 (N_2392,N_1190,N_1654);
or U2393 (N_2393,N_1757,N_1763);
nand U2394 (N_2394,N_1366,N_1340);
nand U2395 (N_2395,N_1996,N_1344);
nor U2396 (N_2396,N_1064,N_1006);
nand U2397 (N_2397,N_1893,N_1353);
nor U2398 (N_2398,N_1525,N_1778);
or U2399 (N_2399,N_1418,N_1680);
nand U2400 (N_2400,N_1255,N_1518);
xnor U2401 (N_2401,N_1308,N_1067);
and U2402 (N_2402,N_1298,N_1828);
nor U2403 (N_2403,N_1454,N_1709);
xor U2404 (N_2404,N_1786,N_1972);
xor U2405 (N_2405,N_1467,N_1329);
or U2406 (N_2406,N_1589,N_1485);
or U2407 (N_2407,N_1752,N_1515);
or U2408 (N_2408,N_1284,N_1631);
xnor U2409 (N_2409,N_1079,N_1976);
nor U2410 (N_2410,N_1857,N_1056);
nor U2411 (N_2411,N_1764,N_1235);
xor U2412 (N_2412,N_1185,N_1165);
nor U2413 (N_2413,N_1926,N_1579);
xor U2414 (N_2414,N_1929,N_1207);
nand U2415 (N_2415,N_1349,N_1282);
or U2416 (N_2416,N_1254,N_1559);
xnor U2417 (N_2417,N_1121,N_1934);
xor U2418 (N_2418,N_1289,N_1232);
nor U2419 (N_2419,N_1641,N_1661);
or U2420 (N_2420,N_1967,N_1259);
nand U2421 (N_2421,N_1877,N_1690);
or U2422 (N_2422,N_1798,N_1229);
nand U2423 (N_2423,N_1899,N_1151);
and U2424 (N_2424,N_1554,N_1703);
nor U2425 (N_2425,N_1480,N_1818);
xnor U2426 (N_2426,N_1726,N_1922);
or U2427 (N_2427,N_1114,N_1343);
nand U2428 (N_2428,N_1497,N_1960);
and U2429 (N_2429,N_1437,N_1543);
nor U2430 (N_2430,N_1186,N_1672);
and U2431 (N_2431,N_1077,N_1236);
or U2432 (N_2432,N_1488,N_1486);
nor U2433 (N_2433,N_1174,N_1345);
xnor U2434 (N_2434,N_1580,N_1886);
xnor U2435 (N_2435,N_1319,N_1011);
nand U2436 (N_2436,N_1802,N_1230);
or U2437 (N_2437,N_1889,N_1040);
nor U2438 (N_2438,N_1849,N_1435);
xor U2439 (N_2439,N_1919,N_1438);
nand U2440 (N_2440,N_1833,N_1371);
nor U2441 (N_2441,N_1141,N_1555);
nand U2442 (N_2442,N_1111,N_1706);
nand U2443 (N_2443,N_1762,N_1930);
nor U2444 (N_2444,N_1091,N_1130);
xor U2445 (N_2445,N_1495,N_1311);
and U2446 (N_2446,N_1720,N_1214);
or U2447 (N_2447,N_1084,N_1576);
and U2448 (N_2448,N_1374,N_1242);
or U2449 (N_2449,N_1388,N_1369);
nand U2450 (N_2450,N_1175,N_1397);
xnor U2451 (N_2451,N_1722,N_1776);
nor U2452 (N_2452,N_1855,N_1617);
nand U2453 (N_2453,N_1841,N_1983);
or U2454 (N_2454,N_1637,N_1303);
or U2455 (N_2455,N_1657,N_1842);
nor U2456 (N_2456,N_1450,N_1791);
nand U2457 (N_2457,N_1938,N_1096);
xor U2458 (N_2458,N_1177,N_1457);
xnor U2459 (N_2459,N_1167,N_1513);
or U2460 (N_2460,N_1507,N_1781);
or U2461 (N_2461,N_1010,N_1646);
or U2462 (N_2462,N_1699,N_1149);
and U2463 (N_2463,N_1428,N_1219);
nand U2464 (N_2464,N_1677,N_1357);
nand U2465 (N_2465,N_1950,N_1238);
and U2466 (N_2466,N_1028,N_1172);
xor U2467 (N_2467,N_1280,N_1601);
or U2468 (N_2468,N_1233,N_1608);
nand U2469 (N_2469,N_1640,N_1386);
xnor U2470 (N_2470,N_1746,N_1536);
nor U2471 (N_2471,N_1192,N_1420);
xor U2472 (N_2472,N_1607,N_1546);
or U2473 (N_2473,N_1578,N_1741);
xor U2474 (N_2474,N_1957,N_1405);
and U2475 (N_2475,N_1773,N_1356);
and U2476 (N_2476,N_1351,N_1016);
nor U2477 (N_2477,N_1025,N_1080);
nand U2478 (N_2478,N_1073,N_1571);
or U2479 (N_2479,N_1027,N_1493);
xnor U2480 (N_2480,N_1582,N_1246);
or U2481 (N_2481,N_1965,N_1707);
nor U2482 (N_2482,N_1876,N_1188);
nand U2483 (N_2483,N_1854,N_1312);
nor U2484 (N_2484,N_1052,N_1249);
xor U2485 (N_2485,N_1419,N_1529);
or U2486 (N_2486,N_1502,N_1359);
or U2487 (N_2487,N_1429,N_1826);
nor U2488 (N_2488,N_1029,N_1247);
nand U2489 (N_2489,N_1126,N_1313);
nor U2490 (N_2490,N_1496,N_1804);
or U2491 (N_2491,N_1449,N_1150);
or U2492 (N_2492,N_1179,N_1484);
and U2493 (N_2493,N_1869,N_1602);
or U2494 (N_2494,N_1118,N_1644);
and U2495 (N_2495,N_1634,N_1473);
or U2496 (N_2496,N_1609,N_1583);
nand U2497 (N_2497,N_1032,N_1274);
nor U2498 (N_2498,N_1612,N_1775);
and U2499 (N_2499,N_1700,N_1257);
nor U2500 (N_2500,N_1852,N_1188);
xnor U2501 (N_2501,N_1652,N_1671);
xor U2502 (N_2502,N_1575,N_1682);
nor U2503 (N_2503,N_1954,N_1378);
nor U2504 (N_2504,N_1102,N_1918);
or U2505 (N_2505,N_1646,N_1923);
nand U2506 (N_2506,N_1546,N_1525);
and U2507 (N_2507,N_1104,N_1355);
or U2508 (N_2508,N_1092,N_1392);
and U2509 (N_2509,N_1551,N_1155);
or U2510 (N_2510,N_1435,N_1067);
xnor U2511 (N_2511,N_1270,N_1874);
nand U2512 (N_2512,N_1348,N_1444);
and U2513 (N_2513,N_1226,N_1295);
nand U2514 (N_2514,N_1913,N_1224);
nand U2515 (N_2515,N_1001,N_1723);
nor U2516 (N_2516,N_1304,N_1742);
nand U2517 (N_2517,N_1781,N_1063);
or U2518 (N_2518,N_1799,N_1023);
nor U2519 (N_2519,N_1465,N_1624);
or U2520 (N_2520,N_1377,N_1128);
and U2521 (N_2521,N_1849,N_1075);
nor U2522 (N_2522,N_1189,N_1211);
nand U2523 (N_2523,N_1323,N_1805);
and U2524 (N_2524,N_1399,N_1651);
or U2525 (N_2525,N_1945,N_1481);
nand U2526 (N_2526,N_1140,N_1108);
nand U2527 (N_2527,N_1443,N_1315);
nand U2528 (N_2528,N_1364,N_1583);
xor U2529 (N_2529,N_1430,N_1569);
xnor U2530 (N_2530,N_1472,N_1811);
xnor U2531 (N_2531,N_1856,N_1916);
or U2532 (N_2532,N_1366,N_1898);
or U2533 (N_2533,N_1004,N_1707);
and U2534 (N_2534,N_1249,N_1635);
and U2535 (N_2535,N_1041,N_1104);
nand U2536 (N_2536,N_1174,N_1068);
xnor U2537 (N_2537,N_1086,N_1491);
and U2538 (N_2538,N_1495,N_1041);
or U2539 (N_2539,N_1269,N_1601);
nand U2540 (N_2540,N_1327,N_1043);
or U2541 (N_2541,N_1963,N_1960);
nand U2542 (N_2542,N_1755,N_1390);
nand U2543 (N_2543,N_1480,N_1207);
nand U2544 (N_2544,N_1902,N_1915);
xnor U2545 (N_2545,N_1946,N_1283);
or U2546 (N_2546,N_1944,N_1384);
nand U2547 (N_2547,N_1047,N_1868);
or U2548 (N_2548,N_1107,N_1600);
and U2549 (N_2549,N_1547,N_1637);
or U2550 (N_2550,N_1175,N_1131);
xnor U2551 (N_2551,N_1937,N_1700);
xor U2552 (N_2552,N_1107,N_1921);
nor U2553 (N_2553,N_1337,N_1296);
or U2554 (N_2554,N_1246,N_1700);
xor U2555 (N_2555,N_1429,N_1641);
or U2556 (N_2556,N_1924,N_1542);
and U2557 (N_2557,N_1604,N_1740);
nor U2558 (N_2558,N_1236,N_1841);
nor U2559 (N_2559,N_1305,N_1188);
and U2560 (N_2560,N_1819,N_1022);
nor U2561 (N_2561,N_1877,N_1560);
and U2562 (N_2562,N_1399,N_1753);
nor U2563 (N_2563,N_1057,N_1035);
nor U2564 (N_2564,N_1516,N_1919);
xor U2565 (N_2565,N_1856,N_1983);
or U2566 (N_2566,N_1958,N_1436);
nor U2567 (N_2567,N_1282,N_1501);
and U2568 (N_2568,N_1740,N_1651);
or U2569 (N_2569,N_1760,N_1058);
or U2570 (N_2570,N_1037,N_1557);
xor U2571 (N_2571,N_1492,N_1519);
and U2572 (N_2572,N_1582,N_1194);
nand U2573 (N_2573,N_1083,N_1380);
xor U2574 (N_2574,N_1790,N_1146);
nand U2575 (N_2575,N_1916,N_1850);
nand U2576 (N_2576,N_1507,N_1954);
nand U2577 (N_2577,N_1345,N_1247);
nor U2578 (N_2578,N_1206,N_1013);
or U2579 (N_2579,N_1896,N_1249);
nand U2580 (N_2580,N_1091,N_1694);
or U2581 (N_2581,N_1661,N_1407);
and U2582 (N_2582,N_1199,N_1390);
and U2583 (N_2583,N_1073,N_1513);
xnor U2584 (N_2584,N_1153,N_1719);
xor U2585 (N_2585,N_1570,N_1217);
nor U2586 (N_2586,N_1481,N_1121);
and U2587 (N_2587,N_1535,N_1593);
nand U2588 (N_2588,N_1167,N_1932);
and U2589 (N_2589,N_1632,N_1893);
nor U2590 (N_2590,N_1640,N_1011);
xor U2591 (N_2591,N_1228,N_1743);
and U2592 (N_2592,N_1627,N_1214);
and U2593 (N_2593,N_1319,N_1828);
nand U2594 (N_2594,N_1915,N_1073);
and U2595 (N_2595,N_1857,N_1208);
nand U2596 (N_2596,N_1112,N_1909);
nor U2597 (N_2597,N_1943,N_1872);
or U2598 (N_2598,N_1556,N_1220);
nor U2599 (N_2599,N_1910,N_1713);
or U2600 (N_2600,N_1838,N_1828);
or U2601 (N_2601,N_1211,N_1992);
nand U2602 (N_2602,N_1450,N_1203);
xor U2603 (N_2603,N_1695,N_1275);
xor U2604 (N_2604,N_1913,N_1477);
or U2605 (N_2605,N_1400,N_1527);
nand U2606 (N_2606,N_1073,N_1540);
nor U2607 (N_2607,N_1890,N_1263);
nor U2608 (N_2608,N_1275,N_1670);
or U2609 (N_2609,N_1932,N_1257);
nand U2610 (N_2610,N_1928,N_1435);
and U2611 (N_2611,N_1986,N_1809);
xnor U2612 (N_2612,N_1537,N_1411);
or U2613 (N_2613,N_1446,N_1151);
nor U2614 (N_2614,N_1964,N_1359);
or U2615 (N_2615,N_1016,N_1488);
nor U2616 (N_2616,N_1344,N_1742);
nand U2617 (N_2617,N_1620,N_1300);
nand U2618 (N_2618,N_1218,N_1857);
xor U2619 (N_2619,N_1769,N_1310);
nor U2620 (N_2620,N_1011,N_1198);
nor U2621 (N_2621,N_1614,N_1554);
nand U2622 (N_2622,N_1663,N_1900);
nor U2623 (N_2623,N_1835,N_1569);
or U2624 (N_2624,N_1371,N_1825);
nand U2625 (N_2625,N_1301,N_1125);
and U2626 (N_2626,N_1945,N_1061);
nand U2627 (N_2627,N_1561,N_1095);
and U2628 (N_2628,N_1610,N_1577);
and U2629 (N_2629,N_1631,N_1759);
nand U2630 (N_2630,N_1084,N_1022);
nor U2631 (N_2631,N_1422,N_1797);
and U2632 (N_2632,N_1197,N_1974);
xnor U2633 (N_2633,N_1019,N_1558);
nor U2634 (N_2634,N_1914,N_1039);
nor U2635 (N_2635,N_1416,N_1003);
nor U2636 (N_2636,N_1462,N_1820);
and U2637 (N_2637,N_1139,N_1559);
nor U2638 (N_2638,N_1550,N_1552);
xor U2639 (N_2639,N_1050,N_1549);
xnor U2640 (N_2640,N_1575,N_1404);
or U2641 (N_2641,N_1223,N_1129);
xor U2642 (N_2642,N_1488,N_1806);
xnor U2643 (N_2643,N_1923,N_1121);
nand U2644 (N_2644,N_1048,N_1921);
and U2645 (N_2645,N_1991,N_1955);
nand U2646 (N_2646,N_1869,N_1153);
nor U2647 (N_2647,N_1353,N_1546);
xnor U2648 (N_2648,N_1270,N_1953);
nor U2649 (N_2649,N_1242,N_1549);
or U2650 (N_2650,N_1880,N_1547);
and U2651 (N_2651,N_1480,N_1226);
nor U2652 (N_2652,N_1249,N_1098);
nand U2653 (N_2653,N_1896,N_1696);
nand U2654 (N_2654,N_1795,N_1222);
xnor U2655 (N_2655,N_1069,N_1052);
xnor U2656 (N_2656,N_1822,N_1128);
and U2657 (N_2657,N_1281,N_1181);
and U2658 (N_2658,N_1737,N_1986);
xor U2659 (N_2659,N_1935,N_1714);
nand U2660 (N_2660,N_1002,N_1262);
and U2661 (N_2661,N_1952,N_1640);
xor U2662 (N_2662,N_1047,N_1965);
nor U2663 (N_2663,N_1030,N_1981);
and U2664 (N_2664,N_1148,N_1735);
xor U2665 (N_2665,N_1878,N_1776);
nand U2666 (N_2666,N_1869,N_1552);
xor U2667 (N_2667,N_1165,N_1597);
xor U2668 (N_2668,N_1856,N_1520);
xor U2669 (N_2669,N_1342,N_1414);
or U2670 (N_2670,N_1144,N_1399);
or U2671 (N_2671,N_1426,N_1773);
xor U2672 (N_2672,N_1403,N_1424);
or U2673 (N_2673,N_1437,N_1709);
and U2674 (N_2674,N_1528,N_1016);
and U2675 (N_2675,N_1451,N_1400);
nor U2676 (N_2676,N_1186,N_1930);
and U2677 (N_2677,N_1147,N_1307);
nor U2678 (N_2678,N_1019,N_1317);
xnor U2679 (N_2679,N_1109,N_1634);
nand U2680 (N_2680,N_1442,N_1569);
and U2681 (N_2681,N_1340,N_1976);
nand U2682 (N_2682,N_1216,N_1374);
nand U2683 (N_2683,N_1408,N_1667);
nand U2684 (N_2684,N_1165,N_1179);
or U2685 (N_2685,N_1442,N_1134);
or U2686 (N_2686,N_1955,N_1319);
xnor U2687 (N_2687,N_1642,N_1622);
and U2688 (N_2688,N_1351,N_1955);
or U2689 (N_2689,N_1913,N_1191);
or U2690 (N_2690,N_1460,N_1831);
and U2691 (N_2691,N_1381,N_1636);
and U2692 (N_2692,N_1148,N_1237);
and U2693 (N_2693,N_1240,N_1373);
or U2694 (N_2694,N_1851,N_1976);
nand U2695 (N_2695,N_1964,N_1844);
and U2696 (N_2696,N_1239,N_1145);
and U2697 (N_2697,N_1857,N_1706);
nor U2698 (N_2698,N_1346,N_1030);
and U2699 (N_2699,N_1039,N_1132);
xor U2700 (N_2700,N_1573,N_1431);
xnor U2701 (N_2701,N_1787,N_1803);
and U2702 (N_2702,N_1923,N_1939);
nor U2703 (N_2703,N_1113,N_1139);
or U2704 (N_2704,N_1003,N_1820);
or U2705 (N_2705,N_1784,N_1431);
xnor U2706 (N_2706,N_1592,N_1528);
xnor U2707 (N_2707,N_1770,N_1816);
and U2708 (N_2708,N_1246,N_1692);
xnor U2709 (N_2709,N_1322,N_1389);
or U2710 (N_2710,N_1730,N_1470);
xnor U2711 (N_2711,N_1536,N_1607);
xor U2712 (N_2712,N_1916,N_1872);
nor U2713 (N_2713,N_1792,N_1034);
nand U2714 (N_2714,N_1556,N_1078);
nand U2715 (N_2715,N_1927,N_1012);
or U2716 (N_2716,N_1602,N_1788);
nor U2717 (N_2717,N_1656,N_1882);
and U2718 (N_2718,N_1703,N_1663);
or U2719 (N_2719,N_1331,N_1160);
nand U2720 (N_2720,N_1469,N_1126);
xnor U2721 (N_2721,N_1303,N_1313);
xor U2722 (N_2722,N_1506,N_1538);
nor U2723 (N_2723,N_1977,N_1437);
nor U2724 (N_2724,N_1403,N_1297);
nor U2725 (N_2725,N_1501,N_1600);
or U2726 (N_2726,N_1860,N_1487);
and U2727 (N_2727,N_1161,N_1619);
and U2728 (N_2728,N_1129,N_1298);
xnor U2729 (N_2729,N_1206,N_1316);
or U2730 (N_2730,N_1322,N_1467);
or U2731 (N_2731,N_1270,N_1274);
or U2732 (N_2732,N_1627,N_1354);
or U2733 (N_2733,N_1285,N_1048);
and U2734 (N_2734,N_1830,N_1048);
nor U2735 (N_2735,N_1131,N_1640);
nor U2736 (N_2736,N_1627,N_1910);
nor U2737 (N_2737,N_1810,N_1342);
or U2738 (N_2738,N_1560,N_1507);
xor U2739 (N_2739,N_1083,N_1635);
and U2740 (N_2740,N_1620,N_1592);
nor U2741 (N_2741,N_1137,N_1096);
and U2742 (N_2742,N_1362,N_1638);
xor U2743 (N_2743,N_1312,N_1493);
or U2744 (N_2744,N_1741,N_1675);
nor U2745 (N_2745,N_1973,N_1241);
and U2746 (N_2746,N_1408,N_1542);
or U2747 (N_2747,N_1921,N_1908);
or U2748 (N_2748,N_1427,N_1526);
nor U2749 (N_2749,N_1719,N_1406);
and U2750 (N_2750,N_1604,N_1668);
or U2751 (N_2751,N_1937,N_1856);
and U2752 (N_2752,N_1911,N_1190);
nand U2753 (N_2753,N_1585,N_1980);
and U2754 (N_2754,N_1390,N_1792);
nand U2755 (N_2755,N_1640,N_1821);
nor U2756 (N_2756,N_1392,N_1211);
and U2757 (N_2757,N_1754,N_1400);
nor U2758 (N_2758,N_1749,N_1875);
and U2759 (N_2759,N_1255,N_1165);
or U2760 (N_2760,N_1428,N_1545);
nor U2761 (N_2761,N_1191,N_1094);
and U2762 (N_2762,N_1853,N_1089);
nor U2763 (N_2763,N_1887,N_1517);
nor U2764 (N_2764,N_1905,N_1789);
nand U2765 (N_2765,N_1713,N_1077);
nor U2766 (N_2766,N_1537,N_1476);
and U2767 (N_2767,N_1969,N_1717);
nand U2768 (N_2768,N_1236,N_1738);
and U2769 (N_2769,N_1278,N_1874);
nor U2770 (N_2770,N_1991,N_1408);
nor U2771 (N_2771,N_1808,N_1860);
xor U2772 (N_2772,N_1186,N_1161);
or U2773 (N_2773,N_1162,N_1128);
nand U2774 (N_2774,N_1544,N_1734);
nor U2775 (N_2775,N_1028,N_1510);
nor U2776 (N_2776,N_1489,N_1987);
and U2777 (N_2777,N_1008,N_1967);
and U2778 (N_2778,N_1420,N_1952);
xor U2779 (N_2779,N_1404,N_1590);
xnor U2780 (N_2780,N_1071,N_1269);
or U2781 (N_2781,N_1816,N_1056);
nor U2782 (N_2782,N_1245,N_1773);
nand U2783 (N_2783,N_1510,N_1334);
and U2784 (N_2784,N_1287,N_1904);
or U2785 (N_2785,N_1577,N_1154);
xnor U2786 (N_2786,N_1028,N_1164);
nor U2787 (N_2787,N_1305,N_1690);
xnor U2788 (N_2788,N_1560,N_1205);
nand U2789 (N_2789,N_1246,N_1673);
and U2790 (N_2790,N_1858,N_1232);
or U2791 (N_2791,N_1719,N_1323);
nand U2792 (N_2792,N_1629,N_1574);
nand U2793 (N_2793,N_1754,N_1804);
and U2794 (N_2794,N_1864,N_1546);
nand U2795 (N_2795,N_1789,N_1230);
xnor U2796 (N_2796,N_1161,N_1617);
and U2797 (N_2797,N_1101,N_1768);
or U2798 (N_2798,N_1753,N_1671);
xor U2799 (N_2799,N_1954,N_1073);
and U2800 (N_2800,N_1158,N_1435);
or U2801 (N_2801,N_1770,N_1604);
nand U2802 (N_2802,N_1403,N_1687);
nand U2803 (N_2803,N_1255,N_1055);
nand U2804 (N_2804,N_1428,N_1534);
xnor U2805 (N_2805,N_1701,N_1828);
and U2806 (N_2806,N_1694,N_1817);
xor U2807 (N_2807,N_1519,N_1323);
nor U2808 (N_2808,N_1217,N_1343);
and U2809 (N_2809,N_1730,N_1929);
nor U2810 (N_2810,N_1445,N_1477);
or U2811 (N_2811,N_1221,N_1315);
and U2812 (N_2812,N_1845,N_1093);
nand U2813 (N_2813,N_1841,N_1636);
or U2814 (N_2814,N_1276,N_1289);
nand U2815 (N_2815,N_1932,N_1720);
nand U2816 (N_2816,N_1095,N_1850);
nand U2817 (N_2817,N_1632,N_1202);
xnor U2818 (N_2818,N_1944,N_1586);
nand U2819 (N_2819,N_1309,N_1074);
or U2820 (N_2820,N_1698,N_1644);
nor U2821 (N_2821,N_1138,N_1396);
xnor U2822 (N_2822,N_1533,N_1277);
nor U2823 (N_2823,N_1120,N_1515);
or U2824 (N_2824,N_1505,N_1955);
or U2825 (N_2825,N_1410,N_1012);
nand U2826 (N_2826,N_1832,N_1740);
xor U2827 (N_2827,N_1197,N_1786);
nand U2828 (N_2828,N_1643,N_1462);
nand U2829 (N_2829,N_1344,N_1986);
nor U2830 (N_2830,N_1569,N_1652);
nor U2831 (N_2831,N_1707,N_1760);
or U2832 (N_2832,N_1474,N_1818);
nor U2833 (N_2833,N_1372,N_1965);
nor U2834 (N_2834,N_1087,N_1868);
nand U2835 (N_2835,N_1900,N_1182);
nor U2836 (N_2836,N_1182,N_1785);
or U2837 (N_2837,N_1303,N_1452);
nand U2838 (N_2838,N_1540,N_1362);
nand U2839 (N_2839,N_1220,N_1838);
nor U2840 (N_2840,N_1794,N_1633);
nand U2841 (N_2841,N_1729,N_1901);
and U2842 (N_2842,N_1944,N_1211);
nand U2843 (N_2843,N_1226,N_1781);
and U2844 (N_2844,N_1654,N_1857);
xor U2845 (N_2845,N_1527,N_1406);
nor U2846 (N_2846,N_1677,N_1634);
nand U2847 (N_2847,N_1717,N_1230);
nor U2848 (N_2848,N_1530,N_1670);
and U2849 (N_2849,N_1030,N_1349);
or U2850 (N_2850,N_1388,N_1196);
nor U2851 (N_2851,N_1837,N_1685);
and U2852 (N_2852,N_1517,N_1676);
nand U2853 (N_2853,N_1168,N_1935);
nor U2854 (N_2854,N_1734,N_1740);
or U2855 (N_2855,N_1708,N_1874);
or U2856 (N_2856,N_1430,N_1163);
nand U2857 (N_2857,N_1998,N_1770);
xnor U2858 (N_2858,N_1397,N_1015);
and U2859 (N_2859,N_1015,N_1848);
nor U2860 (N_2860,N_1345,N_1116);
nor U2861 (N_2861,N_1939,N_1109);
nor U2862 (N_2862,N_1179,N_1163);
nand U2863 (N_2863,N_1260,N_1217);
xnor U2864 (N_2864,N_1399,N_1692);
xnor U2865 (N_2865,N_1563,N_1456);
xor U2866 (N_2866,N_1068,N_1170);
nand U2867 (N_2867,N_1324,N_1013);
or U2868 (N_2868,N_1385,N_1755);
nor U2869 (N_2869,N_1614,N_1399);
and U2870 (N_2870,N_1957,N_1586);
nor U2871 (N_2871,N_1757,N_1139);
nand U2872 (N_2872,N_1891,N_1125);
nand U2873 (N_2873,N_1773,N_1718);
nor U2874 (N_2874,N_1167,N_1454);
nand U2875 (N_2875,N_1040,N_1678);
xor U2876 (N_2876,N_1571,N_1466);
and U2877 (N_2877,N_1677,N_1313);
and U2878 (N_2878,N_1604,N_1510);
nand U2879 (N_2879,N_1990,N_1185);
nor U2880 (N_2880,N_1222,N_1014);
nor U2881 (N_2881,N_1245,N_1685);
xnor U2882 (N_2882,N_1836,N_1711);
xor U2883 (N_2883,N_1971,N_1418);
xnor U2884 (N_2884,N_1537,N_1993);
and U2885 (N_2885,N_1444,N_1119);
nand U2886 (N_2886,N_1732,N_1273);
xnor U2887 (N_2887,N_1798,N_1825);
and U2888 (N_2888,N_1060,N_1353);
nor U2889 (N_2889,N_1394,N_1602);
xor U2890 (N_2890,N_1025,N_1867);
xnor U2891 (N_2891,N_1538,N_1594);
and U2892 (N_2892,N_1911,N_1995);
nor U2893 (N_2893,N_1527,N_1457);
or U2894 (N_2894,N_1044,N_1931);
xor U2895 (N_2895,N_1295,N_1102);
nand U2896 (N_2896,N_1856,N_1731);
or U2897 (N_2897,N_1195,N_1554);
xor U2898 (N_2898,N_1913,N_1857);
xnor U2899 (N_2899,N_1427,N_1024);
or U2900 (N_2900,N_1277,N_1435);
nor U2901 (N_2901,N_1167,N_1686);
nor U2902 (N_2902,N_1601,N_1692);
and U2903 (N_2903,N_1709,N_1697);
nand U2904 (N_2904,N_1713,N_1358);
nand U2905 (N_2905,N_1534,N_1031);
nand U2906 (N_2906,N_1307,N_1915);
nor U2907 (N_2907,N_1276,N_1124);
and U2908 (N_2908,N_1960,N_1600);
nand U2909 (N_2909,N_1367,N_1671);
nor U2910 (N_2910,N_1654,N_1230);
and U2911 (N_2911,N_1193,N_1292);
nand U2912 (N_2912,N_1206,N_1179);
xnor U2913 (N_2913,N_1942,N_1253);
xnor U2914 (N_2914,N_1121,N_1157);
and U2915 (N_2915,N_1411,N_1469);
xnor U2916 (N_2916,N_1659,N_1973);
nand U2917 (N_2917,N_1106,N_1452);
nand U2918 (N_2918,N_1237,N_1338);
nor U2919 (N_2919,N_1704,N_1552);
nor U2920 (N_2920,N_1182,N_1497);
or U2921 (N_2921,N_1013,N_1411);
nand U2922 (N_2922,N_1006,N_1744);
nand U2923 (N_2923,N_1507,N_1007);
nor U2924 (N_2924,N_1772,N_1083);
nor U2925 (N_2925,N_1934,N_1737);
nor U2926 (N_2926,N_1711,N_1623);
or U2927 (N_2927,N_1049,N_1800);
or U2928 (N_2928,N_1280,N_1999);
nand U2929 (N_2929,N_1025,N_1145);
nand U2930 (N_2930,N_1310,N_1196);
or U2931 (N_2931,N_1378,N_1974);
and U2932 (N_2932,N_1188,N_1101);
or U2933 (N_2933,N_1057,N_1333);
xor U2934 (N_2934,N_1814,N_1382);
nand U2935 (N_2935,N_1144,N_1184);
xnor U2936 (N_2936,N_1525,N_1030);
nor U2937 (N_2937,N_1779,N_1943);
nand U2938 (N_2938,N_1942,N_1773);
nand U2939 (N_2939,N_1170,N_1981);
xnor U2940 (N_2940,N_1414,N_1200);
or U2941 (N_2941,N_1905,N_1884);
nor U2942 (N_2942,N_1351,N_1226);
and U2943 (N_2943,N_1459,N_1578);
and U2944 (N_2944,N_1743,N_1776);
nor U2945 (N_2945,N_1605,N_1389);
and U2946 (N_2946,N_1951,N_1572);
nor U2947 (N_2947,N_1125,N_1632);
nor U2948 (N_2948,N_1757,N_1610);
and U2949 (N_2949,N_1582,N_1007);
nor U2950 (N_2950,N_1669,N_1195);
or U2951 (N_2951,N_1759,N_1871);
nand U2952 (N_2952,N_1439,N_1901);
and U2953 (N_2953,N_1079,N_1001);
xnor U2954 (N_2954,N_1214,N_1311);
or U2955 (N_2955,N_1994,N_1597);
nor U2956 (N_2956,N_1930,N_1543);
nor U2957 (N_2957,N_1602,N_1988);
and U2958 (N_2958,N_1337,N_1646);
and U2959 (N_2959,N_1914,N_1804);
xnor U2960 (N_2960,N_1672,N_1559);
and U2961 (N_2961,N_1685,N_1679);
nand U2962 (N_2962,N_1097,N_1000);
xor U2963 (N_2963,N_1229,N_1624);
nand U2964 (N_2964,N_1478,N_1436);
or U2965 (N_2965,N_1449,N_1477);
nand U2966 (N_2966,N_1560,N_1702);
nor U2967 (N_2967,N_1698,N_1402);
nand U2968 (N_2968,N_1918,N_1635);
nor U2969 (N_2969,N_1582,N_1111);
nor U2970 (N_2970,N_1188,N_1121);
nor U2971 (N_2971,N_1196,N_1108);
nand U2972 (N_2972,N_1589,N_1052);
or U2973 (N_2973,N_1499,N_1635);
or U2974 (N_2974,N_1712,N_1821);
and U2975 (N_2975,N_1470,N_1528);
nand U2976 (N_2976,N_1104,N_1236);
xnor U2977 (N_2977,N_1866,N_1820);
and U2978 (N_2978,N_1186,N_1124);
xnor U2979 (N_2979,N_1684,N_1457);
nand U2980 (N_2980,N_1009,N_1356);
nand U2981 (N_2981,N_1631,N_1330);
or U2982 (N_2982,N_1822,N_1174);
xnor U2983 (N_2983,N_1203,N_1653);
nor U2984 (N_2984,N_1475,N_1419);
or U2985 (N_2985,N_1878,N_1579);
and U2986 (N_2986,N_1271,N_1556);
nand U2987 (N_2987,N_1964,N_1064);
nor U2988 (N_2988,N_1182,N_1879);
or U2989 (N_2989,N_1714,N_1938);
nand U2990 (N_2990,N_1979,N_1490);
or U2991 (N_2991,N_1564,N_1935);
xor U2992 (N_2992,N_1109,N_1458);
or U2993 (N_2993,N_1239,N_1448);
nand U2994 (N_2994,N_1838,N_1443);
and U2995 (N_2995,N_1696,N_1353);
nor U2996 (N_2996,N_1275,N_1258);
and U2997 (N_2997,N_1338,N_1875);
nor U2998 (N_2998,N_1381,N_1890);
nand U2999 (N_2999,N_1301,N_1351);
nand U3000 (N_3000,N_2017,N_2158);
and U3001 (N_3001,N_2789,N_2474);
nor U3002 (N_3002,N_2283,N_2078);
xor U3003 (N_3003,N_2256,N_2972);
xnor U3004 (N_3004,N_2291,N_2621);
nor U3005 (N_3005,N_2172,N_2811);
nand U3006 (N_3006,N_2243,N_2346);
xor U3007 (N_3007,N_2877,N_2505);
and U3008 (N_3008,N_2897,N_2774);
nand U3009 (N_3009,N_2241,N_2166);
xnor U3010 (N_3010,N_2205,N_2514);
and U3011 (N_3011,N_2362,N_2295);
nand U3012 (N_3012,N_2983,N_2962);
xnor U3013 (N_3013,N_2784,N_2091);
nor U3014 (N_3014,N_2325,N_2936);
nand U3015 (N_3015,N_2513,N_2799);
xnor U3016 (N_3016,N_2351,N_2976);
and U3017 (N_3017,N_2143,N_2824);
or U3018 (N_3018,N_2562,N_2528);
and U3019 (N_3019,N_2544,N_2566);
nand U3020 (N_3020,N_2451,N_2218);
or U3021 (N_3021,N_2735,N_2367);
or U3022 (N_3022,N_2581,N_2492);
nand U3023 (N_3023,N_2081,N_2374);
xnor U3024 (N_3024,N_2751,N_2048);
nor U3025 (N_3025,N_2371,N_2058);
xnor U3026 (N_3026,N_2155,N_2418);
xnor U3027 (N_3027,N_2586,N_2392);
nor U3028 (N_3028,N_2190,N_2613);
nand U3029 (N_3029,N_2405,N_2272);
or U3030 (N_3030,N_2075,N_2627);
nand U3031 (N_3031,N_2736,N_2404);
or U3032 (N_3032,N_2583,N_2742);
nor U3033 (N_3033,N_2519,N_2746);
and U3034 (N_3034,N_2323,N_2432);
xnor U3035 (N_3035,N_2044,N_2846);
and U3036 (N_3036,N_2138,N_2309);
nor U3037 (N_3037,N_2576,N_2658);
nand U3038 (N_3038,N_2959,N_2357);
nor U3039 (N_3039,N_2217,N_2607);
nand U3040 (N_3040,N_2132,N_2164);
nor U3041 (N_3041,N_2473,N_2468);
nor U3042 (N_3042,N_2297,N_2956);
xor U3043 (N_3043,N_2677,N_2083);
xor U3044 (N_3044,N_2591,N_2171);
nor U3045 (N_3045,N_2604,N_2881);
or U3046 (N_3046,N_2597,N_2643);
xor U3047 (N_3047,N_2728,N_2457);
nor U3048 (N_3048,N_2935,N_2781);
and U3049 (N_3049,N_2648,N_2993);
or U3050 (N_3050,N_2424,N_2675);
nand U3051 (N_3051,N_2395,N_2332);
and U3052 (N_3052,N_2630,N_2699);
and U3053 (N_3053,N_2294,N_2813);
xor U3054 (N_3054,N_2684,N_2456);
or U3055 (N_3055,N_2957,N_2884);
or U3056 (N_3056,N_2944,N_2831);
or U3057 (N_3057,N_2082,N_2796);
nand U3058 (N_3058,N_2015,N_2169);
nand U3059 (N_3059,N_2614,N_2146);
nor U3060 (N_3060,N_2270,N_2790);
xnor U3061 (N_3061,N_2531,N_2317);
nand U3062 (N_3062,N_2449,N_2486);
or U3063 (N_3063,N_2483,N_2919);
and U3064 (N_3064,N_2096,N_2599);
nor U3065 (N_3065,N_2454,N_2899);
and U3066 (N_3066,N_2380,N_2500);
nor U3067 (N_3067,N_2706,N_2147);
nand U3068 (N_3068,N_2996,N_2927);
xnor U3069 (N_3069,N_2772,N_2408);
and U3070 (N_3070,N_2720,N_2240);
or U3071 (N_3071,N_2211,N_2467);
xor U3072 (N_3072,N_2333,N_2741);
or U3073 (N_3073,N_2749,N_2200);
nor U3074 (N_3074,N_2010,N_2232);
or U3075 (N_3075,N_2763,N_2637);
nor U3076 (N_3076,N_2274,N_2777);
or U3077 (N_3077,N_2046,N_2038);
or U3078 (N_3078,N_2924,N_2238);
nor U3079 (N_3079,N_2978,N_2108);
nor U3080 (N_3080,N_2871,N_2328);
xor U3081 (N_3081,N_2131,N_2106);
or U3082 (N_3082,N_2445,N_2506);
nor U3083 (N_3083,N_2565,N_2902);
xor U3084 (N_3084,N_2140,N_2365);
nand U3085 (N_3085,N_2582,N_2753);
and U3086 (N_3086,N_2293,N_2242);
nand U3087 (N_3087,N_2888,N_2536);
or U3088 (N_3088,N_2117,N_2610);
nor U3089 (N_3089,N_2791,N_2471);
nand U3090 (N_3090,N_2119,N_2450);
nand U3091 (N_3091,N_2943,N_2435);
xnor U3092 (N_3092,N_2692,N_2055);
nor U3093 (N_3093,N_2480,N_2535);
nand U3094 (N_3094,N_2191,N_2255);
and U3095 (N_3095,N_2700,N_2246);
nand U3096 (N_3096,N_2768,N_2532);
and U3097 (N_3097,N_2413,N_2624);
nor U3098 (N_3098,N_2496,N_2429);
xor U3099 (N_3099,N_2723,N_2157);
xor U3100 (N_3100,N_2859,N_2909);
or U3101 (N_3101,N_2981,N_2002);
and U3102 (N_3102,N_2175,N_2820);
and U3103 (N_3103,N_2515,N_2690);
nand U3104 (N_3104,N_2012,N_2727);
xor U3105 (N_3105,N_2953,N_2161);
nor U3106 (N_3106,N_2227,N_2244);
nand U3107 (N_3107,N_2137,N_2679);
nor U3108 (N_3108,N_2236,N_2288);
and U3109 (N_3109,N_2014,N_2072);
nor U3110 (N_3110,N_2299,N_2748);
xnor U3111 (N_3111,N_2027,N_2592);
nand U3112 (N_3112,N_2366,N_2856);
xnor U3113 (N_3113,N_2925,N_2298);
and U3114 (N_3114,N_2198,N_2854);
xnor U3115 (N_3115,N_2262,N_2818);
and U3116 (N_3116,N_2303,N_2016);
nor U3117 (N_3117,N_2650,N_2965);
or U3118 (N_3118,N_2215,N_2938);
nand U3119 (N_3119,N_2070,N_2431);
nor U3120 (N_3120,N_2714,N_2989);
xnor U3121 (N_3121,N_2484,N_2141);
and U3122 (N_3122,N_2076,N_2825);
nor U3123 (N_3123,N_2969,N_2701);
or U3124 (N_3124,N_2250,N_2833);
nand U3125 (N_3125,N_2278,N_2767);
or U3126 (N_3126,N_2605,N_2857);
nand U3127 (N_3127,N_2159,N_2381);
and U3128 (N_3128,N_2873,N_2747);
and U3129 (N_3129,N_2419,N_2202);
nand U3130 (N_3130,N_2406,N_2640);
nand U3131 (N_3131,N_2391,N_2337);
nand U3132 (N_3132,N_2370,N_2415);
xor U3133 (N_3133,N_2363,N_2906);
xnor U3134 (N_3134,N_2301,N_2901);
and U3135 (N_3135,N_2130,N_2841);
nand U3136 (N_3136,N_2339,N_2921);
or U3137 (N_3137,N_2320,N_2039);
nand U3138 (N_3138,N_2470,N_2252);
nand U3139 (N_3139,N_2573,N_2187);
xor U3140 (N_3140,N_2882,N_2422);
xor U3141 (N_3141,N_2101,N_2305);
xor U3142 (N_3142,N_2529,N_2281);
nor U3143 (N_3143,N_2122,N_2360);
nand U3144 (N_3144,N_2894,N_2525);
nor U3145 (N_3145,N_2696,N_2606);
and U3146 (N_3146,N_2596,N_2071);
nor U3147 (N_3147,N_2974,N_2446);
and U3148 (N_3148,N_2510,N_2030);
nand U3149 (N_3149,N_2788,N_2886);
nor U3150 (N_3150,N_2835,N_2089);
nor U3151 (N_3151,N_2144,N_2114);
xor U3152 (N_3152,N_2920,N_2847);
nor U3153 (N_3153,N_2633,N_2853);
nand U3154 (N_3154,N_2267,N_2389);
xnor U3155 (N_3155,N_2612,N_2782);
nor U3156 (N_3156,N_2843,N_2798);
nor U3157 (N_3157,N_2534,N_2265);
and U3158 (N_3158,N_2695,N_2386);
or U3159 (N_3159,N_2029,N_2353);
nand U3160 (N_3160,N_2379,N_2358);
xor U3161 (N_3161,N_2290,N_2522);
and U3162 (N_3162,N_2973,N_2098);
xor U3163 (N_3163,N_2276,N_2656);
nand U3164 (N_3164,N_2382,N_2300);
nor U3165 (N_3165,N_2099,N_2923);
or U3166 (N_3166,N_2125,N_2182);
or U3167 (N_3167,N_2403,N_2285);
or U3168 (N_3168,N_2917,N_2307);
nand U3169 (N_3169,N_2863,N_2639);
nor U3170 (N_3170,N_2231,N_2491);
and U3171 (N_3171,N_2100,N_2185);
xnor U3172 (N_3172,N_2546,N_2762);
nor U3173 (N_3173,N_2213,N_2848);
and U3174 (N_3174,N_2930,N_2134);
nand U3175 (N_3175,N_2795,N_2711);
nor U3176 (N_3176,N_2121,N_2839);
nand U3177 (N_3177,N_2942,N_2201);
or U3178 (N_3178,N_2088,N_2752);
and U3179 (N_3179,N_2123,N_2387);
xor U3180 (N_3180,N_2277,N_2951);
or U3181 (N_3181,N_2941,N_2771);
nand U3182 (N_3182,N_2349,N_2964);
nor U3183 (N_3183,N_2129,N_2673);
nand U3184 (N_3184,N_2954,N_2181);
and U3185 (N_3185,N_2685,N_2563);
and U3186 (N_3186,N_2952,N_2322);
xor U3187 (N_3187,N_2672,N_2958);
and U3188 (N_3188,N_2571,N_2442);
and U3189 (N_3189,N_2011,N_2263);
and U3190 (N_3190,N_2682,N_2775);
nand U3191 (N_3191,N_2968,N_2885);
or U3192 (N_3192,N_2092,N_2054);
and U3193 (N_3193,N_2557,N_2876);
nand U3194 (N_3194,N_2223,N_2439);
nor U3195 (N_3195,N_2516,N_2050);
or U3196 (N_3196,N_2127,N_2802);
xor U3197 (N_3197,N_2584,N_2426);
or U3198 (N_3198,N_2869,N_2926);
nor U3199 (N_3199,N_2047,N_2004);
or U3200 (N_3200,N_2345,N_2049);
xnor U3201 (N_3201,N_2173,N_2678);
and U3202 (N_3202,N_2312,N_2718);
nor U3203 (N_3203,N_2864,N_2352);
nor U3204 (N_3204,N_2485,N_2179);
nor U3205 (N_3205,N_2036,N_2879);
and U3206 (N_3206,N_2521,N_2651);
nand U3207 (N_3207,N_2489,N_2397);
nor U3208 (N_3208,N_2388,N_2556);
or U3209 (N_3209,N_2618,N_2588);
xor U3210 (N_3210,N_2154,N_2355);
xor U3211 (N_3211,N_2458,N_2955);
and U3212 (N_3212,N_2033,N_2253);
xor U3213 (N_3213,N_2296,N_2553);
nor U3214 (N_3214,N_2487,N_2688);
nor U3215 (N_3215,N_2103,N_2980);
nor U3216 (N_3216,N_2399,N_2574);
and U3217 (N_3217,N_2773,N_2693);
nor U3218 (N_3218,N_2647,N_2903);
xor U3219 (N_3219,N_2000,N_2235);
xor U3220 (N_3220,N_2937,N_2502);
nor U3221 (N_3221,N_2570,N_2664);
xor U3222 (N_3222,N_2990,N_2947);
nor U3223 (N_3223,N_2611,N_2786);
nand U3224 (N_3224,N_2335,N_2945);
nand U3225 (N_3225,N_2713,N_2644);
nor U3226 (N_3226,N_2828,N_2249);
and U3227 (N_3227,N_2933,N_2616);
xnor U3228 (N_3228,N_2396,N_2538);
xnor U3229 (N_3229,N_2868,N_2511);
and U3230 (N_3230,N_2292,N_2977);
and U3231 (N_3231,N_2006,N_2949);
or U3232 (N_3232,N_2875,N_2725);
nor U3233 (N_3233,N_2372,N_2118);
nand U3234 (N_3234,N_2549,N_2020);
or U3235 (N_3235,N_2539,N_2453);
and U3236 (N_3236,N_2409,N_2602);
nand U3237 (N_3237,N_2259,N_2922);
and U3238 (N_3238,N_2412,N_2109);
or U3239 (N_3239,N_2940,N_2260);
xnor U3240 (N_3240,N_2589,N_2629);
or U3241 (N_3241,N_2934,N_2475);
and U3242 (N_3242,N_2851,N_2237);
or U3243 (N_3243,N_2459,N_2587);
xnor U3244 (N_3244,N_2914,N_2226);
nand U3245 (N_3245,N_2832,N_2359);
or U3246 (N_3246,N_2855,N_2434);
nand U3247 (N_3247,N_2208,N_2575);
nand U3248 (N_3248,N_2135,N_2615);
or U3249 (N_3249,N_2193,N_2660);
nand U3250 (N_3250,N_2269,N_2273);
nor U3251 (N_3251,N_2452,N_2268);
xnor U3252 (N_3252,N_2170,N_2719);
xnor U3253 (N_3253,N_2984,N_2601);
or U3254 (N_3254,N_2074,N_2815);
nor U3255 (N_3255,N_2862,N_2148);
xnor U3256 (N_3256,N_2776,N_2662);
xor U3257 (N_3257,N_2209,N_2478);
xnor U3258 (N_3258,N_2517,N_2378);
xor U3259 (N_3259,N_2160,N_2433);
nand U3260 (N_3260,N_2731,N_2804);
nor U3261 (N_3261,N_2373,N_2056);
or U3262 (N_3262,N_2932,N_2961);
and U3263 (N_3263,N_2622,N_2686);
and U3264 (N_3264,N_2849,N_2830);
or U3265 (N_3265,N_2220,N_2992);
or U3266 (N_3266,N_2997,N_2737);
nor U3267 (N_3267,N_2994,N_2558);
and U3268 (N_3268,N_2115,N_2493);
or U3269 (N_3269,N_2344,N_2668);
xor U3270 (N_3270,N_2655,N_2377);
nor U3271 (N_3271,N_2887,N_2834);
nor U3272 (N_3272,N_2013,N_2598);
xor U3273 (N_3273,N_2628,N_2537);
nand U3274 (N_3274,N_2745,N_2913);
nand U3275 (N_3275,N_2548,N_2022);
or U3276 (N_3276,N_2916,N_2061);
nor U3277 (N_3277,N_2635,N_2165);
xnor U3278 (N_3278,N_2090,N_2991);
xor U3279 (N_3279,N_2948,N_2311);
and U3280 (N_3280,N_2509,N_2266);
or U3281 (N_3281,N_2340,N_2638);
xnor U3282 (N_3282,N_2860,N_2168);
xnor U3283 (N_3283,N_2645,N_2809);
nor U3284 (N_3284,N_2331,N_2721);
nand U3285 (N_3285,N_2021,N_2659);
nor U3286 (N_3286,N_2946,N_2874);
xnor U3287 (N_3287,N_2095,N_2836);
nand U3288 (N_3288,N_2214,N_2866);
nor U3289 (N_3289,N_2180,N_2005);
xnor U3290 (N_3290,N_2907,N_2754);
or U3291 (N_3291,N_2222,N_2670);
xnor U3292 (N_3292,N_2136,N_2219);
xnor U3293 (N_3293,N_2540,N_2816);
or U3294 (N_3294,N_2073,N_2407);
or U3295 (N_3295,N_2654,N_2110);
or U3296 (N_3296,N_2585,N_2765);
and U3297 (N_3297,N_2079,N_2826);
xnor U3298 (N_3298,N_2019,N_2199);
and U3299 (N_3299,N_2858,N_2086);
nor U3300 (N_3300,N_2619,N_2979);
xnor U3301 (N_3301,N_2769,N_2623);
nor U3302 (N_3302,N_2465,N_2560);
or U3303 (N_3303,N_2709,N_2669);
and U3304 (N_3304,N_2987,N_2810);
nor U3305 (N_3305,N_2982,N_2448);
nand U3306 (N_3306,N_2803,N_2840);
or U3307 (N_3307,N_2649,N_2402);
nor U3308 (N_3308,N_2900,N_2488);
xor U3309 (N_3309,N_2463,N_2003);
xnor U3310 (N_3310,N_2376,N_2400);
nand U3311 (N_3311,N_2069,N_2113);
nand U3312 (N_3312,N_2104,N_2183);
xor U3313 (N_3313,N_2212,N_2194);
xor U3314 (N_3314,N_2271,N_2744);
xnor U3315 (N_3315,N_2318,N_2228);
nand U3316 (N_3316,N_2898,N_2393);
nand U3317 (N_3317,N_2334,N_2304);
nand U3318 (N_3318,N_2554,N_2494);
or U3319 (N_3319,N_2908,N_2652);
nor U3320 (N_3320,N_2653,N_2436);
or U3321 (N_3321,N_2893,N_2827);
xnor U3322 (N_3322,N_2755,N_2733);
and U3323 (N_3323,N_2889,N_2438);
or U3324 (N_3324,N_2085,N_2306);
or U3325 (N_3325,N_2911,N_2821);
nand U3326 (N_3326,N_2822,N_2001);
xnor U3327 (N_3327,N_2657,N_2369);
nor U3328 (N_3328,N_2462,N_2233);
xnor U3329 (N_3329,N_2896,N_2910);
and U3330 (N_3330,N_2757,N_2490);
nor U3331 (N_3331,N_2829,N_2915);
and U3332 (N_3332,N_2440,N_2375);
and U3333 (N_3333,N_2551,N_2031);
nand U3334 (N_3334,N_2676,N_2350);
nand U3335 (N_3335,N_2750,N_2112);
nor U3336 (N_3336,N_2356,N_2385);
nand U3337 (N_3337,N_2321,N_2609);
and U3338 (N_3338,N_2145,N_2230);
xnor U3339 (N_3339,N_2729,N_2430);
and U3340 (N_3340,N_2280,N_2087);
and U3341 (N_3341,N_2097,N_2043);
nand U3342 (N_3342,N_2793,N_2975);
nand U3343 (N_3343,N_2880,N_2697);
and U3344 (N_3344,N_2845,N_2667);
nor U3345 (N_3345,N_2567,N_2064);
xnor U3346 (N_3346,N_2569,N_2111);
nand U3347 (N_3347,N_2342,N_2248);
nand U3348 (N_3348,N_2778,N_2279);
xor U3349 (N_3349,N_2258,N_2878);
nor U3350 (N_3350,N_2626,N_2730);
or U3351 (N_3351,N_2518,N_2308);
nor U3352 (N_3352,N_2636,N_2469);
or U3353 (N_3353,N_2336,N_2466);
xnor U3354 (N_3354,N_2162,N_2053);
nor U3355 (N_3355,N_2823,N_2892);
nand U3356 (N_3356,N_2417,N_2837);
and U3357 (N_3357,N_2302,N_2051);
nor U3358 (N_3358,N_2124,N_2133);
xor U3359 (N_3359,N_2313,N_2726);
nand U3360 (N_3360,N_2008,N_2527);
nor U3361 (N_3361,N_2310,N_2414);
xnor U3362 (N_3362,N_2533,N_2608);
nor U3363 (N_3363,N_2530,N_2666);
and U3364 (N_3364,N_2542,N_2423);
nor U3365 (N_3365,N_2819,N_2128);
nor U3366 (N_3366,N_2779,N_2284);
nand U3367 (N_3367,N_2674,N_2764);
and U3368 (N_3368,N_2971,N_2229);
or U3369 (N_3369,N_2364,N_2787);
and U3370 (N_3370,N_2756,N_2671);
nand U3371 (N_3371,N_2870,N_2093);
or U3372 (N_3372,N_2383,N_2526);
xor U3373 (N_3373,N_2476,N_2151);
nand U3374 (N_3374,N_2724,N_2698);
or U3375 (N_3375,N_2929,N_2443);
or U3376 (N_3376,N_2009,N_2420);
nand U3377 (N_3377,N_2632,N_2501);
nor U3378 (N_3378,N_2206,N_2499);
xor U3379 (N_3379,N_2722,N_2316);
xor U3380 (N_3380,N_2028,N_2066);
and U3381 (N_3381,N_2464,N_2572);
nor U3382 (N_3382,N_2807,N_2065);
and U3383 (N_3383,N_2761,N_2985);
nor U3384 (N_3384,N_2261,N_2805);
xnor U3385 (N_3385,N_2504,N_2150);
or U3386 (N_3386,N_2460,N_2703);
nand U3387 (N_3387,N_2107,N_2617);
or U3388 (N_3388,N_2394,N_2286);
nor U3389 (N_3389,N_2681,N_2153);
nor U3390 (N_3390,N_2247,N_2197);
or U3391 (N_3391,N_2928,N_2023);
or U3392 (N_3392,N_2067,N_2105);
and U3393 (N_3393,N_2743,N_2264);
or U3394 (N_3394,N_2760,N_2411);
nor U3395 (N_3395,N_2792,N_2931);
or U3396 (N_3396,N_2497,N_2225);
or U3397 (N_3397,N_2060,N_2080);
xor U3398 (N_3398,N_2057,N_2207);
nand U3399 (N_3399,N_2361,N_2203);
nand U3400 (N_3400,N_2814,N_2094);
and U3401 (N_3401,N_2343,N_2441);
nor U3402 (N_3402,N_2641,N_2806);
nand U3403 (N_3403,N_2196,N_2883);
xor U3404 (N_3404,N_2390,N_2084);
or U3405 (N_3405,N_2221,N_2998);
nand U3406 (N_3406,N_2801,N_2715);
nand U3407 (N_3407,N_2872,N_2708);
or U3408 (N_3408,N_2867,N_2642);
xnor U3409 (N_3409,N_2579,N_2177);
nand U3410 (N_3410,N_2024,N_2188);
nand U3411 (N_3411,N_2368,N_2694);
nand U3412 (N_3412,N_2710,N_2447);
and U3413 (N_3413,N_2738,N_2543);
xnor U3414 (N_3414,N_2865,N_2507);
nor U3415 (N_3415,N_2239,N_2995);
xor U3416 (N_3416,N_2766,N_2319);
or U3417 (N_3417,N_2603,N_2797);
or U3418 (N_3418,N_2590,N_2018);
xor U3419 (N_3419,N_2139,N_2716);
and U3420 (N_3420,N_2508,N_2498);
nor U3421 (N_3421,N_2564,N_2425);
nor U3422 (N_3422,N_2999,N_2663);
and U3423 (N_3423,N_2102,N_2477);
nand U3424 (N_3424,N_2665,N_2547);
nor U3425 (N_3425,N_2245,N_2552);
nand U3426 (N_3426,N_2966,N_2705);
xor U3427 (N_3427,N_2912,N_2347);
nor U3428 (N_3428,N_2568,N_2338);
nor U3429 (N_3429,N_2905,N_2689);
nand U3430 (N_3430,N_2950,N_2026);
xnor U3431 (N_3431,N_2812,N_2437);
nor U3432 (N_3432,N_2739,N_2416);
xor U3433 (N_3433,N_2986,N_2068);
nor U3434 (N_3434,N_2427,N_2126);
or U3435 (N_3435,N_2348,N_2282);
nor U3436 (N_3436,N_2204,N_2580);
or U3437 (N_3437,N_2025,N_2503);
or U3438 (N_3438,N_2890,N_2620);
xnor U3439 (N_3439,N_2341,N_2780);
or U3440 (N_3440,N_2520,N_2523);
nand U3441 (N_3441,N_2192,N_2461);
nand U3442 (N_3442,N_2354,N_2324);
xor U3443 (N_3443,N_2315,N_2210);
nand U3444 (N_3444,N_2257,N_2455);
or U3445 (N_3445,N_2891,N_2495);
and U3446 (N_3446,N_2142,N_2559);
nor U3447 (N_3447,N_2593,N_2524);
xor U3448 (N_3448,N_2398,N_2691);
nand U3449 (N_3449,N_2037,N_2289);
xor U3450 (N_3450,N_2702,N_2555);
or U3451 (N_3451,N_2687,N_2042);
or U3452 (N_3452,N_2712,N_2216);
nor U3453 (N_3453,N_2861,N_2770);
nand U3454 (N_3454,N_2704,N_2330);
nand U3455 (N_3455,N_2040,N_2149);
or U3456 (N_3456,N_2167,N_2410);
xnor U3457 (N_3457,N_2163,N_2577);
and U3458 (N_3458,N_2421,N_2287);
and U3459 (N_3459,N_2428,N_2631);
and U3460 (N_3460,N_2512,N_2254);
and U3461 (N_3461,N_2541,N_2401);
and U3462 (N_3462,N_2251,N_2561);
nand U3463 (N_3463,N_2850,N_2838);
and U3464 (N_3464,N_2680,N_2052);
or U3465 (N_3465,N_2184,N_2967);
nor U3466 (N_3466,N_2234,N_2740);
and U3467 (N_3467,N_2479,N_2482);
nor U3468 (N_3468,N_2963,N_2960);
or U3469 (N_3469,N_2895,N_2007);
or U3470 (N_3470,N_2035,N_2472);
nand U3471 (N_3471,N_2594,N_2174);
and U3472 (N_3472,N_2595,N_2918);
nand U3473 (N_3473,N_2329,N_2578);
nor U3474 (N_3474,N_2314,N_2178);
or U3475 (N_3475,N_2032,N_2550);
nand U3476 (N_3476,N_2970,N_2077);
and U3477 (N_3477,N_2844,N_2817);
xor U3478 (N_3478,N_2732,N_2634);
or U3479 (N_3479,N_2852,N_2327);
nor U3480 (N_3480,N_2224,N_2116);
xnor U3481 (N_3481,N_2758,N_2904);
or U3482 (N_3482,N_2800,N_2734);
xnor U3483 (N_3483,N_2384,N_2600);
nand U3484 (N_3484,N_2063,N_2794);
or U3485 (N_3485,N_2045,N_2156);
nor U3486 (N_3486,N_2481,N_2759);
and U3487 (N_3487,N_2275,N_2444);
nand U3488 (N_3488,N_2988,N_2059);
nand U3489 (N_3489,N_2062,N_2189);
xnor U3490 (N_3490,N_2176,N_2545);
nor U3491 (N_3491,N_2683,N_2646);
nand U3492 (N_3492,N_2842,N_2939);
and U3493 (N_3493,N_2195,N_2120);
nand U3494 (N_3494,N_2707,N_2041);
xnor U3495 (N_3495,N_2625,N_2186);
nand U3496 (N_3496,N_2034,N_2326);
or U3497 (N_3497,N_2808,N_2785);
nor U3498 (N_3498,N_2783,N_2152);
or U3499 (N_3499,N_2717,N_2661);
nand U3500 (N_3500,N_2033,N_2297);
or U3501 (N_3501,N_2385,N_2049);
or U3502 (N_3502,N_2233,N_2348);
nor U3503 (N_3503,N_2956,N_2520);
or U3504 (N_3504,N_2583,N_2832);
and U3505 (N_3505,N_2437,N_2974);
nand U3506 (N_3506,N_2535,N_2277);
or U3507 (N_3507,N_2151,N_2588);
and U3508 (N_3508,N_2776,N_2426);
and U3509 (N_3509,N_2137,N_2783);
or U3510 (N_3510,N_2782,N_2854);
nor U3511 (N_3511,N_2379,N_2977);
nor U3512 (N_3512,N_2016,N_2216);
xnor U3513 (N_3513,N_2538,N_2760);
and U3514 (N_3514,N_2525,N_2984);
nand U3515 (N_3515,N_2538,N_2394);
xor U3516 (N_3516,N_2333,N_2051);
or U3517 (N_3517,N_2395,N_2721);
nand U3518 (N_3518,N_2153,N_2320);
nor U3519 (N_3519,N_2290,N_2125);
nand U3520 (N_3520,N_2705,N_2985);
or U3521 (N_3521,N_2416,N_2058);
and U3522 (N_3522,N_2935,N_2062);
xor U3523 (N_3523,N_2299,N_2612);
or U3524 (N_3524,N_2988,N_2807);
or U3525 (N_3525,N_2603,N_2620);
nand U3526 (N_3526,N_2615,N_2864);
and U3527 (N_3527,N_2400,N_2568);
and U3528 (N_3528,N_2908,N_2208);
or U3529 (N_3529,N_2510,N_2133);
nor U3530 (N_3530,N_2518,N_2053);
or U3531 (N_3531,N_2201,N_2986);
nand U3532 (N_3532,N_2254,N_2258);
and U3533 (N_3533,N_2689,N_2319);
nand U3534 (N_3534,N_2401,N_2678);
nand U3535 (N_3535,N_2193,N_2109);
nor U3536 (N_3536,N_2121,N_2865);
and U3537 (N_3537,N_2975,N_2214);
nor U3538 (N_3538,N_2478,N_2838);
and U3539 (N_3539,N_2247,N_2577);
and U3540 (N_3540,N_2194,N_2044);
nor U3541 (N_3541,N_2562,N_2617);
nor U3542 (N_3542,N_2577,N_2338);
nor U3543 (N_3543,N_2187,N_2944);
and U3544 (N_3544,N_2096,N_2683);
nand U3545 (N_3545,N_2081,N_2444);
nand U3546 (N_3546,N_2149,N_2212);
nor U3547 (N_3547,N_2616,N_2538);
nor U3548 (N_3548,N_2588,N_2911);
nor U3549 (N_3549,N_2875,N_2661);
xor U3550 (N_3550,N_2464,N_2167);
nand U3551 (N_3551,N_2656,N_2788);
nor U3552 (N_3552,N_2789,N_2775);
nand U3553 (N_3553,N_2865,N_2593);
xor U3554 (N_3554,N_2883,N_2110);
and U3555 (N_3555,N_2963,N_2783);
and U3556 (N_3556,N_2385,N_2380);
xor U3557 (N_3557,N_2569,N_2291);
xor U3558 (N_3558,N_2519,N_2220);
nor U3559 (N_3559,N_2767,N_2381);
nand U3560 (N_3560,N_2994,N_2778);
nand U3561 (N_3561,N_2998,N_2014);
or U3562 (N_3562,N_2180,N_2332);
nand U3563 (N_3563,N_2520,N_2071);
xnor U3564 (N_3564,N_2854,N_2377);
or U3565 (N_3565,N_2732,N_2666);
or U3566 (N_3566,N_2335,N_2341);
or U3567 (N_3567,N_2337,N_2953);
or U3568 (N_3568,N_2701,N_2779);
xor U3569 (N_3569,N_2062,N_2043);
nor U3570 (N_3570,N_2637,N_2388);
nand U3571 (N_3571,N_2239,N_2445);
or U3572 (N_3572,N_2202,N_2582);
nand U3573 (N_3573,N_2099,N_2909);
xor U3574 (N_3574,N_2169,N_2768);
and U3575 (N_3575,N_2284,N_2920);
nand U3576 (N_3576,N_2392,N_2979);
xnor U3577 (N_3577,N_2939,N_2751);
xor U3578 (N_3578,N_2607,N_2991);
or U3579 (N_3579,N_2202,N_2132);
nand U3580 (N_3580,N_2730,N_2171);
xnor U3581 (N_3581,N_2233,N_2766);
nor U3582 (N_3582,N_2699,N_2358);
nor U3583 (N_3583,N_2105,N_2435);
or U3584 (N_3584,N_2816,N_2141);
nor U3585 (N_3585,N_2417,N_2154);
nand U3586 (N_3586,N_2800,N_2284);
nand U3587 (N_3587,N_2217,N_2191);
xor U3588 (N_3588,N_2244,N_2743);
or U3589 (N_3589,N_2034,N_2111);
nand U3590 (N_3590,N_2943,N_2854);
xnor U3591 (N_3591,N_2505,N_2181);
nor U3592 (N_3592,N_2141,N_2154);
nand U3593 (N_3593,N_2827,N_2708);
nor U3594 (N_3594,N_2812,N_2867);
and U3595 (N_3595,N_2784,N_2001);
and U3596 (N_3596,N_2401,N_2584);
or U3597 (N_3597,N_2114,N_2619);
or U3598 (N_3598,N_2687,N_2459);
xnor U3599 (N_3599,N_2504,N_2512);
nand U3600 (N_3600,N_2070,N_2958);
and U3601 (N_3601,N_2315,N_2340);
and U3602 (N_3602,N_2538,N_2236);
nand U3603 (N_3603,N_2444,N_2493);
or U3604 (N_3604,N_2884,N_2363);
or U3605 (N_3605,N_2528,N_2995);
nor U3606 (N_3606,N_2388,N_2907);
and U3607 (N_3607,N_2135,N_2981);
nand U3608 (N_3608,N_2826,N_2104);
or U3609 (N_3609,N_2079,N_2141);
or U3610 (N_3610,N_2075,N_2887);
nand U3611 (N_3611,N_2534,N_2040);
xor U3612 (N_3612,N_2546,N_2433);
nand U3613 (N_3613,N_2795,N_2760);
nand U3614 (N_3614,N_2878,N_2526);
nor U3615 (N_3615,N_2056,N_2290);
or U3616 (N_3616,N_2251,N_2621);
nor U3617 (N_3617,N_2059,N_2983);
nand U3618 (N_3618,N_2179,N_2415);
nor U3619 (N_3619,N_2097,N_2477);
nand U3620 (N_3620,N_2844,N_2895);
xor U3621 (N_3621,N_2109,N_2925);
and U3622 (N_3622,N_2089,N_2543);
xnor U3623 (N_3623,N_2931,N_2275);
nor U3624 (N_3624,N_2523,N_2251);
and U3625 (N_3625,N_2746,N_2664);
nor U3626 (N_3626,N_2472,N_2836);
nand U3627 (N_3627,N_2653,N_2416);
nor U3628 (N_3628,N_2215,N_2404);
or U3629 (N_3629,N_2816,N_2562);
and U3630 (N_3630,N_2712,N_2084);
nor U3631 (N_3631,N_2711,N_2886);
nor U3632 (N_3632,N_2588,N_2107);
nand U3633 (N_3633,N_2299,N_2624);
nor U3634 (N_3634,N_2727,N_2702);
nor U3635 (N_3635,N_2118,N_2620);
or U3636 (N_3636,N_2576,N_2841);
nor U3637 (N_3637,N_2685,N_2819);
and U3638 (N_3638,N_2120,N_2705);
nand U3639 (N_3639,N_2224,N_2528);
nand U3640 (N_3640,N_2380,N_2043);
nand U3641 (N_3641,N_2097,N_2459);
or U3642 (N_3642,N_2346,N_2178);
or U3643 (N_3643,N_2107,N_2523);
nor U3644 (N_3644,N_2166,N_2540);
nand U3645 (N_3645,N_2979,N_2461);
or U3646 (N_3646,N_2116,N_2934);
nor U3647 (N_3647,N_2594,N_2928);
or U3648 (N_3648,N_2723,N_2149);
nand U3649 (N_3649,N_2113,N_2378);
and U3650 (N_3650,N_2804,N_2721);
nand U3651 (N_3651,N_2523,N_2282);
xor U3652 (N_3652,N_2667,N_2220);
nand U3653 (N_3653,N_2147,N_2333);
nand U3654 (N_3654,N_2974,N_2365);
xor U3655 (N_3655,N_2983,N_2229);
and U3656 (N_3656,N_2887,N_2022);
and U3657 (N_3657,N_2014,N_2092);
or U3658 (N_3658,N_2407,N_2290);
and U3659 (N_3659,N_2499,N_2020);
and U3660 (N_3660,N_2480,N_2093);
or U3661 (N_3661,N_2246,N_2934);
nand U3662 (N_3662,N_2317,N_2509);
or U3663 (N_3663,N_2518,N_2562);
nand U3664 (N_3664,N_2477,N_2765);
nor U3665 (N_3665,N_2665,N_2404);
nor U3666 (N_3666,N_2663,N_2877);
nand U3667 (N_3667,N_2581,N_2269);
nand U3668 (N_3668,N_2062,N_2394);
or U3669 (N_3669,N_2388,N_2764);
nor U3670 (N_3670,N_2830,N_2555);
xnor U3671 (N_3671,N_2908,N_2602);
nor U3672 (N_3672,N_2928,N_2140);
nand U3673 (N_3673,N_2546,N_2304);
and U3674 (N_3674,N_2727,N_2909);
nor U3675 (N_3675,N_2498,N_2688);
xnor U3676 (N_3676,N_2313,N_2003);
and U3677 (N_3677,N_2029,N_2446);
nor U3678 (N_3678,N_2085,N_2025);
or U3679 (N_3679,N_2197,N_2729);
and U3680 (N_3680,N_2236,N_2459);
or U3681 (N_3681,N_2904,N_2453);
nand U3682 (N_3682,N_2590,N_2217);
nor U3683 (N_3683,N_2664,N_2282);
or U3684 (N_3684,N_2801,N_2202);
and U3685 (N_3685,N_2472,N_2928);
or U3686 (N_3686,N_2160,N_2456);
xnor U3687 (N_3687,N_2390,N_2606);
nor U3688 (N_3688,N_2392,N_2085);
nand U3689 (N_3689,N_2102,N_2181);
xnor U3690 (N_3690,N_2036,N_2784);
nand U3691 (N_3691,N_2896,N_2313);
and U3692 (N_3692,N_2339,N_2548);
nand U3693 (N_3693,N_2918,N_2861);
and U3694 (N_3694,N_2724,N_2049);
and U3695 (N_3695,N_2478,N_2574);
and U3696 (N_3696,N_2165,N_2713);
and U3697 (N_3697,N_2183,N_2387);
nand U3698 (N_3698,N_2256,N_2307);
and U3699 (N_3699,N_2798,N_2780);
nand U3700 (N_3700,N_2108,N_2364);
or U3701 (N_3701,N_2706,N_2646);
nor U3702 (N_3702,N_2245,N_2136);
or U3703 (N_3703,N_2761,N_2675);
nor U3704 (N_3704,N_2032,N_2555);
and U3705 (N_3705,N_2838,N_2250);
nand U3706 (N_3706,N_2734,N_2307);
or U3707 (N_3707,N_2575,N_2644);
and U3708 (N_3708,N_2172,N_2029);
or U3709 (N_3709,N_2863,N_2334);
xnor U3710 (N_3710,N_2971,N_2905);
nand U3711 (N_3711,N_2644,N_2953);
or U3712 (N_3712,N_2628,N_2786);
and U3713 (N_3713,N_2951,N_2660);
xor U3714 (N_3714,N_2119,N_2038);
and U3715 (N_3715,N_2715,N_2588);
nor U3716 (N_3716,N_2494,N_2686);
nand U3717 (N_3717,N_2604,N_2367);
nor U3718 (N_3718,N_2172,N_2304);
or U3719 (N_3719,N_2243,N_2784);
nor U3720 (N_3720,N_2942,N_2561);
and U3721 (N_3721,N_2378,N_2699);
nand U3722 (N_3722,N_2629,N_2260);
or U3723 (N_3723,N_2251,N_2562);
nand U3724 (N_3724,N_2200,N_2524);
and U3725 (N_3725,N_2440,N_2198);
nor U3726 (N_3726,N_2757,N_2837);
and U3727 (N_3727,N_2359,N_2120);
or U3728 (N_3728,N_2360,N_2237);
nand U3729 (N_3729,N_2744,N_2685);
or U3730 (N_3730,N_2267,N_2834);
nor U3731 (N_3731,N_2299,N_2541);
nand U3732 (N_3732,N_2919,N_2893);
and U3733 (N_3733,N_2673,N_2798);
nand U3734 (N_3734,N_2066,N_2981);
and U3735 (N_3735,N_2396,N_2190);
nand U3736 (N_3736,N_2484,N_2256);
nor U3737 (N_3737,N_2498,N_2117);
or U3738 (N_3738,N_2480,N_2753);
xor U3739 (N_3739,N_2361,N_2766);
xnor U3740 (N_3740,N_2371,N_2658);
nor U3741 (N_3741,N_2792,N_2852);
or U3742 (N_3742,N_2295,N_2048);
and U3743 (N_3743,N_2979,N_2077);
nand U3744 (N_3744,N_2186,N_2491);
nor U3745 (N_3745,N_2224,N_2567);
xnor U3746 (N_3746,N_2968,N_2535);
and U3747 (N_3747,N_2825,N_2883);
or U3748 (N_3748,N_2813,N_2714);
nor U3749 (N_3749,N_2491,N_2917);
nand U3750 (N_3750,N_2075,N_2653);
and U3751 (N_3751,N_2816,N_2650);
nand U3752 (N_3752,N_2639,N_2084);
nor U3753 (N_3753,N_2594,N_2991);
xor U3754 (N_3754,N_2039,N_2835);
xor U3755 (N_3755,N_2409,N_2191);
nor U3756 (N_3756,N_2739,N_2951);
xnor U3757 (N_3757,N_2800,N_2642);
and U3758 (N_3758,N_2126,N_2277);
or U3759 (N_3759,N_2802,N_2854);
nand U3760 (N_3760,N_2311,N_2682);
or U3761 (N_3761,N_2045,N_2077);
or U3762 (N_3762,N_2368,N_2472);
nand U3763 (N_3763,N_2035,N_2808);
nor U3764 (N_3764,N_2679,N_2288);
or U3765 (N_3765,N_2735,N_2476);
or U3766 (N_3766,N_2159,N_2302);
nand U3767 (N_3767,N_2017,N_2844);
and U3768 (N_3768,N_2786,N_2300);
xor U3769 (N_3769,N_2332,N_2374);
or U3770 (N_3770,N_2269,N_2080);
xor U3771 (N_3771,N_2437,N_2697);
xor U3772 (N_3772,N_2550,N_2232);
and U3773 (N_3773,N_2139,N_2396);
nand U3774 (N_3774,N_2618,N_2959);
nor U3775 (N_3775,N_2604,N_2339);
and U3776 (N_3776,N_2202,N_2573);
xor U3777 (N_3777,N_2805,N_2122);
nor U3778 (N_3778,N_2092,N_2901);
nor U3779 (N_3779,N_2919,N_2748);
nor U3780 (N_3780,N_2196,N_2429);
or U3781 (N_3781,N_2254,N_2100);
xnor U3782 (N_3782,N_2697,N_2527);
xnor U3783 (N_3783,N_2043,N_2625);
and U3784 (N_3784,N_2865,N_2882);
nor U3785 (N_3785,N_2597,N_2373);
nor U3786 (N_3786,N_2244,N_2182);
xnor U3787 (N_3787,N_2137,N_2381);
xor U3788 (N_3788,N_2869,N_2875);
nand U3789 (N_3789,N_2685,N_2251);
and U3790 (N_3790,N_2336,N_2716);
nand U3791 (N_3791,N_2957,N_2484);
nor U3792 (N_3792,N_2546,N_2564);
xor U3793 (N_3793,N_2514,N_2406);
and U3794 (N_3794,N_2052,N_2120);
xnor U3795 (N_3795,N_2699,N_2213);
nor U3796 (N_3796,N_2045,N_2410);
xor U3797 (N_3797,N_2613,N_2943);
nor U3798 (N_3798,N_2782,N_2772);
or U3799 (N_3799,N_2546,N_2388);
nand U3800 (N_3800,N_2792,N_2787);
xor U3801 (N_3801,N_2666,N_2657);
nor U3802 (N_3802,N_2558,N_2465);
xnor U3803 (N_3803,N_2283,N_2517);
xor U3804 (N_3804,N_2192,N_2649);
nand U3805 (N_3805,N_2409,N_2599);
or U3806 (N_3806,N_2357,N_2229);
and U3807 (N_3807,N_2235,N_2705);
or U3808 (N_3808,N_2618,N_2682);
nor U3809 (N_3809,N_2053,N_2727);
and U3810 (N_3810,N_2922,N_2688);
nand U3811 (N_3811,N_2945,N_2226);
nor U3812 (N_3812,N_2893,N_2235);
nor U3813 (N_3813,N_2939,N_2269);
xnor U3814 (N_3814,N_2882,N_2517);
xor U3815 (N_3815,N_2669,N_2704);
nor U3816 (N_3816,N_2623,N_2102);
xnor U3817 (N_3817,N_2347,N_2955);
xor U3818 (N_3818,N_2918,N_2331);
nor U3819 (N_3819,N_2112,N_2203);
nand U3820 (N_3820,N_2451,N_2457);
and U3821 (N_3821,N_2340,N_2022);
nor U3822 (N_3822,N_2513,N_2243);
or U3823 (N_3823,N_2517,N_2899);
and U3824 (N_3824,N_2665,N_2521);
nor U3825 (N_3825,N_2890,N_2553);
or U3826 (N_3826,N_2147,N_2768);
nor U3827 (N_3827,N_2989,N_2985);
nor U3828 (N_3828,N_2211,N_2395);
nor U3829 (N_3829,N_2328,N_2286);
xnor U3830 (N_3830,N_2336,N_2693);
and U3831 (N_3831,N_2239,N_2002);
nor U3832 (N_3832,N_2720,N_2746);
and U3833 (N_3833,N_2870,N_2056);
xnor U3834 (N_3834,N_2175,N_2080);
xnor U3835 (N_3835,N_2843,N_2351);
or U3836 (N_3836,N_2373,N_2378);
xor U3837 (N_3837,N_2458,N_2159);
nor U3838 (N_3838,N_2855,N_2308);
and U3839 (N_3839,N_2947,N_2378);
and U3840 (N_3840,N_2495,N_2769);
nand U3841 (N_3841,N_2978,N_2197);
xor U3842 (N_3842,N_2446,N_2899);
or U3843 (N_3843,N_2710,N_2004);
and U3844 (N_3844,N_2904,N_2726);
xor U3845 (N_3845,N_2630,N_2365);
nor U3846 (N_3846,N_2740,N_2611);
nor U3847 (N_3847,N_2402,N_2229);
and U3848 (N_3848,N_2958,N_2595);
nor U3849 (N_3849,N_2035,N_2741);
nor U3850 (N_3850,N_2463,N_2639);
or U3851 (N_3851,N_2868,N_2993);
and U3852 (N_3852,N_2503,N_2141);
nand U3853 (N_3853,N_2863,N_2244);
nor U3854 (N_3854,N_2862,N_2290);
and U3855 (N_3855,N_2222,N_2561);
and U3856 (N_3856,N_2405,N_2803);
nand U3857 (N_3857,N_2529,N_2292);
xor U3858 (N_3858,N_2024,N_2015);
and U3859 (N_3859,N_2616,N_2066);
xnor U3860 (N_3860,N_2809,N_2506);
or U3861 (N_3861,N_2744,N_2747);
and U3862 (N_3862,N_2563,N_2474);
xnor U3863 (N_3863,N_2015,N_2951);
or U3864 (N_3864,N_2209,N_2143);
xor U3865 (N_3865,N_2227,N_2359);
nand U3866 (N_3866,N_2315,N_2647);
or U3867 (N_3867,N_2743,N_2458);
nor U3868 (N_3868,N_2472,N_2796);
nand U3869 (N_3869,N_2792,N_2797);
nand U3870 (N_3870,N_2288,N_2613);
xnor U3871 (N_3871,N_2951,N_2919);
and U3872 (N_3872,N_2747,N_2046);
nor U3873 (N_3873,N_2547,N_2320);
and U3874 (N_3874,N_2897,N_2378);
nand U3875 (N_3875,N_2741,N_2548);
nor U3876 (N_3876,N_2631,N_2179);
and U3877 (N_3877,N_2593,N_2294);
nand U3878 (N_3878,N_2643,N_2249);
nand U3879 (N_3879,N_2913,N_2217);
nand U3880 (N_3880,N_2986,N_2818);
xor U3881 (N_3881,N_2927,N_2296);
or U3882 (N_3882,N_2151,N_2149);
and U3883 (N_3883,N_2487,N_2383);
and U3884 (N_3884,N_2142,N_2197);
and U3885 (N_3885,N_2063,N_2792);
xor U3886 (N_3886,N_2126,N_2755);
nand U3887 (N_3887,N_2134,N_2497);
and U3888 (N_3888,N_2850,N_2156);
xor U3889 (N_3889,N_2572,N_2512);
nand U3890 (N_3890,N_2245,N_2174);
nand U3891 (N_3891,N_2773,N_2135);
nand U3892 (N_3892,N_2977,N_2101);
xnor U3893 (N_3893,N_2071,N_2287);
xor U3894 (N_3894,N_2247,N_2515);
and U3895 (N_3895,N_2286,N_2545);
xor U3896 (N_3896,N_2571,N_2498);
and U3897 (N_3897,N_2888,N_2501);
nor U3898 (N_3898,N_2245,N_2323);
or U3899 (N_3899,N_2579,N_2451);
and U3900 (N_3900,N_2395,N_2242);
and U3901 (N_3901,N_2109,N_2052);
nand U3902 (N_3902,N_2691,N_2884);
nand U3903 (N_3903,N_2568,N_2580);
and U3904 (N_3904,N_2477,N_2498);
xor U3905 (N_3905,N_2990,N_2192);
and U3906 (N_3906,N_2132,N_2893);
nand U3907 (N_3907,N_2483,N_2817);
and U3908 (N_3908,N_2046,N_2769);
nand U3909 (N_3909,N_2685,N_2432);
xor U3910 (N_3910,N_2775,N_2332);
xnor U3911 (N_3911,N_2465,N_2932);
or U3912 (N_3912,N_2945,N_2023);
nor U3913 (N_3913,N_2681,N_2862);
or U3914 (N_3914,N_2526,N_2569);
nand U3915 (N_3915,N_2870,N_2585);
and U3916 (N_3916,N_2785,N_2154);
xnor U3917 (N_3917,N_2439,N_2950);
and U3918 (N_3918,N_2946,N_2072);
or U3919 (N_3919,N_2391,N_2366);
or U3920 (N_3920,N_2319,N_2141);
nor U3921 (N_3921,N_2854,N_2347);
and U3922 (N_3922,N_2140,N_2705);
nor U3923 (N_3923,N_2465,N_2392);
and U3924 (N_3924,N_2847,N_2673);
xnor U3925 (N_3925,N_2289,N_2113);
or U3926 (N_3926,N_2599,N_2650);
nor U3927 (N_3927,N_2010,N_2443);
and U3928 (N_3928,N_2113,N_2590);
and U3929 (N_3929,N_2152,N_2028);
xor U3930 (N_3930,N_2226,N_2075);
and U3931 (N_3931,N_2567,N_2331);
nor U3932 (N_3932,N_2156,N_2780);
nand U3933 (N_3933,N_2585,N_2705);
or U3934 (N_3934,N_2342,N_2295);
and U3935 (N_3935,N_2416,N_2952);
and U3936 (N_3936,N_2056,N_2928);
and U3937 (N_3937,N_2842,N_2692);
and U3938 (N_3938,N_2657,N_2300);
and U3939 (N_3939,N_2292,N_2161);
nor U3940 (N_3940,N_2318,N_2380);
xor U3941 (N_3941,N_2938,N_2689);
nor U3942 (N_3942,N_2157,N_2092);
and U3943 (N_3943,N_2805,N_2142);
nor U3944 (N_3944,N_2603,N_2464);
nor U3945 (N_3945,N_2977,N_2454);
nand U3946 (N_3946,N_2200,N_2118);
nor U3947 (N_3947,N_2820,N_2666);
xor U3948 (N_3948,N_2929,N_2676);
nand U3949 (N_3949,N_2459,N_2309);
or U3950 (N_3950,N_2518,N_2862);
and U3951 (N_3951,N_2286,N_2951);
and U3952 (N_3952,N_2428,N_2524);
xnor U3953 (N_3953,N_2750,N_2033);
or U3954 (N_3954,N_2794,N_2193);
or U3955 (N_3955,N_2999,N_2329);
and U3956 (N_3956,N_2969,N_2662);
nor U3957 (N_3957,N_2186,N_2913);
and U3958 (N_3958,N_2484,N_2635);
and U3959 (N_3959,N_2144,N_2211);
and U3960 (N_3960,N_2410,N_2383);
nand U3961 (N_3961,N_2285,N_2761);
or U3962 (N_3962,N_2678,N_2964);
xor U3963 (N_3963,N_2790,N_2435);
or U3964 (N_3964,N_2176,N_2334);
or U3965 (N_3965,N_2314,N_2293);
or U3966 (N_3966,N_2928,N_2361);
nor U3967 (N_3967,N_2086,N_2392);
nor U3968 (N_3968,N_2143,N_2761);
or U3969 (N_3969,N_2019,N_2965);
or U3970 (N_3970,N_2096,N_2355);
nand U3971 (N_3971,N_2106,N_2001);
or U3972 (N_3972,N_2525,N_2251);
nand U3973 (N_3973,N_2075,N_2429);
xor U3974 (N_3974,N_2781,N_2837);
xor U3975 (N_3975,N_2435,N_2292);
xor U3976 (N_3976,N_2549,N_2887);
or U3977 (N_3977,N_2453,N_2620);
and U3978 (N_3978,N_2267,N_2258);
or U3979 (N_3979,N_2853,N_2580);
nand U3980 (N_3980,N_2745,N_2929);
nand U3981 (N_3981,N_2821,N_2411);
and U3982 (N_3982,N_2097,N_2177);
and U3983 (N_3983,N_2936,N_2762);
nand U3984 (N_3984,N_2936,N_2659);
or U3985 (N_3985,N_2931,N_2734);
nand U3986 (N_3986,N_2958,N_2731);
nand U3987 (N_3987,N_2567,N_2202);
xnor U3988 (N_3988,N_2529,N_2683);
and U3989 (N_3989,N_2843,N_2121);
nor U3990 (N_3990,N_2781,N_2263);
or U3991 (N_3991,N_2691,N_2762);
and U3992 (N_3992,N_2299,N_2944);
and U3993 (N_3993,N_2719,N_2127);
and U3994 (N_3994,N_2032,N_2589);
nand U3995 (N_3995,N_2756,N_2629);
xor U3996 (N_3996,N_2462,N_2650);
nor U3997 (N_3997,N_2423,N_2892);
nand U3998 (N_3998,N_2536,N_2566);
or U3999 (N_3999,N_2215,N_2577);
xnor U4000 (N_4000,N_3380,N_3034);
nor U4001 (N_4001,N_3867,N_3441);
nand U4002 (N_4002,N_3763,N_3125);
and U4003 (N_4003,N_3201,N_3445);
nand U4004 (N_4004,N_3951,N_3435);
and U4005 (N_4005,N_3624,N_3744);
and U4006 (N_4006,N_3946,N_3560);
and U4007 (N_4007,N_3578,N_3818);
nand U4008 (N_4008,N_3926,N_3796);
nor U4009 (N_4009,N_3154,N_3456);
nor U4010 (N_4010,N_3277,N_3257);
and U4011 (N_4011,N_3110,N_3907);
nor U4012 (N_4012,N_3056,N_3516);
nand U4013 (N_4013,N_3359,N_3647);
and U4014 (N_4014,N_3054,N_3439);
or U4015 (N_4015,N_3065,N_3303);
xor U4016 (N_4016,N_3734,N_3904);
xnor U4017 (N_4017,N_3640,N_3613);
and U4018 (N_4018,N_3750,N_3851);
nor U4019 (N_4019,N_3238,N_3780);
or U4020 (N_4020,N_3124,N_3007);
nand U4021 (N_4021,N_3333,N_3714);
nor U4022 (N_4022,N_3950,N_3683);
and U4023 (N_4023,N_3520,N_3292);
nor U4024 (N_4024,N_3461,N_3067);
or U4025 (N_4025,N_3944,N_3166);
or U4026 (N_4026,N_3972,N_3331);
and U4027 (N_4027,N_3934,N_3343);
nand U4028 (N_4028,N_3369,N_3535);
nand U4029 (N_4029,N_3163,N_3383);
nand U4030 (N_4030,N_3595,N_3409);
xnor U4031 (N_4031,N_3675,N_3894);
nand U4032 (N_4032,N_3430,N_3008);
xor U4033 (N_4033,N_3475,N_3116);
nand U4034 (N_4034,N_3316,N_3623);
nand U4035 (N_4035,N_3919,N_3255);
nor U4036 (N_4036,N_3226,N_3345);
xnor U4037 (N_4037,N_3498,N_3442);
nor U4038 (N_4038,N_3768,N_3283);
nor U4039 (N_4039,N_3853,N_3577);
nor U4040 (N_4040,N_3385,N_3572);
nor U4041 (N_4041,N_3284,N_3378);
xor U4042 (N_4042,N_3381,N_3726);
xnor U4043 (N_4043,N_3455,N_3499);
or U4044 (N_4044,N_3061,N_3270);
and U4045 (N_4045,N_3155,N_3846);
nor U4046 (N_4046,N_3178,N_3622);
or U4047 (N_4047,N_3957,N_3326);
and U4048 (N_4048,N_3458,N_3738);
and U4049 (N_4049,N_3421,N_3285);
nor U4050 (N_4050,N_3569,N_3694);
nor U4051 (N_4051,N_3874,N_3252);
nand U4052 (N_4052,N_3674,N_3684);
nand U4053 (N_4053,N_3899,N_3229);
nand U4054 (N_4054,N_3481,N_3393);
xor U4055 (N_4055,N_3519,N_3510);
or U4056 (N_4056,N_3123,N_3996);
nor U4057 (N_4057,N_3398,N_3183);
or U4058 (N_4058,N_3993,N_3011);
or U4059 (N_4059,N_3876,N_3440);
and U4060 (N_4060,N_3882,N_3296);
or U4061 (N_4061,N_3096,N_3702);
xnor U4062 (N_4062,N_3731,N_3718);
or U4063 (N_4063,N_3666,N_3689);
or U4064 (N_4064,N_3099,N_3809);
nor U4065 (N_4065,N_3823,N_3098);
and U4066 (N_4066,N_3453,N_3754);
xnor U4067 (N_4067,N_3676,N_3888);
xnor U4068 (N_4068,N_3737,N_3810);
and U4069 (N_4069,N_3749,N_3928);
xnor U4070 (N_4070,N_3949,N_3638);
or U4071 (N_4071,N_3133,N_3999);
and U4072 (N_4072,N_3969,N_3959);
nor U4073 (N_4073,N_3661,N_3566);
nand U4074 (N_4074,N_3747,N_3087);
and U4075 (N_4075,N_3088,N_3792);
and U4076 (N_4076,N_3690,N_3571);
or U4077 (N_4077,N_3653,N_3134);
xnor U4078 (N_4078,N_3606,N_3799);
or U4079 (N_4079,N_3873,N_3554);
xor U4080 (N_4080,N_3587,N_3095);
nor U4081 (N_4081,N_3740,N_3827);
nand U4082 (N_4082,N_3299,N_3289);
or U4083 (N_4083,N_3309,N_3663);
and U4084 (N_4084,N_3035,N_3507);
nor U4085 (N_4085,N_3018,N_3091);
or U4086 (N_4086,N_3982,N_3839);
nand U4087 (N_4087,N_3512,N_3093);
nand U4088 (N_4088,N_3148,N_3161);
xor U4089 (N_4089,N_3408,N_3086);
and U4090 (N_4090,N_3636,N_3621);
nor U4091 (N_4091,N_3245,N_3649);
or U4092 (N_4092,N_3070,N_3930);
or U4093 (N_4093,N_3149,N_3174);
and U4094 (N_4094,N_3826,N_3915);
nor U4095 (N_4095,N_3495,N_3457);
nand U4096 (N_4096,N_3772,N_3527);
and U4097 (N_4097,N_3135,N_3937);
nor U4098 (N_4098,N_3616,N_3650);
nor U4099 (N_4099,N_3964,N_3274);
nor U4100 (N_4100,N_3231,N_3513);
nor U4101 (N_4101,N_3199,N_3175);
and U4102 (N_4102,N_3139,N_3480);
and U4103 (N_4103,N_3487,N_3269);
and U4104 (N_4104,N_3364,N_3619);
xnor U4105 (N_4105,N_3691,N_3464);
xnor U4106 (N_4106,N_3195,N_3041);
nor U4107 (N_4107,N_3544,N_3902);
nand U4108 (N_4108,N_3806,N_3465);
nor U4109 (N_4109,N_3762,N_3643);
nand U4110 (N_4110,N_3153,N_3479);
or U4111 (N_4111,N_3294,N_3076);
or U4112 (N_4112,N_3221,N_3373);
or U4113 (N_4113,N_3751,N_3743);
or U4114 (N_4114,N_3916,N_3488);
nand U4115 (N_4115,N_3366,N_3119);
nand U4116 (N_4116,N_3049,N_3720);
nand U4117 (N_4117,N_3844,N_3576);
or U4118 (N_4118,N_3805,N_3173);
and U4119 (N_4119,N_3412,N_3489);
xnor U4120 (N_4120,N_3971,N_3109);
and U4121 (N_4121,N_3868,N_3525);
and U4122 (N_4122,N_3586,N_3454);
and U4123 (N_4123,N_3908,N_3822);
or U4124 (N_4124,N_3137,N_3781);
nor U4125 (N_4125,N_3790,N_3633);
xnor U4126 (N_4126,N_3290,N_3552);
nor U4127 (N_4127,N_3236,N_3377);
nor U4128 (N_4128,N_3992,N_3813);
or U4129 (N_4129,N_3043,N_3987);
or U4130 (N_4130,N_3942,N_3047);
nor U4131 (N_4131,N_3074,N_3497);
or U4132 (N_4132,N_3769,N_3042);
or U4133 (N_4133,N_3319,N_3561);
xnor U4134 (N_4134,N_3699,N_3205);
nand U4135 (N_4135,N_3835,N_3528);
nor U4136 (N_4136,N_3058,N_3594);
xor U4137 (N_4137,N_3778,N_3077);
nand U4138 (N_4138,N_3005,N_3798);
nor U4139 (N_4139,N_3697,N_3609);
nand U4140 (N_4140,N_3462,N_3884);
nand U4141 (N_4141,N_3977,N_3436);
and U4142 (N_4142,N_3526,N_3838);
or U4143 (N_4143,N_3390,N_3797);
xor U4144 (N_4144,N_3418,N_3128);
xor U4145 (N_4145,N_3898,N_3776);
nor U4146 (N_4146,N_3046,N_3320);
nor U4147 (N_4147,N_3816,N_3931);
and U4148 (N_4148,N_3686,N_3237);
or U4149 (N_4149,N_3673,N_3985);
and U4150 (N_4150,N_3910,N_3228);
nand U4151 (N_4151,N_3524,N_3431);
and U4152 (N_4152,N_3272,N_3815);
or U4153 (N_4153,N_3280,N_3502);
or U4154 (N_4154,N_3962,N_3538);
or U4155 (N_4155,N_3695,N_3997);
or U4156 (N_4156,N_3176,N_3618);
nor U4157 (N_4157,N_3515,N_3830);
xnor U4158 (N_4158,N_3313,N_3909);
and U4159 (N_4159,N_3534,N_3786);
and U4160 (N_4160,N_3917,N_3596);
and U4161 (N_4161,N_3306,N_3793);
nor U4162 (N_4162,N_3395,N_3546);
or U4163 (N_4163,N_3376,N_3896);
nor U4164 (N_4164,N_3384,N_3933);
or U4165 (N_4165,N_3521,N_3387);
or U4166 (N_4166,N_3328,N_3388);
xor U4167 (N_4167,N_3533,N_3104);
and U4168 (N_4168,N_3753,N_3886);
xnor U4169 (N_4169,N_3438,N_3113);
or U4170 (N_4170,N_3672,N_3282);
nand U4171 (N_4171,N_3869,N_3644);
or U4172 (N_4172,N_3020,N_3048);
xnor U4173 (N_4173,N_3836,N_3021);
nor U4174 (N_4174,N_3870,N_3471);
or U4175 (N_4175,N_3703,N_3016);
xnor U4176 (N_4176,N_3182,N_3967);
or U4177 (N_4177,N_3925,N_3954);
nand U4178 (N_4178,N_3019,N_3185);
xnor U4179 (N_4179,N_3975,N_3062);
nand U4180 (N_4180,N_3474,N_3045);
or U4181 (N_4181,N_3834,N_3730);
or U4182 (N_4182,N_3989,N_3260);
nand U4183 (N_4183,N_3652,N_3208);
nor U4184 (N_4184,N_3444,N_3311);
nor U4185 (N_4185,N_3463,N_3540);
and U4186 (N_4186,N_3230,N_3591);
and U4187 (N_4187,N_3670,N_3298);
and U4188 (N_4188,N_3103,N_3582);
or U4189 (N_4189,N_3028,N_3852);
nand U4190 (N_4190,N_3847,N_3550);
nor U4191 (N_4191,N_3404,N_3355);
nand U4192 (N_4192,N_3181,N_3801);
nand U4193 (N_4193,N_3746,N_3217);
or U4194 (N_4194,N_3476,N_3363);
nor U4195 (N_4195,N_3685,N_3988);
or U4196 (N_4196,N_3064,N_3548);
xnor U4197 (N_4197,N_3562,N_3850);
nand U4198 (N_4198,N_3317,N_3914);
nor U4199 (N_4199,N_3211,N_3143);
or U4200 (N_4200,N_3227,N_3518);
nand U4201 (N_4201,N_3551,N_3820);
or U4202 (N_4202,N_3825,N_3681);
or U4203 (N_4203,N_3129,N_3422);
nor U4204 (N_4204,N_3913,N_3529);
xor U4205 (N_4205,N_3994,N_3938);
and U4206 (N_4206,N_3607,N_3642);
nor U4207 (N_4207,N_3770,N_3010);
nor U4208 (N_4208,N_3553,N_3761);
nand U4209 (N_4209,N_3105,N_3027);
nand U4210 (N_4210,N_3878,N_3563);
and U4211 (N_4211,N_3308,N_3943);
and U4212 (N_4212,N_3955,N_3541);
or U4213 (N_4213,N_3581,N_3953);
nand U4214 (N_4214,N_3482,N_3402);
xor U4215 (N_4215,N_3648,N_3947);
nor U4216 (N_4216,N_3242,N_3322);
nor U4217 (N_4217,N_3278,N_3263);
xnor U4218 (N_4218,N_3705,N_3031);
and U4219 (N_4219,N_3984,N_3060);
and U4220 (N_4220,N_3452,N_3592);
nor U4221 (N_4221,N_3244,N_3759);
nor U4222 (N_4222,N_3239,N_3615);
xor U4223 (N_4223,N_3156,N_3940);
xor U4224 (N_4224,N_3117,N_3542);
nor U4225 (N_4225,N_3433,N_3141);
nor U4226 (N_4226,N_3234,N_3371);
and U4227 (N_4227,N_3523,N_3410);
and U4228 (N_4228,N_3849,N_3789);
xor U4229 (N_4229,N_3579,N_3094);
nor U4230 (N_4230,N_3503,N_3118);
nor U4231 (N_4231,N_3122,N_3680);
and U4232 (N_4232,N_3921,N_3817);
and U4233 (N_4233,N_3708,N_3501);
or U4234 (N_4234,N_3437,N_3036);
nand U4235 (N_4235,N_3396,N_3108);
nor U4236 (N_4236,N_3083,N_3192);
nor U4237 (N_4237,N_3202,N_3449);
nor U4238 (N_4238,N_3078,N_3918);
nor U4239 (N_4239,N_3980,N_3669);
or U4240 (N_4240,N_3427,N_3875);
and U4241 (N_4241,N_3434,N_3981);
and U4242 (N_4242,N_3583,N_3698);
nand U4243 (N_4243,N_3812,N_3291);
or U4244 (N_4244,N_3127,N_3267);
nand U4245 (N_4245,N_3679,N_3017);
xor U4246 (N_4246,N_3911,N_3171);
and U4247 (N_4247,N_3106,N_3459);
nand U4248 (N_4248,N_3920,N_3511);
nand U4249 (N_4249,N_3531,N_3353);
xnor U4250 (N_4250,N_3811,N_3991);
xnor U4251 (N_4251,N_3871,N_3700);
or U4252 (N_4252,N_3146,N_3138);
nor U4253 (N_4253,N_3030,N_3415);
nor U4254 (N_4254,N_3614,N_3120);
xnor U4255 (N_4255,N_3351,N_3370);
nand U4256 (N_4256,N_3903,N_3250);
xor U4257 (N_4257,N_3053,N_3262);
and U4258 (N_4258,N_3314,N_3411);
or U4259 (N_4259,N_3634,N_3855);
nor U4260 (N_4260,N_3736,N_3960);
or U4261 (N_4261,N_3469,N_3025);
or U4262 (N_4262,N_3145,N_3575);
nand U4263 (N_4263,N_3814,N_3391);
nand U4264 (N_4264,N_3216,N_3704);
nor U4265 (N_4265,N_3342,N_3241);
nor U4266 (N_4266,N_3608,N_3808);
nand U4267 (N_4267,N_3349,N_3100);
or U4268 (N_4268,N_3764,N_3573);
and U4269 (N_4269,N_3968,N_3382);
and U4270 (N_4270,N_3630,N_3420);
nand U4271 (N_4271,N_3413,N_3733);
and U4272 (N_4272,N_3246,N_3824);
and U4273 (N_4273,N_3361,N_3939);
nor U4274 (N_4274,N_3490,N_3678);
nand U4275 (N_4275,N_3522,N_3492);
xor U4276 (N_4276,N_3073,N_3861);
nor U4277 (N_4277,N_3215,N_3641);
xor U4278 (N_4278,N_3767,N_3900);
xor U4279 (N_4279,N_3929,N_3115);
and U4280 (N_4280,N_3788,N_3131);
and U4281 (N_4281,N_3998,N_3325);
nand U4282 (N_4282,N_3995,N_3159);
nand U4283 (N_4283,N_3033,N_3549);
nor U4284 (N_4284,N_3629,N_3745);
xnor U4285 (N_4285,N_3374,N_3038);
and U4286 (N_4286,N_3865,N_3170);
or U4287 (N_4287,N_3610,N_3662);
and U4288 (N_4288,N_3240,N_3080);
or U4289 (N_4289,N_3728,N_3039);
nor U4290 (N_4290,N_3843,N_3771);
nor U4291 (N_4291,N_3978,N_3539);
and U4292 (N_4292,N_3198,N_3601);
nor U4293 (N_4293,N_3318,N_3766);
nor U4294 (N_4294,N_3254,N_3264);
nor U4295 (N_4295,N_3777,N_3286);
nor U4296 (N_4296,N_3574,N_3256);
nor U4297 (N_4297,N_3785,N_3002);
nor U4298 (N_4298,N_3187,N_3639);
or U4299 (N_4299,N_3271,N_3169);
nor U4300 (N_4300,N_3783,N_3090);
or U4301 (N_4301,N_3713,N_3179);
or U4302 (N_4302,N_3935,N_3625);
xor U4303 (N_4303,N_3258,N_3547);
or U4304 (N_4304,N_3321,N_3451);
nand U4305 (N_4305,N_3660,N_3514);
and U4306 (N_4306,N_3696,N_3952);
nand U4307 (N_4307,N_3188,N_3506);
or U4308 (N_4308,N_3446,N_3426);
nor U4309 (N_4309,N_3190,N_3687);
xor U4310 (N_4310,N_3140,N_3779);
xor U4311 (N_4311,N_3668,N_3339);
and U4312 (N_4312,N_3787,N_3840);
xor U4313 (N_4313,N_3079,N_3379);
xnor U4314 (N_4314,N_3302,N_3219);
xor U4315 (N_4315,N_3253,N_3247);
xnor U4316 (N_4316,N_3288,N_3829);
nor U4317 (N_4317,N_3348,N_3715);
or U4318 (N_4318,N_3013,N_3860);
nor U4319 (N_4319,N_3037,N_3032);
xor U4320 (N_4320,N_3213,N_3248);
nor U4321 (N_4321,N_3722,N_3602);
or U4322 (N_4322,N_3890,N_3323);
xor U4323 (N_4323,N_3279,N_3448);
xor U4324 (N_4324,N_3347,N_3617);
nor U4325 (N_4325,N_3611,N_3880);
and U4326 (N_4326,N_3665,N_3329);
xor U4327 (N_4327,N_3259,N_3559);
nor U4328 (N_4328,N_3367,N_3191);
or U4329 (N_4329,N_3932,N_3948);
or U4330 (N_4330,N_3121,N_3417);
nand U4331 (N_4331,N_3877,N_3428);
nand U4332 (N_4332,N_3837,N_3832);
nor U4333 (N_4333,N_3389,N_3494);
and U4334 (N_4334,N_3450,N_3335);
or U4335 (N_4335,N_3407,N_3414);
or U4336 (N_4336,N_3416,N_3209);
xnor U4337 (N_4337,N_3655,N_3337);
nor U4338 (N_4338,N_3599,N_3147);
and U4339 (N_4339,N_3168,N_3397);
nor U4340 (N_4340,N_3249,N_3297);
nand U4341 (N_4341,N_3470,N_3004);
nor U4342 (N_4342,N_3082,N_3848);
or U4343 (N_4343,N_3530,N_3084);
and U4344 (N_4344,N_3775,N_3075);
and U4345 (N_4345,N_3177,N_3399);
nor U4346 (N_4346,N_3941,N_3265);
and U4347 (N_4347,N_3107,N_3375);
nand U4348 (N_4348,N_3210,N_3891);
nor U4349 (N_4349,N_3301,N_3558);
nand U4350 (N_4350,N_3637,N_3986);
nor U4351 (N_4351,N_3483,N_3859);
and U4352 (N_4352,N_3627,N_3312);
nand U4353 (N_4353,N_3597,N_3620);
nor U4354 (N_4354,N_3556,N_3424);
or U4355 (N_4355,N_3220,N_3307);
xor U4356 (N_4356,N_3102,N_3612);
and U4357 (N_4357,N_3287,N_3719);
nand U4358 (N_4358,N_3365,N_3752);
and U4359 (N_4359,N_3332,N_3631);
xnor U4360 (N_4360,N_3200,N_3493);
nand U4361 (N_4361,N_3132,N_3701);
xnor U4362 (N_4362,N_3782,N_3203);
xor U4363 (N_4363,N_3895,N_3905);
and U4364 (N_4364,N_3567,N_3945);
nor U4365 (N_4365,N_3261,N_3727);
nor U4366 (N_4366,N_3589,N_3310);
xor U4367 (N_4367,N_3757,N_3545);
or U4368 (N_4368,N_3057,N_3197);
and U4369 (N_4369,N_3026,N_3887);
nor U4370 (N_4370,N_3923,N_3273);
nand U4371 (N_4371,N_3225,N_3509);
nand U4372 (N_4372,N_3965,N_3707);
nor U4373 (N_4373,N_3063,N_3425);
nand U4374 (N_4374,N_3906,N_3496);
and U4375 (N_4375,N_3305,N_3406);
nor U4376 (N_4376,N_3092,N_3144);
nand U4377 (N_4377,N_3664,N_3350);
nand U4378 (N_4378,N_3603,N_3330);
and U4379 (N_4379,N_3646,N_3341);
and U4380 (N_4380,N_3023,N_3114);
nor U4381 (N_4381,N_3344,N_3739);
nand U4382 (N_4382,N_3774,N_3963);
or U4383 (N_4383,N_3006,N_3354);
nor U4384 (N_4384,N_3845,N_3863);
and U4385 (N_4385,N_3568,N_3150);
nor U4386 (N_4386,N_3543,N_3508);
xnor U4387 (N_4387,N_3158,N_3628);
xor U4388 (N_4388,N_3447,N_3748);
nor U4389 (N_4389,N_3632,N_3866);
nand U4390 (N_4390,N_3276,N_3912);
nor U4391 (N_4391,N_3677,N_3505);
and U4392 (N_4392,N_3651,N_3142);
nand U4393 (N_4393,N_3765,N_3165);
xnor U4394 (N_4394,N_3710,N_3266);
nand U4395 (N_4395,N_3214,N_3394);
nand U4396 (N_4396,N_3386,N_3883);
and U4397 (N_4397,N_3467,N_3184);
xnor U4398 (N_4398,N_3059,N_3012);
nor U4399 (N_4399,N_3725,N_3066);
nand U4400 (N_4400,N_3983,N_3593);
and U4401 (N_4401,N_3657,N_3819);
nand U4402 (N_4402,N_3500,N_3001);
nand U4403 (N_4403,N_3040,N_3468);
xor U4404 (N_4404,N_3485,N_3961);
nor U4405 (N_4405,N_3072,N_3218);
xnor U4406 (N_4406,N_3052,N_3716);
and U4407 (N_4407,N_3709,N_3207);
nand U4408 (N_4408,N_3491,N_3590);
or U4409 (N_4409,N_3659,N_3517);
and U4410 (N_4410,N_3189,N_3532);
nand U4411 (N_4411,N_3976,N_3854);
nand U4412 (N_4412,N_3164,N_3862);
nor U4413 (N_4413,N_3014,N_3403);
or U4414 (N_4414,N_3055,N_3268);
xnor U4415 (N_4415,N_3232,N_3804);
xnor U4416 (N_4416,N_3717,N_3802);
and U4417 (N_4417,N_3372,N_3966);
or U4418 (N_4418,N_3791,N_3224);
and U4419 (N_4419,N_3885,N_3243);
xnor U4420 (N_4420,N_3600,N_3443);
and U4421 (N_4421,N_3022,N_3085);
xnor U4422 (N_4422,N_3927,N_3688);
or U4423 (N_4423,N_3473,N_3193);
or U4424 (N_4424,N_3024,N_3828);
and U4425 (N_4425,N_3741,N_3223);
or U4426 (N_4426,N_3429,N_3295);
xnor U4427 (N_4427,N_3009,N_3857);
nor U4428 (N_4428,N_3300,N_3340);
nor U4429 (N_4429,N_3588,N_3605);
nor U4430 (N_4430,N_3901,N_3864);
xnor U4431 (N_4431,N_3357,N_3758);
nor U4432 (N_4432,N_3069,N_3212);
nor U4433 (N_4433,N_3101,N_3356);
nor U4434 (N_4434,N_3570,N_3186);
xor U4435 (N_4435,N_3841,N_3979);
and U4436 (N_4436,N_3784,N_3706);
nand U4437 (N_4437,N_3327,N_3821);
nand U4438 (N_4438,N_3856,N_3275);
and U4439 (N_4439,N_3233,N_3051);
and U4440 (N_4440,N_3029,N_3050);
nor U4441 (N_4441,N_3405,N_3922);
or U4442 (N_4442,N_3654,N_3881);
xor U4443 (N_4443,N_3112,N_3111);
and U4444 (N_4444,N_3478,N_3831);
and U4445 (N_4445,N_3729,N_3157);
nand U4446 (N_4446,N_3897,N_3251);
nor U4447 (N_4447,N_3973,N_3315);
xor U4448 (N_4448,N_3162,N_3504);
or U4449 (N_4449,N_3564,N_3097);
and U4450 (N_4450,N_3484,N_3742);
xnor U4451 (N_4451,N_3760,N_3537);
nor U4452 (N_4452,N_3151,N_3721);
or U4453 (N_4453,N_3194,N_3723);
nand U4454 (N_4454,N_3368,N_3172);
and U4455 (N_4455,N_3803,N_3071);
or U4456 (N_4456,N_3180,N_3800);
and U4457 (N_4457,N_3152,N_3756);
xor U4458 (N_4458,N_3711,N_3842);
or U4459 (N_4459,N_3336,N_3585);
or U4460 (N_4460,N_3580,N_3324);
nor U4461 (N_4461,N_3735,N_3423);
nand U4462 (N_4462,N_3126,N_3858);
or U4463 (N_4463,N_3724,N_3773);
or U4464 (N_4464,N_3352,N_3626);
and U4465 (N_4465,N_3555,N_3432);
nand U4466 (N_4466,N_3712,N_3206);
nand U4467 (N_4467,N_3362,N_3732);
nor U4468 (N_4468,N_3892,N_3003);
nand U4469 (N_4469,N_3936,N_3604);
and U4470 (N_4470,N_3130,N_3807);
and U4471 (N_4471,N_3956,N_3879);
and U4472 (N_4472,N_3346,N_3833);
or U4473 (N_4473,N_3281,N_3068);
or U4474 (N_4474,N_3645,N_3692);
or U4475 (N_4475,N_3667,N_3682);
nor U4476 (N_4476,N_3160,N_3401);
and U4477 (N_4477,N_3460,N_3477);
nand U4478 (N_4478,N_3755,N_3958);
nand U4479 (N_4479,N_3472,N_3338);
and U4480 (N_4480,N_3671,N_3893);
xor U4481 (N_4481,N_3656,N_3990);
nand U4482 (N_4482,N_3044,N_3584);
nor U4483 (N_4483,N_3794,N_3974);
xnor U4484 (N_4484,N_3196,N_3081);
nand U4485 (N_4485,N_3000,N_3304);
xnor U4486 (N_4486,N_3222,N_3872);
xor U4487 (N_4487,N_3598,N_3486);
nand U4488 (N_4488,N_3400,N_3970);
nor U4489 (N_4489,N_3565,N_3924);
nor U4490 (N_4490,N_3360,N_3204);
xor U4491 (N_4491,N_3795,N_3167);
and U4492 (N_4492,N_3693,N_3658);
or U4493 (N_4493,N_3358,N_3557);
xor U4494 (N_4494,N_3466,N_3419);
and U4495 (N_4495,N_3089,N_3334);
nand U4496 (N_4496,N_3889,N_3136);
xor U4497 (N_4497,N_3235,N_3015);
nand U4498 (N_4498,N_3536,N_3293);
nor U4499 (N_4499,N_3635,N_3392);
or U4500 (N_4500,N_3598,N_3335);
nor U4501 (N_4501,N_3077,N_3803);
or U4502 (N_4502,N_3333,N_3182);
or U4503 (N_4503,N_3975,N_3940);
or U4504 (N_4504,N_3627,N_3464);
and U4505 (N_4505,N_3465,N_3855);
and U4506 (N_4506,N_3864,N_3071);
xor U4507 (N_4507,N_3901,N_3768);
and U4508 (N_4508,N_3092,N_3930);
or U4509 (N_4509,N_3265,N_3817);
xnor U4510 (N_4510,N_3918,N_3578);
or U4511 (N_4511,N_3638,N_3951);
and U4512 (N_4512,N_3174,N_3755);
and U4513 (N_4513,N_3909,N_3048);
xnor U4514 (N_4514,N_3881,N_3220);
nor U4515 (N_4515,N_3037,N_3858);
or U4516 (N_4516,N_3630,N_3352);
and U4517 (N_4517,N_3173,N_3728);
xnor U4518 (N_4518,N_3575,N_3456);
xnor U4519 (N_4519,N_3349,N_3126);
nand U4520 (N_4520,N_3282,N_3205);
and U4521 (N_4521,N_3486,N_3842);
nor U4522 (N_4522,N_3399,N_3210);
nand U4523 (N_4523,N_3244,N_3449);
nand U4524 (N_4524,N_3264,N_3135);
or U4525 (N_4525,N_3491,N_3087);
and U4526 (N_4526,N_3602,N_3570);
and U4527 (N_4527,N_3449,N_3294);
and U4528 (N_4528,N_3486,N_3707);
nor U4529 (N_4529,N_3601,N_3595);
and U4530 (N_4530,N_3885,N_3273);
and U4531 (N_4531,N_3414,N_3246);
nand U4532 (N_4532,N_3434,N_3193);
xor U4533 (N_4533,N_3751,N_3797);
nand U4534 (N_4534,N_3915,N_3422);
and U4535 (N_4535,N_3317,N_3934);
nor U4536 (N_4536,N_3527,N_3245);
nand U4537 (N_4537,N_3989,N_3528);
nand U4538 (N_4538,N_3763,N_3605);
and U4539 (N_4539,N_3719,N_3681);
and U4540 (N_4540,N_3113,N_3161);
nand U4541 (N_4541,N_3154,N_3340);
nor U4542 (N_4542,N_3689,N_3320);
nand U4543 (N_4543,N_3001,N_3412);
nor U4544 (N_4544,N_3355,N_3703);
or U4545 (N_4545,N_3342,N_3349);
nand U4546 (N_4546,N_3534,N_3307);
or U4547 (N_4547,N_3976,N_3280);
xor U4548 (N_4548,N_3362,N_3617);
or U4549 (N_4549,N_3165,N_3877);
and U4550 (N_4550,N_3129,N_3179);
or U4551 (N_4551,N_3779,N_3765);
nand U4552 (N_4552,N_3433,N_3554);
or U4553 (N_4553,N_3661,N_3808);
nor U4554 (N_4554,N_3796,N_3880);
xor U4555 (N_4555,N_3980,N_3526);
xor U4556 (N_4556,N_3454,N_3472);
xor U4557 (N_4557,N_3326,N_3338);
nor U4558 (N_4558,N_3251,N_3031);
and U4559 (N_4559,N_3138,N_3604);
or U4560 (N_4560,N_3659,N_3063);
nand U4561 (N_4561,N_3203,N_3291);
xor U4562 (N_4562,N_3723,N_3638);
and U4563 (N_4563,N_3280,N_3579);
or U4564 (N_4564,N_3498,N_3122);
and U4565 (N_4565,N_3213,N_3251);
and U4566 (N_4566,N_3459,N_3464);
nand U4567 (N_4567,N_3533,N_3392);
nor U4568 (N_4568,N_3642,N_3709);
nand U4569 (N_4569,N_3725,N_3199);
xnor U4570 (N_4570,N_3505,N_3236);
or U4571 (N_4571,N_3608,N_3641);
nor U4572 (N_4572,N_3704,N_3230);
or U4573 (N_4573,N_3712,N_3101);
xor U4574 (N_4574,N_3521,N_3598);
nor U4575 (N_4575,N_3659,N_3528);
or U4576 (N_4576,N_3763,N_3584);
or U4577 (N_4577,N_3228,N_3753);
xor U4578 (N_4578,N_3247,N_3075);
nor U4579 (N_4579,N_3771,N_3262);
nand U4580 (N_4580,N_3977,N_3849);
nand U4581 (N_4581,N_3772,N_3421);
nor U4582 (N_4582,N_3226,N_3369);
nor U4583 (N_4583,N_3584,N_3622);
nand U4584 (N_4584,N_3406,N_3757);
nand U4585 (N_4585,N_3129,N_3331);
or U4586 (N_4586,N_3611,N_3675);
nand U4587 (N_4587,N_3213,N_3527);
and U4588 (N_4588,N_3753,N_3204);
xor U4589 (N_4589,N_3288,N_3011);
nand U4590 (N_4590,N_3197,N_3050);
or U4591 (N_4591,N_3224,N_3777);
or U4592 (N_4592,N_3960,N_3737);
xnor U4593 (N_4593,N_3277,N_3370);
xor U4594 (N_4594,N_3259,N_3656);
and U4595 (N_4595,N_3014,N_3557);
and U4596 (N_4596,N_3221,N_3520);
or U4597 (N_4597,N_3319,N_3270);
nor U4598 (N_4598,N_3924,N_3348);
or U4599 (N_4599,N_3299,N_3083);
nand U4600 (N_4600,N_3368,N_3957);
nand U4601 (N_4601,N_3714,N_3823);
xnor U4602 (N_4602,N_3061,N_3756);
xor U4603 (N_4603,N_3338,N_3374);
nand U4604 (N_4604,N_3524,N_3220);
nand U4605 (N_4605,N_3791,N_3455);
nor U4606 (N_4606,N_3390,N_3784);
nor U4607 (N_4607,N_3293,N_3788);
or U4608 (N_4608,N_3077,N_3123);
nor U4609 (N_4609,N_3779,N_3237);
or U4610 (N_4610,N_3214,N_3295);
and U4611 (N_4611,N_3543,N_3204);
xnor U4612 (N_4612,N_3469,N_3010);
xor U4613 (N_4613,N_3529,N_3336);
xor U4614 (N_4614,N_3845,N_3775);
nand U4615 (N_4615,N_3415,N_3515);
nand U4616 (N_4616,N_3401,N_3988);
or U4617 (N_4617,N_3069,N_3724);
and U4618 (N_4618,N_3845,N_3715);
nand U4619 (N_4619,N_3431,N_3757);
or U4620 (N_4620,N_3947,N_3775);
nor U4621 (N_4621,N_3639,N_3274);
or U4622 (N_4622,N_3823,N_3347);
nand U4623 (N_4623,N_3487,N_3634);
nand U4624 (N_4624,N_3855,N_3221);
and U4625 (N_4625,N_3037,N_3263);
nor U4626 (N_4626,N_3622,N_3403);
nand U4627 (N_4627,N_3203,N_3866);
nand U4628 (N_4628,N_3117,N_3151);
or U4629 (N_4629,N_3499,N_3734);
or U4630 (N_4630,N_3150,N_3297);
nand U4631 (N_4631,N_3071,N_3907);
nand U4632 (N_4632,N_3270,N_3417);
nand U4633 (N_4633,N_3632,N_3518);
and U4634 (N_4634,N_3516,N_3456);
and U4635 (N_4635,N_3018,N_3636);
or U4636 (N_4636,N_3877,N_3787);
nand U4637 (N_4637,N_3063,N_3905);
and U4638 (N_4638,N_3877,N_3467);
nand U4639 (N_4639,N_3918,N_3721);
nor U4640 (N_4640,N_3945,N_3626);
or U4641 (N_4641,N_3220,N_3092);
nor U4642 (N_4642,N_3526,N_3237);
or U4643 (N_4643,N_3961,N_3638);
nand U4644 (N_4644,N_3053,N_3560);
xor U4645 (N_4645,N_3808,N_3812);
nand U4646 (N_4646,N_3160,N_3119);
or U4647 (N_4647,N_3936,N_3636);
or U4648 (N_4648,N_3505,N_3899);
nor U4649 (N_4649,N_3872,N_3202);
or U4650 (N_4650,N_3105,N_3795);
nand U4651 (N_4651,N_3887,N_3272);
or U4652 (N_4652,N_3445,N_3317);
and U4653 (N_4653,N_3902,N_3987);
or U4654 (N_4654,N_3142,N_3936);
nand U4655 (N_4655,N_3060,N_3514);
xor U4656 (N_4656,N_3071,N_3912);
nand U4657 (N_4657,N_3180,N_3354);
or U4658 (N_4658,N_3752,N_3466);
nand U4659 (N_4659,N_3296,N_3630);
nor U4660 (N_4660,N_3271,N_3043);
or U4661 (N_4661,N_3669,N_3428);
nor U4662 (N_4662,N_3800,N_3211);
xnor U4663 (N_4663,N_3500,N_3211);
nor U4664 (N_4664,N_3825,N_3281);
xor U4665 (N_4665,N_3555,N_3605);
and U4666 (N_4666,N_3357,N_3844);
xor U4667 (N_4667,N_3745,N_3929);
nand U4668 (N_4668,N_3851,N_3201);
xor U4669 (N_4669,N_3894,N_3029);
xor U4670 (N_4670,N_3858,N_3096);
nor U4671 (N_4671,N_3863,N_3328);
nand U4672 (N_4672,N_3227,N_3718);
and U4673 (N_4673,N_3357,N_3950);
or U4674 (N_4674,N_3851,N_3743);
nand U4675 (N_4675,N_3383,N_3236);
nor U4676 (N_4676,N_3169,N_3440);
and U4677 (N_4677,N_3030,N_3625);
xnor U4678 (N_4678,N_3307,N_3005);
or U4679 (N_4679,N_3652,N_3288);
nand U4680 (N_4680,N_3889,N_3844);
and U4681 (N_4681,N_3031,N_3784);
nand U4682 (N_4682,N_3468,N_3718);
or U4683 (N_4683,N_3861,N_3193);
and U4684 (N_4684,N_3726,N_3195);
nor U4685 (N_4685,N_3594,N_3610);
and U4686 (N_4686,N_3794,N_3091);
nor U4687 (N_4687,N_3741,N_3685);
and U4688 (N_4688,N_3672,N_3027);
nand U4689 (N_4689,N_3526,N_3891);
or U4690 (N_4690,N_3023,N_3510);
and U4691 (N_4691,N_3859,N_3986);
or U4692 (N_4692,N_3712,N_3775);
xor U4693 (N_4693,N_3578,N_3376);
xnor U4694 (N_4694,N_3907,N_3436);
or U4695 (N_4695,N_3459,N_3275);
nand U4696 (N_4696,N_3159,N_3624);
nor U4697 (N_4697,N_3929,N_3529);
nor U4698 (N_4698,N_3204,N_3927);
nand U4699 (N_4699,N_3635,N_3654);
or U4700 (N_4700,N_3970,N_3128);
xor U4701 (N_4701,N_3900,N_3295);
or U4702 (N_4702,N_3501,N_3460);
nand U4703 (N_4703,N_3179,N_3627);
nand U4704 (N_4704,N_3608,N_3384);
xnor U4705 (N_4705,N_3842,N_3679);
or U4706 (N_4706,N_3076,N_3656);
nor U4707 (N_4707,N_3449,N_3163);
and U4708 (N_4708,N_3431,N_3555);
or U4709 (N_4709,N_3254,N_3721);
nor U4710 (N_4710,N_3650,N_3126);
nand U4711 (N_4711,N_3637,N_3184);
nor U4712 (N_4712,N_3453,N_3722);
nor U4713 (N_4713,N_3157,N_3012);
and U4714 (N_4714,N_3795,N_3802);
xor U4715 (N_4715,N_3137,N_3007);
or U4716 (N_4716,N_3535,N_3184);
nand U4717 (N_4717,N_3177,N_3873);
nor U4718 (N_4718,N_3862,N_3055);
or U4719 (N_4719,N_3166,N_3077);
xor U4720 (N_4720,N_3451,N_3627);
xor U4721 (N_4721,N_3116,N_3669);
nor U4722 (N_4722,N_3082,N_3192);
and U4723 (N_4723,N_3188,N_3809);
or U4724 (N_4724,N_3403,N_3426);
nor U4725 (N_4725,N_3905,N_3792);
xor U4726 (N_4726,N_3046,N_3310);
nand U4727 (N_4727,N_3087,N_3809);
nor U4728 (N_4728,N_3908,N_3339);
nand U4729 (N_4729,N_3172,N_3746);
xnor U4730 (N_4730,N_3877,N_3435);
nor U4731 (N_4731,N_3289,N_3251);
nand U4732 (N_4732,N_3490,N_3605);
nand U4733 (N_4733,N_3204,N_3631);
nor U4734 (N_4734,N_3994,N_3822);
xor U4735 (N_4735,N_3898,N_3021);
nand U4736 (N_4736,N_3513,N_3743);
or U4737 (N_4737,N_3933,N_3418);
nand U4738 (N_4738,N_3085,N_3008);
nor U4739 (N_4739,N_3627,N_3791);
or U4740 (N_4740,N_3537,N_3627);
and U4741 (N_4741,N_3155,N_3048);
xnor U4742 (N_4742,N_3956,N_3084);
xnor U4743 (N_4743,N_3319,N_3404);
or U4744 (N_4744,N_3345,N_3815);
nor U4745 (N_4745,N_3508,N_3820);
xor U4746 (N_4746,N_3707,N_3083);
or U4747 (N_4747,N_3935,N_3216);
nand U4748 (N_4748,N_3796,N_3505);
nor U4749 (N_4749,N_3790,N_3203);
and U4750 (N_4750,N_3818,N_3412);
nor U4751 (N_4751,N_3946,N_3263);
nand U4752 (N_4752,N_3491,N_3728);
nor U4753 (N_4753,N_3621,N_3205);
and U4754 (N_4754,N_3614,N_3345);
or U4755 (N_4755,N_3612,N_3261);
nand U4756 (N_4756,N_3266,N_3177);
or U4757 (N_4757,N_3128,N_3042);
and U4758 (N_4758,N_3511,N_3423);
nor U4759 (N_4759,N_3654,N_3524);
nor U4760 (N_4760,N_3939,N_3194);
and U4761 (N_4761,N_3904,N_3855);
nand U4762 (N_4762,N_3565,N_3990);
and U4763 (N_4763,N_3044,N_3602);
xor U4764 (N_4764,N_3188,N_3421);
nand U4765 (N_4765,N_3267,N_3312);
nand U4766 (N_4766,N_3287,N_3524);
nand U4767 (N_4767,N_3758,N_3316);
or U4768 (N_4768,N_3374,N_3303);
xnor U4769 (N_4769,N_3401,N_3818);
xor U4770 (N_4770,N_3762,N_3249);
nor U4771 (N_4771,N_3476,N_3365);
xnor U4772 (N_4772,N_3150,N_3102);
xnor U4773 (N_4773,N_3603,N_3637);
or U4774 (N_4774,N_3874,N_3683);
nand U4775 (N_4775,N_3508,N_3873);
nand U4776 (N_4776,N_3547,N_3229);
or U4777 (N_4777,N_3171,N_3370);
nor U4778 (N_4778,N_3664,N_3082);
and U4779 (N_4779,N_3920,N_3566);
nor U4780 (N_4780,N_3383,N_3199);
and U4781 (N_4781,N_3372,N_3736);
xor U4782 (N_4782,N_3681,N_3255);
xor U4783 (N_4783,N_3934,N_3517);
and U4784 (N_4784,N_3668,N_3370);
and U4785 (N_4785,N_3980,N_3466);
xor U4786 (N_4786,N_3151,N_3747);
and U4787 (N_4787,N_3176,N_3576);
and U4788 (N_4788,N_3534,N_3225);
nor U4789 (N_4789,N_3460,N_3395);
xor U4790 (N_4790,N_3287,N_3000);
and U4791 (N_4791,N_3011,N_3545);
nor U4792 (N_4792,N_3991,N_3578);
xnor U4793 (N_4793,N_3636,N_3542);
nand U4794 (N_4794,N_3671,N_3301);
xnor U4795 (N_4795,N_3837,N_3592);
xnor U4796 (N_4796,N_3917,N_3111);
nor U4797 (N_4797,N_3042,N_3067);
nor U4798 (N_4798,N_3011,N_3686);
xnor U4799 (N_4799,N_3443,N_3199);
nor U4800 (N_4800,N_3658,N_3493);
xnor U4801 (N_4801,N_3191,N_3728);
nand U4802 (N_4802,N_3291,N_3429);
xor U4803 (N_4803,N_3412,N_3657);
nand U4804 (N_4804,N_3614,N_3908);
xnor U4805 (N_4805,N_3104,N_3470);
nor U4806 (N_4806,N_3765,N_3800);
or U4807 (N_4807,N_3325,N_3475);
and U4808 (N_4808,N_3010,N_3666);
nand U4809 (N_4809,N_3779,N_3927);
xnor U4810 (N_4810,N_3708,N_3301);
nor U4811 (N_4811,N_3629,N_3082);
xnor U4812 (N_4812,N_3798,N_3732);
xor U4813 (N_4813,N_3052,N_3506);
or U4814 (N_4814,N_3879,N_3253);
nand U4815 (N_4815,N_3267,N_3039);
nand U4816 (N_4816,N_3705,N_3292);
nand U4817 (N_4817,N_3050,N_3984);
or U4818 (N_4818,N_3485,N_3605);
and U4819 (N_4819,N_3686,N_3303);
nor U4820 (N_4820,N_3640,N_3918);
xnor U4821 (N_4821,N_3246,N_3313);
and U4822 (N_4822,N_3855,N_3076);
nor U4823 (N_4823,N_3582,N_3905);
nor U4824 (N_4824,N_3394,N_3586);
nor U4825 (N_4825,N_3311,N_3761);
nor U4826 (N_4826,N_3874,N_3592);
or U4827 (N_4827,N_3598,N_3314);
nand U4828 (N_4828,N_3746,N_3259);
xnor U4829 (N_4829,N_3542,N_3053);
nor U4830 (N_4830,N_3603,N_3540);
xor U4831 (N_4831,N_3566,N_3271);
nor U4832 (N_4832,N_3166,N_3097);
or U4833 (N_4833,N_3700,N_3858);
or U4834 (N_4834,N_3962,N_3633);
or U4835 (N_4835,N_3809,N_3406);
nor U4836 (N_4836,N_3028,N_3537);
or U4837 (N_4837,N_3016,N_3486);
nor U4838 (N_4838,N_3061,N_3297);
xor U4839 (N_4839,N_3490,N_3302);
or U4840 (N_4840,N_3877,N_3155);
nand U4841 (N_4841,N_3516,N_3043);
nand U4842 (N_4842,N_3891,N_3191);
nor U4843 (N_4843,N_3276,N_3074);
and U4844 (N_4844,N_3899,N_3044);
nor U4845 (N_4845,N_3458,N_3161);
nand U4846 (N_4846,N_3968,N_3667);
and U4847 (N_4847,N_3177,N_3430);
nand U4848 (N_4848,N_3980,N_3519);
nand U4849 (N_4849,N_3779,N_3708);
nand U4850 (N_4850,N_3927,N_3893);
and U4851 (N_4851,N_3260,N_3492);
and U4852 (N_4852,N_3631,N_3352);
or U4853 (N_4853,N_3099,N_3996);
nand U4854 (N_4854,N_3456,N_3268);
and U4855 (N_4855,N_3909,N_3175);
nor U4856 (N_4856,N_3835,N_3858);
xnor U4857 (N_4857,N_3578,N_3256);
nor U4858 (N_4858,N_3361,N_3532);
and U4859 (N_4859,N_3183,N_3988);
or U4860 (N_4860,N_3368,N_3074);
nor U4861 (N_4861,N_3909,N_3257);
nand U4862 (N_4862,N_3609,N_3500);
xnor U4863 (N_4863,N_3944,N_3760);
and U4864 (N_4864,N_3859,N_3957);
and U4865 (N_4865,N_3355,N_3817);
xor U4866 (N_4866,N_3438,N_3972);
nor U4867 (N_4867,N_3656,N_3202);
nand U4868 (N_4868,N_3236,N_3729);
nor U4869 (N_4869,N_3698,N_3671);
and U4870 (N_4870,N_3074,N_3648);
and U4871 (N_4871,N_3616,N_3659);
or U4872 (N_4872,N_3453,N_3632);
xnor U4873 (N_4873,N_3258,N_3635);
xnor U4874 (N_4874,N_3577,N_3763);
xnor U4875 (N_4875,N_3438,N_3268);
xnor U4876 (N_4876,N_3692,N_3799);
xor U4877 (N_4877,N_3258,N_3684);
nand U4878 (N_4878,N_3341,N_3332);
or U4879 (N_4879,N_3594,N_3284);
or U4880 (N_4880,N_3235,N_3340);
xnor U4881 (N_4881,N_3340,N_3585);
nor U4882 (N_4882,N_3958,N_3015);
or U4883 (N_4883,N_3475,N_3172);
nand U4884 (N_4884,N_3037,N_3497);
or U4885 (N_4885,N_3308,N_3791);
nor U4886 (N_4886,N_3145,N_3038);
nor U4887 (N_4887,N_3521,N_3740);
or U4888 (N_4888,N_3769,N_3952);
or U4889 (N_4889,N_3579,N_3139);
or U4890 (N_4890,N_3099,N_3268);
and U4891 (N_4891,N_3380,N_3141);
or U4892 (N_4892,N_3619,N_3674);
nor U4893 (N_4893,N_3851,N_3624);
nand U4894 (N_4894,N_3789,N_3865);
and U4895 (N_4895,N_3756,N_3128);
and U4896 (N_4896,N_3413,N_3654);
xor U4897 (N_4897,N_3916,N_3689);
and U4898 (N_4898,N_3648,N_3036);
and U4899 (N_4899,N_3196,N_3562);
nand U4900 (N_4900,N_3361,N_3224);
or U4901 (N_4901,N_3975,N_3279);
nor U4902 (N_4902,N_3740,N_3040);
and U4903 (N_4903,N_3109,N_3973);
or U4904 (N_4904,N_3055,N_3793);
nand U4905 (N_4905,N_3686,N_3281);
or U4906 (N_4906,N_3264,N_3939);
nand U4907 (N_4907,N_3715,N_3956);
xor U4908 (N_4908,N_3930,N_3685);
and U4909 (N_4909,N_3484,N_3009);
nor U4910 (N_4910,N_3020,N_3347);
xor U4911 (N_4911,N_3963,N_3967);
xnor U4912 (N_4912,N_3872,N_3601);
nand U4913 (N_4913,N_3945,N_3630);
xnor U4914 (N_4914,N_3784,N_3956);
xnor U4915 (N_4915,N_3554,N_3300);
nand U4916 (N_4916,N_3783,N_3185);
or U4917 (N_4917,N_3750,N_3263);
and U4918 (N_4918,N_3998,N_3565);
xnor U4919 (N_4919,N_3949,N_3511);
and U4920 (N_4920,N_3829,N_3070);
nor U4921 (N_4921,N_3924,N_3047);
and U4922 (N_4922,N_3301,N_3107);
nand U4923 (N_4923,N_3008,N_3644);
or U4924 (N_4924,N_3758,N_3703);
or U4925 (N_4925,N_3788,N_3013);
nand U4926 (N_4926,N_3292,N_3217);
nand U4927 (N_4927,N_3803,N_3805);
nor U4928 (N_4928,N_3744,N_3850);
and U4929 (N_4929,N_3275,N_3387);
xor U4930 (N_4930,N_3284,N_3812);
xnor U4931 (N_4931,N_3604,N_3361);
xnor U4932 (N_4932,N_3344,N_3714);
nand U4933 (N_4933,N_3676,N_3359);
or U4934 (N_4934,N_3153,N_3087);
nand U4935 (N_4935,N_3014,N_3328);
nor U4936 (N_4936,N_3918,N_3100);
and U4937 (N_4937,N_3492,N_3495);
nor U4938 (N_4938,N_3431,N_3052);
xnor U4939 (N_4939,N_3301,N_3526);
xnor U4940 (N_4940,N_3670,N_3434);
and U4941 (N_4941,N_3522,N_3778);
xor U4942 (N_4942,N_3333,N_3465);
and U4943 (N_4943,N_3577,N_3562);
nor U4944 (N_4944,N_3965,N_3375);
nor U4945 (N_4945,N_3257,N_3197);
and U4946 (N_4946,N_3970,N_3492);
xor U4947 (N_4947,N_3083,N_3945);
nand U4948 (N_4948,N_3768,N_3338);
or U4949 (N_4949,N_3892,N_3984);
nor U4950 (N_4950,N_3247,N_3150);
nand U4951 (N_4951,N_3810,N_3455);
nor U4952 (N_4952,N_3068,N_3798);
and U4953 (N_4953,N_3672,N_3840);
xor U4954 (N_4954,N_3713,N_3555);
nor U4955 (N_4955,N_3735,N_3540);
or U4956 (N_4956,N_3690,N_3854);
nor U4957 (N_4957,N_3959,N_3069);
nand U4958 (N_4958,N_3417,N_3787);
and U4959 (N_4959,N_3459,N_3332);
or U4960 (N_4960,N_3557,N_3367);
or U4961 (N_4961,N_3682,N_3206);
or U4962 (N_4962,N_3404,N_3323);
nand U4963 (N_4963,N_3149,N_3799);
xor U4964 (N_4964,N_3073,N_3021);
or U4965 (N_4965,N_3390,N_3648);
nor U4966 (N_4966,N_3007,N_3650);
or U4967 (N_4967,N_3460,N_3290);
nor U4968 (N_4968,N_3529,N_3136);
nand U4969 (N_4969,N_3921,N_3493);
nand U4970 (N_4970,N_3515,N_3354);
or U4971 (N_4971,N_3460,N_3920);
nand U4972 (N_4972,N_3908,N_3403);
xnor U4973 (N_4973,N_3960,N_3669);
and U4974 (N_4974,N_3303,N_3685);
or U4975 (N_4975,N_3683,N_3073);
and U4976 (N_4976,N_3455,N_3057);
or U4977 (N_4977,N_3474,N_3085);
nor U4978 (N_4978,N_3151,N_3578);
and U4979 (N_4979,N_3125,N_3958);
nor U4980 (N_4980,N_3284,N_3418);
nand U4981 (N_4981,N_3435,N_3626);
nand U4982 (N_4982,N_3667,N_3156);
and U4983 (N_4983,N_3900,N_3844);
xor U4984 (N_4984,N_3064,N_3029);
nor U4985 (N_4985,N_3283,N_3186);
nand U4986 (N_4986,N_3135,N_3933);
xor U4987 (N_4987,N_3593,N_3603);
nor U4988 (N_4988,N_3861,N_3541);
xnor U4989 (N_4989,N_3718,N_3914);
nor U4990 (N_4990,N_3723,N_3564);
or U4991 (N_4991,N_3756,N_3504);
nor U4992 (N_4992,N_3467,N_3235);
xnor U4993 (N_4993,N_3777,N_3830);
xnor U4994 (N_4994,N_3513,N_3168);
xor U4995 (N_4995,N_3477,N_3517);
nand U4996 (N_4996,N_3447,N_3727);
nor U4997 (N_4997,N_3528,N_3187);
nand U4998 (N_4998,N_3825,N_3988);
nand U4999 (N_4999,N_3041,N_3816);
nand U5000 (N_5000,N_4906,N_4675);
nor U5001 (N_5001,N_4192,N_4188);
xor U5002 (N_5002,N_4376,N_4184);
nor U5003 (N_5003,N_4018,N_4146);
nor U5004 (N_5004,N_4263,N_4652);
or U5005 (N_5005,N_4265,N_4239);
nand U5006 (N_5006,N_4278,N_4824);
xnor U5007 (N_5007,N_4819,N_4346);
nand U5008 (N_5008,N_4934,N_4875);
or U5009 (N_5009,N_4455,N_4913);
nor U5010 (N_5010,N_4161,N_4432);
nand U5011 (N_5011,N_4220,N_4201);
or U5012 (N_5012,N_4320,N_4958);
nor U5013 (N_5013,N_4366,N_4830);
and U5014 (N_5014,N_4488,N_4310);
nor U5015 (N_5015,N_4673,N_4690);
nand U5016 (N_5016,N_4294,N_4525);
nor U5017 (N_5017,N_4223,N_4345);
xor U5018 (N_5018,N_4617,N_4340);
xnor U5019 (N_5019,N_4999,N_4597);
xor U5020 (N_5020,N_4742,N_4465);
or U5021 (N_5021,N_4833,N_4554);
or U5022 (N_5022,N_4419,N_4250);
and U5023 (N_5023,N_4307,N_4347);
nand U5024 (N_5024,N_4799,N_4952);
xor U5025 (N_5025,N_4963,N_4701);
or U5026 (N_5026,N_4474,N_4193);
or U5027 (N_5027,N_4247,N_4771);
nand U5028 (N_5028,N_4500,N_4748);
or U5029 (N_5029,N_4152,N_4684);
nand U5030 (N_5030,N_4632,N_4905);
or U5031 (N_5031,N_4526,N_4887);
nor U5032 (N_5032,N_4976,N_4922);
and U5033 (N_5033,N_4497,N_4890);
nand U5034 (N_5034,N_4537,N_4168);
xnor U5035 (N_5035,N_4202,N_4761);
or U5036 (N_5036,N_4815,N_4016);
xor U5037 (N_5037,N_4739,N_4687);
nor U5038 (N_5038,N_4475,N_4923);
nor U5039 (N_5039,N_4928,N_4048);
xnor U5040 (N_5040,N_4249,N_4206);
nor U5041 (N_5041,N_4494,N_4831);
nor U5042 (N_5042,N_4164,N_4495);
and U5043 (N_5043,N_4400,N_4492);
and U5044 (N_5044,N_4795,N_4702);
and U5045 (N_5045,N_4343,N_4522);
nand U5046 (N_5046,N_4626,N_4036);
and U5047 (N_5047,N_4172,N_4292);
nor U5048 (N_5048,N_4079,N_4352);
or U5049 (N_5049,N_4736,N_4924);
or U5050 (N_5050,N_4588,N_4792);
or U5051 (N_5051,N_4829,N_4023);
or U5052 (N_5052,N_4000,N_4843);
nor U5053 (N_5053,N_4769,N_4452);
nand U5054 (N_5054,N_4274,N_4169);
nor U5055 (N_5055,N_4431,N_4893);
and U5056 (N_5056,N_4364,N_4966);
xnor U5057 (N_5057,N_4938,N_4695);
nor U5058 (N_5058,N_4037,N_4723);
and U5059 (N_5059,N_4101,N_4804);
and U5060 (N_5060,N_4859,N_4003);
and U5061 (N_5061,N_4167,N_4926);
or U5062 (N_5062,N_4296,N_4106);
nor U5063 (N_5063,N_4911,N_4425);
and U5064 (N_5064,N_4219,N_4153);
nor U5065 (N_5065,N_4987,N_4468);
and U5066 (N_5066,N_4543,N_4803);
nand U5067 (N_5067,N_4147,N_4403);
and U5068 (N_5068,N_4094,N_4752);
xor U5069 (N_5069,N_4162,N_4787);
xor U5070 (N_5070,N_4888,N_4845);
xor U5071 (N_5071,N_4199,N_4629);
nand U5072 (N_5072,N_4145,N_4342);
or U5073 (N_5073,N_4257,N_4204);
xnor U5074 (N_5074,N_4714,N_4892);
and U5075 (N_5075,N_4160,N_4104);
and U5076 (N_5076,N_4559,N_4885);
nor U5077 (N_5077,N_4844,N_4649);
nor U5078 (N_5078,N_4024,N_4808);
nor U5079 (N_5079,N_4625,N_4996);
xnor U5080 (N_5080,N_4594,N_4897);
or U5081 (N_5081,N_4654,N_4754);
and U5082 (N_5082,N_4740,N_4117);
or U5083 (N_5083,N_4020,N_4076);
or U5084 (N_5084,N_4679,N_4322);
and U5085 (N_5085,N_4074,N_4213);
and U5086 (N_5086,N_4997,N_4384);
nor U5087 (N_5087,N_4744,N_4004);
nor U5088 (N_5088,N_4643,N_4084);
nor U5089 (N_5089,N_4354,N_4461);
xor U5090 (N_5090,N_4667,N_4760);
nand U5091 (N_5091,N_4705,N_4470);
or U5092 (N_5092,N_4648,N_4448);
or U5093 (N_5093,N_4991,N_4937);
nand U5094 (N_5094,N_4584,N_4668);
nand U5095 (N_5095,N_4399,N_4772);
or U5096 (N_5096,N_4089,N_4699);
and U5097 (N_5097,N_4434,N_4176);
nor U5098 (N_5098,N_4300,N_4511);
nand U5099 (N_5099,N_4598,N_4010);
nor U5100 (N_5100,N_4225,N_4585);
or U5101 (N_5101,N_4590,N_4515);
nand U5102 (N_5102,N_4931,N_4916);
nor U5103 (N_5103,N_4917,N_4103);
xor U5104 (N_5104,N_4421,N_4118);
or U5105 (N_5105,N_4582,N_4130);
and U5106 (N_5106,N_4569,N_4719);
xor U5107 (N_5107,N_4878,N_4535);
and U5108 (N_5108,N_4043,N_4170);
and U5109 (N_5109,N_4990,N_4866);
and U5110 (N_5110,N_4194,N_4746);
or U5111 (N_5111,N_4077,N_4908);
and U5112 (N_5112,N_4373,N_4639);
nand U5113 (N_5113,N_4258,N_4339);
nand U5114 (N_5114,N_4853,N_4809);
and U5115 (N_5115,N_4344,N_4027);
or U5116 (N_5116,N_4717,N_4062);
nor U5117 (N_5117,N_4960,N_4589);
nand U5118 (N_5118,N_4472,N_4676);
nor U5119 (N_5119,N_4596,N_4747);
or U5120 (N_5120,N_4788,N_4513);
xor U5121 (N_5121,N_4724,N_4180);
nand U5122 (N_5122,N_4238,N_4396);
and U5123 (N_5123,N_4127,N_4749);
and U5124 (N_5124,N_4564,N_4682);
and U5125 (N_5125,N_4880,N_4750);
and U5126 (N_5126,N_4031,N_4816);
nor U5127 (N_5127,N_4388,N_4694);
xor U5128 (N_5128,N_4441,N_4323);
or U5129 (N_5129,N_4367,N_4698);
or U5130 (N_5130,N_4650,N_4557);
and U5131 (N_5131,N_4454,N_4600);
xnor U5132 (N_5132,N_4614,N_4841);
and U5133 (N_5133,N_4186,N_4802);
and U5134 (N_5134,N_4435,N_4707);
nand U5135 (N_5135,N_4041,N_4418);
nor U5136 (N_5136,N_4979,N_4381);
nand U5137 (N_5137,N_4150,N_4575);
nor U5138 (N_5138,N_4409,N_4969);
and U5139 (N_5139,N_4456,N_4026);
and U5140 (N_5140,N_4657,N_4826);
nor U5141 (N_5141,N_4112,N_4471);
nand U5142 (N_5142,N_4759,N_4858);
or U5143 (N_5143,N_4414,N_4581);
and U5144 (N_5144,N_4411,N_4510);
and U5145 (N_5145,N_4097,N_4974);
xor U5146 (N_5146,N_4734,N_4688);
nor U5147 (N_5147,N_4610,N_4189);
xor U5148 (N_5148,N_4408,N_4218);
xnor U5149 (N_5149,N_4067,N_4357);
and U5150 (N_5150,N_4116,N_4828);
nor U5151 (N_5151,N_4523,N_4786);
and U5152 (N_5152,N_4375,N_4224);
nor U5153 (N_5153,N_4449,N_4889);
nor U5154 (N_5154,N_4896,N_4704);
or U5155 (N_5155,N_4727,N_4132);
nand U5156 (N_5156,N_4835,N_4646);
nor U5157 (N_5157,N_4546,N_4313);
and U5158 (N_5158,N_4134,N_4302);
and U5159 (N_5159,N_4528,N_4797);
or U5160 (N_5160,N_4601,N_4603);
and U5161 (N_5161,N_4539,N_4361);
nor U5162 (N_5162,N_4262,N_4315);
xnor U5163 (N_5163,N_4463,N_4940);
nand U5164 (N_5164,N_4064,N_4426);
nor U5165 (N_5165,N_4834,N_4267);
nor U5166 (N_5166,N_4832,N_4618);
nor U5167 (N_5167,N_4195,N_4593);
nor U5168 (N_5168,N_4281,N_4233);
nand U5169 (N_5169,N_4653,N_4563);
nor U5170 (N_5170,N_4166,N_4818);
xnor U5171 (N_5171,N_4131,N_4827);
and U5172 (N_5172,N_4964,N_4236);
nand U5173 (N_5173,N_4254,N_4847);
nor U5174 (N_5174,N_4430,N_4241);
and U5175 (N_5175,N_4521,N_4856);
and U5176 (N_5176,N_4288,N_4123);
nand U5177 (N_5177,N_4159,N_4336);
nand U5178 (N_5178,N_4686,N_4033);
nand U5179 (N_5179,N_4825,N_4333);
and U5180 (N_5180,N_4807,N_4737);
nand U5181 (N_5181,N_4226,N_4640);
nand U5182 (N_5182,N_4385,N_4237);
nor U5183 (N_5183,N_4209,N_4013);
xnor U5184 (N_5184,N_4731,N_4605);
nand U5185 (N_5185,N_4273,N_4993);
nor U5186 (N_5186,N_4630,N_4138);
or U5187 (N_5187,N_4945,N_4946);
nand U5188 (N_5188,N_4052,N_4898);
or U5189 (N_5189,N_4527,N_4370);
or U5190 (N_5190,N_4360,N_4284);
xor U5191 (N_5191,N_4139,N_4785);
nand U5192 (N_5192,N_4277,N_4395);
nand U5193 (N_5193,N_4493,N_4351);
nor U5194 (N_5194,N_4072,N_4711);
or U5195 (N_5195,N_4729,N_4082);
nand U5196 (N_5196,N_4136,N_4613);
xnor U5197 (N_5197,N_4607,N_4245);
xor U5198 (N_5198,N_4285,N_4536);
or U5199 (N_5199,N_4604,N_4297);
nor U5200 (N_5200,N_4087,N_4457);
nor U5201 (N_5201,N_4222,N_4390);
or U5202 (N_5202,N_4895,N_4114);
nand U5203 (N_5203,N_4460,N_4524);
nand U5204 (N_5204,N_4155,N_4846);
nor U5205 (N_5205,N_4633,N_4207);
and U5206 (N_5206,N_4002,N_4022);
nand U5207 (N_5207,N_4291,N_4369);
or U5208 (N_5208,N_4619,N_4365);
nand U5209 (N_5209,N_4276,N_4915);
nor U5210 (N_5210,N_4720,N_4205);
nor U5211 (N_5211,N_4040,N_4635);
nor U5212 (N_5212,N_4019,N_4975);
nand U5213 (N_5213,N_4781,N_4417);
nor U5214 (N_5214,N_4075,N_4133);
and U5215 (N_5215,N_4349,N_4382);
nor U5216 (N_5216,N_4623,N_4995);
and U5217 (N_5217,N_4756,N_4548);
xnor U5218 (N_5218,N_4110,N_4732);
xnor U5219 (N_5219,N_4374,N_4156);
xnor U5220 (N_5220,N_4534,N_4058);
and U5221 (N_5221,N_4469,N_4083);
nand U5222 (N_5222,N_4986,N_4341);
nand U5223 (N_5223,N_4726,N_4801);
nor U5224 (N_5224,N_4124,N_4459);
nand U5225 (N_5225,N_4392,N_4095);
nand U5226 (N_5226,N_4587,N_4311);
xor U5227 (N_5227,N_4337,N_4871);
nand U5228 (N_5228,N_4044,N_4666);
and U5229 (N_5229,N_4105,N_4243);
or U5230 (N_5230,N_4259,N_4091);
or U5231 (N_5231,N_4778,N_4948);
and U5232 (N_5232,N_4935,N_4674);
nand U5233 (N_5233,N_4289,N_4255);
nand U5234 (N_5234,N_4063,N_4178);
nand U5235 (N_5235,N_4586,N_4822);
nor U5236 (N_5236,N_4071,N_4864);
xor U5237 (N_5237,N_4198,N_4485);
nand U5238 (N_5238,N_4715,N_4009);
nand U5239 (N_5239,N_4085,N_4932);
nand U5240 (N_5240,N_4440,N_4907);
xor U5241 (N_5241,N_4232,N_4394);
xor U5242 (N_5242,N_4942,N_4122);
nor U5243 (N_5243,N_4627,N_4268);
nand U5244 (N_5244,N_4933,N_4775);
nand U5245 (N_5245,N_4054,N_4305);
nand U5246 (N_5246,N_4516,N_4529);
xnor U5247 (N_5247,N_4899,N_4661);
nand U5248 (N_5248,N_4280,N_4253);
nand U5249 (N_5249,N_4006,N_4580);
and U5250 (N_5250,N_4068,N_4069);
and U5251 (N_5251,N_4573,N_4174);
and U5252 (N_5252,N_4279,N_4282);
xnor U5253 (N_5253,N_4450,N_4185);
nand U5254 (N_5254,N_4894,N_4725);
xnor U5255 (N_5255,N_4439,N_4275);
or U5256 (N_5256,N_4025,N_4216);
xnor U5257 (N_5257,N_4318,N_4356);
nand U5258 (N_5258,N_4883,N_4608);
xor U5259 (N_5259,N_4314,N_4696);
or U5260 (N_5260,N_4854,N_4109);
nand U5261 (N_5261,N_4776,N_4697);
and U5262 (N_5262,N_4599,N_4212);
nor U5263 (N_5263,N_4316,N_4955);
and U5264 (N_5264,N_4865,N_4609);
nand U5265 (N_5265,N_4055,N_4716);
nor U5266 (N_5266,N_4304,N_4936);
nand U5267 (N_5267,N_4283,N_4927);
and U5268 (N_5268,N_4959,N_4738);
nand U5269 (N_5269,N_4709,N_4480);
nor U5270 (N_5270,N_4484,N_4944);
nand U5271 (N_5271,N_4148,N_4820);
or U5272 (N_5272,N_4879,N_4857);
or U5273 (N_5273,N_4780,N_4165);
nand U5274 (N_5274,N_4217,N_4957);
nor U5275 (N_5275,N_4228,N_4287);
xor U5276 (N_5276,N_4397,N_4290);
or U5277 (N_5277,N_4479,N_4230);
nor U5278 (N_5278,N_4863,N_4355);
nand U5279 (N_5279,N_4299,N_4773);
nand U5280 (N_5280,N_4177,N_4505);
xor U5281 (N_5281,N_4246,N_4542);
nor U5282 (N_5282,N_4900,N_4532);
nor U5283 (N_5283,N_4047,N_4514);
nand U5284 (N_5284,N_4200,N_4644);
and U5285 (N_5285,N_4001,N_4681);
nand U5286 (N_5286,N_4503,N_4757);
and U5287 (N_5287,N_4141,N_4840);
nor U5288 (N_5288,N_4850,N_4547);
nand U5289 (N_5289,N_4540,N_4665);
nand U5290 (N_5290,N_4743,N_4173);
and U5291 (N_5291,N_4446,N_4487);
and U5292 (N_5292,N_4359,N_4327);
nor U5293 (N_5293,N_4121,N_4606);
nor U5294 (N_5294,N_4545,N_4501);
nand U5295 (N_5295,N_4651,N_4579);
or U5296 (N_5296,N_4142,N_4994);
nor U5297 (N_5297,N_4507,N_4777);
nand U5298 (N_5298,N_4647,N_4144);
nor U5299 (N_5299,N_4904,N_4903);
and U5300 (N_5300,N_4229,N_4555);
and U5301 (N_5301,N_4443,N_4140);
nand U5302 (N_5302,N_4353,N_4591);
xnor U5303 (N_5303,N_4961,N_4332);
nand U5304 (N_5304,N_4008,N_4753);
xnor U5305 (N_5305,N_4358,N_4458);
nor U5306 (N_5306,N_4252,N_4572);
xor U5307 (N_5307,N_4240,N_4518);
xnor U5308 (N_5308,N_4096,N_4508);
nor U5309 (N_5309,N_4386,N_4324);
nor U5310 (N_5310,N_4046,N_4902);
xnor U5311 (N_5311,N_4837,N_4870);
nand U5312 (N_5312,N_4549,N_4424);
nand U5313 (N_5313,N_4793,N_4442);
nor U5314 (N_5314,N_4641,N_4473);
nand U5315 (N_5315,N_4334,N_4881);
nor U5316 (N_5316,N_4663,N_4973);
and U5317 (N_5317,N_4143,N_4416);
xor U5318 (N_5318,N_4982,N_4005);
nand U5319 (N_5319,N_4306,N_4574);
and U5320 (N_5320,N_4483,N_4852);
nand U5321 (N_5321,N_4842,N_4486);
and U5322 (N_5322,N_4693,N_4891);
and U5323 (N_5323,N_4377,N_4860);
nor U5324 (N_5324,N_4691,N_4677);
or U5325 (N_5325,N_4912,N_4298);
xnor U5326 (N_5326,N_4766,N_4774);
nor U5327 (N_5327,N_4953,N_4135);
or U5328 (N_5328,N_4444,N_4102);
and U5329 (N_5329,N_4631,N_4919);
nor U5330 (N_5330,N_4989,N_4700);
nand U5331 (N_5331,N_4462,N_4406);
xnor U5332 (N_5332,N_4851,N_4078);
and U5333 (N_5333,N_4560,N_4558);
and U5334 (N_5334,N_4293,N_4798);
or U5335 (N_5335,N_4645,N_4490);
or U5336 (N_5336,N_4423,N_4149);
nand U5337 (N_5337,N_4628,N_4197);
nor U5338 (N_5338,N_4556,N_4983);
nor U5339 (N_5339,N_4562,N_4295);
xor U5340 (N_5340,N_4190,N_4791);
or U5341 (N_5341,N_4119,N_4678);
or U5342 (N_5342,N_4489,N_4956);
nor U5343 (N_5343,N_4595,N_4427);
and U5344 (N_5344,N_4925,N_4874);
xnor U5345 (N_5345,N_4429,N_4271);
nand U5346 (N_5346,N_4393,N_4583);
nand U5347 (N_5347,N_4042,N_4502);
nor U5348 (N_5348,N_4751,N_4466);
nand U5349 (N_5349,N_4971,N_4420);
nor U5350 (N_5350,N_4034,N_4261);
xnor U5351 (N_5351,N_4477,N_4007);
and U5352 (N_5352,N_4531,N_4918);
xor U5353 (N_5353,N_4806,N_4762);
xnor U5354 (N_5354,N_4437,N_4115);
and U5355 (N_5355,N_4301,N_4764);
and U5356 (N_5356,N_4093,N_4038);
nor U5357 (N_5357,N_4553,N_4796);
xnor U5358 (N_5358,N_4615,N_4208);
nor U5359 (N_5359,N_4943,N_4992);
nor U5360 (N_5360,N_4810,N_4445);
or U5361 (N_5361,N_4967,N_4972);
and U5362 (N_5362,N_4685,N_4482);
and U5363 (N_5363,N_4624,N_4566);
nor U5364 (N_5364,N_4158,N_4498);
xor U5365 (N_5365,N_4947,N_4378);
or U5366 (N_5366,N_4057,N_4988);
and U5367 (N_5367,N_4476,N_4187);
xnor U5368 (N_5368,N_4861,N_4519);
nand U5369 (N_5369,N_4520,N_4950);
and U5370 (N_5370,N_4453,N_4789);
xor U5371 (N_5371,N_4721,N_4869);
nand U5372 (N_5372,N_4049,N_4552);
and U5373 (N_5373,N_4438,N_4642);
xor U5374 (N_5374,N_4380,N_4921);
nand U5375 (N_5375,N_4984,N_4413);
or U5376 (N_5376,N_4151,N_4985);
nor U5377 (N_5377,N_4794,N_4855);
or U5378 (N_5378,N_4568,N_4015);
nor U5379 (N_5379,N_4128,N_4447);
nand U5380 (N_5380,N_4326,N_4836);
nor U5381 (N_5381,N_4065,N_4372);
xnor U5382 (N_5382,N_4538,N_4672);
nor U5383 (N_5383,N_4066,N_4722);
and U5384 (N_5384,N_4713,N_4061);
nor U5385 (N_5385,N_4658,N_4730);
and U5386 (N_5386,N_4839,N_4512);
nor U5387 (N_5387,N_4876,N_4081);
xor U5388 (N_5388,N_4692,N_4090);
xnor U5389 (N_5389,N_4108,N_4478);
nor U5390 (N_5390,N_4602,N_4312);
and U5391 (N_5391,N_4264,N_4350);
or U5392 (N_5392,N_4708,N_4060);
or U5393 (N_5393,N_4028,N_4882);
xor U5394 (N_5394,N_4886,N_4570);
xor U5395 (N_5395,N_4611,N_4561);
xor U5396 (N_5396,N_4733,N_4422);
xor U5397 (N_5397,N_4612,N_4286);
nor U5398 (N_5398,N_4059,N_4578);
or U5399 (N_5399,N_4506,N_4571);
nor U5400 (N_5400,N_4379,N_4029);
nand U5401 (N_5401,N_4317,N_4662);
nor U5402 (N_5402,N_4873,N_4428);
or U5403 (N_5403,N_4032,N_4660);
or U5404 (N_5404,N_4765,N_4211);
and U5405 (N_5405,N_4391,N_4655);
nor U5406 (N_5406,N_4741,N_4182);
nor U5407 (N_5407,N_4929,N_4868);
nand U5408 (N_5408,N_4544,N_4227);
and U5409 (N_5409,N_4621,N_4039);
xnor U5410 (N_5410,N_4183,N_4683);
or U5411 (N_5411,N_4415,N_4813);
and U5412 (N_5412,N_4260,N_4407);
xor U5413 (N_5413,N_4949,N_4954);
nor U5414 (N_5414,N_4451,N_4035);
nand U5415 (N_5415,N_4970,N_4405);
nand U5416 (N_5416,N_4745,N_4812);
nand U5417 (N_5417,N_4877,N_4763);
or U5418 (N_5418,N_4331,N_4070);
nor U5419 (N_5419,N_4017,N_4387);
and U5420 (N_5420,N_4755,N_4410);
nand U5421 (N_5421,N_4080,N_4541);
nor U5422 (N_5422,N_4266,N_4179);
and U5423 (N_5423,N_4129,N_4251);
xnor U5424 (N_5424,N_4113,N_4620);
nand U5425 (N_5425,N_4436,N_4530);
nor U5426 (N_5426,N_4163,N_4256);
and U5427 (N_5427,N_4120,N_4638);
nor U5428 (N_5428,N_4767,N_4965);
and U5429 (N_5429,N_4242,N_4056);
xor U5430 (N_5430,N_4303,N_4328);
xor U5431 (N_5431,N_4014,N_4718);
nand U5432 (N_5432,N_4782,N_4664);
nor U5433 (N_5433,N_4977,N_4951);
or U5434 (N_5434,N_4805,N_4823);
or U5435 (N_5435,N_4867,N_4616);
xor U5436 (N_5436,N_4884,N_4330);
nor U5437 (N_5437,N_4800,N_4551);
xor U5438 (N_5438,N_4814,N_4728);
or U5439 (N_5439,N_4499,N_4401);
nor U5440 (N_5440,N_4231,N_4030);
xor U5441 (N_5441,N_4669,N_4784);
nor U5442 (N_5442,N_4978,N_4053);
and U5443 (N_5443,N_4221,N_4768);
and U5444 (N_5444,N_4710,N_4248);
nand U5445 (N_5445,N_4939,N_4758);
or U5446 (N_5446,N_4215,N_4636);
nor U5447 (N_5447,N_4706,N_4550);
xnor U5448 (N_5448,N_4175,N_4504);
or U5449 (N_5449,N_4404,N_4021);
xor U5450 (N_5450,N_4998,N_4481);
nor U5451 (N_5451,N_4203,N_4348);
nand U5452 (N_5452,N_4099,N_4517);
xor U5453 (N_5453,N_4637,N_4098);
and U5454 (N_5454,N_4329,N_4092);
or U5455 (N_5455,N_4930,N_4671);
xor U5456 (N_5456,N_4191,N_4171);
or U5457 (N_5457,N_4234,N_4088);
nor U5458 (N_5458,N_4086,N_4308);
or U5459 (N_5459,N_4689,N_4412);
nor U5460 (N_5460,N_4111,N_4073);
and U5461 (N_5461,N_4901,N_4680);
or U5462 (N_5462,N_4214,N_4849);
nor U5463 (N_5463,N_4567,N_4045);
xor U5464 (N_5464,N_4011,N_4981);
xor U5465 (N_5465,N_4670,N_4196);
nor U5466 (N_5466,N_4272,N_4910);
nand U5467 (N_5467,N_4270,N_4433);
and U5468 (N_5468,N_4811,N_4656);
nand U5469 (N_5469,N_4577,N_4783);
xnor U5470 (N_5470,N_4389,N_4565);
or U5471 (N_5471,N_4137,N_4770);
or U5472 (N_5472,N_4634,N_4980);
or U5473 (N_5473,N_4319,N_4712);
or U5474 (N_5474,N_4848,N_4496);
xor U5475 (N_5475,N_4210,N_4909);
and U5476 (N_5476,N_4467,N_4622);
and U5477 (N_5477,N_4309,N_4321);
nor U5478 (N_5478,N_4659,N_4464);
xnor U5479 (N_5479,N_4533,N_4872);
nor U5480 (N_5480,N_4051,N_4371);
or U5481 (N_5481,N_4914,N_4368);
xor U5482 (N_5482,N_4154,N_4968);
nor U5483 (N_5483,N_4335,N_4100);
or U5484 (N_5484,N_4235,N_4269);
xor U5485 (N_5485,N_4838,N_4817);
xor U5486 (N_5486,N_4592,N_4050);
or U5487 (N_5487,N_4491,N_4920);
or U5488 (N_5488,N_4107,N_4790);
nor U5489 (N_5489,N_4157,N_4779);
or U5490 (N_5490,N_4402,N_4821);
or U5491 (N_5491,N_4362,N_4941);
and U5492 (N_5492,N_4338,N_4012);
or U5493 (N_5493,N_4862,N_4181);
and U5494 (N_5494,N_4125,N_4126);
xor U5495 (N_5495,N_4735,N_4962);
or U5496 (N_5496,N_4398,N_4576);
xnor U5497 (N_5497,N_4383,N_4363);
and U5498 (N_5498,N_4244,N_4325);
or U5499 (N_5499,N_4703,N_4509);
nor U5500 (N_5500,N_4052,N_4817);
nor U5501 (N_5501,N_4705,N_4906);
nand U5502 (N_5502,N_4441,N_4643);
or U5503 (N_5503,N_4411,N_4577);
nand U5504 (N_5504,N_4689,N_4776);
or U5505 (N_5505,N_4660,N_4669);
and U5506 (N_5506,N_4674,N_4005);
xor U5507 (N_5507,N_4201,N_4697);
and U5508 (N_5508,N_4901,N_4089);
xor U5509 (N_5509,N_4713,N_4505);
or U5510 (N_5510,N_4332,N_4882);
and U5511 (N_5511,N_4462,N_4784);
xnor U5512 (N_5512,N_4792,N_4278);
nand U5513 (N_5513,N_4080,N_4545);
and U5514 (N_5514,N_4961,N_4864);
or U5515 (N_5515,N_4602,N_4937);
or U5516 (N_5516,N_4175,N_4611);
and U5517 (N_5517,N_4079,N_4878);
and U5518 (N_5518,N_4589,N_4679);
xnor U5519 (N_5519,N_4394,N_4544);
and U5520 (N_5520,N_4467,N_4073);
nor U5521 (N_5521,N_4097,N_4114);
nand U5522 (N_5522,N_4135,N_4171);
or U5523 (N_5523,N_4850,N_4355);
nor U5524 (N_5524,N_4221,N_4782);
nand U5525 (N_5525,N_4619,N_4658);
and U5526 (N_5526,N_4602,N_4729);
and U5527 (N_5527,N_4644,N_4078);
xor U5528 (N_5528,N_4331,N_4415);
and U5529 (N_5529,N_4041,N_4405);
or U5530 (N_5530,N_4670,N_4454);
xor U5531 (N_5531,N_4896,N_4605);
nand U5532 (N_5532,N_4683,N_4132);
xor U5533 (N_5533,N_4661,N_4110);
or U5534 (N_5534,N_4218,N_4286);
nor U5535 (N_5535,N_4550,N_4695);
nor U5536 (N_5536,N_4176,N_4631);
nor U5537 (N_5537,N_4468,N_4132);
nand U5538 (N_5538,N_4823,N_4912);
and U5539 (N_5539,N_4133,N_4339);
nand U5540 (N_5540,N_4248,N_4949);
xor U5541 (N_5541,N_4369,N_4523);
xnor U5542 (N_5542,N_4130,N_4407);
or U5543 (N_5543,N_4950,N_4041);
nor U5544 (N_5544,N_4487,N_4253);
or U5545 (N_5545,N_4161,N_4254);
or U5546 (N_5546,N_4522,N_4502);
nand U5547 (N_5547,N_4177,N_4467);
nor U5548 (N_5548,N_4881,N_4421);
nand U5549 (N_5549,N_4078,N_4033);
or U5550 (N_5550,N_4758,N_4424);
nand U5551 (N_5551,N_4497,N_4251);
or U5552 (N_5552,N_4007,N_4456);
and U5553 (N_5553,N_4474,N_4034);
xnor U5554 (N_5554,N_4377,N_4811);
nand U5555 (N_5555,N_4168,N_4158);
nand U5556 (N_5556,N_4939,N_4788);
nand U5557 (N_5557,N_4217,N_4912);
or U5558 (N_5558,N_4699,N_4297);
and U5559 (N_5559,N_4672,N_4783);
or U5560 (N_5560,N_4437,N_4121);
nor U5561 (N_5561,N_4480,N_4213);
or U5562 (N_5562,N_4753,N_4449);
nor U5563 (N_5563,N_4251,N_4085);
and U5564 (N_5564,N_4032,N_4333);
and U5565 (N_5565,N_4721,N_4353);
nand U5566 (N_5566,N_4947,N_4846);
or U5567 (N_5567,N_4289,N_4356);
nor U5568 (N_5568,N_4313,N_4783);
nand U5569 (N_5569,N_4164,N_4544);
and U5570 (N_5570,N_4570,N_4696);
xor U5571 (N_5571,N_4211,N_4935);
nand U5572 (N_5572,N_4809,N_4921);
nor U5573 (N_5573,N_4329,N_4290);
xor U5574 (N_5574,N_4266,N_4347);
and U5575 (N_5575,N_4016,N_4397);
xor U5576 (N_5576,N_4201,N_4591);
nand U5577 (N_5577,N_4984,N_4235);
or U5578 (N_5578,N_4008,N_4604);
xor U5579 (N_5579,N_4124,N_4050);
and U5580 (N_5580,N_4459,N_4374);
xnor U5581 (N_5581,N_4898,N_4599);
and U5582 (N_5582,N_4699,N_4487);
or U5583 (N_5583,N_4244,N_4256);
or U5584 (N_5584,N_4148,N_4718);
nand U5585 (N_5585,N_4756,N_4067);
or U5586 (N_5586,N_4011,N_4073);
xor U5587 (N_5587,N_4997,N_4075);
or U5588 (N_5588,N_4011,N_4053);
and U5589 (N_5589,N_4350,N_4685);
xnor U5590 (N_5590,N_4562,N_4888);
and U5591 (N_5591,N_4701,N_4069);
and U5592 (N_5592,N_4716,N_4518);
xnor U5593 (N_5593,N_4434,N_4790);
or U5594 (N_5594,N_4916,N_4433);
and U5595 (N_5595,N_4825,N_4935);
or U5596 (N_5596,N_4101,N_4246);
xnor U5597 (N_5597,N_4653,N_4398);
nor U5598 (N_5598,N_4071,N_4244);
and U5599 (N_5599,N_4091,N_4345);
nand U5600 (N_5600,N_4983,N_4318);
nor U5601 (N_5601,N_4848,N_4747);
nor U5602 (N_5602,N_4626,N_4709);
nor U5603 (N_5603,N_4450,N_4508);
and U5604 (N_5604,N_4503,N_4282);
or U5605 (N_5605,N_4075,N_4406);
xnor U5606 (N_5606,N_4760,N_4542);
xnor U5607 (N_5607,N_4650,N_4481);
or U5608 (N_5608,N_4795,N_4988);
or U5609 (N_5609,N_4862,N_4555);
or U5610 (N_5610,N_4834,N_4982);
and U5611 (N_5611,N_4998,N_4621);
xnor U5612 (N_5612,N_4568,N_4993);
nor U5613 (N_5613,N_4169,N_4809);
nor U5614 (N_5614,N_4862,N_4468);
nor U5615 (N_5615,N_4295,N_4195);
nor U5616 (N_5616,N_4165,N_4460);
nand U5617 (N_5617,N_4684,N_4800);
nor U5618 (N_5618,N_4475,N_4454);
nand U5619 (N_5619,N_4975,N_4314);
or U5620 (N_5620,N_4257,N_4448);
and U5621 (N_5621,N_4554,N_4195);
xor U5622 (N_5622,N_4491,N_4826);
and U5623 (N_5623,N_4209,N_4482);
xnor U5624 (N_5624,N_4450,N_4303);
nor U5625 (N_5625,N_4256,N_4632);
and U5626 (N_5626,N_4764,N_4324);
or U5627 (N_5627,N_4008,N_4434);
or U5628 (N_5628,N_4654,N_4427);
nor U5629 (N_5629,N_4007,N_4576);
and U5630 (N_5630,N_4596,N_4410);
xor U5631 (N_5631,N_4095,N_4896);
and U5632 (N_5632,N_4438,N_4887);
nand U5633 (N_5633,N_4231,N_4936);
and U5634 (N_5634,N_4728,N_4919);
xnor U5635 (N_5635,N_4215,N_4127);
and U5636 (N_5636,N_4711,N_4871);
xnor U5637 (N_5637,N_4705,N_4571);
or U5638 (N_5638,N_4486,N_4516);
nor U5639 (N_5639,N_4265,N_4016);
or U5640 (N_5640,N_4127,N_4446);
or U5641 (N_5641,N_4654,N_4421);
nor U5642 (N_5642,N_4263,N_4053);
nor U5643 (N_5643,N_4506,N_4257);
nor U5644 (N_5644,N_4489,N_4342);
nor U5645 (N_5645,N_4744,N_4073);
and U5646 (N_5646,N_4715,N_4622);
and U5647 (N_5647,N_4853,N_4072);
nand U5648 (N_5648,N_4042,N_4469);
nand U5649 (N_5649,N_4974,N_4481);
or U5650 (N_5650,N_4310,N_4083);
or U5651 (N_5651,N_4479,N_4905);
nand U5652 (N_5652,N_4671,N_4344);
nor U5653 (N_5653,N_4564,N_4188);
xnor U5654 (N_5654,N_4639,N_4967);
and U5655 (N_5655,N_4504,N_4636);
nand U5656 (N_5656,N_4491,N_4991);
nor U5657 (N_5657,N_4435,N_4816);
and U5658 (N_5658,N_4286,N_4310);
xnor U5659 (N_5659,N_4964,N_4272);
nor U5660 (N_5660,N_4789,N_4454);
or U5661 (N_5661,N_4040,N_4470);
nand U5662 (N_5662,N_4174,N_4508);
and U5663 (N_5663,N_4971,N_4498);
xor U5664 (N_5664,N_4659,N_4994);
nand U5665 (N_5665,N_4456,N_4226);
nand U5666 (N_5666,N_4162,N_4568);
nor U5667 (N_5667,N_4219,N_4957);
and U5668 (N_5668,N_4074,N_4401);
nand U5669 (N_5669,N_4322,N_4781);
or U5670 (N_5670,N_4615,N_4701);
and U5671 (N_5671,N_4628,N_4481);
nor U5672 (N_5672,N_4838,N_4371);
xor U5673 (N_5673,N_4736,N_4669);
nor U5674 (N_5674,N_4272,N_4622);
and U5675 (N_5675,N_4020,N_4120);
or U5676 (N_5676,N_4472,N_4263);
nand U5677 (N_5677,N_4512,N_4170);
and U5678 (N_5678,N_4255,N_4829);
xnor U5679 (N_5679,N_4887,N_4497);
nor U5680 (N_5680,N_4715,N_4360);
nor U5681 (N_5681,N_4313,N_4285);
and U5682 (N_5682,N_4337,N_4854);
nor U5683 (N_5683,N_4914,N_4482);
and U5684 (N_5684,N_4115,N_4818);
and U5685 (N_5685,N_4649,N_4218);
xor U5686 (N_5686,N_4501,N_4924);
xor U5687 (N_5687,N_4222,N_4173);
nand U5688 (N_5688,N_4848,N_4905);
nand U5689 (N_5689,N_4434,N_4652);
nor U5690 (N_5690,N_4994,N_4407);
nor U5691 (N_5691,N_4103,N_4527);
nand U5692 (N_5692,N_4139,N_4017);
xor U5693 (N_5693,N_4063,N_4282);
nand U5694 (N_5694,N_4873,N_4869);
nand U5695 (N_5695,N_4437,N_4701);
nor U5696 (N_5696,N_4585,N_4917);
nand U5697 (N_5697,N_4579,N_4630);
xnor U5698 (N_5698,N_4344,N_4611);
or U5699 (N_5699,N_4568,N_4609);
xnor U5700 (N_5700,N_4882,N_4462);
and U5701 (N_5701,N_4329,N_4922);
nor U5702 (N_5702,N_4154,N_4387);
nor U5703 (N_5703,N_4759,N_4651);
and U5704 (N_5704,N_4480,N_4602);
xor U5705 (N_5705,N_4686,N_4911);
nor U5706 (N_5706,N_4154,N_4422);
and U5707 (N_5707,N_4983,N_4432);
or U5708 (N_5708,N_4367,N_4298);
nor U5709 (N_5709,N_4733,N_4047);
xor U5710 (N_5710,N_4422,N_4696);
nor U5711 (N_5711,N_4768,N_4924);
or U5712 (N_5712,N_4093,N_4918);
xor U5713 (N_5713,N_4456,N_4811);
xnor U5714 (N_5714,N_4841,N_4503);
or U5715 (N_5715,N_4202,N_4426);
or U5716 (N_5716,N_4428,N_4487);
xnor U5717 (N_5717,N_4059,N_4277);
nor U5718 (N_5718,N_4724,N_4702);
and U5719 (N_5719,N_4821,N_4456);
and U5720 (N_5720,N_4450,N_4883);
nor U5721 (N_5721,N_4003,N_4953);
nand U5722 (N_5722,N_4049,N_4897);
nand U5723 (N_5723,N_4588,N_4318);
or U5724 (N_5724,N_4006,N_4961);
nand U5725 (N_5725,N_4005,N_4523);
or U5726 (N_5726,N_4136,N_4875);
xnor U5727 (N_5727,N_4718,N_4380);
and U5728 (N_5728,N_4256,N_4515);
xnor U5729 (N_5729,N_4544,N_4993);
and U5730 (N_5730,N_4972,N_4992);
nor U5731 (N_5731,N_4495,N_4431);
nand U5732 (N_5732,N_4845,N_4079);
nor U5733 (N_5733,N_4573,N_4959);
and U5734 (N_5734,N_4067,N_4576);
nor U5735 (N_5735,N_4778,N_4722);
xor U5736 (N_5736,N_4758,N_4204);
nor U5737 (N_5737,N_4725,N_4602);
xnor U5738 (N_5738,N_4527,N_4634);
and U5739 (N_5739,N_4625,N_4023);
nor U5740 (N_5740,N_4264,N_4098);
nor U5741 (N_5741,N_4734,N_4135);
nor U5742 (N_5742,N_4334,N_4668);
or U5743 (N_5743,N_4077,N_4051);
nor U5744 (N_5744,N_4923,N_4306);
nand U5745 (N_5745,N_4285,N_4627);
nand U5746 (N_5746,N_4014,N_4249);
nor U5747 (N_5747,N_4616,N_4427);
or U5748 (N_5748,N_4567,N_4445);
nor U5749 (N_5749,N_4371,N_4407);
nand U5750 (N_5750,N_4266,N_4891);
or U5751 (N_5751,N_4409,N_4106);
and U5752 (N_5752,N_4179,N_4226);
nand U5753 (N_5753,N_4413,N_4638);
xnor U5754 (N_5754,N_4589,N_4306);
nor U5755 (N_5755,N_4755,N_4221);
nor U5756 (N_5756,N_4694,N_4114);
or U5757 (N_5757,N_4084,N_4896);
nor U5758 (N_5758,N_4058,N_4517);
and U5759 (N_5759,N_4499,N_4797);
nand U5760 (N_5760,N_4355,N_4823);
or U5761 (N_5761,N_4315,N_4182);
nor U5762 (N_5762,N_4302,N_4655);
xnor U5763 (N_5763,N_4963,N_4125);
and U5764 (N_5764,N_4226,N_4888);
nor U5765 (N_5765,N_4181,N_4644);
xnor U5766 (N_5766,N_4075,N_4638);
xor U5767 (N_5767,N_4586,N_4642);
and U5768 (N_5768,N_4583,N_4407);
nor U5769 (N_5769,N_4952,N_4348);
or U5770 (N_5770,N_4917,N_4726);
xor U5771 (N_5771,N_4789,N_4246);
and U5772 (N_5772,N_4598,N_4413);
and U5773 (N_5773,N_4466,N_4345);
or U5774 (N_5774,N_4356,N_4278);
xnor U5775 (N_5775,N_4173,N_4105);
xnor U5776 (N_5776,N_4287,N_4652);
nand U5777 (N_5777,N_4487,N_4664);
nand U5778 (N_5778,N_4146,N_4944);
nor U5779 (N_5779,N_4181,N_4165);
nor U5780 (N_5780,N_4799,N_4168);
or U5781 (N_5781,N_4895,N_4230);
nand U5782 (N_5782,N_4502,N_4801);
and U5783 (N_5783,N_4980,N_4286);
nor U5784 (N_5784,N_4023,N_4262);
and U5785 (N_5785,N_4040,N_4846);
or U5786 (N_5786,N_4281,N_4056);
or U5787 (N_5787,N_4018,N_4847);
nor U5788 (N_5788,N_4499,N_4672);
and U5789 (N_5789,N_4874,N_4792);
nor U5790 (N_5790,N_4447,N_4001);
nor U5791 (N_5791,N_4824,N_4968);
nand U5792 (N_5792,N_4099,N_4259);
and U5793 (N_5793,N_4551,N_4814);
or U5794 (N_5794,N_4248,N_4450);
and U5795 (N_5795,N_4284,N_4504);
xor U5796 (N_5796,N_4945,N_4870);
nand U5797 (N_5797,N_4742,N_4579);
and U5798 (N_5798,N_4736,N_4705);
or U5799 (N_5799,N_4511,N_4430);
nor U5800 (N_5800,N_4434,N_4755);
xnor U5801 (N_5801,N_4462,N_4997);
nor U5802 (N_5802,N_4526,N_4125);
xor U5803 (N_5803,N_4036,N_4552);
and U5804 (N_5804,N_4234,N_4029);
or U5805 (N_5805,N_4783,N_4275);
or U5806 (N_5806,N_4511,N_4128);
or U5807 (N_5807,N_4289,N_4816);
and U5808 (N_5808,N_4844,N_4431);
xor U5809 (N_5809,N_4381,N_4501);
xnor U5810 (N_5810,N_4382,N_4213);
or U5811 (N_5811,N_4424,N_4068);
or U5812 (N_5812,N_4040,N_4219);
nor U5813 (N_5813,N_4027,N_4959);
nand U5814 (N_5814,N_4717,N_4266);
nor U5815 (N_5815,N_4175,N_4336);
xor U5816 (N_5816,N_4715,N_4445);
xnor U5817 (N_5817,N_4489,N_4265);
or U5818 (N_5818,N_4985,N_4816);
nand U5819 (N_5819,N_4653,N_4771);
or U5820 (N_5820,N_4046,N_4675);
or U5821 (N_5821,N_4273,N_4452);
nor U5822 (N_5822,N_4654,N_4593);
or U5823 (N_5823,N_4481,N_4879);
or U5824 (N_5824,N_4030,N_4203);
nor U5825 (N_5825,N_4142,N_4524);
or U5826 (N_5826,N_4661,N_4319);
nand U5827 (N_5827,N_4898,N_4252);
or U5828 (N_5828,N_4228,N_4639);
xor U5829 (N_5829,N_4039,N_4156);
or U5830 (N_5830,N_4084,N_4212);
xor U5831 (N_5831,N_4454,N_4056);
nand U5832 (N_5832,N_4649,N_4377);
nand U5833 (N_5833,N_4904,N_4428);
and U5834 (N_5834,N_4726,N_4258);
and U5835 (N_5835,N_4441,N_4660);
and U5836 (N_5836,N_4592,N_4600);
and U5837 (N_5837,N_4409,N_4079);
nor U5838 (N_5838,N_4736,N_4310);
nand U5839 (N_5839,N_4199,N_4379);
xnor U5840 (N_5840,N_4201,N_4889);
xnor U5841 (N_5841,N_4320,N_4982);
and U5842 (N_5842,N_4631,N_4332);
and U5843 (N_5843,N_4075,N_4152);
nand U5844 (N_5844,N_4374,N_4829);
nor U5845 (N_5845,N_4462,N_4310);
nand U5846 (N_5846,N_4419,N_4201);
or U5847 (N_5847,N_4879,N_4147);
or U5848 (N_5848,N_4068,N_4899);
nand U5849 (N_5849,N_4771,N_4382);
and U5850 (N_5850,N_4159,N_4905);
nor U5851 (N_5851,N_4310,N_4937);
xnor U5852 (N_5852,N_4766,N_4443);
nand U5853 (N_5853,N_4842,N_4520);
nor U5854 (N_5854,N_4607,N_4390);
nor U5855 (N_5855,N_4158,N_4655);
xnor U5856 (N_5856,N_4893,N_4755);
nor U5857 (N_5857,N_4847,N_4737);
and U5858 (N_5858,N_4758,N_4293);
nand U5859 (N_5859,N_4660,N_4903);
nor U5860 (N_5860,N_4913,N_4853);
nand U5861 (N_5861,N_4615,N_4484);
or U5862 (N_5862,N_4548,N_4281);
and U5863 (N_5863,N_4964,N_4433);
or U5864 (N_5864,N_4940,N_4603);
nand U5865 (N_5865,N_4111,N_4406);
xnor U5866 (N_5866,N_4194,N_4748);
and U5867 (N_5867,N_4352,N_4579);
or U5868 (N_5868,N_4436,N_4434);
nor U5869 (N_5869,N_4892,N_4190);
nor U5870 (N_5870,N_4237,N_4812);
nor U5871 (N_5871,N_4642,N_4722);
and U5872 (N_5872,N_4612,N_4968);
nor U5873 (N_5873,N_4942,N_4012);
or U5874 (N_5874,N_4171,N_4972);
xnor U5875 (N_5875,N_4175,N_4793);
or U5876 (N_5876,N_4102,N_4193);
or U5877 (N_5877,N_4058,N_4648);
nor U5878 (N_5878,N_4234,N_4020);
xnor U5879 (N_5879,N_4031,N_4860);
nand U5880 (N_5880,N_4923,N_4876);
xor U5881 (N_5881,N_4056,N_4970);
xor U5882 (N_5882,N_4598,N_4145);
or U5883 (N_5883,N_4648,N_4101);
and U5884 (N_5884,N_4307,N_4206);
and U5885 (N_5885,N_4951,N_4202);
nand U5886 (N_5886,N_4338,N_4685);
or U5887 (N_5887,N_4386,N_4853);
nor U5888 (N_5888,N_4239,N_4242);
nor U5889 (N_5889,N_4641,N_4357);
and U5890 (N_5890,N_4599,N_4124);
nor U5891 (N_5891,N_4241,N_4164);
and U5892 (N_5892,N_4583,N_4867);
or U5893 (N_5893,N_4952,N_4379);
xnor U5894 (N_5894,N_4560,N_4349);
or U5895 (N_5895,N_4710,N_4923);
nand U5896 (N_5896,N_4548,N_4481);
and U5897 (N_5897,N_4385,N_4595);
and U5898 (N_5898,N_4425,N_4134);
xor U5899 (N_5899,N_4691,N_4074);
xor U5900 (N_5900,N_4634,N_4108);
nand U5901 (N_5901,N_4892,N_4111);
and U5902 (N_5902,N_4452,N_4409);
and U5903 (N_5903,N_4164,N_4905);
nor U5904 (N_5904,N_4093,N_4278);
and U5905 (N_5905,N_4342,N_4944);
xor U5906 (N_5906,N_4931,N_4292);
or U5907 (N_5907,N_4306,N_4460);
or U5908 (N_5908,N_4018,N_4401);
xor U5909 (N_5909,N_4440,N_4077);
nand U5910 (N_5910,N_4381,N_4874);
nand U5911 (N_5911,N_4445,N_4015);
nor U5912 (N_5912,N_4523,N_4935);
xnor U5913 (N_5913,N_4211,N_4200);
or U5914 (N_5914,N_4467,N_4708);
nor U5915 (N_5915,N_4283,N_4114);
xor U5916 (N_5916,N_4019,N_4030);
nor U5917 (N_5917,N_4793,N_4453);
xor U5918 (N_5918,N_4208,N_4629);
nand U5919 (N_5919,N_4828,N_4553);
xnor U5920 (N_5920,N_4256,N_4355);
and U5921 (N_5921,N_4604,N_4570);
or U5922 (N_5922,N_4726,N_4866);
and U5923 (N_5923,N_4228,N_4968);
xor U5924 (N_5924,N_4809,N_4305);
and U5925 (N_5925,N_4198,N_4089);
xnor U5926 (N_5926,N_4166,N_4397);
nor U5927 (N_5927,N_4854,N_4174);
xor U5928 (N_5928,N_4546,N_4308);
or U5929 (N_5929,N_4703,N_4916);
or U5930 (N_5930,N_4426,N_4920);
or U5931 (N_5931,N_4365,N_4499);
nand U5932 (N_5932,N_4475,N_4215);
xnor U5933 (N_5933,N_4561,N_4905);
and U5934 (N_5934,N_4050,N_4852);
xnor U5935 (N_5935,N_4244,N_4026);
or U5936 (N_5936,N_4092,N_4164);
xnor U5937 (N_5937,N_4222,N_4324);
or U5938 (N_5938,N_4947,N_4731);
or U5939 (N_5939,N_4955,N_4709);
xnor U5940 (N_5940,N_4266,N_4138);
nand U5941 (N_5941,N_4979,N_4690);
or U5942 (N_5942,N_4392,N_4288);
xnor U5943 (N_5943,N_4761,N_4907);
or U5944 (N_5944,N_4093,N_4578);
and U5945 (N_5945,N_4469,N_4773);
nor U5946 (N_5946,N_4429,N_4000);
nor U5947 (N_5947,N_4190,N_4405);
xnor U5948 (N_5948,N_4412,N_4224);
and U5949 (N_5949,N_4281,N_4024);
or U5950 (N_5950,N_4540,N_4580);
and U5951 (N_5951,N_4062,N_4872);
nand U5952 (N_5952,N_4002,N_4211);
or U5953 (N_5953,N_4411,N_4871);
or U5954 (N_5954,N_4049,N_4615);
xnor U5955 (N_5955,N_4467,N_4319);
nand U5956 (N_5956,N_4937,N_4066);
nor U5957 (N_5957,N_4464,N_4603);
xor U5958 (N_5958,N_4200,N_4577);
and U5959 (N_5959,N_4416,N_4581);
nor U5960 (N_5960,N_4778,N_4852);
or U5961 (N_5961,N_4726,N_4709);
and U5962 (N_5962,N_4293,N_4985);
and U5963 (N_5963,N_4199,N_4424);
xor U5964 (N_5964,N_4752,N_4277);
nand U5965 (N_5965,N_4192,N_4458);
and U5966 (N_5966,N_4735,N_4399);
and U5967 (N_5967,N_4126,N_4769);
xor U5968 (N_5968,N_4860,N_4841);
or U5969 (N_5969,N_4919,N_4271);
xnor U5970 (N_5970,N_4949,N_4186);
nand U5971 (N_5971,N_4175,N_4217);
nor U5972 (N_5972,N_4577,N_4268);
nand U5973 (N_5973,N_4188,N_4624);
nor U5974 (N_5974,N_4158,N_4636);
and U5975 (N_5975,N_4523,N_4987);
or U5976 (N_5976,N_4957,N_4372);
nand U5977 (N_5977,N_4848,N_4588);
xor U5978 (N_5978,N_4586,N_4242);
nand U5979 (N_5979,N_4133,N_4313);
nor U5980 (N_5980,N_4155,N_4902);
and U5981 (N_5981,N_4525,N_4052);
nand U5982 (N_5982,N_4089,N_4835);
or U5983 (N_5983,N_4839,N_4604);
or U5984 (N_5984,N_4795,N_4061);
or U5985 (N_5985,N_4391,N_4275);
nor U5986 (N_5986,N_4058,N_4684);
or U5987 (N_5987,N_4298,N_4160);
nor U5988 (N_5988,N_4286,N_4535);
and U5989 (N_5989,N_4282,N_4491);
xnor U5990 (N_5990,N_4702,N_4851);
nor U5991 (N_5991,N_4916,N_4334);
xor U5992 (N_5992,N_4778,N_4025);
nor U5993 (N_5993,N_4252,N_4294);
and U5994 (N_5994,N_4139,N_4315);
or U5995 (N_5995,N_4596,N_4528);
xor U5996 (N_5996,N_4432,N_4103);
nor U5997 (N_5997,N_4703,N_4348);
nand U5998 (N_5998,N_4287,N_4800);
and U5999 (N_5999,N_4970,N_4291);
nor U6000 (N_6000,N_5155,N_5115);
and U6001 (N_6001,N_5995,N_5837);
or U6002 (N_6002,N_5522,N_5693);
and U6003 (N_6003,N_5930,N_5603);
nand U6004 (N_6004,N_5337,N_5910);
xor U6005 (N_6005,N_5034,N_5542);
and U6006 (N_6006,N_5183,N_5209);
nor U6007 (N_6007,N_5913,N_5415);
and U6008 (N_6008,N_5564,N_5560);
nand U6009 (N_6009,N_5315,N_5336);
and U6010 (N_6010,N_5375,N_5140);
nand U6011 (N_6011,N_5187,N_5486);
nand U6012 (N_6012,N_5577,N_5214);
or U6013 (N_6013,N_5865,N_5885);
nand U6014 (N_6014,N_5591,N_5710);
or U6015 (N_6015,N_5765,N_5749);
and U6016 (N_6016,N_5733,N_5616);
and U6017 (N_6017,N_5556,N_5005);
or U6018 (N_6018,N_5354,N_5648);
nand U6019 (N_6019,N_5017,N_5117);
nor U6020 (N_6020,N_5088,N_5418);
xor U6021 (N_6021,N_5386,N_5543);
or U6022 (N_6022,N_5359,N_5960);
and U6023 (N_6023,N_5978,N_5135);
or U6024 (N_6024,N_5043,N_5816);
or U6025 (N_6025,N_5179,N_5176);
or U6026 (N_6026,N_5771,N_5655);
and U6027 (N_6027,N_5219,N_5470);
and U6028 (N_6028,N_5847,N_5841);
and U6029 (N_6029,N_5658,N_5364);
nor U6030 (N_6030,N_5672,N_5300);
nand U6031 (N_6031,N_5356,N_5881);
nand U6032 (N_6032,N_5783,N_5138);
or U6033 (N_6033,N_5035,N_5168);
or U6034 (N_6034,N_5487,N_5391);
or U6035 (N_6035,N_5262,N_5961);
and U6036 (N_6036,N_5645,N_5157);
nor U6037 (N_6037,N_5149,N_5498);
and U6038 (N_6038,N_5854,N_5875);
and U6039 (N_6039,N_5372,N_5795);
xor U6040 (N_6040,N_5633,N_5849);
and U6041 (N_6041,N_5943,N_5549);
and U6042 (N_6042,N_5212,N_5036);
or U6043 (N_6043,N_5946,N_5481);
xor U6044 (N_6044,N_5734,N_5191);
nor U6045 (N_6045,N_5442,N_5095);
or U6046 (N_6046,N_5263,N_5936);
nand U6047 (N_6047,N_5096,N_5724);
nor U6048 (N_6048,N_5067,N_5644);
xnor U6049 (N_6049,N_5351,N_5144);
and U6050 (N_6050,N_5388,N_5220);
or U6051 (N_6051,N_5215,N_5305);
nand U6052 (N_6052,N_5124,N_5150);
nand U6053 (N_6053,N_5868,N_5864);
or U6054 (N_6054,N_5285,N_5694);
and U6055 (N_6055,N_5980,N_5905);
or U6056 (N_6056,N_5696,N_5573);
and U6057 (N_6057,N_5147,N_5712);
xnor U6058 (N_6058,N_5713,N_5226);
nor U6059 (N_6059,N_5477,N_5353);
nand U6060 (N_6060,N_5731,N_5678);
and U6061 (N_6061,N_5866,N_5079);
nor U6062 (N_6062,N_5082,N_5892);
nor U6063 (N_6063,N_5075,N_5662);
and U6064 (N_6064,N_5950,N_5965);
and U6065 (N_6065,N_5118,N_5202);
xor U6066 (N_6066,N_5076,N_5654);
and U6067 (N_6067,N_5130,N_5248);
nand U6068 (N_6068,N_5538,N_5106);
and U6069 (N_6069,N_5039,N_5152);
and U6070 (N_6070,N_5921,N_5751);
or U6071 (N_6071,N_5829,N_5363);
or U6072 (N_6072,N_5396,N_5318);
or U6073 (N_6073,N_5283,N_5730);
nor U6074 (N_6074,N_5899,N_5265);
xor U6075 (N_6075,N_5066,N_5196);
and U6076 (N_6076,N_5527,N_5022);
and U6077 (N_6077,N_5873,N_5981);
and U6078 (N_6078,N_5843,N_5643);
nand U6079 (N_6079,N_5876,N_5906);
and U6080 (N_6080,N_5113,N_5797);
or U6081 (N_6081,N_5977,N_5764);
xnor U6082 (N_6082,N_5735,N_5234);
and U6083 (N_6083,N_5755,N_5680);
and U6084 (N_6084,N_5621,N_5988);
and U6085 (N_6085,N_5878,N_5100);
and U6086 (N_6086,N_5282,N_5446);
xor U6087 (N_6087,N_5193,N_5695);
nand U6088 (N_6088,N_5178,N_5330);
nand U6089 (N_6089,N_5170,N_5613);
nor U6090 (N_6090,N_5935,N_5275);
and U6091 (N_6091,N_5671,N_5623);
xnor U6092 (N_6092,N_5939,N_5790);
xor U6093 (N_6093,N_5244,N_5456);
or U6094 (N_6094,N_5473,N_5929);
or U6095 (N_6095,N_5334,N_5483);
or U6096 (N_6096,N_5582,N_5227);
and U6097 (N_6097,N_5862,N_5000);
and U6098 (N_6098,N_5041,N_5801);
nor U6099 (N_6099,N_5412,N_5016);
and U6100 (N_6100,N_5125,N_5008);
xor U6101 (N_6101,N_5387,N_5989);
and U6102 (N_6102,N_5600,N_5224);
nand U6103 (N_6103,N_5894,N_5833);
nor U6104 (N_6104,N_5649,N_5681);
and U6105 (N_6105,N_5421,N_5010);
and U6106 (N_6106,N_5116,N_5120);
xnor U6107 (N_6107,N_5101,N_5539);
nor U6108 (N_6108,N_5126,N_5347);
and U6109 (N_6109,N_5907,N_5314);
xnor U6110 (N_6110,N_5682,N_5871);
and U6111 (N_6111,N_5601,N_5964);
nor U6112 (N_6112,N_5758,N_5465);
and U6113 (N_6113,N_5333,N_5172);
or U6114 (N_6114,N_5518,N_5690);
nor U6115 (N_6115,N_5235,N_5799);
nand U6116 (N_6116,N_5842,N_5812);
xor U6117 (N_6117,N_5872,N_5493);
and U6118 (N_6118,N_5617,N_5018);
and U6119 (N_6119,N_5427,N_5380);
nor U6120 (N_6120,N_5312,N_5225);
xor U6121 (N_6121,N_5827,N_5177);
or U6122 (N_6122,N_5970,N_5851);
nand U6123 (N_6123,N_5944,N_5579);
and U6124 (N_6124,N_5122,N_5651);
nor U6125 (N_6125,N_5256,N_5302);
and U6126 (N_6126,N_5503,N_5973);
nor U6127 (N_6127,N_5171,N_5932);
xor U6128 (N_6128,N_5141,N_5182);
or U6129 (N_6129,N_5917,N_5107);
and U6130 (N_6130,N_5666,N_5565);
and U6131 (N_6131,N_5194,N_5546);
or U6132 (N_6132,N_5787,N_5698);
nand U6133 (N_6133,N_5774,N_5626);
or U6134 (N_6134,N_5555,N_5858);
and U6135 (N_6135,N_5725,N_5540);
nor U6136 (N_6136,N_5986,N_5667);
nand U6137 (N_6137,N_5408,N_5055);
nand U6138 (N_6138,N_5139,N_5021);
or U6139 (N_6139,N_5954,N_5015);
or U6140 (N_6140,N_5349,N_5810);
nor U6141 (N_6141,N_5326,N_5567);
xnor U6142 (N_6142,N_5641,N_5278);
nand U6143 (N_6143,N_5821,N_5423);
nor U6144 (N_6144,N_5718,N_5846);
xnor U6145 (N_6145,N_5893,N_5948);
nand U6146 (N_6146,N_5791,N_5609);
or U6147 (N_6147,N_5515,N_5453);
nor U6148 (N_6148,N_5258,N_5597);
nand U6149 (N_6149,N_5319,N_5089);
nor U6150 (N_6150,N_5478,N_5531);
nand U6151 (N_6151,N_5311,N_5399);
or U6152 (N_6152,N_5232,N_5632);
nand U6153 (N_6153,N_5335,N_5009);
or U6154 (N_6154,N_5697,N_5629);
or U6155 (N_6155,N_5668,N_5385);
or U6156 (N_6156,N_5966,N_5584);
nor U6157 (N_6157,N_5506,N_5392);
nor U6158 (N_6158,N_5128,N_5982);
nand U6159 (N_6159,N_5709,N_5112);
nor U6160 (N_6160,N_5998,N_5451);
xor U6161 (N_6161,N_5611,N_5061);
nand U6162 (N_6162,N_5653,N_5761);
nor U6163 (N_6163,N_5085,N_5437);
and U6164 (N_6164,N_5622,N_5042);
or U6165 (N_6165,N_5708,N_5373);
xor U6166 (N_6166,N_5729,N_5230);
xnor U6167 (N_6167,N_5519,N_5742);
xnor U6168 (N_6168,N_5119,N_5745);
xnor U6169 (N_6169,N_5753,N_5958);
or U6170 (N_6170,N_5902,N_5571);
xnor U6171 (N_6171,N_5925,N_5254);
nand U6172 (N_6172,N_5967,N_5239);
xnor U6173 (N_6173,N_5246,N_5911);
nand U6174 (N_6174,N_5502,N_5722);
and U6175 (N_6175,N_5806,N_5114);
nand U6176 (N_6176,N_5264,N_5877);
nand U6177 (N_6177,N_5165,N_5707);
or U6178 (N_6178,N_5298,N_5635);
and U6179 (N_6179,N_5647,N_5077);
nor U6180 (N_6180,N_5475,N_5886);
nand U6181 (N_6181,N_5510,N_5661);
nor U6182 (N_6182,N_5675,N_5204);
nand U6183 (N_6183,N_5142,N_5975);
nor U6184 (N_6184,N_5535,N_5389);
nor U6185 (N_6185,N_5838,N_5901);
and U6186 (N_6186,N_5360,N_5304);
nor U6187 (N_6187,N_5217,N_5993);
nand U6188 (N_6188,N_5517,N_5832);
and U6189 (N_6189,N_5439,N_5741);
or U6190 (N_6190,N_5092,N_5024);
or U6191 (N_6191,N_5188,N_5860);
or U6192 (N_6192,N_5688,N_5628);
or U6193 (N_6193,N_5702,N_5863);
nand U6194 (N_6194,N_5541,N_5378);
nor U6195 (N_6195,N_5547,N_5383);
nand U6196 (N_6196,N_5164,N_5460);
and U6197 (N_6197,N_5684,N_5445);
or U6198 (N_6198,N_5721,N_5156);
xor U6199 (N_6199,N_5595,N_5201);
or U6200 (N_6200,N_5277,N_5365);
nor U6201 (N_6201,N_5428,N_5501);
and U6202 (N_6202,N_5819,N_5401);
nand U6203 (N_6203,N_5804,N_5454);
or U6204 (N_6204,N_5715,N_5181);
nor U6205 (N_6205,N_5480,N_5777);
nor U6206 (N_6206,N_5236,N_5509);
nand U6207 (N_6207,N_5080,N_5443);
xor U6208 (N_6208,N_5968,N_5683);
nor U6209 (N_6209,N_5736,N_5476);
and U6210 (N_6210,N_5781,N_5110);
or U6211 (N_6211,N_5516,N_5430);
nor U6212 (N_6212,N_5381,N_5020);
or U6213 (N_6213,N_5342,N_5425);
and U6214 (N_6214,N_5468,N_5945);
nor U6215 (N_6215,N_5033,N_5450);
and U6216 (N_6216,N_5316,N_5037);
and U6217 (N_6217,N_5025,N_5250);
and U6218 (N_6218,N_5794,N_5711);
xor U6219 (N_6219,N_5580,N_5784);
or U6220 (N_6220,N_5290,N_5469);
nor U6221 (N_6221,N_5956,N_5382);
nor U6222 (N_6222,N_5652,N_5770);
or U6223 (N_6223,N_5922,N_5490);
nand U6224 (N_6224,N_5590,N_5433);
nand U6225 (N_6225,N_5007,N_5508);
and U6226 (N_6226,N_5604,N_5362);
nand U6227 (N_6227,N_5971,N_5402);
nand U6228 (N_6228,N_5288,N_5151);
or U6229 (N_6229,N_5775,N_5291);
nor U6230 (N_6230,N_5216,N_5521);
xnor U6231 (N_6231,N_5959,N_5814);
and U6232 (N_6232,N_5247,N_5714);
nor U6233 (N_6233,N_5757,N_5023);
or U6234 (N_6234,N_5384,N_5789);
nand U6235 (N_6235,N_5659,N_5340);
nand U6236 (N_6236,N_5780,N_5405);
nor U6237 (N_6237,N_5572,N_5459);
nor U6238 (N_6238,N_5419,N_5148);
xor U6239 (N_6239,N_5103,N_5669);
xor U6240 (N_6240,N_5371,N_5313);
xor U6241 (N_6241,N_5438,N_5321);
xnor U6242 (N_6242,N_5192,N_5213);
nand U6243 (N_6243,N_5497,N_5826);
nor U6244 (N_6244,N_5308,N_5820);
and U6245 (N_6245,N_5650,N_5562);
nor U6246 (N_6246,N_5608,N_5802);
nand U6247 (N_6247,N_5552,N_5586);
or U6248 (N_6248,N_5134,N_5937);
nand U6249 (N_6249,N_5673,N_5404);
and U6250 (N_6250,N_5520,N_5500);
xor U6251 (N_6251,N_5570,N_5545);
or U6252 (N_6252,N_5064,N_5537);
and U6253 (N_6253,N_5146,N_5292);
nand U6254 (N_6254,N_5358,N_5689);
or U6255 (N_6255,N_5491,N_5637);
and U6256 (N_6256,N_5811,N_5665);
or U6257 (N_6257,N_5482,N_5274);
nand U6258 (N_6258,N_5824,N_5703);
and U6259 (N_6259,N_5489,N_5271);
or U6260 (N_6260,N_5084,N_5003);
and U6261 (N_6261,N_5704,N_5926);
or U6262 (N_6262,N_5815,N_5636);
or U6263 (N_6263,N_5086,N_5848);
and U6264 (N_6264,N_5727,N_5897);
and U6265 (N_6265,N_5369,N_5471);
xnor U6266 (N_6266,N_5479,N_5348);
and U6267 (N_6267,N_5257,N_5422);
nor U6268 (N_6268,N_5448,N_5557);
nand U6269 (N_6269,N_5090,N_5123);
nand U6270 (N_6270,N_5638,N_5259);
nor U6271 (N_6271,N_5768,N_5197);
xor U6272 (N_6272,N_5207,N_5228);
or U6273 (N_6273,N_5762,N_5295);
nand U6274 (N_6274,N_5406,N_5807);
and U6275 (N_6275,N_5994,N_5432);
xnor U6276 (N_6276,N_5566,N_5779);
nand U6277 (N_6277,N_5624,N_5203);
xnor U6278 (N_6278,N_5287,N_5625);
or U6279 (N_6279,N_5058,N_5990);
or U6280 (N_6280,N_5109,N_5706);
nand U6281 (N_6281,N_5281,N_5548);
nor U6282 (N_6282,N_5900,N_5198);
xor U6283 (N_6283,N_5286,N_5743);
nor U6284 (N_6284,N_5159,N_5798);
xnor U6285 (N_6285,N_5748,N_5161);
and U6286 (N_6286,N_5133,N_5435);
and U6287 (N_6287,N_5507,N_5485);
nand U6288 (N_6288,N_5320,N_5132);
nand U6289 (N_6289,N_5883,N_5154);
nor U6290 (N_6290,N_5676,N_5610);
nor U6291 (N_6291,N_5909,N_5185);
and U6292 (N_6292,N_5208,N_5184);
nand U6293 (N_6293,N_5912,N_5803);
xor U6294 (N_6294,N_5440,N_5924);
and U6295 (N_6295,N_5550,N_5525);
nand U6296 (N_6296,N_5813,N_5575);
and U6297 (N_6297,N_5822,N_5029);
xor U6298 (N_6298,N_5720,N_5098);
nor U6299 (N_6299,N_5051,N_5346);
and U6300 (N_6300,N_5266,N_5136);
nor U6301 (N_6301,N_5111,N_5394);
and U6302 (N_6302,N_5805,N_5940);
xnor U6303 (N_6303,N_5800,N_5766);
xnor U6304 (N_6304,N_5524,N_5856);
nand U6305 (N_6305,N_5488,N_5788);
nand U6306 (N_6306,N_5568,N_5467);
xor U6307 (N_6307,N_5011,N_5317);
and U6308 (N_6308,N_5569,N_5370);
nand U6309 (N_6309,N_5642,N_5366);
nand U6310 (N_6310,N_5344,N_5963);
and U6311 (N_6311,N_5068,N_5409);
xnor U6312 (N_6312,N_5447,N_5424);
xnor U6313 (N_6313,N_5294,N_5823);
or U6314 (N_6314,N_5646,N_5162);
xnor U6315 (N_6315,N_5289,N_5097);
xnor U6316 (N_6316,N_5004,N_5328);
nand U6317 (N_6317,N_5461,N_5195);
xnor U6318 (N_6318,N_5189,N_5047);
or U6319 (N_6319,N_5592,N_5931);
or U6320 (N_6320,N_5561,N_5825);
or U6321 (N_6321,N_5327,N_5331);
or U6322 (N_6322,N_5938,N_5857);
nand U6323 (N_6323,N_5436,N_5143);
xor U6324 (N_6324,N_5882,N_5692);
nand U6325 (N_6325,N_5072,N_5747);
or U6326 (N_6326,N_5280,N_5231);
nand U6327 (N_6327,N_5726,N_5127);
xor U6328 (N_6328,N_5513,N_5972);
xnor U6329 (N_6329,N_5657,N_5466);
nand U6330 (N_6330,N_5121,N_5056);
and U6331 (N_6331,N_5723,N_5410);
nor U6332 (N_6332,N_5411,N_5458);
and U6333 (N_6333,N_5105,N_5691);
nand U6334 (N_6334,N_5677,N_5889);
or U6335 (N_6335,N_5329,N_5083);
or U6336 (N_6336,N_5953,N_5769);
and U6337 (N_6337,N_5045,N_5840);
nor U6338 (N_6338,N_5376,N_5589);
and U6339 (N_6339,N_5763,N_5390);
xor U6340 (N_6340,N_5639,N_5260);
nand U6341 (N_6341,N_5514,N_5587);
nor U6342 (N_6342,N_5338,N_5904);
nand U6343 (N_6343,N_5532,N_5026);
and U6344 (N_6344,N_5737,N_5379);
and U6345 (N_6345,N_5786,N_5752);
nand U6346 (N_6346,N_5526,N_5002);
and U6347 (N_6347,N_5229,N_5420);
or U6348 (N_6348,N_5942,N_5057);
or U6349 (N_6349,N_5104,N_5974);
nor U6350 (N_6350,N_5393,N_5355);
xor U6351 (N_6351,N_5914,N_5270);
and U6352 (N_6352,N_5307,N_5293);
nor U6353 (N_6353,N_5048,N_5245);
nand U6354 (N_6354,N_5001,N_5014);
and U6355 (N_6355,N_5377,N_5740);
xor U6356 (N_6356,N_5828,N_5046);
xnor U6357 (N_6357,N_5744,N_5941);
nand U6358 (N_6358,N_5063,N_5867);
nor U6359 (N_6359,N_5028,N_5173);
xnor U6360 (N_6360,N_5240,N_5332);
or U6361 (N_6361,N_5620,N_5992);
nor U6362 (N_6362,N_5836,N_5071);
nor U6363 (N_6363,N_5153,N_5760);
and U6364 (N_6364,N_5928,N_5504);
xor U6365 (N_6365,N_5920,N_5494);
or U6366 (N_6366,N_5053,N_5558);
nor U6367 (N_6367,N_5492,N_5462);
nor U6368 (N_6368,N_5888,N_5324);
nor U6369 (N_6369,N_5599,N_5615);
nand U6370 (N_6370,N_5607,N_5574);
or U6371 (N_6371,N_5630,N_5299);
or U6372 (N_6372,N_5218,N_5773);
and U6373 (N_6373,N_5255,N_5160);
or U6374 (N_6374,N_5158,N_5962);
and U6375 (N_6375,N_5598,N_5027);
or U6376 (N_6376,N_5918,N_5243);
nor U6377 (N_6377,N_5553,N_5339);
nand U6378 (N_6378,N_5403,N_5284);
or U6379 (N_6379,N_5983,N_5852);
xnor U6380 (N_6380,N_5065,N_5221);
or U6381 (N_6381,N_5434,N_5073);
xnor U6382 (N_6382,N_5596,N_5374);
xor U6383 (N_6383,N_5474,N_5903);
or U6384 (N_6384,N_5426,N_5576);
and U6385 (N_6385,N_5441,N_5728);
nand U6386 (N_6386,N_5544,N_5674);
or U6387 (N_6387,N_5272,N_5223);
and U6388 (N_6388,N_5038,N_5581);
or U6389 (N_6389,N_5533,N_5679);
nor U6390 (N_6390,N_5767,N_5606);
nor U6391 (N_6391,N_5785,N_5163);
or U6392 (N_6392,N_5301,N_5352);
nor U6393 (N_6393,N_5251,N_5129);
nor U6394 (N_6394,N_5844,N_5782);
nand U6395 (N_6395,N_5252,N_5870);
xor U6396 (N_6396,N_5927,N_5303);
nor U6397 (N_6397,N_5554,N_5809);
and U6398 (N_6398,N_5078,N_5414);
or U6399 (N_6399,N_5484,N_5361);
or U6400 (N_6400,N_5869,N_5060);
or U6401 (N_6401,N_5052,N_5952);
xor U6402 (N_6402,N_5431,N_5407);
xor U6403 (N_6403,N_5323,N_5523);
nor U6404 (N_6404,N_5776,N_5818);
and U6405 (N_6405,N_5772,N_5705);
or U6406 (N_6406,N_5839,N_5594);
xor U6407 (N_6407,N_5670,N_5884);
or U6408 (N_6408,N_5357,N_5701);
nor U6409 (N_6409,N_5174,N_5457);
nand U6410 (N_6410,N_5261,N_5368);
nand U6411 (N_6411,N_5588,N_5031);
nand U6412 (N_6412,N_5979,N_5269);
nor U6413 (N_6413,N_5756,N_5253);
nor U6414 (N_6414,N_5242,N_5859);
xor U6415 (N_6415,N_5322,N_5297);
nand U6416 (N_6416,N_5618,N_5957);
nand U6417 (N_6417,N_5093,N_5070);
or U6418 (N_6418,N_5634,N_5455);
nand U6419 (N_6419,N_5310,N_5131);
or U6420 (N_6420,N_5969,N_5074);
nand U6421 (N_6421,N_5210,N_5233);
and U6422 (N_6422,N_5754,N_5343);
nand U6423 (N_6423,N_5663,N_5719);
nand U6424 (N_6424,N_5180,N_5874);
nand U6425 (N_6425,N_5044,N_5585);
nand U6426 (N_6426,N_5593,N_5397);
xnor U6427 (N_6427,N_5619,N_5627);
or U6428 (N_6428,N_5559,N_5429);
xnor U6429 (N_6429,N_5536,N_5341);
xor U6430 (N_6430,N_5267,N_5325);
xor U6431 (N_6431,N_5835,N_5463);
and U6432 (N_6432,N_5413,N_5934);
xor U6433 (N_6433,N_5040,N_5850);
nand U6434 (N_6434,N_5916,N_5296);
nor U6435 (N_6435,N_5853,N_5563);
and U6436 (N_6436,N_5660,N_5099);
nand U6437 (N_6437,N_5495,N_5551);
xor U6438 (N_6438,N_5996,N_5241);
nor U6439 (N_6439,N_5793,N_5534);
nand U6440 (N_6440,N_5612,N_5464);
xnor U6441 (N_6441,N_5614,N_5880);
xnor U6442 (N_6442,N_5059,N_5955);
nand U6443 (N_6443,N_5032,N_5738);
nor U6444 (N_6444,N_5717,N_5512);
xor U6445 (N_6445,N_5583,N_5309);
or U6446 (N_6446,N_5102,N_5999);
nor U6447 (N_6447,N_5211,N_5687);
and U6448 (N_6448,N_5087,N_5452);
xor U6449 (N_6449,N_5656,N_5896);
nor U6450 (N_6450,N_5831,N_5834);
nand U6451 (N_6451,N_5169,N_5529);
nor U6452 (N_6452,N_5273,N_5530);
xor U6453 (N_6453,N_5746,N_5947);
or U6454 (N_6454,N_5222,N_5345);
or U6455 (N_6455,N_5013,N_5716);
and U6456 (N_6456,N_5915,N_5167);
or U6457 (N_6457,N_5206,N_5528);
xor U6458 (N_6458,N_5175,N_5985);
or U6459 (N_6459,N_5602,N_5237);
and U6460 (N_6460,N_5700,N_5199);
xnor U6461 (N_6461,N_5472,N_5987);
and U6462 (N_6462,N_5306,N_5279);
xor U6463 (N_6463,N_5778,N_5792);
xor U6464 (N_6464,N_5449,N_5933);
nand U6465 (N_6465,N_5054,N_5511);
or U6466 (N_6466,N_5991,N_5732);
nand U6467 (N_6467,N_5808,N_5006);
xnor U6468 (N_6468,N_5830,N_5062);
nand U6469 (N_6469,N_5817,N_5417);
or U6470 (N_6470,N_5049,N_5898);
and U6471 (N_6471,N_5919,N_5759);
nand U6472 (N_6472,N_5069,N_5444);
and U6473 (N_6473,N_5350,N_5699);
or U6474 (N_6474,N_5081,N_5268);
and U6475 (N_6475,N_5499,N_5879);
and U6476 (N_6476,N_5137,N_5891);
and U6477 (N_6477,N_5205,N_5505);
nor U6478 (N_6478,N_5030,N_5997);
or U6479 (N_6479,N_5895,N_5796);
xor U6480 (N_6480,N_5496,N_5923);
nor U6481 (N_6481,N_5664,N_5845);
xnor U6482 (N_6482,N_5750,N_5019);
and U6483 (N_6483,N_5984,N_5400);
or U6484 (N_6484,N_5949,N_5012);
nand U6485 (N_6485,N_5166,N_5976);
nand U6486 (N_6486,N_5855,N_5398);
and U6487 (N_6487,N_5908,N_5050);
or U6488 (N_6488,N_5091,N_5890);
xor U6489 (N_6489,N_5367,N_5605);
xnor U6490 (N_6490,N_5861,N_5094);
nor U6491 (N_6491,N_5145,N_5578);
nor U6492 (N_6492,N_5686,N_5416);
xnor U6493 (N_6493,N_5276,N_5249);
xor U6494 (N_6494,N_5887,N_5739);
or U6495 (N_6495,N_5631,N_5395);
xnor U6496 (N_6496,N_5640,N_5108);
nor U6497 (N_6497,N_5951,N_5685);
xor U6498 (N_6498,N_5200,N_5238);
and U6499 (N_6499,N_5190,N_5186);
nor U6500 (N_6500,N_5018,N_5634);
and U6501 (N_6501,N_5055,N_5430);
or U6502 (N_6502,N_5606,N_5919);
xnor U6503 (N_6503,N_5666,N_5530);
xnor U6504 (N_6504,N_5001,N_5257);
nand U6505 (N_6505,N_5682,N_5257);
or U6506 (N_6506,N_5719,N_5750);
or U6507 (N_6507,N_5422,N_5537);
nand U6508 (N_6508,N_5399,N_5306);
and U6509 (N_6509,N_5327,N_5782);
and U6510 (N_6510,N_5422,N_5743);
or U6511 (N_6511,N_5763,N_5864);
and U6512 (N_6512,N_5450,N_5152);
or U6513 (N_6513,N_5877,N_5065);
xor U6514 (N_6514,N_5450,N_5791);
xnor U6515 (N_6515,N_5977,N_5233);
and U6516 (N_6516,N_5076,N_5186);
or U6517 (N_6517,N_5097,N_5058);
nor U6518 (N_6518,N_5061,N_5575);
or U6519 (N_6519,N_5776,N_5504);
or U6520 (N_6520,N_5645,N_5840);
or U6521 (N_6521,N_5035,N_5818);
and U6522 (N_6522,N_5395,N_5934);
xor U6523 (N_6523,N_5533,N_5511);
nor U6524 (N_6524,N_5906,N_5755);
nand U6525 (N_6525,N_5341,N_5075);
xnor U6526 (N_6526,N_5315,N_5638);
nand U6527 (N_6527,N_5576,N_5805);
nor U6528 (N_6528,N_5942,N_5694);
nor U6529 (N_6529,N_5607,N_5727);
and U6530 (N_6530,N_5270,N_5041);
and U6531 (N_6531,N_5258,N_5723);
nand U6532 (N_6532,N_5456,N_5042);
xnor U6533 (N_6533,N_5768,N_5352);
nor U6534 (N_6534,N_5089,N_5025);
xnor U6535 (N_6535,N_5759,N_5332);
nor U6536 (N_6536,N_5645,N_5433);
nand U6537 (N_6537,N_5747,N_5706);
xnor U6538 (N_6538,N_5466,N_5969);
and U6539 (N_6539,N_5645,N_5934);
xor U6540 (N_6540,N_5465,N_5880);
and U6541 (N_6541,N_5365,N_5895);
or U6542 (N_6542,N_5169,N_5914);
and U6543 (N_6543,N_5700,N_5039);
xor U6544 (N_6544,N_5153,N_5688);
nor U6545 (N_6545,N_5347,N_5188);
or U6546 (N_6546,N_5648,N_5909);
nand U6547 (N_6547,N_5976,N_5389);
nor U6548 (N_6548,N_5231,N_5942);
and U6549 (N_6549,N_5677,N_5527);
or U6550 (N_6550,N_5361,N_5337);
nand U6551 (N_6551,N_5777,N_5937);
nand U6552 (N_6552,N_5976,N_5592);
nand U6553 (N_6553,N_5081,N_5134);
xnor U6554 (N_6554,N_5178,N_5901);
xnor U6555 (N_6555,N_5356,N_5669);
xor U6556 (N_6556,N_5414,N_5968);
or U6557 (N_6557,N_5978,N_5232);
and U6558 (N_6558,N_5967,N_5116);
and U6559 (N_6559,N_5090,N_5971);
or U6560 (N_6560,N_5201,N_5108);
nor U6561 (N_6561,N_5020,N_5137);
xnor U6562 (N_6562,N_5304,N_5440);
and U6563 (N_6563,N_5432,N_5524);
nand U6564 (N_6564,N_5781,N_5452);
nand U6565 (N_6565,N_5592,N_5693);
nor U6566 (N_6566,N_5143,N_5434);
nand U6567 (N_6567,N_5769,N_5330);
nand U6568 (N_6568,N_5929,N_5399);
nand U6569 (N_6569,N_5336,N_5229);
xnor U6570 (N_6570,N_5885,N_5347);
and U6571 (N_6571,N_5099,N_5581);
nor U6572 (N_6572,N_5332,N_5502);
nor U6573 (N_6573,N_5681,N_5301);
nand U6574 (N_6574,N_5733,N_5137);
nor U6575 (N_6575,N_5745,N_5157);
or U6576 (N_6576,N_5447,N_5078);
nand U6577 (N_6577,N_5665,N_5784);
nand U6578 (N_6578,N_5540,N_5580);
nor U6579 (N_6579,N_5803,N_5623);
xor U6580 (N_6580,N_5467,N_5828);
or U6581 (N_6581,N_5731,N_5607);
nor U6582 (N_6582,N_5863,N_5785);
and U6583 (N_6583,N_5703,N_5380);
nor U6584 (N_6584,N_5963,N_5036);
xor U6585 (N_6585,N_5811,N_5683);
nor U6586 (N_6586,N_5382,N_5571);
xor U6587 (N_6587,N_5734,N_5118);
xnor U6588 (N_6588,N_5541,N_5430);
nand U6589 (N_6589,N_5089,N_5951);
xnor U6590 (N_6590,N_5659,N_5799);
xnor U6591 (N_6591,N_5439,N_5314);
nor U6592 (N_6592,N_5782,N_5581);
and U6593 (N_6593,N_5437,N_5968);
xor U6594 (N_6594,N_5857,N_5670);
xor U6595 (N_6595,N_5735,N_5774);
or U6596 (N_6596,N_5356,N_5211);
nor U6597 (N_6597,N_5373,N_5309);
or U6598 (N_6598,N_5547,N_5739);
nor U6599 (N_6599,N_5879,N_5341);
nand U6600 (N_6600,N_5041,N_5293);
nand U6601 (N_6601,N_5328,N_5348);
or U6602 (N_6602,N_5147,N_5732);
nor U6603 (N_6603,N_5975,N_5576);
and U6604 (N_6604,N_5062,N_5328);
and U6605 (N_6605,N_5662,N_5854);
and U6606 (N_6606,N_5574,N_5006);
nand U6607 (N_6607,N_5043,N_5734);
xor U6608 (N_6608,N_5896,N_5422);
xnor U6609 (N_6609,N_5543,N_5224);
nand U6610 (N_6610,N_5009,N_5870);
or U6611 (N_6611,N_5591,N_5445);
nand U6612 (N_6612,N_5455,N_5011);
and U6613 (N_6613,N_5102,N_5215);
xor U6614 (N_6614,N_5896,N_5094);
nor U6615 (N_6615,N_5845,N_5073);
or U6616 (N_6616,N_5875,N_5282);
or U6617 (N_6617,N_5049,N_5422);
nand U6618 (N_6618,N_5005,N_5641);
and U6619 (N_6619,N_5455,N_5227);
nand U6620 (N_6620,N_5359,N_5384);
xnor U6621 (N_6621,N_5906,N_5665);
nand U6622 (N_6622,N_5378,N_5603);
and U6623 (N_6623,N_5881,N_5748);
nor U6624 (N_6624,N_5660,N_5201);
xnor U6625 (N_6625,N_5414,N_5250);
and U6626 (N_6626,N_5991,N_5664);
xnor U6627 (N_6627,N_5580,N_5497);
nand U6628 (N_6628,N_5294,N_5573);
nand U6629 (N_6629,N_5636,N_5476);
or U6630 (N_6630,N_5037,N_5059);
xnor U6631 (N_6631,N_5303,N_5272);
nor U6632 (N_6632,N_5296,N_5469);
xnor U6633 (N_6633,N_5290,N_5256);
nor U6634 (N_6634,N_5981,N_5320);
nor U6635 (N_6635,N_5611,N_5383);
xnor U6636 (N_6636,N_5645,N_5705);
nand U6637 (N_6637,N_5253,N_5969);
nand U6638 (N_6638,N_5918,N_5139);
nor U6639 (N_6639,N_5741,N_5988);
and U6640 (N_6640,N_5782,N_5788);
nor U6641 (N_6641,N_5929,N_5395);
and U6642 (N_6642,N_5569,N_5652);
nand U6643 (N_6643,N_5873,N_5017);
or U6644 (N_6644,N_5324,N_5936);
nand U6645 (N_6645,N_5542,N_5355);
and U6646 (N_6646,N_5247,N_5141);
nand U6647 (N_6647,N_5867,N_5043);
or U6648 (N_6648,N_5272,N_5225);
xnor U6649 (N_6649,N_5012,N_5819);
nor U6650 (N_6650,N_5260,N_5676);
nand U6651 (N_6651,N_5606,N_5036);
xnor U6652 (N_6652,N_5509,N_5454);
nor U6653 (N_6653,N_5945,N_5297);
nand U6654 (N_6654,N_5617,N_5210);
nor U6655 (N_6655,N_5383,N_5416);
or U6656 (N_6656,N_5233,N_5945);
or U6657 (N_6657,N_5866,N_5490);
nand U6658 (N_6658,N_5488,N_5732);
nand U6659 (N_6659,N_5424,N_5603);
nor U6660 (N_6660,N_5501,N_5302);
xnor U6661 (N_6661,N_5914,N_5848);
nor U6662 (N_6662,N_5204,N_5697);
xor U6663 (N_6663,N_5176,N_5014);
xor U6664 (N_6664,N_5188,N_5670);
or U6665 (N_6665,N_5368,N_5296);
xnor U6666 (N_6666,N_5067,N_5834);
nand U6667 (N_6667,N_5601,N_5421);
and U6668 (N_6668,N_5239,N_5206);
nand U6669 (N_6669,N_5375,N_5480);
or U6670 (N_6670,N_5979,N_5014);
nand U6671 (N_6671,N_5935,N_5054);
xor U6672 (N_6672,N_5933,N_5705);
nor U6673 (N_6673,N_5420,N_5981);
nor U6674 (N_6674,N_5609,N_5119);
xnor U6675 (N_6675,N_5797,N_5610);
nand U6676 (N_6676,N_5790,N_5138);
nor U6677 (N_6677,N_5245,N_5643);
or U6678 (N_6678,N_5752,N_5081);
and U6679 (N_6679,N_5505,N_5967);
nor U6680 (N_6680,N_5209,N_5146);
nand U6681 (N_6681,N_5552,N_5882);
or U6682 (N_6682,N_5624,N_5703);
or U6683 (N_6683,N_5677,N_5633);
nand U6684 (N_6684,N_5381,N_5158);
and U6685 (N_6685,N_5101,N_5983);
or U6686 (N_6686,N_5643,N_5856);
nand U6687 (N_6687,N_5501,N_5147);
nand U6688 (N_6688,N_5539,N_5821);
xnor U6689 (N_6689,N_5692,N_5242);
or U6690 (N_6690,N_5240,N_5747);
nand U6691 (N_6691,N_5774,N_5210);
xnor U6692 (N_6692,N_5334,N_5419);
nand U6693 (N_6693,N_5547,N_5385);
nand U6694 (N_6694,N_5234,N_5104);
xnor U6695 (N_6695,N_5123,N_5184);
or U6696 (N_6696,N_5022,N_5168);
nand U6697 (N_6697,N_5250,N_5189);
or U6698 (N_6698,N_5123,N_5468);
nand U6699 (N_6699,N_5693,N_5871);
nand U6700 (N_6700,N_5408,N_5325);
nand U6701 (N_6701,N_5359,N_5770);
and U6702 (N_6702,N_5625,N_5873);
or U6703 (N_6703,N_5790,N_5599);
and U6704 (N_6704,N_5450,N_5874);
and U6705 (N_6705,N_5947,N_5065);
or U6706 (N_6706,N_5623,N_5915);
and U6707 (N_6707,N_5957,N_5212);
or U6708 (N_6708,N_5507,N_5857);
or U6709 (N_6709,N_5350,N_5351);
nor U6710 (N_6710,N_5641,N_5461);
xor U6711 (N_6711,N_5957,N_5643);
nor U6712 (N_6712,N_5706,N_5694);
xor U6713 (N_6713,N_5526,N_5171);
nor U6714 (N_6714,N_5016,N_5619);
xnor U6715 (N_6715,N_5147,N_5314);
and U6716 (N_6716,N_5839,N_5056);
nand U6717 (N_6717,N_5295,N_5810);
nand U6718 (N_6718,N_5091,N_5540);
nor U6719 (N_6719,N_5315,N_5196);
nor U6720 (N_6720,N_5990,N_5344);
xor U6721 (N_6721,N_5096,N_5894);
and U6722 (N_6722,N_5088,N_5076);
or U6723 (N_6723,N_5783,N_5687);
xor U6724 (N_6724,N_5921,N_5869);
xor U6725 (N_6725,N_5874,N_5603);
nand U6726 (N_6726,N_5400,N_5651);
xnor U6727 (N_6727,N_5500,N_5700);
and U6728 (N_6728,N_5744,N_5507);
xor U6729 (N_6729,N_5543,N_5785);
nand U6730 (N_6730,N_5970,N_5679);
nand U6731 (N_6731,N_5608,N_5893);
and U6732 (N_6732,N_5255,N_5044);
nand U6733 (N_6733,N_5709,N_5300);
or U6734 (N_6734,N_5264,N_5846);
nor U6735 (N_6735,N_5458,N_5188);
nor U6736 (N_6736,N_5306,N_5096);
or U6737 (N_6737,N_5640,N_5642);
nor U6738 (N_6738,N_5915,N_5662);
or U6739 (N_6739,N_5269,N_5919);
nand U6740 (N_6740,N_5245,N_5698);
nand U6741 (N_6741,N_5478,N_5071);
nand U6742 (N_6742,N_5867,N_5905);
xor U6743 (N_6743,N_5147,N_5931);
nor U6744 (N_6744,N_5270,N_5992);
nor U6745 (N_6745,N_5416,N_5402);
or U6746 (N_6746,N_5173,N_5250);
nand U6747 (N_6747,N_5724,N_5568);
xor U6748 (N_6748,N_5910,N_5399);
nand U6749 (N_6749,N_5300,N_5731);
nand U6750 (N_6750,N_5753,N_5858);
nand U6751 (N_6751,N_5263,N_5179);
or U6752 (N_6752,N_5268,N_5350);
and U6753 (N_6753,N_5910,N_5986);
xor U6754 (N_6754,N_5912,N_5144);
or U6755 (N_6755,N_5648,N_5708);
xnor U6756 (N_6756,N_5267,N_5798);
and U6757 (N_6757,N_5758,N_5163);
xnor U6758 (N_6758,N_5902,N_5634);
xor U6759 (N_6759,N_5209,N_5831);
and U6760 (N_6760,N_5232,N_5458);
nand U6761 (N_6761,N_5604,N_5471);
xnor U6762 (N_6762,N_5832,N_5059);
nand U6763 (N_6763,N_5521,N_5670);
nand U6764 (N_6764,N_5243,N_5930);
and U6765 (N_6765,N_5264,N_5975);
and U6766 (N_6766,N_5910,N_5531);
nor U6767 (N_6767,N_5881,N_5707);
or U6768 (N_6768,N_5520,N_5710);
nor U6769 (N_6769,N_5963,N_5594);
or U6770 (N_6770,N_5737,N_5088);
xor U6771 (N_6771,N_5210,N_5395);
nand U6772 (N_6772,N_5018,N_5109);
nor U6773 (N_6773,N_5334,N_5465);
or U6774 (N_6774,N_5601,N_5006);
nor U6775 (N_6775,N_5222,N_5217);
nor U6776 (N_6776,N_5204,N_5515);
nor U6777 (N_6777,N_5712,N_5543);
xnor U6778 (N_6778,N_5784,N_5482);
nand U6779 (N_6779,N_5032,N_5034);
and U6780 (N_6780,N_5894,N_5434);
and U6781 (N_6781,N_5726,N_5883);
or U6782 (N_6782,N_5041,N_5371);
and U6783 (N_6783,N_5264,N_5736);
nand U6784 (N_6784,N_5793,N_5838);
nand U6785 (N_6785,N_5284,N_5044);
or U6786 (N_6786,N_5485,N_5593);
nand U6787 (N_6787,N_5338,N_5637);
and U6788 (N_6788,N_5327,N_5607);
nand U6789 (N_6789,N_5955,N_5957);
and U6790 (N_6790,N_5296,N_5634);
or U6791 (N_6791,N_5640,N_5249);
nand U6792 (N_6792,N_5897,N_5561);
and U6793 (N_6793,N_5040,N_5076);
nand U6794 (N_6794,N_5562,N_5688);
nand U6795 (N_6795,N_5975,N_5966);
nand U6796 (N_6796,N_5810,N_5780);
xor U6797 (N_6797,N_5409,N_5325);
and U6798 (N_6798,N_5183,N_5790);
and U6799 (N_6799,N_5026,N_5068);
or U6800 (N_6800,N_5526,N_5945);
nor U6801 (N_6801,N_5626,N_5436);
or U6802 (N_6802,N_5970,N_5766);
nor U6803 (N_6803,N_5868,N_5107);
nand U6804 (N_6804,N_5743,N_5395);
or U6805 (N_6805,N_5934,N_5307);
xnor U6806 (N_6806,N_5263,N_5316);
nand U6807 (N_6807,N_5480,N_5148);
and U6808 (N_6808,N_5767,N_5936);
xor U6809 (N_6809,N_5204,N_5229);
and U6810 (N_6810,N_5857,N_5256);
and U6811 (N_6811,N_5584,N_5282);
or U6812 (N_6812,N_5567,N_5786);
and U6813 (N_6813,N_5101,N_5812);
xor U6814 (N_6814,N_5483,N_5235);
or U6815 (N_6815,N_5508,N_5279);
and U6816 (N_6816,N_5533,N_5242);
and U6817 (N_6817,N_5247,N_5098);
xnor U6818 (N_6818,N_5163,N_5969);
nand U6819 (N_6819,N_5316,N_5219);
and U6820 (N_6820,N_5258,N_5782);
and U6821 (N_6821,N_5777,N_5271);
and U6822 (N_6822,N_5579,N_5032);
and U6823 (N_6823,N_5818,N_5873);
xnor U6824 (N_6824,N_5559,N_5165);
or U6825 (N_6825,N_5658,N_5430);
xor U6826 (N_6826,N_5525,N_5271);
and U6827 (N_6827,N_5520,N_5756);
nor U6828 (N_6828,N_5710,N_5529);
nand U6829 (N_6829,N_5332,N_5902);
or U6830 (N_6830,N_5829,N_5635);
nor U6831 (N_6831,N_5033,N_5819);
and U6832 (N_6832,N_5115,N_5837);
nor U6833 (N_6833,N_5026,N_5519);
and U6834 (N_6834,N_5791,N_5643);
nor U6835 (N_6835,N_5993,N_5967);
nor U6836 (N_6836,N_5669,N_5908);
or U6837 (N_6837,N_5396,N_5931);
and U6838 (N_6838,N_5879,N_5762);
xor U6839 (N_6839,N_5575,N_5440);
or U6840 (N_6840,N_5166,N_5088);
nand U6841 (N_6841,N_5120,N_5910);
and U6842 (N_6842,N_5226,N_5257);
xor U6843 (N_6843,N_5602,N_5791);
nor U6844 (N_6844,N_5136,N_5662);
or U6845 (N_6845,N_5859,N_5130);
nand U6846 (N_6846,N_5589,N_5625);
and U6847 (N_6847,N_5621,N_5406);
xor U6848 (N_6848,N_5136,N_5204);
nand U6849 (N_6849,N_5845,N_5355);
or U6850 (N_6850,N_5780,N_5947);
or U6851 (N_6851,N_5725,N_5489);
nor U6852 (N_6852,N_5198,N_5547);
nand U6853 (N_6853,N_5644,N_5907);
or U6854 (N_6854,N_5300,N_5735);
and U6855 (N_6855,N_5531,N_5152);
nor U6856 (N_6856,N_5434,N_5205);
or U6857 (N_6857,N_5888,N_5749);
nand U6858 (N_6858,N_5151,N_5507);
nor U6859 (N_6859,N_5180,N_5371);
xor U6860 (N_6860,N_5015,N_5945);
nor U6861 (N_6861,N_5839,N_5218);
xor U6862 (N_6862,N_5157,N_5374);
xor U6863 (N_6863,N_5164,N_5433);
xnor U6864 (N_6864,N_5504,N_5580);
xor U6865 (N_6865,N_5123,N_5831);
nor U6866 (N_6866,N_5551,N_5334);
nand U6867 (N_6867,N_5201,N_5772);
xnor U6868 (N_6868,N_5519,N_5628);
nand U6869 (N_6869,N_5530,N_5659);
nand U6870 (N_6870,N_5659,N_5134);
and U6871 (N_6871,N_5400,N_5443);
nor U6872 (N_6872,N_5193,N_5183);
and U6873 (N_6873,N_5712,N_5906);
or U6874 (N_6874,N_5490,N_5852);
xnor U6875 (N_6875,N_5728,N_5208);
or U6876 (N_6876,N_5128,N_5824);
nor U6877 (N_6877,N_5876,N_5119);
nor U6878 (N_6878,N_5937,N_5446);
or U6879 (N_6879,N_5142,N_5765);
or U6880 (N_6880,N_5677,N_5999);
nor U6881 (N_6881,N_5993,N_5526);
xnor U6882 (N_6882,N_5646,N_5486);
and U6883 (N_6883,N_5257,N_5967);
or U6884 (N_6884,N_5241,N_5181);
and U6885 (N_6885,N_5381,N_5956);
or U6886 (N_6886,N_5672,N_5280);
or U6887 (N_6887,N_5518,N_5656);
xnor U6888 (N_6888,N_5115,N_5568);
or U6889 (N_6889,N_5464,N_5965);
and U6890 (N_6890,N_5950,N_5641);
xor U6891 (N_6891,N_5669,N_5127);
nand U6892 (N_6892,N_5517,N_5458);
or U6893 (N_6893,N_5167,N_5134);
nor U6894 (N_6894,N_5914,N_5515);
nor U6895 (N_6895,N_5683,N_5881);
xnor U6896 (N_6896,N_5701,N_5187);
nor U6897 (N_6897,N_5327,N_5979);
and U6898 (N_6898,N_5242,N_5752);
xor U6899 (N_6899,N_5632,N_5181);
xnor U6900 (N_6900,N_5520,N_5237);
and U6901 (N_6901,N_5609,N_5074);
nor U6902 (N_6902,N_5862,N_5679);
xor U6903 (N_6903,N_5155,N_5329);
nor U6904 (N_6904,N_5786,N_5726);
and U6905 (N_6905,N_5836,N_5182);
and U6906 (N_6906,N_5675,N_5825);
and U6907 (N_6907,N_5854,N_5683);
or U6908 (N_6908,N_5937,N_5471);
and U6909 (N_6909,N_5026,N_5145);
and U6910 (N_6910,N_5022,N_5062);
and U6911 (N_6911,N_5680,N_5895);
and U6912 (N_6912,N_5401,N_5946);
or U6913 (N_6913,N_5054,N_5432);
or U6914 (N_6914,N_5820,N_5601);
or U6915 (N_6915,N_5022,N_5200);
or U6916 (N_6916,N_5112,N_5969);
xnor U6917 (N_6917,N_5253,N_5396);
and U6918 (N_6918,N_5264,N_5742);
or U6919 (N_6919,N_5649,N_5085);
nor U6920 (N_6920,N_5307,N_5180);
and U6921 (N_6921,N_5563,N_5390);
xnor U6922 (N_6922,N_5621,N_5824);
and U6923 (N_6923,N_5327,N_5323);
nor U6924 (N_6924,N_5764,N_5909);
or U6925 (N_6925,N_5499,N_5702);
or U6926 (N_6926,N_5579,N_5103);
or U6927 (N_6927,N_5210,N_5489);
nand U6928 (N_6928,N_5422,N_5467);
nand U6929 (N_6929,N_5215,N_5314);
xor U6930 (N_6930,N_5412,N_5986);
or U6931 (N_6931,N_5362,N_5260);
or U6932 (N_6932,N_5111,N_5399);
nand U6933 (N_6933,N_5928,N_5722);
xor U6934 (N_6934,N_5741,N_5835);
or U6935 (N_6935,N_5988,N_5070);
or U6936 (N_6936,N_5598,N_5579);
xor U6937 (N_6937,N_5227,N_5004);
xnor U6938 (N_6938,N_5713,N_5261);
xnor U6939 (N_6939,N_5357,N_5741);
xor U6940 (N_6940,N_5900,N_5480);
nand U6941 (N_6941,N_5658,N_5504);
nor U6942 (N_6942,N_5616,N_5453);
nand U6943 (N_6943,N_5796,N_5894);
or U6944 (N_6944,N_5290,N_5462);
xnor U6945 (N_6945,N_5839,N_5394);
and U6946 (N_6946,N_5118,N_5878);
and U6947 (N_6947,N_5998,N_5280);
nor U6948 (N_6948,N_5984,N_5611);
or U6949 (N_6949,N_5110,N_5755);
nand U6950 (N_6950,N_5871,N_5214);
nand U6951 (N_6951,N_5871,N_5552);
nor U6952 (N_6952,N_5013,N_5106);
xnor U6953 (N_6953,N_5731,N_5578);
nor U6954 (N_6954,N_5449,N_5137);
and U6955 (N_6955,N_5165,N_5016);
xnor U6956 (N_6956,N_5291,N_5727);
nor U6957 (N_6957,N_5794,N_5439);
nor U6958 (N_6958,N_5395,N_5949);
and U6959 (N_6959,N_5751,N_5167);
or U6960 (N_6960,N_5925,N_5568);
or U6961 (N_6961,N_5290,N_5289);
or U6962 (N_6962,N_5081,N_5961);
nor U6963 (N_6963,N_5543,N_5878);
nand U6964 (N_6964,N_5311,N_5419);
nand U6965 (N_6965,N_5999,N_5235);
nor U6966 (N_6966,N_5725,N_5928);
and U6967 (N_6967,N_5489,N_5188);
nand U6968 (N_6968,N_5033,N_5998);
and U6969 (N_6969,N_5548,N_5533);
or U6970 (N_6970,N_5546,N_5598);
or U6971 (N_6971,N_5813,N_5915);
and U6972 (N_6972,N_5206,N_5542);
and U6973 (N_6973,N_5850,N_5101);
nor U6974 (N_6974,N_5956,N_5248);
xnor U6975 (N_6975,N_5126,N_5048);
and U6976 (N_6976,N_5962,N_5336);
nor U6977 (N_6977,N_5727,N_5957);
or U6978 (N_6978,N_5309,N_5483);
nand U6979 (N_6979,N_5403,N_5989);
or U6980 (N_6980,N_5111,N_5264);
nor U6981 (N_6981,N_5838,N_5451);
or U6982 (N_6982,N_5784,N_5742);
nor U6983 (N_6983,N_5501,N_5406);
nor U6984 (N_6984,N_5195,N_5526);
and U6985 (N_6985,N_5371,N_5694);
and U6986 (N_6986,N_5442,N_5816);
or U6987 (N_6987,N_5203,N_5735);
and U6988 (N_6988,N_5014,N_5142);
or U6989 (N_6989,N_5522,N_5531);
and U6990 (N_6990,N_5360,N_5395);
xnor U6991 (N_6991,N_5349,N_5071);
nand U6992 (N_6992,N_5672,N_5702);
nor U6993 (N_6993,N_5229,N_5457);
or U6994 (N_6994,N_5801,N_5645);
or U6995 (N_6995,N_5875,N_5081);
and U6996 (N_6996,N_5228,N_5076);
xnor U6997 (N_6997,N_5436,N_5252);
nand U6998 (N_6998,N_5355,N_5044);
nor U6999 (N_6999,N_5799,N_5076);
or U7000 (N_7000,N_6325,N_6090);
xor U7001 (N_7001,N_6746,N_6542);
and U7002 (N_7002,N_6328,N_6705);
xnor U7003 (N_7003,N_6394,N_6477);
and U7004 (N_7004,N_6471,N_6534);
xnor U7005 (N_7005,N_6482,N_6064);
nor U7006 (N_7006,N_6178,N_6146);
nor U7007 (N_7007,N_6889,N_6073);
nor U7008 (N_7008,N_6019,N_6526);
xor U7009 (N_7009,N_6290,N_6958);
nand U7010 (N_7010,N_6005,N_6969);
or U7011 (N_7011,N_6934,N_6404);
nand U7012 (N_7012,N_6143,N_6628);
and U7013 (N_7013,N_6784,N_6110);
or U7014 (N_7014,N_6540,N_6268);
nor U7015 (N_7015,N_6140,N_6931);
nor U7016 (N_7016,N_6393,N_6108);
or U7017 (N_7017,N_6646,N_6311);
and U7018 (N_7018,N_6704,N_6864);
xor U7019 (N_7019,N_6687,N_6085);
nor U7020 (N_7020,N_6608,N_6500);
or U7021 (N_7021,N_6484,N_6677);
nand U7022 (N_7022,N_6047,N_6385);
nor U7023 (N_7023,N_6868,N_6811);
and U7024 (N_7024,N_6314,N_6298);
or U7025 (N_7025,N_6456,N_6932);
nand U7026 (N_7026,N_6904,N_6375);
nand U7027 (N_7027,N_6539,N_6643);
nand U7028 (N_7028,N_6610,N_6360);
xnor U7029 (N_7029,N_6246,N_6755);
and U7030 (N_7030,N_6693,N_6873);
xnor U7031 (N_7031,N_6149,N_6997);
xor U7032 (N_7032,N_6288,N_6816);
or U7033 (N_7033,N_6415,N_6176);
xor U7034 (N_7034,N_6479,N_6720);
nand U7035 (N_7035,N_6545,N_6383);
xor U7036 (N_7036,N_6758,N_6406);
or U7037 (N_7037,N_6035,N_6434);
xnor U7038 (N_7038,N_6236,N_6147);
or U7039 (N_7039,N_6772,N_6858);
and U7040 (N_7040,N_6212,N_6763);
nor U7041 (N_7041,N_6538,N_6478);
or U7042 (N_7042,N_6095,N_6967);
nor U7043 (N_7043,N_6613,N_6657);
nor U7044 (N_7044,N_6558,N_6387);
nand U7045 (N_7045,N_6674,N_6446);
xor U7046 (N_7046,N_6962,N_6381);
or U7047 (N_7047,N_6269,N_6900);
xor U7048 (N_7048,N_6217,N_6177);
or U7049 (N_7049,N_6709,N_6376);
nand U7050 (N_7050,N_6285,N_6592);
or U7051 (N_7051,N_6468,N_6903);
and U7052 (N_7052,N_6812,N_6039);
nor U7053 (N_7053,N_6204,N_6091);
nor U7054 (N_7054,N_6626,N_6320);
xnor U7055 (N_7055,N_6295,N_6711);
nor U7056 (N_7056,N_6825,N_6422);
nor U7057 (N_7057,N_6839,N_6106);
and U7058 (N_7058,N_6507,N_6906);
nor U7059 (N_7059,N_6627,N_6065);
xor U7060 (N_7060,N_6745,N_6525);
nor U7061 (N_7061,N_6447,N_6378);
and U7062 (N_7062,N_6304,N_6848);
and U7063 (N_7063,N_6276,N_6027);
and U7064 (N_7064,N_6896,N_6250);
xnor U7065 (N_7065,N_6944,N_6136);
or U7066 (N_7066,N_6976,N_6609);
nand U7067 (N_7067,N_6154,N_6390);
nor U7068 (N_7068,N_6803,N_6856);
nor U7069 (N_7069,N_6157,N_6552);
nor U7070 (N_7070,N_6122,N_6637);
nor U7071 (N_7071,N_6949,N_6201);
nand U7072 (N_7072,N_6749,N_6145);
xor U7073 (N_7073,N_6913,N_6193);
or U7074 (N_7074,N_6403,N_6286);
and U7075 (N_7075,N_6046,N_6901);
nor U7076 (N_7076,N_6729,N_6142);
nand U7077 (N_7077,N_6853,N_6547);
nor U7078 (N_7078,N_6611,N_6882);
xnor U7079 (N_7079,N_6194,N_6683);
and U7080 (N_7080,N_6678,N_6570);
nor U7081 (N_7081,N_6871,N_6564);
nor U7082 (N_7082,N_6053,N_6412);
or U7083 (N_7083,N_6211,N_6851);
nand U7084 (N_7084,N_6981,N_6866);
nor U7085 (N_7085,N_6453,N_6777);
xor U7086 (N_7086,N_6009,N_6503);
and U7087 (N_7087,N_6041,N_6079);
nand U7088 (N_7088,N_6028,N_6228);
or U7089 (N_7089,N_6884,N_6089);
nand U7090 (N_7090,N_6952,N_6363);
nand U7091 (N_7091,N_6060,N_6076);
nor U7092 (N_7092,N_6912,N_6030);
xor U7093 (N_7093,N_6826,N_6413);
or U7094 (N_7094,N_6681,N_6072);
xnor U7095 (N_7095,N_6441,N_6530);
nor U7096 (N_7096,N_6834,N_6162);
nand U7097 (N_7097,N_6580,N_6245);
nand U7098 (N_7098,N_6215,N_6277);
or U7099 (N_7099,N_6818,N_6672);
or U7100 (N_7100,N_6401,N_6649);
or U7101 (N_7101,N_6303,N_6038);
or U7102 (N_7102,N_6813,N_6577);
nand U7103 (N_7103,N_6721,N_6890);
or U7104 (N_7104,N_6362,N_6400);
nor U7105 (N_7105,N_6827,N_6671);
xor U7106 (N_7106,N_6237,N_6894);
and U7107 (N_7107,N_6461,N_6751);
or U7108 (N_7108,N_6593,N_6379);
and U7109 (N_7109,N_6020,N_6659);
nor U7110 (N_7110,N_6684,N_6275);
and U7111 (N_7111,N_6980,N_6126);
and U7112 (N_7112,N_6752,N_6954);
and U7113 (N_7113,N_6759,N_6569);
xor U7114 (N_7114,N_6597,N_6828);
or U7115 (N_7115,N_6801,N_6975);
xor U7116 (N_7116,N_6537,N_6271);
nor U7117 (N_7117,N_6113,N_6621);
nor U7118 (N_7118,N_6937,N_6062);
and U7119 (N_7119,N_6874,N_6596);
nand U7120 (N_7120,N_6778,N_6452);
xor U7121 (N_7121,N_6058,N_6052);
nand U7122 (N_7122,N_6947,N_6776);
and U7123 (N_7123,N_6377,N_6210);
nor U7124 (N_7124,N_6226,N_6425);
nand U7125 (N_7125,N_6111,N_6370);
nand U7126 (N_7126,N_6491,N_6444);
nor U7127 (N_7127,N_6862,N_6940);
and U7128 (N_7128,N_6270,N_6492);
nand U7129 (N_7129,N_6760,N_6652);
nand U7130 (N_7130,N_6417,N_6734);
and U7131 (N_7131,N_6831,N_6790);
and U7132 (N_7132,N_6647,N_6159);
xnor U7133 (N_7133,N_6893,N_6830);
or U7134 (N_7134,N_6883,N_6435);
nand U7135 (N_7135,N_6302,N_6057);
nand U7136 (N_7136,N_6249,N_6914);
and U7137 (N_7137,N_6521,N_6996);
nor U7138 (N_7138,N_6483,N_6727);
nor U7139 (N_7139,N_6523,N_6287);
nand U7140 (N_7140,N_6040,N_6833);
or U7141 (N_7141,N_6765,N_6368);
nor U7142 (N_7142,N_6710,N_6587);
or U7143 (N_7143,N_6667,N_6187);
xor U7144 (N_7144,N_6129,N_6802);
nand U7145 (N_7145,N_6518,N_6104);
nand U7146 (N_7146,N_6702,N_6829);
nor U7147 (N_7147,N_6156,N_6023);
nand U7148 (N_7148,N_6308,N_6574);
and U7149 (N_7149,N_6029,N_6207);
xor U7150 (N_7150,N_6714,N_6179);
and U7151 (N_7151,N_6465,N_6118);
nor U7152 (N_7152,N_6432,N_6941);
nor U7153 (N_7153,N_6965,N_6445);
xor U7154 (N_7154,N_6169,N_6725);
nor U7155 (N_7155,N_6664,N_6791);
or U7156 (N_7156,N_6520,N_6730);
xor U7157 (N_7157,N_6353,N_6757);
and U7158 (N_7158,N_6402,N_6408);
nand U7159 (N_7159,N_6988,N_6679);
nand U7160 (N_7160,N_6566,N_6472);
and U7161 (N_7161,N_6423,N_6151);
nand U7162 (N_7162,N_6232,N_6589);
or U7163 (N_7163,N_6950,N_6563);
or U7164 (N_7164,N_6731,N_6257);
or U7165 (N_7165,N_6407,N_6867);
nand U7166 (N_7166,N_6634,N_6620);
nor U7167 (N_7167,N_6037,N_6296);
nand U7168 (N_7168,N_6094,N_6733);
xnor U7169 (N_7169,N_6280,N_6183);
xnor U7170 (N_7170,N_6810,N_6234);
or U7171 (N_7171,N_6910,N_6054);
and U7172 (N_7172,N_6330,N_6636);
xor U7173 (N_7173,N_6253,N_6255);
nor U7174 (N_7174,N_6498,N_6220);
and U7175 (N_7175,N_6568,N_6392);
or U7176 (N_7176,N_6097,N_6265);
nand U7177 (N_7177,N_6860,N_6123);
nor U7178 (N_7178,N_6281,N_6336);
nand U7179 (N_7179,N_6063,N_6093);
or U7180 (N_7180,N_6279,N_6875);
nand U7181 (N_7181,N_6656,N_6496);
and U7182 (N_7182,N_6015,N_6956);
or U7183 (N_7183,N_6102,N_6986);
and U7184 (N_7184,N_6529,N_6554);
or U7185 (N_7185,N_6662,N_6968);
or U7186 (N_7186,N_6886,N_6992);
xnor U7187 (N_7187,N_6259,N_6511);
and U7188 (N_7188,N_6036,N_6532);
and U7189 (N_7189,N_6092,N_6930);
nor U7190 (N_7190,N_6148,N_6604);
and U7191 (N_7191,N_6533,N_6779);
and U7192 (N_7192,N_6132,N_6443);
or U7193 (N_7193,N_6294,N_6691);
xnor U7194 (N_7194,N_6809,N_6514);
nor U7195 (N_7195,N_6859,N_6824);
nand U7196 (N_7196,N_6274,N_6324);
xnor U7197 (N_7197,N_6723,N_6476);
nand U7198 (N_7198,N_6562,N_6945);
and U7199 (N_7199,N_6099,N_6224);
xor U7200 (N_7200,N_6431,N_6556);
and U7201 (N_7201,N_6137,N_6042);
nor U7202 (N_7202,N_6354,N_6876);
or U7203 (N_7203,N_6499,N_6134);
xnor U7204 (N_7204,N_6789,N_6116);
nor U7205 (N_7205,N_6488,N_6963);
or U7206 (N_7206,N_6513,N_6966);
nor U7207 (N_7207,N_6541,N_6318);
nand U7208 (N_7208,N_6202,N_6891);
nand U7209 (N_7209,N_6524,N_6384);
xnor U7210 (N_7210,N_6805,N_6619);
nor U7211 (N_7211,N_6497,N_6645);
xnor U7212 (N_7212,N_6773,N_6206);
nand U7213 (N_7213,N_6689,N_6832);
and U7214 (N_7214,N_6473,N_6291);
and U7215 (N_7215,N_6821,N_6388);
and U7216 (N_7216,N_6675,N_6424);
xnor U7217 (N_7217,N_6305,N_6462);
or U7218 (N_7218,N_6048,N_6050);
nand U7219 (N_7219,N_6133,N_6077);
nor U7220 (N_7220,N_6138,N_6326);
and U7221 (N_7221,N_6925,N_6395);
and U7222 (N_7222,N_6084,N_6034);
and U7223 (N_7223,N_6292,N_6567);
nor U7224 (N_7224,N_6045,N_6951);
xor U7225 (N_7225,N_6756,N_6155);
nand U7226 (N_7226,N_6317,N_6528);
nand U7227 (N_7227,N_6241,N_6289);
nor U7228 (N_7228,N_6258,N_6707);
nand U7229 (N_7229,N_6991,N_6300);
nor U7230 (N_7230,N_6333,N_6850);
nand U7231 (N_7231,N_6722,N_6744);
or U7232 (N_7232,N_6244,N_6895);
xnor U7233 (N_7233,N_6660,N_6650);
or U7234 (N_7234,N_6440,N_6316);
nor U7235 (N_7235,N_6124,N_6261);
or U7236 (N_7236,N_6855,N_6780);
or U7237 (N_7237,N_6835,N_6819);
nor U7238 (N_7238,N_6168,N_6219);
xnor U7239 (N_7239,N_6586,N_6315);
nor U7240 (N_7240,N_6854,N_6227);
nand U7241 (N_7241,N_6495,N_6439);
and U7242 (N_7242,N_6663,N_6284);
nor U7243 (N_7243,N_6214,N_6666);
and U7244 (N_7244,N_6069,N_6939);
and U7245 (N_7245,N_6229,N_6414);
xor U7246 (N_7246,N_6869,N_6487);
nand U7247 (N_7247,N_6190,N_6373);
nor U7248 (N_7248,N_6706,N_6175);
and U7249 (N_7249,N_6358,N_6557);
xnor U7250 (N_7250,N_6021,N_6357);
xor U7251 (N_7251,N_6238,N_6669);
and U7252 (N_7252,N_6033,N_6017);
xor U7253 (N_7253,N_6141,N_6782);
and U7254 (N_7254,N_6203,N_6999);
xor U7255 (N_7255,N_6615,N_6716);
xnor U7256 (N_7256,N_6160,N_6885);
xnor U7257 (N_7257,N_6135,N_6127);
xnor U7258 (N_7258,N_6512,N_6648);
or U7259 (N_7259,N_6121,N_6852);
or U7260 (N_7260,N_6724,N_6209);
nor U7261 (N_7261,N_6908,N_6536);
nand U7262 (N_7262,N_6369,N_6008);
xor U7263 (N_7263,N_6251,N_6849);
nor U7264 (N_7264,N_6463,N_6125);
xnor U7265 (N_7265,N_6139,N_6920);
nand U7266 (N_7266,N_6486,N_6911);
nor U7267 (N_7267,N_6485,N_6708);
nand U7268 (N_7268,N_6973,N_6522);
nor U7269 (N_7269,N_6355,N_6924);
or U7270 (N_7270,N_6612,N_6051);
nand U7271 (N_7271,N_6785,N_6323);
and U7272 (N_7272,N_6011,N_6605);
xnor U7273 (N_7273,N_6365,N_6936);
nand U7274 (N_7274,N_6682,N_6233);
or U7275 (N_7275,N_6712,N_6916);
nor U7276 (N_7276,N_6591,N_6748);
nand U7277 (N_7277,N_6128,N_6519);
xnor U7278 (N_7278,N_6927,N_6510);
nand U7279 (N_7279,N_6205,N_6565);
and U7280 (N_7280,N_6075,N_6459);
xnor U7281 (N_7281,N_6366,N_6929);
and U7282 (N_7282,N_6971,N_6942);
nor U7283 (N_7283,N_6032,N_6685);
xnor U7284 (N_7284,N_6583,N_6195);
and U7285 (N_7285,N_6775,N_6979);
nand U7286 (N_7286,N_6310,N_6359);
and U7287 (N_7287,N_6616,N_6598);
nor U7288 (N_7288,N_6080,N_6736);
or U7289 (N_7289,N_6761,N_6614);
nand U7290 (N_7290,N_6467,N_6770);
or U7291 (N_7291,N_6517,N_6016);
nor U7292 (N_7292,N_6665,N_6429);
xnor U7293 (N_7293,N_6559,N_6546);
nor U7294 (N_7294,N_6350,N_6961);
nor U7295 (N_7295,N_6332,N_6396);
xnor U7296 (N_7296,N_6345,N_6571);
and U7297 (N_7297,N_6256,N_6083);
nor U7298 (N_7298,N_6576,N_6668);
nand U7299 (N_7299,N_6426,N_6055);
xnor U7300 (N_7300,N_6673,N_6638);
and U7301 (N_7301,N_6888,N_6977);
or U7302 (N_7302,N_6166,N_6242);
nor U7303 (N_7303,N_6918,N_6235);
and U7304 (N_7304,N_6306,N_6715);
xor U7305 (N_7305,N_6692,N_6293);
xnor U7306 (N_7306,N_6152,N_6347);
xnor U7307 (N_7307,N_6700,N_6098);
or U7308 (N_7308,N_6987,N_6264);
xnor U7309 (N_7309,N_6516,N_6184);
nand U7310 (N_7310,N_6625,N_6225);
xnor U7311 (N_7311,N_6909,N_6696);
xnor U7312 (N_7312,N_6380,N_6278);
nand U7313 (N_7313,N_6766,N_6501);
nor U7314 (N_7314,N_6405,N_6254);
xor U7315 (N_7315,N_6594,N_6985);
and U7316 (N_7316,N_6240,N_6998);
nand U7317 (N_7317,N_6170,N_6340);
and U7318 (N_7318,N_6694,N_6031);
and U7319 (N_7319,N_6337,N_6197);
or U7320 (N_7320,N_6630,N_6792);
xor U7321 (N_7321,N_6438,N_6120);
nand U7322 (N_7322,N_6013,N_6732);
and U7323 (N_7323,N_6252,N_6535);
nand U7324 (N_7324,N_6658,N_6319);
xnor U7325 (N_7325,N_6272,N_6181);
nor U7326 (N_7326,N_6470,N_6820);
or U7327 (N_7327,N_6329,N_6356);
and U7328 (N_7328,N_6167,N_6301);
nand U7329 (N_7329,N_6982,N_6865);
and U7330 (N_7330,N_6561,N_6798);
xnor U7331 (N_7331,N_6068,N_6633);
or U7332 (N_7332,N_6059,N_6153);
xnor U7333 (N_7333,N_6282,N_6464);
xnor U7334 (N_7334,N_6655,N_6793);
and U7335 (N_7335,N_6795,N_6448);
nand U7336 (N_7336,N_6907,N_6974);
nand U7337 (N_7337,N_6364,N_6505);
or U7338 (N_7338,N_6575,N_6845);
nor U7339 (N_7339,N_6905,N_6807);
or U7340 (N_7340,N_6001,N_6703);
nor U7341 (N_7341,N_6836,N_6840);
nand U7342 (N_7342,N_6640,N_6343);
or U7343 (N_7343,N_6188,N_6631);
nor U7344 (N_7344,N_6972,N_6010);
nor U7345 (N_7345,N_6398,N_6946);
nand U7346 (N_7346,N_6739,N_6603);
or U7347 (N_7347,N_6391,N_6957);
xnor U7348 (N_7348,N_6196,N_6107);
and U7349 (N_7349,N_6781,N_6322);
or U7350 (N_7350,N_6044,N_6935);
and U7351 (N_7351,N_6984,N_6573);
xnor U7352 (N_7352,N_6466,N_6171);
nand U7353 (N_7353,N_6230,N_6312);
and U7354 (N_7354,N_6349,N_6103);
xnor U7355 (N_7355,N_6457,N_6144);
xnor U7356 (N_7356,N_6644,N_6515);
xnor U7357 (N_7357,N_6796,N_6474);
or U7358 (N_7358,N_6794,N_6460);
and U7359 (N_7359,N_6437,N_6728);
nor U7360 (N_7360,N_6185,N_6553);
or U7361 (N_7361,N_6455,N_6105);
xor U7362 (N_7362,N_6026,N_6416);
nand U7363 (N_7363,N_6014,N_6676);
nor U7364 (N_7364,N_6313,N_6191);
xnor U7365 (N_7365,N_6964,N_6071);
nand U7366 (N_7366,N_6374,N_6247);
xor U7367 (N_7367,N_6718,N_6953);
or U7368 (N_7368,N_6297,N_6003);
nor U7369 (N_7369,N_6680,N_6786);
nand U7370 (N_7370,N_6878,N_6231);
xor U7371 (N_7371,N_6877,N_6622);
nand U7372 (N_7372,N_6411,N_6698);
xor U7373 (N_7373,N_6582,N_6004);
or U7374 (N_7374,N_6600,N_6983);
nor U7375 (N_7375,N_6837,N_6506);
nand U7376 (N_7376,N_6007,N_6218);
nand U7377 (N_7377,N_6857,N_6442);
and U7378 (N_7378,N_6970,N_6165);
and U7379 (N_7379,N_6022,N_6420);
or U7380 (N_7380,N_6067,N_6814);
nor U7381 (N_7381,N_6049,N_6960);
or U7382 (N_7382,N_6509,N_6342);
nand U7383 (N_7383,N_6726,N_6933);
xor U7384 (N_7384,N_6579,N_6815);
and U7385 (N_7385,N_6754,N_6601);
or U7386 (N_7386,N_6747,N_6263);
and U7387 (N_7387,N_6490,N_6078);
xor U7388 (N_7388,N_6738,N_6959);
or U7389 (N_7389,N_6607,N_6131);
nor U7390 (N_7390,N_6267,N_6892);
nand U7391 (N_7391,N_6938,N_6389);
xnor U7392 (N_7392,N_6870,N_6012);
or U7393 (N_7393,N_6096,N_6713);
nand U7394 (N_7394,N_6804,N_6213);
and U7395 (N_7395,N_6719,N_6743);
nor U7396 (N_7396,N_6843,N_6688);
nand U7397 (N_7397,N_6182,N_6436);
nor U7398 (N_7398,N_6299,N_6086);
and U7399 (N_7399,N_6762,N_6243);
and U7400 (N_7400,N_6887,N_6771);
xnor U7401 (N_7401,N_6025,N_6585);
and U7402 (N_7402,N_6341,N_6695);
and U7403 (N_7403,N_6923,N_6639);
xor U7404 (N_7404,N_6881,N_6764);
nand U7405 (N_7405,N_6921,N_6481);
xor U7406 (N_7406,N_6578,N_6897);
or U7407 (N_7407,N_6361,N_6061);
or U7408 (N_7408,N_6115,N_6449);
or U7409 (N_7409,N_6180,N_6993);
nor U7410 (N_7410,N_6418,N_6783);
or U7411 (N_7411,N_6100,N_6409);
or U7412 (N_7412,N_6172,N_6189);
xnor U7413 (N_7413,N_6872,N_6548);
xnor U7414 (N_7414,N_6797,N_6430);
xnor U7415 (N_7415,N_6978,N_6428);
and U7416 (N_7416,N_6163,N_6590);
nand U7417 (N_7417,N_6690,N_6344);
nor U7418 (N_7418,N_6130,N_6847);
nand U7419 (N_7419,N_6024,N_6158);
xor U7420 (N_7420,N_6800,N_6216);
nor U7421 (N_7421,N_6581,N_6551);
nor U7422 (N_7422,N_6427,N_6651);
nand U7423 (N_7423,N_6919,N_6742);
xnor U7424 (N_7424,N_6768,N_6469);
or U7425 (N_7425,N_6686,N_6697);
or U7426 (N_7426,N_6266,N_6531);
and U7427 (N_7427,N_6372,N_6995);
nand U7428 (N_7428,N_6846,N_6624);
xnor U7429 (N_7429,N_6382,N_6262);
nor U7430 (N_7430,N_6248,N_6117);
or U7431 (N_7431,N_6502,N_6955);
nor U7432 (N_7432,N_6618,N_6348);
xnor U7433 (N_7433,N_6841,N_6451);
xnor U7434 (N_7434,N_6994,N_6543);
xor U7435 (N_7435,N_6174,N_6880);
nand U7436 (N_7436,N_6200,N_6629);
or U7437 (N_7437,N_6642,N_6352);
or U7438 (N_7438,N_6454,N_6922);
or U7439 (N_7439,N_6989,N_6737);
and U7440 (N_7440,N_6371,N_6602);
or U7441 (N_7441,N_6899,N_6808);
and U7442 (N_7442,N_6806,N_6753);
xnor U7443 (N_7443,N_6397,N_6863);
or U7444 (N_7444,N_6741,N_6043);
xor U7445 (N_7445,N_6101,N_6081);
xor U7446 (N_7446,N_6788,N_6898);
nor U7447 (N_7447,N_6339,N_6321);
xor U7448 (N_7448,N_6822,N_6208);
nor U7449 (N_7449,N_6494,N_6335);
or U7450 (N_7450,N_6817,N_6221);
and U7451 (N_7451,N_6699,N_6006);
xor U7452 (N_7452,N_6799,N_6769);
or U7453 (N_7453,N_6112,N_6489);
xor U7454 (N_7454,N_6056,N_6928);
or U7455 (N_7455,N_6199,N_6327);
or U7456 (N_7456,N_6717,N_6735);
nor U7457 (N_7457,N_6572,N_6018);
and U7458 (N_7458,N_6948,N_6002);
or U7459 (N_7459,N_6173,N_6351);
or U7460 (N_7460,N_6164,N_6338);
and U7461 (N_7461,N_6588,N_6223);
nor U7462 (N_7462,N_6606,N_6273);
and U7463 (N_7463,N_6066,N_6861);
nor U7464 (N_7464,N_6109,N_6902);
xnor U7465 (N_7465,N_6331,N_6990);
xor U7466 (N_7466,N_6087,N_6260);
and U7467 (N_7467,N_6838,N_6309);
or U7468 (N_7468,N_6433,N_6599);
xor U7469 (N_7469,N_6480,N_6787);
or U7470 (N_7470,N_6879,N_6150);
and U7471 (N_7471,N_6493,N_6088);
or U7472 (N_7472,N_6070,N_6555);
xnor U7473 (N_7473,N_6222,N_6198);
or U7474 (N_7474,N_6421,N_6767);
and U7475 (N_7475,N_6632,N_6823);
and U7476 (N_7476,N_6475,N_6450);
nand U7477 (N_7477,N_6504,N_6670);
xnor U7478 (N_7478,N_6508,N_6926);
or U7479 (N_7479,N_6635,N_6386);
nor U7480 (N_7480,N_6943,N_6419);
nand U7481 (N_7481,N_6074,N_6584);
or U7482 (N_7482,N_6119,N_6000);
or U7483 (N_7483,N_6842,N_6186);
or U7484 (N_7484,N_6740,N_6544);
or U7485 (N_7485,N_6334,N_6346);
xnor U7486 (N_7486,N_6844,N_6623);
or U7487 (N_7487,N_6192,N_6410);
nor U7488 (N_7488,N_6701,N_6595);
xor U7489 (N_7489,N_6641,N_6750);
nand U7490 (N_7490,N_6239,N_6550);
and U7491 (N_7491,N_6399,N_6654);
nand U7492 (N_7492,N_6917,N_6307);
nor U7493 (N_7493,N_6653,N_6560);
nand U7494 (N_7494,N_6458,N_6549);
nand U7495 (N_7495,N_6367,N_6082);
xnor U7496 (N_7496,N_6161,N_6774);
and U7497 (N_7497,N_6527,N_6915);
xor U7498 (N_7498,N_6283,N_6114);
xor U7499 (N_7499,N_6617,N_6661);
and U7500 (N_7500,N_6640,N_6737);
and U7501 (N_7501,N_6515,N_6683);
or U7502 (N_7502,N_6695,N_6070);
and U7503 (N_7503,N_6659,N_6241);
and U7504 (N_7504,N_6055,N_6748);
or U7505 (N_7505,N_6999,N_6901);
xnor U7506 (N_7506,N_6226,N_6703);
nand U7507 (N_7507,N_6340,N_6188);
or U7508 (N_7508,N_6659,N_6053);
nor U7509 (N_7509,N_6133,N_6976);
nor U7510 (N_7510,N_6382,N_6792);
nor U7511 (N_7511,N_6657,N_6033);
or U7512 (N_7512,N_6724,N_6737);
nand U7513 (N_7513,N_6743,N_6968);
nand U7514 (N_7514,N_6538,N_6700);
or U7515 (N_7515,N_6735,N_6861);
nor U7516 (N_7516,N_6336,N_6122);
or U7517 (N_7517,N_6151,N_6328);
xnor U7518 (N_7518,N_6690,N_6197);
or U7519 (N_7519,N_6315,N_6714);
xor U7520 (N_7520,N_6895,N_6192);
xor U7521 (N_7521,N_6488,N_6113);
xor U7522 (N_7522,N_6152,N_6141);
xnor U7523 (N_7523,N_6051,N_6565);
or U7524 (N_7524,N_6139,N_6960);
nand U7525 (N_7525,N_6511,N_6810);
or U7526 (N_7526,N_6375,N_6465);
xor U7527 (N_7527,N_6151,N_6239);
or U7528 (N_7528,N_6240,N_6255);
or U7529 (N_7529,N_6999,N_6750);
xor U7530 (N_7530,N_6900,N_6507);
xor U7531 (N_7531,N_6101,N_6305);
nor U7532 (N_7532,N_6991,N_6209);
and U7533 (N_7533,N_6250,N_6362);
and U7534 (N_7534,N_6411,N_6978);
nand U7535 (N_7535,N_6417,N_6860);
nand U7536 (N_7536,N_6558,N_6563);
and U7537 (N_7537,N_6721,N_6234);
nor U7538 (N_7538,N_6027,N_6032);
nand U7539 (N_7539,N_6066,N_6633);
xor U7540 (N_7540,N_6502,N_6470);
xnor U7541 (N_7541,N_6856,N_6028);
xnor U7542 (N_7542,N_6331,N_6750);
nor U7543 (N_7543,N_6099,N_6776);
or U7544 (N_7544,N_6330,N_6612);
nor U7545 (N_7545,N_6971,N_6393);
nor U7546 (N_7546,N_6711,N_6390);
nand U7547 (N_7547,N_6575,N_6390);
or U7548 (N_7548,N_6513,N_6036);
nand U7549 (N_7549,N_6696,N_6264);
nand U7550 (N_7550,N_6343,N_6614);
or U7551 (N_7551,N_6732,N_6791);
and U7552 (N_7552,N_6363,N_6303);
and U7553 (N_7553,N_6683,N_6238);
and U7554 (N_7554,N_6465,N_6124);
nand U7555 (N_7555,N_6637,N_6146);
xor U7556 (N_7556,N_6619,N_6020);
and U7557 (N_7557,N_6623,N_6481);
xor U7558 (N_7558,N_6166,N_6196);
nor U7559 (N_7559,N_6003,N_6138);
nor U7560 (N_7560,N_6970,N_6398);
xnor U7561 (N_7561,N_6058,N_6020);
nand U7562 (N_7562,N_6913,N_6151);
nor U7563 (N_7563,N_6334,N_6300);
and U7564 (N_7564,N_6661,N_6450);
or U7565 (N_7565,N_6001,N_6418);
xnor U7566 (N_7566,N_6381,N_6889);
nor U7567 (N_7567,N_6183,N_6698);
nand U7568 (N_7568,N_6418,N_6707);
and U7569 (N_7569,N_6950,N_6245);
or U7570 (N_7570,N_6632,N_6503);
xnor U7571 (N_7571,N_6944,N_6825);
nand U7572 (N_7572,N_6405,N_6303);
or U7573 (N_7573,N_6800,N_6398);
nor U7574 (N_7574,N_6783,N_6591);
or U7575 (N_7575,N_6403,N_6256);
and U7576 (N_7576,N_6934,N_6939);
or U7577 (N_7577,N_6663,N_6905);
xor U7578 (N_7578,N_6801,N_6320);
nand U7579 (N_7579,N_6882,N_6793);
and U7580 (N_7580,N_6883,N_6226);
or U7581 (N_7581,N_6582,N_6202);
or U7582 (N_7582,N_6371,N_6818);
and U7583 (N_7583,N_6386,N_6770);
nand U7584 (N_7584,N_6307,N_6325);
nor U7585 (N_7585,N_6040,N_6188);
nor U7586 (N_7586,N_6500,N_6823);
nand U7587 (N_7587,N_6002,N_6813);
or U7588 (N_7588,N_6957,N_6160);
or U7589 (N_7589,N_6144,N_6394);
nand U7590 (N_7590,N_6535,N_6917);
and U7591 (N_7591,N_6361,N_6844);
nor U7592 (N_7592,N_6575,N_6987);
xor U7593 (N_7593,N_6921,N_6651);
or U7594 (N_7594,N_6763,N_6069);
nand U7595 (N_7595,N_6081,N_6413);
xor U7596 (N_7596,N_6852,N_6619);
xor U7597 (N_7597,N_6944,N_6148);
and U7598 (N_7598,N_6193,N_6243);
xnor U7599 (N_7599,N_6606,N_6352);
xor U7600 (N_7600,N_6176,N_6618);
nor U7601 (N_7601,N_6040,N_6330);
or U7602 (N_7602,N_6909,N_6138);
and U7603 (N_7603,N_6851,N_6249);
nand U7604 (N_7604,N_6338,N_6865);
or U7605 (N_7605,N_6712,N_6438);
or U7606 (N_7606,N_6385,N_6319);
nand U7607 (N_7607,N_6840,N_6417);
xnor U7608 (N_7608,N_6582,N_6025);
or U7609 (N_7609,N_6313,N_6146);
nand U7610 (N_7610,N_6968,N_6618);
and U7611 (N_7611,N_6875,N_6037);
or U7612 (N_7612,N_6565,N_6054);
xnor U7613 (N_7613,N_6642,N_6728);
and U7614 (N_7614,N_6764,N_6501);
or U7615 (N_7615,N_6751,N_6529);
or U7616 (N_7616,N_6118,N_6899);
xor U7617 (N_7617,N_6136,N_6102);
or U7618 (N_7618,N_6412,N_6326);
nor U7619 (N_7619,N_6547,N_6401);
nand U7620 (N_7620,N_6458,N_6290);
or U7621 (N_7621,N_6937,N_6011);
nor U7622 (N_7622,N_6408,N_6104);
nor U7623 (N_7623,N_6298,N_6270);
and U7624 (N_7624,N_6154,N_6073);
xnor U7625 (N_7625,N_6287,N_6332);
xor U7626 (N_7626,N_6736,N_6348);
nand U7627 (N_7627,N_6672,N_6317);
or U7628 (N_7628,N_6988,N_6107);
or U7629 (N_7629,N_6543,N_6260);
nand U7630 (N_7630,N_6716,N_6056);
xnor U7631 (N_7631,N_6179,N_6265);
xnor U7632 (N_7632,N_6867,N_6959);
or U7633 (N_7633,N_6975,N_6228);
nor U7634 (N_7634,N_6217,N_6148);
xor U7635 (N_7635,N_6796,N_6083);
xnor U7636 (N_7636,N_6234,N_6456);
or U7637 (N_7637,N_6225,N_6386);
or U7638 (N_7638,N_6071,N_6141);
or U7639 (N_7639,N_6729,N_6260);
or U7640 (N_7640,N_6816,N_6815);
and U7641 (N_7641,N_6871,N_6767);
or U7642 (N_7642,N_6559,N_6319);
nor U7643 (N_7643,N_6844,N_6566);
xor U7644 (N_7644,N_6819,N_6545);
or U7645 (N_7645,N_6643,N_6188);
nand U7646 (N_7646,N_6855,N_6498);
nand U7647 (N_7647,N_6432,N_6452);
nor U7648 (N_7648,N_6976,N_6577);
nand U7649 (N_7649,N_6707,N_6080);
or U7650 (N_7650,N_6559,N_6253);
nand U7651 (N_7651,N_6092,N_6761);
xor U7652 (N_7652,N_6600,N_6851);
xnor U7653 (N_7653,N_6959,N_6764);
or U7654 (N_7654,N_6476,N_6057);
and U7655 (N_7655,N_6566,N_6034);
or U7656 (N_7656,N_6770,N_6132);
xnor U7657 (N_7657,N_6600,N_6083);
xnor U7658 (N_7658,N_6047,N_6412);
nor U7659 (N_7659,N_6086,N_6552);
or U7660 (N_7660,N_6355,N_6420);
or U7661 (N_7661,N_6529,N_6257);
or U7662 (N_7662,N_6599,N_6940);
xor U7663 (N_7663,N_6683,N_6622);
nor U7664 (N_7664,N_6112,N_6397);
or U7665 (N_7665,N_6654,N_6423);
or U7666 (N_7666,N_6770,N_6598);
and U7667 (N_7667,N_6349,N_6662);
nor U7668 (N_7668,N_6569,N_6326);
nand U7669 (N_7669,N_6031,N_6199);
and U7670 (N_7670,N_6194,N_6587);
and U7671 (N_7671,N_6302,N_6946);
nand U7672 (N_7672,N_6825,N_6429);
nand U7673 (N_7673,N_6120,N_6695);
nor U7674 (N_7674,N_6908,N_6887);
nor U7675 (N_7675,N_6581,N_6181);
or U7676 (N_7676,N_6799,N_6982);
nor U7677 (N_7677,N_6540,N_6842);
and U7678 (N_7678,N_6150,N_6410);
and U7679 (N_7679,N_6675,N_6257);
xnor U7680 (N_7680,N_6279,N_6991);
nand U7681 (N_7681,N_6412,N_6124);
and U7682 (N_7682,N_6397,N_6415);
nand U7683 (N_7683,N_6118,N_6759);
or U7684 (N_7684,N_6047,N_6638);
xor U7685 (N_7685,N_6492,N_6539);
xor U7686 (N_7686,N_6736,N_6167);
nand U7687 (N_7687,N_6506,N_6286);
nand U7688 (N_7688,N_6971,N_6396);
and U7689 (N_7689,N_6332,N_6054);
or U7690 (N_7690,N_6997,N_6455);
xnor U7691 (N_7691,N_6738,N_6701);
or U7692 (N_7692,N_6245,N_6814);
and U7693 (N_7693,N_6435,N_6774);
xnor U7694 (N_7694,N_6843,N_6347);
xor U7695 (N_7695,N_6008,N_6504);
and U7696 (N_7696,N_6836,N_6593);
nor U7697 (N_7697,N_6791,N_6159);
nor U7698 (N_7698,N_6869,N_6077);
nor U7699 (N_7699,N_6761,N_6890);
and U7700 (N_7700,N_6171,N_6231);
xor U7701 (N_7701,N_6981,N_6704);
nand U7702 (N_7702,N_6478,N_6819);
xor U7703 (N_7703,N_6349,N_6536);
nand U7704 (N_7704,N_6874,N_6250);
or U7705 (N_7705,N_6994,N_6018);
nand U7706 (N_7706,N_6467,N_6080);
nor U7707 (N_7707,N_6569,N_6980);
nor U7708 (N_7708,N_6517,N_6238);
xor U7709 (N_7709,N_6538,N_6172);
and U7710 (N_7710,N_6360,N_6246);
nor U7711 (N_7711,N_6489,N_6986);
and U7712 (N_7712,N_6311,N_6223);
or U7713 (N_7713,N_6135,N_6524);
nor U7714 (N_7714,N_6315,N_6227);
and U7715 (N_7715,N_6696,N_6117);
or U7716 (N_7716,N_6340,N_6546);
and U7717 (N_7717,N_6320,N_6313);
xnor U7718 (N_7718,N_6277,N_6562);
nor U7719 (N_7719,N_6292,N_6534);
xnor U7720 (N_7720,N_6023,N_6547);
xor U7721 (N_7721,N_6640,N_6542);
nor U7722 (N_7722,N_6345,N_6568);
nand U7723 (N_7723,N_6638,N_6924);
xor U7724 (N_7724,N_6520,N_6891);
xor U7725 (N_7725,N_6754,N_6622);
nor U7726 (N_7726,N_6656,N_6594);
nand U7727 (N_7727,N_6601,N_6068);
xnor U7728 (N_7728,N_6121,N_6064);
nor U7729 (N_7729,N_6295,N_6832);
nor U7730 (N_7730,N_6338,N_6917);
xor U7731 (N_7731,N_6705,N_6473);
nor U7732 (N_7732,N_6798,N_6186);
and U7733 (N_7733,N_6701,N_6792);
nor U7734 (N_7734,N_6063,N_6936);
or U7735 (N_7735,N_6908,N_6143);
nor U7736 (N_7736,N_6883,N_6863);
or U7737 (N_7737,N_6476,N_6657);
and U7738 (N_7738,N_6066,N_6828);
nor U7739 (N_7739,N_6973,N_6868);
and U7740 (N_7740,N_6202,N_6917);
or U7741 (N_7741,N_6064,N_6473);
or U7742 (N_7742,N_6887,N_6304);
nand U7743 (N_7743,N_6186,N_6449);
nor U7744 (N_7744,N_6879,N_6677);
and U7745 (N_7745,N_6142,N_6448);
or U7746 (N_7746,N_6553,N_6928);
or U7747 (N_7747,N_6587,N_6530);
xnor U7748 (N_7748,N_6533,N_6825);
xor U7749 (N_7749,N_6096,N_6952);
and U7750 (N_7750,N_6155,N_6047);
nand U7751 (N_7751,N_6621,N_6546);
xnor U7752 (N_7752,N_6335,N_6959);
nand U7753 (N_7753,N_6991,N_6098);
nor U7754 (N_7754,N_6101,N_6733);
xor U7755 (N_7755,N_6000,N_6022);
nand U7756 (N_7756,N_6599,N_6894);
nand U7757 (N_7757,N_6024,N_6915);
nor U7758 (N_7758,N_6034,N_6892);
or U7759 (N_7759,N_6148,N_6766);
or U7760 (N_7760,N_6223,N_6973);
xnor U7761 (N_7761,N_6134,N_6126);
nor U7762 (N_7762,N_6523,N_6443);
nand U7763 (N_7763,N_6707,N_6407);
and U7764 (N_7764,N_6060,N_6903);
nor U7765 (N_7765,N_6550,N_6142);
or U7766 (N_7766,N_6471,N_6899);
xnor U7767 (N_7767,N_6163,N_6359);
nor U7768 (N_7768,N_6389,N_6941);
or U7769 (N_7769,N_6613,N_6816);
xnor U7770 (N_7770,N_6275,N_6858);
xnor U7771 (N_7771,N_6072,N_6444);
nand U7772 (N_7772,N_6094,N_6185);
nor U7773 (N_7773,N_6913,N_6743);
or U7774 (N_7774,N_6948,N_6488);
nor U7775 (N_7775,N_6501,N_6677);
nand U7776 (N_7776,N_6632,N_6191);
or U7777 (N_7777,N_6044,N_6004);
xnor U7778 (N_7778,N_6364,N_6659);
nand U7779 (N_7779,N_6565,N_6576);
nand U7780 (N_7780,N_6725,N_6756);
and U7781 (N_7781,N_6727,N_6572);
and U7782 (N_7782,N_6106,N_6111);
nor U7783 (N_7783,N_6226,N_6508);
and U7784 (N_7784,N_6939,N_6980);
and U7785 (N_7785,N_6620,N_6991);
xnor U7786 (N_7786,N_6333,N_6129);
or U7787 (N_7787,N_6575,N_6474);
xor U7788 (N_7788,N_6586,N_6072);
nand U7789 (N_7789,N_6267,N_6386);
or U7790 (N_7790,N_6794,N_6129);
or U7791 (N_7791,N_6685,N_6733);
nor U7792 (N_7792,N_6618,N_6085);
or U7793 (N_7793,N_6626,N_6925);
or U7794 (N_7794,N_6048,N_6188);
and U7795 (N_7795,N_6137,N_6954);
nor U7796 (N_7796,N_6687,N_6928);
and U7797 (N_7797,N_6107,N_6915);
or U7798 (N_7798,N_6862,N_6520);
and U7799 (N_7799,N_6113,N_6412);
and U7800 (N_7800,N_6867,N_6935);
nor U7801 (N_7801,N_6502,N_6581);
nand U7802 (N_7802,N_6850,N_6205);
nor U7803 (N_7803,N_6519,N_6235);
nor U7804 (N_7804,N_6273,N_6729);
xor U7805 (N_7805,N_6817,N_6568);
nand U7806 (N_7806,N_6346,N_6797);
xnor U7807 (N_7807,N_6176,N_6011);
and U7808 (N_7808,N_6663,N_6136);
and U7809 (N_7809,N_6279,N_6646);
nor U7810 (N_7810,N_6803,N_6534);
nand U7811 (N_7811,N_6379,N_6306);
and U7812 (N_7812,N_6128,N_6026);
and U7813 (N_7813,N_6528,N_6091);
and U7814 (N_7814,N_6340,N_6440);
and U7815 (N_7815,N_6229,N_6373);
nor U7816 (N_7816,N_6980,N_6204);
and U7817 (N_7817,N_6075,N_6691);
xnor U7818 (N_7818,N_6024,N_6622);
or U7819 (N_7819,N_6735,N_6757);
and U7820 (N_7820,N_6143,N_6744);
xnor U7821 (N_7821,N_6299,N_6409);
xnor U7822 (N_7822,N_6498,N_6571);
and U7823 (N_7823,N_6487,N_6081);
xor U7824 (N_7824,N_6670,N_6477);
and U7825 (N_7825,N_6445,N_6129);
and U7826 (N_7826,N_6668,N_6064);
xor U7827 (N_7827,N_6511,N_6138);
nor U7828 (N_7828,N_6774,N_6120);
xor U7829 (N_7829,N_6276,N_6333);
xnor U7830 (N_7830,N_6145,N_6231);
nand U7831 (N_7831,N_6123,N_6962);
xnor U7832 (N_7832,N_6034,N_6955);
or U7833 (N_7833,N_6628,N_6305);
nor U7834 (N_7834,N_6784,N_6219);
xor U7835 (N_7835,N_6964,N_6067);
nor U7836 (N_7836,N_6655,N_6036);
nand U7837 (N_7837,N_6300,N_6765);
and U7838 (N_7838,N_6083,N_6959);
nor U7839 (N_7839,N_6791,N_6521);
or U7840 (N_7840,N_6285,N_6953);
or U7841 (N_7841,N_6147,N_6757);
nand U7842 (N_7842,N_6891,N_6830);
nor U7843 (N_7843,N_6682,N_6922);
xnor U7844 (N_7844,N_6574,N_6281);
nand U7845 (N_7845,N_6149,N_6373);
and U7846 (N_7846,N_6782,N_6904);
and U7847 (N_7847,N_6955,N_6109);
nand U7848 (N_7848,N_6866,N_6345);
and U7849 (N_7849,N_6954,N_6908);
and U7850 (N_7850,N_6338,N_6819);
and U7851 (N_7851,N_6824,N_6049);
or U7852 (N_7852,N_6030,N_6470);
xnor U7853 (N_7853,N_6236,N_6821);
xor U7854 (N_7854,N_6548,N_6896);
xor U7855 (N_7855,N_6531,N_6444);
xnor U7856 (N_7856,N_6896,N_6533);
nor U7857 (N_7857,N_6907,N_6993);
and U7858 (N_7858,N_6921,N_6757);
xor U7859 (N_7859,N_6634,N_6952);
nand U7860 (N_7860,N_6985,N_6595);
nor U7861 (N_7861,N_6378,N_6993);
and U7862 (N_7862,N_6003,N_6613);
nor U7863 (N_7863,N_6434,N_6284);
or U7864 (N_7864,N_6771,N_6733);
and U7865 (N_7865,N_6058,N_6184);
and U7866 (N_7866,N_6655,N_6911);
xor U7867 (N_7867,N_6689,N_6612);
and U7868 (N_7868,N_6522,N_6117);
and U7869 (N_7869,N_6615,N_6548);
and U7870 (N_7870,N_6821,N_6572);
or U7871 (N_7871,N_6272,N_6602);
and U7872 (N_7872,N_6559,N_6771);
xnor U7873 (N_7873,N_6893,N_6767);
and U7874 (N_7874,N_6268,N_6446);
and U7875 (N_7875,N_6003,N_6264);
xnor U7876 (N_7876,N_6380,N_6181);
xnor U7877 (N_7877,N_6827,N_6898);
xnor U7878 (N_7878,N_6852,N_6057);
or U7879 (N_7879,N_6896,N_6753);
nand U7880 (N_7880,N_6626,N_6953);
xnor U7881 (N_7881,N_6791,N_6650);
xnor U7882 (N_7882,N_6767,N_6488);
or U7883 (N_7883,N_6620,N_6503);
nand U7884 (N_7884,N_6879,N_6153);
nor U7885 (N_7885,N_6100,N_6590);
nand U7886 (N_7886,N_6843,N_6094);
nand U7887 (N_7887,N_6691,N_6756);
xnor U7888 (N_7888,N_6758,N_6905);
xor U7889 (N_7889,N_6272,N_6051);
nand U7890 (N_7890,N_6933,N_6693);
or U7891 (N_7891,N_6863,N_6712);
nor U7892 (N_7892,N_6884,N_6741);
xnor U7893 (N_7893,N_6074,N_6989);
or U7894 (N_7894,N_6248,N_6734);
nor U7895 (N_7895,N_6257,N_6824);
nand U7896 (N_7896,N_6628,N_6867);
and U7897 (N_7897,N_6301,N_6801);
or U7898 (N_7898,N_6645,N_6911);
xor U7899 (N_7899,N_6371,N_6213);
nand U7900 (N_7900,N_6662,N_6834);
xnor U7901 (N_7901,N_6009,N_6188);
or U7902 (N_7902,N_6550,N_6618);
nor U7903 (N_7903,N_6761,N_6723);
and U7904 (N_7904,N_6047,N_6054);
nor U7905 (N_7905,N_6208,N_6501);
or U7906 (N_7906,N_6758,N_6591);
nor U7907 (N_7907,N_6729,N_6786);
and U7908 (N_7908,N_6070,N_6853);
or U7909 (N_7909,N_6514,N_6146);
and U7910 (N_7910,N_6412,N_6102);
and U7911 (N_7911,N_6994,N_6907);
xnor U7912 (N_7912,N_6373,N_6883);
nor U7913 (N_7913,N_6060,N_6489);
nand U7914 (N_7914,N_6706,N_6124);
nand U7915 (N_7915,N_6890,N_6754);
xnor U7916 (N_7916,N_6550,N_6891);
xor U7917 (N_7917,N_6739,N_6226);
xor U7918 (N_7918,N_6673,N_6531);
xor U7919 (N_7919,N_6705,N_6447);
nor U7920 (N_7920,N_6458,N_6366);
nand U7921 (N_7921,N_6485,N_6766);
nand U7922 (N_7922,N_6664,N_6498);
nand U7923 (N_7923,N_6610,N_6074);
and U7924 (N_7924,N_6594,N_6850);
and U7925 (N_7925,N_6840,N_6693);
nor U7926 (N_7926,N_6588,N_6583);
nand U7927 (N_7927,N_6428,N_6923);
or U7928 (N_7928,N_6252,N_6972);
nor U7929 (N_7929,N_6095,N_6433);
nor U7930 (N_7930,N_6539,N_6801);
nor U7931 (N_7931,N_6611,N_6353);
and U7932 (N_7932,N_6819,N_6975);
nor U7933 (N_7933,N_6068,N_6337);
nor U7934 (N_7934,N_6104,N_6295);
nand U7935 (N_7935,N_6686,N_6867);
nand U7936 (N_7936,N_6403,N_6128);
and U7937 (N_7937,N_6581,N_6195);
nand U7938 (N_7938,N_6010,N_6880);
or U7939 (N_7939,N_6378,N_6120);
or U7940 (N_7940,N_6736,N_6441);
or U7941 (N_7941,N_6175,N_6279);
nor U7942 (N_7942,N_6636,N_6651);
nor U7943 (N_7943,N_6507,N_6549);
or U7944 (N_7944,N_6021,N_6439);
nand U7945 (N_7945,N_6107,N_6011);
nand U7946 (N_7946,N_6057,N_6060);
and U7947 (N_7947,N_6618,N_6375);
nand U7948 (N_7948,N_6292,N_6747);
nor U7949 (N_7949,N_6214,N_6942);
nor U7950 (N_7950,N_6789,N_6748);
xor U7951 (N_7951,N_6036,N_6299);
and U7952 (N_7952,N_6190,N_6034);
and U7953 (N_7953,N_6633,N_6941);
and U7954 (N_7954,N_6036,N_6747);
nand U7955 (N_7955,N_6416,N_6971);
and U7956 (N_7956,N_6507,N_6500);
nand U7957 (N_7957,N_6879,N_6644);
xnor U7958 (N_7958,N_6962,N_6182);
xor U7959 (N_7959,N_6244,N_6277);
or U7960 (N_7960,N_6794,N_6810);
nand U7961 (N_7961,N_6295,N_6272);
and U7962 (N_7962,N_6013,N_6857);
nand U7963 (N_7963,N_6432,N_6100);
xor U7964 (N_7964,N_6773,N_6278);
nor U7965 (N_7965,N_6468,N_6382);
nand U7966 (N_7966,N_6734,N_6964);
nor U7967 (N_7967,N_6354,N_6585);
and U7968 (N_7968,N_6908,N_6823);
nor U7969 (N_7969,N_6472,N_6352);
nand U7970 (N_7970,N_6468,N_6391);
nand U7971 (N_7971,N_6938,N_6366);
and U7972 (N_7972,N_6998,N_6967);
xor U7973 (N_7973,N_6864,N_6725);
xor U7974 (N_7974,N_6752,N_6602);
nor U7975 (N_7975,N_6326,N_6460);
nor U7976 (N_7976,N_6845,N_6329);
xor U7977 (N_7977,N_6723,N_6700);
xor U7978 (N_7978,N_6434,N_6314);
xnor U7979 (N_7979,N_6549,N_6447);
nor U7980 (N_7980,N_6956,N_6202);
and U7981 (N_7981,N_6332,N_6368);
nor U7982 (N_7982,N_6157,N_6725);
nor U7983 (N_7983,N_6429,N_6436);
nor U7984 (N_7984,N_6315,N_6782);
and U7985 (N_7985,N_6765,N_6054);
or U7986 (N_7986,N_6622,N_6436);
xor U7987 (N_7987,N_6460,N_6818);
and U7988 (N_7988,N_6252,N_6219);
and U7989 (N_7989,N_6013,N_6902);
xor U7990 (N_7990,N_6001,N_6523);
and U7991 (N_7991,N_6118,N_6386);
or U7992 (N_7992,N_6356,N_6027);
nand U7993 (N_7993,N_6753,N_6157);
or U7994 (N_7994,N_6927,N_6774);
nor U7995 (N_7995,N_6552,N_6454);
and U7996 (N_7996,N_6761,N_6360);
xnor U7997 (N_7997,N_6488,N_6574);
xor U7998 (N_7998,N_6265,N_6569);
nor U7999 (N_7999,N_6777,N_6182);
xnor U8000 (N_8000,N_7953,N_7951);
nand U8001 (N_8001,N_7217,N_7976);
and U8002 (N_8002,N_7949,N_7159);
xnor U8003 (N_8003,N_7535,N_7143);
nor U8004 (N_8004,N_7222,N_7815);
nor U8005 (N_8005,N_7154,N_7673);
and U8006 (N_8006,N_7403,N_7347);
and U8007 (N_8007,N_7350,N_7515);
or U8008 (N_8008,N_7959,N_7634);
nor U8009 (N_8009,N_7050,N_7832);
xor U8010 (N_8010,N_7916,N_7896);
nand U8011 (N_8011,N_7726,N_7731);
nor U8012 (N_8012,N_7840,N_7266);
or U8013 (N_8013,N_7869,N_7259);
xor U8014 (N_8014,N_7683,N_7556);
nor U8015 (N_8015,N_7824,N_7493);
xnor U8016 (N_8016,N_7190,N_7590);
nor U8017 (N_8017,N_7453,N_7199);
or U8018 (N_8018,N_7390,N_7473);
nand U8019 (N_8019,N_7382,N_7823);
and U8020 (N_8020,N_7408,N_7298);
nand U8021 (N_8021,N_7311,N_7447);
nor U8022 (N_8022,N_7293,N_7448);
nand U8023 (N_8023,N_7530,N_7970);
or U8024 (N_8024,N_7985,N_7723);
or U8025 (N_8025,N_7569,N_7081);
xnor U8026 (N_8026,N_7601,N_7341);
xor U8027 (N_8027,N_7269,N_7006);
nand U8028 (N_8028,N_7317,N_7602);
xnor U8029 (N_8029,N_7559,N_7302);
nand U8030 (N_8030,N_7044,N_7391);
or U8031 (N_8031,N_7172,N_7284);
or U8032 (N_8032,N_7520,N_7964);
or U8033 (N_8033,N_7123,N_7054);
or U8034 (N_8034,N_7801,N_7682);
nor U8035 (N_8035,N_7924,N_7454);
or U8036 (N_8036,N_7499,N_7254);
and U8037 (N_8037,N_7129,N_7336);
nor U8038 (N_8038,N_7645,N_7605);
xnor U8039 (N_8039,N_7374,N_7288);
nand U8040 (N_8040,N_7607,N_7544);
and U8041 (N_8041,N_7240,N_7704);
nor U8042 (N_8042,N_7622,N_7082);
nor U8043 (N_8043,N_7641,N_7722);
and U8044 (N_8044,N_7435,N_7466);
and U8045 (N_8045,N_7911,N_7920);
nand U8046 (N_8046,N_7234,N_7517);
xnor U8047 (N_8047,N_7277,N_7105);
or U8048 (N_8048,N_7210,N_7656);
nor U8049 (N_8049,N_7021,N_7078);
nor U8050 (N_8050,N_7136,N_7904);
xor U8051 (N_8051,N_7402,N_7810);
nand U8052 (N_8052,N_7863,N_7065);
nand U8053 (N_8053,N_7371,N_7780);
and U8054 (N_8054,N_7087,N_7836);
nand U8055 (N_8055,N_7119,N_7411);
or U8056 (N_8056,N_7040,N_7670);
or U8057 (N_8057,N_7680,N_7899);
or U8058 (N_8058,N_7508,N_7902);
xor U8059 (N_8059,N_7507,N_7060);
nor U8060 (N_8060,N_7183,N_7464);
nor U8061 (N_8061,N_7686,N_7460);
xor U8062 (N_8062,N_7197,N_7853);
or U8063 (N_8063,N_7735,N_7662);
nor U8064 (N_8064,N_7271,N_7474);
or U8065 (N_8065,N_7330,N_7106);
nand U8066 (N_8066,N_7525,N_7000);
or U8067 (N_8067,N_7676,N_7173);
xnor U8068 (N_8068,N_7618,N_7191);
nand U8069 (N_8069,N_7063,N_7459);
xnor U8070 (N_8070,N_7431,N_7773);
xor U8071 (N_8071,N_7113,N_7725);
and U8072 (N_8072,N_7692,N_7931);
or U8073 (N_8073,N_7762,N_7884);
xor U8074 (N_8074,N_7619,N_7788);
nor U8075 (N_8075,N_7872,N_7224);
xnor U8076 (N_8076,N_7068,N_7938);
xor U8077 (N_8077,N_7555,N_7351);
nand U8078 (N_8078,N_7481,N_7945);
xor U8079 (N_8079,N_7839,N_7895);
nor U8080 (N_8080,N_7609,N_7230);
nand U8081 (N_8081,N_7069,N_7398);
nand U8082 (N_8082,N_7175,N_7978);
or U8083 (N_8083,N_7015,N_7480);
nand U8084 (N_8084,N_7881,N_7080);
nand U8085 (N_8085,N_7498,N_7642);
and U8086 (N_8086,N_7548,N_7135);
nor U8087 (N_8087,N_7316,N_7873);
nor U8088 (N_8088,N_7756,N_7308);
and U8089 (N_8089,N_7410,N_7306);
nand U8090 (N_8090,N_7344,N_7373);
or U8091 (N_8091,N_7192,N_7061);
or U8092 (N_8092,N_7227,N_7261);
and U8093 (N_8093,N_7637,N_7636);
and U8094 (N_8094,N_7130,N_7971);
nand U8095 (N_8095,N_7941,N_7358);
and U8096 (N_8096,N_7760,N_7467);
nand U8097 (N_8097,N_7355,N_7303);
or U8098 (N_8098,N_7007,N_7857);
or U8099 (N_8099,N_7084,N_7991);
or U8100 (N_8100,N_7223,N_7456);
or U8101 (N_8101,N_7663,N_7797);
nand U8102 (N_8102,N_7189,N_7606);
or U8103 (N_8103,N_7998,N_7596);
xor U8104 (N_8104,N_7378,N_7621);
nand U8105 (N_8105,N_7386,N_7772);
or U8106 (N_8106,N_7237,N_7580);
and U8107 (N_8107,N_7141,N_7458);
nor U8108 (N_8108,N_7935,N_7108);
and U8109 (N_8109,N_7558,N_7203);
xnor U8110 (N_8110,N_7965,N_7418);
and U8111 (N_8111,N_7029,N_7258);
nand U8112 (N_8112,N_7013,N_7434);
and U8113 (N_8113,N_7030,N_7887);
or U8114 (N_8114,N_7455,N_7765);
xnor U8115 (N_8115,N_7443,N_7811);
and U8116 (N_8116,N_7724,N_7281);
or U8117 (N_8117,N_7919,N_7890);
xor U8118 (N_8118,N_7048,N_7100);
nand U8119 (N_8119,N_7501,N_7714);
nand U8120 (N_8120,N_7235,N_7687);
and U8121 (N_8121,N_7956,N_7574);
or U8122 (N_8122,N_7085,N_7362);
nor U8123 (N_8123,N_7343,N_7334);
nand U8124 (N_8124,N_7784,N_7462);
or U8125 (N_8125,N_7326,N_7977);
nand U8126 (N_8126,N_7888,N_7101);
xor U8127 (N_8127,N_7201,N_7388);
nand U8128 (N_8128,N_7655,N_7587);
nor U8129 (N_8129,N_7339,N_7929);
nor U8130 (N_8130,N_7167,N_7875);
nor U8131 (N_8131,N_7174,N_7097);
or U8132 (N_8132,N_7116,N_7504);
xnor U8133 (N_8133,N_7290,N_7543);
nor U8134 (N_8134,N_7653,N_7878);
xnor U8135 (N_8135,N_7648,N_7755);
and U8136 (N_8136,N_7109,N_7425);
nor U8137 (N_8137,N_7250,N_7743);
and U8138 (N_8138,N_7521,N_7565);
nor U8139 (N_8139,N_7208,N_7107);
nand U8140 (N_8140,N_7990,N_7727);
xor U8141 (N_8141,N_7251,N_7786);
nor U8142 (N_8142,N_7318,N_7879);
and U8143 (N_8143,N_7830,N_7128);
or U8144 (N_8144,N_7630,N_7769);
or U8145 (N_8145,N_7289,N_7059);
nand U8146 (N_8146,N_7996,N_7551);
and U8147 (N_8147,N_7286,N_7180);
and U8148 (N_8148,N_7171,N_7575);
nand U8149 (N_8149,N_7323,N_7522);
and U8150 (N_8150,N_7685,N_7534);
and U8151 (N_8151,N_7793,N_7588);
nand U8152 (N_8152,N_7110,N_7342);
or U8153 (N_8153,N_7913,N_7294);
and U8154 (N_8154,N_7471,N_7276);
xor U8155 (N_8155,N_7209,N_7690);
and U8156 (N_8156,N_7452,N_7248);
or U8157 (N_8157,N_7672,N_7491);
xor U8158 (N_8158,N_7668,N_7694);
xnor U8159 (N_8159,N_7376,N_7427);
or U8160 (N_8160,N_7489,N_7002);
nor U8161 (N_8161,N_7239,N_7972);
nand U8162 (N_8162,N_7885,N_7018);
and U8163 (N_8163,N_7337,N_7028);
nand U8164 (N_8164,N_7958,N_7360);
nand U8165 (N_8165,N_7581,N_7406);
xnor U8166 (N_8166,N_7541,N_7791);
and U8167 (N_8167,N_7843,N_7436);
nand U8168 (N_8168,N_7592,N_7862);
or U8169 (N_8169,N_7554,N_7893);
nand U8170 (N_8170,N_7450,N_7093);
xnor U8171 (N_8171,N_7001,N_7829);
and U8172 (N_8172,N_7688,N_7265);
nand U8173 (N_8173,N_7967,N_7741);
nand U8174 (N_8174,N_7616,N_7738);
xor U8175 (N_8175,N_7632,N_7485);
nand U8176 (N_8176,N_7218,N_7202);
and U8177 (N_8177,N_7708,N_7272);
xnor U8178 (N_8178,N_7055,N_7463);
xnor U8179 (N_8179,N_7075,N_7274);
and U8180 (N_8180,N_7858,N_7927);
xnor U8181 (N_8181,N_7661,N_7961);
or U8182 (N_8182,N_7500,N_7940);
xnor U8183 (N_8183,N_7200,N_7761);
and U8184 (N_8184,N_7903,N_7695);
xnor U8185 (N_8185,N_7312,N_7273);
and U8186 (N_8186,N_7763,N_7946);
or U8187 (N_8187,N_7948,N_7345);
or U8188 (N_8188,N_7138,N_7803);
and U8189 (N_8189,N_7379,N_7943);
nand U8190 (N_8190,N_7363,N_7338);
and U8191 (N_8191,N_7368,N_7086);
and U8192 (N_8192,N_7072,N_7417);
nand U8193 (N_8193,N_7721,N_7986);
xor U8194 (N_8194,N_7912,N_7891);
or U8195 (N_8195,N_7533,N_7992);
or U8196 (N_8196,N_7357,N_7660);
nand U8197 (N_8197,N_7512,N_7297);
nand U8198 (N_8198,N_7092,N_7827);
or U8199 (N_8199,N_7322,N_7187);
and U8200 (N_8200,N_7229,N_7428);
nand U8201 (N_8201,N_7936,N_7492);
and U8202 (N_8202,N_7283,N_7650);
nor U8203 (N_8203,N_7538,N_7974);
nand U8204 (N_8204,N_7540,N_7262);
nand U8205 (N_8205,N_7939,N_7833);
nor U8206 (N_8206,N_7795,N_7659);
nor U8207 (N_8207,N_7077,N_7693);
and U8208 (N_8208,N_7781,N_7400);
or U8209 (N_8209,N_7487,N_7184);
nor U8210 (N_8210,N_7654,N_7325);
or U8211 (N_8211,N_7383,N_7825);
or U8212 (N_8212,N_7518,N_7744);
nand U8213 (N_8213,N_7354,N_7812);
xor U8214 (N_8214,N_7871,N_7212);
nand U8215 (N_8215,N_7560,N_7665);
and U8216 (N_8216,N_7153,N_7268);
xor U8217 (N_8217,N_7291,N_7635);
nand U8218 (N_8218,N_7300,N_7805);
nor U8219 (N_8219,N_7145,N_7897);
nand U8220 (N_8220,N_7926,N_7319);
nand U8221 (N_8221,N_7578,N_7349);
nor U8222 (N_8222,N_7134,N_7031);
xnor U8223 (N_8223,N_7429,N_7516);
xnor U8224 (N_8224,N_7754,N_7664);
and U8225 (N_8225,N_7442,N_7667);
xnor U8226 (N_8226,N_7421,N_7757);
and U8227 (N_8227,N_7639,N_7828);
and U8228 (N_8228,N_7915,N_7917);
nor U8229 (N_8229,N_7073,N_7838);
or U8230 (N_8230,N_7594,N_7238);
or U8231 (N_8231,N_7674,N_7122);
or U8232 (N_8232,N_7571,N_7163);
and U8233 (N_8233,N_7851,N_7717);
xor U8234 (N_8234,N_7745,N_7742);
nand U8235 (N_8235,N_7177,N_7035);
nand U8236 (N_8236,N_7707,N_7027);
or U8237 (N_8237,N_7999,N_7599);
and U8238 (N_8238,N_7033,N_7156);
or U8239 (N_8239,N_7292,N_7090);
nand U8240 (N_8240,N_7937,N_7583);
xnor U8241 (N_8241,N_7994,N_7011);
and U8242 (N_8242,N_7132,N_7979);
or U8243 (N_8243,N_7880,N_7993);
nand U8244 (N_8244,N_7207,N_7257);
and U8245 (N_8245,N_7758,N_7285);
xnor U8246 (N_8246,N_7249,N_7367);
and U8247 (N_8247,N_7528,N_7196);
or U8248 (N_8248,N_7779,N_7389);
nor U8249 (N_8249,N_7346,N_7506);
nor U8250 (N_8250,N_7553,N_7557);
and U8251 (N_8251,N_7279,N_7987);
and U8252 (N_8252,N_7385,N_7807);
nor U8253 (N_8253,N_7729,N_7603);
nor U8254 (N_8254,N_7989,N_7861);
nor U8255 (N_8255,N_7882,N_7296);
xnor U8256 (N_8256,N_7465,N_7394);
and U8257 (N_8257,N_7352,N_7681);
nand U8258 (N_8258,N_7867,N_7988);
or U8259 (N_8259,N_7395,N_7572);
xnor U8260 (N_8260,N_7894,N_7980);
and U8261 (N_8261,N_7914,N_7503);
nor U8262 (N_8262,N_7247,N_7009);
and U8263 (N_8263,N_7562,N_7211);
or U8264 (N_8264,N_7524,N_7014);
and U8265 (N_8265,N_7168,N_7537);
nor U8266 (N_8266,N_7675,N_7550);
and U8267 (N_8267,N_7901,N_7445);
nand U8268 (N_8268,N_7124,N_7438);
nor U8269 (N_8269,N_7188,N_7270);
nand U8270 (N_8270,N_7933,N_7928);
nor U8271 (N_8271,N_7563,N_7749);
nand U8272 (N_8272,N_7866,N_7133);
or U8273 (N_8273,N_7115,N_7652);
nand U8274 (N_8274,N_7963,N_7221);
or U8275 (N_8275,N_7709,N_7094);
nand U8276 (N_8276,N_7424,N_7127);
nor U8277 (N_8277,N_7620,N_7178);
and U8278 (N_8278,N_7321,N_7865);
nand U8279 (N_8279,N_7969,N_7204);
xnor U8280 (N_8280,N_7399,N_7246);
or U8281 (N_8281,N_7706,N_7483);
or U8282 (N_8282,N_7377,N_7275);
or U8283 (N_8283,N_7091,N_7739);
nand U8284 (N_8284,N_7472,N_7906);
or U8285 (N_8285,N_7611,N_7102);
and U8286 (N_8286,N_7042,N_7020);
nor U8287 (N_8287,N_7767,N_7245);
nor U8288 (N_8288,N_7396,N_7814);
nor U8289 (N_8289,N_7004,N_7730);
nand U8290 (N_8290,N_7118,N_7039);
xor U8291 (N_8291,N_7886,N_7701);
xnor U8292 (N_8292,N_7817,N_7822);
and U8293 (N_8293,N_7638,N_7629);
xnor U8294 (N_8294,N_7697,N_7612);
or U8295 (N_8295,N_7740,N_7095);
xor U8296 (N_8296,N_7647,N_7658);
nor U8297 (N_8297,N_7225,N_7752);
and U8298 (N_8298,N_7407,N_7328);
and U8299 (N_8299,N_7478,N_7733);
or U8300 (N_8300,N_7753,N_7151);
and U8301 (N_8301,N_7778,N_7950);
xnor U8302 (N_8302,N_7324,N_7846);
nor U8303 (N_8303,N_7327,N_7148);
nand U8304 (N_8304,N_7719,N_7103);
and U8305 (N_8305,N_7140,N_7045);
nand U8306 (N_8306,N_7718,N_7484);
nand U8307 (N_8307,N_7278,N_7526);
and U8308 (N_8308,N_7008,N_7984);
nor U8309 (N_8309,N_7305,N_7513);
nor U8310 (N_8310,N_7155,N_7161);
or U8311 (N_8311,N_7633,N_7019);
or U8312 (N_8312,N_7214,N_7195);
or U8313 (N_8313,N_7691,N_7461);
xor U8314 (N_8314,N_7205,N_7868);
and U8315 (N_8315,N_7139,N_7051);
nor U8316 (N_8316,N_7058,N_7255);
or U8317 (N_8317,N_7372,N_7955);
and U8318 (N_8318,N_7164,N_7333);
and U8319 (N_8319,N_7071,N_7837);
nand U8320 (N_8320,N_7981,N_7313);
nand U8321 (N_8321,N_7856,N_7005);
nor U8322 (N_8322,N_7568,N_7567);
and U8323 (N_8323,N_7287,N_7185);
nand U8324 (N_8324,N_7111,N_7074);
nor U8325 (N_8325,N_7671,N_7220);
and U8326 (N_8326,N_7315,N_7790);
xor U8327 (N_8327,N_7446,N_7831);
xnor U8328 (N_8328,N_7819,N_7842);
nand U8329 (N_8329,N_7966,N_7420);
nor U8330 (N_8330,N_7366,N_7468);
nand U8331 (N_8331,N_7598,N_7393);
nand U8332 (N_8332,N_7549,N_7295);
nand U8333 (N_8333,N_7835,N_7152);
or U8334 (N_8334,N_7610,N_7510);
xor U8335 (N_8335,N_7043,N_7231);
xnor U8336 (N_8336,N_7527,N_7877);
or U8337 (N_8337,N_7046,N_7962);
or U8338 (N_8338,N_7944,N_7826);
and U8339 (N_8339,N_7617,N_7536);
nor U8340 (N_8340,N_7908,N_7041);
nand U8341 (N_8341,N_7475,N_7047);
and U8342 (N_8342,N_7012,N_7870);
or U8343 (N_8343,N_7038,N_7802);
nand U8344 (N_8344,N_7808,N_7206);
nand U8345 (N_8345,N_7158,N_7960);
nor U8346 (N_8346,N_7451,N_7748);
and U8347 (N_8347,N_7126,N_7573);
nand U8348 (N_8348,N_7799,N_7056);
and U8349 (N_8349,N_7734,N_7649);
and U8350 (N_8350,N_7643,N_7626);
or U8351 (N_8351,N_7282,N_7120);
nor U8352 (N_8352,N_7490,N_7957);
nand U8353 (N_8353,N_7502,N_7244);
xnor U8354 (N_8354,N_7181,N_7432);
xor U8355 (N_8355,N_7523,N_7702);
and U8356 (N_8356,N_7820,N_7444);
nor U8357 (N_8357,N_7062,N_7713);
or U8358 (N_8358,N_7413,N_7604);
and U8359 (N_8359,N_7854,N_7098);
nor U8360 (N_8360,N_7792,N_7785);
nand U8361 (N_8361,N_7215,N_7096);
or U8362 (N_8362,N_7025,N_7646);
and U8363 (N_8363,N_7975,N_7783);
or U8364 (N_8364,N_7678,N_7874);
nand U8365 (N_8365,N_7728,N_7364);
nand U8366 (N_8366,N_7750,N_7712);
nand U8367 (N_8367,N_7479,N_7776);
xor U8368 (N_8368,N_7737,N_7179);
nor U8369 (N_8369,N_7625,N_7859);
nand U8370 (N_8370,N_7699,N_7770);
and U8371 (N_8371,N_7022,N_7566);
nor U8372 (N_8372,N_7705,N_7099);
nand U8373 (N_8373,N_7932,N_7934);
nand U8374 (N_8374,N_7213,N_7157);
xnor U8375 (N_8375,N_7796,N_7684);
nand U8376 (N_8376,N_7804,N_7582);
and U8377 (N_8377,N_7023,N_7160);
nand U8378 (N_8378,N_7076,N_7593);
and U8379 (N_8379,N_7083,N_7798);
and U8380 (N_8380,N_7243,N_7057);
nand U8381 (N_8381,N_7923,N_7586);
xor U8382 (N_8382,N_7651,N_7380);
nor U8383 (N_8383,N_7834,N_7310);
xor U8384 (N_8384,N_7314,N_7905);
or U8385 (N_8385,N_7552,N_7585);
nand U8386 (N_8386,N_7532,N_7644);
and U8387 (N_8387,N_7117,N_7064);
nand U8388 (N_8388,N_7608,N_7666);
or U8389 (N_8389,N_7369,N_7497);
or U8390 (N_8390,N_7470,N_7782);
xor U8391 (N_8391,N_7412,N_7301);
and U8392 (N_8392,N_7623,N_7561);
and U8393 (N_8393,N_7010,N_7361);
and U8394 (N_8394,N_7716,N_7079);
or U8395 (N_8395,N_7488,N_7182);
nor U8396 (N_8396,N_7876,N_7165);
or U8397 (N_8397,N_7631,N_7356);
nand U8398 (N_8398,N_7017,N_7348);
or U8399 (N_8399,N_7775,N_7968);
xnor U8400 (N_8400,N_7026,N_7925);
nand U8401 (N_8401,N_7365,N_7253);
and U8402 (N_8402,N_7024,N_7067);
xnor U8403 (N_8403,N_7787,N_7392);
and U8404 (N_8404,N_7496,N_7628);
nand U8405 (N_8405,N_7053,N_7600);
nand U8406 (N_8406,N_7844,N_7732);
nor U8407 (N_8407,N_7242,N_7613);
nor U8408 (N_8408,N_7511,N_7304);
or U8409 (N_8409,N_7711,N_7267);
xnor U8410 (N_8410,N_7766,N_7669);
nand U8411 (N_8411,N_7845,N_7627);
nor U8412 (N_8412,N_7370,N_7439);
nand U8413 (N_8413,N_7307,N_7494);
or U8414 (N_8414,N_7700,N_7794);
xnor U8415 (N_8415,N_7457,N_7864);
nand U8416 (N_8416,N_7260,N_7768);
nand U8417 (N_8417,N_7907,N_7774);
nand U8418 (N_8418,N_7764,N_7909);
nand U8419 (N_8419,N_7147,N_7264);
and U8420 (N_8420,N_7529,N_7003);
nor U8421 (N_8421,N_7892,N_7353);
nand U8422 (N_8422,N_7137,N_7759);
nor U8423 (N_8423,N_7034,N_7469);
nand U8424 (N_8424,N_7016,N_7850);
and U8425 (N_8425,N_7146,N_7104);
and U8426 (N_8426,N_7900,N_7545);
nor U8427 (N_8427,N_7514,N_7495);
xor U8428 (N_8428,N_7689,N_7409);
or U8429 (N_8429,N_7777,N_7589);
or U8430 (N_8430,N_7049,N_7806);
xor U8431 (N_8431,N_7415,N_7449);
nor U8432 (N_8432,N_7821,N_7430);
xor U8433 (N_8433,N_7952,N_7800);
and U8434 (N_8434,N_7849,N_7226);
and U8435 (N_8435,N_7889,N_7070);
nor U8436 (N_8436,N_7150,N_7997);
xor U8437 (N_8437,N_7036,N_7162);
or U8438 (N_8438,N_7579,N_7232);
nand U8439 (N_8439,N_7614,N_7309);
nand U8440 (N_8440,N_7883,N_7112);
xor U8441 (N_8441,N_7404,N_7125);
or U8442 (N_8442,N_7983,N_7089);
xnor U8443 (N_8443,N_7921,N_7263);
nand U8444 (N_8444,N_7252,N_7696);
or U8445 (N_8445,N_7698,N_7898);
and U8446 (N_8446,N_7414,N_7852);
nor U8447 (N_8447,N_7624,N_7847);
nor U8448 (N_8448,N_7280,N_7228);
xnor U8449 (N_8449,N_7597,N_7359);
nand U8450 (N_8450,N_7615,N_7816);
and U8451 (N_8451,N_7677,N_7416);
nor U8452 (N_8452,N_7922,N_7751);
or U8453 (N_8453,N_7746,N_7547);
nor U8454 (N_8454,N_7332,N_7703);
nor U8455 (N_8455,N_7423,N_7789);
xor U8456 (N_8456,N_7576,N_7144);
and U8457 (N_8457,N_7942,N_7771);
nor U8458 (N_8458,N_7595,N_7397);
nor U8459 (N_8459,N_7570,N_7419);
nand U8460 (N_8460,N_7375,N_7584);
nand U8461 (N_8461,N_7947,N_7331);
or U8462 (N_8462,N_7422,N_7329);
and U8463 (N_8463,N_7486,N_7169);
and U8464 (N_8464,N_7170,N_7405);
and U8465 (N_8465,N_7509,N_7973);
nor U8466 (N_8466,N_7131,N_7720);
xnor U8467 (N_8467,N_7381,N_7505);
xor U8468 (N_8468,N_7747,N_7982);
nand U8469 (N_8469,N_7860,N_7149);
and U8470 (N_8470,N_7114,N_7679);
nand U8471 (N_8471,N_7052,N_7066);
or U8472 (N_8472,N_7193,N_7256);
nor U8473 (N_8473,N_7531,N_7387);
nor U8474 (N_8474,N_7166,N_7216);
nor U8475 (N_8475,N_7476,N_7037);
and U8476 (N_8476,N_7441,N_7320);
nand U8477 (N_8477,N_7426,N_7433);
or U8478 (N_8478,N_7910,N_7142);
and U8479 (N_8479,N_7198,N_7219);
and U8480 (N_8480,N_7546,N_7437);
or U8481 (N_8481,N_7657,N_7335);
xnor U8482 (N_8482,N_7539,N_7564);
nor U8483 (N_8483,N_7194,N_7176);
nand U8484 (N_8484,N_7809,N_7241);
or U8485 (N_8485,N_7233,N_7482);
xnor U8486 (N_8486,N_7930,N_7918);
nand U8487 (N_8487,N_7186,N_7340);
or U8488 (N_8488,N_7591,N_7818);
xor U8489 (N_8489,N_7848,N_7121);
nand U8490 (N_8490,N_7813,N_7577);
nand U8491 (N_8491,N_7032,N_7384);
xnor U8492 (N_8492,N_7841,N_7995);
xnor U8493 (N_8493,N_7299,N_7477);
or U8494 (N_8494,N_7640,N_7736);
nand U8495 (N_8495,N_7440,N_7542);
nor U8496 (N_8496,N_7710,N_7401);
nor U8497 (N_8497,N_7954,N_7715);
xnor U8498 (N_8498,N_7519,N_7236);
and U8499 (N_8499,N_7088,N_7855);
nand U8500 (N_8500,N_7049,N_7230);
nor U8501 (N_8501,N_7968,N_7064);
or U8502 (N_8502,N_7177,N_7280);
xor U8503 (N_8503,N_7800,N_7837);
nor U8504 (N_8504,N_7915,N_7649);
xnor U8505 (N_8505,N_7312,N_7796);
nor U8506 (N_8506,N_7095,N_7986);
nor U8507 (N_8507,N_7103,N_7415);
or U8508 (N_8508,N_7971,N_7284);
nor U8509 (N_8509,N_7084,N_7593);
nor U8510 (N_8510,N_7210,N_7594);
and U8511 (N_8511,N_7971,N_7370);
nand U8512 (N_8512,N_7559,N_7878);
nand U8513 (N_8513,N_7288,N_7986);
nor U8514 (N_8514,N_7229,N_7114);
and U8515 (N_8515,N_7857,N_7009);
xor U8516 (N_8516,N_7763,N_7422);
and U8517 (N_8517,N_7750,N_7934);
or U8518 (N_8518,N_7423,N_7080);
nand U8519 (N_8519,N_7916,N_7643);
or U8520 (N_8520,N_7538,N_7516);
and U8521 (N_8521,N_7910,N_7713);
nor U8522 (N_8522,N_7203,N_7730);
nor U8523 (N_8523,N_7631,N_7323);
nand U8524 (N_8524,N_7068,N_7973);
nor U8525 (N_8525,N_7589,N_7191);
nand U8526 (N_8526,N_7882,N_7416);
or U8527 (N_8527,N_7504,N_7264);
nor U8528 (N_8528,N_7087,N_7190);
nand U8529 (N_8529,N_7874,N_7565);
xor U8530 (N_8530,N_7399,N_7807);
xnor U8531 (N_8531,N_7540,N_7146);
nand U8532 (N_8532,N_7812,N_7613);
nor U8533 (N_8533,N_7467,N_7097);
nand U8534 (N_8534,N_7050,N_7211);
nor U8535 (N_8535,N_7799,N_7037);
and U8536 (N_8536,N_7087,N_7789);
or U8537 (N_8537,N_7963,N_7140);
and U8538 (N_8538,N_7092,N_7101);
nand U8539 (N_8539,N_7303,N_7927);
or U8540 (N_8540,N_7057,N_7138);
nand U8541 (N_8541,N_7674,N_7153);
nand U8542 (N_8542,N_7053,N_7481);
nand U8543 (N_8543,N_7921,N_7619);
or U8544 (N_8544,N_7254,N_7554);
or U8545 (N_8545,N_7055,N_7948);
nor U8546 (N_8546,N_7652,N_7582);
or U8547 (N_8547,N_7397,N_7157);
nand U8548 (N_8548,N_7069,N_7361);
or U8549 (N_8549,N_7976,N_7587);
xnor U8550 (N_8550,N_7618,N_7930);
nor U8551 (N_8551,N_7129,N_7523);
and U8552 (N_8552,N_7040,N_7693);
and U8553 (N_8553,N_7784,N_7573);
nand U8554 (N_8554,N_7314,N_7422);
nand U8555 (N_8555,N_7856,N_7832);
or U8556 (N_8556,N_7703,N_7152);
nand U8557 (N_8557,N_7685,N_7962);
and U8558 (N_8558,N_7564,N_7025);
nand U8559 (N_8559,N_7653,N_7813);
or U8560 (N_8560,N_7323,N_7508);
and U8561 (N_8561,N_7965,N_7492);
nand U8562 (N_8562,N_7759,N_7366);
and U8563 (N_8563,N_7900,N_7802);
xnor U8564 (N_8564,N_7689,N_7608);
xnor U8565 (N_8565,N_7449,N_7482);
nand U8566 (N_8566,N_7935,N_7565);
xnor U8567 (N_8567,N_7313,N_7756);
or U8568 (N_8568,N_7217,N_7372);
and U8569 (N_8569,N_7863,N_7703);
nor U8570 (N_8570,N_7034,N_7761);
nand U8571 (N_8571,N_7980,N_7420);
xor U8572 (N_8572,N_7943,N_7976);
xor U8573 (N_8573,N_7526,N_7086);
and U8574 (N_8574,N_7826,N_7112);
xnor U8575 (N_8575,N_7417,N_7975);
or U8576 (N_8576,N_7257,N_7178);
nor U8577 (N_8577,N_7768,N_7569);
or U8578 (N_8578,N_7286,N_7129);
nor U8579 (N_8579,N_7045,N_7457);
xor U8580 (N_8580,N_7958,N_7590);
nor U8581 (N_8581,N_7440,N_7205);
or U8582 (N_8582,N_7727,N_7942);
and U8583 (N_8583,N_7631,N_7071);
and U8584 (N_8584,N_7755,N_7789);
and U8585 (N_8585,N_7218,N_7152);
or U8586 (N_8586,N_7234,N_7159);
nand U8587 (N_8587,N_7925,N_7280);
nand U8588 (N_8588,N_7021,N_7268);
nand U8589 (N_8589,N_7503,N_7928);
or U8590 (N_8590,N_7725,N_7541);
xor U8591 (N_8591,N_7520,N_7629);
nor U8592 (N_8592,N_7102,N_7723);
or U8593 (N_8593,N_7991,N_7245);
or U8594 (N_8594,N_7701,N_7052);
or U8595 (N_8595,N_7887,N_7311);
nor U8596 (N_8596,N_7359,N_7619);
nand U8597 (N_8597,N_7531,N_7182);
and U8598 (N_8598,N_7563,N_7983);
and U8599 (N_8599,N_7741,N_7921);
xnor U8600 (N_8600,N_7936,N_7344);
nand U8601 (N_8601,N_7743,N_7906);
or U8602 (N_8602,N_7444,N_7603);
or U8603 (N_8603,N_7761,N_7705);
nand U8604 (N_8604,N_7281,N_7323);
and U8605 (N_8605,N_7101,N_7655);
nand U8606 (N_8606,N_7315,N_7984);
nor U8607 (N_8607,N_7352,N_7123);
or U8608 (N_8608,N_7524,N_7720);
or U8609 (N_8609,N_7568,N_7770);
xnor U8610 (N_8610,N_7060,N_7544);
or U8611 (N_8611,N_7348,N_7446);
and U8612 (N_8612,N_7010,N_7533);
nand U8613 (N_8613,N_7138,N_7463);
xnor U8614 (N_8614,N_7510,N_7390);
nor U8615 (N_8615,N_7155,N_7656);
nand U8616 (N_8616,N_7048,N_7273);
or U8617 (N_8617,N_7130,N_7650);
nor U8618 (N_8618,N_7990,N_7289);
or U8619 (N_8619,N_7533,N_7756);
or U8620 (N_8620,N_7719,N_7137);
or U8621 (N_8621,N_7216,N_7562);
xor U8622 (N_8622,N_7377,N_7139);
and U8623 (N_8623,N_7892,N_7975);
and U8624 (N_8624,N_7176,N_7786);
nor U8625 (N_8625,N_7803,N_7817);
nand U8626 (N_8626,N_7207,N_7975);
nand U8627 (N_8627,N_7999,N_7880);
or U8628 (N_8628,N_7510,N_7647);
or U8629 (N_8629,N_7876,N_7347);
and U8630 (N_8630,N_7011,N_7292);
xor U8631 (N_8631,N_7320,N_7045);
and U8632 (N_8632,N_7690,N_7858);
and U8633 (N_8633,N_7005,N_7680);
nand U8634 (N_8634,N_7789,N_7184);
xnor U8635 (N_8635,N_7875,N_7199);
xor U8636 (N_8636,N_7300,N_7818);
and U8637 (N_8637,N_7049,N_7218);
nor U8638 (N_8638,N_7455,N_7314);
xnor U8639 (N_8639,N_7969,N_7889);
or U8640 (N_8640,N_7967,N_7597);
nand U8641 (N_8641,N_7121,N_7029);
nor U8642 (N_8642,N_7755,N_7965);
xnor U8643 (N_8643,N_7900,N_7555);
and U8644 (N_8644,N_7345,N_7723);
or U8645 (N_8645,N_7397,N_7893);
nand U8646 (N_8646,N_7676,N_7040);
nor U8647 (N_8647,N_7650,N_7890);
xor U8648 (N_8648,N_7027,N_7313);
xor U8649 (N_8649,N_7489,N_7418);
nor U8650 (N_8650,N_7965,N_7071);
nor U8651 (N_8651,N_7063,N_7197);
nand U8652 (N_8652,N_7527,N_7760);
nor U8653 (N_8653,N_7722,N_7623);
nor U8654 (N_8654,N_7573,N_7214);
nand U8655 (N_8655,N_7610,N_7058);
nand U8656 (N_8656,N_7391,N_7899);
and U8657 (N_8657,N_7808,N_7415);
xor U8658 (N_8658,N_7183,N_7069);
or U8659 (N_8659,N_7355,N_7025);
and U8660 (N_8660,N_7765,N_7346);
and U8661 (N_8661,N_7095,N_7021);
nor U8662 (N_8662,N_7536,N_7301);
and U8663 (N_8663,N_7423,N_7069);
xor U8664 (N_8664,N_7508,N_7321);
and U8665 (N_8665,N_7580,N_7200);
and U8666 (N_8666,N_7174,N_7975);
xnor U8667 (N_8667,N_7398,N_7604);
xnor U8668 (N_8668,N_7015,N_7978);
xor U8669 (N_8669,N_7875,N_7485);
nor U8670 (N_8670,N_7571,N_7765);
or U8671 (N_8671,N_7067,N_7496);
xor U8672 (N_8672,N_7491,N_7961);
xor U8673 (N_8673,N_7206,N_7191);
or U8674 (N_8674,N_7038,N_7153);
nand U8675 (N_8675,N_7690,N_7974);
nor U8676 (N_8676,N_7643,N_7871);
nor U8677 (N_8677,N_7362,N_7712);
and U8678 (N_8678,N_7393,N_7585);
xor U8679 (N_8679,N_7037,N_7106);
or U8680 (N_8680,N_7433,N_7025);
and U8681 (N_8681,N_7835,N_7034);
or U8682 (N_8682,N_7683,N_7389);
and U8683 (N_8683,N_7807,N_7182);
xor U8684 (N_8684,N_7779,N_7618);
or U8685 (N_8685,N_7922,N_7149);
nand U8686 (N_8686,N_7734,N_7984);
xor U8687 (N_8687,N_7967,N_7529);
xor U8688 (N_8688,N_7993,N_7953);
xnor U8689 (N_8689,N_7529,N_7322);
nand U8690 (N_8690,N_7803,N_7224);
xor U8691 (N_8691,N_7733,N_7923);
nand U8692 (N_8692,N_7550,N_7077);
nand U8693 (N_8693,N_7571,N_7403);
and U8694 (N_8694,N_7425,N_7852);
or U8695 (N_8695,N_7722,N_7784);
and U8696 (N_8696,N_7601,N_7377);
or U8697 (N_8697,N_7964,N_7297);
or U8698 (N_8698,N_7476,N_7295);
and U8699 (N_8699,N_7756,N_7585);
nor U8700 (N_8700,N_7836,N_7496);
or U8701 (N_8701,N_7953,N_7212);
or U8702 (N_8702,N_7737,N_7891);
xor U8703 (N_8703,N_7713,N_7197);
xnor U8704 (N_8704,N_7223,N_7917);
xor U8705 (N_8705,N_7828,N_7265);
nand U8706 (N_8706,N_7619,N_7878);
nor U8707 (N_8707,N_7142,N_7754);
and U8708 (N_8708,N_7085,N_7882);
nor U8709 (N_8709,N_7142,N_7678);
and U8710 (N_8710,N_7864,N_7462);
and U8711 (N_8711,N_7299,N_7584);
xnor U8712 (N_8712,N_7843,N_7282);
or U8713 (N_8713,N_7694,N_7473);
nand U8714 (N_8714,N_7191,N_7488);
xnor U8715 (N_8715,N_7690,N_7412);
or U8716 (N_8716,N_7134,N_7999);
or U8717 (N_8717,N_7134,N_7970);
nand U8718 (N_8718,N_7769,N_7857);
nor U8719 (N_8719,N_7093,N_7517);
or U8720 (N_8720,N_7291,N_7632);
nand U8721 (N_8721,N_7508,N_7693);
xor U8722 (N_8722,N_7977,N_7604);
or U8723 (N_8723,N_7579,N_7117);
or U8724 (N_8724,N_7231,N_7358);
or U8725 (N_8725,N_7325,N_7042);
xor U8726 (N_8726,N_7542,N_7218);
nand U8727 (N_8727,N_7823,N_7989);
or U8728 (N_8728,N_7379,N_7763);
and U8729 (N_8729,N_7836,N_7963);
nor U8730 (N_8730,N_7302,N_7637);
nor U8731 (N_8731,N_7248,N_7076);
or U8732 (N_8732,N_7458,N_7933);
nand U8733 (N_8733,N_7961,N_7580);
nand U8734 (N_8734,N_7516,N_7137);
nor U8735 (N_8735,N_7224,N_7696);
or U8736 (N_8736,N_7321,N_7837);
nor U8737 (N_8737,N_7392,N_7377);
nor U8738 (N_8738,N_7653,N_7299);
nand U8739 (N_8739,N_7220,N_7067);
nand U8740 (N_8740,N_7354,N_7155);
and U8741 (N_8741,N_7871,N_7973);
nand U8742 (N_8742,N_7074,N_7673);
xnor U8743 (N_8743,N_7602,N_7269);
or U8744 (N_8744,N_7355,N_7502);
or U8745 (N_8745,N_7332,N_7633);
nand U8746 (N_8746,N_7679,N_7318);
nand U8747 (N_8747,N_7396,N_7002);
nor U8748 (N_8748,N_7499,N_7900);
nor U8749 (N_8749,N_7694,N_7729);
nor U8750 (N_8750,N_7564,N_7081);
or U8751 (N_8751,N_7199,N_7404);
nand U8752 (N_8752,N_7201,N_7477);
or U8753 (N_8753,N_7456,N_7230);
or U8754 (N_8754,N_7356,N_7096);
nand U8755 (N_8755,N_7054,N_7666);
nor U8756 (N_8756,N_7316,N_7453);
xor U8757 (N_8757,N_7785,N_7360);
nand U8758 (N_8758,N_7112,N_7843);
nor U8759 (N_8759,N_7084,N_7930);
and U8760 (N_8760,N_7592,N_7239);
and U8761 (N_8761,N_7795,N_7175);
or U8762 (N_8762,N_7399,N_7489);
and U8763 (N_8763,N_7578,N_7553);
and U8764 (N_8764,N_7819,N_7878);
nand U8765 (N_8765,N_7920,N_7261);
nor U8766 (N_8766,N_7229,N_7884);
xor U8767 (N_8767,N_7962,N_7285);
xnor U8768 (N_8768,N_7610,N_7957);
nand U8769 (N_8769,N_7650,N_7946);
nor U8770 (N_8770,N_7335,N_7582);
nand U8771 (N_8771,N_7590,N_7435);
and U8772 (N_8772,N_7901,N_7886);
nand U8773 (N_8773,N_7890,N_7366);
xor U8774 (N_8774,N_7101,N_7854);
nand U8775 (N_8775,N_7196,N_7108);
nand U8776 (N_8776,N_7626,N_7935);
and U8777 (N_8777,N_7587,N_7750);
and U8778 (N_8778,N_7061,N_7951);
and U8779 (N_8779,N_7039,N_7605);
nor U8780 (N_8780,N_7449,N_7681);
xor U8781 (N_8781,N_7773,N_7264);
xnor U8782 (N_8782,N_7111,N_7906);
and U8783 (N_8783,N_7198,N_7744);
and U8784 (N_8784,N_7811,N_7960);
nor U8785 (N_8785,N_7035,N_7903);
xor U8786 (N_8786,N_7179,N_7344);
nand U8787 (N_8787,N_7928,N_7188);
nor U8788 (N_8788,N_7182,N_7760);
nor U8789 (N_8789,N_7075,N_7824);
nand U8790 (N_8790,N_7589,N_7507);
or U8791 (N_8791,N_7522,N_7495);
nand U8792 (N_8792,N_7007,N_7095);
xor U8793 (N_8793,N_7689,N_7432);
and U8794 (N_8794,N_7294,N_7959);
and U8795 (N_8795,N_7579,N_7888);
and U8796 (N_8796,N_7909,N_7512);
nor U8797 (N_8797,N_7185,N_7752);
nor U8798 (N_8798,N_7148,N_7780);
nand U8799 (N_8799,N_7202,N_7461);
or U8800 (N_8800,N_7813,N_7486);
and U8801 (N_8801,N_7272,N_7468);
nor U8802 (N_8802,N_7656,N_7592);
nor U8803 (N_8803,N_7513,N_7244);
xnor U8804 (N_8804,N_7859,N_7448);
xnor U8805 (N_8805,N_7214,N_7927);
or U8806 (N_8806,N_7293,N_7575);
or U8807 (N_8807,N_7308,N_7959);
xor U8808 (N_8808,N_7730,N_7627);
nand U8809 (N_8809,N_7781,N_7733);
nand U8810 (N_8810,N_7867,N_7921);
nor U8811 (N_8811,N_7811,N_7484);
nor U8812 (N_8812,N_7517,N_7668);
xor U8813 (N_8813,N_7030,N_7878);
nor U8814 (N_8814,N_7860,N_7725);
and U8815 (N_8815,N_7267,N_7992);
and U8816 (N_8816,N_7411,N_7223);
xor U8817 (N_8817,N_7525,N_7925);
nand U8818 (N_8818,N_7894,N_7621);
xnor U8819 (N_8819,N_7995,N_7143);
and U8820 (N_8820,N_7774,N_7030);
xor U8821 (N_8821,N_7688,N_7139);
or U8822 (N_8822,N_7032,N_7797);
nand U8823 (N_8823,N_7134,N_7787);
and U8824 (N_8824,N_7456,N_7824);
nor U8825 (N_8825,N_7976,N_7228);
nand U8826 (N_8826,N_7037,N_7806);
nor U8827 (N_8827,N_7824,N_7737);
xnor U8828 (N_8828,N_7362,N_7650);
nand U8829 (N_8829,N_7012,N_7577);
nand U8830 (N_8830,N_7934,N_7482);
nand U8831 (N_8831,N_7481,N_7141);
nor U8832 (N_8832,N_7260,N_7546);
or U8833 (N_8833,N_7136,N_7306);
nor U8834 (N_8834,N_7932,N_7097);
xnor U8835 (N_8835,N_7932,N_7349);
or U8836 (N_8836,N_7706,N_7726);
nand U8837 (N_8837,N_7613,N_7443);
xnor U8838 (N_8838,N_7108,N_7686);
nor U8839 (N_8839,N_7090,N_7696);
and U8840 (N_8840,N_7163,N_7733);
nand U8841 (N_8841,N_7431,N_7031);
nand U8842 (N_8842,N_7607,N_7519);
xor U8843 (N_8843,N_7191,N_7926);
nor U8844 (N_8844,N_7049,N_7020);
and U8845 (N_8845,N_7551,N_7637);
xor U8846 (N_8846,N_7191,N_7946);
and U8847 (N_8847,N_7361,N_7771);
or U8848 (N_8848,N_7874,N_7522);
nand U8849 (N_8849,N_7075,N_7381);
and U8850 (N_8850,N_7911,N_7472);
and U8851 (N_8851,N_7652,N_7507);
nor U8852 (N_8852,N_7281,N_7123);
xnor U8853 (N_8853,N_7916,N_7790);
nor U8854 (N_8854,N_7790,N_7873);
or U8855 (N_8855,N_7120,N_7564);
or U8856 (N_8856,N_7675,N_7420);
nor U8857 (N_8857,N_7168,N_7295);
xnor U8858 (N_8858,N_7404,N_7970);
or U8859 (N_8859,N_7601,N_7487);
and U8860 (N_8860,N_7607,N_7987);
nand U8861 (N_8861,N_7499,N_7971);
and U8862 (N_8862,N_7701,N_7759);
and U8863 (N_8863,N_7485,N_7187);
or U8864 (N_8864,N_7768,N_7513);
nor U8865 (N_8865,N_7660,N_7929);
xnor U8866 (N_8866,N_7589,N_7804);
xnor U8867 (N_8867,N_7030,N_7643);
or U8868 (N_8868,N_7468,N_7686);
or U8869 (N_8869,N_7227,N_7471);
or U8870 (N_8870,N_7027,N_7556);
nand U8871 (N_8871,N_7179,N_7416);
xor U8872 (N_8872,N_7940,N_7571);
and U8873 (N_8873,N_7538,N_7872);
nand U8874 (N_8874,N_7676,N_7971);
nand U8875 (N_8875,N_7982,N_7513);
and U8876 (N_8876,N_7775,N_7836);
nor U8877 (N_8877,N_7124,N_7878);
and U8878 (N_8878,N_7668,N_7852);
xnor U8879 (N_8879,N_7509,N_7868);
and U8880 (N_8880,N_7026,N_7892);
and U8881 (N_8881,N_7527,N_7618);
or U8882 (N_8882,N_7839,N_7723);
nand U8883 (N_8883,N_7801,N_7226);
and U8884 (N_8884,N_7472,N_7049);
nand U8885 (N_8885,N_7349,N_7235);
nor U8886 (N_8886,N_7649,N_7474);
or U8887 (N_8887,N_7228,N_7147);
or U8888 (N_8888,N_7658,N_7365);
xnor U8889 (N_8889,N_7516,N_7958);
and U8890 (N_8890,N_7228,N_7622);
or U8891 (N_8891,N_7852,N_7779);
nor U8892 (N_8892,N_7290,N_7811);
xnor U8893 (N_8893,N_7806,N_7760);
xor U8894 (N_8894,N_7830,N_7564);
nor U8895 (N_8895,N_7013,N_7509);
nand U8896 (N_8896,N_7567,N_7903);
nand U8897 (N_8897,N_7410,N_7099);
nor U8898 (N_8898,N_7732,N_7428);
nor U8899 (N_8899,N_7847,N_7206);
nand U8900 (N_8900,N_7019,N_7796);
and U8901 (N_8901,N_7579,N_7671);
xnor U8902 (N_8902,N_7772,N_7192);
or U8903 (N_8903,N_7801,N_7586);
and U8904 (N_8904,N_7493,N_7884);
and U8905 (N_8905,N_7867,N_7520);
nor U8906 (N_8906,N_7503,N_7324);
nor U8907 (N_8907,N_7937,N_7507);
nor U8908 (N_8908,N_7947,N_7084);
or U8909 (N_8909,N_7189,N_7147);
nor U8910 (N_8910,N_7948,N_7808);
nor U8911 (N_8911,N_7102,N_7188);
xnor U8912 (N_8912,N_7641,N_7850);
nor U8913 (N_8913,N_7982,N_7298);
nor U8914 (N_8914,N_7568,N_7463);
nor U8915 (N_8915,N_7533,N_7474);
nand U8916 (N_8916,N_7914,N_7314);
nor U8917 (N_8917,N_7551,N_7173);
nand U8918 (N_8918,N_7120,N_7808);
and U8919 (N_8919,N_7799,N_7588);
and U8920 (N_8920,N_7385,N_7364);
or U8921 (N_8921,N_7506,N_7320);
and U8922 (N_8922,N_7823,N_7172);
or U8923 (N_8923,N_7713,N_7107);
or U8924 (N_8924,N_7429,N_7040);
xnor U8925 (N_8925,N_7592,N_7791);
or U8926 (N_8926,N_7848,N_7980);
or U8927 (N_8927,N_7624,N_7962);
nor U8928 (N_8928,N_7459,N_7222);
or U8929 (N_8929,N_7541,N_7918);
and U8930 (N_8930,N_7390,N_7535);
and U8931 (N_8931,N_7553,N_7083);
and U8932 (N_8932,N_7736,N_7554);
nand U8933 (N_8933,N_7139,N_7424);
and U8934 (N_8934,N_7737,N_7856);
nand U8935 (N_8935,N_7571,N_7900);
nor U8936 (N_8936,N_7109,N_7964);
nand U8937 (N_8937,N_7350,N_7015);
nor U8938 (N_8938,N_7028,N_7293);
nand U8939 (N_8939,N_7733,N_7654);
xnor U8940 (N_8940,N_7569,N_7950);
xor U8941 (N_8941,N_7209,N_7926);
nand U8942 (N_8942,N_7797,N_7322);
and U8943 (N_8943,N_7326,N_7989);
or U8944 (N_8944,N_7508,N_7088);
and U8945 (N_8945,N_7277,N_7167);
xor U8946 (N_8946,N_7750,N_7087);
or U8947 (N_8947,N_7371,N_7099);
and U8948 (N_8948,N_7937,N_7252);
nand U8949 (N_8949,N_7737,N_7017);
xnor U8950 (N_8950,N_7720,N_7912);
and U8951 (N_8951,N_7222,N_7483);
nor U8952 (N_8952,N_7203,N_7277);
nor U8953 (N_8953,N_7694,N_7259);
or U8954 (N_8954,N_7956,N_7552);
nor U8955 (N_8955,N_7751,N_7649);
nand U8956 (N_8956,N_7593,N_7095);
nand U8957 (N_8957,N_7185,N_7569);
nor U8958 (N_8958,N_7457,N_7057);
xnor U8959 (N_8959,N_7556,N_7704);
nor U8960 (N_8960,N_7195,N_7761);
and U8961 (N_8961,N_7819,N_7448);
or U8962 (N_8962,N_7590,N_7777);
and U8963 (N_8963,N_7870,N_7389);
or U8964 (N_8964,N_7657,N_7144);
or U8965 (N_8965,N_7339,N_7902);
nor U8966 (N_8966,N_7590,N_7279);
and U8967 (N_8967,N_7952,N_7301);
and U8968 (N_8968,N_7835,N_7326);
or U8969 (N_8969,N_7085,N_7068);
and U8970 (N_8970,N_7193,N_7025);
or U8971 (N_8971,N_7787,N_7772);
and U8972 (N_8972,N_7854,N_7882);
nand U8973 (N_8973,N_7618,N_7033);
xnor U8974 (N_8974,N_7001,N_7789);
or U8975 (N_8975,N_7844,N_7184);
xnor U8976 (N_8976,N_7489,N_7144);
and U8977 (N_8977,N_7491,N_7040);
or U8978 (N_8978,N_7957,N_7915);
xor U8979 (N_8979,N_7734,N_7509);
nor U8980 (N_8980,N_7607,N_7793);
nand U8981 (N_8981,N_7729,N_7171);
xor U8982 (N_8982,N_7076,N_7217);
and U8983 (N_8983,N_7126,N_7606);
and U8984 (N_8984,N_7973,N_7168);
and U8985 (N_8985,N_7786,N_7741);
or U8986 (N_8986,N_7107,N_7728);
or U8987 (N_8987,N_7527,N_7848);
and U8988 (N_8988,N_7271,N_7161);
and U8989 (N_8989,N_7907,N_7187);
or U8990 (N_8990,N_7995,N_7197);
nand U8991 (N_8991,N_7528,N_7539);
nor U8992 (N_8992,N_7795,N_7437);
nand U8993 (N_8993,N_7218,N_7036);
and U8994 (N_8994,N_7713,N_7112);
and U8995 (N_8995,N_7036,N_7815);
nand U8996 (N_8996,N_7162,N_7945);
and U8997 (N_8997,N_7443,N_7501);
nand U8998 (N_8998,N_7061,N_7054);
xor U8999 (N_8999,N_7453,N_7822);
nand U9000 (N_9000,N_8920,N_8158);
nor U9001 (N_9001,N_8754,N_8237);
and U9002 (N_9002,N_8236,N_8492);
nand U9003 (N_9003,N_8428,N_8577);
and U9004 (N_9004,N_8047,N_8285);
xnor U9005 (N_9005,N_8957,N_8634);
nand U9006 (N_9006,N_8548,N_8891);
or U9007 (N_9007,N_8629,N_8355);
and U9008 (N_9008,N_8288,N_8838);
and U9009 (N_9009,N_8547,N_8823);
and U9010 (N_9010,N_8145,N_8804);
or U9011 (N_9011,N_8259,N_8636);
xnor U9012 (N_9012,N_8928,N_8533);
xnor U9013 (N_9013,N_8349,N_8739);
and U9014 (N_9014,N_8734,N_8850);
nand U9015 (N_9015,N_8263,N_8280);
nor U9016 (N_9016,N_8654,N_8282);
or U9017 (N_9017,N_8019,N_8029);
nor U9018 (N_9018,N_8855,N_8726);
and U9019 (N_9019,N_8300,N_8925);
xor U9020 (N_9020,N_8779,N_8065);
xnor U9021 (N_9021,N_8796,N_8187);
or U9022 (N_9022,N_8767,N_8657);
and U9023 (N_9023,N_8458,N_8879);
and U9024 (N_9024,N_8315,N_8388);
and U9025 (N_9025,N_8277,N_8619);
or U9026 (N_9026,N_8747,N_8030);
or U9027 (N_9027,N_8111,N_8421);
and U9028 (N_9028,N_8916,N_8055);
xor U9029 (N_9029,N_8875,N_8929);
xor U9030 (N_9030,N_8893,N_8057);
and U9031 (N_9031,N_8614,N_8602);
xor U9032 (N_9032,N_8364,N_8094);
xor U9033 (N_9033,N_8782,N_8971);
nor U9034 (N_9034,N_8402,N_8665);
or U9035 (N_9035,N_8487,N_8085);
and U9036 (N_9036,N_8616,N_8507);
and U9037 (N_9037,N_8161,N_8563);
and U9038 (N_9038,N_8670,N_8105);
and U9039 (N_9039,N_8358,N_8289);
xnor U9040 (N_9040,N_8382,N_8174);
and U9041 (N_9041,N_8213,N_8522);
nor U9042 (N_9042,N_8933,N_8902);
xnor U9043 (N_9043,N_8895,N_8535);
and U9044 (N_9044,N_8760,N_8110);
xor U9045 (N_9045,N_8699,N_8196);
xnor U9046 (N_9046,N_8653,N_8203);
xor U9047 (N_9047,N_8440,N_8718);
and U9048 (N_9048,N_8419,N_8673);
nor U9049 (N_9049,N_8150,N_8633);
nand U9050 (N_9050,N_8183,N_8341);
xnor U9051 (N_9051,N_8171,N_8239);
and U9052 (N_9052,N_8301,N_8869);
nand U9053 (N_9053,N_8207,N_8177);
and U9054 (N_9054,N_8095,N_8870);
or U9055 (N_9055,N_8595,N_8041);
nor U9056 (N_9056,N_8587,N_8296);
and U9057 (N_9057,N_8609,N_8214);
and U9058 (N_9058,N_8143,N_8409);
nand U9059 (N_9059,N_8276,N_8938);
or U9060 (N_9060,N_8186,N_8346);
nor U9061 (N_9061,N_8042,N_8475);
and U9062 (N_9062,N_8156,N_8062);
or U9063 (N_9063,N_8255,N_8700);
xnor U9064 (N_9064,N_8827,N_8520);
nor U9065 (N_9065,N_8218,N_8676);
or U9066 (N_9066,N_8993,N_8119);
xor U9067 (N_9067,N_8627,N_8082);
and U9068 (N_9068,N_8710,N_8674);
or U9069 (N_9069,N_8903,N_8572);
nor U9070 (N_9070,N_8864,N_8652);
nor U9071 (N_9071,N_8248,N_8446);
nor U9072 (N_9072,N_8148,N_8694);
xor U9073 (N_9073,N_8774,N_8284);
xnor U9074 (N_9074,N_8374,N_8025);
nand U9075 (N_9075,N_8818,N_8687);
or U9076 (N_9076,N_8287,N_8232);
xor U9077 (N_9077,N_8939,N_8594);
and U9078 (N_9078,N_8045,N_8155);
or U9079 (N_9079,N_8641,N_8299);
nor U9080 (N_9080,N_8112,N_8354);
or U9081 (N_9081,N_8684,N_8337);
nor U9082 (N_9082,N_8224,N_8473);
nor U9083 (N_9083,N_8467,N_8021);
nand U9084 (N_9084,N_8540,N_8560);
and U9085 (N_9085,N_8116,N_8182);
or U9086 (N_9086,N_8778,N_8840);
nand U9087 (N_9087,N_8940,N_8262);
or U9088 (N_9088,N_8539,N_8833);
or U9089 (N_9089,N_8621,N_8012);
or U9090 (N_9090,N_8815,N_8886);
and U9091 (N_9091,N_8672,N_8521);
nor U9092 (N_9092,N_8705,N_8848);
nand U9093 (N_9093,N_8080,N_8486);
or U9094 (N_9094,N_8841,N_8471);
nand U9095 (N_9095,N_8666,N_8427);
nor U9096 (N_9096,N_8347,N_8046);
and U9097 (N_9097,N_8789,N_8575);
or U9098 (N_9098,N_8089,N_8311);
nand U9099 (N_9099,N_8704,N_8215);
nand U9100 (N_9100,N_8510,N_8418);
xor U9101 (N_9101,N_8439,N_8530);
and U9102 (N_9102,N_8728,N_8561);
or U9103 (N_9103,N_8137,N_8892);
or U9104 (N_9104,N_8541,N_8585);
xnor U9105 (N_9105,N_8274,N_8820);
or U9106 (N_9106,N_8909,N_8733);
nand U9107 (N_9107,N_8783,N_8332);
xor U9108 (N_9108,N_8872,N_8251);
nor U9109 (N_9109,N_8067,N_8984);
nor U9110 (N_9110,N_8593,N_8292);
xor U9111 (N_9111,N_8442,N_8570);
or U9112 (N_9112,N_8389,N_8400);
and U9113 (N_9113,N_8922,N_8958);
nand U9114 (N_9114,N_8556,N_8759);
or U9115 (N_9115,N_8640,N_8352);
or U9116 (N_9116,N_8240,N_8596);
or U9117 (N_9117,N_8859,N_8873);
nand U9118 (N_9118,N_8983,N_8888);
nand U9119 (N_9119,N_8342,N_8153);
nand U9120 (N_9120,N_8317,N_8201);
nand U9121 (N_9121,N_8954,N_8429);
or U9122 (N_9122,N_8788,N_8549);
and U9123 (N_9123,N_8081,N_8076);
or U9124 (N_9124,N_8669,N_8499);
or U9125 (N_9125,N_8582,N_8321);
and U9126 (N_9126,N_8776,N_8298);
nor U9127 (N_9127,N_8612,N_8613);
xnor U9128 (N_9128,N_8949,N_8795);
nand U9129 (N_9129,N_8688,N_8787);
xnor U9130 (N_9130,N_8597,N_8506);
xor U9131 (N_9131,N_8573,N_8966);
or U9132 (N_9132,N_8412,N_8786);
nand U9133 (N_9133,N_8511,N_8777);
nand U9134 (N_9134,N_8134,N_8310);
and U9135 (N_9135,N_8508,N_8509);
or U9136 (N_9136,N_8987,N_8588);
and U9137 (N_9137,N_8675,N_8191);
nor U9138 (N_9138,N_8106,N_8632);
or U9139 (N_9139,N_8905,N_8569);
or U9140 (N_9140,N_8927,N_8297);
nand U9141 (N_9141,N_8264,N_8845);
xnor U9142 (N_9142,N_8740,N_8142);
and U9143 (N_9143,N_8279,N_8562);
and U9144 (N_9144,N_8498,N_8557);
nor U9145 (N_9145,N_8189,N_8396);
nor U9146 (N_9146,N_8491,N_8554);
nand U9147 (N_9147,N_8960,N_8951);
xnor U9148 (N_9148,N_8680,N_8483);
or U9149 (N_9149,N_8398,N_8260);
and U9150 (N_9150,N_8455,N_8496);
xnor U9151 (N_9151,N_8559,N_8885);
and U9152 (N_9152,N_8843,N_8581);
nand U9153 (N_9153,N_8743,N_8384);
nor U9154 (N_9154,N_8459,N_8635);
nand U9155 (N_9155,N_8008,N_8646);
xor U9156 (N_9156,N_8985,N_8791);
and U9157 (N_9157,N_8469,N_8825);
nor U9158 (N_9158,N_8121,N_8417);
nand U9159 (N_9159,N_8371,N_8188);
and U9160 (N_9160,N_8628,N_8713);
or U9161 (N_9161,N_8480,N_8265);
nor U9162 (N_9162,N_8645,N_8500);
nand U9163 (N_9163,N_8617,N_8069);
nand U9164 (N_9164,N_8146,N_8436);
nand U9165 (N_9165,N_8749,N_8387);
nand U9166 (N_9166,N_8399,N_8824);
xnor U9167 (N_9167,N_8915,N_8338);
nand U9168 (N_9168,N_8431,N_8200);
nand U9169 (N_9169,N_8519,N_8307);
nand U9170 (N_9170,N_8424,N_8878);
nor U9171 (N_9171,N_8720,N_8172);
xnor U9172 (N_9172,N_8644,N_8147);
or U9173 (N_9173,N_8322,N_8009);
or U9174 (N_9174,N_8553,N_8844);
and U9175 (N_9175,N_8972,N_8751);
and U9176 (N_9176,N_8752,N_8862);
xnor U9177 (N_9177,N_8977,N_8166);
nor U9178 (N_9178,N_8851,N_8717);
and U9179 (N_9179,N_8835,N_8910);
nor U9180 (N_9180,N_8136,N_8798);
or U9181 (N_9181,N_8981,N_8536);
and U9182 (N_9182,N_8441,N_8222);
or U9183 (N_9183,N_8999,N_8742);
nor U9184 (N_9184,N_8501,N_8370);
or U9185 (N_9185,N_8220,N_8772);
nand U9186 (N_9186,N_8775,N_8626);
xor U9187 (N_9187,N_8810,N_8714);
nand U9188 (N_9188,N_8378,N_8638);
or U9189 (N_9189,N_8980,N_8883);
nor U9190 (N_9190,N_8765,N_8231);
xor U9191 (N_9191,N_8329,N_8416);
or U9192 (N_9192,N_8286,N_8668);
xnor U9193 (N_9193,N_8730,N_8324);
nor U9194 (N_9194,N_8525,N_8357);
xnor U9195 (N_9195,N_8408,N_8488);
or U9196 (N_9196,N_8472,N_8502);
or U9197 (N_9197,N_8071,N_8725);
and U9198 (N_9198,N_8495,N_8805);
nand U9199 (N_9199,N_8120,N_8591);
or U9200 (N_9200,N_8123,N_8233);
xnor U9201 (N_9201,N_8662,N_8132);
and U9202 (N_9202,N_8216,N_8624);
nand U9203 (N_9203,N_8195,N_8550);
xnor U9204 (N_9204,N_8639,N_8576);
nor U9205 (N_9205,N_8366,N_8066);
nor U9206 (N_9206,N_8505,N_8452);
nand U9207 (N_9207,N_8061,N_8103);
and U9208 (N_9208,N_8917,N_8974);
nand U9209 (N_9209,N_8997,N_8852);
nor U9210 (N_9210,N_8133,N_8308);
xor U9211 (N_9211,N_8567,N_8865);
and U9212 (N_9212,N_8434,N_8242);
and U9213 (N_9213,N_8345,N_8839);
nor U9214 (N_9214,N_8244,N_8160);
xor U9215 (N_9215,N_8184,N_8650);
or U9216 (N_9216,N_8149,N_8011);
and U9217 (N_9217,N_8190,N_8866);
xnor U9218 (N_9218,N_8955,N_8275);
or U9219 (N_9219,N_8392,N_8053);
nor U9220 (N_9220,N_8328,N_8208);
and U9221 (N_9221,N_8127,N_8001);
nor U9222 (N_9222,N_8024,N_8901);
xor U9223 (N_9223,N_8748,N_8438);
or U9224 (N_9224,N_8258,N_8686);
xor U9225 (N_9225,N_8278,N_8016);
xnor U9226 (N_9226,N_8316,N_8537);
and U9227 (N_9227,N_8649,N_8701);
nor U9228 (N_9228,N_8163,N_8990);
nor U9229 (N_9229,N_8179,N_8982);
nand U9230 (N_9230,N_8719,N_8088);
nand U9231 (N_9231,N_8454,N_8528);
nand U9232 (N_9232,N_8745,N_8181);
or U9233 (N_9233,N_8584,N_8994);
and U9234 (N_9234,N_8766,N_8527);
nand U9235 (N_9235,N_8115,N_8962);
nand U9236 (N_9236,N_8755,N_8494);
xnor U9237 (N_9237,N_8631,N_8685);
or U9238 (N_9238,N_8661,N_8959);
xnor U9239 (N_9239,N_8093,N_8314);
xor U9240 (N_9240,N_8003,N_8219);
nor U9241 (N_9241,N_8969,N_8794);
and U9242 (N_9242,N_8139,N_8294);
nand U9243 (N_9243,N_8853,N_8269);
xor U9244 (N_9244,N_8038,N_8225);
nor U9245 (N_9245,N_8395,N_8946);
nand U9246 (N_9246,N_8026,N_8604);
xor U9247 (N_9247,N_8758,N_8814);
and U9248 (N_9248,N_8780,N_8663);
xor U9249 (N_9249,N_8658,N_8868);
or U9250 (N_9250,N_8468,N_8154);
and U9251 (N_9251,N_8401,N_8044);
nand U9252 (N_9252,N_8555,N_8114);
and U9253 (N_9253,N_8302,N_8808);
nand U9254 (N_9254,N_8462,N_8151);
xnor U9255 (N_9255,N_8882,N_8461);
nand U9256 (N_9256,N_8813,N_8963);
and U9257 (N_9257,N_8503,N_8822);
or U9258 (N_9258,N_8175,N_8546);
xnor U9259 (N_9259,N_8543,N_8574);
or U9260 (N_9260,N_8565,N_8943);
nor U9261 (N_9261,N_8247,N_8385);
nand U9262 (N_9262,N_8423,N_8456);
or U9263 (N_9263,N_8253,N_8159);
and U9264 (N_9264,N_8359,N_8790);
or U9265 (N_9265,N_8415,N_8377);
or U9266 (N_9266,N_8464,N_8857);
or U9267 (N_9267,N_8031,N_8611);
and U9268 (N_9268,N_8601,N_8598);
xor U9269 (N_9269,N_8010,N_8005);
or U9270 (N_9270,N_8463,N_8211);
and U9271 (N_9271,N_8202,N_8165);
or U9272 (N_9272,N_8290,N_8169);
or U9273 (N_9273,N_8967,N_8552);
and U9274 (N_9274,N_8579,N_8821);
or U9275 (N_9275,N_8318,N_8817);
xor U9276 (N_9276,N_8380,N_8926);
nor U9277 (N_9277,N_8693,N_8542);
or U9278 (N_9278,N_8319,N_8013);
and U9279 (N_9279,N_8027,N_8829);
and U9280 (N_9280,N_8283,N_8070);
or U9281 (N_9281,N_8932,N_8975);
nor U9282 (N_9282,N_8204,N_8691);
xnor U9283 (N_9283,N_8724,N_8083);
xor U9284 (N_9284,N_8889,N_8096);
or U9285 (N_9285,N_8339,N_8534);
xor U9286 (N_9286,N_8489,N_8526);
xnor U9287 (N_9287,N_8167,N_8090);
nand U9288 (N_9288,N_8518,N_8948);
xor U9289 (N_9289,N_8871,N_8605);
xor U9290 (N_9290,N_8444,N_8532);
xor U9291 (N_9291,N_8887,N_8152);
or U9292 (N_9292,N_8696,N_8375);
xnor U9293 (N_9293,N_8599,N_8199);
or U9294 (N_9294,N_8784,N_8422);
xnor U9295 (N_9295,N_8092,N_8447);
nand U9296 (N_9296,N_8603,N_8135);
and U9297 (N_9297,N_8986,N_8768);
or U9298 (N_9298,N_8330,N_8226);
nand U9299 (N_9299,N_8372,N_8270);
nor U9300 (N_9300,N_8268,N_8898);
nor U9301 (N_9301,N_8086,N_8770);
xnor U9302 (N_9302,N_8406,N_8664);
or U9303 (N_9303,N_8750,N_8970);
xnor U9304 (N_9304,N_8809,N_8578);
nand U9305 (N_9305,N_8140,N_8708);
or U9306 (N_9306,N_8937,N_8138);
nor U9307 (N_9307,N_8647,N_8432);
nand U9308 (N_9308,N_8217,N_8800);
and U9309 (N_9309,N_8529,N_8781);
nand U9310 (N_9310,N_8060,N_8426);
and U9311 (N_9311,N_8945,N_8978);
xor U9312 (N_9312,N_8326,N_8411);
nand U9313 (N_9313,N_8968,N_8303);
xnor U9314 (N_9314,N_8723,N_8538);
or U9315 (N_9315,N_8325,N_8731);
xor U9316 (N_9316,N_8470,N_8097);
or U9317 (N_9317,N_8837,N_8369);
xor U9318 (N_9318,N_8004,N_8908);
xor U9319 (N_9319,N_8018,N_8104);
or U9320 (N_9320,N_8703,N_8445);
xnor U9321 (N_9321,N_8620,N_8998);
nand U9322 (N_9322,N_8034,N_8764);
and U9323 (N_9323,N_8266,N_8515);
or U9324 (N_9324,N_8101,N_8098);
or U9325 (N_9325,N_8753,N_8435);
nand U9326 (N_9326,N_8033,N_8679);
and U9327 (N_9327,N_8157,N_8168);
and U9328 (N_9328,N_8403,N_8028);
or U9329 (N_9329,N_8918,N_8973);
nand U9330 (N_9330,N_8124,N_8801);
or U9331 (N_9331,N_8517,N_8900);
nand U9332 (N_9332,N_8642,N_8331);
or U9333 (N_9333,N_8757,N_8059);
or U9334 (N_9334,N_8072,N_8058);
or U9335 (N_9335,N_8039,N_8906);
and U9336 (N_9336,N_8709,N_8677);
nand U9337 (N_9337,N_8727,N_8589);
nor U9338 (N_9338,N_8697,N_8257);
and U9339 (N_9339,N_8320,N_8249);
and U9340 (N_9340,N_8206,N_8413);
or U9341 (N_9341,N_8015,N_8911);
and U9342 (N_9342,N_8773,N_8363);
xor U9343 (N_9343,N_8936,N_8544);
nor U9344 (N_9344,N_8414,N_8861);
nor U9345 (N_9345,N_8129,N_8450);
xor U9346 (N_9346,N_8109,N_8651);
nand U9347 (N_9347,N_8711,N_8625);
nand U9348 (N_9348,N_8695,N_8924);
nand U9349 (N_9349,N_8077,N_8032);
or U9350 (N_9350,N_8923,N_8193);
and U9351 (N_9351,N_8131,N_8681);
and U9352 (N_9352,N_8209,N_8323);
or U9353 (N_9353,N_8881,N_8246);
or U9354 (N_9354,N_8630,N_8763);
nor U9355 (N_9355,N_8344,N_8433);
or U9356 (N_9356,N_8729,N_8656);
or U9357 (N_9357,N_8988,N_8919);
nor U9358 (N_9358,N_8391,N_8453);
nor U9359 (N_9359,N_8942,N_8683);
nand U9360 (N_9360,N_8128,N_8064);
and U9361 (N_9361,N_8803,N_8682);
xor U9362 (N_9362,N_8113,N_8716);
or U9363 (N_9363,N_8607,N_8022);
nor U9364 (N_9364,N_8944,N_8637);
nand U9365 (N_9365,N_8953,N_8449);
and U9366 (N_9366,N_8272,N_8036);
and U9367 (N_9367,N_8457,N_8828);
nor U9368 (N_9368,N_8309,N_8856);
or U9369 (N_9369,N_8736,N_8223);
nand U9370 (N_9370,N_8295,N_8880);
nand U9371 (N_9371,N_8722,N_8245);
nand U9372 (N_9372,N_8792,N_8049);
nor U9373 (N_9373,N_8051,N_8466);
nand U9374 (N_9374,N_8583,N_8368);
and U9375 (N_9375,N_8074,N_8950);
nor U9376 (N_9376,N_8425,N_8874);
nor U9377 (N_9377,N_8176,N_8312);
nand U9378 (N_9378,N_8035,N_8007);
nand U9379 (N_9379,N_8834,N_8580);
xnor U9380 (N_9380,N_8867,N_8293);
and U9381 (N_9381,N_8390,N_8485);
and U9382 (N_9382,N_8474,N_8712);
nor U9383 (N_9383,N_8381,N_8221);
or U9384 (N_9384,N_8379,N_8079);
nand U9385 (N_9385,N_8671,N_8568);
nor U9386 (N_9386,N_8192,N_8858);
nand U9387 (N_9387,N_8238,N_8860);
nand U9388 (N_9388,N_8118,N_8523);
xor U9389 (N_9389,N_8930,N_8799);
nor U9390 (N_9390,N_8514,N_8407);
and U9391 (N_9391,N_8048,N_8545);
nand U9392 (N_9392,N_8430,N_8126);
and U9393 (N_9393,N_8241,N_8437);
or U9394 (N_9394,N_8707,N_8173);
or U9395 (N_9395,N_8478,N_8976);
and U9396 (N_9396,N_8000,N_8989);
nand U9397 (N_9397,N_8830,N_8386);
nor U9398 (N_9398,N_8504,N_8490);
or U9399 (N_9399,N_8648,N_8897);
nand U9400 (N_9400,N_8912,N_8306);
or U9401 (N_9401,N_8234,N_8846);
nand U9402 (N_9402,N_8913,N_8335);
nand U9403 (N_9403,N_8037,N_8979);
and U9404 (N_9404,N_8590,N_8566);
or U9405 (N_9405,N_8002,N_8194);
nand U9406 (N_9406,N_8210,N_8965);
and U9407 (N_9407,N_8655,N_8043);
xor U9408 (N_9408,N_8144,N_8404);
xnor U9409 (N_9409,N_8849,N_8493);
or U9410 (N_9410,N_8305,N_8056);
and U9411 (N_9411,N_8513,N_8420);
nor U9412 (N_9412,N_8465,N_8659);
xnor U9413 (N_9413,N_8690,N_8229);
and U9414 (N_9414,N_8376,N_8689);
nor U9415 (N_9415,N_8842,N_8484);
and U9416 (N_9416,N_8622,N_8564);
nor U9417 (N_9417,N_8360,N_8460);
nand U9418 (N_9418,N_8876,N_8052);
and U9419 (N_9419,N_8721,N_8351);
nor U9420 (N_9420,N_8512,N_8762);
xor U9421 (N_9421,N_8756,N_8281);
or U9422 (N_9422,N_8235,N_8586);
or U9423 (N_9423,N_8608,N_8558);
nand U9424 (N_9424,N_8941,N_8353);
nor U9425 (N_9425,N_8907,N_8746);
nand U9426 (N_9426,N_8227,N_8667);
or U9427 (N_9427,N_8078,N_8826);
and U9428 (N_9428,N_8606,N_8702);
xor U9429 (N_9429,N_8761,N_8271);
and U9430 (N_9430,N_8397,N_8313);
or U9431 (N_9431,N_8890,N_8117);
xnor U9432 (N_9432,N_8482,N_8660);
and U9433 (N_9433,N_8185,N_8099);
nor U9434 (N_9434,N_8243,N_8198);
xnor U9435 (N_9435,N_8054,N_8084);
or U9436 (N_9436,N_8267,N_8205);
xnor U9437 (N_9437,N_8020,N_8884);
nand U9438 (N_9438,N_8102,N_8068);
nor U9439 (N_9439,N_8348,N_8164);
nor U9440 (N_9440,N_8995,N_8170);
nor U9441 (N_9441,N_8836,N_8479);
nor U9442 (N_9442,N_8643,N_8212);
and U9443 (N_9443,N_8847,N_8812);
and U9444 (N_9444,N_8956,N_8100);
xnor U9445 (N_9445,N_8934,N_8615);
xnor U9446 (N_9446,N_8797,N_8996);
nand U9447 (N_9447,N_8075,N_8162);
or U9448 (N_9448,N_8340,N_8254);
or U9449 (N_9449,N_8741,N_8122);
xnor U9450 (N_9450,N_8250,N_8336);
nor U9451 (N_9451,N_8832,N_8592);
nor U9452 (N_9452,N_8356,N_8947);
or U9453 (N_9453,N_8623,N_8831);
or U9454 (N_9454,N_8230,N_8261);
or U9455 (N_9455,N_8014,N_8476);
and U9456 (N_9456,N_8273,N_8785);
nand U9457 (N_9457,N_8087,N_8863);
and U9458 (N_9458,N_8551,N_8410);
or U9459 (N_9459,N_8334,N_8715);
nand U9460 (N_9460,N_8291,N_8811);
xnor U9461 (N_9461,N_8531,N_8516);
nand U9462 (N_9462,N_8771,N_8373);
xor U9463 (N_9463,N_8992,N_8017);
and U9464 (N_9464,N_8023,N_8904);
nand U9465 (N_9465,N_8732,N_8393);
xor U9466 (N_9466,N_8443,N_8807);
nand U9467 (N_9467,N_8405,N_8252);
and U9468 (N_9468,N_8692,N_8497);
and U9469 (N_9469,N_8367,N_8816);
nor U9470 (N_9470,N_8819,N_8678);
xor U9471 (N_9471,N_8141,N_8178);
and U9472 (N_9472,N_8394,N_8793);
nor U9473 (N_9473,N_8180,N_8040);
nor U9474 (N_9474,N_8921,N_8802);
and U9475 (N_9475,N_8333,N_8744);
nor U9476 (N_9476,N_8361,N_8931);
nor U9477 (N_9477,N_8769,N_8006);
xor U9478 (N_9478,N_8383,N_8961);
nor U9479 (N_9479,N_8571,N_8343);
nand U9480 (N_9480,N_8197,N_8350);
nor U9481 (N_9481,N_8524,N_8451);
or U9482 (N_9482,N_8952,N_8108);
xnor U9483 (N_9483,N_8964,N_8304);
nor U9484 (N_9484,N_8362,N_8935);
and U9485 (N_9485,N_8365,N_8618);
nor U9486 (N_9486,N_8477,N_8894);
nor U9487 (N_9487,N_8063,N_8698);
xor U9488 (N_9488,N_8806,N_8706);
or U9489 (N_9489,N_8914,N_8899);
nand U9490 (N_9490,N_8481,N_8327);
xor U9491 (N_9491,N_8091,N_8854);
nand U9492 (N_9492,N_8448,N_8073);
nor U9493 (N_9493,N_8600,N_8228);
or U9494 (N_9494,N_8896,N_8125);
nand U9495 (N_9495,N_8877,N_8050);
or U9496 (N_9496,N_8256,N_8735);
and U9497 (N_9497,N_8107,N_8130);
and U9498 (N_9498,N_8610,N_8737);
nand U9499 (N_9499,N_8738,N_8991);
and U9500 (N_9500,N_8539,N_8812);
nand U9501 (N_9501,N_8795,N_8957);
nand U9502 (N_9502,N_8510,N_8881);
nand U9503 (N_9503,N_8624,N_8399);
or U9504 (N_9504,N_8518,N_8271);
and U9505 (N_9505,N_8796,N_8105);
nand U9506 (N_9506,N_8314,N_8197);
and U9507 (N_9507,N_8843,N_8379);
xnor U9508 (N_9508,N_8439,N_8713);
nand U9509 (N_9509,N_8419,N_8789);
nor U9510 (N_9510,N_8526,N_8999);
and U9511 (N_9511,N_8630,N_8609);
and U9512 (N_9512,N_8708,N_8704);
and U9513 (N_9513,N_8574,N_8435);
xnor U9514 (N_9514,N_8572,N_8185);
and U9515 (N_9515,N_8508,N_8332);
or U9516 (N_9516,N_8222,N_8696);
and U9517 (N_9517,N_8983,N_8553);
nand U9518 (N_9518,N_8012,N_8691);
nor U9519 (N_9519,N_8952,N_8717);
nor U9520 (N_9520,N_8158,N_8019);
nor U9521 (N_9521,N_8567,N_8589);
nand U9522 (N_9522,N_8914,N_8327);
and U9523 (N_9523,N_8867,N_8346);
or U9524 (N_9524,N_8307,N_8531);
nand U9525 (N_9525,N_8873,N_8070);
or U9526 (N_9526,N_8343,N_8107);
xor U9527 (N_9527,N_8599,N_8489);
xor U9528 (N_9528,N_8130,N_8281);
nor U9529 (N_9529,N_8125,N_8482);
nor U9530 (N_9530,N_8051,N_8374);
xnor U9531 (N_9531,N_8115,N_8343);
nand U9532 (N_9532,N_8728,N_8184);
nand U9533 (N_9533,N_8754,N_8949);
nand U9534 (N_9534,N_8283,N_8586);
or U9535 (N_9535,N_8810,N_8031);
nand U9536 (N_9536,N_8128,N_8364);
nand U9537 (N_9537,N_8760,N_8951);
xnor U9538 (N_9538,N_8796,N_8985);
nor U9539 (N_9539,N_8487,N_8117);
nor U9540 (N_9540,N_8507,N_8217);
nand U9541 (N_9541,N_8418,N_8040);
or U9542 (N_9542,N_8999,N_8961);
xor U9543 (N_9543,N_8310,N_8869);
nand U9544 (N_9544,N_8616,N_8902);
nor U9545 (N_9545,N_8560,N_8513);
and U9546 (N_9546,N_8161,N_8483);
or U9547 (N_9547,N_8822,N_8236);
and U9548 (N_9548,N_8308,N_8854);
and U9549 (N_9549,N_8879,N_8972);
nor U9550 (N_9550,N_8633,N_8755);
nand U9551 (N_9551,N_8140,N_8315);
xor U9552 (N_9552,N_8553,N_8941);
xnor U9553 (N_9553,N_8788,N_8321);
nand U9554 (N_9554,N_8783,N_8053);
xor U9555 (N_9555,N_8837,N_8655);
xor U9556 (N_9556,N_8041,N_8712);
or U9557 (N_9557,N_8240,N_8829);
nand U9558 (N_9558,N_8443,N_8984);
xor U9559 (N_9559,N_8173,N_8078);
nor U9560 (N_9560,N_8472,N_8397);
xor U9561 (N_9561,N_8022,N_8073);
and U9562 (N_9562,N_8213,N_8474);
xnor U9563 (N_9563,N_8174,N_8315);
xnor U9564 (N_9564,N_8644,N_8711);
nand U9565 (N_9565,N_8472,N_8897);
or U9566 (N_9566,N_8757,N_8650);
or U9567 (N_9567,N_8090,N_8905);
xnor U9568 (N_9568,N_8167,N_8940);
nor U9569 (N_9569,N_8976,N_8150);
xnor U9570 (N_9570,N_8708,N_8378);
and U9571 (N_9571,N_8608,N_8572);
nor U9572 (N_9572,N_8641,N_8187);
xor U9573 (N_9573,N_8428,N_8018);
or U9574 (N_9574,N_8712,N_8441);
nand U9575 (N_9575,N_8765,N_8613);
and U9576 (N_9576,N_8936,N_8438);
nand U9577 (N_9577,N_8188,N_8993);
xor U9578 (N_9578,N_8423,N_8686);
and U9579 (N_9579,N_8759,N_8962);
nor U9580 (N_9580,N_8795,N_8425);
xnor U9581 (N_9581,N_8283,N_8217);
nand U9582 (N_9582,N_8395,N_8228);
and U9583 (N_9583,N_8825,N_8411);
and U9584 (N_9584,N_8757,N_8067);
nor U9585 (N_9585,N_8342,N_8971);
nor U9586 (N_9586,N_8918,N_8268);
and U9587 (N_9587,N_8041,N_8955);
and U9588 (N_9588,N_8669,N_8819);
nand U9589 (N_9589,N_8355,N_8174);
or U9590 (N_9590,N_8398,N_8761);
or U9591 (N_9591,N_8791,N_8285);
nor U9592 (N_9592,N_8994,N_8222);
nor U9593 (N_9593,N_8916,N_8640);
xnor U9594 (N_9594,N_8796,N_8405);
nor U9595 (N_9595,N_8687,N_8405);
and U9596 (N_9596,N_8318,N_8200);
nor U9597 (N_9597,N_8900,N_8622);
and U9598 (N_9598,N_8784,N_8523);
and U9599 (N_9599,N_8307,N_8816);
xnor U9600 (N_9600,N_8165,N_8534);
nand U9601 (N_9601,N_8306,N_8661);
xor U9602 (N_9602,N_8289,N_8159);
and U9603 (N_9603,N_8007,N_8966);
or U9604 (N_9604,N_8897,N_8559);
and U9605 (N_9605,N_8886,N_8556);
nor U9606 (N_9606,N_8392,N_8945);
nor U9607 (N_9607,N_8558,N_8936);
or U9608 (N_9608,N_8284,N_8475);
nor U9609 (N_9609,N_8758,N_8968);
nand U9610 (N_9610,N_8564,N_8285);
nor U9611 (N_9611,N_8756,N_8224);
or U9612 (N_9612,N_8013,N_8678);
and U9613 (N_9613,N_8567,N_8387);
and U9614 (N_9614,N_8357,N_8732);
nand U9615 (N_9615,N_8089,N_8687);
nor U9616 (N_9616,N_8309,N_8148);
nor U9617 (N_9617,N_8127,N_8153);
nand U9618 (N_9618,N_8340,N_8946);
or U9619 (N_9619,N_8580,N_8450);
nor U9620 (N_9620,N_8175,N_8256);
nor U9621 (N_9621,N_8034,N_8749);
or U9622 (N_9622,N_8487,N_8574);
or U9623 (N_9623,N_8547,N_8240);
or U9624 (N_9624,N_8700,N_8213);
or U9625 (N_9625,N_8610,N_8979);
nor U9626 (N_9626,N_8894,N_8201);
nor U9627 (N_9627,N_8628,N_8265);
nand U9628 (N_9628,N_8994,N_8524);
xor U9629 (N_9629,N_8469,N_8219);
nand U9630 (N_9630,N_8118,N_8289);
and U9631 (N_9631,N_8687,N_8401);
and U9632 (N_9632,N_8520,N_8869);
xor U9633 (N_9633,N_8028,N_8514);
xnor U9634 (N_9634,N_8569,N_8728);
xor U9635 (N_9635,N_8492,N_8090);
nor U9636 (N_9636,N_8116,N_8560);
xnor U9637 (N_9637,N_8064,N_8724);
nand U9638 (N_9638,N_8894,N_8963);
or U9639 (N_9639,N_8138,N_8972);
nor U9640 (N_9640,N_8342,N_8055);
and U9641 (N_9641,N_8714,N_8068);
or U9642 (N_9642,N_8950,N_8543);
nand U9643 (N_9643,N_8553,N_8234);
and U9644 (N_9644,N_8815,N_8094);
nand U9645 (N_9645,N_8921,N_8306);
nor U9646 (N_9646,N_8447,N_8636);
and U9647 (N_9647,N_8685,N_8888);
nand U9648 (N_9648,N_8048,N_8584);
and U9649 (N_9649,N_8877,N_8488);
nand U9650 (N_9650,N_8170,N_8684);
xor U9651 (N_9651,N_8552,N_8746);
or U9652 (N_9652,N_8638,N_8904);
and U9653 (N_9653,N_8671,N_8199);
xnor U9654 (N_9654,N_8159,N_8714);
nor U9655 (N_9655,N_8445,N_8270);
nand U9656 (N_9656,N_8719,N_8595);
or U9657 (N_9657,N_8267,N_8328);
nor U9658 (N_9658,N_8207,N_8732);
xnor U9659 (N_9659,N_8678,N_8655);
or U9660 (N_9660,N_8344,N_8214);
and U9661 (N_9661,N_8890,N_8708);
or U9662 (N_9662,N_8994,N_8758);
nand U9663 (N_9663,N_8164,N_8128);
nor U9664 (N_9664,N_8147,N_8645);
and U9665 (N_9665,N_8804,N_8721);
nor U9666 (N_9666,N_8591,N_8183);
and U9667 (N_9667,N_8120,N_8982);
and U9668 (N_9668,N_8676,N_8585);
nor U9669 (N_9669,N_8787,N_8126);
or U9670 (N_9670,N_8024,N_8034);
nand U9671 (N_9671,N_8155,N_8944);
nor U9672 (N_9672,N_8654,N_8169);
or U9673 (N_9673,N_8649,N_8408);
nand U9674 (N_9674,N_8185,N_8129);
nand U9675 (N_9675,N_8082,N_8071);
or U9676 (N_9676,N_8773,N_8770);
and U9677 (N_9677,N_8782,N_8632);
xor U9678 (N_9678,N_8460,N_8681);
and U9679 (N_9679,N_8635,N_8390);
or U9680 (N_9680,N_8578,N_8774);
or U9681 (N_9681,N_8222,N_8226);
xnor U9682 (N_9682,N_8642,N_8134);
nor U9683 (N_9683,N_8228,N_8993);
or U9684 (N_9684,N_8778,N_8839);
nand U9685 (N_9685,N_8936,N_8858);
nor U9686 (N_9686,N_8624,N_8436);
nand U9687 (N_9687,N_8538,N_8172);
or U9688 (N_9688,N_8511,N_8962);
xor U9689 (N_9689,N_8291,N_8116);
and U9690 (N_9690,N_8339,N_8801);
nor U9691 (N_9691,N_8480,N_8818);
nand U9692 (N_9692,N_8629,N_8001);
nor U9693 (N_9693,N_8384,N_8218);
and U9694 (N_9694,N_8459,N_8085);
or U9695 (N_9695,N_8018,N_8921);
nor U9696 (N_9696,N_8158,N_8986);
or U9697 (N_9697,N_8439,N_8586);
xnor U9698 (N_9698,N_8349,N_8561);
or U9699 (N_9699,N_8409,N_8448);
nor U9700 (N_9700,N_8484,N_8070);
xor U9701 (N_9701,N_8075,N_8455);
xnor U9702 (N_9702,N_8739,N_8477);
xnor U9703 (N_9703,N_8027,N_8784);
nand U9704 (N_9704,N_8139,N_8213);
xor U9705 (N_9705,N_8071,N_8794);
or U9706 (N_9706,N_8478,N_8523);
or U9707 (N_9707,N_8980,N_8426);
nand U9708 (N_9708,N_8421,N_8675);
and U9709 (N_9709,N_8220,N_8628);
or U9710 (N_9710,N_8987,N_8888);
and U9711 (N_9711,N_8751,N_8789);
and U9712 (N_9712,N_8452,N_8439);
nand U9713 (N_9713,N_8539,N_8988);
nor U9714 (N_9714,N_8255,N_8427);
nor U9715 (N_9715,N_8337,N_8651);
and U9716 (N_9716,N_8399,N_8900);
xor U9717 (N_9717,N_8777,N_8730);
nor U9718 (N_9718,N_8884,N_8572);
nor U9719 (N_9719,N_8355,N_8035);
or U9720 (N_9720,N_8457,N_8034);
or U9721 (N_9721,N_8564,N_8153);
xnor U9722 (N_9722,N_8986,N_8925);
xnor U9723 (N_9723,N_8249,N_8445);
and U9724 (N_9724,N_8964,N_8380);
nor U9725 (N_9725,N_8809,N_8803);
nand U9726 (N_9726,N_8876,N_8745);
nand U9727 (N_9727,N_8160,N_8546);
xnor U9728 (N_9728,N_8008,N_8468);
and U9729 (N_9729,N_8052,N_8396);
nand U9730 (N_9730,N_8509,N_8355);
nand U9731 (N_9731,N_8820,N_8088);
nand U9732 (N_9732,N_8323,N_8380);
and U9733 (N_9733,N_8914,N_8455);
nor U9734 (N_9734,N_8178,N_8303);
nand U9735 (N_9735,N_8214,N_8856);
xor U9736 (N_9736,N_8297,N_8497);
nor U9737 (N_9737,N_8855,N_8487);
xor U9738 (N_9738,N_8971,N_8430);
nand U9739 (N_9739,N_8417,N_8834);
xnor U9740 (N_9740,N_8497,N_8997);
nor U9741 (N_9741,N_8421,N_8347);
and U9742 (N_9742,N_8690,N_8277);
xnor U9743 (N_9743,N_8249,N_8814);
or U9744 (N_9744,N_8454,N_8565);
nand U9745 (N_9745,N_8722,N_8050);
nor U9746 (N_9746,N_8901,N_8767);
nor U9747 (N_9747,N_8059,N_8459);
and U9748 (N_9748,N_8546,N_8933);
nand U9749 (N_9749,N_8953,N_8591);
xor U9750 (N_9750,N_8165,N_8066);
nand U9751 (N_9751,N_8294,N_8846);
or U9752 (N_9752,N_8833,N_8943);
and U9753 (N_9753,N_8419,N_8455);
nand U9754 (N_9754,N_8271,N_8592);
nand U9755 (N_9755,N_8478,N_8695);
xnor U9756 (N_9756,N_8988,N_8052);
and U9757 (N_9757,N_8073,N_8881);
nor U9758 (N_9758,N_8295,N_8986);
nor U9759 (N_9759,N_8637,N_8923);
nor U9760 (N_9760,N_8825,N_8368);
xnor U9761 (N_9761,N_8020,N_8956);
xnor U9762 (N_9762,N_8790,N_8287);
and U9763 (N_9763,N_8103,N_8181);
or U9764 (N_9764,N_8295,N_8572);
or U9765 (N_9765,N_8956,N_8916);
nor U9766 (N_9766,N_8232,N_8415);
nand U9767 (N_9767,N_8313,N_8436);
nand U9768 (N_9768,N_8805,N_8729);
or U9769 (N_9769,N_8892,N_8827);
nor U9770 (N_9770,N_8731,N_8709);
xor U9771 (N_9771,N_8028,N_8198);
nor U9772 (N_9772,N_8028,N_8337);
and U9773 (N_9773,N_8779,N_8858);
and U9774 (N_9774,N_8508,N_8311);
or U9775 (N_9775,N_8051,N_8332);
and U9776 (N_9776,N_8318,N_8791);
nand U9777 (N_9777,N_8051,N_8426);
and U9778 (N_9778,N_8887,N_8820);
xnor U9779 (N_9779,N_8773,N_8439);
nor U9780 (N_9780,N_8255,N_8125);
and U9781 (N_9781,N_8042,N_8669);
nor U9782 (N_9782,N_8970,N_8638);
or U9783 (N_9783,N_8757,N_8349);
xnor U9784 (N_9784,N_8042,N_8236);
and U9785 (N_9785,N_8000,N_8020);
nor U9786 (N_9786,N_8325,N_8773);
and U9787 (N_9787,N_8835,N_8005);
xor U9788 (N_9788,N_8329,N_8724);
and U9789 (N_9789,N_8007,N_8798);
and U9790 (N_9790,N_8339,N_8076);
nor U9791 (N_9791,N_8940,N_8468);
nand U9792 (N_9792,N_8191,N_8130);
nand U9793 (N_9793,N_8638,N_8376);
xnor U9794 (N_9794,N_8103,N_8748);
nor U9795 (N_9795,N_8662,N_8746);
or U9796 (N_9796,N_8297,N_8627);
and U9797 (N_9797,N_8612,N_8205);
xnor U9798 (N_9798,N_8037,N_8101);
and U9799 (N_9799,N_8855,N_8119);
nor U9800 (N_9800,N_8884,N_8231);
and U9801 (N_9801,N_8733,N_8837);
nor U9802 (N_9802,N_8634,N_8686);
nand U9803 (N_9803,N_8979,N_8836);
nand U9804 (N_9804,N_8636,N_8870);
nor U9805 (N_9805,N_8785,N_8746);
xnor U9806 (N_9806,N_8817,N_8241);
xor U9807 (N_9807,N_8206,N_8501);
nand U9808 (N_9808,N_8631,N_8834);
or U9809 (N_9809,N_8392,N_8773);
or U9810 (N_9810,N_8914,N_8446);
nand U9811 (N_9811,N_8255,N_8702);
nand U9812 (N_9812,N_8320,N_8948);
or U9813 (N_9813,N_8865,N_8104);
nor U9814 (N_9814,N_8001,N_8549);
xnor U9815 (N_9815,N_8063,N_8029);
and U9816 (N_9816,N_8265,N_8712);
nand U9817 (N_9817,N_8736,N_8590);
xor U9818 (N_9818,N_8566,N_8150);
xor U9819 (N_9819,N_8140,N_8170);
or U9820 (N_9820,N_8781,N_8636);
and U9821 (N_9821,N_8530,N_8071);
nand U9822 (N_9822,N_8526,N_8122);
xor U9823 (N_9823,N_8232,N_8204);
or U9824 (N_9824,N_8014,N_8423);
and U9825 (N_9825,N_8003,N_8222);
and U9826 (N_9826,N_8918,N_8799);
nor U9827 (N_9827,N_8879,N_8200);
nor U9828 (N_9828,N_8265,N_8077);
xor U9829 (N_9829,N_8825,N_8841);
xor U9830 (N_9830,N_8580,N_8424);
nand U9831 (N_9831,N_8707,N_8541);
nand U9832 (N_9832,N_8345,N_8861);
and U9833 (N_9833,N_8101,N_8271);
and U9834 (N_9834,N_8167,N_8146);
or U9835 (N_9835,N_8822,N_8862);
and U9836 (N_9836,N_8343,N_8184);
xor U9837 (N_9837,N_8864,N_8059);
and U9838 (N_9838,N_8836,N_8629);
nand U9839 (N_9839,N_8682,N_8655);
nor U9840 (N_9840,N_8462,N_8587);
nor U9841 (N_9841,N_8627,N_8912);
and U9842 (N_9842,N_8644,N_8991);
xnor U9843 (N_9843,N_8516,N_8310);
and U9844 (N_9844,N_8824,N_8934);
nor U9845 (N_9845,N_8735,N_8186);
or U9846 (N_9846,N_8886,N_8814);
xor U9847 (N_9847,N_8065,N_8246);
nor U9848 (N_9848,N_8436,N_8156);
nor U9849 (N_9849,N_8242,N_8117);
and U9850 (N_9850,N_8300,N_8997);
nand U9851 (N_9851,N_8726,N_8524);
nand U9852 (N_9852,N_8045,N_8519);
nand U9853 (N_9853,N_8579,N_8887);
nand U9854 (N_9854,N_8029,N_8812);
xor U9855 (N_9855,N_8529,N_8456);
nand U9856 (N_9856,N_8050,N_8499);
nor U9857 (N_9857,N_8521,N_8258);
and U9858 (N_9858,N_8232,N_8586);
xor U9859 (N_9859,N_8712,N_8058);
or U9860 (N_9860,N_8202,N_8112);
and U9861 (N_9861,N_8750,N_8422);
xor U9862 (N_9862,N_8450,N_8279);
nand U9863 (N_9863,N_8535,N_8859);
or U9864 (N_9864,N_8640,N_8744);
nor U9865 (N_9865,N_8533,N_8779);
nand U9866 (N_9866,N_8580,N_8887);
and U9867 (N_9867,N_8120,N_8361);
xnor U9868 (N_9868,N_8744,N_8963);
or U9869 (N_9869,N_8352,N_8047);
nor U9870 (N_9870,N_8538,N_8695);
nand U9871 (N_9871,N_8602,N_8597);
nand U9872 (N_9872,N_8737,N_8077);
nor U9873 (N_9873,N_8431,N_8377);
and U9874 (N_9874,N_8825,N_8471);
xnor U9875 (N_9875,N_8641,N_8276);
or U9876 (N_9876,N_8891,N_8444);
nand U9877 (N_9877,N_8426,N_8087);
nor U9878 (N_9878,N_8643,N_8769);
nor U9879 (N_9879,N_8827,N_8168);
nor U9880 (N_9880,N_8821,N_8442);
xnor U9881 (N_9881,N_8245,N_8581);
nand U9882 (N_9882,N_8577,N_8983);
and U9883 (N_9883,N_8393,N_8210);
xnor U9884 (N_9884,N_8657,N_8588);
xnor U9885 (N_9885,N_8155,N_8759);
nand U9886 (N_9886,N_8158,N_8759);
or U9887 (N_9887,N_8658,N_8134);
nor U9888 (N_9888,N_8721,N_8371);
xor U9889 (N_9889,N_8502,N_8782);
nor U9890 (N_9890,N_8828,N_8398);
nand U9891 (N_9891,N_8057,N_8446);
nor U9892 (N_9892,N_8500,N_8942);
xor U9893 (N_9893,N_8358,N_8728);
nor U9894 (N_9894,N_8911,N_8640);
and U9895 (N_9895,N_8631,N_8170);
xnor U9896 (N_9896,N_8751,N_8137);
nand U9897 (N_9897,N_8152,N_8943);
nor U9898 (N_9898,N_8531,N_8220);
and U9899 (N_9899,N_8778,N_8311);
xor U9900 (N_9900,N_8746,N_8799);
nor U9901 (N_9901,N_8022,N_8035);
nor U9902 (N_9902,N_8617,N_8003);
and U9903 (N_9903,N_8451,N_8153);
nand U9904 (N_9904,N_8098,N_8282);
xnor U9905 (N_9905,N_8876,N_8649);
or U9906 (N_9906,N_8183,N_8758);
and U9907 (N_9907,N_8426,N_8417);
and U9908 (N_9908,N_8519,N_8272);
nand U9909 (N_9909,N_8095,N_8160);
or U9910 (N_9910,N_8721,N_8418);
or U9911 (N_9911,N_8345,N_8737);
xor U9912 (N_9912,N_8899,N_8837);
nand U9913 (N_9913,N_8245,N_8153);
xnor U9914 (N_9914,N_8637,N_8645);
xnor U9915 (N_9915,N_8710,N_8778);
nor U9916 (N_9916,N_8639,N_8049);
nand U9917 (N_9917,N_8789,N_8934);
xnor U9918 (N_9918,N_8765,N_8647);
nor U9919 (N_9919,N_8103,N_8738);
or U9920 (N_9920,N_8595,N_8879);
xor U9921 (N_9921,N_8847,N_8166);
or U9922 (N_9922,N_8646,N_8645);
nand U9923 (N_9923,N_8878,N_8554);
nor U9924 (N_9924,N_8675,N_8608);
nand U9925 (N_9925,N_8154,N_8045);
nor U9926 (N_9926,N_8126,N_8197);
nand U9927 (N_9927,N_8586,N_8739);
nand U9928 (N_9928,N_8060,N_8105);
and U9929 (N_9929,N_8462,N_8804);
nand U9930 (N_9930,N_8961,N_8885);
nor U9931 (N_9931,N_8067,N_8692);
nand U9932 (N_9932,N_8388,N_8597);
and U9933 (N_9933,N_8089,N_8833);
and U9934 (N_9934,N_8396,N_8063);
nand U9935 (N_9935,N_8135,N_8517);
and U9936 (N_9936,N_8085,N_8116);
or U9937 (N_9937,N_8915,N_8590);
and U9938 (N_9938,N_8054,N_8223);
and U9939 (N_9939,N_8612,N_8280);
nand U9940 (N_9940,N_8242,N_8874);
xor U9941 (N_9941,N_8364,N_8785);
or U9942 (N_9942,N_8643,N_8844);
nor U9943 (N_9943,N_8658,N_8889);
xor U9944 (N_9944,N_8535,N_8745);
or U9945 (N_9945,N_8712,N_8475);
xnor U9946 (N_9946,N_8955,N_8326);
xnor U9947 (N_9947,N_8759,N_8383);
and U9948 (N_9948,N_8385,N_8582);
or U9949 (N_9949,N_8725,N_8711);
nor U9950 (N_9950,N_8428,N_8231);
or U9951 (N_9951,N_8544,N_8440);
and U9952 (N_9952,N_8436,N_8093);
or U9953 (N_9953,N_8651,N_8661);
or U9954 (N_9954,N_8976,N_8208);
nor U9955 (N_9955,N_8634,N_8151);
and U9956 (N_9956,N_8841,N_8349);
nor U9957 (N_9957,N_8263,N_8838);
xor U9958 (N_9958,N_8705,N_8640);
xor U9959 (N_9959,N_8963,N_8347);
or U9960 (N_9960,N_8709,N_8826);
nand U9961 (N_9961,N_8418,N_8962);
or U9962 (N_9962,N_8913,N_8729);
xor U9963 (N_9963,N_8446,N_8994);
nand U9964 (N_9964,N_8577,N_8766);
nor U9965 (N_9965,N_8651,N_8006);
or U9966 (N_9966,N_8325,N_8690);
xnor U9967 (N_9967,N_8724,N_8715);
xor U9968 (N_9968,N_8257,N_8686);
nand U9969 (N_9969,N_8942,N_8469);
xor U9970 (N_9970,N_8664,N_8904);
xnor U9971 (N_9971,N_8838,N_8889);
xor U9972 (N_9972,N_8439,N_8126);
or U9973 (N_9973,N_8867,N_8254);
nand U9974 (N_9974,N_8030,N_8907);
xor U9975 (N_9975,N_8308,N_8154);
xor U9976 (N_9976,N_8959,N_8004);
xnor U9977 (N_9977,N_8074,N_8538);
or U9978 (N_9978,N_8871,N_8704);
and U9979 (N_9979,N_8908,N_8378);
nor U9980 (N_9980,N_8659,N_8992);
nor U9981 (N_9981,N_8626,N_8472);
xnor U9982 (N_9982,N_8840,N_8135);
and U9983 (N_9983,N_8262,N_8726);
nand U9984 (N_9984,N_8180,N_8819);
nor U9985 (N_9985,N_8928,N_8925);
or U9986 (N_9986,N_8000,N_8544);
nor U9987 (N_9987,N_8237,N_8705);
or U9988 (N_9988,N_8430,N_8726);
nand U9989 (N_9989,N_8115,N_8967);
xnor U9990 (N_9990,N_8324,N_8781);
or U9991 (N_9991,N_8755,N_8375);
or U9992 (N_9992,N_8239,N_8929);
xor U9993 (N_9993,N_8554,N_8070);
nand U9994 (N_9994,N_8339,N_8527);
nand U9995 (N_9995,N_8662,N_8570);
nand U9996 (N_9996,N_8764,N_8083);
nor U9997 (N_9997,N_8375,N_8125);
xor U9998 (N_9998,N_8247,N_8388);
nand U9999 (N_9999,N_8978,N_8862);
xnor U10000 (N_10000,N_9815,N_9814);
xor U10001 (N_10001,N_9995,N_9497);
xnor U10002 (N_10002,N_9928,N_9415);
or U10003 (N_10003,N_9936,N_9177);
xor U10004 (N_10004,N_9161,N_9571);
xor U10005 (N_10005,N_9195,N_9651);
or U10006 (N_10006,N_9566,N_9961);
xnor U10007 (N_10007,N_9860,N_9862);
xor U10008 (N_10008,N_9238,N_9383);
nor U10009 (N_10009,N_9715,N_9431);
xnor U10010 (N_10010,N_9938,N_9468);
xor U10011 (N_10011,N_9118,N_9285);
and U10012 (N_10012,N_9922,N_9451);
xor U10013 (N_10013,N_9706,N_9012);
nor U10014 (N_10014,N_9899,N_9037);
nor U10015 (N_10015,N_9626,N_9018);
or U10016 (N_10016,N_9467,N_9439);
nand U10017 (N_10017,N_9186,N_9799);
nor U10018 (N_10018,N_9108,N_9833);
nand U10019 (N_10019,N_9463,N_9099);
xnor U10020 (N_10020,N_9386,N_9168);
xnor U10021 (N_10021,N_9137,N_9920);
or U10022 (N_10022,N_9091,N_9424);
and U10023 (N_10023,N_9380,N_9194);
xnor U10024 (N_10024,N_9054,N_9629);
nor U10025 (N_10025,N_9941,N_9311);
nor U10026 (N_10026,N_9314,N_9734);
or U10027 (N_10027,N_9660,N_9900);
nor U10028 (N_10028,N_9109,N_9917);
xnor U10029 (N_10029,N_9374,N_9363);
nor U10030 (N_10030,N_9034,N_9990);
nand U10031 (N_10031,N_9350,N_9332);
or U10032 (N_10032,N_9391,N_9616);
nor U10033 (N_10033,N_9760,N_9965);
xnor U10034 (N_10034,N_9614,N_9838);
nand U10035 (N_10035,N_9071,N_9329);
nand U10036 (N_10036,N_9894,N_9952);
xor U10037 (N_10037,N_9066,N_9130);
and U10038 (N_10038,N_9681,N_9373);
and U10039 (N_10039,N_9261,N_9646);
nor U10040 (N_10040,N_9971,N_9946);
nor U10041 (N_10041,N_9477,N_9306);
nand U10042 (N_10042,N_9086,N_9029);
nor U10043 (N_10043,N_9065,N_9281);
nand U10044 (N_10044,N_9709,N_9419);
nand U10045 (N_10045,N_9169,N_9714);
xnor U10046 (N_10046,N_9693,N_9335);
xor U10047 (N_10047,N_9475,N_9542);
nor U10048 (N_10048,N_9901,N_9111);
xor U10049 (N_10049,N_9540,N_9077);
xor U10050 (N_10050,N_9942,N_9047);
or U10051 (N_10051,N_9509,N_9736);
nor U10052 (N_10052,N_9413,N_9339);
nand U10053 (N_10053,N_9556,N_9960);
nand U10054 (N_10054,N_9215,N_9144);
xnor U10055 (N_10055,N_9817,N_9000);
nand U10056 (N_10056,N_9212,N_9934);
nor U10057 (N_10057,N_9915,N_9425);
nand U10058 (N_10058,N_9871,N_9807);
nor U10059 (N_10059,N_9097,N_9672);
nor U10060 (N_10060,N_9820,N_9800);
nand U10061 (N_10061,N_9684,N_9581);
or U10062 (N_10062,N_9241,N_9909);
xor U10063 (N_10063,N_9361,N_9661);
and U10064 (N_10064,N_9305,N_9919);
and U10065 (N_10065,N_9765,N_9489);
nor U10066 (N_10066,N_9121,N_9666);
nor U10067 (N_10067,N_9787,N_9187);
and U10068 (N_10068,N_9641,N_9006);
xnor U10069 (N_10069,N_9623,N_9893);
or U10070 (N_10070,N_9867,N_9272);
xor U10071 (N_10071,N_9810,N_9764);
or U10072 (N_10072,N_9412,N_9404);
and U10073 (N_10073,N_9989,N_9676);
or U10074 (N_10074,N_9576,N_9014);
nand U10075 (N_10075,N_9779,N_9058);
nand U10076 (N_10076,N_9527,N_9007);
nor U10077 (N_10077,N_9247,N_9310);
or U10078 (N_10078,N_9338,N_9352);
and U10079 (N_10079,N_9520,N_9443);
or U10080 (N_10080,N_9945,N_9165);
nand U10081 (N_10081,N_9392,N_9859);
nor U10082 (N_10082,N_9784,N_9789);
or U10083 (N_10083,N_9745,N_9129);
nand U10084 (N_10084,N_9470,N_9173);
nor U10085 (N_10085,N_9795,N_9019);
nor U10086 (N_10086,N_9251,N_9143);
xor U10087 (N_10087,N_9320,N_9634);
nand U10088 (N_10088,N_9223,N_9600);
nand U10089 (N_10089,N_9858,N_9549);
nand U10090 (N_10090,N_9368,N_9943);
and U10091 (N_10091,N_9399,N_9589);
and U10092 (N_10092,N_9385,N_9691);
xnor U10093 (N_10093,N_9515,N_9429);
and U10094 (N_10094,N_9481,N_9348);
xnor U10095 (N_10095,N_9737,N_9216);
nor U10096 (N_10096,N_9585,N_9035);
xnor U10097 (N_10097,N_9023,N_9716);
xnor U10098 (N_10098,N_9028,N_9975);
nand U10099 (N_10099,N_9752,N_9876);
nand U10100 (N_10100,N_9135,N_9450);
and U10101 (N_10101,N_9844,N_9030);
nand U10102 (N_10102,N_9868,N_9382);
nor U10103 (N_10103,N_9610,N_9983);
nor U10104 (N_10104,N_9703,N_9484);
nand U10105 (N_10105,N_9558,N_9897);
nor U10106 (N_10106,N_9448,N_9776);
and U10107 (N_10107,N_9080,N_9300);
nand U10108 (N_10108,N_9211,N_9466);
nand U10109 (N_10109,N_9455,N_9724);
nor U10110 (N_10110,N_9770,N_9822);
xnor U10111 (N_10111,N_9732,N_9297);
xnor U10112 (N_10112,N_9994,N_9988);
nor U10113 (N_10113,N_9498,N_9793);
nand U10114 (N_10114,N_9541,N_9016);
or U10115 (N_10115,N_9819,N_9355);
xnor U10116 (N_10116,N_9128,N_9171);
and U10117 (N_10117,N_9544,N_9831);
xor U10118 (N_10118,N_9125,N_9127);
or U10119 (N_10119,N_9523,N_9689);
nand U10120 (N_10120,N_9166,N_9202);
xnor U10121 (N_10121,N_9505,N_9525);
xor U10122 (N_10122,N_9444,N_9698);
nor U10123 (N_10123,N_9325,N_9997);
nand U10124 (N_10124,N_9278,N_9292);
and U10125 (N_10125,N_9309,N_9738);
and U10126 (N_10126,N_9156,N_9557);
xnor U10127 (N_10127,N_9387,N_9347);
or U10128 (N_10128,N_9632,N_9697);
nand U10129 (N_10129,N_9149,N_9153);
nor U10130 (N_10130,N_9530,N_9598);
or U10131 (N_10131,N_9287,N_9089);
xor U10132 (N_10132,N_9460,N_9974);
nand U10133 (N_10133,N_9160,N_9771);
xnor U10134 (N_10134,N_9956,N_9617);
nand U10135 (N_10135,N_9196,N_9577);
nand U10136 (N_10136,N_9553,N_9828);
and U10137 (N_10137,N_9701,N_9925);
xor U10138 (N_10138,N_9865,N_9662);
and U10139 (N_10139,N_9298,N_9639);
nor U10140 (N_10140,N_9704,N_9905);
nor U10141 (N_10141,N_9654,N_9461);
or U10142 (N_10142,N_9718,N_9853);
nor U10143 (N_10143,N_9864,N_9762);
nand U10144 (N_10144,N_9020,N_9514);
xor U10145 (N_10145,N_9422,N_9322);
and U10146 (N_10146,N_9735,N_9083);
and U10147 (N_10147,N_9794,N_9596);
xnor U10148 (N_10148,N_9755,N_9818);
nor U10149 (N_10149,N_9611,N_9122);
or U10150 (N_10150,N_9478,N_9277);
nand U10151 (N_10151,N_9213,N_9562);
nand U10152 (N_10152,N_9220,N_9655);
and U10153 (N_10153,N_9367,N_9090);
nand U10154 (N_10154,N_9578,N_9147);
and U10155 (N_10155,N_9979,N_9184);
nand U10156 (N_10156,N_9049,N_9206);
nor U10157 (N_10157,N_9843,N_9146);
and U10158 (N_10158,N_9102,N_9438);
xor U10159 (N_10159,N_9189,N_9039);
nand U10160 (N_10160,N_9243,N_9908);
nand U10161 (N_10161,N_9804,N_9085);
xnor U10162 (N_10162,N_9878,N_9044);
and U10163 (N_10163,N_9265,N_9264);
xnor U10164 (N_10164,N_9955,N_9313);
nor U10165 (N_10165,N_9229,N_9837);
and U10166 (N_10166,N_9939,N_9637);
xor U10167 (N_10167,N_9087,N_9914);
xnor U10168 (N_10168,N_9002,N_9235);
xnor U10169 (N_10169,N_9331,N_9685);
xnor U10170 (N_10170,N_9648,N_9671);
or U10171 (N_10171,N_9407,N_9032);
or U10172 (N_10172,N_9686,N_9402);
nor U10173 (N_10173,N_9494,N_9741);
nor U10174 (N_10174,N_9188,N_9063);
nand U10175 (N_10175,N_9279,N_9887);
nand U10176 (N_10176,N_9668,N_9801);
nand U10177 (N_10177,N_9403,N_9883);
nor U10178 (N_10178,N_9437,N_9948);
and U10179 (N_10179,N_9531,N_9694);
xor U10180 (N_10180,N_9778,N_9396);
and U10181 (N_10181,N_9921,N_9008);
and U10182 (N_10182,N_9116,N_9051);
or U10183 (N_10183,N_9895,N_9711);
nand U10184 (N_10184,N_9885,N_9053);
or U10185 (N_10185,N_9758,N_9472);
and U10186 (N_10186,N_9185,N_9432);
and U10187 (N_10187,N_9809,N_9554);
nor U10188 (N_10188,N_9256,N_9120);
xor U10189 (N_10189,N_9259,N_9501);
nand U10190 (N_10190,N_9015,N_9835);
or U10191 (N_10191,N_9645,N_9785);
and U10192 (N_10192,N_9647,N_9733);
nor U10193 (N_10193,N_9713,N_9245);
or U10194 (N_10194,N_9201,N_9286);
or U10195 (N_10195,N_9075,N_9172);
or U10196 (N_10196,N_9746,N_9095);
and U10197 (N_10197,N_9163,N_9565);
or U10198 (N_10198,N_9638,N_9931);
nor U10199 (N_10199,N_9533,N_9276);
nand U10200 (N_10200,N_9234,N_9110);
and U10201 (N_10201,N_9896,N_9115);
nor U10202 (N_10202,N_9070,N_9138);
nand U10203 (N_10203,N_9673,N_9517);
nand U10204 (N_10204,N_9364,N_9993);
nor U10205 (N_10205,N_9708,N_9369);
xnor U10206 (N_10206,N_9548,N_9359);
and U10207 (N_10207,N_9124,N_9690);
nand U10208 (N_10208,N_9246,N_9469);
nor U10209 (N_10209,N_9567,N_9376);
and U10210 (N_10210,N_9230,N_9927);
and U10211 (N_10211,N_9888,N_9010);
or U10212 (N_10212,N_9912,N_9255);
or U10213 (N_10213,N_9145,N_9688);
or U10214 (N_10214,N_9093,N_9603);
or U10215 (N_10215,N_9606,N_9487);
or U10216 (N_10216,N_9214,N_9710);
and U10217 (N_10217,N_9178,N_9663);
xnor U10218 (N_10218,N_9197,N_9707);
and U10219 (N_10219,N_9748,N_9495);
or U10220 (N_10220,N_9290,N_9107);
xor U10221 (N_10221,N_9340,N_9604);
or U10222 (N_10222,N_9537,N_9408);
nor U10223 (N_10223,N_9420,N_9210);
nor U10224 (N_10224,N_9826,N_9417);
nor U10225 (N_10225,N_9845,N_9275);
xor U10226 (N_10226,N_9579,N_9608);
nand U10227 (N_10227,N_9959,N_9154);
nand U10228 (N_10228,N_9303,N_9052);
nor U10229 (N_10229,N_9117,N_9782);
and U10230 (N_10230,N_9076,N_9267);
and U10231 (N_10231,N_9114,N_9846);
and U10232 (N_10232,N_9280,N_9635);
nor U10233 (N_10233,N_9547,N_9360);
nand U10234 (N_10234,N_9394,N_9913);
xnor U10235 (N_10235,N_9739,N_9729);
and U10236 (N_10236,N_9569,N_9209);
and U10237 (N_10237,N_9696,N_9048);
nand U10238 (N_10238,N_9191,N_9239);
xnor U10239 (N_10239,N_9806,N_9861);
nor U10240 (N_10240,N_9119,N_9958);
xnor U10241 (N_10241,N_9937,N_9082);
xor U10242 (N_10242,N_9848,N_9870);
xor U10243 (N_10243,N_9236,N_9502);
nand U10244 (N_10244,N_9378,N_9823);
xnor U10245 (N_10245,N_9538,N_9199);
and U10246 (N_10246,N_9642,N_9084);
and U10247 (N_10247,N_9966,N_9321);
nand U10248 (N_10248,N_9510,N_9038);
nand U10249 (N_10249,N_9774,N_9808);
xnor U10250 (N_10250,N_9252,N_9754);
or U10251 (N_10251,N_9193,N_9319);
xor U10252 (N_10252,N_9333,N_9574);
nand U10253 (N_10253,N_9410,N_9643);
or U10254 (N_10254,N_9855,N_9398);
xor U10255 (N_10255,N_9057,N_9678);
and U10256 (N_10256,N_9283,N_9174);
nor U10257 (N_10257,N_9854,N_9106);
nand U10258 (N_10258,N_9307,N_9842);
and U10259 (N_10259,N_9788,N_9140);
or U10260 (N_10260,N_9605,N_9851);
or U10261 (N_10261,N_9059,N_9929);
nor U10262 (N_10262,N_9088,N_9656);
nor U10263 (N_10263,N_9358,N_9204);
nor U10264 (N_10264,N_9098,N_9777);
and U10265 (N_10265,N_9282,N_9379);
or U10266 (N_10266,N_9418,N_9056);
xor U10267 (N_10267,N_9674,N_9653);
xnor U10268 (N_10268,N_9744,N_9260);
nand U10269 (N_10269,N_9249,N_9263);
xor U10270 (N_10270,N_9262,N_9977);
nand U10271 (N_10271,N_9316,N_9873);
nand U10272 (N_10272,N_9042,N_9136);
or U10273 (N_10273,N_9254,N_9257);
nor U10274 (N_10274,N_9772,N_9176);
nand U10275 (N_10275,N_9414,N_9101);
or U10276 (N_10276,N_9198,N_9304);
and U10277 (N_10277,N_9840,N_9511);
xnor U10278 (N_10278,N_9486,N_9657);
nor U10279 (N_10279,N_9750,N_9930);
or U10280 (N_10280,N_9872,N_9503);
nand U10281 (N_10281,N_9442,N_9456);
nor U10282 (N_10282,N_9421,N_9874);
xnor U10283 (N_10283,N_9406,N_9550);
xor U10284 (N_10284,N_9968,N_9649);
nand U10285 (N_10285,N_9081,N_9667);
nor U10286 (N_10286,N_9613,N_9768);
nand U10287 (N_10287,N_9344,N_9602);
nand U10288 (N_10288,N_9231,N_9683);
and U10289 (N_10289,N_9395,N_9516);
or U10290 (N_10290,N_9167,N_9731);
or U10291 (N_10291,N_9397,N_9411);
nor U10292 (N_10292,N_9227,N_9123);
nor U10293 (N_10293,N_9426,N_9863);
xnor U10294 (N_10294,N_9464,N_9474);
or U10295 (N_10295,N_9366,N_9192);
nand U10296 (N_10296,N_9473,N_9471);
and U10297 (N_10297,N_9624,N_9628);
or U10298 (N_10298,N_9769,N_9781);
xnor U10299 (N_10299,N_9354,N_9248);
or U10300 (N_10300,N_9518,N_9428);
nand U10301 (N_10301,N_9832,N_9796);
or U10302 (N_10302,N_9775,N_9522);
nor U10303 (N_10303,N_9291,N_9999);
nand U10304 (N_10304,N_9423,N_9933);
or U10305 (N_10305,N_9595,N_9222);
nor U10306 (N_10306,N_9712,N_9162);
or U10307 (N_10307,N_9824,N_9951);
xor U10308 (N_10308,N_9005,N_9009);
nand U10309 (N_10309,N_9892,N_9126);
or U10310 (N_10310,N_9142,N_9926);
and U10311 (N_10311,N_9969,N_9659);
xor U10312 (N_10312,N_9986,N_9205);
or U10313 (N_10313,N_9232,N_9786);
or U10314 (N_10314,N_9458,N_9441);
and U10315 (N_10315,N_9727,N_9695);
xnor U10316 (N_10316,N_9719,N_9982);
or U10317 (N_10317,N_9105,N_9024);
and U10318 (N_10318,N_9886,N_9535);
or U10319 (N_10319,N_9670,N_9992);
nand U10320 (N_10320,N_9022,N_9375);
xor U10321 (N_10321,N_9011,N_9593);
nand U10322 (N_10322,N_9725,N_9543);
and U10323 (N_10323,N_9625,N_9652);
xnor U10324 (N_10324,N_9377,N_9545);
or U10325 (N_10325,N_9390,N_9200);
nor U10326 (N_10326,N_9295,N_9803);
nor U10327 (N_10327,N_9268,N_9219);
xor U10328 (N_10328,N_9175,N_9452);
xor U10329 (N_10329,N_9092,N_9839);
nand U10330 (N_10330,N_9274,N_9618);
and U10331 (N_10331,N_9962,N_9620);
nor U10332 (N_10332,N_9067,N_9324);
xor U10333 (N_10333,N_9273,N_9270);
nand U10334 (N_10334,N_9534,N_9113);
and U10335 (N_10335,N_9330,N_9299);
or U10336 (N_10336,N_9296,N_9866);
nand U10337 (N_10337,N_9449,N_9759);
and U10338 (N_10338,N_9491,N_9869);
and U10339 (N_10339,N_9747,N_9342);
and U10340 (N_10340,N_9301,N_9879);
nor U10341 (N_10341,N_9017,N_9680);
nor U10342 (N_10342,N_9633,N_9644);
nand U10343 (N_10343,N_9346,N_9798);
and U10344 (N_10344,N_9207,N_9372);
or U10345 (N_10345,N_9001,N_9250);
xor U10346 (N_10346,N_9880,N_9155);
nor U10347 (N_10347,N_9302,N_9987);
xnor U10348 (N_10348,N_9217,N_9665);
nand U10349 (N_10349,N_9294,N_9190);
or U10350 (N_10350,N_9284,N_9766);
or U10351 (N_10351,N_9476,N_9447);
xor U10352 (N_10352,N_9454,N_9208);
xnor U10353 (N_10353,N_9742,N_9151);
nor U10354 (N_10354,N_9349,N_9182);
and U10355 (N_10355,N_9004,N_9756);
or U10356 (N_10356,N_9590,N_9271);
xor U10357 (N_10357,N_9722,N_9170);
or U10358 (N_10358,N_9584,N_9910);
nand U10359 (N_10359,N_9357,N_9244);
nand U10360 (N_10360,N_9792,N_9561);
nor U10361 (N_10361,N_9805,N_9749);
and U10362 (N_10362,N_9327,N_9492);
nor U10363 (N_10363,N_9508,N_9984);
nor U10364 (N_10364,N_9730,N_9978);
nand U10365 (N_10365,N_9062,N_9046);
xnor U10366 (N_10366,N_9773,N_9524);
xnor U10367 (N_10367,N_9890,N_9991);
nor U10368 (N_10368,N_9753,N_9027);
xor U10369 (N_10369,N_9388,N_9221);
nor U10370 (N_10370,N_9159,N_9705);
nor U10371 (N_10371,N_9228,N_9315);
nor U10372 (N_10372,N_9055,N_9763);
nor U10373 (N_10373,N_9026,N_9677);
and U10374 (N_10374,N_9343,N_9907);
or U10375 (N_10375,N_9446,N_9507);
and U10376 (N_10376,N_9949,N_9336);
or U10377 (N_10377,N_9401,N_9218);
or U10378 (N_10378,N_9060,N_9630);
nand U10379 (N_10379,N_9356,N_9967);
nor U10380 (N_10380,N_9033,N_9841);
or U10381 (N_10381,N_9061,N_9699);
xnor U10382 (N_10382,N_9045,N_9073);
and U10383 (N_10383,N_9717,N_9591);
nor U10384 (N_10384,N_9852,N_9973);
nand U10385 (N_10385,N_9555,N_9233);
or U10386 (N_10386,N_9622,N_9069);
nand U10387 (N_10387,N_9821,N_9963);
or U10388 (N_10388,N_9499,N_9743);
and U10389 (N_10389,N_9877,N_9580);
or U10390 (N_10390,N_9370,N_9761);
nand U10391 (N_10391,N_9783,N_9607);
or U10392 (N_10392,N_9950,N_9640);
or U10393 (N_10393,N_9797,N_9751);
and U10394 (N_10394,N_9539,N_9827);
nor U10395 (N_10395,N_9582,N_9180);
and U10396 (N_10396,N_9692,N_9836);
xor U10397 (N_10397,N_9985,N_9568);
xor U10398 (N_10398,N_9957,N_9479);
or U10399 (N_10399,N_9148,N_9592);
and U10400 (N_10400,N_9970,N_9911);
or U10401 (N_10401,N_9400,N_9650);
nand U10402 (N_10402,N_9588,N_9627);
or U10403 (N_10403,N_9924,N_9308);
nor U10404 (N_10404,N_9980,N_9050);
or U10405 (N_10405,N_9152,N_9181);
nor U10406 (N_10406,N_9679,N_9312);
nand U10407 (N_10407,N_9601,N_9675);
xnor U10408 (N_10408,N_9318,N_9882);
xnor U10409 (N_10409,N_9068,N_9043);
nor U10410 (N_10410,N_9953,N_9563);
nand U10411 (N_10411,N_9462,N_9881);
or U10412 (N_10412,N_9500,N_9040);
nor U10413 (N_10413,N_9767,N_9133);
and U10414 (N_10414,N_9253,N_9013);
nand U10415 (N_10415,N_9700,N_9619);
or U10416 (N_10416,N_9512,N_9621);
nand U10417 (N_10417,N_9546,N_9337);
or U10418 (N_10418,N_9536,N_9096);
nor U10419 (N_10419,N_9998,N_9519);
nand U10420 (N_10420,N_9903,N_9371);
nand U10421 (N_10421,N_9720,N_9780);
nor U10422 (N_10422,N_9485,N_9904);
and U10423 (N_10423,N_9664,N_9317);
nand U10424 (N_10424,N_9112,N_9740);
and U10425 (N_10425,N_9183,N_9488);
and U10426 (N_10426,N_9889,N_9636);
nor U10427 (N_10427,N_9726,N_9572);
and U10428 (N_10428,N_9074,N_9141);
xnor U10429 (N_10429,N_9457,N_9079);
and U10430 (N_10430,N_9834,N_9480);
nor U10431 (N_10431,N_9434,N_9445);
nand U10432 (N_10432,N_9345,N_9856);
and U10433 (N_10433,N_9669,N_9224);
xnor U10434 (N_10434,N_9918,N_9078);
nand U10435 (N_10435,N_9226,N_9139);
nor U10436 (N_10436,N_9552,N_9427);
or U10437 (N_10437,N_9728,N_9560);
xor U10438 (N_10438,N_9587,N_9790);
xnor U10439 (N_10439,N_9682,N_9351);
nand U10440 (N_10440,N_9334,N_9496);
xnor U10441 (N_10441,N_9157,N_9594);
xnor U10442 (N_10442,N_9528,N_9094);
xor U10443 (N_10443,N_9813,N_9811);
xnor U10444 (N_10444,N_9025,N_9240);
and U10445 (N_10445,N_9416,N_9849);
nor U10446 (N_10446,N_9430,N_9526);
xnor U10447 (N_10447,N_9440,N_9954);
or U10448 (N_10448,N_9916,N_9513);
and U10449 (N_10449,N_9898,N_9323);
xor U10450 (N_10450,N_9944,N_9288);
nor U10451 (N_10451,N_9179,N_9612);
xor U10452 (N_10452,N_9850,N_9150);
and U10453 (N_10453,N_9064,N_9289);
nand U10454 (N_10454,N_9393,N_9493);
nor U10455 (N_10455,N_9702,N_9459);
or U10456 (N_10456,N_9104,N_9389);
or U10457 (N_10457,N_9829,N_9615);
xor U10458 (N_10458,N_9564,N_9435);
nor U10459 (N_10459,N_9964,N_9599);
nand U10460 (N_10460,N_9723,N_9164);
and U10461 (N_10461,N_9103,N_9326);
and U10462 (N_10462,N_9072,N_9258);
nand U10463 (N_10463,N_9490,N_9940);
xor U10464 (N_10464,N_9532,N_9132);
or U10465 (N_10465,N_9972,N_9976);
or U10466 (N_10466,N_9100,N_9757);
and U10467 (N_10467,N_9947,N_9875);
or U10468 (N_10468,N_9981,N_9609);
nor U10469 (N_10469,N_9847,N_9293);
nand U10470 (N_10470,N_9269,N_9631);
or U10471 (N_10471,N_9529,N_9802);
nand U10472 (N_10472,N_9405,N_9041);
nand U10473 (N_10473,N_9816,N_9384);
nand U10474 (N_10474,N_9031,N_9483);
nand U10475 (N_10475,N_9551,N_9891);
nor U10476 (N_10476,N_9381,N_9812);
and U10477 (N_10477,N_9506,N_9996);
or U10478 (N_10478,N_9203,N_9884);
nor U10479 (N_10479,N_9721,N_9242);
and U10480 (N_10480,N_9573,N_9328);
xor U10481 (N_10481,N_9353,N_9830);
and U10482 (N_10482,N_9237,N_9902);
and U10483 (N_10483,N_9658,N_9266);
xnor U10484 (N_10484,N_9036,N_9570);
or U10485 (N_10485,N_9003,N_9341);
nand U10486 (N_10486,N_9365,N_9687);
nor U10487 (N_10487,N_9482,N_9409);
or U10488 (N_10488,N_9021,N_9131);
or U10489 (N_10489,N_9158,N_9935);
nor U10490 (N_10490,N_9857,N_9362);
or U10491 (N_10491,N_9433,N_9597);
and U10492 (N_10492,N_9906,N_9436);
nand U10493 (N_10493,N_9134,N_9583);
nor U10494 (N_10494,N_9825,N_9453);
and U10495 (N_10495,N_9465,N_9923);
nand U10496 (N_10496,N_9932,N_9791);
and U10497 (N_10497,N_9504,N_9586);
xnor U10498 (N_10498,N_9225,N_9575);
xor U10499 (N_10499,N_9559,N_9521);
nand U10500 (N_10500,N_9302,N_9608);
nand U10501 (N_10501,N_9451,N_9759);
and U10502 (N_10502,N_9010,N_9358);
nand U10503 (N_10503,N_9023,N_9526);
xnor U10504 (N_10504,N_9319,N_9613);
and U10505 (N_10505,N_9650,N_9421);
or U10506 (N_10506,N_9726,N_9779);
nor U10507 (N_10507,N_9673,N_9954);
nand U10508 (N_10508,N_9914,N_9729);
or U10509 (N_10509,N_9064,N_9943);
and U10510 (N_10510,N_9493,N_9378);
and U10511 (N_10511,N_9418,N_9069);
or U10512 (N_10512,N_9206,N_9851);
and U10513 (N_10513,N_9216,N_9412);
xor U10514 (N_10514,N_9480,N_9599);
and U10515 (N_10515,N_9777,N_9564);
nand U10516 (N_10516,N_9533,N_9958);
and U10517 (N_10517,N_9586,N_9696);
nor U10518 (N_10518,N_9690,N_9409);
or U10519 (N_10519,N_9409,N_9360);
and U10520 (N_10520,N_9154,N_9799);
and U10521 (N_10521,N_9699,N_9996);
or U10522 (N_10522,N_9472,N_9889);
and U10523 (N_10523,N_9553,N_9857);
nand U10524 (N_10524,N_9078,N_9034);
nand U10525 (N_10525,N_9503,N_9918);
nor U10526 (N_10526,N_9289,N_9759);
nor U10527 (N_10527,N_9158,N_9329);
nand U10528 (N_10528,N_9461,N_9012);
nor U10529 (N_10529,N_9506,N_9345);
and U10530 (N_10530,N_9858,N_9890);
nor U10531 (N_10531,N_9830,N_9963);
nor U10532 (N_10532,N_9124,N_9254);
nor U10533 (N_10533,N_9186,N_9442);
xor U10534 (N_10534,N_9092,N_9983);
and U10535 (N_10535,N_9054,N_9058);
and U10536 (N_10536,N_9950,N_9537);
xor U10537 (N_10537,N_9325,N_9580);
xor U10538 (N_10538,N_9952,N_9597);
or U10539 (N_10539,N_9877,N_9581);
nand U10540 (N_10540,N_9187,N_9163);
nor U10541 (N_10541,N_9923,N_9016);
nand U10542 (N_10542,N_9199,N_9772);
xnor U10543 (N_10543,N_9793,N_9358);
and U10544 (N_10544,N_9598,N_9439);
or U10545 (N_10545,N_9089,N_9876);
nor U10546 (N_10546,N_9112,N_9299);
nor U10547 (N_10547,N_9121,N_9871);
nor U10548 (N_10548,N_9833,N_9586);
and U10549 (N_10549,N_9084,N_9413);
and U10550 (N_10550,N_9853,N_9709);
xor U10551 (N_10551,N_9542,N_9154);
and U10552 (N_10552,N_9786,N_9528);
nand U10553 (N_10553,N_9241,N_9857);
nand U10554 (N_10554,N_9924,N_9541);
or U10555 (N_10555,N_9472,N_9237);
nor U10556 (N_10556,N_9986,N_9735);
or U10557 (N_10557,N_9328,N_9226);
or U10558 (N_10558,N_9517,N_9946);
or U10559 (N_10559,N_9470,N_9733);
or U10560 (N_10560,N_9056,N_9557);
nand U10561 (N_10561,N_9676,N_9106);
xnor U10562 (N_10562,N_9879,N_9426);
xor U10563 (N_10563,N_9537,N_9066);
nor U10564 (N_10564,N_9047,N_9666);
xnor U10565 (N_10565,N_9159,N_9752);
xor U10566 (N_10566,N_9432,N_9696);
nor U10567 (N_10567,N_9127,N_9722);
nor U10568 (N_10568,N_9338,N_9836);
and U10569 (N_10569,N_9368,N_9369);
xor U10570 (N_10570,N_9755,N_9804);
or U10571 (N_10571,N_9632,N_9881);
and U10572 (N_10572,N_9787,N_9074);
xor U10573 (N_10573,N_9103,N_9398);
xor U10574 (N_10574,N_9987,N_9231);
xnor U10575 (N_10575,N_9308,N_9217);
nand U10576 (N_10576,N_9628,N_9636);
nor U10577 (N_10577,N_9905,N_9097);
and U10578 (N_10578,N_9532,N_9423);
and U10579 (N_10579,N_9896,N_9831);
nor U10580 (N_10580,N_9948,N_9904);
xor U10581 (N_10581,N_9680,N_9625);
xor U10582 (N_10582,N_9451,N_9096);
or U10583 (N_10583,N_9339,N_9398);
or U10584 (N_10584,N_9106,N_9218);
or U10585 (N_10585,N_9243,N_9060);
nor U10586 (N_10586,N_9606,N_9308);
and U10587 (N_10587,N_9324,N_9035);
and U10588 (N_10588,N_9393,N_9929);
nor U10589 (N_10589,N_9129,N_9823);
and U10590 (N_10590,N_9518,N_9101);
or U10591 (N_10591,N_9738,N_9477);
xor U10592 (N_10592,N_9238,N_9108);
xnor U10593 (N_10593,N_9976,N_9595);
xnor U10594 (N_10594,N_9747,N_9357);
xnor U10595 (N_10595,N_9725,N_9573);
and U10596 (N_10596,N_9235,N_9612);
and U10597 (N_10597,N_9567,N_9087);
and U10598 (N_10598,N_9647,N_9722);
xor U10599 (N_10599,N_9132,N_9963);
nor U10600 (N_10600,N_9876,N_9193);
and U10601 (N_10601,N_9673,N_9631);
nor U10602 (N_10602,N_9117,N_9823);
xor U10603 (N_10603,N_9998,N_9749);
nor U10604 (N_10604,N_9875,N_9845);
and U10605 (N_10605,N_9869,N_9552);
or U10606 (N_10606,N_9156,N_9359);
and U10607 (N_10607,N_9915,N_9966);
and U10608 (N_10608,N_9744,N_9342);
xnor U10609 (N_10609,N_9284,N_9959);
nor U10610 (N_10610,N_9334,N_9892);
and U10611 (N_10611,N_9970,N_9626);
nor U10612 (N_10612,N_9253,N_9255);
and U10613 (N_10613,N_9284,N_9299);
and U10614 (N_10614,N_9159,N_9630);
nor U10615 (N_10615,N_9893,N_9940);
nor U10616 (N_10616,N_9769,N_9768);
nor U10617 (N_10617,N_9887,N_9002);
nand U10618 (N_10618,N_9989,N_9937);
xor U10619 (N_10619,N_9550,N_9441);
nor U10620 (N_10620,N_9535,N_9336);
nor U10621 (N_10621,N_9912,N_9150);
or U10622 (N_10622,N_9073,N_9732);
or U10623 (N_10623,N_9739,N_9342);
xnor U10624 (N_10624,N_9717,N_9752);
xor U10625 (N_10625,N_9315,N_9470);
or U10626 (N_10626,N_9027,N_9469);
nor U10627 (N_10627,N_9583,N_9863);
nor U10628 (N_10628,N_9697,N_9669);
nand U10629 (N_10629,N_9787,N_9444);
nand U10630 (N_10630,N_9908,N_9840);
xor U10631 (N_10631,N_9223,N_9584);
xnor U10632 (N_10632,N_9595,N_9081);
nor U10633 (N_10633,N_9271,N_9046);
or U10634 (N_10634,N_9011,N_9991);
or U10635 (N_10635,N_9104,N_9658);
and U10636 (N_10636,N_9326,N_9504);
nor U10637 (N_10637,N_9422,N_9958);
and U10638 (N_10638,N_9396,N_9100);
nor U10639 (N_10639,N_9800,N_9879);
and U10640 (N_10640,N_9360,N_9795);
or U10641 (N_10641,N_9355,N_9587);
and U10642 (N_10642,N_9045,N_9047);
or U10643 (N_10643,N_9061,N_9882);
or U10644 (N_10644,N_9720,N_9986);
or U10645 (N_10645,N_9061,N_9425);
nor U10646 (N_10646,N_9009,N_9364);
nor U10647 (N_10647,N_9299,N_9373);
xnor U10648 (N_10648,N_9777,N_9581);
nand U10649 (N_10649,N_9524,N_9724);
xnor U10650 (N_10650,N_9691,N_9539);
and U10651 (N_10651,N_9176,N_9749);
and U10652 (N_10652,N_9593,N_9573);
xor U10653 (N_10653,N_9832,N_9586);
or U10654 (N_10654,N_9039,N_9922);
or U10655 (N_10655,N_9006,N_9337);
nand U10656 (N_10656,N_9310,N_9512);
nor U10657 (N_10657,N_9842,N_9237);
or U10658 (N_10658,N_9961,N_9451);
xnor U10659 (N_10659,N_9625,N_9818);
or U10660 (N_10660,N_9969,N_9648);
nand U10661 (N_10661,N_9382,N_9723);
nor U10662 (N_10662,N_9919,N_9024);
nor U10663 (N_10663,N_9990,N_9969);
and U10664 (N_10664,N_9125,N_9651);
nand U10665 (N_10665,N_9279,N_9185);
or U10666 (N_10666,N_9212,N_9182);
xnor U10667 (N_10667,N_9476,N_9882);
or U10668 (N_10668,N_9113,N_9544);
xnor U10669 (N_10669,N_9098,N_9248);
and U10670 (N_10670,N_9067,N_9015);
xnor U10671 (N_10671,N_9766,N_9654);
nand U10672 (N_10672,N_9857,N_9560);
or U10673 (N_10673,N_9041,N_9878);
nor U10674 (N_10674,N_9177,N_9397);
xnor U10675 (N_10675,N_9591,N_9734);
nor U10676 (N_10676,N_9527,N_9807);
xor U10677 (N_10677,N_9384,N_9300);
or U10678 (N_10678,N_9066,N_9713);
xor U10679 (N_10679,N_9865,N_9941);
nand U10680 (N_10680,N_9044,N_9948);
xnor U10681 (N_10681,N_9568,N_9484);
nand U10682 (N_10682,N_9040,N_9790);
or U10683 (N_10683,N_9303,N_9919);
xnor U10684 (N_10684,N_9790,N_9608);
nor U10685 (N_10685,N_9392,N_9080);
or U10686 (N_10686,N_9250,N_9025);
nand U10687 (N_10687,N_9764,N_9663);
nor U10688 (N_10688,N_9699,N_9286);
xnor U10689 (N_10689,N_9865,N_9272);
or U10690 (N_10690,N_9230,N_9054);
nor U10691 (N_10691,N_9538,N_9561);
and U10692 (N_10692,N_9451,N_9783);
xnor U10693 (N_10693,N_9183,N_9072);
nor U10694 (N_10694,N_9432,N_9069);
or U10695 (N_10695,N_9495,N_9326);
or U10696 (N_10696,N_9786,N_9998);
nand U10697 (N_10697,N_9362,N_9973);
nor U10698 (N_10698,N_9487,N_9899);
and U10699 (N_10699,N_9500,N_9013);
nor U10700 (N_10700,N_9817,N_9276);
and U10701 (N_10701,N_9112,N_9536);
and U10702 (N_10702,N_9176,N_9115);
xor U10703 (N_10703,N_9497,N_9087);
or U10704 (N_10704,N_9747,N_9116);
nor U10705 (N_10705,N_9062,N_9281);
nand U10706 (N_10706,N_9424,N_9837);
and U10707 (N_10707,N_9107,N_9144);
or U10708 (N_10708,N_9565,N_9938);
xor U10709 (N_10709,N_9376,N_9276);
nand U10710 (N_10710,N_9189,N_9097);
xnor U10711 (N_10711,N_9474,N_9414);
and U10712 (N_10712,N_9627,N_9563);
nor U10713 (N_10713,N_9050,N_9583);
xor U10714 (N_10714,N_9690,N_9761);
nand U10715 (N_10715,N_9088,N_9925);
and U10716 (N_10716,N_9594,N_9227);
or U10717 (N_10717,N_9476,N_9054);
nand U10718 (N_10718,N_9962,N_9395);
or U10719 (N_10719,N_9583,N_9920);
nand U10720 (N_10720,N_9893,N_9253);
and U10721 (N_10721,N_9337,N_9393);
nand U10722 (N_10722,N_9855,N_9448);
nor U10723 (N_10723,N_9553,N_9616);
xor U10724 (N_10724,N_9336,N_9530);
xnor U10725 (N_10725,N_9328,N_9161);
nand U10726 (N_10726,N_9061,N_9439);
or U10727 (N_10727,N_9255,N_9732);
or U10728 (N_10728,N_9254,N_9604);
nor U10729 (N_10729,N_9979,N_9560);
xor U10730 (N_10730,N_9870,N_9525);
nor U10731 (N_10731,N_9115,N_9752);
nand U10732 (N_10732,N_9361,N_9633);
nor U10733 (N_10733,N_9178,N_9351);
xnor U10734 (N_10734,N_9897,N_9116);
or U10735 (N_10735,N_9920,N_9919);
nor U10736 (N_10736,N_9503,N_9093);
or U10737 (N_10737,N_9528,N_9690);
nand U10738 (N_10738,N_9605,N_9020);
nand U10739 (N_10739,N_9371,N_9567);
and U10740 (N_10740,N_9714,N_9679);
or U10741 (N_10741,N_9535,N_9840);
or U10742 (N_10742,N_9010,N_9932);
and U10743 (N_10743,N_9101,N_9265);
nand U10744 (N_10744,N_9140,N_9873);
nor U10745 (N_10745,N_9032,N_9992);
nand U10746 (N_10746,N_9946,N_9675);
and U10747 (N_10747,N_9703,N_9908);
and U10748 (N_10748,N_9361,N_9764);
xor U10749 (N_10749,N_9230,N_9188);
nand U10750 (N_10750,N_9064,N_9481);
and U10751 (N_10751,N_9307,N_9261);
and U10752 (N_10752,N_9859,N_9833);
or U10753 (N_10753,N_9846,N_9175);
and U10754 (N_10754,N_9428,N_9292);
nand U10755 (N_10755,N_9052,N_9030);
nand U10756 (N_10756,N_9840,N_9752);
or U10757 (N_10757,N_9515,N_9030);
xor U10758 (N_10758,N_9264,N_9622);
nand U10759 (N_10759,N_9796,N_9477);
nor U10760 (N_10760,N_9033,N_9301);
xnor U10761 (N_10761,N_9786,N_9041);
or U10762 (N_10762,N_9883,N_9626);
or U10763 (N_10763,N_9123,N_9028);
nor U10764 (N_10764,N_9391,N_9383);
xnor U10765 (N_10765,N_9047,N_9322);
nor U10766 (N_10766,N_9916,N_9546);
and U10767 (N_10767,N_9388,N_9410);
nor U10768 (N_10768,N_9887,N_9119);
and U10769 (N_10769,N_9333,N_9356);
or U10770 (N_10770,N_9961,N_9719);
or U10771 (N_10771,N_9241,N_9538);
nand U10772 (N_10772,N_9868,N_9745);
xor U10773 (N_10773,N_9261,N_9538);
nor U10774 (N_10774,N_9392,N_9508);
xnor U10775 (N_10775,N_9368,N_9306);
nor U10776 (N_10776,N_9095,N_9422);
nor U10777 (N_10777,N_9365,N_9419);
xor U10778 (N_10778,N_9896,N_9394);
xor U10779 (N_10779,N_9695,N_9556);
xor U10780 (N_10780,N_9567,N_9979);
nand U10781 (N_10781,N_9073,N_9661);
xnor U10782 (N_10782,N_9720,N_9519);
and U10783 (N_10783,N_9936,N_9270);
or U10784 (N_10784,N_9245,N_9357);
and U10785 (N_10785,N_9314,N_9096);
nor U10786 (N_10786,N_9904,N_9828);
and U10787 (N_10787,N_9017,N_9320);
xnor U10788 (N_10788,N_9040,N_9485);
nand U10789 (N_10789,N_9990,N_9502);
nor U10790 (N_10790,N_9275,N_9334);
nor U10791 (N_10791,N_9709,N_9010);
xnor U10792 (N_10792,N_9547,N_9076);
nand U10793 (N_10793,N_9931,N_9973);
xnor U10794 (N_10794,N_9866,N_9047);
nor U10795 (N_10795,N_9991,N_9607);
or U10796 (N_10796,N_9115,N_9384);
or U10797 (N_10797,N_9075,N_9321);
xor U10798 (N_10798,N_9366,N_9959);
nor U10799 (N_10799,N_9891,N_9532);
and U10800 (N_10800,N_9581,N_9486);
and U10801 (N_10801,N_9108,N_9878);
or U10802 (N_10802,N_9975,N_9088);
nor U10803 (N_10803,N_9770,N_9170);
nor U10804 (N_10804,N_9493,N_9325);
and U10805 (N_10805,N_9422,N_9591);
or U10806 (N_10806,N_9858,N_9224);
nand U10807 (N_10807,N_9368,N_9499);
and U10808 (N_10808,N_9467,N_9333);
or U10809 (N_10809,N_9913,N_9507);
or U10810 (N_10810,N_9672,N_9134);
nor U10811 (N_10811,N_9710,N_9090);
nand U10812 (N_10812,N_9510,N_9549);
and U10813 (N_10813,N_9713,N_9568);
or U10814 (N_10814,N_9063,N_9084);
and U10815 (N_10815,N_9318,N_9084);
and U10816 (N_10816,N_9380,N_9239);
nand U10817 (N_10817,N_9473,N_9625);
or U10818 (N_10818,N_9599,N_9901);
nor U10819 (N_10819,N_9302,N_9847);
or U10820 (N_10820,N_9268,N_9201);
xor U10821 (N_10821,N_9725,N_9759);
xor U10822 (N_10822,N_9992,N_9892);
nor U10823 (N_10823,N_9604,N_9608);
and U10824 (N_10824,N_9090,N_9785);
xor U10825 (N_10825,N_9111,N_9983);
and U10826 (N_10826,N_9611,N_9697);
xor U10827 (N_10827,N_9154,N_9296);
and U10828 (N_10828,N_9694,N_9526);
xor U10829 (N_10829,N_9578,N_9195);
nand U10830 (N_10830,N_9658,N_9892);
or U10831 (N_10831,N_9667,N_9828);
and U10832 (N_10832,N_9914,N_9368);
or U10833 (N_10833,N_9037,N_9684);
and U10834 (N_10834,N_9340,N_9625);
and U10835 (N_10835,N_9564,N_9380);
nand U10836 (N_10836,N_9132,N_9177);
nand U10837 (N_10837,N_9598,N_9305);
nor U10838 (N_10838,N_9496,N_9557);
xnor U10839 (N_10839,N_9738,N_9677);
xnor U10840 (N_10840,N_9281,N_9306);
or U10841 (N_10841,N_9626,N_9322);
nand U10842 (N_10842,N_9697,N_9152);
or U10843 (N_10843,N_9690,N_9423);
nand U10844 (N_10844,N_9506,N_9720);
nand U10845 (N_10845,N_9857,N_9675);
xnor U10846 (N_10846,N_9934,N_9790);
nand U10847 (N_10847,N_9288,N_9620);
xnor U10848 (N_10848,N_9267,N_9581);
and U10849 (N_10849,N_9541,N_9721);
or U10850 (N_10850,N_9656,N_9000);
and U10851 (N_10851,N_9548,N_9222);
or U10852 (N_10852,N_9957,N_9435);
or U10853 (N_10853,N_9608,N_9492);
and U10854 (N_10854,N_9827,N_9221);
nor U10855 (N_10855,N_9641,N_9624);
and U10856 (N_10856,N_9980,N_9637);
or U10857 (N_10857,N_9237,N_9277);
or U10858 (N_10858,N_9593,N_9719);
xnor U10859 (N_10859,N_9958,N_9942);
xor U10860 (N_10860,N_9009,N_9635);
nand U10861 (N_10861,N_9319,N_9309);
xnor U10862 (N_10862,N_9313,N_9500);
nand U10863 (N_10863,N_9608,N_9523);
and U10864 (N_10864,N_9731,N_9842);
xor U10865 (N_10865,N_9977,N_9641);
nand U10866 (N_10866,N_9726,N_9752);
xnor U10867 (N_10867,N_9196,N_9134);
and U10868 (N_10868,N_9155,N_9239);
xnor U10869 (N_10869,N_9187,N_9773);
nor U10870 (N_10870,N_9171,N_9820);
nand U10871 (N_10871,N_9805,N_9566);
or U10872 (N_10872,N_9575,N_9690);
nor U10873 (N_10873,N_9591,N_9225);
and U10874 (N_10874,N_9054,N_9150);
or U10875 (N_10875,N_9497,N_9653);
nand U10876 (N_10876,N_9338,N_9916);
xor U10877 (N_10877,N_9880,N_9680);
or U10878 (N_10878,N_9388,N_9153);
nand U10879 (N_10879,N_9056,N_9215);
xor U10880 (N_10880,N_9804,N_9921);
xnor U10881 (N_10881,N_9844,N_9027);
nor U10882 (N_10882,N_9478,N_9519);
and U10883 (N_10883,N_9071,N_9564);
xor U10884 (N_10884,N_9775,N_9860);
nor U10885 (N_10885,N_9398,N_9919);
xnor U10886 (N_10886,N_9203,N_9695);
or U10887 (N_10887,N_9077,N_9548);
nor U10888 (N_10888,N_9441,N_9509);
or U10889 (N_10889,N_9535,N_9110);
and U10890 (N_10890,N_9065,N_9892);
xor U10891 (N_10891,N_9777,N_9802);
or U10892 (N_10892,N_9544,N_9488);
or U10893 (N_10893,N_9616,N_9100);
xor U10894 (N_10894,N_9485,N_9463);
or U10895 (N_10895,N_9118,N_9497);
and U10896 (N_10896,N_9579,N_9265);
nand U10897 (N_10897,N_9114,N_9242);
nand U10898 (N_10898,N_9556,N_9568);
nor U10899 (N_10899,N_9314,N_9250);
nor U10900 (N_10900,N_9795,N_9654);
or U10901 (N_10901,N_9019,N_9486);
nor U10902 (N_10902,N_9315,N_9974);
or U10903 (N_10903,N_9502,N_9550);
or U10904 (N_10904,N_9061,N_9857);
nor U10905 (N_10905,N_9437,N_9069);
nand U10906 (N_10906,N_9975,N_9063);
nor U10907 (N_10907,N_9654,N_9250);
or U10908 (N_10908,N_9082,N_9696);
nor U10909 (N_10909,N_9972,N_9299);
and U10910 (N_10910,N_9917,N_9321);
xnor U10911 (N_10911,N_9283,N_9846);
nor U10912 (N_10912,N_9509,N_9623);
xor U10913 (N_10913,N_9079,N_9901);
and U10914 (N_10914,N_9360,N_9916);
nand U10915 (N_10915,N_9954,N_9796);
and U10916 (N_10916,N_9433,N_9011);
xnor U10917 (N_10917,N_9181,N_9661);
xor U10918 (N_10918,N_9741,N_9321);
or U10919 (N_10919,N_9357,N_9891);
and U10920 (N_10920,N_9717,N_9515);
and U10921 (N_10921,N_9182,N_9907);
and U10922 (N_10922,N_9023,N_9090);
or U10923 (N_10923,N_9562,N_9315);
or U10924 (N_10924,N_9980,N_9185);
nor U10925 (N_10925,N_9686,N_9212);
and U10926 (N_10926,N_9843,N_9134);
xnor U10927 (N_10927,N_9037,N_9288);
nand U10928 (N_10928,N_9781,N_9194);
and U10929 (N_10929,N_9707,N_9261);
or U10930 (N_10930,N_9586,N_9872);
xor U10931 (N_10931,N_9580,N_9781);
nand U10932 (N_10932,N_9101,N_9844);
nand U10933 (N_10933,N_9312,N_9038);
and U10934 (N_10934,N_9065,N_9593);
nand U10935 (N_10935,N_9473,N_9651);
or U10936 (N_10936,N_9575,N_9523);
xnor U10937 (N_10937,N_9732,N_9799);
and U10938 (N_10938,N_9829,N_9188);
nand U10939 (N_10939,N_9711,N_9902);
xnor U10940 (N_10940,N_9877,N_9469);
nand U10941 (N_10941,N_9545,N_9229);
nor U10942 (N_10942,N_9790,N_9275);
xor U10943 (N_10943,N_9899,N_9193);
or U10944 (N_10944,N_9614,N_9920);
nand U10945 (N_10945,N_9796,N_9585);
and U10946 (N_10946,N_9099,N_9927);
nand U10947 (N_10947,N_9897,N_9450);
xor U10948 (N_10948,N_9542,N_9452);
xor U10949 (N_10949,N_9378,N_9522);
nor U10950 (N_10950,N_9654,N_9175);
nand U10951 (N_10951,N_9232,N_9176);
xor U10952 (N_10952,N_9140,N_9105);
nor U10953 (N_10953,N_9659,N_9018);
and U10954 (N_10954,N_9668,N_9920);
nor U10955 (N_10955,N_9765,N_9185);
nor U10956 (N_10956,N_9256,N_9738);
nand U10957 (N_10957,N_9004,N_9097);
and U10958 (N_10958,N_9514,N_9340);
and U10959 (N_10959,N_9931,N_9927);
and U10960 (N_10960,N_9550,N_9586);
nor U10961 (N_10961,N_9688,N_9398);
nand U10962 (N_10962,N_9946,N_9673);
and U10963 (N_10963,N_9881,N_9519);
and U10964 (N_10964,N_9250,N_9565);
nand U10965 (N_10965,N_9401,N_9420);
nand U10966 (N_10966,N_9116,N_9704);
xnor U10967 (N_10967,N_9497,N_9015);
xnor U10968 (N_10968,N_9067,N_9431);
nand U10969 (N_10969,N_9867,N_9754);
nor U10970 (N_10970,N_9138,N_9836);
or U10971 (N_10971,N_9407,N_9759);
or U10972 (N_10972,N_9284,N_9532);
xor U10973 (N_10973,N_9612,N_9416);
and U10974 (N_10974,N_9319,N_9168);
xnor U10975 (N_10975,N_9379,N_9336);
xor U10976 (N_10976,N_9816,N_9890);
or U10977 (N_10977,N_9740,N_9634);
nand U10978 (N_10978,N_9273,N_9733);
nand U10979 (N_10979,N_9926,N_9247);
nor U10980 (N_10980,N_9543,N_9149);
or U10981 (N_10981,N_9751,N_9692);
or U10982 (N_10982,N_9682,N_9861);
nand U10983 (N_10983,N_9810,N_9943);
nor U10984 (N_10984,N_9077,N_9020);
nand U10985 (N_10985,N_9429,N_9330);
nor U10986 (N_10986,N_9980,N_9447);
and U10987 (N_10987,N_9056,N_9110);
nand U10988 (N_10988,N_9577,N_9874);
nor U10989 (N_10989,N_9116,N_9925);
or U10990 (N_10990,N_9597,N_9815);
and U10991 (N_10991,N_9877,N_9314);
and U10992 (N_10992,N_9129,N_9133);
and U10993 (N_10993,N_9929,N_9293);
or U10994 (N_10994,N_9072,N_9292);
nor U10995 (N_10995,N_9965,N_9250);
nand U10996 (N_10996,N_9883,N_9348);
or U10997 (N_10997,N_9494,N_9012);
nor U10998 (N_10998,N_9425,N_9510);
xnor U10999 (N_10999,N_9120,N_9887);
or U11000 (N_11000,N_10378,N_10542);
xnor U11001 (N_11001,N_10335,N_10725);
nand U11002 (N_11002,N_10122,N_10007);
or U11003 (N_11003,N_10191,N_10065);
or U11004 (N_11004,N_10402,N_10879);
and U11005 (N_11005,N_10983,N_10736);
nor U11006 (N_11006,N_10767,N_10946);
nor U11007 (N_11007,N_10538,N_10233);
and U11008 (N_11008,N_10118,N_10570);
xnor U11009 (N_11009,N_10059,N_10374);
and U11010 (N_11010,N_10091,N_10670);
nand U11011 (N_11011,N_10762,N_10565);
and U11012 (N_11012,N_10809,N_10087);
or U11013 (N_11013,N_10868,N_10174);
nand U11014 (N_11014,N_10349,N_10436);
xor U11015 (N_11015,N_10110,N_10265);
nand U11016 (N_11016,N_10236,N_10443);
and U11017 (N_11017,N_10874,N_10893);
xor U11018 (N_11018,N_10856,N_10627);
and U11019 (N_11019,N_10653,N_10389);
xnor U11020 (N_11020,N_10372,N_10268);
xor U11021 (N_11021,N_10970,N_10495);
or U11022 (N_11022,N_10786,N_10084);
nand U11023 (N_11023,N_10985,N_10644);
or U11024 (N_11024,N_10535,N_10224);
nand U11025 (N_11025,N_10253,N_10184);
nand U11026 (N_11026,N_10938,N_10036);
or U11027 (N_11027,N_10602,N_10482);
or U11028 (N_11028,N_10775,N_10485);
nor U11029 (N_11029,N_10547,N_10305);
nor U11030 (N_11030,N_10697,N_10537);
or U11031 (N_11031,N_10857,N_10380);
xor U11032 (N_11032,N_10309,N_10613);
nor U11033 (N_11033,N_10832,N_10971);
and U11034 (N_11034,N_10039,N_10450);
xnor U11035 (N_11035,N_10444,N_10416);
nor U11036 (N_11036,N_10667,N_10422);
nor U11037 (N_11037,N_10238,N_10223);
nor U11038 (N_11038,N_10536,N_10962);
nor U11039 (N_11039,N_10556,N_10650);
nor U11040 (N_11040,N_10600,N_10201);
nand U11041 (N_11041,N_10215,N_10753);
and U11042 (N_11042,N_10111,N_10493);
nor U11043 (N_11043,N_10630,N_10000);
nor U11044 (N_11044,N_10993,N_10735);
xnor U11045 (N_11045,N_10280,N_10514);
nor U11046 (N_11046,N_10251,N_10811);
nand U11047 (N_11047,N_10665,N_10205);
nor U11048 (N_11048,N_10321,N_10581);
and U11049 (N_11049,N_10439,N_10513);
or U11050 (N_11050,N_10186,N_10323);
nand U11051 (N_11051,N_10724,N_10834);
nand U11052 (N_11052,N_10203,N_10197);
nor U11053 (N_11053,N_10249,N_10069);
xor U11054 (N_11054,N_10803,N_10225);
xor U11055 (N_11055,N_10030,N_10707);
and U11056 (N_11056,N_10620,N_10204);
xor U11057 (N_11057,N_10107,N_10660);
nand U11058 (N_11058,N_10234,N_10540);
nand U11059 (N_11059,N_10413,N_10796);
or U11060 (N_11060,N_10755,N_10569);
or U11061 (N_11061,N_10700,N_10176);
and U11062 (N_11062,N_10506,N_10876);
nand U11063 (N_11063,N_10781,N_10453);
or U11064 (N_11064,N_10144,N_10130);
xnor U11065 (N_11065,N_10766,N_10793);
and U11066 (N_11066,N_10524,N_10768);
xor U11067 (N_11067,N_10454,N_10751);
or U11068 (N_11068,N_10326,N_10312);
nand U11069 (N_11069,N_10752,N_10286);
xnor U11070 (N_11070,N_10999,N_10270);
and U11071 (N_11071,N_10490,N_10633);
or U11072 (N_11072,N_10515,N_10292);
nor U11073 (N_11073,N_10348,N_10659);
or U11074 (N_11074,N_10629,N_10071);
or U11075 (N_11075,N_10440,N_10988);
or U11076 (N_11076,N_10584,N_10391);
or U11077 (N_11077,N_10934,N_10098);
nand U11078 (N_11078,N_10928,N_10310);
and U11079 (N_11079,N_10330,N_10998);
xnor U11080 (N_11080,N_10239,N_10940);
xor U11081 (N_11081,N_10479,N_10702);
nand U11082 (N_11082,N_10703,N_10854);
nor U11083 (N_11083,N_10279,N_10100);
nor U11084 (N_11084,N_10727,N_10362);
nor U11085 (N_11085,N_10587,N_10193);
nor U11086 (N_11086,N_10229,N_10738);
and U11087 (N_11087,N_10077,N_10188);
or U11088 (N_11088,N_10123,N_10561);
nor U11089 (N_11089,N_10133,N_10941);
nand U11090 (N_11090,N_10282,N_10520);
and U11091 (N_11091,N_10820,N_10115);
nand U11092 (N_11092,N_10414,N_10977);
xnor U11093 (N_11093,N_10745,N_10083);
nor U11094 (N_11094,N_10331,N_10257);
xnor U11095 (N_11095,N_10340,N_10390);
nand U11096 (N_11096,N_10687,N_10711);
xnor U11097 (N_11097,N_10746,N_10099);
nand U11098 (N_11098,N_10638,N_10956);
nor U11099 (N_11099,N_10149,N_10783);
nor U11100 (N_11100,N_10597,N_10498);
xor U11101 (N_11101,N_10301,N_10849);
or U11102 (N_11102,N_10325,N_10045);
and U11103 (N_11103,N_10145,N_10079);
or U11104 (N_11104,N_10332,N_10829);
and U11105 (N_11105,N_10392,N_10882);
or U11106 (N_11106,N_10258,N_10168);
nand U11107 (N_11107,N_10858,N_10915);
xnor U11108 (N_11108,N_10139,N_10343);
xnor U11109 (N_11109,N_10241,N_10823);
and U11110 (N_11110,N_10002,N_10120);
or U11111 (N_11111,N_10911,N_10161);
nand U11112 (N_11112,N_10012,N_10929);
xnor U11113 (N_11113,N_10539,N_10973);
nor U11114 (N_11114,N_10966,N_10690);
or U11115 (N_11115,N_10626,N_10812);
xor U11116 (N_11116,N_10445,N_10471);
nand U11117 (N_11117,N_10029,N_10798);
or U11118 (N_11118,N_10995,N_10109);
or U11119 (N_11119,N_10954,N_10612);
xnor U11120 (N_11120,N_10965,N_10532);
nand U11121 (N_11121,N_10042,N_10360);
and U11122 (N_11122,N_10760,N_10943);
and U11123 (N_11123,N_10470,N_10619);
or U11124 (N_11124,N_10463,N_10642);
nor U11125 (N_11125,N_10737,N_10299);
nand U11126 (N_11126,N_10624,N_10712);
xor U11127 (N_11127,N_10554,N_10723);
or U11128 (N_11128,N_10958,N_10676);
nor U11129 (N_11129,N_10648,N_10405);
xnor U11130 (N_11130,N_10418,N_10319);
and U11131 (N_11131,N_10064,N_10541);
xor U11132 (N_11132,N_10592,N_10231);
nand U11133 (N_11133,N_10936,N_10884);
or U11134 (N_11134,N_10932,N_10713);
nand U11135 (N_11135,N_10827,N_10086);
xnor U11136 (N_11136,N_10226,N_10574);
nor U11137 (N_11137,N_10371,N_10222);
and U11138 (N_11138,N_10865,N_10183);
or U11139 (N_11139,N_10281,N_10106);
xnor U11140 (N_11140,N_10860,N_10549);
xor U11141 (N_11141,N_10035,N_10246);
and U11142 (N_11142,N_10433,N_10489);
nand U11143 (N_11143,N_10156,N_10992);
xnor U11144 (N_11144,N_10873,N_10864);
nand U11145 (N_11145,N_10160,N_10169);
nand U11146 (N_11146,N_10023,N_10611);
and U11147 (N_11147,N_10285,N_10949);
nand U11148 (N_11148,N_10682,N_10788);
nand U11149 (N_11149,N_10428,N_10244);
nor U11150 (N_11150,N_10779,N_10082);
or U11151 (N_11151,N_10434,N_10076);
nor U11152 (N_11152,N_10774,N_10604);
xnor U11153 (N_11153,N_10385,N_10322);
and U11154 (N_11154,N_10232,N_10870);
nor U11155 (N_11155,N_10997,N_10780);
nor U11156 (N_11156,N_10656,N_10698);
nand U11157 (N_11157,N_10488,N_10664);
and U11158 (N_11158,N_10840,N_10072);
and U11159 (N_11159,N_10345,N_10990);
nor U11160 (N_11160,N_10128,N_10112);
or U11161 (N_11161,N_10741,N_10897);
and U11162 (N_11162,N_10119,N_10852);
nor U11163 (N_11163,N_10294,N_10763);
nor U11164 (N_11164,N_10705,N_10138);
and U11165 (N_11165,N_10274,N_10333);
or U11166 (N_11166,N_10913,N_10919);
nand U11167 (N_11167,N_10987,N_10757);
and U11168 (N_11168,N_10375,N_10734);
xnor U11169 (N_11169,N_10887,N_10591);
xor U11170 (N_11170,N_10177,N_10399);
nand U11171 (N_11171,N_10363,N_10314);
xnor U11172 (N_11172,N_10804,N_10484);
nand U11173 (N_11173,N_10228,N_10533);
nor U11174 (N_11174,N_10930,N_10959);
xnor U11175 (N_11175,N_10442,N_10105);
xor U11176 (N_11176,N_10551,N_10866);
nor U11177 (N_11177,N_10015,N_10625);
nand U11178 (N_11178,N_10066,N_10770);
nand U11179 (N_11179,N_10057,N_10568);
nor U11180 (N_11180,N_10437,N_10743);
nor U11181 (N_11181,N_10383,N_10481);
nand U11182 (N_11182,N_10802,N_10869);
nand U11183 (N_11183,N_10609,N_10825);
or U11184 (N_11184,N_10606,N_10353);
or U11185 (N_11185,N_10589,N_10978);
xnor U11186 (N_11186,N_10837,N_10933);
nand U11187 (N_11187,N_10486,N_10179);
nand U11188 (N_11188,N_10821,N_10557);
or U11189 (N_11189,N_10469,N_10769);
xnor U11190 (N_11190,N_10267,N_10103);
or U11191 (N_11191,N_10338,N_10021);
or U11192 (N_11192,N_10276,N_10447);
or U11193 (N_11193,N_10510,N_10907);
and U11194 (N_11194,N_10318,N_10839);
nor U11195 (N_11195,N_10902,N_10594);
xor U11196 (N_11196,N_10792,N_10657);
nand U11197 (N_11197,N_10019,N_10598);
or U11198 (N_11198,N_10585,N_10679);
and U11199 (N_11199,N_10218,N_10875);
or U11200 (N_11200,N_10038,N_10908);
nor U11201 (N_11201,N_10635,N_10491);
or U11202 (N_11202,N_10032,N_10688);
nor U11203 (N_11203,N_10061,N_10474);
nand U11204 (N_11204,N_10708,N_10068);
or U11205 (N_11205,N_10423,N_10354);
xor U11206 (N_11206,N_10003,N_10634);
nor U11207 (N_11207,N_10369,N_10221);
or U11208 (N_11208,N_10189,N_10843);
nand U11209 (N_11209,N_10302,N_10808);
or U11210 (N_11210,N_10050,N_10216);
and U11211 (N_11211,N_10980,N_10847);
and U11212 (N_11212,N_10262,N_10129);
xor U11213 (N_11213,N_10078,N_10455);
xnor U11214 (N_11214,N_10277,N_10555);
xnor U11215 (N_11215,N_10994,N_10334);
or U11216 (N_11216,N_10028,N_10164);
xor U11217 (N_11217,N_10534,N_10344);
or U11218 (N_11218,N_10607,N_10717);
xor U11219 (N_11219,N_10548,N_10576);
xnor U11220 (N_11220,N_10347,N_10947);
nand U11221 (N_11221,N_10976,N_10773);
or U11222 (N_11222,N_10170,N_10148);
nand U11223 (N_11223,N_10939,N_10298);
or U11224 (N_11224,N_10850,N_10867);
and U11225 (N_11225,N_10904,N_10173);
xnor U11226 (N_11226,N_10945,N_10521);
or U11227 (N_11227,N_10674,N_10394);
nand U11228 (N_11228,N_10181,N_10255);
and U11229 (N_11229,N_10503,N_10208);
nand U11230 (N_11230,N_10646,N_10043);
nor U11231 (N_11231,N_10706,N_10899);
or U11232 (N_11232,N_10272,N_10153);
and U11233 (N_11233,N_10715,N_10951);
and U11234 (N_11234,N_10288,N_10888);
nand U11235 (N_11235,N_10242,N_10311);
xnor U11236 (N_11236,N_10639,N_10652);
nand U11237 (N_11237,N_10252,N_10579);
xor U11238 (N_11238,N_10681,N_10158);
or U11239 (N_11239,N_10154,N_10608);
nor U11240 (N_11240,N_10134,N_10694);
and U11241 (N_11241,N_10531,N_10718);
and U11242 (N_11242,N_10795,N_10826);
and U11243 (N_11243,N_10141,N_10563);
or U11244 (N_11244,N_10601,N_10283);
and U11245 (N_11245,N_10878,N_10461);
xor U11246 (N_11246,N_10235,N_10778);
xor U11247 (N_11247,N_10157,N_10580);
nand U11248 (N_11248,N_10001,N_10341);
nor U11249 (N_11249,N_10230,N_10517);
xor U11250 (N_11250,N_10836,N_10500);
nor U11251 (N_11251,N_10684,N_10142);
xor U11252 (N_11252,N_10784,N_10614);
xnor U11253 (N_11253,N_10658,N_10008);
nor U11254 (N_11254,N_10031,N_10421);
nor U11255 (N_11255,N_10883,N_10048);
and U11256 (N_11256,N_10572,N_10906);
or U11257 (N_11257,N_10957,N_10357);
and U11258 (N_11258,N_10605,N_10182);
nand U11259 (N_11259,N_10009,N_10689);
nor U11260 (N_11260,N_10449,N_10801);
xnor U11261 (N_11261,N_10575,N_10448);
nand U11262 (N_11262,N_10944,N_10400);
nand U11263 (N_11263,N_10508,N_10617);
nor U11264 (N_11264,N_10213,N_10814);
and U11265 (N_11265,N_10497,N_10942);
nand U11266 (N_11266,N_10663,N_10441);
or U11267 (N_11267,N_10830,N_10126);
xnor U11268 (N_11268,N_10645,N_10473);
or U11269 (N_11269,N_10742,N_10996);
and U11270 (N_11270,N_10914,N_10004);
xnor U11271 (N_11271,N_10260,N_10761);
and U11272 (N_11272,N_10458,N_10668);
xor U11273 (N_11273,N_10926,N_10404);
nor U11274 (N_11274,N_10917,N_10599);
nand U11275 (N_11275,N_10088,N_10296);
nor U11276 (N_11276,N_10200,N_10284);
and U11277 (N_11277,N_10628,N_10398);
nor U11278 (N_11278,N_10196,N_10430);
nand U11279 (N_11279,N_10673,N_10198);
nor U11280 (N_11280,N_10351,N_10336);
nand U11281 (N_11281,N_10227,N_10456);
nor U11282 (N_11282,N_10162,N_10545);
or U11283 (N_11283,N_10452,N_10451);
nand U11284 (N_11284,N_10699,N_10528);
and U11285 (N_11285,N_10910,N_10799);
nand U11286 (N_11286,N_10370,N_10859);
or U11287 (N_11287,N_10135,N_10838);
or U11288 (N_11288,N_10806,N_10982);
nor U11289 (N_11289,N_10955,N_10127);
xnor U11290 (N_11290,N_10693,N_10492);
or U11291 (N_11291,N_10683,N_10046);
nand U11292 (N_11292,N_10155,N_10662);
nor U11293 (N_11293,N_10805,N_10677);
xor U11294 (N_11294,N_10559,N_10337);
or U11295 (N_11295,N_10163,N_10765);
and U11296 (N_11296,N_10195,N_10546);
nor U11297 (N_11297,N_10494,N_10327);
xor U11298 (N_11298,N_10759,N_10016);
or U11299 (N_11299,N_10691,N_10905);
nor U11300 (N_11300,N_10948,N_10150);
xor U11301 (N_11301,N_10263,N_10113);
and U11302 (N_11302,N_10364,N_10790);
xor U11303 (N_11303,N_10243,N_10863);
nor U11304 (N_11304,N_10872,N_10975);
and U11305 (N_11305,N_10395,N_10352);
or U11306 (N_11306,N_10438,N_10467);
or U11307 (N_11307,N_10206,N_10373);
or U11308 (N_11308,N_10496,N_10041);
nand U11309 (N_11309,N_10217,N_10603);
xor U11310 (N_11310,N_10307,N_10080);
nor U11311 (N_11311,N_10695,N_10219);
or U11312 (N_11312,N_10101,N_10530);
and U11313 (N_11313,N_10610,N_10961);
xnor U11314 (N_11314,N_10721,N_10049);
and U11315 (N_11315,N_10317,N_10081);
xnor U11316 (N_11316,N_10409,N_10654);
xor U11317 (N_11317,N_10502,N_10807);
xnor U11318 (N_11318,N_10631,N_10748);
xor U11319 (N_11319,N_10297,N_10845);
and U11320 (N_11320,N_10117,N_10058);
nor U11321 (N_11321,N_10828,N_10512);
nand U11322 (N_11322,N_10543,N_10671);
nand U11323 (N_11323,N_10507,N_10468);
xnor U11324 (N_11324,N_10641,N_10726);
or U11325 (N_11325,N_10810,N_10295);
nand U11326 (N_11326,N_10056,N_10655);
nor U11327 (N_11327,N_10220,N_10709);
or U11328 (N_11328,N_10722,N_10732);
xnor U11329 (N_11329,N_10719,N_10720);
nand U11330 (N_11330,N_10367,N_10480);
or U11331 (N_11331,N_10381,N_10637);
nor U11332 (N_11332,N_10925,N_10037);
and U11333 (N_11333,N_10842,N_10782);
nand U11334 (N_11334,N_10393,N_10397);
xor U11335 (N_11335,N_10147,N_10892);
nor U11336 (N_11336,N_10237,N_10178);
or U11337 (N_11337,N_10026,N_10483);
and U11338 (N_11338,N_10025,N_10901);
nand U11339 (N_11339,N_10509,N_10552);
nor U11340 (N_11340,N_10979,N_10504);
or U11341 (N_11341,N_10207,N_10131);
or U11342 (N_11342,N_10921,N_10643);
nand U11343 (N_11343,N_10647,N_10747);
or U11344 (N_11344,N_10010,N_10387);
nor U11345 (N_11345,N_10254,N_10593);
or U11346 (N_11346,N_10287,N_10935);
nor U11347 (N_11347,N_10187,N_10478);
nand U11348 (N_11348,N_10920,N_10240);
xor U11349 (N_11349,N_10202,N_10818);
or U11350 (N_11350,N_10984,N_10791);
and U11351 (N_11351,N_10005,N_10855);
xnor U11352 (N_11352,N_10516,N_10819);
xnor U11353 (N_11353,N_10590,N_10462);
xnor U11354 (N_11354,N_10419,N_10020);
or U11355 (N_11355,N_10640,N_10896);
nor U11356 (N_11356,N_10623,N_10339);
and U11357 (N_11357,N_10143,N_10313);
nor U11358 (N_11358,N_10388,N_10034);
or U11359 (N_11359,N_10680,N_10096);
and U11360 (N_11360,N_10578,N_10562);
and U11361 (N_11361,N_10716,N_10909);
nor U11362 (N_11362,N_10040,N_10527);
nor U11363 (N_11363,N_10417,N_10379);
xor U11364 (N_11364,N_10560,N_10848);
nand U11365 (N_11365,N_10269,N_10881);
nand U11366 (N_11366,N_10089,N_10022);
or U11367 (N_11367,N_10733,N_10501);
nand U11368 (N_11368,N_10675,N_10583);
or U11369 (N_11369,N_10476,N_10211);
xor U11370 (N_11370,N_10425,N_10114);
and U11371 (N_11371,N_10090,N_10800);
nand U11372 (N_11372,N_10816,N_10877);
nor U11373 (N_11373,N_10885,N_10359);
nor U11374 (N_11374,N_10407,N_10927);
and U11375 (N_11375,N_10011,N_10410);
and U11376 (N_11376,N_10558,N_10710);
or U11377 (N_11377,N_10446,N_10475);
nand U11378 (N_11378,N_10092,N_10797);
nor U11379 (N_11379,N_10986,N_10964);
nor U11380 (N_11380,N_10018,N_10776);
and U11381 (N_11381,N_10764,N_10194);
nand U11382 (N_11382,N_10014,N_10406);
or U11383 (N_11383,N_10073,N_10756);
and U11384 (N_11384,N_10749,N_10054);
nor U11385 (N_11385,N_10853,N_10924);
or U11386 (N_11386,N_10027,N_10271);
or U11387 (N_11387,N_10894,N_10912);
nor U11388 (N_11388,N_10324,N_10886);
nor U11389 (N_11389,N_10596,N_10895);
nand U11390 (N_11390,N_10124,N_10006);
xor U11391 (N_11391,N_10328,N_10871);
and U11392 (N_11392,N_10097,N_10431);
nand U11393 (N_11393,N_10291,N_10567);
or U11394 (N_11394,N_10952,N_10315);
nand U11395 (N_11395,N_10408,N_10731);
nor U11396 (N_11396,N_10518,N_10308);
nor U11397 (N_11397,N_10140,N_10465);
nand U11398 (N_11398,N_10396,N_10382);
xor U11399 (N_11399,N_10714,N_10304);
nor U11400 (N_11400,N_10316,N_10519);
and U11401 (N_11401,N_10963,N_10055);
nor U11402 (N_11402,N_10972,N_10991);
or U11403 (N_11403,N_10772,N_10686);
and U11404 (N_11404,N_10728,N_10771);
or U11405 (N_11405,N_10365,N_10136);
and U11406 (N_11406,N_10861,N_10550);
and U11407 (N_11407,N_10175,N_10047);
nor U11408 (N_11408,N_10116,N_10420);
or U11409 (N_11409,N_10210,N_10487);
nand U11410 (N_11410,N_10429,N_10377);
nand U11411 (N_11411,N_10358,N_10566);
or U11412 (N_11412,N_10320,N_10151);
nand U11413 (N_11413,N_10074,N_10616);
nor U11414 (N_11414,N_10900,N_10744);
and U11415 (N_11415,N_10132,N_10167);
xor U11416 (N_11416,N_10787,N_10666);
nand U11417 (N_11417,N_10967,N_10146);
nand U11418 (N_11418,N_10435,N_10137);
or U11419 (N_11419,N_10033,N_10386);
or U11420 (N_11420,N_10922,N_10261);
xnor U11421 (N_11421,N_10248,N_10190);
nand U11422 (N_11422,N_10355,N_10851);
xnor U11423 (N_11423,N_10044,N_10729);
nor U11424 (N_11424,N_10366,N_10582);
nor U11425 (N_11425,N_10636,N_10649);
and U11426 (N_11426,N_10511,N_10075);
xor U11427 (N_11427,N_10460,N_10070);
xor U11428 (N_11428,N_10815,N_10245);
xor U11429 (N_11429,N_10953,N_10477);
and U11430 (N_11430,N_10529,N_10165);
and U11431 (N_11431,N_10180,N_10415);
or U11432 (N_11432,N_10172,N_10466);
xnor U11433 (N_11433,N_10824,N_10290);
and U11434 (N_11434,N_10661,N_10696);
nor U11435 (N_11435,N_10356,N_10063);
nor U11436 (N_11436,N_10692,N_10817);
and U11437 (N_11437,N_10121,N_10342);
nand U11438 (N_11438,N_10199,N_10350);
nand U11439 (N_11439,N_10432,N_10166);
and U11440 (N_11440,N_10024,N_10785);
and U11441 (N_11441,N_10758,N_10013);
nand U11442 (N_11442,N_10891,N_10577);
nand U11443 (N_11443,N_10621,N_10678);
nor U11444 (N_11444,N_10017,N_10505);
nor U11445 (N_11445,N_10701,N_10672);
and U11446 (N_11446,N_10171,N_10152);
nor U11447 (N_11447,N_10095,N_10403);
xor U11448 (N_11448,N_10185,N_10739);
nor U11449 (N_11449,N_10256,N_10968);
or U11450 (N_11450,N_10586,N_10969);
and U11451 (N_11451,N_10632,N_10361);
nand U11452 (N_11452,N_10499,N_10669);
nor U11453 (N_11453,N_10250,N_10835);
nand U11454 (N_11454,N_10052,N_10411);
nand U11455 (N_11455,N_10813,N_10368);
nor U11456 (N_11456,N_10651,N_10974);
or U11457 (N_11457,N_10424,N_10264);
xnor U11458 (N_11458,N_10831,N_10571);
or U11459 (N_11459,N_10426,N_10329);
xnor U11460 (N_11460,N_10740,N_10553);
nand U11461 (N_11461,N_10053,N_10525);
xor U11462 (N_11462,N_10918,N_10192);
nand U11463 (N_11463,N_10062,N_10085);
xor U11464 (N_11464,N_10472,N_10916);
xnor U11465 (N_11465,N_10789,N_10412);
xor U11466 (N_11466,N_10989,N_10889);
xnor U11467 (N_11467,N_10950,N_10862);
or U11468 (N_11468,N_10833,N_10464);
and U11469 (N_11469,N_10777,N_10459);
or U11470 (N_11470,N_10273,N_10457);
nor U11471 (N_11471,N_10588,N_10104);
nand U11472 (N_11472,N_10937,N_10564);
nor U11473 (N_11473,N_10401,N_10523);
nand U11474 (N_11474,N_10384,N_10522);
or U11475 (N_11475,N_10209,N_10846);
xnor U11476 (N_11476,N_10427,N_10841);
or U11477 (N_11477,N_10060,N_10125);
xnor U11478 (N_11478,N_10247,N_10303);
nand U11479 (N_11479,N_10880,N_10289);
nand U11480 (N_11480,N_10595,N_10376);
or U11481 (N_11481,N_10931,N_10898);
and U11482 (N_11482,N_10259,N_10822);
or U11483 (N_11483,N_10266,N_10102);
or U11484 (N_11484,N_10981,N_10306);
nor U11485 (N_11485,N_10214,N_10754);
and U11486 (N_11486,N_10544,N_10615);
nand U11487 (N_11487,N_10108,N_10159);
and U11488 (N_11488,N_10051,N_10300);
and U11489 (N_11489,N_10526,N_10903);
xor U11490 (N_11490,N_10293,N_10573);
nand U11491 (N_11491,N_10622,N_10923);
nand U11492 (N_11492,N_10960,N_10278);
nor U11493 (N_11493,N_10067,N_10890);
or U11494 (N_11494,N_10685,N_10844);
nand U11495 (N_11495,N_10346,N_10730);
nor U11496 (N_11496,N_10750,N_10093);
xnor U11497 (N_11497,N_10094,N_10704);
xor U11498 (N_11498,N_10618,N_10212);
nand U11499 (N_11499,N_10794,N_10275);
nor U11500 (N_11500,N_10390,N_10296);
xnor U11501 (N_11501,N_10162,N_10071);
nand U11502 (N_11502,N_10080,N_10473);
nor U11503 (N_11503,N_10292,N_10615);
and U11504 (N_11504,N_10669,N_10012);
and U11505 (N_11505,N_10855,N_10581);
or U11506 (N_11506,N_10806,N_10367);
xor U11507 (N_11507,N_10123,N_10474);
nor U11508 (N_11508,N_10245,N_10754);
or U11509 (N_11509,N_10190,N_10612);
and U11510 (N_11510,N_10939,N_10192);
or U11511 (N_11511,N_10381,N_10074);
nor U11512 (N_11512,N_10984,N_10801);
or U11513 (N_11513,N_10754,N_10576);
and U11514 (N_11514,N_10817,N_10359);
nand U11515 (N_11515,N_10934,N_10994);
nand U11516 (N_11516,N_10309,N_10004);
and U11517 (N_11517,N_10247,N_10105);
and U11518 (N_11518,N_10941,N_10063);
and U11519 (N_11519,N_10699,N_10643);
nor U11520 (N_11520,N_10732,N_10602);
nand U11521 (N_11521,N_10125,N_10502);
nand U11522 (N_11522,N_10799,N_10902);
and U11523 (N_11523,N_10032,N_10216);
nand U11524 (N_11524,N_10809,N_10265);
and U11525 (N_11525,N_10031,N_10674);
nor U11526 (N_11526,N_10420,N_10437);
or U11527 (N_11527,N_10242,N_10758);
nand U11528 (N_11528,N_10251,N_10857);
nor U11529 (N_11529,N_10222,N_10167);
nor U11530 (N_11530,N_10622,N_10039);
nor U11531 (N_11531,N_10613,N_10173);
nand U11532 (N_11532,N_10663,N_10886);
and U11533 (N_11533,N_10274,N_10770);
nor U11534 (N_11534,N_10654,N_10018);
nor U11535 (N_11535,N_10528,N_10297);
and U11536 (N_11536,N_10407,N_10395);
xnor U11537 (N_11537,N_10791,N_10713);
xnor U11538 (N_11538,N_10473,N_10757);
or U11539 (N_11539,N_10873,N_10208);
nor U11540 (N_11540,N_10759,N_10326);
and U11541 (N_11541,N_10609,N_10396);
xnor U11542 (N_11542,N_10975,N_10934);
nand U11543 (N_11543,N_10990,N_10413);
nand U11544 (N_11544,N_10199,N_10946);
nand U11545 (N_11545,N_10134,N_10655);
or U11546 (N_11546,N_10710,N_10676);
xor U11547 (N_11547,N_10783,N_10053);
nor U11548 (N_11548,N_10949,N_10200);
nand U11549 (N_11549,N_10401,N_10185);
xor U11550 (N_11550,N_10060,N_10704);
nor U11551 (N_11551,N_10475,N_10854);
xor U11552 (N_11552,N_10975,N_10244);
xnor U11553 (N_11553,N_10809,N_10410);
and U11554 (N_11554,N_10657,N_10439);
nor U11555 (N_11555,N_10298,N_10673);
and U11556 (N_11556,N_10192,N_10419);
and U11557 (N_11557,N_10461,N_10784);
and U11558 (N_11558,N_10532,N_10598);
or U11559 (N_11559,N_10683,N_10787);
or U11560 (N_11560,N_10286,N_10597);
xnor U11561 (N_11561,N_10680,N_10013);
or U11562 (N_11562,N_10909,N_10796);
and U11563 (N_11563,N_10780,N_10864);
or U11564 (N_11564,N_10270,N_10417);
nor U11565 (N_11565,N_10100,N_10943);
and U11566 (N_11566,N_10926,N_10991);
xor U11567 (N_11567,N_10681,N_10709);
or U11568 (N_11568,N_10337,N_10709);
or U11569 (N_11569,N_10322,N_10618);
or U11570 (N_11570,N_10673,N_10737);
nand U11571 (N_11571,N_10078,N_10935);
or U11572 (N_11572,N_10511,N_10365);
nor U11573 (N_11573,N_10586,N_10872);
and U11574 (N_11574,N_10734,N_10799);
xor U11575 (N_11575,N_10954,N_10987);
nor U11576 (N_11576,N_10285,N_10813);
nor U11577 (N_11577,N_10550,N_10633);
or U11578 (N_11578,N_10591,N_10205);
nor U11579 (N_11579,N_10076,N_10572);
xor U11580 (N_11580,N_10501,N_10122);
nor U11581 (N_11581,N_10426,N_10119);
nand U11582 (N_11582,N_10782,N_10455);
nand U11583 (N_11583,N_10986,N_10631);
nor U11584 (N_11584,N_10714,N_10068);
and U11585 (N_11585,N_10827,N_10963);
xnor U11586 (N_11586,N_10747,N_10088);
or U11587 (N_11587,N_10419,N_10685);
or U11588 (N_11588,N_10762,N_10351);
nor U11589 (N_11589,N_10966,N_10150);
or U11590 (N_11590,N_10988,N_10477);
nand U11591 (N_11591,N_10638,N_10516);
and U11592 (N_11592,N_10298,N_10460);
and U11593 (N_11593,N_10481,N_10938);
xor U11594 (N_11594,N_10896,N_10428);
nor U11595 (N_11595,N_10918,N_10553);
and U11596 (N_11596,N_10412,N_10648);
nand U11597 (N_11597,N_10114,N_10015);
nand U11598 (N_11598,N_10425,N_10150);
or U11599 (N_11599,N_10437,N_10213);
and U11600 (N_11600,N_10818,N_10986);
or U11601 (N_11601,N_10282,N_10878);
xnor U11602 (N_11602,N_10502,N_10338);
nand U11603 (N_11603,N_10488,N_10761);
or U11604 (N_11604,N_10291,N_10740);
xnor U11605 (N_11605,N_10863,N_10747);
nor U11606 (N_11606,N_10424,N_10325);
nand U11607 (N_11607,N_10559,N_10374);
nor U11608 (N_11608,N_10661,N_10185);
xor U11609 (N_11609,N_10602,N_10938);
nor U11610 (N_11610,N_10717,N_10103);
xnor U11611 (N_11611,N_10298,N_10085);
and U11612 (N_11612,N_10976,N_10790);
xor U11613 (N_11613,N_10378,N_10041);
or U11614 (N_11614,N_10298,N_10053);
or U11615 (N_11615,N_10854,N_10620);
and U11616 (N_11616,N_10266,N_10742);
xnor U11617 (N_11617,N_10127,N_10628);
or U11618 (N_11618,N_10008,N_10101);
and U11619 (N_11619,N_10118,N_10862);
nand U11620 (N_11620,N_10658,N_10810);
or U11621 (N_11621,N_10283,N_10955);
nor U11622 (N_11622,N_10971,N_10282);
and U11623 (N_11623,N_10699,N_10447);
and U11624 (N_11624,N_10910,N_10260);
and U11625 (N_11625,N_10336,N_10520);
or U11626 (N_11626,N_10232,N_10155);
or U11627 (N_11627,N_10962,N_10075);
nand U11628 (N_11628,N_10528,N_10079);
and U11629 (N_11629,N_10134,N_10843);
or U11630 (N_11630,N_10342,N_10400);
or U11631 (N_11631,N_10086,N_10798);
xor U11632 (N_11632,N_10464,N_10110);
nand U11633 (N_11633,N_10870,N_10438);
or U11634 (N_11634,N_10152,N_10333);
and U11635 (N_11635,N_10672,N_10942);
nor U11636 (N_11636,N_10486,N_10562);
xor U11637 (N_11637,N_10191,N_10102);
xnor U11638 (N_11638,N_10008,N_10859);
xor U11639 (N_11639,N_10727,N_10397);
and U11640 (N_11640,N_10708,N_10304);
nand U11641 (N_11641,N_10674,N_10048);
nor U11642 (N_11642,N_10674,N_10897);
or U11643 (N_11643,N_10690,N_10906);
and U11644 (N_11644,N_10765,N_10776);
or U11645 (N_11645,N_10659,N_10878);
xor U11646 (N_11646,N_10064,N_10809);
and U11647 (N_11647,N_10250,N_10382);
nor U11648 (N_11648,N_10290,N_10556);
nor U11649 (N_11649,N_10556,N_10087);
and U11650 (N_11650,N_10867,N_10291);
and U11651 (N_11651,N_10703,N_10244);
nor U11652 (N_11652,N_10424,N_10192);
or U11653 (N_11653,N_10416,N_10102);
nand U11654 (N_11654,N_10856,N_10982);
nor U11655 (N_11655,N_10875,N_10685);
xnor U11656 (N_11656,N_10983,N_10867);
nand U11657 (N_11657,N_10534,N_10193);
xor U11658 (N_11658,N_10126,N_10072);
nand U11659 (N_11659,N_10421,N_10512);
or U11660 (N_11660,N_10783,N_10457);
and U11661 (N_11661,N_10568,N_10585);
and U11662 (N_11662,N_10373,N_10476);
and U11663 (N_11663,N_10471,N_10935);
xor U11664 (N_11664,N_10282,N_10244);
and U11665 (N_11665,N_10466,N_10332);
xnor U11666 (N_11666,N_10402,N_10577);
or U11667 (N_11667,N_10673,N_10019);
or U11668 (N_11668,N_10949,N_10624);
and U11669 (N_11669,N_10220,N_10382);
nor U11670 (N_11670,N_10258,N_10188);
or U11671 (N_11671,N_10126,N_10102);
or U11672 (N_11672,N_10283,N_10895);
nand U11673 (N_11673,N_10672,N_10818);
and U11674 (N_11674,N_10533,N_10379);
or U11675 (N_11675,N_10746,N_10840);
or U11676 (N_11676,N_10562,N_10725);
nand U11677 (N_11677,N_10752,N_10619);
nand U11678 (N_11678,N_10954,N_10679);
xnor U11679 (N_11679,N_10434,N_10258);
xor U11680 (N_11680,N_10713,N_10304);
xor U11681 (N_11681,N_10314,N_10882);
nor U11682 (N_11682,N_10580,N_10908);
or U11683 (N_11683,N_10650,N_10851);
and U11684 (N_11684,N_10481,N_10387);
xnor U11685 (N_11685,N_10652,N_10039);
nor U11686 (N_11686,N_10428,N_10471);
nor U11687 (N_11687,N_10292,N_10409);
nand U11688 (N_11688,N_10564,N_10821);
xor U11689 (N_11689,N_10158,N_10191);
xnor U11690 (N_11690,N_10138,N_10356);
xnor U11691 (N_11691,N_10791,N_10516);
and U11692 (N_11692,N_10759,N_10543);
or U11693 (N_11693,N_10844,N_10825);
xnor U11694 (N_11694,N_10514,N_10873);
nor U11695 (N_11695,N_10749,N_10941);
and U11696 (N_11696,N_10075,N_10578);
nor U11697 (N_11697,N_10032,N_10135);
xor U11698 (N_11698,N_10944,N_10505);
xnor U11699 (N_11699,N_10921,N_10523);
nand U11700 (N_11700,N_10906,N_10542);
nand U11701 (N_11701,N_10427,N_10177);
nor U11702 (N_11702,N_10997,N_10992);
nor U11703 (N_11703,N_10742,N_10616);
or U11704 (N_11704,N_10910,N_10263);
nor U11705 (N_11705,N_10603,N_10630);
or U11706 (N_11706,N_10191,N_10090);
and U11707 (N_11707,N_10487,N_10453);
and U11708 (N_11708,N_10096,N_10597);
xor U11709 (N_11709,N_10473,N_10172);
and U11710 (N_11710,N_10962,N_10769);
nand U11711 (N_11711,N_10742,N_10769);
xor U11712 (N_11712,N_10973,N_10911);
nor U11713 (N_11713,N_10214,N_10769);
nand U11714 (N_11714,N_10303,N_10298);
xor U11715 (N_11715,N_10794,N_10568);
xnor U11716 (N_11716,N_10008,N_10997);
xnor U11717 (N_11717,N_10026,N_10385);
xnor U11718 (N_11718,N_10561,N_10950);
xnor U11719 (N_11719,N_10033,N_10074);
nand U11720 (N_11720,N_10309,N_10024);
nor U11721 (N_11721,N_10359,N_10957);
and U11722 (N_11722,N_10358,N_10495);
and U11723 (N_11723,N_10051,N_10318);
xor U11724 (N_11724,N_10444,N_10737);
nand U11725 (N_11725,N_10394,N_10618);
or U11726 (N_11726,N_10957,N_10083);
or U11727 (N_11727,N_10398,N_10744);
nor U11728 (N_11728,N_10558,N_10254);
nand U11729 (N_11729,N_10779,N_10538);
xnor U11730 (N_11730,N_10418,N_10257);
and U11731 (N_11731,N_10162,N_10647);
and U11732 (N_11732,N_10597,N_10795);
or U11733 (N_11733,N_10257,N_10723);
and U11734 (N_11734,N_10572,N_10077);
and U11735 (N_11735,N_10362,N_10918);
nor U11736 (N_11736,N_10307,N_10905);
and U11737 (N_11737,N_10893,N_10813);
or U11738 (N_11738,N_10449,N_10322);
nand U11739 (N_11739,N_10110,N_10391);
or U11740 (N_11740,N_10424,N_10971);
or U11741 (N_11741,N_10709,N_10285);
and U11742 (N_11742,N_10282,N_10432);
or U11743 (N_11743,N_10452,N_10915);
and U11744 (N_11744,N_10379,N_10423);
nor U11745 (N_11745,N_10011,N_10279);
and U11746 (N_11746,N_10911,N_10520);
nor U11747 (N_11747,N_10715,N_10933);
and U11748 (N_11748,N_10435,N_10605);
or U11749 (N_11749,N_10374,N_10356);
and U11750 (N_11750,N_10953,N_10547);
nor U11751 (N_11751,N_10685,N_10767);
xnor U11752 (N_11752,N_10395,N_10775);
nand U11753 (N_11753,N_10747,N_10726);
or U11754 (N_11754,N_10088,N_10865);
or U11755 (N_11755,N_10643,N_10029);
and U11756 (N_11756,N_10871,N_10065);
nor U11757 (N_11757,N_10791,N_10369);
nor U11758 (N_11758,N_10506,N_10055);
or U11759 (N_11759,N_10097,N_10479);
and U11760 (N_11760,N_10115,N_10166);
and U11761 (N_11761,N_10514,N_10958);
nand U11762 (N_11762,N_10252,N_10673);
nand U11763 (N_11763,N_10960,N_10902);
xor U11764 (N_11764,N_10499,N_10335);
nand U11765 (N_11765,N_10404,N_10359);
and U11766 (N_11766,N_10388,N_10772);
or U11767 (N_11767,N_10937,N_10258);
nor U11768 (N_11768,N_10652,N_10873);
or U11769 (N_11769,N_10943,N_10901);
nand U11770 (N_11770,N_10105,N_10549);
or U11771 (N_11771,N_10465,N_10692);
nor U11772 (N_11772,N_10986,N_10871);
nor U11773 (N_11773,N_10733,N_10414);
xor U11774 (N_11774,N_10125,N_10484);
or U11775 (N_11775,N_10344,N_10360);
nor U11776 (N_11776,N_10049,N_10433);
and U11777 (N_11777,N_10657,N_10840);
or U11778 (N_11778,N_10175,N_10482);
and U11779 (N_11779,N_10912,N_10958);
xnor U11780 (N_11780,N_10971,N_10793);
and U11781 (N_11781,N_10713,N_10814);
xnor U11782 (N_11782,N_10633,N_10788);
nor U11783 (N_11783,N_10958,N_10830);
xor U11784 (N_11784,N_10806,N_10499);
and U11785 (N_11785,N_10036,N_10966);
nand U11786 (N_11786,N_10815,N_10976);
xor U11787 (N_11787,N_10740,N_10536);
nand U11788 (N_11788,N_10294,N_10708);
nand U11789 (N_11789,N_10509,N_10500);
or U11790 (N_11790,N_10838,N_10890);
nor U11791 (N_11791,N_10328,N_10004);
nand U11792 (N_11792,N_10609,N_10498);
xor U11793 (N_11793,N_10079,N_10373);
or U11794 (N_11794,N_10677,N_10291);
nor U11795 (N_11795,N_10528,N_10170);
nand U11796 (N_11796,N_10529,N_10729);
xor U11797 (N_11797,N_10512,N_10472);
or U11798 (N_11798,N_10132,N_10046);
xnor U11799 (N_11799,N_10189,N_10269);
and U11800 (N_11800,N_10304,N_10098);
and U11801 (N_11801,N_10373,N_10251);
nor U11802 (N_11802,N_10152,N_10570);
nor U11803 (N_11803,N_10560,N_10051);
xnor U11804 (N_11804,N_10579,N_10502);
or U11805 (N_11805,N_10384,N_10898);
nor U11806 (N_11806,N_10771,N_10830);
xnor U11807 (N_11807,N_10744,N_10572);
or U11808 (N_11808,N_10584,N_10263);
and U11809 (N_11809,N_10268,N_10174);
or U11810 (N_11810,N_10870,N_10628);
nand U11811 (N_11811,N_10413,N_10124);
nor U11812 (N_11812,N_10588,N_10489);
nand U11813 (N_11813,N_10488,N_10273);
nand U11814 (N_11814,N_10666,N_10352);
nand U11815 (N_11815,N_10119,N_10973);
nand U11816 (N_11816,N_10404,N_10011);
or U11817 (N_11817,N_10073,N_10522);
and U11818 (N_11818,N_10741,N_10495);
nor U11819 (N_11819,N_10610,N_10606);
or U11820 (N_11820,N_10792,N_10390);
nor U11821 (N_11821,N_10064,N_10179);
or U11822 (N_11822,N_10138,N_10533);
nand U11823 (N_11823,N_10596,N_10382);
and U11824 (N_11824,N_10325,N_10467);
nand U11825 (N_11825,N_10508,N_10842);
or U11826 (N_11826,N_10219,N_10330);
or U11827 (N_11827,N_10020,N_10553);
and U11828 (N_11828,N_10904,N_10774);
nor U11829 (N_11829,N_10257,N_10982);
xor U11830 (N_11830,N_10705,N_10697);
nor U11831 (N_11831,N_10618,N_10416);
or U11832 (N_11832,N_10311,N_10002);
nand U11833 (N_11833,N_10528,N_10679);
nor U11834 (N_11834,N_10973,N_10486);
or U11835 (N_11835,N_10479,N_10934);
or U11836 (N_11836,N_10672,N_10644);
and U11837 (N_11837,N_10232,N_10390);
nand U11838 (N_11838,N_10464,N_10287);
and U11839 (N_11839,N_10150,N_10016);
xnor U11840 (N_11840,N_10982,N_10220);
xnor U11841 (N_11841,N_10636,N_10816);
or U11842 (N_11842,N_10493,N_10903);
or U11843 (N_11843,N_10411,N_10732);
nand U11844 (N_11844,N_10991,N_10953);
or U11845 (N_11845,N_10403,N_10872);
nand U11846 (N_11846,N_10270,N_10298);
and U11847 (N_11847,N_10169,N_10185);
nor U11848 (N_11848,N_10040,N_10115);
xor U11849 (N_11849,N_10460,N_10343);
nand U11850 (N_11850,N_10238,N_10770);
xnor U11851 (N_11851,N_10324,N_10018);
nor U11852 (N_11852,N_10543,N_10686);
nor U11853 (N_11853,N_10075,N_10913);
xor U11854 (N_11854,N_10232,N_10927);
nor U11855 (N_11855,N_10500,N_10381);
nand U11856 (N_11856,N_10328,N_10988);
xor U11857 (N_11857,N_10955,N_10781);
or U11858 (N_11858,N_10222,N_10543);
nand U11859 (N_11859,N_10958,N_10708);
or U11860 (N_11860,N_10962,N_10483);
and U11861 (N_11861,N_10689,N_10709);
or U11862 (N_11862,N_10379,N_10325);
nor U11863 (N_11863,N_10803,N_10742);
xor U11864 (N_11864,N_10028,N_10566);
or U11865 (N_11865,N_10921,N_10878);
nor U11866 (N_11866,N_10174,N_10694);
xor U11867 (N_11867,N_10446,N_10629);
or U11868 (N_11868,N_10686,N_10787);
nand U11869 (N_11869,N_10245,N_10352);
xnor U11870 (N_11870,N_10576,N_10763);
xnor U11871 (N_11871,N_10029,N_10669);
nor U11872 (N_11872,N_10981,N_10468);
xor U11873 (N_11873,N_10692,N_10053);
or U11874 (N_11874,N_10631,N_10358);
or U11875 (N_11875,N_10034,N_10008);
nor U11876 (N_11876,N_10802,N_10685);
xnor U11877 (N_11877,N_10824,N_10920);
nor U11878 (N_11878,N_10558,N_10514);
and U11879 (N_11879,N_10692,N_10710);
or U11880 (N_11880,N_10466,N_10437);
xor U11881 (N_11881,N_10253,N_10371);
xor U11882 (N_11882,N_10092,N_10492);
nand U11883 (N_11883,N_10956,N_10909);
or U11884 (N_11884,N_10036,N_10775);
nand U11885 (N_11885,N_10911,N_10742);
xor U11886 (N_11886,N_10420,N_10506);
xor U11887 (N_11887,N_10906,N_10266);
nand U11888 (N_11888,N_10385,N_10771);
or U11889 (N_11889,N_10941,N_10354);
or U11890 (N_11890,N_10896,N_10843);
nor U11891 (N_11891,N_10754,N_10749);
or U11892 (N_11892,N_10287,N_10148);
xnor U11893 (N_11893,N_10821,N_10580);
xor U11894 (N_11894,N_10022,N_10224);
and U11895 (N_11895,N_10775,N_10616);
and U11896 (N_11896,N_10298,N_10731);
and U11897 (N_11897,N_10365,N_10446);
or U11898 (N_11898,N_10789,N_10510);
and U11899 (N_11899,N_10482,N_10686);
and U11900 (N_11900,N_10105,N_10794);
and U11901 (N_11901,N_10361,N_10372);
nor U11902 (N_11902,N_10626,N_10421);
xnor U11903 (N_11903,N_10613,N_10456);
nor U11904 (N_11904,N_10909,N_10761);
and U11905 (N_11905,N_10537,N_10607);
or U11906 (N_11906,N_10330,N_10362);
nor U11907 (N_11907,N_10731,N_10908);
xor U11908 (N_11908,N_10433,N_10887);
or U11909 (N_11909,N_10263,N_10755);
xnor U11910 (N_11910,N_10980,N_10516);
and U11911 (N_11911,N_10627,N_10389);
nor U11912 (N_11912,N_10974,N_10663);
xnor U11913 (N_11913,N_10747,N_10266);
nor U11914 (N_11914,N_10642,N_10834);
and U11915 (N_11915,N_10893,N_10208);
nand U11916 (N_11916,N_10209,N_10196);
or U11917 (N_11917,N_10872,N_10750);
xor U11918 (N_11918,N_10348,N_10987);
xor U11919 (N_11919,N_10291,N_10739);
or U11920 (N_11920,N_10837,N_10301);
or U11921 (N_11921,N_10034,N_10046);
and U11922 (N_11922,N_10784,N_10847);
xnor U11923 (N_11923,N_10612,N_10851);
and U11924 (N_11924,N_10043,N_10609);
and U11925 (N_11925,N_10673,N_10280);
and U11926 (N_11926,N_10523,N_10928);
nand U11927 (N_11927,N_10937,N_10839);
nor U11928 (N_11928,N_10571,N_10266);
nand U11929 (N_11929,N_10611,N_10270);
nor U11930 (N_11930,N_10421,N_10670);
or U11931 (N_11931,N_10141,N_10983);
xnor U11932 (N_11932,N_10416,N_10540);
nand U11933 (N_11933,N_10133,N_10510);
nor U11934 (N_11934,N_10834,N_10955);
or U11935 (N_11935,N_10955,N_10520);
and U11936 (N_11936,N_10039,N_10000);
nand U11937 (N_11937,N_10777,N_10174);
and U11938 (N_11938,N_10384,N_10365);
and U11939 (N_11939,N_10604,N_10711);
nand U11940 (N_11940,N_10326,N_10760);
nand U11941 (N_11941,N_10932,N_10031);
nand U11942 (N_11942,N_10658,N_10530);
and U11943 (N_11943,N_10347,N_10350);
or U11944 (N_11944,N_10105,N_10811);
nor U11945 (N_11945,N_10162,N_10283);
xnor U11946 (N_11946,N_10440,N_10423);
nand U11947 (N_11947,N_10929,N_10984);
nand U11948 (N_11948,N_10307,N_10448);
and U11949 (N_11949,N_10465,N_10170);
or U11950 (N_11950,N_10447,N_10116);
and U11951 (N_11951,N_10235,N_10699);
nand U11952 (N_11952,N_10739,N_10628);
xor U11953 (N_11953,N_10432,N_10065);
and U11954 (N_11954,N_10720,N_10951);
nand U11955 (N_11955,N_10236,N_10234);
nor U11956 (N_11956,N_10970,N_10829);
and U11957 (N_11957,N_10310,N_10253);
xnor U11958 (N_11958,N_10855,N_10418);
nor U11959 (N_11959,N_10384,N_10198);
or U11960 (N_11960,N_10135,N_10768);
nand U11961 (N_11961,N_10381,N_10657);
and U11962 (N_11962,N_10550,N_10501);
or U11963 (N_11963,N_10833,N_10888);
and U11964 (N_11964,N_10538,N_10724);
nand U11965 (N_11965,N_10622,N_10455);
nor U11966 (N_11966,N_10429,N_10871);
nor U11967 (N_11967,N_10241,N_10048);
nor U11968 (N_11968,N_10726,N_10206);
xor U11969 (N_11969,N_10345,N_10481);
xnor U11970 (N_11970,N_10225,N_10078);
xnor U11971 (N_11971,N_10342,N_10890);
or U11972 (N_11972,N_10361,N_10160);
and U11973 (N_11973,N_10473,N_10990);
and U11974 (N_11974,N_10730,N_10961);
nor U11975 (N_11975,N_10877,N_10586);
xnor U11976 (N_11976,N_10482,N_10281);
or U11977 (N_11977,N_10956,N_10393);
xnor U11978 (N_11978,N_10810,N_10407);
xor U11979 (N_11979,N_10842,N_10804);
or U11980 (N_11980,N_10351,N_10745);
and U11981 (N_11981,N_10967,N_10656);
nand U11982 (N_11982,N_10270,N_10377);
and U11983 (N_11983,N_10359,N_10084);
nand U11984 (N_11984,N_10838,N_10928);
or U11985 (N_11985,N_10231,N_10250);
nor U11986 (N_11986,N_10097,N_10346);
nand U11987 (N_11987,N_10184,N_10284);
nor U11988 (N_11988,N_10464,N_10307);
xnor U11989 (N_11989,N_10978,N_10213);
and U11990 (N_11990,N_10709,N_10947);
and U11991 (N_11991,N_10798,N_10648);
nor U11992 (N_11992,N_10174,N_10902);
nand U11993 (N_11993,N_10790,N_10486);
nand U11994 (N_11994,N_10167,N_10558);
xor U11995 (N_11995,N_10132,N_10112);
nand U11996 (N_11996,N_10149,N_10667);
or U11997 (N_11997,N_10494,N_10095);
nand U11998 (N_11998,N_10210,N_10362);
xnor U11999 (N_11999,N_10670,N_10807);
xor U12000 (N_12000,N_11562,N_11905);
or U12001 (N_12001,N_11211,N_11785);
xor U12002 (N_12002,N_11838,N_11157);
and U12003 (N_12003,N_11930,N_11218);
xnor U12004 (N_12004,N_11715,N_11660);
nor U12005 (N_12005,N_11603,N_11226);
or U12006 (N_12006,N_11529,N_11279);
or U12007 (N_12007,N_11516,N_11429);
or U12008 (N_12008,N_11418,N_11917);
and U12009 (N_12009,N_11617,N_11551);
and U12010 (N_12010,N_11809,N_11553);
and U12011 (N_12011,N_11100,N_11408);
nand U12012 (N_12012,N_11171,N_11077);
nand U12013 (N_12013,N_11861,N_11445);
nor U12014 (N_12014,N_11751,N_11452);
or U12015 (N_12015,N_11354,N_11752);
nor U12016 (N_12016,N_11756,N_11963);
nand U12017 (N_12017,N_11256,N_11629);
nand U12018 (N_12018,N_11319,N_11244);
nand U12019 (N_12019,N_11866,N_11458);
and U12020 (N_12020,N_11833,N_11870);
or U12021 (N_12021,N_11827,N_11151);
or U12022 (N_12022,N_11823,N_11178);
nor U12023 (N_12023,N_11337,N_11273);
and U12024 (N_12024,N_11058,N_11806);
nand U12025 (N_12025,N_11851,N_11261);
xnor U12026 (N_12026,N_11667,N_11110);
or U12027 (N_12027,N_11788,N_11965);
and U12028 (N_12028,N_11060,N_11444);
or U12029 (N_12029,N_11493,N_11491);
xor U12030 (N_12030,N_11031,N_11441);
or U12031 (N_12031,N_11394,N_11257);
xnor U12032 (N_12032,N_11800,N_11313);
nor U12033 (N_12033,N_11084,N_11767);
nand U12034 (N_12034,N_11694,N_11766);
nand U12035 (N_12035,N_11947,N_11297);
nand U12036 (N_12036,N_11978,N_11545);
nand U12037 (N_12037,N_11386,N_11798);
nand U12038 (N_12038,N_11682,N_11604);
nor U12039 (N_12039,N_11001,N_11831);
and U12040 (N_12040,N_11489,N_11234);
and U12041 (N_12041,N_11461,N_11799);
or U12042 (N_12042,N_11816,N_11586);
nand U12043 (N_12043,N_11787,N_11263);
or U12044 (N_12044,N_11731,N_11690);
or U12045 (N_12045,N_11403,N_11236);
nand U12046 (N_12046,N_11262,N_11306);
and U12047 (N_12047,N_11534,N_11579);
nor U12048 (N_12048,N_11705,N_11755);
xor U12049 (N_12049,N_11958,N_11074);
and U12050 (N_12050,N_11185,N_11162);
nand U12051 (N_12051,N_11343,N_11713);
nand U12052 (N_12052,N_11083,N_11832);
or U12053 (N_12053,N_11710,N_11747);
nand U12054 (N_12054,N_11204,N_11375);
xor U12055 (N_12055,N_11164,N_11381);
nand U12056 (N_12056,N_11404,N_11672);
and U12057 (N_12057,N_11396,N_11335);
or U12058 (N_12058,N_11032,N_11321);
nand U12059 (N_12059,N_11049,N_11650);
nor U12060 (N_12060,N_11893,N_11775);
xnor U12061 (N_12061,N_11406,N_11305);
or U12062 (N_12062,N_11366,N_11307);
nand U12063 (N_12063,N_11535,N_11997);
or U12064 (N_12064,N_11308,N_11585);
and U12065 (N_12065,N_11665,N_11810);
and U12066 (N_12066,N_11248,N_11043);
or U12067 (N_12067,N_11777,N_11931);
or U12068 (N_12068,N_11186,N_11383);
and U12069 (N_12069,N_11175,N_11523);
nand U12070 (N_12070,N_11587,N_11447);
nor U12071 (N_12071,N_11134,N_11428);
xor U12072 (N_12072,N_11760,N_11974);
nand U12073 (N_12073,N_11150,N_11317);
nand U12074 (N_12074,N_11314,N_11829);
nand U12075 (N_12075,N_11808,N_11664);
xnor U12076 (N_12076,N_11129,N_11781);
nand U12077 (N_12077,N_11907,N_11653);
xor U12078 (N_12078,N_11764,N_11568);
nand U12079 (N_12079,N_11464,N_11599);
nand U12080 (N_12080,N_11388,N_11245);
nand U12081 (N_12081,N_11399,N_11901);
and U12082 (N_12082,N_11737,N_11675);
nor U12083 (N_12083,N_11413,N_11374);
nand U12084 (N_12084,N_11594,N_11888);
nand U12085 (N_12085,N_11423,N_11023);
nor U12086 (N_12086,N_11082,N_11143);
nor U12087 (N_12087,N_11841,N_11886);
xnor U12088 (N_12088,N_11221,N_11251);
xor U12089 (N_12089,N_11229,N_11814);
or U12090 (N_12090,N_11140,N_11050);
or U12091 (N_12091,N_11486,N_11398);
xnor U12092 (N_12092,N_11144,N_11584);
or U12093 (N_12093,N_11079,N_11385);
and U12094 (N_12094,N_11995,N_11472);
and U12095 (N_12095,N_11304,N_11509);
and U12096 (N_12096,N_11002,N_11910);
nor U12097 (N_12097,N_11582,N_11322);
xor U12098 (N_12098,N_11061,N_11651);
nand U12099 (N_12099,N_11911,N_11680);
nand U12100 (N_12100,N_11174,N_11260);
nor U12101 (N_12101,N_11889,N_11525);
xor U12102 (N_12102,N_11357,N_11044);
or U12103 (N_12103,N_11576,N_11719);
nor U12104 (N_12104,N_11591,N_11644);
and U12105 (N_12105,N_11819,N_11750);
nand U12106 (N_12106,N_11607,N_11853);
and U12107 (N_12107,N_11239,N_11674);
nand U12108 (N_12108,N_11108,N_11419);
or U12109 (N_12109,N_11287,N_11501);
nor U12110 (N_12110,N_11720,N_11700);
xor U12111 (N_12111,N_11479,N_11511);
and U12112 (N_12112,N_11902,N_11205);
xor U12113 (N_12113,N_11527,N_11985);
nand U12114 (N_12114,N_11272,N_11512);
xor U12115 (N_12115,N_11003,N_11506);
nand U12116 (N_12116,N_11432,N_11620);
or U12117 (N_12117,N_11361,N_11359);
or U12118 (N_12118,N_11820,N_11302);
xor U12119 (N_12119,N_11451,N_11275);
nor U12120 (N_12120,N_11064,N_11367);
nand U12121 (N_12121,N_11111,N_11513);
xor U12122 (N_12122,N_11497,N_11934);
and U12123 (N_12123,N_11789,N_11547);
nand U12124 (N_12124,N_11455,N_11540);
and U12125 (N_12125,N_11254,N_11805);
or U12126 (N_12126,N_11928,N_11906);
or U12127 (N_12127,N_11938,N_11740);
and U12128 (N_12128,N_11400,N_11633);
or U12129 (N_12129,N_11241,N_11711);
xnor U12130 (N_12130,N_11964,N_11492);
nor U12131 (N_12131,N_11727,N_11065);
or U12132 (N_12132,N_11015,N_11278);
or U12133 (N_12133,N_11242,N_11701);
and U12134 (N_12134,N_11167,N_11643);
xor U12135 (N_12135,N_11152,N_11608);
xor U12136 (N_12136,N_11942,N_11970);
nor U12137 (N_12137,N_11117,N_11703);
or U12138 (N_12138,N_11219,N_11372);
xor U12139 (N_12139,N_11133,N_11678);
nor U12140 (N_12140,N_11932,N_11474);
xnor U12141 (N_12141,N_11011,N_11939);
or U12142 (N_12142,N_11768,N_11336);
or U12143 (N_12143,N_11783,N_11807);
or U12144 (N_12144,N_11293,N_11858);
xnor U12145 (N_12145,N_11193,N_11648);
xor U12146 (N_12146,N_11803,N_11884);
and U12147 (N_12147,N_11087,N_11733);
nor U12148 (N_12148,N_11877,N_11225);
xor U12149 (N_12149,N_11860,N_11835);
xor U12150 (N_12150,N_11342,N_11093);
or U12151 (N_12151,N_11941,N_11796);
and U12152 (N_12152,N_11035,N_11548);
xor U12153 (N_12153,N_11228,N_11954);
nor U12154 (N_12154,N_11136,N_11786);
or U12155 (N_12155,N_11933,N_11704);
and U12156 (N_12156,N_11004,N_11330);
nor U12157 (N_12157,N_11736,N_11776);
and U12158 (N_12158,N_11341,N_11948);
and U12159 (N_12159,N_11887,N_11801);
and U12160 (N_12160,N_11190,N_11616);
or U12161 (N_12161,N_11131,N_11331);
or U12162 (N_12162,N_11602,N_11613);
nand U12163 (N_12163,N_11033,N_11303);
xnor U12164 (N_12164,N_11977,N_11334);
and U12165 (N_12165,N_11181,N_11988);
nand U12166 (N_12166,N_11687,N_11983);
and U12167 (N_12167,N_11908,N_11377);
nand U12168 (N_12168,N_11379,N_11748);
xor U12169 (N_12169,N_11056,N_11417);
nor U12170 (N_12170,N_11630,N_11161);
xnor U12171 (N_12171,N_11233,N_11846);
nor U12172 (N_12172,N_11580,N_11642);
nor U12173 (N_12173,N_11600,N_11348);
xnor U12174 (N_12174,N_11007,N_11344);
nand U12175 (N_12175,N_11916,N_11231);
nand U12176 (N_12176,N_11825,N_11109);
nor U12177 (N_12177,N_11728,N_11328);
or U12178 (N_12178,N_11338,N_11726);
nand U12179 (N_12179,N_11583,N_11096);
nand U12180 (N_12180,N_11188,N_11420);
and U12181 (N_12181,N_11826,N_11949);
or U12182 (N_12182,N_11757,N_11165);
xor U12183 (N_12183,N_11666,N_11876);
nand U12184 (N_12184,N_11252,N_11951);
nand U12185 (N_12185,N_11350,N_11378);
or U12186 (N_12186,N_11623,N_11349);
and U12187 (N_12187,N_11663,N_11542);
or U12188 (N_12188,N_11073,N_11029);
and U12189 (N_12189,N_11688,N_11495);
nor U12190 (N_12190,N_11010,N_11159);
xor U12191 (N_12191,N_11284,N_11890);
nand U12192 (N_12192,N_11924,N_11707);
nor U12193 (N_12193,N_11194,N_11734);
and U12194 (N_12194,N_11993,N_11518);
and U12195 (N_12195,N_11561,N_11067);
nor U12196 (N_12196,N_11972,N_11395);
and U12197 (N_12197,N_11026,N_11119);
xor U12198 (N_12198,N_11028,N_11609);
nand U12199 (N_12199,N_11191,N_11494);
xor U12200 (N_12200,N_11255,N_11327);
nand U12201 (N_12201,N_11173,N_11196);
nand U12202 (N_12202,N_11697,N_11968);
nand U12203 (N_12203,N_11480,N_11457);
nand U12204 (N_12204,N_11891,N_11462);
and U12205 (N_12205,N_11201,N_11019);
nor U12206 (N_12206,N_11006,N_11612);
and U12207 (N_12207,N_11309,N_11828);
nand U12208 (N_12208,N_11448,N_11325);
nand U12209 (N_12209,N_11515,N_11048);
and U12210 (N_12210,N_11440,N_11944);
nor U12211 (N_12211,N_11316,N_11095);
or U12212 (N_12212,N_11224,N_11869);
and U12213 (N_12213,N_11559,N_11619);
xnor U12214 (N_12214,N_11596,N_11363);
nor U12215 (N_12215,N_11976,N_11635);
and U12216 (N_12216,N_11097,N_11209);
nand U12217 (N_12217,N_11546,N_11759);
nor U12218 (N_12218,N_11681,N_11268);
nand U12219 (N_12219,N_11955,N_11702);
nand U12220 (N_12220,N_11957,N_11892);
or U12221 (N_12221,N_11923,N_11519);
nand U12222 (N_12222,N_11645,N_11282);
and U12223 (N_12223,N_11470,N_11514);
nand U12224 (N_12224,N_11856,N_11104);
xor U12225 (N_12225,N_11961,N_11863);
and U12226 (N_12226,N_11691,N_11160);
xnor U12227 (N_12227,N_11054,N_11679);
nand U12228 (N_12228,N_11311,N_11742);
and U12229 (N_12229,N_11299,N_11634);
xor U12230 (N_12230,N_11145,N_11230);
xor U12231 (N_12231,N_11431,N_11821);
nand U12232 (N_12232,N_11744,N_11926);
or U12233 (N_12233,N_11848,N_11802);
or U12234 (N_12234,N_11882,N_11574);
nor U12235 (N_12235,N_11318,N_11564);
nor U12236 (N_12236,N_11971,N_11956);
or U12237 (N_12237,N_11724,N_11477);
or U12238 (N_12238,N_11427,N_11389);
and U12239 (N_12239,N_11765,N_11125);
and U12240 (N_12240,N_11824,N_11240);
and U12241 (N_12241,N_11391,N_11794);
or U12242 (N_12242,N_11692,N_11871);
and U12243 (N_12243,N_11370,N_11080);
and U12244 (N_12244,N_11270,N_11088);
nor U12245 (N_12245,N_11078,N_11855);
xnor U12246 (N_12246,N_11723,N_11771);
nand U12247 (N_12247,N_11132,N_11469);
xnor U12248 (N_12248,N_11792,N_11536);
and U12249 (N_12249,N_11661,N_11845);
xnor U12250 (N_12250,N_11929,N_11034);
and U12251 (N_12251,N_11137,N_11722);
or U12252 (N_12252,N_11927,N_11880);
nand U12253 (N_12253,N_11543,N_11421);
xnor U12254 (N_12254,N_11000,N_11813);
nor U12255 (N_12255,N_11281,N_11639);
and U12256 (N_12256,N_11655,N_11184);
xnor U12257 (N_12257,N_11605,N_11994);
and U12258 (N_12258,N_11528,N_11405);
xnor U12259 (N_12259,N_11286,N_11741);
nor U12260 (N_12260,N_11089,N_11038);
nand U12261 (N_12261,N_11091,N_11166);
or U12262 (N_12262,N_11463,N_11356);
nor U12263 (N_12263,N_11524,N_11991);
nor U12264 (N_12264,N_11062,N_11358);
nand U12265 (N_12265,N_11761,N_11641);
or U12266 (N_12266,N_11659,N_11817);
xnor U12267 (N_12267,N_11123,N_11267);
nand U12268 (N_12268,N_11039,N_11005);
nand U12269 (N_12269,N_11854,N_11502);
and U12270 (N_12270,N_11059,N_11818);
nor U12271 (N_12271,N_11510,N_11392);
nor U12272 (N_12272,N_11153,N_11735);
nand U12273 (N_12273,N_11793,N_11867);
nor U12274 (N_12274,N_11565,N_11790);
or U12275 (N_12275,N_11042,N_11481);
and U12276 (N_12276,N_11081,N_11778);
and U12277 (N_12277,N_11769,N_11120);
xnor U12278 (N_12278,N_11671,N_11259);
nor U12279 (N_12279,N_11412,N_11537);
and U12280 (N_12280,N_11683,N_11291);
nor U12281 (N_12281,N_11076,N_11371);
nor U12282 (N_12282,N_11124,N_11557);
xnor U12283 (N_12283,N_11149,N_11990);
nand U12284 (N_12284,N_11217,N_11158);
nor U12285 (N_12285,N_11857,N_11085);
or U12286 (N_12286,N_11333,N_11182);
and U12287 (N_12287,N_11830,N_11782);
nand U12288 (N_12288,N_11589,N_11323);
nand U12289 (N_12289,N_11953,N_11677);
xor U12290 (N_12290,N_11895,N_11436);
nand U12291 (N_12291,N_11266,N_11066);
or U12292 (N_12292,N_11521,N_11758);
nor U12293 (N_12293,N_11207,N_11689);
nor U12294 (N_12294,N_11555,N_11092);
and U12295 (N_12295,N_11069,N_11453);
nand U12296 (N_12296,N_11285,N_11936);
or U12297 (N_12297,N_11714,N_11116);
xor U12298 (N_12298,N_11815,N_11626);
nand U12299 (N_12299,N_11347,N_11393);
and U12300 (N_12300,N_11146,N_11496);
xnor U12301 (N_12301,N_11770,N_11187);
xnor U12302 (N_12302,N_11526,N_11364);
or U12303 (N_12303,N_11189,N_11113);
xnor U12304 (N_12304,N_11484,N_11987);
or U12305 (N_12305,N_11315,N_11433);
xor U12306 (N_12306,N_11490,N_11873);
and U12307 (N_12307,N_11558,N_11141);
and U12308 (N_12308,N_11025,N_11746);
or U12309 (N_12309,N_11578,N_11365);
xnor U12310 (N_12310,N_11590,N_11549);
and U12311 (N_12311,N_11435,N_11552);
nand U12312 (N_12312,N_11220,N_11312);
and U12313 (N_12313,N_11508,N_11581);
or U12314 (N_12314,N_11142,N_11696);
xor U12315 (N_12315,N_11914,N_11407);
nor U12316 (N_12316,N_11718,N_11258);
nand U12317 (N_12317,N_11637,N_11169);
and U12318 (N_12318,N_11631,N_11105);
nor U12319 (N_12319,N_11601,N_11246);
nor U12320 (N_12320,N_11402,N_11121);
nor U12321 (N_12321,N_11271,N_11449);
and U12322 (N_12322,N_11657,N_11872);
xnor U12323 (N_12323,N_11532,N_11176);
or U12324 (N_12324,N_11898,N_11439);
nor U12325 (N_12325,N_11979,N_11301);
xor U12326 (N_12326,N_11847,N_11446);
and U12327 (N_12327,N_11966,N_11739);
or U12328 (N_12328,N_11772,N_11530);
and U12329 (N_12329,N_11422,N_11541);
xor U12330 (N_12330,N_11288,N_11454);
and U12331 (N_12331,N_11022,N_11852);
nand U12332 (N_12332,N_11868,N_11018);
and U12333 (N_12333,N_11126,N_11476);
nand U12334 (N_12334,N_11636,N_11068);
nor U12335 (N_12335,N_11183,N_11329);
nand U12336 (N_12336,N_11415,N_11897);
nor U12337 (N_12337,N_11397,N_11243);
nand U12338 (N_12338,N_11570,N_11249);
or U12339 (N_12339,N_11738,N_11465);
and U12340 (N_12340,N_11622,N_11409);
nand U12341 (N_12341,N_11215,N_11036);
or U12342 (N_12342,N_11216,N_11982);
xnor U12343 (N_12343,N_11883,N_11483);
nand U12344 (N_12344,N_11300,N_11382);
nand U12345 (N_12345,N_11717,N_11203);
xnor U12346 (N_12346,N_11811,N_11981);
and U12347 (N_12347,N_11984,N_11139);
nand U12348 (N_12348,N_11904,N_11859);
and U12349 (N_12349,N_11352,N_11638);
or U12350 (N_12350,N_11763,N_11684);
and U12351 (N_12351,N_11045,N_11780);
nand U12352 (N_12352,N_11416,N_11206);
nand U12353 (N_12353,N_11567,N_11471);
or U12354 (N_12354,N_11712,N_11430);
and U12355 (N_12355,N_11037,N_11875);
xnor U12356 (N_12356,N_11959,N_11114);
xor U12357 (N_12357,N_11573,N_11843);
and U12358 (N_12358,N_11560,N_11920);
and U12359 (N_12359,N_11885,N_11269);
xor U12360 (N_12360,N_11369,N_11588);
and U12361 (N_12361,N_11615,N_11122);
nor U12362 (N_12362,N_11238,N_11339);
and U12363 (N_12363,N_11292,N_11373);
and U12364 (N_12364,N_11592,N_11012);
nand U12365 (N_12365,N_11130,N_11438);
and U12366 (N_12366,N_11232,N_11921);
and U12367 (N_12367,N_11686,N_11102);
nand U12368 (N_12368,N_11414,N_11086);
xnor U12369 (N_12369,N_11063,N_11909);
nor U12370 (N_12370,N_11380,N_11695);
or U12371 (N_12371,N_11346,N_11214);
or U12372 (N_12372,N_11879,N_11784);
xnor U12373 (N_12373,N_11708,N_11253);
xnor U12374 (N_12374,N_11384,N_11053);
xor U12375 (N_12375,N_11024,N_11566);
xor U12376 (N_12376,N_11101,N_11155);
xnor U12377 (N_12377,N_11355,N_11345);
nand U12378 (N_12378,N_11351,N_11522);
and U12379 (N_12379,N_11554,N_11625);
nor U12380 (N_12380,N_11274,N_11989);
nor U12381 (N_12381,N_11544,N_11670);
xor U12382 (N_12382,N_11969,N_11721);
or U12383 (N_12383,N_11202,N_11112);
and U12384 (N_12384,N_11047,N_11676);
nand U12385 (N_12385,N_11698,N_11999);
xnor U12386 (N_12386,N_11839,N_11646);
nor U12387 (N_12387,N_11467,N_11915);
or U12388 (N_12388,N_11569,N_11919);
or U12389 (N_12389,N_11410,N_11353);
nand U12390 (N_12390,N_11652,N_11894);
nand U12391 (N_12391,N_11265,N_11837);
nor U12392 (N_12392,N_11170,N_11745);
or U12393 (N_12393,N_11498,N_11289);
or U12394 (N_12394,N_11070,N_11992);
nor U12395 (N_12395,N_11030,N_11250);
and U12396 (N_12396,N_11390,N_11055);
and U12397 (N_12397,N_11450,N_11235);
or U12398 (N_12398,N_11135,N_11795);
or U12399 (N_12399,N_11147,N_11693);
and U12400 (N_12400,N_11197,N_11709);
and U12401 (N_12401,N_11531,N_11975);
nor U12402 (N_12402,N_11836,N_11550);
nand U12403 (N_12403,N_11918,N_11654);
and U12404 (N_12404,N_11980,N_11326);
xor U12405 (N_12405,N_11621,N_11115);
and U12406 (N_12406,N_11812,N_11387);
xor U12407 (N_12407,N_11099,N_11725);
nand U12408 (N_12408,N_11168,N_11940);
and U12409 (N_12409,N_11503,N_11401);
xor U12410 (N_12410,N_11656,N_11276);
nand U12411 (N_12411,N_11842,N_11459);
and U12412 (N_12412,N_11294,N_11647);
and U12413 (N_12413,N_11849,N_11172);
or U12414 (N_12414,N_11706,N_11107);
xor U12415 (N_12415,N_11822,N_11685);
nor U12416 (N_12416,N_11075,N_11505);
nor U12417 (N_12417,N_11632,N_11195);
nor U12418 (N_12418,N_11426,N_11797);
and U12419 (N_12419,N_11507,N_11618);
and U12420 (N_12420,N_11208,N_11013);
nand U12421 (N_12421,N_11485,N_11952);
and U12422 (N_12422,N_11499,N_11850);
nor U12423 (N_12423,N_11874,N_11669);
nand U12424 (N_12424,N_11922,N_11699);
nor U12425 (N_12425,N_11340,N_11290);
or U12426 (N_12426,N_11791,N_11051);
nand U12427 (N_12427,N_11606,N_11106);
or U12428 (N_12428,N_11227,N_11027);
nor U12429 (N_12429,N_11071,N_11572);
nor U12430 (N_12430,N_11016,N_11320);
or U12431 (N_12431,N_11732,N_11324);
or U12432 (N_12432,N_11624,N_11598);
xor U12433 (N_12433,N_11310,N_11774);
nor U12434 (N_12434,N_11017,N_11834);
or U12435 (N_12435,N_11743,N_11881);
xor U12436 (N_12436,N_11094,N_11437);
nor U12437 (N_12437,N_11154,N_11864);
or U12438 (N_12438,N_11473,N_11640);
nor U12439 (N_12439,N_11804,N_11500);
and U12440 (N_12440,N_11593,N_11199);
nor U12441 (N_12441,N_11996,N_11716);
nor U12442 (N_12442,N_11899,N_11237);
nor U12443 (N_12443,N_11180,N_11468);
xnor U12444 (N_12444,N_11280,N_11950);
xor U12445 (N_12445,N_11945,N_11138);
or U12446 (N_12446,N_11376,N_11434);
or U12447 (N_12447,N_11729,N_11614);
or U12448 (N_12448,N_11040,N_11925);
xnor U12449 (N_12449,N_11103,N_11556);
nand U12450 (N_12450,N_11962,N_11753);
and U12451 (N_12451,N_11862,N_11475);
nand U12452 (N_12452,N_11442,N_11960);
nor U12453 (N_12453,N_11443,N_11021);
and U12454 (N_12454,N_11896,N_11460);
xor U12455 (N_12455,N_11673,N_11563);
and U12456 (N_12456,N_11192,N_11538);
or U12457 (N_12457,N_11840,N_11487);
nor U12458 (N_12458,N_11967,N_11425);
xnor U12459 (N_12459,N_11730,N_11627);
and U12460 (N_12460,N_11118,N_11520);
and U12461 (N_12461,N_11986,N_11998);
nand U12462 (N_12462,N_11912,N_11773);
and U12463 (N_12463,N_11946,N_11179);
xor U12464 (N_12464,N_11128,N_11935);
or U12465 (N_12465,N_11210,N_11296);
or U12466 (N_12466,N_11456,N_11779);
nand U12467 (N_12467,N_11865,N_11098);
nor U12468 (N_12468,N_11575,N_11277);
xnor U12469 (N_12469,N_11668,N_11482);
nand U12470 (N_12470,N_11900,N_11571);
nand U12471 (N_12471,N_11488,N_11424);
and U12472 (N_12472,N_11212,N_11163);
and U12473 (N_12473,N_11020,N_11628);
nand U12474 (N_12474,N_11148,N_11878);
nand U12475 (N_12475,N_11213,N_11973);
nor U12476 (N_12476,N_11283,N_11200);
or U12477 (N_12477,N_11466,N_11595);
nor U12478 (N_12478,N_11247,N_11072);
nand U12479 (N_12479,N_11844,N_11662);
nor U12480 (N_12480,N_11610,N_11222);
nor U12481 (N_12481,N_11943,N_11597);
or U12482 (N_12482,N_11295,N_11362);
xnor U12483 (N_12483,N_11223,N_11298);
nand U12484 (N_12484,N_11156,N_11903);
xnor U12485 (N_12485,N_11008,N_11014);
nor U12486 (N_12486,N_11264,N_11090);
and U12487 (N_12487,N_11577,N_11127);
or U12488 (N_12488,N_11332,N_11913);
nand U12489 (N_12489,N_11749,N_11539);
nand U12490 (N_12490,N_11009,N_11041);
or U12491 (N_12491,N_11360,N_11052);
or U12492 (N_12492,N_11198,N_11754);
or U12493 (N_12493,N_11478,N_11368);
xor U12494 (N_12494,N_11649,N_11611);
or U12495 (N_12495,N_11517,N_11177);
nor U12496 (N_12496,N_11057,N_11411);
nor U12497 (N_12497,N_11504,N_11762);
xor U12498 (N_12498,N_11533,N_11658);
or U12499 (N_12499,N_11046,N_11937);
and U12500 (N_12500,N_11608,N_11819);
or U12501 (N_12501,N_11424,N_11400);
nand U12502 (N_12502,N_11961,N_11075);
and U12503 (N_12503,N_11883,N_11930);
or U12504 (N_12504,N_11294,N_11982);
nand U12505 (N_12505,N_11043,N_11655);
xnor U12506 (N_12506,N_11503,N_11894);
or U12507 (N_12507,N_11375,N_11685);
nor U12508 (N_12508,N_11733,N_11683);
and U12509 (N_12509,N_11229,N_11244);
xor U12510 (N_12510,N_11820,N_11646);
and U12511 (N_12511,N_11435,N_11945);
or U12512 (N_12512,N_11553,N_11242);
and U12513 (N_12513,N_11503,N_11861);
nand U12514 (N_12514,N_11226,N_11327);
nand U12515 (N_12515,N_11904,N_11381);
or U12516 (N_12516,N_11487,N_11238);
xnor U12517 (N_12517,N_11786,N_11721);
and U12518 (N_12518,N_11307,N_11689);
nor U12519 (N_12519,N_11540,N_11401);
nor U12520 (N_12520,N_11236,N_11624);
nand U12521 (N_12521,N_11569,N_11698);
nand U12522 (N_12522,N_11719,N_11750);
xor U12523 (N_12523,N_11454,N_11057);
or U12524 (N_12524,N_11053,N_11276);
nand U12525 (N_12525,N_11519,N_11555);
nor U12526 (N_12526,N_11054,N_11222);
nor U12527 (N_12527,N_11089,N_11021);
nand U12528 (N_12528,N_11605,N_11049);
and U12529 (N_12529,N_11741,N_11990);
nand U12530 (N_12530,N_11127,N_11491);
or U12531 (N_12531,N_11752,N_11255);
nor U12532 (N_12532,N_11317,N_11882);
nor U12533 (N_12533,N_11361,N_11871);
nor U12534 (N_12534,N_11355,N_11145);
or U12535 (N_12535,N_11282,N_11734);
xnor U12536 (N_12536,N_11295,N_11686);
nand U12537 (N_12537,N_11444,N_11932);
and U12538 (N_12538,N_11968,N_11822);
xnor U12539 (N_12539,N_11674,N_11959);
nand U12540 (N_12540,N_11583,N_11087);
or U12541 (N_12541,N_11453,N_11454);
xor U12542 (N_12542,N_11180,N_11793);
nor U12543 (N_12543,N_11061,N_11367);
nor U12544 (N_12544,N_11603,N_11147);
nand U12545 (N_12545,N_11132,N_11276);
nand U12546 (N_12546,N_11885,N_11198);
or U12547 (N_12547,N_11396,N_11267);
or U12548 (N_12548,N_11518,N_11435);
xnor U12549 (N_12549,N_11415,N_11202);
nand U12550 (N_12550,N_11546,N_11920);
or U12551 (N_12551,N_11239,N_11262);
xor U12552 (N_12552,N_11276,N_11187);
xor U12553 (N_12553,N_11990,N_11693);
nand U12554 (N_12554,N_11717,N_11781);
xor U12555 (N_12555,N_11549,N_11142);
or U12556 (N_12556,N_11115,N_11597);
nor U12557 (N_12557,N_11255,N_11893);
nor U12558 (N_12558,N_11882,N_11524);
nand U12559 (N_12559,N_11782,N_11502);
nor U12560 (N_12560,N_11153,N_11530);
or U12561 (N_12561,N_11037,N_11131);
and U12562 (N_12562,N_11998,N_11164);
xor U12563 (N_12563,N_11520,N_11434);
xor U12564 (N_12564,N_11900,N_11771);
and U12565 (N_12565,N_11590,N_11544);
or U12566 (N_12566,N_11028,N_11530);
or U12567 (N_12567,N_11248,N_11333);
nand U12568 (N_12568,N_11223,N_11447);
nand U12569 (N_12569,N_11914,N_11755);
nand U12570 (N_12570,N_11330,N_11447);
nor U12571 (N_12571,N_11189,N_11765);
and U12572 (N_12572,N_11466,N_11088);
or U12573 (N_12573,N_11359,N_11895);
xor U12574 (N_12574,N_11884,N_11931);
or U12575 (N_12575,N_11620,N_11961);
nand U12576 (N_12576,N_11106,N_11511);
and U12577 (N_12577,N_11848,N_11604);
nor U12578 (N_12578,N_11626,N_11678);
xnor U12579 (N_12579,N_11909,N_11126);
and U12580 (N_12580,N_11624,N_11693);
or U12581 (N_12581,N_11179,N_11061);
xor U12582 (N_12582,N_11289,N_11778);
nor U12583 (N_12583,N_11846,N_11647);
nor U12584 (N_12584,N_11102,N_11050);
or U12585 (N_12585,N_11155,N_11760);
xor U12586 (N_12586,N_11584,N_11449);
nand U12587 (N_12587,N_11931,N_11182);
xnor U12588 (N_12588,N_11100,N_11976);
nor U12589 (N_12589,N_11480,N_11437);
nor U12590 (N_12590,N_11626,N_11484);
nor U12591 (N_12591,N_11671,N_11150);
and U12592 (N_12592,N_11562,N_11891);
nor U12593 (N_12593,N_11053,N_11046);
nor U12594 (N_12594,N_11057,N_11402);
or U12595 (N_12595,N_11151,N_11770);
nor U12596 (N_12596,N_11544,N_11826);
xnor U12597 (N_12597,N_11029,N_11002);
or U12598 (N_12598,N_11555,N_11039);
and U12599 (N_12599,N_11389,N_11334);
nor U12600 (N_12600,N_11728,N_11517);
and U12601 (N_12601,N_11344,N_11059);
xnor U12602 (N_12602,N_11780,N_11696);
or U12603 (N_12603,N_11717,N_11570);
xor U12604 (N_12604,N_11034,N_11580);
and U12605 (N_12605,N_11315,N_11650);
nand U12606 (N_12606,N_11710,N_11656);
nor U12607 (N_12607,N_11939,N_11631);
nor U12608 (N_12608,N_11023,N_11884);
xnor U12609 (N_12609,N_11449,N_11643);
nor U12610 (N_12610,N_11040,N_11973);
or U12611 (N_12611,N_11486,N_11134);
xnor U12612 (N_12612,N_11125,N_11907);
nand U12613 (N_12613,N_11518,N_11054);
and U12614 (N_12614,N_11333,N_11448);
or U12615 (N_12615,N_11830,N_11289);
and U12616 (N_12616,N_11780,N_11370);
xor U12617 (N_12617,N_11909,N_11417);
or U12618 (N_12618,N_11805,N_11887);
nor U12619 (N_12619,N_11222,N_11311);
nand U12620 (N_12620,N_11513,N_11569);
nand U12621 (N_12621,N_11719,N_11138);
and U12622 (N_12622,N_11333,N_11446);
xnor U12623 (N_12623,N_11922,N_11178);
xnor U12624 (N_12624,N_11145,N_11835);
and U12625 (N_12625,N_11017,N_11751);
nand U12626 (N_12626,N_11381,N_11147);
nor U12627 (N_12627,N_11126,N_11489);
xor U12628 (N_12628,N_11767,N_11418);
nand U12629 (N_12629,N_11612,N_11449);
and U12630 (N_12630,N_11383,N_11755);
or U12631 (N_12631,N_11527,N_11201);
nand U12632 (N_12632,N_11146,N_11453);
or U12633 (N_12633,N_11659,N_11194);
or U12634 (N_12634,N_11143,N_11102);
nand U12635 (N_12635,N_11404,N_11889);
or U12636 (N_12636,N_11580,N_11085);
nor U12637 (N_12637,N_11669,N_11412);
nand U12638 (N_12638,N_11317,N_11681);
nand U12639 (N_12639,N_11422,N_11037);
nand U12640 (N_12640,N_11606,N_11178);
nor U12641 (N_12641,N_11223,N_11088);
and U12642 (N_12642,N_11058,N_11322);
or U12643 (N_12643,N_11273,N_11360);
and U12644 (N_12644,N_11022,N_11194);
xnor U12645 (N_12645,N_11868,N_11948);
or U12646 (N_12646,N_11630,N_11830);
nor U12647 (N_12647,N_11464,N_11395);
or U12648 (N_12648,N_11160,N_11856);
nor U12649 (N_12649,N_11651,N_11871);
xor U12650 (N_12650,N_11887,N_11051);
nor U12651 (N_12651,N_11176,N_11704);
nor U12652 (N_12652,N_11832,N_11683);
nor U12653 (N_12653,N_11283,N_11994);
and U12654 (N_12654,N_11650,N_11545);
and U12655 (N_12655,N_11987,N_11251);
xor U12656 (N_12656,N_11083,N_11575);
or U12657 (N_12657,N_11174,N_11888);
or U12658 (N_12658,N_11789,N_11231);
xor U12659 (N_12659,N_11236,N_11555);
xor U12660 (N_12660,N_11086,N_11698);
nand U12661 (N_12661,N_11723,N_11151);
or U12662 (N_12662,N_11864,N_11420);
and U12663 (N_12663,N_11239,N_11066);
nor U12664 (N_12664,N_11494,N_11281);
nor U12665 (N_12665,N_11416,N_11303);
xnor U12666 (N_12666,N_11007,N_11849);
nor U12667 (N_12667,N_11416,N_11179);
xnor U12668 (N_12668,N_11303,N_11104);
and U12669 (N_12669,N_11953,N_11440);
nand U12670 (N_12670,N_11875,N_11126);
nand U12671 (N_12671,N_11659,N_11961);
and U12672 (N_12672,N_11282,N_11833);
nand U12673 (N_12673,N_11991,N_11597);
or U12674 (N_12674,N_11908,N_11616);
nand U12675 (N_12675,N_11931,N_11960);
nor U12676 (N_12676,N_11243,N_11429);
nand U12677 (N_12677,N_11938,N_11319);
nand U12678 (N_12678,N_11430,N_11271);
or U12679 (N_12679,N_11074,N_11862);
and U12680 (N_12680,N_11249,N_11288);
and U12681 (N_12681,N_11934,N_11804);
xor U12682 (N_12682,N_11836,N_11028);
xnor U12683 (N_12683,N_11501,N_11529);
nor U12684 (N_12684,N_11628,N_11739);
and U12685 (N_12685,N_11211,N_11088);
and U12686 (N_12686,N_11947,N_11969);
xor U12687 (N_12687,N_11925,N_11710);
and U12688 (N_12688,N_11506,N_11186);
xor U12689 (N_12689,N_11132,N_11902);
or U12690 (N_12690,N_11266,N_11295);
or U12691 (N_12691,N_11761,N_11123);
nor U12692 (N_12692,N_11280,N_11295);
nand U12693 (N_12693,N_11379,N_11394);
xnor U12694 (N_12694,N_11572,N_11574);
nand U12695 (N_12695,N_11292,N_11182);
nor U12696 (N_12696,N_11334,N_11833);
xor U12697 (N_12697,N_11778,N_11820);
or U12698 (N_12698,N_11745,N_11132);
or U12699 (N_12699,N_11178,N_11147);
xor U12700 (N_12700,N_11223,N_11945);
nor U12701 (N_12701,N_11014,N_11716);
and U12702 (N_12702,N_11217,N_11353);
nor U12703 (N_12703,N_11721,N_11057);
xnor U12704 (N_12704,N_11147,N_11239);
nor U12705 (N_12705,N_11669,N_11424);
xor U12706 (N_12706,N_11547,N_11643);
nor U12707 (N_12707,N_11227,N_11811);
nand U12708 (N_12708,N_11383,N_11704);
or U12709 (N_12709,N_11654,N_11060);
xor U12710 (N_12710,N_11620,N_11754);
nor U12711 (N_12711,N_11888,N_11772);
xnor U12712 (N_12712,N_11638,N_11771);
nand U12713 (N_12713,N_11990,N_11142);
or U12714 (N_12714,N_11399,N_11101);
nor U12715 (N_12715,N_11970,N_11735);
and U12716 (N_12716,N_11500,N_11245);
nand U12717 (N_12717,N_11267,N_11811);
or U12718 (N_12718,N_11750,N_11006);
xor U12719 (N_12719,N_11776,N_11108);
nor U12720 (N_12720,N_11369,N_11158);
xnor U12721 (N_12721,N_11696,N_11281);
nand U12722 (N_12722,N_11754,N_11517);
or U12723 (N_12723,N_11538,N_11957);
nor U12724 (N_12724,N_11673,N_11662);
or U12725 (N_12725,N_11886,N_11734);
nor U12726 (N_12726,N_11607,N_11940);
or U12727 (N_12727,N_11339,N_11751);
and U12728 (N_12728,N_11564,N_11860);
and U12729 (N_12729,N_11496,N_11940);
xnor U12730 (N_12730,N_11526,N_11889);
and U12731 (N_12731,N_11084,N_11985);
or U12732 (N_12732,N_11783,N_11879);
nand U12733 (N_12733,N_11193,N_11506);
nand U12734 (N_12734,N_11602,N_11441);
xor U12735 (N_12735,N_11487,N_11403);
nand U12736 (N_12736,N_11262,N_11060);
and U12737 (N_12737,N_11735,N_11479);
or U12738 (N_12738,N_11877,N_11669);
xor U12739 (N_12739,N_11309,N_11369);
or U12740 (N_12740,N_11985,N_11591);
or U12741 (N_12741,N_11420,N_11490);
nor U12742 (N_12742,N_11705,N_11679);
xnor U12743 (N_12743,N_11639,N_11153);
or U12744 (N_12744,N_11445,N_11737);
xnor U12745 (N_12745,N_11593,N_11003);
xnor U12746 (N_12746,N_11504,N_11075);
nand U12747 (N_12747,N_11928,N_11456);
nand U12748 (N_12748,N_11430,N_11954);
or U12749 (N_12749,N_11023,N_11900);
nand U12750 (N_12750,N_11603,N_11491);
and U12751 (N_12751,N_11694,N_11777);
nand U12752 (N_12752,N_11880,N_11896);
or U12753 (N_12753,N_11391,N_11278);
or U12754 (N_12754,N_11746,N_11781);
nand U12755 (N_12755,N_11646,N_11906);
nand U12756 (N_12756,N_11850,N_11208);
xor U12757 (N_12757,N_11357,N_11320);
and U12758 (N_12758,N_11564,N_11057);
or U12759 (N_12759,N_11049,N_11527);
nor U12760 (N_12760,N_11894,N_11068);
nor U12761 (N_12761,N_11227,N_11859);
or U12762 (N_12762,N_11780,N_11707);
or U12763 (N_12763,N_11379,N_11112);
and U12764 (N_12764,N_11229,N_11252);
nor U12765 (N_12765,N_11855,N_11900);
nor U12766 (N_12766,N_11706,N_11336);
and U12767 (N_12767,N_11556,N_11454);
nor U12768 (N_12768,N_11927,N_11513);
nand U12769 (N_12769,N_11551,N_11910);
and U12770 (N_12770,N_11578,N_11425);
nand U12771 (N_12771,N_11277,N_11187);
nor U12772 (N_12772,N_11191,N_11295);
nand U12773 (N_12773,N_11803,N_11173);
or U12774 (N_12774,N_11991,N_11204);
or U12775 (N_12775,N_11267,N_11759);
xnor U12776 (N_12776,N_11757,N_11577);
xnor U12777 (N_12777,N_11620,N_11798);
nor U12778 (N_12778,N_11413,N_11937);
or U12779 (N_12779,N_11600,N_11615);
xor U12780 (N_12780,N_11372,N_11963);
nor U12781 (N_12781,N_11756,N_11527);
or U12782 (N_12782,N_11331,N_11168);
nor U12783 (N_12783,N_11976,N_11775);
xnor U12784 (N_12784,N_11925,N_11757);
nor U12785 (N_12785,N_11852,N_11816);
nor U12786 (N_12786,N_11447,N_11663);
xnor U12787 (N_12787,N_11677,N_11053);
or U12788 (N_12788,N_11322,N_11335);
nor U12789 (N_12789,N_11941,N_11904);
xnor U12790 (N_12790,N_11603,N_11285);
nor U12791 (N_12791,N_11523,N_11127);
nand U12792 (N_12792,N_11817,N_11121);
or U12793 (N_12793,N_11116,N_11898);
xor U12794 (N_12794,N_11008,N_11761);
nor U12795 (N_12795,N_11546,N_11285);
and U12796 (N_12796,N_11327,N_11755);
or U12797 (N_12797,N_11193,N_11195);
xor U12798 (N_12798,N_11249,N_11669);
nor U12799 (N_12799,N_11363,N_11794);
nor U12800 (N_12800,N_11545,N_11938);
or U12801 (N_12801,N_11762,N_11653);
xnor U12802 (N_12802,N_11701,N_11279);
xnor U12803 (N_12803,N_11234,N_11688);
xor U12804 (N_12804,N_11135,N_11661);
or U12805 (N_12805,N_11555,N_11495);
or U12806 (N_12806,N_11905,N_11020);
and U12807 (N_12807,N_11643,N_11455);
or U12808 (N_12808,N_11060,N_11473);
and U12809 (N_12809,N_11953,N_11260);
xor U12810 (N_12810,N_11561,N_11718);
xnor U12811 (N_12811,N_11718,N_11283);
and U12812 (N_12812,N_11193,N_11733);
or U12813 (N_12813,N_11886,N_11079);
and U12814 (N_12814,N_11505,N_11787);
and U12815 (N_12815,N_11236,N_11832);
or U12816 (N_12816,N_11610,N_11531);
xnor U12817 (N_12817,N_11109,N_11858);
nand U12818 (N_12818,N_11337,N_11535);
nor U12819 (N_12819,N_11180,N_11839);
xor U12820 (N_12820,N_11807,N_11248);
nor U12821 (N_12821,N_11029,N_11740);
and U12822 (N_12822,N_11807,N_11423);
nor U12823 (N_12823,N_11862,N_11047);
or U12824 (N_12824,N_11316,N_11525);
xnor U12825 (N_12825,N_11264,N_11971);
xnor U12826 (N_12826,N_11479,N_11397);
xor U12827 (N_12827,N_11264,N_11695);
and U12828 (N_12828,N_11429,N_11044);
nand U12829 (N_12829,N_11995,N_11600);
nand U12830 (N_12830,N_11753,N_11328);
nand U12831 (N_12831,N_11179,N_11690);
or U12832 (N_12832,N_11954,N_11054);
nand U12833 (N_12833,N_11211,N_11306);
xor U12834 (N_12834,N_11529,N_11342);
and U12835 (N_12835,N_11461,N_11243);
nand U12836 (N_12836,N_11929,N_11269);
and U12837 (N_12837,N_11715,N_11173);
xor U12838 (N_12838,N_11100,N_11450);
nand U12839 (N_12839,N_11951,N_11702);
nor U12840 (N_12840,N_11916,N_11473);
and U12841 (N_12841,N_11355,N_11973);
xor U12842 (N_12842,N_11255,N_11940);
and U12843 (N_12843,N_11541,N_11494);
and U12844 (N_12844,N_11110,N_11483);
or U12845 (N_12845,N_11585,N_11456);
xor U12846 (N_12846,N_11393,N_11597);
or U12847 (N_12847,N_11396,N_11351);
nand U12848 (N_12848,N_11299,N_11666);
or U12849 (N_12849,N_11388,N_11719);
and U12850 (N_12850,N_11004,N_11386);
and U12851 (N_12851,N_11664,N_11496);
nand U12852 (N_12852,N_11874,N_11479);
nor U12853 (N_12853,N_11888,N_11562);
and U12854 (N_12854,N_11875,N_11015);
xnor U12855 (N_12855,N_11190,N_11532);
nand U12856 (N_12856,N_11455,N_11571);
xor U12857 (N_12857,N_11070,N_11624);
nor U12858 (N_12858,N_11849,N_11099);
nor U12859 (N_12859,N_11502,N_11364);
xor U12860 (N_12860,N_11745,N_11280);
and U12861 (N_12861,N_11633,N_11017);
xor U12862 (N_12862,N_11649,N_11837);
nor U12863 (N_12863,N_11818,N_11826);
and U12864 (N_12864,N_11829,N_11078);
or U12865 (N_12865,N_11948,N_11795);
nor U12866 (N_12866,N_11635,N_11062);
and U12867 (N_12867,N_11547,N_11391);
nor U12868 (N_12868,N_11026,N_11656);
and U12869 (N_12869,N_11358,N_11275);
or U12870 (N_12870,N_11835,N_11802);
nand U12871 (N_12871,N_11525,N_11001);
nand U12872 (N_12872,N_11365,N_11730);
nand U12873 (N_12873,N_11230,N_11373);
or U12874 (N_12874,N_11575,N_11813);
xnor U12875 (N_12875,N_11751,N_11790);
nand U12876 (N_12876,N_11848,N_11146);
xnor U12877 (N_12877,N_11958,N_11486);
or U12878 (N_12878,N_11513,N_11065);
nor U12879 (N_12879,N_11614,N_11005);
nand U12880 (N_12880,N_11130,N_11105);
nor U12881 (N_12881,N_11866,N_11163);
or U12882 (N_12882,N_11953,N_11667);
or U12883 (N_12883,N_11041,N_11596);
and U12884 (N_12884,N_11438,N_11024);
nor U12885 (N_12885,N_11406,N_11091);
xor U12886 (N_12886,N_11626,N_11265);
nand U12887 (N_12887,N_11196,N_11164);
nand U12888 (N_12888,N_11234,N_11980);
or U12889 (N_12889,N_11979,N_11240);
nor U12890 (N_12890,N_11752,N_11613);
nand U12891 (N_12891,N_11916,N_11275);
xnor U12892 (N_12892,N_11311,N_11778);
xnor U12893 (N_12893,N_11037,N_11532);
nand U12894 (N_12894,N_11379,N_11272);
nor U12895 (N_12895,N_11975,N_11997);
and U12896 (N_12896,N_11148,N_11916);
or U12897 (N_12897,N_11461,N_11744);
and U12898 (N_12898,N_11589,N_11566);
xor U12899 (N_12899,N_11616,N_11481);
or U12900 (N_12900,N_11945,N_11161);
xor U12901 (N_12901,N_11778,N_11952);
or U12902 (N_12902,N_11962,N_11534);
nor U12903 (N_12903,N_11693,N_11501);
or U12904 (N_12904,N_11600,N_11643);
nand U12905 (N_12905,N_11411,N_11899);
or U12906 (N_12906,N_11437,N_11354);
or U12907 (N_12907,N_11050,N_11469);
and U12908 (N_12908,N_11735,N_11265);
xor U12909 (N_12909,N_11911,N_11792);
or U12910 (N_12910,N_11603,N_11985);
xnor U12911 (N_12911,N_11273,N_11643);
or U12912 (N_12912,N_11559,N_11571);
or U12913 (N_12913,N_11072,N_11232);
nor U12914 (N_12914,N_11850,N_11489);
nor U12915 (N_12915,N_11260,N_11457);
or U12916 (N_12916,N_11144,N_11929);
or U12917 (N_12917,N_11913,N_11150);
nand U12918 (N_12918,N_11725,N_11536);
or U12919 (N_12919,N_11310,N_11503);
xnor U12920 (N_12920,N_11611,N_11605);
nand U12921 (N_12921,N_11354,N_11298);
and U12922 (N_12922,N_11743,N_11986);
and U12923 (N_12923,N_11588,N_11498);
nand U12924 (N_12924,N_11261,N_11522);
nor U12925 (N_12925,N_11980,N_11297);
or U12926 (N_12926,N_11475,N_11699);
xnor U12927 (N_12927,N_11677,N_11143);
nor U12928 (N_12928,N_11329,N_11276);
nand U12929 (N_12929,N_11639,N_11157);
and U12930 (N_12930,N_11246,N_11739);
nand U12931 (N_12931,N_11002,N_11453);
and U12932 (N_12932,N_11020,N_11672);
nor U12933 (N_12933,N_11877,N_11411);
nand U12934 (N_12934,N_11828,N_11656);
nor U12935 (N_12935,N_11383,N_11358);
nand U12936 (N_12936,N_11164,N_11075);
or U12937 (N_12937,N_11972,N_11895);
nor U12938 (N_12938,N_11758,N_11048);
nor U12939 (N_12939,N_11372,N_11180);
and U12940 (N_12940,N_11381,N_11102);
xor U12941 (N_12941,N_11283,N_11700);
or U12942 (N_12942,N_11712,N_11293);
nor U12943 (N_12943,N_11534,N_11771);
xnor U12944 (N_12944,N_11502,N_11910);
and U12945 (N_12945,N_11341,N_11140);
and U12946 (N_12946,N_11395,N_11943);
or U12947 (N_12947,N_11983,N_11741);
nand U12948 (N_12948,N_11689,N_11717);
and U12949 (N_12949,N_11059,N_11680);
xor U12950 (N_12950,N_11724,N_11684);
and U12951 (N_12951,N_11767,N_11559);
nor U12952 (N_12952,N_11871,N_11155);
or U12953 (N_12953,N_11199,N_11211);
xnor U12954 (N_12954,N_11620,N_11242);
or U12955 (N_12955,N_11775,N_11453);
xor U12956 (N_12956,N_11762,N_11998);
or U12957 (N_12957,N_11993,N_11526);
and U12958 (N_12958,N_11187,N_11903);
and U12959 (N_12959,N_11550,N_11538);
and U12960 (N_12960,N_11511,N_11595);
and U12961 (N_12961,N_11002,N_11668);
nor U12962 (N_12962,N_11414,N_11079);
and U12963 (N_12963,N_11772,N_11147);
nand U12964 (N_12964,N_11334,N_11069);
nor U12965 (N_12965,N_11683,N_11014);
nand U12966 (N_12966,N_11694,N_11768);
nor U12967 (N_12967,N_11432,N_11989);
xnor U12968 (N_12968,N_11892,N_11069);
xnor U12969 (N_12969,N_11425,N_11136);
nor U12970 (N_12970,N_11109,N_11707);
or U12971 (N_12971,N_11628,N_11300);
and U12972 (N_12972,N_11796,N_11092);
or U12973 (N_12973,N_11178,N_11811);
nor U12974 (N_12974,N_11944,N_11521);
or U12975 (N_12975,N_11596,N_11097);
nor U12976 (N_12976,N_11323,N_11286);
and U12977 (N_12977,N_11943,N_11564);
nand U12978 (N_12978,N_11899,N_11274);
and U12979 (N_12979,N_11658,N_11668);
or U12980 (N_12980,N_11332,N_11357);
or U12981 (N_12981,N_11367,N_11043);
nor U12982 (N_12982,N_11919,N_11063);
and U12983 (N_12983,N_11034,N_11904);
xor U12984 (N_12984,N_11365,N_11268);
nand U12985 (N_12985,N_11270,N_11447);
and U12986 (N_12986,N_11367,N_11258);
nand U12987 (N_12987,N_11774,N_11977);
and U12988 (N_12988,N_11929,N_11346);
xnor U12989 (N_12989,N_11444,N_11104);
or U12990 (N_12990,N_11154,N_11849);
and U12991 (N_12991,N_11911,N_11262);
or U12992 (N_12992,N_11813,N_11069);
nor U12993 (N_12993,N_11298,N_11953);
or U12994 (N_12994,N_11082,N_11946);
nor U12995 (N_12995,N_11213,N_11998);
xnor U12996 (N_12996,N_11102,N_11458);
or U12997 (N_12997,N_11929,N_11348);
and U12998 (N_12998,N_11400,N_11851);
or U12999 (N_12999,N_11354,N_11826);
or U13000 (N_13000,N_12447,N_12649);
nand U13001 (N_13001,N_12458,N_12273);
nor U13002 (N_13002,N_12655,N_12350);
xnor U13003 (N_13003,N_12677,N_12910);
xnor U13004 (N_13004,N_12881,N_12294);
xnor U13005 (N_13005,N_12626,N_12150);
nand U13006 (N_13006,N_12112,N_12564);
xnor U13007 (N_13007,N_12025,N_12091);
and U13008 (N_13008,N_12045,N_12977);
or U13009 (N_13009,N_12650,N_12597);
nand U13010 (N_13010,N_12386,N_12179);
nand U13011 (N_13011,N_12252,N_12737);
xor U13012 (N_13012,N_12444,N_12763);
or U13013 (N_13013,N_12725,N_12586);
and U13014 (N_13014,N_12746,N_12728);
or U13015 (N_13015,N_12871,N_12792);
nand U13016 (N_13016,N_12063,N_12611);
nor U13017 (N_13017,N_12408,N_12799);
or U13018 (N_13018,N_12516,N_12837);
and U13019 (N_13019,N_12071,N_12341);
or U13020 (N_13020,N_12125,N_12151);
nor U13021 (N_13021,N_12018,N_12998);
or U13022 (N_13022,N_12777,N_12664);
xor U13023 (N_13023,N_12358,N_12322);
or U13024 (N_13024,N_12654,N_12304);
nand U13025 (N_13025,N_12566,N_12550);
nor U13026 (N_13026,N_12944,N_12781);
nand U13027 (N_13027,N_12807,N_12852);
and U13028 (N_13028,N_12308,N_12765);
xnor U13029 (N_13029,N_12920,N_12375);
xnor U13030 (N_13030,N_12412,N_12607);
nor U13031 (N_13031,N_12318,N_12571);
or U13032 (N_13032,N_12744,N_12190);
and U13033 (N_13033,N_12676,N_12971);
or U13034 (N_13034,N_12320,N_12061);
nand U13035 (N_13035,N_12614,N_12577);
nor U13036 (N_13036,N_12531,N_12848);
xor U13037 (N_13037,N_12689,N_12263);
xor U13038 (N_13038,N_12834,N_12145);
xor U13039 (N_13039,N_12030,N_12931);
and U13040 (N_13040,N_12508,N_12489);
nand U13041 (N_13041,N_12115,N_12438);
xor U13042 (N_13042,N_12682,N_12104);
nand U13043 (N_13043,N_12583,N_12835);
xor U13044 (N_13044,N_12478,N_12327);
nor U13045 (N_13045,N_12722,N_12193);
nor U13046 (N_13046,N_12079,N_12058);
nand U13047 (N_13047,N_12203,N_12879);
nor U13048 (N_13048,N_12015,N_12787);
nor U13049 (N_13049,N_12736,N_12169);
or U13050 (N_13050,N_12174,N_12943);
xor U13051 (N_13051,N_12527,N_12209);
or U13052 (N_13052,N_12714,N_12856);
and U13053 (N_13053,N_12289,N_12403);
and U13054 (N_13054,N_12991,N_12078);
nand U13055 (N_13055,N_12376,N_12219);
or U13056 (N_13056,N_12176,N_12225);
nor U13057 (N_13057,N_12361,N_12707);
nand U13058 (N_13058,N_12536,N_12981);
or U13059 (N_13059,N_12790,N_12757);
nor U13060 (N_13060,N_12342,N_12087);
or U13061 (N_13061,N_12978,N_12627);
nor U13062 (N_13062,N_12214,N_12238);
or U13063 (N_13063,N_12926,N_12286);
and U13064 (N_13064,N_12461,N_12565);
and U13065 (N_13065,N_12643,N_12401);
xnor U13066 (N_13066,N_12783,N_12959);
nand U13067 (N_13067,N_12568,N_12929);
and U13068 (N_13068,N_12735,N_12223);
xnor U13069 (N_13069,N_12927,N_12751);
xnor U13070 (N_13070,N_12280,N_12900);
nand U13071 (N_13071,N_12637,N_12892);
xnor U13072 (N_13072,N_12387,N_12084);
nor U13073 (N_13073,N_12505,N_12231);
and U13074 (N_13074,N_12158,N_12641);
nand U13075 (N_13075,N_12086,N_12905);
and U13076 (N_13076,N_12192,N_12945);
nor U13077 (N_13077,N_12004,N_12590);
or U13078 (N_13078,N_12888,N_12165);
and U13079 (N_13079,N_12443,N_12628);
nor U13080 (N_13080,N_12889,N_12396);
nor U13081 (N_13081,N_12237,N_12954);
nand U13082 (N_13082,N_12661,N_12863);
nor U13083 (N_13083,N_12884,N_12081);
nand U13084 (N_13084,N_12213,N_12405);
and U13085 (N_13085,N_12847,N_12742);
or U13086 (N_13086,N_12809,N_12043);
xnor U13087 (N_13087,N_12123,N_12352);
or U13088 (N_13088,N_12349,N_12916);
nor U13089 (N_13089,N_12932,N_12394);
and U13090 (N_13090,N_12930,N_12957);
and U13091 (N_13091,N_12103,N_12357);
nand U13092 (N_13092,N_12317,N_12975);
nor U13093 (N_13093,N_12532,N_12970);
nor U13094 (N_13094,N_12197,N_12064);
or U13095 (N_13095,N_12748,N_12082);
nor U13096 (N_13096,N_12581,N_12268);
and U13097 (N_13097,N_12715,N_12925);
and U13098 (N_13098,N_12230,N_12758);
or U13099 (N_13099,N_12134,N_12982);
nand U13100 (N_13100,N_12874,N_12328);
and U13101 (N_13101,N_12688,N_12582);
nand U13102 (N_13102,N_12028,N_12321);
nor U13103 (N_13103,N_12769,N_12877);
xnor U13104 (N_13104,N_12200,N_12723);
xnor U13105 (N_13105,N_12099,N_12986);
and U13106 (N_13106,N_12496,N_12038);
and U13107 (N_13107,N_12913,N_12974);
nor U13108 (N_13108,N_12906,N_12631);
and U13109 (N_13109,N_12747,N_12760);
nand U13110 (N_13110,N_12094,N_12116);
nand U13111 (N_13111,N_12288,N_12338);
and U13112 (N_13112,N_12096,N_12298);
or U13113 (N_13113,N_12662,N_12029);
nand U13114 (N_13114,N_12698,N_12040);
or U13115 (N_13115,N_12445,N_12561);
or U13116 (N_13116,N_12469,N_12663);
xnor U13117 (N_13117,N_12782,N_12759);
or U13118 (N_13118,N_12152,N_12708);
xor U13119 (N_13119,N_12741,N_12600);
or U13120 (N_13120,N_12014,N_12805);
nand U13121 (N_13121,N_12454,N_12222);
nor U13122 (N_13122,N_12578,N_12784);
or U13123 (N_13123,N_12267,N_12825);
nor U13124 (N_13124,N_12060,N_12316);
xor U13125 (N_13125,N_12514,N_12528);
nand U13126 (N_13126,N_12258,N_12955);
and U13127 (N_13127,N_12857,N_12325);
nor U13128 (N_13128,N_12279,N_12210);
nand U13129 (N_13129,N_12635,N_12425);
nand U13130 (N_13130,N_12181,N_12501);
xnor U13131 (N_13131,N_12265,N_12921);
xnor U13132 (N_13132,N_12126,N_12131);
xnor U13133 (N_13133,N_12333,N_12594);
and U13134 (N_13134,N_12147,N_12031);
and U13135 (N_13135,N_12716,N_12163);
and U13136 (N_13136,N_12901,N_12711);
nor U13137 (N_13137,N_12039,N_12618);
xor U13138 (N_13138,N_12243,N_12605);
or U13139 (N_13139,N_12420,N_12950);
nand U13140 (N_13140,N_12392,N_12699);
nand U13141 (N_13141,N_12453,N_12184);
xor U13142 (N_13142,N_12953,N_12724);
or U13143 (N_13143,N_12657,N_12612);
xnor U13144 (N_13144,N_12359,N_12095);
nor U13145 (N_13145,N_12673,N_12632);
nor U13146 (N_13146,N_12199,N_12823);
and U13147 (N_13147,N_12753,N_12585);
or U13148 (N_13148,N_12068,N_12653);
and U13149 (N_13149,N_12895,N_12819);
and U13150 (N_13150,N_12482,N_12882);
nand U13151 (N_13151,N_12544,N_12264);
nor U13152 (N_13152,N_12755,N_12864);
nand U13153 (N_13153,N_12241,N_12890);
or U13154 (N_13154,N_12355,N_12220);
xor U13155 (N_13155,N_12026,N_12979);
nand U13156 (N_13156,N_12912,N_12395);
and U13157 (N_13157,N_12269,N_12495);
or U13158 (N_13158,N_12615,N_12323);
or U13159 (N_13159,N_12599,N_12511);
xnor U13160 (N_13160,N_12939,N_12849);
nor U13161 (N_13161,N_12667,N_12419);
or U13162 (N_13162,N_12644,N_12307);
xor U13163 (N_13163,N_12178,N_12076);
and U13164 (N_13164,N_12416,N_12907);
or U13165 (N_13165,N_12138,N_12869);
and U13166 (N_13166,N_12827,N_12720);
or U13167 (N_13167,N_12567,N_12659);
nor U13168 (N_13168,N_12132,N_12604);
nor U13169 (N_13169,N_12646,N_12460);
or U13170 (N_13170,N_12917,N_12775);
nand U13171 (N_13171,N_12051,N_12171);
or U13172 (N_13172,N_12113,N_12162);
xor U13173 (N_13173,N_12250,N_12694);
nor U13174 (N_13174,N_12382,N_12485);
and U13175 (N_13175,N_12674,N_12154);
xnor U13176 (N_13176,N_12842,N_12666);
or U13177 (N_13177,N_12833,N_12009);
or U13178 (N_13178,N_12232,N_12148);
xnor U13179 (N_13179,N_12384,N_12455);
and U13180 (N_13180,N_12185,N_12924);
nor U13181 (N_13181,N_12236,N_12845);
or U13182 (N_13182,N_12940,N_12011);
nand U13183 (N_13183,N_12065,N_12483);
or U13184 (N_13184,N_12196,N_12817);
or U13185 (N_13185,N_12701,N_12534);
nand U13186 (N_13186,N_12128,N_12140);
or U13187 (N_13187,N_12703,N_12885);
nand U13188 (N_13188,N_12191,N_12397);
xnor U13189 (N_13189,N_12985,N_12980);
xnor U13190 (N_13190,N_12398,N_12348);
xor U13191 (N_13191,N_12537,N_12442);
xor U13192 (N_13192,N_12865,N_12306);
xnor U13193 (N_13193,N_12923,N_12013);
and U13194 (N_13194,N_12297,N_12303);
xnor U13195 (N_13195,N_12343,N_12276);
xor U13196 (N_13196,N_12786,N_12434);
nor U13197 (N_13197,N_12378,N_12969);
nand U13198 (N_13198,N_12066,N_12549);
xnor U13199 (N_13199,N_12972,N_12570);
and U13200 (N_13200,N_12391,N_12774);
xnor U13201 (N_13201,N_12617,N_12771);
and U13202 (N_13202,N_12996,N_12610);
or U13203 (N_13203,N_12616,N_12691);
or U13204 (N_13204,N_12356,N_12545);
and U13205 (N_13205,N_12168,N_12976);
nor U13206 (N_13206,N_12421,N_12602);
and U13207 (N_13207,N_12936,N_12413);
or U13208 (N_13208,N_12839,N_12105);
xor U13209 (N_13209,N_12731,N_12999);
and U13210 (N_13210,N_12451,N_12800);
nor U13211 (N_13211,N_12933,N_12205);
and U13212 (N_13212,N_12021,N_12056);
or U13213 (N_13213,N_12876,N_12629);
nor U13214 (N_13214,N_12942,N_12326);
or U13215 (N_13215,N_12207,N_12843);
nand U13216 (N_13216,N_12499,N_12872);
xnor U13217 (N_13217,N_12388,N_12409);
nor U13218 (N_13218,N_12291,N_12563);
and U13219 (N_13219,N_12177,N_12656);
nand U13220 (N_13220,N_12201,N_12172);
or U13221 (N_13221,N_12354,N_12141);
and U13222 (N_13222,N_12475,N_12070);
nand U13223 (N_13223,N_12853,N_12194);
or U13224 (N_13224,N_12486,N_12133);
nor U13225 (N_13225,N_12640,N_12430);
or U13226 (N_13226,N_12389,N_12779);
or U13227 (N_13227,N_12719,N_12363);
xor U13228 (N_13228,N_12353,N_12858);
and U13229 (N_13229,N_12958,N_12949);
nand U13230 (N_13230,N_12217,N_12365);
nand U13231 (N_13231,N_12813,N_12457);
or U13232 (N_13232,N_12149,N_12449);
nor U13233 (N_13233,N_12752,N_12860);
nand U13234 (N_13234,N_12780,N_12732);
nor U13235 (N_13235,N_12313,N_12639);
and U13236 (N_13236,N_12248,N_12255);
or U13237 (N_13237,N_12880,N_12198);
nand U13238 (N_13238,N_12346,N_12399);
or U13239 (N_13239,N_12624,N_12471);
nor U13240 (N_13240,N_12681,N_12883);
xnor U13241 (N_13241,N_12216,N_12767);
nand U13242 (N_13242,N_12000,N_12832);
or U13243 (N_13243,N_12902,N_12793);
nor U13244 (N_13244,N_12796,N_12299);
xnor U13245 (N_13245,N_12504,N_12810);
nand U13246 (N_13246,N_12085,N_12776);
nand U13247 (N_13247,N_12117,N_12558);
or U13248 (N_13248,N_12464,N_12107);
xor U13249 (N_13249,N_12282,N_12239);
nand U13250 (N_13250,N_12315,N_12592);
and U13251 (N_13251,N_12543,N_12756);
nor U13252 (N_13252,N_12973,N_12588);
nor U13253 (N_13253,N_12334,N_12642);
and U13254 (N_13254,N_12859,N_12111);
and U13255 (N_13255,N_12645,N_12702);
and U13256 (N_13256,N_12696,N_12142);
nor U13257 (N_13257,N_12685,N_12452);
or U13258 (N_13258,N_12136,N_12006);
and U13259 (N_13259,N_12789,N_12608);
xnor U13260 (N_13260,N_12838,N_12101);
nand U13261 (N_13261,N_12120,N_12329);
and U13262 (N_13262,N_12740,N_12046);
nand U13263 (N_13263,N_12274,N_12773);
xnor U13264 (N_13264,N_12754,N_12952);
nand U13265 (N_13265,N_12240,N_12795);
xnor U13266 (N_13266,N_12287,N_12922);
or U13267 (N_13267,N_12670,N_12426);
and U13268 (N_13268,N_12552,N_12831);
or U13269 (N_13269,N_12814,N_12480);
nand U13270 (N_13270,N_12024,N_12050);
or U13271 (N_13271,N_12470,N_12705);
nor U13272 (N_13272,N_12556,N_12547);
xor U13273 (N_13273,N_12344,N_12467);
or U13274 (N_13274,N_12652,N_12233);
xnor U13275 (N_13275,N_12048,N_12235);
or U13276 (N_13276,N_12494,N_12512);
or U13277 (N_13277,N_12032,N_12156);
or U13278 (N_13278,N_12366,N_12224);
xor U13279 (N_13279,N_12429,N_12821);
or U13280 (N_13280,N_12428,N_12054);
xor U13281 (N_13281,N_12538,N_12301);
or U13282 (N_13282,N_12557,N_12381);
nor U13283 (N_13283,N_12373,N_12803);
and U13284 (N_13284,N_12533,N_12946);
and U13285 (N_13285,N_12347,N_12539);
xnor U13286 (N_13286,N_12770,N_12651);
or U13287 (N_13287,N_12266,N_12129);
nand U13288 (N_13288,N_12794,N_12330);
and U13289 (N_13289,N_12840,N_12820);
nor U13290 (N_13290,N_12003,N_12569);
and U13291 (N_13291,N_12414,N_12717);
or U13292 (N_13292,N_12816,N_12098);
or U13293 (N_13293,N_12437,N_12992);
and U13294 (N_13294,N_12622,N_12672);
nand U13295 (N_13295,N_12370,N_12878);
or U13296 (N_13296,N_12130,N_12285);
or U13297 (N_13297,N_12402,N_12909);
nand U13298 (N_13298,N_12540,N_12498);
or U13299 (N_13299,N_12053,N_12693);
and U13300 (N_13300,N_12424,N_12075);
nand U13301 (N_13301,N_12122,N_12182);
nor U13302 (N_13302,N_12124,N_12801);
and U13303 (N_13303,N_12340,N_12351);
or U13304 (N_13304,N_12027,N_12706);
xor U13305 (N_13305,N_12868,N_12671);
xor U13306 (N_13306,N_12309,N_12658);
nand U13307 (N_13307,N_12897,N_12180);
xnor U13308 (N_13308,N_12143,N_12433);
and U13309 (N_13309,N_12743,N_12368);
nor U13310 (N_13310,N_12983,N_12580);
or U13311 (N_13311,N_12680,N_12862);
nand U13312 (N_13312,N_12490,N_12683);
xor U13313 (N_13313,N_12886,N_12811);
xnor U13314 (N_13314,N_12961,N_12367);
nor U13315 (N_13315,N_12968,N_12293);
nand U13316 (N_13316,N_12385,N_12146);
nand U13317 (N_13317,N_12155,N_12899);
or U13318 (N_13318,N_12894,N_12074);
or U13319 (N_13319,N_12523,N_12687);
nand U13320 (N_13320,N_12606,N_12477);
or U13321 (N_13321,N_12553,N_12422);
nand U13322 (N_13322,N_12587,N_12476);
and U13323 (N_13323,N_12515,N_12484);
and U13324 (N_13324,N_12559,N_12530);
and U13325 (N_13325,N_12620,N_12634);
xnor U13326 (N_13326,N_12984,N_12067);
and U13327 (N_13327,N_12047,N_12690);
xnor U13328 (N_13328,N_12941,N_12345);
nor U13329 (N_13329,N_12797,N_12844);
nor U13330 (N_13330,N_12911,N_12069);
or U13331 (N_13331,N_12601,N_12187);
nor U13332 (N_13332,N_12001,N_12830);
and U13333 (N_13333,N_12314,N_12492);
nand U13334 (N_13334,N_12709,N_12818);
or U13335 (N_13335,N_12679,N_12675);
nand U13336 (N_13336,N_12007,N_12948);
and U13337 (N_13337,N_12097,N_12745);
or U13338 (N_13338,N_12406,N_12546);
or U13339 (N_13339,N_12102,N_12555);
or U13340 (N_13340,N_12541,N_12463);
nor U13341 (N_13341,N_12609,N_12665);
xnor U13342 (N_13342,N_12491,N_12144);
nand U13343 (N_13343,N_12251,N_12695);
nand U13344 (N_13344,N_12603,N_12826);
and U13345 (N_13345,N_12383,N_12296);
xor U13346 (N_13346,N_12410,N_12619);
and U13347 (N_13347,N_12059,N_12427);
xnor U13348 (N_13348,N_12440,N_12589);
nor U13349 (N_13349,N_12034,N_12822);
xnor U13350 (N_13350,N_12850,N_12204);
xor U13351 (N_13351,N_12551,N_12254);
nand U13352 (N_13352,N_12554,N_12016);
nand U13353 (N_13353,N_12808,N_12517);
and U13354 (N_13354,N_12507,N_12560);
nand U13355 (N_13355,N_12915,N_12211);
nand U13356 (N_13356,N_12260,N_12037);
or U13357 (N_13357,N_12188,N_12022);
xnor U13358 (N_13358,N_12372,N_12290);
and U13359 (N_13359,N_12764,N_12183);
or U13360 (N_13360,N_12121,N_12228);
nor U13361 (N_13361,N_12374,N_12311);
and U13362 (N_13362,N_12520,N_12019);
xnor U13363 (N_13363,N_12989,N_12167);
nor U13364 (N_13364,N_12215,N_12033);
nand U13365 (N_13365,N_12573,N_12562);
nor U13366 (N_13366,N_12990,N_12093);
or U13367 (N_13367,N_12500,N_12778);
or U13368 (N_13368,N_12513,N_12170);
xor U13369 (N_13369,N_12896,N_12278);
or U13370 (N_13370,N_12815,N_12503);
nor U13371 (N_13371,N_12727,N_12415);
and U13372 (N_13372,N_12008,N_12023);
or U13373 (N_13373,N_12854,N_12791);
nor U13374 (N_13374,N_12903,N_12474);
nand U13375 (N_13375,N_12281,N_12904);
and U13376 (N_13376,N_12468,N_12479);
xor U13377 (N_13377,N_12108,N_12529);
or U13378 (N_13378,N_12497,N_12456);
or U13379 (N_13379,N_12035,N_12522);
nor U13380 (N_13380,N_12488,N_12855);
and U13381 (N_13381,N_12057,N_12481);
or U13382 (N_13382,N_12431,N_12244);
nor U13383 (N_13383,N_12017,N_12947);
nand U13384 (N_13384,N_12083,N_12221);
and U13385 (N_13385,N_12502,N_12089);
or U13386 (N_13386,N_12119,N_12668);
nor U13387 (N_13387,N_12118,N_12613);
and U13388 (N_13388,N_12647,N_12772);
or U13389 (N_13389,N_12153,N_12377);
nand U13390 (N_13390,N_12242,N_12020);
xor U13391 (N_13391,N_12055,N_12284);
nor U13392 (N_13392,N_12465,N_12730);
xnor U13393 (N_13393,N_12202,N_12630);
nand U13394 (N_13394,N_12127,N_12466);
and U13395 (N_13395,N_12621,N_12506);
and U13396 (N_13396,N_12110,N_12312);
xnor U13397 (N_13397,N_12336,N_12369);
or U13398 (N_13398,N_12684,N_12319);
nand U13399 (N_13399,N_12261,N_12305);
or U13400 (N_13400,N_12472,N_12012);
or U13401 (N_13401,N_12393,N_12548);
and U13402 (N_13402,N_12166,N_12697);
nor U13403 (N_13403,N_12524,N_12462);
nand U13404 (N_13404,N_12960,N_12951);
nor U13405 (N_13405,N_12788,N_12535);
nand U13406 (N_13406,N_12824,N_12212);
nor U13407 (N_13407,N_12812,N_12851);
xor U13408 (N_13408,N_12994,N_12189);
nor U13409 (N_13409,N_12870,N_12195);
nor U13410 (N_13410,N_12302,N_12928);
or U13411 (N_13411,N_12114,N_12249);
xnor U13412 (N_13412,N_12283,N_12660);
and U13413 (N_13413,N_12160,N_12584);
xor U13414 (N_13414,N_12161,N_12247);
and U13415 (N_13415,N_12400,N_12432);
nand U13416 (N_13416,N_12253,N_12270);
nand U13417 (N_13417,N_12487,N_12245);
or U13418 (N_13418,N_12712,N_12967);
xor U13419 (N_13419,N_12893,N_12234);
and U13420 (N_13420,N_12339,N_12914);
xnor U13421 (N_13421,N_12766,N_12829);
nor U13422 (N_13422,N_12988,N_12875);
nor U13423 (N_13423,N_12246,N_12137);
nand U13424 (N_13424,N_12411,N_12519);
xor U13425 (N_13425,N_12841,N_12077);
nand U13426 (N_13426,N_12718,N_12785);
nand U13427 (N_13427,N_12935,N_12934);
xor U13428 (N_13428,N_12277,N_12997);
or U13429 (N_13429,N_12729,N_12633);
nor U13430 (N_13430,N_12518,N_12836);
and U13431 (N_13431,N_12157,N_12956);
or U13432 (N_13432,N_12139,N_12937);
xnor U13433 (N_13433,N_12572,N_12739);
or U13434 (N_13434,N_12257,N_12423);
nor U13435 (N_13435,N_12768,N_12435);
or U13436 (N_13436,N_12750,N_12186);
xnor U13437 (N_13437,N_12762,N_12272);
xnor U13438 (N_13438,N_12073,N_12275);
xnor U13439 (N_13439,N_12227,N_12579);
and U13440 (N_13440,N_12595,N_12090);
xnor U13441 (N_13441,N_12407,N_12828);
or U13442 (N_13442,N_12390,N_12576);
and U13443 (N_13443,N_12404,N_12072);
or U13444 (N_13444,N_12526,N_12987);
or U13445 (N_13445,N_12638,N_12337);
xor U13446 (N_13446,N_12159,N_12798);
xnor U13447 (N_13447,N_12436,N_12648);
and U13448 (N_13448,N_12574,N_12379);
nand U13449 (N_13449,N_12259,N_12713);
nand U13450 (N_13450,N_12625,N_12861);
and U13451 (N_13451,N_12510,N_12866);
and U13452 (N_13452,N_12206,N_12229);
xor U13453 (N_13453,N_12598,N_12300);
nor U13454 (N_13454,N_12088,N_12908);
xnor U13455 (N_13455,N_12686,N_12010);
nor U13456 (N_13456,N_12459,N_12439);
nand U13457 (N_13457,N_12575,N_12591);
and U13458 (N_13458,N_12036,N_12310);
or U13459 (N_13459,N_12963,N_12804);
nor U13460 (N_13460,N_12802,N_12734);
nor U13461 (N_13461,N_12898,N_12100);
nor U13462 (N_13462,N_12335,N_12761);
nor U13463 (N_13463,N_12593,N_12173);
or U13464 (N_13464,N_12324,N_12380);
nor U13465 (N_13465,N_12473,N_12596);
nand U13466 (N_13466,N_12919,N_12509);
or U13467 (N_13467,N_12262,N_12005);
xnor U13468 (N_13468,N_12891,N_12623);
and U13469 (N_13469,N_12636,N_12041);
or U13470 (N_13470,N_12710,N_12042);
xnor U13471 (N_13471,N_12867,N_12806);
and U13472 (N_13472,N_12873,N_12738);
and U13473 (N_13473,N_12704,N_12441);
nand U13474 (N_13474,N_12292,N_12700);
xor U13475 (N_13475,N_12846,N_12678);
nand U13476 (N_13476,N_12962,N_12542);
xor U13477 (N_13477,N_12993,N_12938);
nand U13478 (N_13478,N_12049,N_12175);
and U13479 (N_13479,N_12295,N_12446);
xor U13480 (N_13480,N_12164,N_12721);
and U13481 (N_13481,N_12052,N_12362);
or U13482 (N_13482,N_12106,N_12525);
and U13483 (N_13483,N_12733,N_12450);
xor U13484 (N_13484,N_12332,N_12418);
nor U13485 (N_13485,N_12371,N_12218);
and U13486 (N_13486,N_12092,N_12726);
nor U13487 (N_13487,N_12964,N_12448);
or U13488 (N_13488,N_12002,N_12360);
or U13489 (N_13489,N_12995,N_12109);
nor U13490 (N_13490,N_12669,N_12080);
or U13491 (N_13491,N_12208,N_12493);
nand U13492 (N_13492,N_12692,N_12364);
nor U13493 (N_13493,N_12135,N_12887);
nor U13494 (N_13494,N_12044,N_12271);
or U13495 (N_13495,N_12331,N_12062);
and U13496 (N_13496,N_12226,N_12966);
xor U13497 (N_13497,N_12749,N_12521);
and U13498 (N_13498,N_12965,N_12256);
xnor U13499 (N_13499,N_12918,N_12417);
xnor U13500 (N_13500,N_12474,N_12971);
nor U13501 (N_13501,N_12185,N_12797);
and U13502 (N_13502,N_12797,N_12302);
nand U13503 (N_13503,N_12736,N_12887);
or U13504 (N_13504,N_12480,N_12198);
or U13505 (N_13505,N_12556,N_12452);
or U13506 (N_13506,N_12321,N_12836);
nand U13507 (N_13507,N_12743,N_12170);
or U13508 (N_13508,N_12914,N_12371);
nand U13509 (N_13509,N_12223,N_12752);
nor U13510 (N_13510,N_12408,N_12662);
nand U13511 (N_13511,N_12942,N_12748);
and U13512 (N_13512,N_12929,N_12723);
and U13513 (N_13513,N_12229,N_12312);
or U13514 (N_13514,N_12111,N_12482);
xor U13515 (N_13515,N_12683,N_12357);
and U13516 (N_13516,N_12149,N_12137);
nor U13517 (N_13517,N_12569,N_12358);
and U13518 (N_13518,N_12122,N_12188);
and U13519 (N_13519,N_12716,N_12957);
nand U13520 (N_13520,N_12553,N_12629);
xnor U13521 (N_13521,N_12819,N_12435);
nand U13522 (N_13522,N_12601,N_12027);
xnor U13523 (N_13523,N_12259,N_12893);
and U13524 (N_13524,N_12109,N_12838);
or U13525 (N_13525,N_12792,N_12880);
nor U13526 (N_13526,N_12331,N_12119);
xor U13527 (N_13527,N_12337,N_12349);
nor U13528 (N_13528,N_12026,N_12425);
nor U13529 (N_13529,N_12765,N_12444);
and U13530 (N_13530,N_12082,N_12261);
nor U13531 (N_13531,N_12998,N_12031);
and U13532 (N_13532,N_12354,N_12508);
xnor U13533 (N_13533,N_12473,N_12470);
nand U13534 (N_13534,N_12078,N_12329);
nand U13535 (N_13535,N_12635,N_12416);
and U13536 (N_13536,N_12338,N_12712);
and U13537 (N_13537,N_12034,N_12809);
nand U13538 (N_13538,N_12555,N_12838);
nand U13539 (N_13539,N_12101,N_12926);
nor U13540 (N_13540,N_12441,N_12608);
and U13541 (N_13541,N_12940,N_12825);
xnor U13542 (N_13542,N_12728,N_12499);
and U13543 (N_13543,N_12345,N_12711);
nor U13544 (N_13544,N_12215,N_12122);
and U13545 (N_13545,N_12705,N_12136);
xnor U13546 (N_13546,N_12652,N_12572);
xnor U13547 (N_13547,N_12794,N_12506);
xnor U13548 (N_13548,N_12790,N_12127);
xor U13549 (N_13549,N_12669,N_12769);
xor U13550 (N_13550,N_12531,N_12275);
xor U13551 (N_13551,N_12651,N_12997);
xor U13552 (N_13552,N_12316,N_12428);
xnor U13553 (N_13553,N_12853,N_12609);
nand U13554 (N_13554,N_12713,N_12759);
xor U13555 (N_13555,N_12396,N_12799);
nor U13556 (N_13556,N_12898,N_12240);
xnor U13557 (N_13557,N_12788,N_12278);
xnor U13558 (N_13558,N_12871,N_12134);
xor U13559 (N_13559,N_12834,N_12898);
nor U13560 (N_13560,N_12772,N_12155);
nor U13561 (N_13561,N_12486,N_12125);
or U13562 (N_13562,N_12406,N_12400);
nor U13563 (N_13563,N_12150,N_12596);
nor U13564 (N_13564,N_12941,N_12321);
nor U13565 (N_13565,N_12463,N_12389);
and U13566 (N_13566,N_12225,N_12013);
and U13567 (N_13567,N_12753,N_12656);
xnor U13568 (N_13568,N_12108,N_12221);
xnor U13569 (N_13569,N_12269,N_12831);
nand U13570 (N_13570,N_12522,N_12890);
nand U13571 (N_13571,N_12401,N_12805);
xnor U13572 (N_13572,N_12503,N_12023);
xnor U13573 (N_13573,N_12808,N_12235);
and U13574 (N_13574,N_12123,N_12856);
and U13575 (N_13575,N_12746,N_12794);
or U13576 (N_13576,N_12691,N_12956);
nor U13577 (N_13577,N_12001,N_12852);
xnor U13578 (N_13578,N_12108,N_12389);
xnor U13579 (N_13579,N_12916,N_12667);
nand U13580 (N_13580,N_12816,N_12383);
nor U13581 (N_13581,N_12582,N_12865);
and U13582 (N_13582,N_12701,N_12786);
or U13583 (N_13583,N_12290,N_12196);
or U13584 (N_13584,N_12773,N_12437);
nor U13585 (N_13585,N_12031,N_12017);
and U13586 (N_13586,N_12597,N_12673);
and U13587 (N_13587,N_12885,N_12655);
nand U13588 (N_13588,N_12582,N_12833);
nor U13589 (N_13589,N_12249,N_12739);
nand U13590 (N_13590,N_12035,N_12910);
and U13591 (N_13591,N_12418,N_12504);
nor U13592 (N_13592,N_12103,N_12485);
nand U13593 (N_13593,N_12066,N_12014);
or U13594 (N_13594,N_12149,N_12809);
and U13595 (N_13595,N_12946,N_12244);
nor U13596 (N_13596,N_12286,N_12921);
nor U13597 (N_13597,N_12374,N_12812);
and U13598 (N_13598,N_12738,N_12845);
or U13599 (N_13599,N_12422,N_12488);
nor U13600 (N_13600,N_12710,N_12238);
or U13601 (N_13601,N_12919,N_12218);
xnor U13602 (N_13602,N_12129,N_12529);
nor U13603 (N_13603,N_12450,N_12807);
or U13604 (N_13604,N_12601,N_12378);
or U13605 (N_13605,N_12210,N_12608);
and U13606 (N_13606,N_12164,N_12370);
and U13607 (N_13607,N_12821,N_12011);
or U13608 (N_13608,N_12121,N_12469);
nand U13609 (N_13609,N_12895,N_12566);
nand U13610 (N_13610,N_12891,N_12399);
and U13611 (N_13611,N_12420,N_12442);
nor U13612 (N_13612,N_12837,N_12246);
and U13613 (N_13613,N_12626,N_12474);
and U13614 (N_13614,N_12764,N_12841);
or U13615 (N_13615,N_12508,N_12415);
xor U13616 (N_13616,N_12179,N_12263);
nand U13617 (N_13617,N_12254,N_12484);
and U13618 (N_13618,N_12349,N_12624);
nand U13619 (N_13619,N_12089,N_12786);
nor U13620 (N_13620,N_12084,N_12104);
nand U13621 (N_13621,N_12875,N_12169);
nand U13622 (N_13622,N_12159,N_12700);
nand U13623 (N_13623,N_12917,N_12969);
nand U13624 (N_13624,N_12063,N_12868);
xnor U13625 (N_13625,N_12331,N_12894);
and U13626 (N_13626,N_12627,N_12968);
nand U13627 (N_13627,N_12097,N_12854);
nand U13628 (N_13628,N_12735,N_12693);
xor U13629 (N_13629,N_12228,N_12096);
xnor U13630 (N_13630,N_12630,N_12991);
nor U13631 (N_13631,N_12538,N_12304);
nand U13632 (N_13632,N_12429,N_12492);
or U13633 (N_13633,N_12342,N_12289);
nor U13634 (N_13634,N_12089,N_12396);
xor U13635 (N_13635,N_12043,N_12645);
nor U13636 (N_13636,N_12687,N_12467);
nor U13637 (N_13637,N_12171,N_12614);
xnor U13638 (N_13638,N_12091,N_12276);
nand U13639 (N_13639,N_12628,N_12648);
or U13640 (N_13640,N_12563,N_12468);
and U13641 (N_13641,N_12774,N_12186);
xnor U13642 (N_13642,N_12477,N_12167);
xnor U13643 (N_13643,N_12920,N_12024);
nand U13644 (N_13644,N_12668,N_12472);
and U13645 (N_13645,N_12015,N_12707);
or U13646 (N_13646,N_12625,N_12690);
nor U13647 (N_13647,N_12231,N_12521);
nor U13648 (N_13648,N_12315,N_12284);
xnor U13649 (N_13649,N_12660,N_12232);
nor U13650 (N_13650,N_12120,N_12962);
and U13651 (N_13651,N_12512,N_12624);
and U13652 (N_13652,N_12052,N_12991);
nand U13653 (N_13653,N_12662,N_12502);
nor U13654 (N_13654,N_12145,N_12408);
or U13655 (N_13655,N_12607,N_12887);
nand U13656 (N_13656,N_12564,N_12051);
and U13657 (N_13657,N_12044,N_12269);
and U13658 (N_13658,N_12880,N_12866);
xor U13659 (N_13659,N_12068,N_12316);
xor U13660 (N_13660,N_12786,N_12482);
or U13661 (N_13661,N_12446,N_12703);
nor U13662 (N_13662,N_12970,N_12480);
or U13663 (N_13663,N_12183,N_12880);
xnor U13664 (N_13664,N_12050,N_12228);
nor U13665 (N_13665,N_12598,N_12526);
or U13666 (N_13666,N_12422,N_12457);
nor U13667 (N_13667,N_12043,N_12685);
and U13668 (N_13668,N_12875,N_12954);
and U13669 (N_13669,N_12845,N_12156);
nor U13670 (N_13670,N_12990,N_12339);
or U13671 (N_13671,N_12691,N_12750);
and U13672 (N_13672,N_12131,N_12094);
nor U13673 (N_13673,N_12855,N_12413);
and U13674 (N_13674,N_12610,N_12781);
nand U13675 (N_13675,N_12556,N_12759);
nor U13676 (N_13676,N_12110,N_12834);
and U13677 (N_13677,N_12980,N_12253);
nor U13678 (N_13678,N_12479,N_12201);
nor U13679 (N_13679,N_12953,N_12904);
nand U13680 (N_13680,N_12142,N_12209);
and U13681 (N_13681,N_12703,N_12728);
and U13682 (N_13682,N_12538,N_12713);
xor U13683 (N_13683,N_12541,N_12108);
nand U13684 (N_13684,N_12272,N_12295);
nand U13685 (N_13685,N_12517,N_12098);
nor U13686 (N_13686,N_12192,N_12525);
xor U13687 (N_13687,N_12457,N_12037);
or U13688 (N_13688,N_12341,N_12984);
and U13689 (N_13689,N_12170,N_12335);
nand U13690 (N_13690,N_12856,N_12397);
nor U13691 (N_13691,N_12933,N_12878);
nand U13692 (N_13692,N_12477,N_12994);
and U13693 (N_13693,N_12582,N_12316);
or U13694 (N_13694,N_12303,N_12059);
nor U13695 (N_13695,N_12959,N_12432);
nand U13696 (N_13696,N_12063,N_12530);
nor U13697 (N_13697,N_12925,N_12690);
and U13698 (N_13698,N_12840,N_12403);
nand U13699 (N_13699,N_12817,N_12970);
or U13700 (N_13700,N_12755,N_12353);
nand U13701 (N_13701,N_12827,N_12190);
nand U13702 (N_13702,N_12191,N_12530);
xor U13703 (N_13703,N_12723,N_12469);
and U13704 (N_13704,N_12368,N_12307);
nand U13705 (N_13705,N_12292,N_12842);
nand U13706 (N_13706,N_12093,N_12666);
or U13707 (N_13707,N_12486,N_12973);
nand U13708 (N_13708,N_12382,N_12798);
xnor U13709 (N_13709,N_12947,N_12613);
nor U13710 (N_13710,N_12122,N_12831);
xnor U13711 (N_13711,N_12830,N_12112);
nor U13712 (N_13712,N_12973,N_12273);
nand U13713 (N_13713,N_12380,N_12622);
and U13714 (N_13714,N_12549,N_12588);
nor U13715 (N_13715,N_12410,N_12109);
nor U13716 (N_13716,N_12873,N_12896);
or U13717 (N_13717,N_12412,N_12571);
or U13718 (N_13718,N_12470,N_12371);
nor U13719 (N_13719,N_12053,N_12957);
nand U13720 (N_13720,N_12995,N_12484);
and U13721 (N_13721,N_12807,N_12256);
and U13722 (N_13722,N_12635,N_12218);
nand U13723 (N_13723,N_12323,N_12289);
xor U13724 (N_13724,N_12147,N_12412);
nor U13725 (N_13725,N_12055,N_12218);
and U13726 (N_13726,N_12334,N_12458);
and U13727 (N_13727,N_12092,N_12046);
nor U13728 (N_13728,N_12456,N_12178);
and U13729 (N_13729,N_12549,N_12816);
xor U13730 (N_13730,N_12284,N_12187);
nor U13731 (N_13731,N_12547,N_12508);
or U13732 (N_13732,N_12425,N_12182);
or U13733 (N_13733,N_12122,N_12472);
nor U13734 (N_13734,N_12095,N_12125);
and U13735 (N_13735,N_12096,N_12724);
xnor U13736 (N_13736,N_12073,N_12891);
nand U13737 (N_13737,N_12567,N_12775);
xor U13738 (N_13738,N_12728,N_12677);
or U13739 (N_13739,N_12140,N_12381);
or U13740 (N_13740,N_12507,N_12116);
nor U13741 (N_13741,N_12700,N_12514);
xnor U13742 (N_13742,N_12558,N_12603);
nor U13743 (N_13743,N_12512,N_12262);
xnor U13744 (N_13744,N_12906,N_12826);
xor U13745 (N_13745,N_12549,N_12525);
or U13746 (N_13746,N_12717,N_12326);
and U13747 (N_13747,N_12866,N_12720);
xor U13748 (N_13748,N_12778,N_12234);
nor U13749 (N_13749,N_12493,N_12692);
xnor U13750 (N_13750,N_12106,N_12758);
nand U13751 (N_13751,N_12971,N_12714);
xnor U13752 (N_13752,N_12090,N_12905);
nand U13753 (N_13753,N_12604,N_12328);
xor U13754 (N_13754,N_12382,N_12141);
nor U13755 (N_13755,N_12249,N_12272);
and U13756 (N_13756,N_12483,N_12861);
xor U13757 (N_13757,N_12101,N_12276);
nand U13758 (N_13758,N_12169,N_12403);
or U13759 (N_13759,N_12432,N_12255);
or U13760 (N_13760,N_12785,N_12807);
or U13761 (N_13761,N_12963,N_12802);
nand U13762 (N_13762,N_12992,N_12867);
and U13763 (N_13763,N_12034,N_12459);
nor U13764 (N_13764,N_12628,N_12516);
nand U13765 (N_13765,N_12050,N_12977);
or U13766 (N_13766,N_12162,N_12268);
nand U13767 (N_13767,N_12971,N_12013);
or U13768 (N_13768,N_12929,N_12263);
nor U13769 (N_13769,N_12383,N_12039);
nor U13770 (N_13770,N_12419,N_12040);
and U13771 (N_13771,N_12725,N_12694);
or U13772 (N_13772,N_12146,N_12800);
nand U13773 (N_13773,N_12557,N_12769);
nand U13774 (N_13774,N_12689,N_12709);
or U13775 (N_13775,N_12781,N_12319);
and U13776 (N_13776,N_12299,N_12966);
nand U13777 (N_13777,N_12029,N_12462);
xnor U13778 (N_13778,N_12256,N_12833);
or U13779 (N_13779,N_12563,N_12757);
nand U13780 (N_13780,N_12469,N_12770);
nand U13781 (N_13781,N_12678,N_12729);
xor U13782 (N_13782,N_12671,N_12080);
and U13783 (N_13783,N_12819,N_12521);
nand U13784 (N_13784,N_12002,N_12489);
or U13785 (N_13785,N_12577,N_12835);
nor U13786 (N_13786,N_12206,N_12618);
xnor U13787 (N_13787,N_12469,N_12712);
xnor U13788 (N_13788,N_12711,N_12050);
or U13789 (N_13789,N_12450,N_12276);
xnor U13790 (N_13790,N_12353,N_12458);
nand U13791 (N_13791,N_12552,N_12176);
nand U13792 (N_13792,N_12154,N_12774);
and U13793 (N_13793,N_12350,N_12750);
nor U13794 (N_13794,N_12083,N_12941);
and U13795 (N_13795,N_12273,N_12854);
xnor U13796 (N_13796,N_12906,N_12084);
nand U13797 (N_13797,N_12484,N_12629);
nor U13798 (N_13798,N_12791,N_12921);
and U13799 (N_13799,N_12980,N_12586);
and U13800 (N_13800,N_12443,N_12766);
nor U13801 (N_13801,N_12199,N_12830);
or U13802 (N_13802,N_12859,N_12635);
xor U13803 (N_13803,N_12038,N_12607);
nor U13804 (N_13804,N_12284,N_12384);
or U13805 (N_13805,N_12213,N_12307);
xnor U13806 (N_13806,N_12098,N_12364);
nand U13807 (N_13807,N_12718,N_12742);
and U13808 (N_13808,N_12824,N_12765);
and U13809 (N_13809,N_12240,N_12942);
or U13810 (N_13810,N_12114,N_12721);
nand U13811 (N_13811,N_12795,N_12631);
or U13812 (N_13812,N_12102,N_12925);
nand U13813 (N_13813,N_12911,N_12927);
xor U13814 (N_13814,N_12387,N_12983);
nor U13815 (N_13815,N_12318,N_12306);
or U13816 (N_13816,N_12247,N_12542);
or U13817 (N_13817,N_12577,N_12036);
or U13818 (N_13818,N_12986,N_12811);
and U13819 (N_13819,N_12085,N_12500);
xor U13820 (N_13820,N_12794,N_12879);
and U13821 (N_13821,N_12823,N_12502);
xnor U13822 (N_13822,N_12664,N_12912);
nand U13823 (N_13823,N_12921,N_12799);
xnor U13824 (N_13824,N_12450,N_12378);
nor U13825 (N_13825,N_12161,N_12638);
and U13826 (N_13826,N_12928,N_12782);
xnor U13827 (N_13827,N_12876,N_12103);
xor U13828 (N_13828,N_12603,N_12507);
nor U13829 (N_13829,N_12454,N_12244);
nor U13830 (N_13830,N_12067,N_12433);
nand U13831 (N_13831,N_12723,N_12179);
nand U13832 (N_13832,N_12716,N_12596);
xor U13833 (N_13833,N_12323,N_12602);
nor U13834 (N_13834,N_12939,N_12740);
nand U13835 (N_13835,N_12003,N_12477);
nand U13836 (N_13836,N_12538,N_12933);
nor U13837 (N_13837,N_12773,N_12223);
or U13838 (N_13838,N_12226,N_12631);
and U13839 (N_13839,N_12988,N_12143);
and U13840 (N_13840,N_12562,N_12757);
nor U13841 (N_13841,N_12543,N_12467);
nor U13842 (N_13842,N_12831,N_12517);
nor U13843 (N_13843,N_12452,N_12910);
xnor U13844 (N_13844,N_12345,N_12201);
nand U13845 (N_13845,N_12457,N_12642);
nand U13846 (N_13846,N_12585,N_12144);
xor U13847 (N_13847,N_12758,N_12030);
nor U13848 (N_13848,N_12967,N_12289);
or U13849 (N_13849,N_12292,N_12277);
nor U13850 (N_13850,N_12133,N_12183);
nand U13851 (N_13851,N_12711,N_12565);
xor U13852 (N_13852,N_12260,N_12601);
and U13853 (N_13853,N_12170,N_12152);
and U13854 (N_13854,N_12521,N_12596);
or U13855 (N_13855,N_12045,N_12555);
and U13856 (N_13856,N_12220,N_12420);
nor U13857 (N_13857,N_12007,N_12220);
nand U13858 (N_13858,N_12974,N_12534);
xor U13859 (N_13859,N_12359,N_12637);
and U13860 (N_13860,N_12841,N_12711);
xnor U13861 (N_13861,N_12036,N_12823);
xor U13862 (N_13862,N_12432,N_12689);
nand U13863 (N_13863,N_12115,N_12727);
and U13864 (N_13864,N_12740,N_12015);
and U13865 (N_13865,N_12758,N_12163);
nor U13866 (N_13866,N_12077,N_12778);
and U13867 (N_13867,N_12998,N_12228);
and U13868 (N_13868,N_12270,N_12729);
nand U13869 (N_13869,N_12394,N_12600);
xor U13870 (N_13870,N_12510,N_12212);
or U13871 (N_13871,N_12608,N_12584);
and U13872 (N_13872,N_12100,N_12713);
nand U13873 (N_13873,N_12035,N_12198);
xnor U13874 (N_13874,N_12346,N_12440);
nand U13875 (N_13875,N_12269,N_12153);
nor U13876 (N_13876,N_12912,N_12368);
or U13877 (N_13877,N_12809,N_12279);
nor U13878 (N_13878,N_12728,N_12031);
xnor U13879 (N_13879,N_12612,N_12348);
nand U13880 (N_13880,N_12249,N_12458);
xor U13881 (N_13881,N_12133,N_12843);
nand U13882 (N_13882,N_12665,N_12758);
xor U13883 (N_13883,N_12943,N_12437);
xor U13884 (N_13884,N_12356,N_12208);
nor U13885 (N_13885,N_12043,N_12866);
nor U13886 (N_13886,N_12370,N_12469);
nand U13887 (N_13887,N_12540,N_12293);
and U13888 (N_13888,N_12886,N_12101);
or U13889 (N_13889,N_12255,N_12584);
nor U13890 (N_13890,N_12592,N_12543);
or U13891 (N_13891,N_12215,N_12226);
or U13892 (N_13892,N_12095,N_12210);
nor U13893 (N_13893,N_12239,N_12837);
nor U13894 (N_13894,N_12965,N_12094);
nand U13895 (N_13895,N_12574,N_12567);
xnor U13896 (N_13896,N_12580,N_12428);
or U13897 (N_13897,N_12291,N_12877);
nand U13898 (N_13898,N_12444,N_12324);
nor U13899 (N_13899,N_12407,N_12392);
nand U13900 (N_13900,N_12221,N_12796);
nor U13901 (N_13901,N_12473,N_12074);
or U13902 (N_13902,N_12414,N_12757);
and U13903 (N_13903,N_12814,N_12609);
nor U13904 (N_13904,N_12561,N_12736);
xor U13905 (N_13905,N_12389,N_12170);
xor U13906 (N_13906,N_12210,N_12714);
xnor U13907 (N_13907,N_12286,N_12303);
or U13908 (N_13908,N_12356,N_12744);
nor U13909 (N_13909,N_12336,N_12374);
or U13910 (N_13910,N_12592,N_12850);
xnor U13911 (N_13911,N_12900,N_12507);
and U13912 (N_13912,N_12737,N_12560);
and U13913 (N_13913,N_12124,N_12806);
xnor U13914 (N_13914,N_12422,N_12145);
xnor U13915 (N_13915,N_12143,N_12557);
and U13916 (N_13916,N_12020,N_12872);
or U13917 (N_13917,N_12632,N_12654);
and U13918 (N_13918,N_12756,N_12216);
nand U13919 (N_13919,N_12739,N_12263);
and U13920 (N_13920,N_12265,N_12185);
nor U13921 (N_13921,N_12157,N_12810);
xnor U13922 (N_13922,N_12491,N_12068);
nor U13923 (N_13923,N_12425,N_12385);
nor U13924 (N_13924,N_12146,N_12343);
and U13925 (N_13925,N_12553,N_12158);
nand U13926 (N_13926,N_12369,N_12716);
and U13927 (N_13927,N_12119,N_12257);
xnor U13928 (N_13928,N_12058,N_12432);
and U13929 (N_13929,N_12365,N_12854);
xnor U13930 (N_13930,N_12329,N_12448);
nand U13931 (N_13931,N_12675,N_12026);
nand U13932 (N_13932,N_12658,N_12153);
nor U13933 (N_13933,N_12164,N_12419);
nor U13934 (N_13934,N_12477,N_12568);
and U13935 (N_13935,N_12802,N_12605);
nand U13936 (N_13936,N_12932,N_12983);
and U13937 (N_13937,N_12908,N_12903);
xnor U13938 (N_13938,N_12860,N_12257);
or U13939 (N_13939,N_12535,N_12915);
nor U13940 (N_13940,N_12810,N_12028);
nor U13941 (N_13941,N_12016,N_12850);
or U13942 (N_13942,N_12511,N_12150);
xnor U13943 (N_13943,N_12174,N_12813);
and U13944 (N_13944,N_12953,N_12658);
xor U13945 (N_13945,N_12265,N_12408);
nand U13946 (N_13946,N_12736,N_12556);
nor U13947 (N_13947,N_12960,N_12803);
xnor U13948 (N_13948,N_12441,N_12249);
xor U13949 (N_13949,N_12137,N_12138);
nand U13950 (N_13950,N_12312,N_12893);
or U13951 (N_13951,N_12124,N_12530);
and U13952 (N_13952,N_12657,N_12037);
and U13953 (N_13953,N_12082,N_12639);
nand U13954 (N_13954,N_12104,N_12190);
and U13955 (N_13955,N_12167,N_12555);
nor U13956 (N_13956,N_12466,N_12967);
or U13957 (N_13957,N_12558,N_12871);
nor U13958 (N_13958,N_12705,N_12434);
or U13959 (N_13959,N_12711,N_12133);
nor U13960 (N_13960,N_12581,N_12029);
and U13961 (N_13961,N_12608,N_12336);
and U13962 (N_13962,N_12121,N_12254);
nand U13963 (N_13963,N_12852,N_12033);
or U13964 (N_13964,N_12052,N_12943);
nand U13965 (N_13965,N_12672,N_12964);
nor U13966 (N_13966,N_12156,N_12688);
nand U13967 (N_13967,N_12393,N_12101);
xnor U13968 (N_13968,N_12996,N_12647);
nand U13969 (N_13969,N_12089,N_12627);
or U13970 (N_13970,N_12143,N_12966);
and U13971 (N_13971,N_12280,N_12936);
nand U13972 (N_13972,N_12680,N_12229);
or U13973 (N_13973,N_12962,N_12077);
nor U13974 (N_13974,N_12325,N_12236);
xor U13975 (N_13975,N_12909,N_12134);
and U13976 (N_13976,N_12297,N_12003);
or U13977 (N_13977,N_12583,N_12484);
nor U13978 (N_13978,N_12368,N_12005);
nand U13979 (N_13979,N_12559,N_12692);
xnor U13980 (N_13980,N_12431,N_12688);
or U13981 (N_13981,N_12941,N_12955);
xnor U13982 (N_13982,N_12038,N_12492);
and U13983 (N_13983,N_12309,N_12187);
nor U13984 (N_13984,N_12483,N_12688);
xnor U13985 (N_13985,N_12926,N_12665);
and U13986 (N_13986,N_12508,N_12372);
nor U13987 (N_13987,N_12041,N_12204);
xor U13988 (N_13988,N_12535,N_12313);
and U13989 (N_13989,N_12358,N_12678);
and U13990 (N_13990,N_12233,N_12148);
nand U13991 (N_13991,N_12834,N_12630);
or U13992 (N_13992,N_12548,N_12212);
nand U13993 (N_13993,N_12896,N_12312);
and U13994 (N_13994,N_12684,N_12933);
or U13995 (N_13995,N_12383,N_12311);
xor U13996 (N_13996,N_12208,N_12160);
xor U13997 (N_13997,N_12618,N_12011);
xor U13998 (N_13998,N_12442,N_12819);
nand U13999 (N_13999,N_12580,N_12595);
nor U14000 (N_14000,N_13176,N_13602);
xor U14001 (N_14001,N_13717,N_13845);
and U14002 (N_14002,N_13023,N_13801);
and U14003 (N_14003,N_13368,N_13103);
nand U14004 (N_14004,N_13210,N_13946);
nor U14005 (N_14005,N_13991,N_13314);
nor U14006 (N_14006,N_13609,N_13182);
xnor U14007 (N_14007,N_13365,N_13100);
nand U14008 (N_14008,N_13105,N_13578);
or U14009 (N_14009,N_13400,N_13265);
nor U14010 (N_14010,N_13215,N_13852);
and U14011 (N_14011,N_13833,N_13360);
and U14012 (N_14012,N_13567,N_13158);
nand U14013 (N_14013,N_13923,N_13018);
or U14014 (N_14014,N_13788,N_13795);
xor U14015 (N_14015,N_13524,N_13255);
xor U14016 (N_14016,N_13986,N_13559);
or U14017 (N_14017,N_13597,N_13995);
or U14018 (N_14018,N_13543,N_13114);
or U14019 (N_14019,N_13761,N_13247);
nand U14020 (N_14020,N_13618,N_13814);
and U14021 (N_14021,N_13532,N_13726);
nor U14022 (N_14022,N_13202,N_13841);
or U14023 (N_14023,N_13533,N_13498);
nor U14024 (N_14024,N_13044,N_13475);
or U14025 (N_14025,N_13484,N_13929);
nand U14026 (N_14026,N_13953,N_13507);
xnor U14027 (N_14027,N_13061,N_13428);
nand U14028 (N_14028,N_13245,N_13577);
xor U14029 (N_14029,N_13350,N_13846);
or U14030 (N_14030,N_13718,N_13009);
and U14031 (N_14031,N_13536,N_13779);
and U14032 (N_14032,N_13756,N_13093);
or U14033 (N_14033,N_13207,N_13688);
or U14034 (N_14034,N_13312,N_13440);
or U14035 (N_14035,N_13831,N_13563);
or U14036 (N_14036,N_13727,N_13722);
or U14037 (N_14037,N_13931,N_13861);
and U14038 (N_14038,N_13917,N_13031);
or U14039 (N_14039,N_13519,N_13523);
nand U14040 (N_14040,N_13141,N_13414);
nor U14041 (N_14041,N_13555,N_13998);
nor U14042 (N_14042,N_13467,N_13634);
xnor U14043 (N_14043,N_13449,N_13893);
nor U14044 (N_14044,N_13283,N_13878);
nor U14045 (N_14045,N_13910,N_13308);
and U14046 (N_14046,N_13331,N_13102);
nor U14047 (N_14047,N_13035,N_13216);
nand U14048 (N_14048,N_13104,N_13352);
xnor U14049 (N_14049,N_13032,N_13847);
and U14050 (N_14050,N_13388,N_13270);
and U14051 (N_14051,N_13658,N_13698);
nor U14052 (N_14052,N_13479,N_13074);
nand U14053 (N_14053,N_13159,N_13227);
or U14054 (N_14054,N_13313,N_13180);
nor U14055 (N_14055,N_13941,N_13165);
nor U14056 (N_14056,N_13939,N_13754);
nor U14057 (N_14057,N_13005,N_13167);
nor U14058 (N_14058,N_13154,N_13059);
and U14059 (N_14059,N_13204,N_13126);
nand U14060 (N_14060,N_13990,N_13709);
nand U14061 (N_14061,N_13409,N_13284);
nor U14062 (N_14062,N_13427,N_13072);
xnor U14063 (N_14063,N_13266,N_13592);
xor U14064 (N_14064,N_13209,N_13144);
nand U14065 (N_14065,N_13511,N_13193);
and U14066 (N_14066,N_13208,N_13187);
and U14067 (N_14067,N_13915,N_13936);
or U14068 (N_14068,N_13185,N_13371);
and U14069 (N_14069,N_13836,N_13025);
nand U14070 (N_14070,N_13528,N_13684);
xnor U14071 (N_14071,N_13812,N_13904);
xor U14072 (N_14072,N_13046,N_13478);
or U14073 (N_14073,N_13913,N_13951);
nor U14074 (N_14074,N_13197,N_13014);
nor U14075 (N_14075,N_13062,N_13749);
nand U14076 (N_14076,N_13622,N_13225);
xor U14077 (N_14077,N_13049,N_13224);
nor U14078 (N_14078,N_13610,N_13474);
xnor U14079 (N_14079,N_13260,N_13254);
nand U14080 (N_14080,N_13891,N_13367);
and U14081 (N_14081,N_13562,N_13963);
xnor U14082 (N_14082,N_13462,N_13730);
xnor U14083 (N_14083,N_13175,N_13095);
xor U14084 (N_14084,N_13908,N_13199);
nor U14085 (N_14085,N_13506,N_13097);
nor U14086 (N_14086,N_13304,N_13011);
and U14087 (N_14087,N_13540,N_13526);
or U14088 (N_14088,N_13439,N_13047);
nand U14089 (N_14089,N_13601,N_13529);
nor U14090 (N_14090,N_13520,N_13111);
and U14091 (N_14091,N_13583,N_13614);
and U14092 (N_14092,N_13599,N_13735);
xor U14093 (N_14093,N_13616,N_13110);
or U14094 (N_14094,N_13556,N_13465);
xor U14095 (N_14095,N_13576,N_13066);
or U14096 (N_14096,N_13553,N_13586);
and U14097 (N_14097,N_13333,N_13402);
nand U14098 (N_14098,N_13149,N_13504);
or U14099 (N_14099,N_13564,N_13223);
nor U14100 (N_14100,N_13890,N_13685);
or U14101 (N_14101,N_13274,N_13017);
nor U14102 (N_14102,N_13826,N_13054);
or U14103 (N_14103,N_13045,N_13594);
nor U14104 (N_14104,N_13593,N_13243);
and U14105 (N_14105,N_13920,N_13370);
and U14106 (N_14106,N_13748,N_13143);
and U14107 (N_14107,N_13067,N_13821);
or U14108 (N_14108,N_13390,N_13757);
xor U14109 (N_14109,N_13220,N_13870);
nor U14110 (N_14110,N_13644,N_13418);
nand U14111 (N_14111,N_13747,N_13482);
or U14112 (N_14112,N_13179,N_13300);
nand U14113 (N_14113,N_13026,N_13119);
nor U14114 (N_14114,N_13437,N_13898);
or U14115 (N_14115,N_13447,N_13956);
nor U14116 (N_14116,N_13868,N_13959);
xnor U14117 (N_14117,N_13369,N_13935);
nor U14118 (N_14118,N_13573,N_13509);
nand U14119 (N_14119,N_13030,N_13854);
nor U14120 (N_14120,N_13560,N_13171);
nor U14121 (N_14121,N_13420,N_13800);
xor U14122 (N_14122,N_13706,N_13351);
and U14123 (N_14123,N_13569,N_13161);
or U14124 (N_14124,N_13774,N_13137);
nand U14125 (N_14125,N_13292,N_13505);
nor U14126 (N_14126,N_13226,N_13624);
xnor U14127 (N_14127,N_13436,N_13106);
or U14128 (N_14128,N_13911,N_13169);
nor U14129 (N_14129,N_13799,N_13746);
and U14130 (N_14130,N_13163,N_13872);
or U14131 (N_14131,N_13636,N_13200);
xor U14132 (N_14132,N_13446,N_13278);
or U14133 (N_14133,N_13002,N_13679);
nor U14134 (N_14134,N_13130,N_13117);
nand U14135 (N_14135,N_13968,N_13924);
and U14136 (N_14136,N_13358,N_13321);
or U14137 (N_14137,N_13584,N_13147);
nand U14138 (N_14138,N_13455,N_13612);
nor U14139 (N_14139,N_13639,N_13464);
nand U14140 (N_14140,N_13345,N_13548);
and U14141 (N_14141,N_13269,N_13557);
nor U14142 (N_14142,N_13109,N_13192);
nand U14143 (N_14143,N_13060,N_13849);
nor U14144 (N_14144,N_13327,N_13785);
or U14145 (N_14145,N_13606,N_13250);
xor U14146 (N_14146,N_13804,N_13657);
or U14147 (N_14147,N_13793,N_13568);
xor U14148 (N_14148,N_13377,N_13297);
and U14149 (N_14149,N_13604,N_13443);
nand U14150 (N_14150,N_13306,N_13751);
nand U14151 (N_14151,N_13319,N_13947);
nor U14152 (N_14152,N_13320,N_13252);
nor U14153 (N_14153,N_13654,N_13448);
nand U14154 (N_14154,N_13912,N_13670);
xor U14155 (N_14155,N_13767,N_13867);
or U14156 (N_14156,N_13595,N_13512);
and U14157 (N_14157,N_13582,N_13473);
xnor U14158 (N_14158,N_13128,N_13777);
and U14159 (N_14159,N_13261,N_13340);
nand U14160 (N_14160,N_13281,N_13343);
nor U14161 (N_14161,N_13974,N_13806);
and U14162 (N_14162,N_13715,N_13457);
nor U14163 (N_14163,N_13240,N_13961);
and U14164 (N_14164,N_13234,N_13742);
and U14165 (N_14165,N_13900,N_13949);
xnor U14166 (N_14166,N_13571,N_13937);
nand U14167 (N_14167,N_13655,N_13286);
or U14168 (N_14168,N_13164,N_13088);
and U14169 (N_14169,N_13431,N_13662);
nand U14170 (N_14170,N_13079,N_13708);
or U14171 (N_14171,N_13648,N_13729);
and U14172 (N_14172,N_13213,N_13676);
nand U14173 (N_14173,N_13982,N_13663);
or U14174 (N_14174,N_13877,N_13395);
xor U14175 (N_14175,N_13341,N_13162);
nor U14176 (N_14176,N_13071,N_13914);
nor U14177 (N_14177,N_13862,N_13098);
xor U14178 (N_14178,N_13116,N_13084);
and U14179 (N_14179,N_13289,N_13744);
and U14180 (N_14180,N_13426,N_13246);
nor U14181 (N_14181,N_13613,N_13191);
nor U14182 (N_14182,N_13019,N_13627);
or U14183 (N_14183,N_13642,N_13575);
and U14184 (N_14184,N_13096,N_13514);
and U14185 (N_14185,N_13127,N_13769);
nand U14186 (N_14186,N_13775,N_13768);
and U14187 (N_14187,N_13628,N_13166);
nor U14188 (N_14188,N_13285,N_13791);
or U14189 (N_14189,N_13605,N_13419);
or U14190 (N_14190,N_13535,N_13256);
and U14191 (N_14191,N_13660,N_13992);
nor U14192 (N_14192,N_13386,N_13083);
xor U14193 (N_14193,N_13344,N_13554);
nand U14194 (N_14194,N_13871,N_13064);
or U14195 (N_14195,N_13690,N_13356);
nor U14196 (N_14196,N_13203,N_13652);
and U14197 (N_14197,N_13566,N_13134);
xor U14198 (N_14198,N_13725,N_13024);
and U14199 (N_14199,N_13491,N_13295);
or U14200 (N_14200,N_13374,N_13434);
and U14201 (N_14201,N_13058,N_13043);
or U14202 (N_14202,N_13750,N_13829);
or U14203 (N_14203,N_13771,N_13010);
nor U14204 (N_14204,N_13808,N_13691);
or U14205 (N_14205,N_13411,N_13268);
nand U14206 (N_14206,N_13952,N_13766);
xnor U14207 (N_14207,N_13036,N_13922);
nor U14208 (N_14208,N_13056,N_13787);
nand U14209 (N_14209,N_13136,N_13738);
nor U14210 (N_14210,N_13206,N_13373);
or U14211 (N_14211,N_13013,N_13581);
or U14212 (N_14212,N_13955,N_13415);
or U14213 (N_14213,N_13493,N_13675);
or U14214 (N_14214,N_13460,N_13550);
nand U14215 (N_14215,N_13611,N_13291);
nor U14216 (N_14216,N_13485,N_13112);
nor U14217 (N_14217,N_13723,N_13970);
xnor U14218 (N_14218,N_13432,N_13755);
or U14219 (N_14219,N_13632,N_13971);
or U14220 (N_14220,N_13542,N_13902);
nand U14221 (N_14221,N_13865,N_13943);
or U14222 (N_14222,N_13444,N_13840);
or U14223 (N_14223,N_13076,N_13366);
xor U14224 (N_14224,N_13063,N_13873);
or U14225 (N_14225,N_13468,N_13324);
and U14226 (N_14226,N_13489,N_13701);
nor U14227 (N_14227,N_13790,N_13798);
xor U14228 (N_14228,N_13574,N_13471);
xor U14229 (N_14229,N_13521,N_13733);
nand U14230 (N_14230,N_13338,N_13229);
xor U14231 (N_14231,N_13572,N_13993);
or U14232 (N_14232,N_13710,N_13681);
and U14233 (N_14233,N_13170,N_13525);
and U14234 (N_14234,N_13359,N_13894);
nand U14235 (N_14235,N_13195,N_13828);
and U14236 (N_14236,N_13570,N_13101);
xor U14237 (N_14237,N_13299,N_13490);
and U14238 (N_14238,N_13976,N_13728);
nor U14239 (N_14239,N_13687,N_13153);
and U14240 (N_14240,N_13824,N_13629);
nand U14241 (N_14241,N_13231,N_13837);
or U14242 (N_14242,N_13277,N_13353);
xnor U14243 (N_14243,N_13355,N_13541);
and U14244 (N_14244,N_13092,N_13714);
or U14245 (N_14245,N_13740,N_13089);
or U14246 (N_14246,N_13819,N_13905);
xnor U14247 (N_14247,N_13934,N_13587);
xnor U14248 (N_14248,N_13930,N_13672);
nand U14249 (N_14249,N_13421,N_13052);
xnor U14250 (N_14250,N_13822,N_13965);
or U14251 (N_14251,N_13707,N_13596);
xnor U14252 (N_14252,N_13181,N_13864);
or U14253 (N_14253,N_13860,N_13157);
nand U14254 (N_14254,N_13977,N_13219);
nor U14255 (N_14255,N_13385,N_13659);
xor U14256 (N_14256,N_13760,N_13372);
xor U14257 (N_14257,N_13481,N_13118);
nor U14258 (N_14258,N_13038,N_13441);
or U14259 (N_14259,N_13194,N_13236);
or U14260 (N_14260,N_13085,N_13257);
or U14261 (N_14261,N_13070,N_13451);
xor U14262 (N_14262,N_13183,N_13459);
nand U14263 (N_14263,N_13336,N_13450);
xor U14264 (N_14264,N_13619,N_13736);
and U14265 (N_14265,N_13994,N_13073);
nand U14266 (N_14266,N_13713,N_13416);
nand U14267 (N_14267,N_13552,N_13262);
nor U14268 (N_14268,N_13695,N_13919);
xnor U14269 (N_14269,N_13656,N_13325);
xnor U14270 (N_14270,N_13724,N_13522);
and U14271 (N_14271,N_13699,N_13809);
nor U14272 (N_14272,N_13813,N_13326);
nor U14273 (N_14273,N_13680,N_13899);
or U14274 (N_14274,N_13702,N_13518);
xnor U14275 (N_14275,N_13410,N_13925);
xnor U14276 (N_14276,N_13916,N_13499);
xnor U14277 (N_14277,N_13907,N_13739);
nor U14278 (N_14278,N_13394,N_13121);
and U14279 (N_14279,N_13776,N_13335);
xnor U14280 (N_14280,N_13721,N_13667);
xor U14281 (N_14281,N_13381,N_13461);
nor U14282 (N_14282,N_13731,N_13984);
nor U14283 (N_14283,N_13275,N_13686);
nand U14284 (N_14284,N_13591,N_13682);
and U14285 (N_14285,N_13753,N_13362);
nor U14286 (N_14286,N_13758,N_13762);
and U14287 (N_14287,N_13933,N_13510);
nor U14288 (N_14288,N_13770,N_13807);
xor U14289 (N_14289,N_13081,N_13830);
nor U14290 (N_14290,N_13323,N_13034);
and U14291 (N_14291,N_13888,N_13389);
nor U14292 (N_14292,N_13501,N_13080);
xor U14293 (N_14293,N_13856,N_13957);
nand U14294 (N_14294,N_13232,N_13021);
nor U14295 (N_14295,N_13875,N_13703);
and U14296 (N_14296,N_13408,N_13029);
nor U14297 (N_14297,N_13950,N_13580);
or U14298 (N_14298,N_13012,N_13361);
or U14299 (N_14299,N_13508,N_13780);
or U14300 (N_14300,N_13789,N_13942);
or U14301 (N_14301,N_13138,N_13810);
and U14302 (N_14302,N_13413,N_13983);
xnor U14303 (N_14303,N_13665,N_13453);
nand U14304 (N_14304,N_13981,N_13125);
xor U14305 (N_14305,N_13889,N_13772);
xnor U14306 (N_14306,N_13228,N_13339);
xor U14307 (N_14307,N_13895,N_13832);
nand U14308 (N_14308,N_13198,N_13075);
and U14309 (N_14309,N_13328,N_13188);
and U14310 (N_14310,N_13235,N_13458);
xor U14311 (N_14311,N_13332,N_13272);
xnor U14312 (N_14312,N_13178,N_13743);
or U14313 (N_14313,N_13705,N_13752);
nor U14314 (N_14314,N_13122,N_13040);
xnor U14315 (N_14315,N_13851,N_13823);
nor U14316 (N_14316,N_13405,N_13435);
xor U14317 (N_14317,N_13671,N_13996);
xnor U14318 (N_14318,N_13940,N_13892);
or U14319 (N_14319,N_13763,N_13249);
xnor U14320 (N_14320,N_13466,N_13379);
or U14321 (N_14321,N_13142,N_13091);
or U14322 (N_14322,N_13588,N_13668);
xor U14323 (N_14323,N_13082,N_13885);
and U14324 (N_14324,N_13839,N_13692);
xnor U14325 (N_14325,N_13843,N_13078);
xnor U14326 (N_14326,N_13927,N_13649);
nand U14327 (N_14327,N_13302,N_13975);
nand U14328 (N_14328,N_13330,N_13069);
nor U14329 (N_14329,N_13003,N_13589);
or U14330 (N_14330,N_13797,N_13494);
and U14331 (N_14331,N_13781,N_13544);
or U14332 (N_14332,N_13293,N_13719);
and U14333 (N_14333,N_13425,N_13879);
xnor U14334 (N_14334,N_13863,N_13251);
xnor U14335 (N_14335,N_13384,N_13697);
nand U14336 (N_14336,N_13623,N_13190);
or U14337 (N_14337,N_13653,N_13186);
nor U14338 (N_14338,N_13683,N_13357);
xor U14339 (N_14339,N_13039,N_13664);
and U14340 (N_14340,N_13311,N_13999);
nand U14341 (N_14341,N_13346,N_13932);
nand U14342 (N_14342,N_13666,N_13057);
nand U14343 (N_14343,N_13579,N_13967);
nand U14344 (N_14344,N_13997,N_13124);
nand U14345 (N_14345,N_13383,N_13037);
or U14346 (N_14346,N_13786,N_13015);
nand U14347 (N_14347,N_13259,N_13438);
or U14348 (N_14348,N_13267,N_13537);
and U14349 (N_14349,N_13765,N_13886);
nor U14350 (N_14350,N_13094,N_13217);
xnor U14351 (N_14351,N_13620,N_13041);
nand U14352 (N_14352,N_13398,N_13033);
or U14353 (N_14353,N_13741,N_13241);
xnor U14354 (N_14354,N_13551,N_13316);
nand U14355 (N_14355,N_13637,N_13315);
nand U14356 (N_14356,N_13113,N_13641);
nand U14357 (N_14357,N_13174,N_13380);
nand U14358 (N_14358,N_13387,N_13486);
and U14359 (N_14359,N_13638,N_13347);
nand U14360 (N_14360,N_13423,N_13858);
nand U14361 (N_14361,N_13784,N_13603);
and U14362 (N_14362,N_13816,N_13087);
xor U14363 (N_14363,N_13237,N_13640);
nor U14364 (N_14364,N_13500,N_13042);
and U14365 (N_14365,N_13962,N_13090);
and U14366 (N_14366,N_13711,N_13201);
and U14367 (N_14367,N_13244,N_13310);
nor U14368 (N_14368,N_13463,N_13276);
and U14369 (N_14369,N_13483,N_13973);
or U14370 (N_14370,N_13318,N_13303);
or U14371 (N_14371,N_13884,N_13549);
and U14372 (N_14372,N_13492,N_13792);
nor U14373 (N_14373,N_13869,N_13205);
nor U14374 (N_14374,N_13513,N_13631);
or U14375 (N_14375,N_13155,N_13972);
and U14376 (N_14376,N_13527,N_13131);
xor U14377 (N_14377,N_13337,N_13397);
or U14378 (N_14378,N_13887,N_13349);
nand U14379 (N_14379,N_13647,N_13253);
nor U14380 (N_14380,N_13827,N_13737);
xnor U14381 (N_14381,N_13516,N_13329);
nand U14382 (N_14382,N_13608,N_13317);
and U14383 (N_14383,N_13053,N_13348);
nor U14384 (N_14384,N_13001,N_13979);
nand U14385 (N_14385,N_13375,N_13517);
or U14386 (N_14386,N_13048,N_13600);
nor U14387 (N_14387,N_13298,N_13433);
nand U14388 (N_14388,N_13248,N_13148);
nand U14389 (N_14389,N_13403,N_13077);
nor U14390 (N_14390,N_13838,N_13065);
or U14391 (N_14391,N_13987,N_13626);
or U14392 (N_14392,N_13538,N_13835);
nand U14393 (N_14393,N_13534,N_13086);
nor U14394 (N_14394,N_13720,N_13222);
xor U14395 (N_14395,N_13734,N_13857);
nor U14396 (N_14396,N_13363,N_13883);
nand U14397 (N_14397,N_13944,N_13264);
or U14398 (N_14398,N_13123,N_13545);
nand U14399 (N_14399,N_13099,N_13497);
or U14400 (N_14400,N_13704,N_13133);
xor U14401 (N_14401,N_13442,N_13590);
xnor U14402 (N_14402,N_13016,N_13495);
or U14403 (N_14403,N_13271,N_13108);
nor U14404 (N_14404,N_13146,N_13669);
xor U14405 (N_14405,N_13004,N_13547);
nand U14406 (N_14406,N_13980,N_13239);
or U14407 (N_14407,N_13661,N_13173);
and U14408 (N_14408,N_13759,N_13646);
or U14409 (N_14409,N_13565,N_13429);
or U14410 (N_14410,N_13635,N_13896);
or U14411 (N_14411,N_13782,N_13853);
or U14412 (N_14412,N_13151,N_13152);
and U14413 (N_14413,N_13392,N_13470);
nor U14414 (N_14414,N_13211,N_13844);
or U14415 (N_14415,N_13585,N_13909);
and U14416 (N_14416,N_13643,N_13160);
xor U14417 (N_14417,N_13645,N_13145);
xnor U14418 (N_14418,N_13184,N_13530);
xor U14419 (N_14419,N_13617,N_13258);
nand U14420 (N_14420,N_13928,N_13903);
or U14421 (N_14421,N_13906,N_13630);
nand U14422 (N_14422,N_13918,N_13140);
or U14423 (N_14423,N_13796,N_13539);
xnor U14424 (N_14424,N_13156,N_13694);
or U14425 (N_14425,N_13818,N_13783);
nor U14426 (N_14426,N_13794,N_13382);
xor U14427 (N_14427,N_13399,N_13135);
nor U14428 (N_14428,N_13007,N_13051);
nor U14429 (N_14429,N_13238,N_13027);
or U14430 (N_14430,N_13712,N_13825);
and U14431 (N_14431,N_13633,N_13454);
nand U14432 (N_14432,N_13120,N_13678);
nand U14433 (N_14433,N_13288,N_13496);
nand U14434 (N_14434,N_13006,N_13848);
nand U14435 (N_14435,N_13716,N_13817);
nor U14436 (N_14436,N_13700,N_13212);
nor U14437 (N_14437,N_13938,N_13650);
nand U14438 (N_14438,N_13988,N_13850);
nand U14439 (N_14439,N_13502,N_13515);
nand U14440 (N_14440,N_13764,N_13301);
xor U14441 (N_14441,N_13000,N_13693);
or U14442 (N_14442,N_13901,N_13958);
nand U14443 (N_14443,N_13842,N_13354);
nand U14444 (N_14444,N_13621,N_13218);
nand U14445 (N_14445,N_13874,N_13598);
xnor U14446 (N_14446,N_13803,N_13815);
nand U14447 (N_14447,N_13342,N_13778);
and U14448 (N_14448,N_13615,N_13773);
or U14449 (N_14449,N_13309,N_13745);
or U14450 (N_14450,N_13811,N_13150);
or U14451 (N_14451,N_13926,N_13050);
or U14452 (N_14452,N_13921,N_13673);
xnor U14453 (N_14453,N_13290,N_13948);
xor U14454 (N_14454,N_13214,N_13294);
and U14455 (N_14455,N_13456,N_13503);
or U14456 (N_14456,N_13978,N_13008);
xnor U14457 (N_14457,N_13531,N_13396);
or U14458 (N_14458,N_13985,N_13625);
nor U14459 (N_14459,N_13859,N_13954);
nand U14460 (N_14460,N_13376,N_13282);
nand U14461 (N_14461,N_13558,N_13412);
or U14462 (N_14462,N_13487,N_13055);
xor U14463 (N_14463,N_13401,N_13732);
and U14464 (N_14464,N_13488,N_13689);
xor U14465 (N_14465,N_13334,N_13422);
nor U14466 (N_14466,N_13280,N_13022);
nand U14467 (N_14467,N_13445,N_13305);
nor U14468 (N_14468,N_13139,N_13263);
and U14469 (N_14469,N_13452,N_13273);
nor U14470 (N_14470,N_13855,N_13651);
or U14471 (N_14471,N_13897,N_13028);
or U14472 (N_14472,N_13674,N_13391);
nand U14473 (N_14473,N_13881,N_13424);
and U14474 (N_14474,N_13802,N_13322);
nand U14475 (N_14475,N_13172,N_13196);
xnor U14476 (N_14476,N_13230,N_13960);
nand U14477 (N_14477,N_13546,N_13677);
xnor U14478 (N_14478,N_13296,N_13472);
and U14479 (N_14479,N_13696,N_13876);
or U14480 (N_14480,N_13287,N_13307);
nor U14481 (N_14481,N_13430,N_13834);
and U14482 (N_14482,N_13020,N_13964);
nor U14483 (N_14483,N_13805,N_13561);
xnor U14484 (N_14484,N_13469,N_13221);
nand U14485 (N_14485,N_13406,N_13945);
and U14486 (N_14486,N_13364,N_13068);
nor U14487 (N_14487,N_13129,N_13107);
and U14488 (N_14488,N_13242,N_13477);
and U14489 (N_14489,N_13393,N_13115);
and U14490 (N_14490,N_13882,N_13866);
xnor U14491 (N_14491,N_13407,N_13168);
nand U14492 (N_14492,N_13177,N_13233);
xnor U14493 (N_14493,N_13820,N_13404);
and U14494 (N_14494,N_13969,N_13378);
xnor U14495 (N_14495,N_13880,N_13476);
xor U14496 (N_14496,N_13966,N_13480);
nand U14497 (N_14497,N_13417,N_13989);
and U14498 (N_14498,N_13607,N_13132);
and U14499 (N_14499,N_13189,N_13279);
or U14500 (N_14500,N_13164,N_13406);
or U14501 (N_14501,N_13221,N_13629);
and U14502 (N_14502,N_13836,N_13430);
and U14503 (N_14503,N_13970,N_13749);
and U14504 (N_14504,N_13299,N_13542);
and U14505 (N_14505,N_13214,N_13222);
or U14506 (N_14506,N_13188,N_13737);
nor U14507 (N_14507,N_13948,N_13635);
or U14508 (N_14508,N_13307,N_13993);
or U14509 (N_14509,N_13754,N_13809);
nand U14510 (N_14510,N_13216,N_13492);
nor U14511 (N_14511,N_13623,N_13822);
and U14512 (N_14512,N_13846,N_13427);
xor U14513 (N_14513,N_13099,N_13820);
xor U14514 (N_14514,N_13050,N_13882);
nand U14515 (N_14515,N_13970,N_13853);
nand U14516 (N_14516,N_13642,N_13196);
xor U14517 (N_14517,N_13665,N_13210);
and U14518 (N_14518,N_13985,N_13982);
and U14519 (N_14519,N_13863,N_13189);
and U14520 (N_14520,N_13520,N_13214);
xor U14521 (N_14521,N_13688,N_13416);
and U14522 (N_14522,N_13195,N_13239);
nor U14523 (N_14523,N_13910,N_13323);
nand U14524 (N_14524,N_13675,N_13977);
nand U14525 (N_14525,N_13197,N_13321);
and U14526 (N_14526,N_13292,N_13311);
nor U14527 (N_14527,N_13280,N_13483);
nor U14528 (N_14528,N_13305,N_13657);
or U14529 (N_14529,N_13839,N_13775);
nor U14530 (N_14530,N_13257,N_13272);
nor U14531 (N_14531,N_13089,N_13769);
xnor U14532 (N_14532,N_13683,N_13259);
nand U14533 (N_14533,N_13750,N_13223);
nor U14534 (N_14534,N_13971,N_13135);
xor U14535 (N_14535,N_13889,N_13253);
and U14536 (N_14536,N_13475,N_13966);
and U14537 (N_14537,N_13571,N_13698);
nand U14538 (N_14538,N_13532,N_13393);
nand U14539 (N_14539,N_13752,N_13479);
and U14540 (N_14540,N_13285,N_13429);
xnor U14541 (N_14541,N_13921,N_13499);
nand U14542 (N_14542,N_13414,N_13485);
xor U14543 (N_14543,N_13451,N_13682);
or U14544 (N_14544,N_13938,N_13415);
nor U14545 (N_14545,N_13612,N_13095);
and U14546 (N_14546,N_13229,N_13378);
xor U14547 (N_14547,N_13168,N_13152);
nor U14548 (N_14548,N_13315,N_13324);
and U14549 (N_14549,N_13307,N_13290);
nand U14550 (N_14550,N_13903,N_13915);
or U14551 (N_14551,N_13963,N_13178);
xnor U14552 (N_14552,N_13471,N_13677);
or U14553 (N_14553,N_13145,N_13812);
nor U14554 (N_14554,N_13909,N_13565);
xnor U14555 (N_14555,N_13960,N_13151);
and U14556 (N_14556,N_13794,N_13006);
xnor U14557 (N_14557,N_13875,N_13063);
and U14558 (N_14558,N_13020,N_13090);
and U14559 (N_14559,N_13543,N_13078);
and U14560 (N_14560,N_13969,N_13352);
nor U14561 (N_14561,N_13357,N_13902);
and U14562 (N_14562,N_13950,N_13019);
nand U14563 (N_14563,N_13648,N_13662);
or U14564 (N_14564,N_13498,N_13066);
nand U14565 (N_14565,N_13360,N_13427);
or U14566 (N_14566,N_13534,N_13807);
xor U14567 (N_14567,N_13433,N_13943);
xor U14568 (N_14568,N_13152,N_13334);
or U14569 (N_14569,N_13728,N_13204);
xor U14570 (N_14570,N_13586,N_13519);
nand U14571 (N_14571,N_13543,N_13846);
xor U14572 (N_14572,N_13853,N_13780);
or U14573 (N_14573,N_13427,N_13011);
nand U14574 (N_14574,N_13366,N_13690);
nor U14575 (N_14575,N_13136,N_13993);
or U14576 (N_14576,N_13191,N_13887);
and U14577 (N_14577,N_13828,N_13330);
xnor U14578 (N_14578,N_13283,N_13375);
and U14579 (N_14579,N_13637,N_13783);
nor U14580 (N_14580,N_13941,N_13643);
and U14581 (N_14581,N_13374,N_13740);
and U14582 (N_14582,N_13931,N_13327);
or U14583 (N_14583,N_13457,N_13945);
nor U14584 (N_14584,N_13420,N_13444);
xnor U14585 (N_14585,N_13406,N_13659);
nor U14586 (N_14586,N_13690,N_13054);
or U14587 (N_14587,N_13204,N_13374);
and U14588 (N_14588,N_13029,N_13550);
xnor U14589 (N_14589,N_13036,N_13586);
and U14590 (N_14590,N_13320,N_13015);
and U14591 (N_14591,N_13578,N_13071);
or U14592 (N_14592,N_13772,N_13418);
and U14593 (N_14593,N_13805,N_13961);
and U14594 (N_14594,N_13507,N_13714);
nand U14595 (N_14595,N_13963,N_13645);
and U14596 (N_14596,N_13910,N_13436);
nand U14597 (N_14597,N_13671,N_13346);
nor U14598 (N_14598,N_13506,N_13619);
nand U14599 (N_14599,N_13901,N_13645);
and U14600 (N_14600,N_13285,N_13981);
and U14601 (N_14601,N_13762,N_13739);
nand U14602 (N_14602,N_13591,N_13619);
or U14603 (N_14603,N_13671,N_13052);
or U14604 (N_14604,N_13979,N_13339);
or U14605 (N_14605,N_13884,N_13029);
and U14606 (N_14606,N_13910,N_13755);
and U14607 (N_14607,N_13226,N_13170);
and U14608 (N_14608,N_13082,N_13025);
nand U14609 (N_14609,N_13995,N_13737);
and U14610 (N_14610,N_13114,N_13530);
nand U14611 (N_14611,N_13728,N_13702);
nand U14612 (N_14612,N_13347,N_13970);
xnor U14613 (N_14613,N_13011,N_13435);
nor U14614 (N_14614,N_13733,N_13141);
xor U14615 (N_14615,N_13140,N_13611);
xor U14616 (N_14616,N_13439,N_13748);
nor U14617 (N_14617,N_13908,N_13820);
nor U14618 (N_14618,N_13028,N_13390);
xor U14619 (N_14619,N_13630,N_13606);
nand U14620 (N_14620,N_13956,N_13869);
xnor U14621 (N_14621,N_13067,N_13384);
xor U14622 (N_14622,N_13080,N_13896);
nor U14623 (N_14623,N_13330,N_13849);
and U14624 (N_14624,N_13198,N_13290);
or U14625 (N_14625,N_13453,N_13921);
and U14626 (N_14626,N_13603,N_13747);
or U14627 (N_14627,N_13459,N_13283);
nor U14628 (N_14628,N_13552,N_13184);
or U14629 (N_14629,N_13968,N_13317);
nand U14630 (N_14630,N_13419,N_13295);
nor U14631 (N_14631,N_13538,N_13276);
nor U14632 (N_14632,N_13686,N_13072);
nand U14633 (N_14633,N_13812,N_13778);
or U14634 (N_14634,N_13075,N_13600);
nand U14635 (N_14635,N_13561,N_13530);
nor U14636 (N_14636,N_13795,N_13707);
and U14637 (N_14637,N_13926,N_13136);
and U14638 (N_14638,N_13291,N_13817);
or U14639 (N_14639,N_13947,N_13474);
and U14640 (N_14640,N_13543,N_13643);
and U14641 (N_14641,N_13618,N_13307);
or U14642 (N_14642,N_13067,N_13534);
nand U14643 (N_14643,N_13111,N_13382);
nor U14644 (N_14644,N_13432,N_13104);
or U14645 (N_14645,N_13301,N_13353);
or U14646 (N_14646,N_13449,N_13986);
xnor U14647 (N_14647,N_13311,N_13905);
nor U14648 (N_14648,N_13492,N_13392);
nand U14649 (N_14649,N_13829,N_13859);
or U14650 (N_14650,N_13128,N_13228);
or U14651 (N_14651,N_13847,N_13439);
xor U14652 (N_14652,N_13930,N_13206);
nand U14653 (N_14653,N_13718,N_13335);
nand U14654 (N_14654,N_13868,N_13349);
or U14655 (N_14655,N_13938,N_13201);
nor U14656 (N_14656,N_13205,N_13742);
nor U14657 (N_14657,N_13982,N_13589);
nand U14658 (N_14658,N_13633,N_13927);
nor U14659 (N_14659,N_13691,N_13162);
and U14660 (N_14660,N_13990,N_13265);
xnor U14661 (N_14661,N_13247,N_13627);
nand U14662 (N_14662,N_13098,N_13722);
and U14663 (N_14663,N_13693,N_13241);
and U14664 (N_14664,N_13188,N_13189);
xnor U14665 (N_14665,N_13172,N_13443);
xor U14666 (N_14666,N_13110,N_13847);
or U14667 (N_14667,N_13288,N_13875);
xor U14668 (N_14668,N_13625,N_13892);
and U14669 (N_14669,N_13711,N_13686);
xnor U14670 (N_14670,N_13699,N_13072);
xor U14671 (N_14671,N_13899,N_13667);
nand U14672 (N_14672,N_13822,N_13178);
and U14673 (N_14673,N_13091,N_13798);
and U14674 (N_14674,N_13849,N_13844);
and U14675 (N_14675,N_13964,N_13682);
nand U14676 (N_14676,N_13828,N_13831);
nand U14677 (N_14677,N_13886,N_13931);
or U14678 (N_14678,N_13545,N_13272);
nand U14679 (N_14679,N_13111,N_13298);
or U14680 (N_14680,N_13181,N_13798);
xnor U14681 (N_14681,N_13803,N_13696);
nor U14682 (N_14682,N_13048,N_13917);
and U14683 (N_14683,N_13608,N_13357);
or U14684 (N_14684,N_13514,N_13316);
nor U14685 (N_14685,N_13411,N_13037);
or U14686 (N_14686,N_13760,N_13956);
nand U14687 (N_14687,N_13055,N_13186);
nand U14688 (N_14688,N_13846,N_13617);
nor U14689 (N_14689,N_13103,N_13093);
nor U14690 (N_14690,N_13584,N_13290);
xor U14691 (N_14691,N_13053,N_13085);
nand U14692 (N_14692,N_13755,N_13720);
and U14693 (N_14693,N_13598,N_13668);
xnor U14694 (N_14694,N_13735,N_13079);
or U14695 (N_14695,N_13901,N_13193);
or U14696 (N_14696,N_13621,N_13355);
nand U14697 (N_14697,N_13902,N_13367);
or U14698 (N_14698,N_13739,N_13422);
and U14699 (N_14699,N_13245,N_13207);
nor U14700 (N_14700,N_13943,N_13538);
xor U14701 (N_14701,N_13572,N_13377);
nor U14702 (N_14702,N_13210,N_13997);
nand U14703 (N_14703,N_13920,N_13200);
xnor U14704 (N_14704,N_13039,N_13854);
or U14705 (N_14705,N_13405,N_13300);
or U14706 (N_14706,N_13859,N_13927);
nand U14707 (N_14707,N_13012,N_13949);
nor U14708 (N_14708,N_13766,N_13034);
xnor U14709 (N_14709,N_13175,N_13749);
and U14710 (N_14710,N_13256,N_13485);
xnor U14711 (N_14711,N_13891,N_13297);
nand U14712 (N_14712,N_13135,N_13684);
xor U14713 (N_14713,N_13847,N_13589);
nor U14714 (N_14714,N_13601,N_13185);
nand U14715 (N_14715,N_13369,N_13159);
nand U14716 (N_14716,N_13011,N_13832);
and U14717 (N_14717,N_13283,N_13877);
nand U14718 (N_14718,N_13685,N_13582);
nor U14719 (N_14719,N_13312,N_13280);
and U14720 (N_14720,N_13487,N_13956);
nand U14721 (N_14721,N_13508,N_13595);
nand U14722 (N_14722,N_13091,N_13679);
nand U14723 (N_14723,N_13400,N_13066);
and U14724 (N_14724,N_13125,N_13276);
nor U14725 (N_14725,N_13157,N_13033);
and U14726 (N_14726,N_13507,N_13296);
or U14727 (N_14727,N_13785,N_13276);
nand U14728 (N_14728,N_13026,N_13934);
nor U14729 (N_14729,N_13854,N_13795);
nor U14730 (N_14730,N_13507,N_13263);
nand U14731 (N_14731,N_13090,N_13909);
or U14732 (N_14732,N_13413,N_13727);
nor U14733 (N_14733,N_13249,N_13016);
xor U14734 (N_14734,N_13572,N_13347);
xor U14735 (N_14735,N_13144,N_13285);
xor U14736 (N_14736,N_13012,N_13571);
xor U14737 (N_14737,N_13327,N_13520);
nor U14738 (N_14738,N_13307,N_13053);
nand U14739 (N_14739,N_13799,N_13242);
xnor U14740 (N_14740,N_13794,N_13538);
nand U14741 (N_14741,N_13701,N_13499);
nor U14742 (N_14742,N_13287,N_13170);
nor U14743 (N_14743,N_13799,N_13648);
xnor U14744 (N_14744,N_13795,N_13993);
nor U14745 (N_14745,N_13805,N_13281);
nor U14746 (N_14746,N_13553,N_13543);
xnor U14747 (N_14747,N_13873,N_13030);
and U14748 (N_14748,N_13939,N_13648);
and U14749 (N_14749,N_13827,N_13170);
nand U14750 (N_14750,N_13841,N_13410);
and U14751 (N_14751,N_13793,N_13538);
nor U14752 (N_14752,N_13077,N_13949);
and U14753 (N_14753,N_13291,N_13851);
or U14754 (N_14754,N_13176,N_13947);
nand U14755 (N_14755,N_13334,N_13424);
or U14756 (N_14756,N_13545,N_13127);
nand U14757 (N_14757,N_13833,N_13272);
or U14758 (N_14758,N_13907,N_13631);
or U14759 (N_14759,N_13726,N_13855);
nand U14760 (N_14760,N_13278,N_13457);
nor U14761 (N_14761,N_13291,N_13871);
nor U14762 (N_14762,N_13688,N_13366);
xor U14763 (N_14763,N_13818,N_13351);
or U14764 (N_14764,N_13032,N_13741);
and U14765 (N_14765,N_13964,N_13646);
and U14766 (N_14766,N_13952,N_13045);
and U14767 (N_14767,N_13032,N_13506);
nand U14768 (N_14768,N_13681,N_13800);
nor U14769 (N_14769,N_13154,N_13127);
xnor U14770 (N_14770,N_13708,N_13105);
nor U14771 (N_14771,N_13983,N_13928);
or U14772 (N_14772,N_13079,N_13564);
or U14773 (N_14773,N_13721,N_13584);
nor U14774 (N_14774,N_13254,N_13496);
nor U14775 (N_14775,N_13213,N_13881);
nand U14776 (N_14776,N_13678,N_13358);
nor U14777 (N_14777,N_13545,N_13807);
nor U14778 (N_14778,N_13599,N_13800);
xnor U14779 (N_14779,N_13696,N_13542);
xor U14780 (N_14780,N_13433,N_13904);
or U14781 (N_14781,N_13260,N_13845);
or U14782 (N_14782,N_13567,N_13847);
xor U14783 (N_14783,N_13900,N_13771);
nor U14784 (N_14784,N_13625,N_13627);
nand U14785 (N_14785,N_13333,N_13056);
and U14786 (N_14786,N_13560,N_13150);
xor U14787 (N_14787,N_13946,N_13821);
nand U14788 (N_14788,N_13833,N_13666);
nor U14789 (N_14789,N_13082,N_13184);
and U14790 (N_14790,N_13271,N_13041);
and U14791 (N_14791,N_13614,N_13985);
nand U14792 (N_14792,N_13270,N_13839);
or U14793 (N_14793,N_13353,N_13150);
nor U14794 (N_14794,N_13272,N_13222);
and U14795 (N_14795,N_13134,N_13627);
and U14796 (N_14796,N_13635,N_13347);
and U14797 (N_14797,N_13102,N_13013);
xnor U14798 (N_14798,N_13216,N_13833);
xnor U14799 (N_14799,N_13747,N_13244);
xnor U14800 (N_14800,N_13579,N_13323);
or U14801 (N_14801,N_13065,N_13313);
or U14802 (N_14802,N_13802,N_13159);
nand U14803 (N_14803,N_13207,N_13582);
or U14804 (N_14804,N_13465,N_13623);
nand U14805 (N_14805,N_13815,N_13302);
or U14806 (N_14806,N_13281,N_13666);
and U14807 (N_14807,N_13871,N_13008);
nand U14808 (N_14808,N_13619,N_13693);
nand U14809 (N_14809,N_13014,N_13819);
nor U14810 (N_14810,N_13401,N_13746);
xor U14811 (N_14811,N_13295,N_13300);
nand U14812 (N_14812,N_13685,N_13152);
or U14813 (N_14813,N_13340,N_13176);
nand U14814 (N_14814,N_13891,N_13098);
and U14815 (N_14815,N_13708,N_13890);
or U14816 (N_14816,N_13336,N_13170);
nor U14817 (N_14817,N_13507,N_13993);
and U14818 (N_14818,N_13342,N_13667);
or U14819 (N_14819,N_13765,N_13144);
nor U14820 (N_14820,N_13195,N_13109);
nand U14821 (N_14821,N_13417,N_13762);
nand U14822 (N_14822,N_13976,N_13031);
nand U14823 (N_14823,N_13722,N_13415);
nand U14824 (N_14824,N_13748,N_13793);
or U14825 (N_14825,N_13087,N_13976);
nor U14826 (N_14826,N_13565,N_13699);
and U14827 (N_14827,N_13936,N_13718);
xor U14828 (N_14828,N_13606,N_13575);
nor U14829 (N_14829,N_13867,N_13200);
and U14830 (N_14830,N_13354,N_13080);
nand U14831 (N_14831,N_13952,N_13333);
or U14832 (N_14832,N_13014,N_13186);
or U14833 (N_14833,N_13369,N_13975);
nor U14834 (N_14834,N_13796,N_13315);
nand U14835 (N_14835,N_13712,N_13032);
and U14836 (N_14836,N_13928,N_13132);
nand U14837 (N_14837,N_13852,N_13708);
nand U14838 (N_14838,N_13267,N_13368);
or U14839 (N_14839,N_13280,N_13544);
or U14840 (N_14840,N_13497,N_13223);
or U14841 (N_14841,N_13331,N_13686);
xnor U14842 (N_14842,N_13348,N_13925);
and U14843 (N_14843,N_13087,N_13034);
and U14844 (N_14844,N_13415,N_13135);
nand U14845 (N_14845,N_13845,N_13902);
xnor U14846 (N_14846,N_13390,N_13347);
nor U14847 (N_14847,N_13877,N_13083);
or U14848 (N_14848,N_13412,N_13858);
and U14849 (N_14849,N_13435,N_13429);
nand U14850 (N_14850,N_13989,N_13179);
and U14851 (N_14851,N_13897,N_13433);
nand U14852 (N_14852,N_13025,N_13516);
xor U14853 (N_14853,N_13640,N_13203);
xnor U14854 (N_14854,N_13621,N_13634);
nand U14855 (N_14855,N_13876,N_13276);
or U14856 (N_14856,N_13878,N_13744);
or U14857 (N_14857,N_13600,N_13500);
and U14858 (N_14858,N_13012,N_13841);
and U14859 (N_14859,N_13576,N_13129);
and U14860 (N_14860,N_13744,N_13918);
nand U14861 (N_14861,N_13901,N_13997);
xor U14862 (N_14862,N_13867,N_13163);
or U14863 (N_14863,N_13330,N_13300);
nor U14864 (N_14864,N_13889,N_13403);
nor U14865 (N_14865,N_13299,N_13596);
and U14866 (N_14866,N_13229,N_13189);
xnor U14867 (N_14867,N_13925,N_13163);
xor U14868 (N_14868,N_13923,N_13661);
and U14869 (N_14869,N_13551,N_13471);
nor U14870 (N_14870,N_13430,N_13054);
or U14871 (N_14871,N_13104,N_13989);
and U14872 (N_14872,N_13097,N_13004);
nand U14873 (N_14873,N_13215,N_13984);
nor U14874 (N_14874,N_13531,N_13836);
and U14875 (N_14875,N_13303,N_13354);
nor U14876 (N_14876,N_13904,N_13715);
nand U14877 (N_14877,N_13620,N_13470);
and U14878 (N_14878,N_13478,N_13830);
and U14879 (N_14879,N_13325,N_13577);
xor U14880 (N_14880,N_13330,N_13100);
nand U14881 (N_14881,N_13793,N_13961);
nor U14882 (N_14882,N_13451,N_13343);
and U14883 (N_14883,N_13212,N_13457);
and U14884 (N_14884,N_13111,N_13757);
nor U14885 (N_14885,N_13600,N_13798);
xnor U14886 (N_14886,N_13886,N_13207);
xor U14887 (N_14887,N_13923,N_13782);
or U14888 (N_14888,N_13376,N_13098);
and U14889 (N_14889,N_13635,N_13026);
and U14890 (N_14890,N_13555,N_13511);
nand U14891 (N_14891,N_13516,N_13565);
nor U14892 (N_14892,N_13371,N_13848);
nor U14893 (N_14893,N_13446,N_13611);
nor U14894 (N_14894,N_13755,N_13487);
or U14895 (N_14895,N_13308,N_13063);
xnor U14896 (N_14896,N_13491,N_13479);
nor U14897 (N_14897,N_13619,N_13870);
and U14898 (N_14898,N_13180,N_13007);
nand U14899 (N_14899,N_13931,N_13114);
nand U14900 (N_14900,N_13026,N_13103);
and U14901 (N_14901,N_13759,N_13494);
nor U14902 (N_14902,N_13895,N_13502);
or U14903 (N_14903,N_13704,N_13905);
or U14904 (N_14904,N_13332,N_13501);
nor U14905 (N_14905,N_13309,N_13890);
nand U14906 (N_14906,N_13649,N_13082);
nor U14907 (N_14907,N_13426,N_13478);
or U14908 (N_14908,N_13888,N_13507);
and U14909 (N_14909,N_13245,N_13037);
nand U14910 (N_14910,N_13567,N_13944);
nor U14911 (N_14911,N_13342,N_13710);
or U14912 (N_14912,N_13622,N_13880);
nand U14913 (N_14913,N_13922,N_13398);
nor U14914 (N_14914,N_13316,N_13165);
and U14915 (N_14915,N_13905,N_13396);
xor U14916 (N_14916,N_13805,N_13608);
xnor U14917 (N_14917,N_13379,N_13669);
or U14918 (N_14918,N_13444,N_13974);
nor U14919 (N_14919,N_13998,N_13692);
xnor U14920 (N_14920,N_13092,N_13069);
and U14921 (N_14921,N_13290,N_13271);
or U14922 (N_14922,N_13007,N_13031);
nor U14923 (N_14923,N_13170,N_13461);
xnor U14924 (N_14924,N_13877,N_13646);
and U14925 (N_14925,N_13181,N_13573);
xor U14926 (N_14926,N_13444,N_13898);
nor U14927 (N_14927,N_13740,N_13813);
and U14928 (N_14928,N_13905,N_13605);
nand U14929 (N_14929,N_13624,N_13966);
or U14930 (N_14930,N_13918,N_13773);
and U14931 (N_14931,N_13846,N_13588);
or U14932 (N_14932,N_13088,N_13509);
nand U14933 (N_14933,N_13788,N_13268);
nor U14934 (N_14934,N_13546,N_13988);
and U14935 (N_14935,N_13838,N_13656);
nand U14936 (N_14936,N_13838,N_13432);
and U14937 (N_14937,N_13619,N_13509);
nor U14938 (N_14938,N_13736,N_13157);
or U14939 (N_14939,N_13667,N_13991);
nor U14940 (N_14940,N_13302,N_13946);
nor U14941 (N_14941,N_13817,N_13653);
or U14942 (N_14942,N_13195,N_13231);
nor U14943 (N_14943,N_13770,N_13522);
nor U14944 (N_14944,N_13732,N_13484);
nor U14945 (N_14945,N_13446,N_13043);
nor U14946 (N_14946,N_13412,N_13532);
nand U14947 (N_14947,N_13155,N_13924);
nand U14948 (N_14948,N_13061,N_13713);
and U14949 (N_14949,N_13582,N_13690);
xor U14950 (N_14950,N_13435,N_13151);
nand U14951 (N_14951,N_13559,N_13563);
xor U14952 (N_14952,N_13342,N_13848);
or U14953 (N_14953,N_13123,N_13395);
and U14954 (N_14954,N_13906,N_13892);
or U14955 (N_14955,N_13448,N_13883);
xnor U14956 (N_14956,N_13949,N_13444);
xor U14957 (N_14957,N_13463,N_13821);
nand U14958 (N_14958,N_13014,N_13323);
or U14959 (N_14959,N_13733,N_13301);
and U14960 (N_14960,N_13606,N_13881);
and U14961 (N_14961,N_13808,N_13076);
nand U14962 (N_14962,N_13627,N_13157);
and U14963 (N_14963,N_13557,N_13894);
nand U14964 (N_14964,N_13150,N_13088);
xnor U14965 (N_14965,N_13404,N_13541);
or U14966 (N_14966,N_13258,N_13578);
nand U14967 (N_14967,N_13750,N_13954);
and U14968 (N_14968,N_13462,N_13474);
nor U14969 (N_14969,N_13637,N_13214);
or U14970 (N_14970,N_13278,N_13154);
nand U14971 (N_14971,N_13765,N_13977);
or U14972 (N_14972,N_13160,N_13826);
xnor U14973 (N_14973,N_13789,N_13631);
xnor U14974 (N_14974,N_13652,N_13583);
nor U14975 (N_14975,N_13827,N_13629);
or U14976 (N_14976,N_13619,N_13646);
nor U14977 (N_14977,N_13790,N_13295);
or U14978 (N_14978,N_13477,N_13959);
nor U14979 (N_14979,N_13182,N_13308);
and U14980 (N_14980,N_13008,N_13466);
and U14981 (N_14981,N_13749,N_13341);
xor U14982 (N_14982,N_13403,N_13061);
nand U14983 (N_14983,N_13368,N_13856);
nor U14984 (N_14984,N_13588,N_13570);
and U14985 (N_14985,N_13432,N_13718);
xor U14986 (N_14986,N_13710,N_13260);
and U14987 (N_14987,N_13218,N_13557);
nor U14988 (N_14988,N_13718,N_13918);
xor U14989 (N_14989,N_13389,N_13171);
xor U14990 (N_14990,N_13203,N_13780);
nand U14991 (N_14991,N_13769,N_13188);
nand U14992 (N_14992,N_13679,N_13992);
and U14993 (N_14993,N_13094,N_13988);
and U14994 (N_14994,N_13883,N_13740);
or U14995 (N_14995,N_13521,N_13146);
and U14996 (N_14996,N_13369,N_13513);
nand U14997 (N_14997,N_13846,N_13867);
or U14998 (N_14998,N_13694,N_13935);
xnor U14999 (N_14999,N_13979,N_13072);
xnor U15000 (N_15000,N_14140,N_14469);
nor U15001 (N_15001,N_14124,N_14129);
nor U15002 (N_15002,N_14725,N_14437);
or U15003 (N_15003,N_14379,N_14371);
and U15004 (N_15004,N_14528,N_14350);
and U15005 (N_15005,N_14650,N_14018);
nor U15006 (N_15006,N_14951,N_14246);
and U15007 (N_15007,N_14507,N_14585);
nor U15008 (N_15008,N_14274,N_14992);
nor U15009 (N_15009,N_14867,N_14556);
or U15010 (N_15010,N_14806,N_14257);
nor U15011 (N_15011,N_14891,N_14519);
nor U15012 (N_15012,N_14597,N_14742);
nor U15013 (N_15013,N_14813,N_14988);
or U15014 (N_15014,N_14835,N_14551);
and U15015 (N_15015,N_14938,N_14561);
xnor U15016 (N_15016,N_14984,N_14253);
nor U15017 (N_15017,N_14588,N_14238);
and U15018 (N_15018,N_14334,N_14996);
nor U15019 (N_15019,N_14213,N_14714);
or U15020 (N_15020,N_14541,N_14694);
nor U15021 (N_15021,N_14903,N_14506);
nor U15022 (N_15022,N_14981,N_14664);
or U15023 (N_15023,N_14530,N_14741);
xor U15024 (N_15024,N_14232,N_14663);
or U15025 (N_15025,N_14757,N_14728);
or U15026 (N_15026,N_14401,N_14746);
or U15027 (N_15027,N_14654,N_14491);
and U15028 (N_15028,N_14440,N_14115);
nand U15029 (N_15029,N_14252,N_14017);
xnor U15030 (N_15030,N_14021,N_14985);
and U15031 (N_15031,N_14127,N_14858);
nand U15032 (N_15032,N_14609,N_14831);
or U15033 (N_15033,N_14766,N_14305);
nor U15034 (N_15034,N_14472,N_14882);
nand U15035 (N_15035,N_14422,N_14655);
and U15036 (N_15036,N_14245,N_14973);
nor U15037 (N_15037,N_14627,N_14415);
or U15038 (N_15038,N_14414,N_14436);
and U15039 (N_15039,N_14780,N_14701);
and U15040 (N_15040,N_14689,N_14263);
and U15041 (N_15041,N_14003,N_14074);
or U15042 (N_15042,N_14395,N_14773);
or U15043 (N_15043,N_14665,N_14764);
xnor U15044 (N_15044,N_14693,N_14898);
and U15045 (N_15045,N_14308,N_14612);
xnor U15046 (N_15046,N_14760,N_14248);
and U15047 (N_15047,N_14575,N_14557);
and U15048 (N_15048,N_14630,N_14347);
nor U15049 (N_15049,N_14893,N_14738);
and U15050 (N_15050,N_14717,N_14463);
nor U15051 (N_15051,N_14567,N_14100);
nor U15052 (N_15052,N_14936,N_14614);
nor U15053 (N_15053,N_14505,N_14119);
or U15054 (N_15054,N_14862,N_14301);
or U15055 (N_15055,N_14323,N_14362);
or U15056 (N_15056,N_14976,N_14811);
xnor U15057 (N_15057,N_14958,N_14964);
and U15058 (N_15058,N_14777,N_14916);
and U15059 (N_15059,N_14358,N_14692);
and U15060 (N_15060,N_14251,N_14816);
or U15061 (N_15061,N_14917,N_14320);
and U15062 (N_15062,N_14312,N_14536);
nor U15063 (N_15063,N_14593,N_14427);
xor U15064 (N_15064,N_14241,N_14433);
and U15065 (N_15065,N_14836,N_14720);
nor U15066 (N_15066,N_14172,N_14486);
nor U15067 (N_15067,N_14118,N_14102);
xnor U15068 (N_15068,N_14933,N_14092);
or U15069 (N_15069,N_14259,N_14311);
and U15070 (N_15070,N_14107,N_14446);
nor U15071 (N_15071,N_14679,N_14577);
xnor U15072 (N_15072,N_14888,N_14887);
nand U15073 (N_15073,N_14032,N_14599);
nand U15074 (N_15074,N_14739,N_14752);
nand U15075 (N_15075,N_14355,N_14041);
nand U15076 (N_15076,N_14829,N_14188);
and U15077 (N_15077,N_14011,N_14130);
nand U15078 (N_15078,N_14591,N_14163);
and U15079 (N_15079,N_14131,N_14518);
nor U15080 (N_15080,N_14133,N_14687);
nor U15081 (N_15081,N_14025,N_14768);
xnor U15082 (N_15082,N_14429,N_14636);
xnor U15083 (N_15083,N_14517,N_14007);
nor U15084 (N_15084,N_14210,N_14456);
nand U15085 (N_15085,N_14834,N_14700);
nand U15086 (N_15086,N_14608,N_14269);
nand U15087 (N_15087,N_14151,N_14135);
or U15088 (N_15088,N_14563,N_14709);
xor U15089 (N_15089,N_14562,N_14897);
xnor U15090 (N_15090,N_14480,N_14657);
nand U15091 (N_15091,N_14382,N_14779);
nor U15092 (N_15092,N_14801,N_14980);
and U15093 (N_15093,N_14559,N_14162);
nand U15094 (N_15094,N_14112,N_14945);
nor U15095 (N_15095,N_14846,N_14059);
nor U15096 (N_15096,N_14703,N_14006);
xnor U15097 (N_15097,N_14158,N_14035);
and U15098 (N_15098,N_14089,N_14105);
nand U15099 (N_15099,N_14617,N_14106);
and U15100 (N_15100,N_14778,N_14474);
xnor U15101 (N_15101,N_14196,N_14789);
or U15102 (N_15102,N_14299,N_14885);
nor U15103 (N_15103,N_14444,N_14082);
or U15104 (N_15104,N_14084,N_14280);
nor U15105 (N_15105,N_14099,N_14791);
nand U15106 (N_15106,N_14616,N_14324);
or U15107 (N_15107,N_14468,N_14619);
nor U15108 (N_15108,N_14868,N_14497);
and U15109 (N_15109,N_14216,N_14383);
and U15110 (N_15110,N_14335,N_14328);
or U15111 (N_15111,N_14549,N_14645);
nand U15112 (N_15112,N_14043,N_14184);
nor U15113 (N_15113,N_14504,N_14808);
xor U15114 (N_15114,N_14351,N_14046);
xor U15115 (N_15115,N_14670,N_14109);
and U15116 (N_15116,N_14596,N_14143);
nor U15117 (N_15117,N_14134,N_14377);
nor U15118 (N_15118,N_14761,N_14496);
xnor U15119 (N_15119,N_14874,N_14521);
or U15120 (N_15120,N_14432,N_14604);
or U15121 (N_15121,N_14870,N_14000);
and U15122 (N_15122,N_14072,N_14750);
or U15123 (N_15123,N_14749,N_14526);
nand U15124 (N_15124,N_14830,N_14843);
xor U15125 (N_15125,N_14175,N_14157);
xnor U15126 (N_15126,N_14721,N_14145);
nand U15127 (N_15127,N_14234,N_14510);
xor U15128 (N_15128,N_14947,N_14576);
nor U15129 (N_15129,N_14851,N_14342);
nand U15130 (N_15130,N_14906,N_14322);
and U15131 (N_15131,N_14008,N_14572);
or U15132 (N_15132,N_14478,N_14641);
xor U15133 (N_15133,N_14441,N_14228);
nand U15134 (N_15134,N_14430,N_14426);
nor U15135 (N_15135,N_14704,N_14990);
and U15136 (N_15136,N_14822,N_14431);
xor U15137 (N_15137,N_14566,N_14681);
or U15138 (N_15138,N_14680,N_14533);
xnor U15139 (N_15139,N_14171,N_14096);
nand U15140 (N_15140,N_14598,N_14971);
or U15141 (N_15141,N_14838,N_14866);
or U15142 (N_15142,N_14818,N_14462);
and U15143 (N_15143,N_14359,N_14333);
xor U15144 (N_15144,N_14573,N_14406);
nand U15145 (N_15145,N_14628,N_14751);
or U15146 (N_15146,N_14982,N_14195);
or U15147 (N_15147,N_14756,N_14989);
nor U15148 (N_15148,N_14178,N_14690);
or U15149 (N_15149,N_14389,N_14343);
nor U15150 (N_15150,N_14297,N_14233);
nor U15151 (N_15151,N_14498,N_14722);
or U15152 (N_15152,N_14209,N_14673);
or U15153 (N_15153,N_14516,N_14772);
nand U15154 (N_15154,N_14423,N_14285);
nor U15155 (N_15155,N_14004,N_14164);
or U15156 (N_15156,N_14602,N_14114);
nor U15157 (N_15157,N_14959,N_14543);
nand U15158 (N_15158,N_14349,N_14144);
nor U15159 (N_15159,N_14592,N_14097);
and U15160 (N_15160,N_14384,N_14070);
nor U15161 (N_15161,N_14261,N_14036);
or U15162 (N_15162,N_14622,N_14674);
nand U15163 (N_15163,N_14219,N_14237);
or U15164 (N_15164,N_14101,N_14428);
and U15165 (N_15165,N_14847,N_14820);
nand U15166 (N_15166,N_14381,N_14170);
and U15167 (N_15167,N_14113,N_14073);
xor U15168 (N_15168,N_14476,N_14108);
and U15169 (N_15169,N_14056,N_14194);
and U15170 (N_15170,N_14077,N_14869);
xor U15171 (N_15171,N_14539,N_14487);
nand U15172 (N_15172,N_14016,N_14790);
nand U15173 (N_15173,N_14523,N_14889);
and U15174 (N_15174,N_14180,N_14946);
nor U15175 (N_15175,N_14057,N_14865);
and U15176 (N_15176,N_14775,N_14805);
nand U15177 (N_15177,N_14361,N_14452);
nand U15178 (N_15178,N_14797,N_14515);
or U15179 (N_15179,N_14438,N_14564);
and U15180 (N_15180,N_14513,N_14277);
nor U15181 (N_15181,N_14028,N_14247);
and U15182 (N_15182,N_14740,N_14642);
or U15183 (N_15183,N_14658,N_14048);
nor U15184 (N_15184,N_14998,N_14719);
or U15185 (N_15185,N_14715,N_14250);
and U15186 (N_15186,N_14753,N_14166);
xnor U15187 (N_15187,N_14705,N_14527);
nand U15188 (N_15188,N_14296,N_14769);
or U15189 (N_15189,N_14921,N_14877);
xor U15190 (N_15190,N_14110,N_14744);
and U15191 (N_15191,N_14603,N_14635);
nor U15192 (N_15192,N_14047,N_14442);
or U15193 (N_15193,N_14337,N_14950);
nand U15194 (N_15194,N_14207,N_14094);
or U15195 (N_15195,N_14221,N_14394);
nor U15196 (N_15196,N_14765,N_14640);
or U15197 (N_15197,N_14123,N_14827);
and U15198 (N_15198,N_14967,N_14483);
and U15199 (N_15199,N_14649,N_14987);
and U15200 (N_15200,N_14373,N_14782);
and U15201 (N_15201,N_14860,N_14538);
nand U15202 (N_15202,N_14999,N_14309);
and U15203 (N_15203,N_14995,N_14883);
nor U15204 (N_15204,N_14416,N_14267);
nand U15205 (N_15205,N_14465,N_14470);
or U15206 (N_15206,N_14339,N_14595);
nor U15207 (N_15207,N_14913,N_14126);
and U15208 (N_15208,N_14182,N_14009);
nand U15209 (N_15209,N_14812,N_14659);
or U15210 (N_15210,N_14369,N_14796);
and U15211 (N_15211,N_14318,N_14065);
xor U15212 (N_15212,N_14661,N_14230);
and U15213 (N_15213,N_14490,N_14409);
nand U15214 (N_15214,N_14859,N_14774);
xnor U15215 (N_15215,N_14249,N_14366);
and U15216 (N_15216,N_14439,N_14391);
nand U15217 (N_15217,N_14810,N_14300);
nor U15218 (N_15218,N_14288,N_14387);
nand U15219 (N_15219,N_14522,N_14943);
and U15220 (N_15220,N_14273,N_14052);
nor U15221 (N_15221,N_14520,N_14589);
and U15222 (N_15222,N_14892,N_14924);
nand U15223 (N_15223,N_14193,N_14168);
or U15224 (N_15224,N_14306,N_14884);
xnor U15225 (N_15225,N_14634,N_14286);
nand U15226 (N_15226,N_14434,N_14871);
nor U15227 (N_15227,N_14696,N_14647);
nand U15228 (N_15228,N_14532,N_14853);
nand U15229 (N_15229,N_14969,N_14907);
or U15230 (N_15230,N_14582,N_14302);
xor U15231 (N_15231,N_14968,N_14159);
nand U15232 (N_15232,N_14198,N_14378);
nand U15233 (N_15233,N_14901,N_14894);
nand U15234 (N_15234,N_14503,N_14828);
or U15235 (N_15235,N_14208,N_14223);
nor U15236 (N_15236,N_14500,N_14881);
nor U15237 (N_15237,N_14067,N_14142);
or U15238 (N_15238,N_14637,N_14511);
and U15239 (N_15239,N_14218,N_14653);
and U15240 (N_15240,N_14909,N_14012);
and U15241 (N_15241,N_14116,N_14844);
and U15242 (N_15242,N_14197,N_14098);
or U15243 (N_15243,N_14393,N_14804);
and U15244 (N_15244,N_14508,N_14443);
and U15245 (N_15245,N_14727,N_14402);
and U15246 (N_15246,N_14632,N_14733);
or U15247 (N_15247,N_14611,N_14939);
nor U15248 (N_15248,N_14878,N_14191);
nor U15249 (N_15249,N_14360,N_14356);
or U15250 (N_15250,N_14179,N_14346);
nor U15251 (N_15251,N_14024,N_14485);
or U15252 (N_15252,N_14660,N_14068);
and U15253 (N_15253,N_14137,N_14857);
and U15254 (N_15254,N_14514,N_14863);
and U15255 (N_15255,N_14716,N_14856);
and U15256 (N_15256,N_14254,N_14590);
nor U15257 (N_15257,N_14282,N_14029);
nand U15258 (N_15258,N_14544,N_14966);
nand U15259 (N_15259,N_14952,N_14581);
xor U15260 (N_15260,N_14932,N_14699);
nand U15261 (N_15261,N_14639,N_14606);
or U15262 (N_15262,N_14149,N_14785);
xnor U15263 (N_15263,N_14671,N_14633);
nand U15264 (N_15264,N_14363,N_14686);
and U15265 (N_15265,N_14060,N_14044);
xnor U15266 (N_15266,N_14919,N_14265);
xor U15267 (N_15267,N_14915,N_14167);
and U15268 (N_15268,N_14150,N_14155);
nand U15269 (N_15269,N_14710,N_14876);
nor U15270 (N_15270,N_14148,N_14918);
nor U15271 (N_15271,N_14450,N_14014);
xor U15272 (N_15272,N_14214,N_14783);
nor U15273 (N_15273,N_14390,N_14819);
xnor U15274 (N_15274,N_14656,N_14737);
nor U15275 (N_15275,N_14392,N_14177);
nor U15276 (N_15276,N_14537,N_14886);
nand U15277 (N_15277,N_14473,N_14880);
and U15278 (N_15278,N_14908,N_14502);
xnor U15279 (N_15279,N_14165,N_14316);
and U15280 (N_15280,N_14186,N_14125);
or U15281 (N_15281,N_14262,N_14678);
xor U15282 (N_15282,N_14552,N_14754);
nor U15283 (N_15283,N_14615,N_14104);
or U15284 (N_15284,N_14090,N_14161);
nand U15285 (N_15285,N_14574,N_14071);
nand U15286 (N_15286,N_14290,N_14281);
or U15287 (N_15287,N_14220,N_14111);
nand U15288 (N_15288,N_14997,N_14956);
xor U15289 (N_15289,N_14902,N_14117);
and U15290 (N_15290,N_14855,N_14817);
nand U15291 (N_15291,N_14944,N_14852);
nand U15292 (N_15292,N_14010,N_14038);
xor U15293 (N_15293,N_14050,N_14403);
nand U15294 (N_15294,N_14509,N_14492);
nor U15295 (N_15295,N_14449,N_14937);
xor U15296 (N_15296,N_14823,N_14957);
or U15297 (N_15297,N_14033,N_14374);
xor U15298 (N_15298,N_14983,N_14138);
nor U15299 (N_15299,N_14467,N_14934);
xor U15300 (N_15300,N_14512,N_14607);
nor U15301 (N_15301,N_14015,N_14310);
xnor U15302 (N_15302,N_14202,N_14648);
nor U15303 (N_15303,N_14698,N_14211);
nor U15304 (N_15304,N_14287,N_14093);
nand U15305 (N_15305,N_14187,N_14529);
nor U15306 (N_15306,N_14240,N_14942);
and U15307 (N_15307,N_14691,N_14019);
nor U15308 (N_15308,N_14289,N_14121);
xor U15309 (N_15309,N_14425,N_14357);
xor U15310 (N_15310,N_14708,N_14571);
nand U15311 (N_15311,N_14466,N_14420);
nor U15312 (N_15312,N_14458,N_14313);
and U15313 (N_15313,N_14341,N_14058);
or U15314 (N_15314,N_14418,N_14183);
xor U15315 (N_15315,N_14156,N_14555);
nor U15316 (N_15316,N_14307,N_14755);
and U15317 (N_15317,N_14718,N_14948);
nor U15318 (N_15318,N_14421,N_14034);
or U15319 (N_15319,N_14873,N_14268);
xor U15320 (N_15320,N_14685,N_14677);
or U15321 (N_15321,N_14479,N_14896);
xor U15322 (N_15322,N_14030,N_14174);
xor U15323 (N_15323,N_14330,N_14875);
nor U15324 (N_15324,N_14136,N_14979);
and U15325 (N_15325,N_14695,N_14554);
xor U15326 (N_15326,N_14457,N_14045);
or U15327 (N_15327,N_14375,N_14325);
or U15328 (N_15328,N_14850,N_14327);
and U15329 (N_15329,N_14153,N_14781);
nor U15330 (N_15330,N_14239,N_14970);
and U15331 (N_15331,N_14455,N_14833);
nor U15332 (N_15332,N_14570,N_14732);
or U15333 (N_15333,N_14173,N_14713);
nor U15334 (N_15334,N_14861,N_14954);
xnor U15335 (N_15335,N_14651,N_14494);
nand U15336 (N_15336,N_14540,N_14329);
xnor U15337 (N_15337,N_14340,N_14410);
xor U15338 (N_15338,N_14922,N_14600);
nor U15339 (N_15339,N_14203,N_14085);
or U15340 (N_15340,N_14075,N_14707);
nand U15341 (N_15341,N_14128,N_14683);
nor U15342 (N_15342,N_14424,N_14352);
nand U15343 (N_15343,N_14548,N_14227);
or U15344 (N_15344,N_14788,N_14493);
nor U15345 (N_15345,N_14594,N_14020);
nand U15346 (N_15346,N_14489,N_14039);
nor U15347 (N_15347,N_14911,N_14925);
and U15348 (N_15348,N_14488,N_14905);
nor U15349 (N_15349,N_14736,N_14303);
nor U15350 (N_15350,N_14978,N_14365);
nor U15351 (N_15351,N_14154,N_14185);
xnor U15352 (N_15352,N_14841,N_14929);
or U15353 (N_15353,N_14293,N_14258);
nand U15354 (N_15354,N_14372,N_14304);
nor U15355 (N_15355,N_14122,N_14826);
and U15356 (N_15356,N_14631,N_14731);
and U15357 (N_15357,N_14613,N_14794);
xnor U15358 (N_15358,N_14798,N_14083);
nor U15359 (N_15359,N_14845,N_14315);
nor U15360 (N_15360,N_14800,N_14879);
nor U15361 (N_15361,N_14348,N_14081);
nor U15362 (N_15362,N_14802,N_14368);
and U15363 (N_15363,N_14338,N_14499);
xnor U15364 (N_15364,N_14026,N_14912);
and U15365 (N_15365,N_14080,N_14941);
nand U15366 (N_15366,N_14629,N_14078);
xor U15367 (N_15367,N_14495,N_14666);
or U15368 (N_15368,N_14965,N_14062);
xor U15369 (N_15369,N_14955,N_14786);
or U15370 (N_15370,N_14275,N_14005);
or U15371 (N_15371,N_14849,N_14336);
nor U15372 (N_15372,N_14795,N_14076);
and U15373 (N_15373,N_14926,N_14899);
nand U15374 (N_15374,N_14146,N_14176);
and U15375 (N_15375,N_14064,N_14579);
nor U15376 (N_15376,N_14200,N_14181);
and U15377 (N_15377,N_14321,N_14279);
and U15378 (N_15378,N_14935,N_14459);
nand U15379 (N_15379,N_14923,N_14266);
nor U15380 (N_15380,N_14260,N_14055);
xnor U15381 (N_15381,N_14224,N_14294);
nand U15382 (N_15382,N_14620,N_14482);
or U15383 (N_15383,N_14688,N_14501);
and U15384 (N_15384,N_14061,N_14484);
or U15385 (N_15385,N_14412,N_14940);
and U15386 (N_15386,N_14991,N_14646);
xor U15387 (N_15387,N_14625,N_14669);
nor U15388 (N_15388,N_14408,N_14762);
and U15389 (N_15389,N_14626,N_14397);
and U15390 (N_15390,N_14475,N_14550);
and U15391 (N_15391,N_14087,N_14994);
nand U15392 (N_15392,N_14023,N_14624);
nand U15393 (N_15393,N_14461,N_14001);
and U15394 (N_15394,N_14792,N_14027);
and U15395 (N_15395,N_14095,N_14832);
nand U15396 (N_15396,N_14776,N_14724);
nand U15397 (N_15397,N_14711,N_14419);
nor U15398 (N_15398,N_14747,N_14037);
xnor U15399 (N_15399,N_14002,N_14545);
nand U15400 (N_15400,N_14726,N_14031);
or U15401 (N_15401,N_14413,N_14837);
and U15402 (N_15402,N_14454,N_14231);
nand U15403 (N_15403,N_14962,N_14895);
nand U15404 (N_15404,N_14580,N_14445);
or U15405 (N_15405,N_14206,N_14364);
and U15406 (N_15406,N_14730,N_14464);
or U15407 (N_15407,N_14236,N_14960);
nand U15408 (N_15408,N_14824,N_14217);
or U15409 (N_15409,N_14793,N_14993);
nand U15410 (N_15410,N_14255,N_14477);
nand U15411 (N_15411,N_14407,N_14481);
or U15412 (N_15412,N_14920,N_14212);
and U15413 (N_15413,N_14767,N_14949);
xor U15414 (N_15414,N_14398,N_14809);
nor U15415 (N_15415,N_14748,N_14723);
xnor U15416 (N_15416,N_14974,N_14558);
or U15417 (N_15417,N_14553,N_14667);
xor U15418 (N_15418,N_14448,N_14388);
nor U15419 (N_15419,N_14049,N_14222);
nor U15420 (N_15420,N_14256,N_14354);
xnor U15421 (N_15421,N_14367,N_14292);
nor U15422 (N_15422,N_14584,N_14215);
and U15423 (N_15423,N_14396,N_14244);
or U15424 (N_15424,N_14525,N_14091);
nand U15425 (N_15425,N_14332,N_14291);
nor U15426 (N_15426,N_14702,N_14063);
xor U15427 (N_15427,N_14840,N_14271);
and U15428 (N_15428,N_14904,N_14839);
or U15429 (N_15429,N_14385,N_14298);
xor U15430 (N_15430,N_14743,N_14623);
and U15431 (N_15431,N_14758,N_14684);
and U15432 (N_15432,N_14417,N_14662);
nor U15433 (N_15433,N_14447,N_14264);
nor U15434 (N_15434,N_14344,N_14225);
nand U15435 (N_15435,N_14147,N_14900);
xnor U15436 (N_15436,N_14242,N_14471);
nor U15437 (N_15437,N_14283,N_14644);
and U15438 (N_15438,N_14546,N_14638);
and U15439 (N_15439,N_14931,N_14815);
nor U15440 (N_15440,N_14201,N_14054);
xor U15441 (N_15441,N_14668,N_14542);
xor U15442 (N_15442,N_14930,N_14069);
or U15443 (N_15443,N_14565,N_14331);
nor U15444 (N_15444,N_14910,N_14120);
nand U15445 (N_15445,N_14848,N_14160);
or U15446 (N_15446,N_14961,N_14854);
or U15447 (N_15447,N_14270,N_14152);
nor U15448 (N_15448,N_14205,N_14411);
and U15449 (N_15449,N_14088,N_14460);
nor U15450 (N_15450,N_14405,N_14547);
nand U15451 (N_15451,N_14814,N_14643);
and U15452 (N_15452,N_14278,N_14169);
or U15453 (N_15453,N_14803,N_14825);
nor U15454 (N_15454,N_14229,N_14928);
and U15455 (N_15455,N_14534,N_14022);
and U15456 (N_15456,N_14053,N_14784);
xnor U15457 (N_15457,N_14086,N_14672);
nor U15458 (N_15458,N_14927,N_14051);
xor U15459 (N_15459,N_14975,N_14353);
nand U15460 (N_15460,N_14986,N_14042);
and U15461 (N_15461,N_14914,N_14189);
nand U15462 (N_15462,N_14963,N_14586);
nand U15463 (N_15463,N_14569,N_14326);
nand U15464 (N_15464,N_14953,N_14807);
nor U15465 (N_15465,N_14842,N_14319);
xnor U15466 (N_15466,N_14745,N_14380);
nor U15467 (N_15467,N_14272,N_14404);
nor U15468 (N_15468,N_14652,N_14226);
or U15469 (N_15469,N_14621,N_14771);
nor U15470 (N_15470,N_14040,N_14370);
and U15471 (N_15471,N_14192,N_14560);
xnor U15472 (N_15472,N_14400,N_14314);
or U15473 (N_15473,N_14729,N_14013);
or U15474 (N_15474,N_14583,N_14735);
and U15475 (N_15475,N_14235,N_14531);
nand U15476 (N_15476,N_14284,N_14103);
nor U15477 (N_15477,N_14799,N_14682);
nor U15478 (N_15478,N_14770,N_14276);
nor U15479 (N_15479,N_14787,N_14190);
or U15480 (N_15480,N_14066,N_14453);
nor U15481 (N_15481,N_14243,N_14675);
xor U15482 (N_15482,N_14141,N_14199);
nand U15483 (N_15483,N_14435,N_14295);
xnor U15484 (N_15484,N_14578,N_14601);
nand U15485 (N_15485,N_14568,N_14864);
nand U15486 (N_15486,N_14697,N_14399);
nor U15487 (N_15487,N_14587,N_14079);
nand U15488 (N_15488,N_14139,N_14345);
or U15489 (N_15489,N_14376,N_14734);
or U15490 (N_15490,N_14386,N_14972);
nand U15491 (N_15491,N_14451,N_14821);
nand U15492 (N_15492,N_14132,N_14872);
and U15493 (N_15493,N_14317,N_14676);
nand U15494 (N_15494,N_14524,N_14618);
or U15495 (N_15495,N_14890,N_14977);
or U15496 (N_15496,N_14605,N_14759);
nand U15497 (N_15497,N_14706,N_14535);
nand U15498 (N_15498,N_14610,N_14763);
or U15499 (N_15499,N_14712,N_14204);
or U15500 (N_15500,N_14824,N_14619);
nand U15501 (N_15501,N_14679,N_14965);
and U15502 (N_15502,N_14247,N_14506);
and U15503 (N_15503,N_14481,N_14343);
and U15504 (N_15504,N_14765,N_14089);
nand U15505 (N_15505,N_14144,N_14764);
nand U15506 (N_15506,N_14590,N_14564);
and U15507 (N_15507,N_14342,N_14574);
nor U15508 (N_15508,N_14141,N_14782);
or U15509 (N_15509,N_14349,N_14648);
xnor U15510 (N_15510,N_14003,N_14787);
xor U15511 (N_15511,N_14148,N_14068);
and U15512 (N_15512,N_14012,N_14168);
nand U15513 (N_15513,N_14363,N_14630);
nor U15514 (N_15514,N_14912,N_14721);
xor U15515 (N_15515,N_14478,N_14387);
nand U15516 (N_15516,N_14392,N_14931);
and U15517 (N_15517,N_14502,N_14651);
xor U15518 (N_15518,N_14669,N_14718);
nand U15519 (N_15519,N_14497,N_14851);
xnor U15520 (N_15520,N_14111,N_14906);
or U15521 (N_15521,N_14134,N_14856);
or U15522 (N_15522,N_14792,N_14041);
or U15523 (N_15523,N_14200,N_14561);
nand U15524 (N_15524,N_14308,N_14222);
or U15525 (N_15525,N_14234,N_14811);
or U15526 (N_15526,N_14771,N_14806);
xnor U15527 (N_15527,N_14472,N_14565);
or U15528 (N_15528,N_14177,N_14958);
nand U15529 (N_15529,N_14020,N_14236);
nand U15530 (N_15530,N_14664,N_14180);
nand U15531 (N_15531,N_14203,N_14171);
nand U15532 (N_15532,N_14486,N_14315);
xor U15533 (N_15533,N_14171,N_14104);
or U15534 (N_15534,N_14920,N_14262);
nor U15535 (N_15535,N_14367,N_14575);
and U15536 (N_15536,N_14839,N_14173);
nand U15537 (N_15537,N_14098,N_14745);
xnor U15538 (N_15538,N_14621,N_14415);
xor U15539 (N_15539,N_14904,N_14167);
or U15540 (N_15540,N_14081,N_14028);
and U15541 (N_15541,N_14156,N_14104);
nor U15542 (N_15542,N_14632,N_14030);
and U15543 (N_15543,N_14821,N_14464);
or U15544 (N_15544,N_14804,N_14378);
or U15545 (N_15545,N_14041,N_14861);
xor U15546 (N_15546,N_14181,N_14474);
or U15547 (N_15547,N_14388,N_14129);
nand U15548 (N_15548,N_14176,N_14029);
xor U15549 (N_15549,N_14228,N_14779);
and U15550 (N_15550,N_14278,N_14119);
and U15551 (N_15551,N_14008,N_14619);
nand U15552 (N_15552,N_14119,N_14522);
nand U15553 (N_15553,N_14287,N_14985);
or U15554 (N_15554,N_14429,N_14140);
xnor U15555 (N_15555,N_14765,N_14663);
nand U15556 (N_15556,N_14810,N_14241);
or U15557 (N_15557,N_14331,N_14454);
nor U15558 (N_15558,N_14681,N_14368);
and U15559 (N_15559,N_14421,N_14044);
nand U15560 (N_15560,N_14247,N_14245);
or U15561 (N_15561,N_14383,N_14351);
nor U15562 (N_15562,N_14245,N_14988);
nor U15563 (N_15563,N_14450,N_14139);
nand U15564 (N_15564,N_14412,N_14610);
nor U15565 (N_15565,N_14072,N_14008);
nand U15566 (N_15566,N_14356,N_14164);
nor U15567 (N_15567,N_14348,N_14543);
nor U15568 (N_15568,N_14556,N_14665);
or U15569 (N_15569,N_14017,N_14734);
nor U15570 (N_15570,N_14329,N_14482);
nand U15571 (N_15571,N_14246,N_14404);
xor U15572 (N_15572,N_14315,N_14225);
and U15573 (N_15573,N_14495,N_14883);
or U15574 (N_15574,N_14645,N_14538);
xor U15575 (N_15575,N_14738,N_14786);
or U15576 (N_15576,N_14390,N_14435);
nand U15577 (N_15577,N_14790,N_14088);
xor U15578 (N_15578,N_14569,N_14273);
or U15579 (N_15579,N_14205,N_14039);
or U15580 (N_15580,N_14059,N_14689);
nor U15581 (N_15581,N_14744,N_14447);
xor U15582 (N_15582,N_14283,N_14177);
nand U15583 (N_15583,N_14665,N_14159);
nand U15584 (N_15584,N_14698,N_14901);
nand U15585 (N_15585,N_14970,N_14276);
or U15586 (N_15586,N_14415,N_14013);
nor U15587 (N_15587,N_14608,N_14858);
nand U15588 (N_15588,N_14473,N_14764);
nand U15589 (N_15589,N_14468,N_14015);
xor U15590 (N_15590,N_14686,N_14464);
nor U15591 (N_15591,N_14776,N_14429);
xnor U15592 (N_15592,N_14495,N_14449);
and U15593 (N_15593,N_14310,N_14789);
and U15594 (N_15594,N_14916,N_14801);
xor U15595 (N_15595,N_14227,N_14391);
and U15596 (N_15596,N_14779,N_14624);
and U15597 (N_15597,N_14804,N_14707);
nand U15598 (N_15598,N_14230,N_14784);
or U15599 (N_15599,N_14212,N_14901);
or U15600 (N_15600,N_14665,N_14194);
and U15601 (N_15601,N_14299,N_14292);
nand U15602 (N_15602,N_14361,N_14994);
nor U15603 (N_15603,N_14910,N_14952);
nor U15604 (N_15604,N_14233,N_14619);
nand U15605 (N_15605,N_14921,N_14157);
nor U15606 (N_15606,N_14459,N_14672);
nand U15607 (N_15607,N_14413,N_14248);
and U15608 (N_15608,N_14349,N_14972);
nand U15609 (N_15609,N_14525,N_14987);
nand U15610 (N_15610,N_14893,N_14160);
nand U15611 (N_15611,N_14231,N_14850);
nand U15612 (N_15612,N_14024,N_14655);
nand U15613 (N_15613,N_14080,N_14587);
or U15614 (N_15614,N_14936,N_14505);
xnor U15615 (N_15615,N_14296,N_14519);
nor U15616 (N_15616,N_14414,N_14058);
or U15617 (N_15617,N_14709,N_14152);
xor U15618 (N_15618,N_14664,N_14918);
xor U15619 (N_15619,N_14849,N_14713);
nand U15620 (N_15620,N_14065,N_14676);
xor U15621 (N_15621,N_14117,N_14382);
nand U15622 (N_15622,N_14178,N_14925);
xnor U15623 (N_15623,N_14870,N_14792);
xor U15624 (N_15624,N_14627,N_14006);
nor U15625 (N_15625,N_14803,N_14284);
nand U15626 (N_15626,N_14956,N_14849);
xnor U15627 (N_15627,N_14404,N_14441);
nand U15628 (N_15628,N_14508,N_14736);
nor U15629 (N_15629,N_14066,N_14430);
or U15630 (N_15630,N_14722,N_14948);
nor U15631 (N_15631,N_14938,N_14653);
or U15632 (N_15632,N_14767,N_14280);
or U15633 (N_15633,N_14604,N_14921);
nand U15634 (N_15634,N_14657,N_14814);
or U15635 (N_15635,N_14203,N_14881);
or U15636 (N_15636,N_14692,N_14485);
or U15637 (N_15637,N_14666,N_14800);
nand U15638 (N_15638,N_14162,N_14881);
nor U15639 (N_15639,N_14555,N_14870);
nand U15640 (N_15640,N_14538,N_14361);
and U15641 (N_15641,N_14530,N_14230);
nand U15642 (N_15642,N_14251,N_14893);
xnor U15643 (N_15643,N_14767,N_14236);
nand U15644 (N_15644,N_14278,N_14214);
nand U15645 (N_15645,N_14658,N_14292);
nor U15646 (N_15646,N_14267,N_14960);
or U15647 (N_15647,N_14749,N_14547);
or U15648 (N_15648,N_14372,N_14048);
or U15649 (N_15649,N_14379,N_14196);
xor U15650 (N_15650,N_14992,N_14126);
or U15651 (N_15651,N_14591,N_14469);
nor U15652 (N_15652,N_14075,N_14650);
or U15653 (N_15653,N_14939,N_14252);
nor U15654 (N_15654,N_14127,N_14442);
or U15655 (N_15655,N_14815,N_14413);
nand U15656 (N_15656,N_14745,N_14698);
or U15657 (N_15657,N_14053,N_14867);
nor U15658 (N_15658,N_14853,N_14933);
and U15659 (N_15659,N_14713,N_14109);
nor U15660 (N_15660,N_14176,N_14793);
nand U15661 (N_15661,N_14984,N_14640);
nand U15662 (N_15662,N_14357,N_14614);
nand U15663 (N_15663,N_14396,N_14873);
xnor U15664 (N_15664,N_14831,N_14139);
nor U15665 (N_15665,N_14201,N_14723);
xnor U15666 (N_15666,N_14656,N_14173);
nor U15667 (N_15667,N_14416,N_14375);
nor U15668 (N_15668,N_14682,N_14164);
xnor U15669 (N_15669,N_14895,N_14847);
xnor U15670 (N_15670,N_14359,N_14278);
nor U15671 (N_15671,N_14606,N_14649);
nor U15672 (N_15672,N_14390,N_14633);
and U15673 (N_15673,N_14176,N_14787);
nand U15674 (N_15674,N_14661,N_14370);
or U15675 (N_15675,N_14279,N_14500);
and U15676 (N_15676,N_14016,N_14657);
and U15677 (N_15677,N_14430,N_14708);
nand U15678 (N_15678,N_14141,N_14965);
or U15679 (N_15679,N_14494,N_14272);
nor U15680 (N_15680,N_14587,N_14894);
xnor U15681 (N_15681,N_14672,N_14777);
nand U15682 (N_15682,N_14044,N_14882);
nand U15683 (N_15683,N_14377,N_14818);
nand U15684 (N_15684,N_14017,N_14031);
nor U15685 (N_15685,N_14978,N_14680);
nor U15686 (N_15686,N_14702,N_14443);
xnor U15687 (N_15687,N_14719,N_14222);
and U15688 (N_15688,N_14160,N_14804);
nor U15689 (N_15689,N_14623,N_14673);
or U15690 (N_15690,N_14090,N_14672);
and U15691 (N_15691,N_14662,N_14752);
nand U15692 (N_15692,N_14110,N_14258);
or U15693 (N_15693,N_14499,N_14062);
or U15694 (N_15694,N_14017,N_14235);
nand U15695 (N_15695,N_14689,N_14003);
or U15696 (N_15696,N_14524,N_14067);
xnor U15697 (N_15697,N_14673,N_14285);
and U15698 (N_15698,N_14288,N_14279);
nand U15699 (N_15699,N_14341,N_14218);
nand U15700 (N_15700,N_14975,N_14021);
or U15701 (N_15701,N_14179,N_14626);
xor U15702 (N_15702,N_14741,N_14966);
nor U15703 (N_15703,N_14218,N_14585);
or U15704 (N_15704,N_14122,N_14249);
nand U15705 (N_15705,N_14714,N_14184);
and U15706 (N_15706,N_14810,N_14945);
or U15707 (N_15707,N_14998,N_14279);
xor U15708 (N_15708,N_14233,N_14177);
xor U15709 (N_15709,N_14060,N_14572);
xnor U15710 (N_15710,N_14505,N_14599);
nor U15711 (N_15711,N_14775,N_14777);
or U15712 (N_15712,N_14584,N_14970);
nand U15713 (N_15713,N_14580,N_14011);
or U15714 (N_15714,N_14000,N_14188);
or U15715 (N_15715,N_14834,N_14001);
or U15716 (N_15716,N_14883,N_14170);
xor U15717 (N_15717,N_14076,N_14264);
or U15718 (N_15718,N_14865,N_14499);
nor U15719 (N_15719,N_14202,N_14942);
and U15720 (N_15720,N_14979,N_14510);
or U15721 (N_15721,N_14751,N_14400);
or U15722 (N_15722,N_14154,N_14076);
or U15723 (N_15723,N_14131,N_14264);
nor U15724 (N_15724,N_14034,N_14790);
nand U15725 (N_15725,N_14495,N_14141);
nor U15726 (N_15726,N_14080,N_14449);
and U15727 (N_15727,N_14109,N_14309);
xnor U15728 (N_15728,N_14081,N_14835);
and U15729 (N_15729,N_14276,N_14238);
xnor U15730 (N_15730,N_14302,N_14248);
or U15731 (N_15731,N_14556,N_14510);
and U15732 (N_15732,N_14985,N_14164);
xor U15733 (N_15733,N_14075,N_14058);
and U15734 (N_15734,N_14135,N_14541);
xor U15735 (N_15735,N_14304,N_14770);
or U15736 (N_15736,N_14101,N_14194);
or U15737 (N_15737,N_14797,N_14833);
xnor U15738 (N_15738,N_14770,N_14319);
xnor U15739 (N_15739,N_14423,N_14000);
xor U15740 (N_15740,N_14233,N_14070);
or U15741 (N_15741,N_14448,N_14624);
nor U15742 (N_15742,N_14512,N_14962);
nand U15743 (N_15743,N_14710,N_14028);
nand U15744 (N_15744,N_14250,N_14473);
xnor U15745 (N_15745,N_14768,N_14229);
nand U15746 (N_15746,N_14044,N_14896);
or U15747 (N_15747,N_14376,N_14485);
xnor U15748 (N_15748,N_14812,N_14212);
nand U15749 (N_15749,N_14023,N_14373);
nand U15750 (N_15750,N_14249,N_14559);
or U15751 (N_15751,N_14032,N_14822);
or U15752 (N_15752,N_14687,N_14891);
nand U15753 (N_15753,N_14727,N_14412);
nand U15754 (N_15754,N_14515,N_14416);
xnor U15755 (N_15755,N_14097,N_14828);
and U15756 (N_15756,N_14509,N_14284);
nor U15757 (N_15757,N_14556,N_14306);
nor U15758 (N_15758,N_14815,N_14990);
xnor U15759 (N_15759,N_14599,N_14481);
xnor U15760 (N_15760,N_14773,N_14414);
nand U15761 (N_15761,N_14304,N_14238);
or U15762 (N_15762,N_14978,N_14483);
nand U15763 (N_15763,N_14156,N_14579);
nand U15764 (N_15764,N_14502,N_14843);
xor U15765 (N_15765,N_14692,N_14228);
nor U15766 (N_15766,N_14439,N_14427);
nor U15767 (N_15767,N_14579,N_14870);
xor U15768 (N_15768,N_14829,N_14066);
and U15769 (N_15769,N_14124,N_14799);
and U15770 (N_15770,N_14976,N_14181);
xnor U15771 (N_15771,N_14349,N_14635);
or U15772 (N_15772,N_14449,N_14497);
nand U15773 (N_15773,N_14531,N_14814);
xnor U15774 (N_15774,N_14630,N_14742);
nor U15775 (N_15775,N_14613,N_14361);
nor U15776 (N_15776,N_14635,N_14213);
nor U15777 (N_15777,N_14678,N_14583);
and U15778 (N_15778,N_14830,N_14588);
or U15779 (N_15779,N_14914,N_14729);
and U15780 (N_15780,N_14390,N_14382);
nor U15781 (N_15781,N_14057,N_14740);
xnor U15782 (N_15782,N_14677,N_14124);
nor U15783 (N_15783,N_14104,N_14052);
nor U15784 (N_15784,N_14491,N_14305);
or U15785 (N_15785,N_14481,N_14255);
nand U15786 (N_15786,N_14936,N_14827);
and U15787 (N_15787,N_14158,N_14796);
xor U15788 (N_15788,N_14225,N_14787);
or U15789 (N_15789,N_14407,N_14581);
xnor U15790 (N_15790,N_14889,N_14133);
nor U15791 (N_15791,N_14629,N_14032);
and U15792 (N_15792,N_14493,N_14008);
nor U15793 (N_15793,N_14339,N_14905);
nor U15794 (N_15794,N_14380,N_14250);
and U15795 (N_15795,N_14098,N_14623);
nand U15796 (N_15796,N_14210,N_14180);
nor U15797 (N_15797,N_14219,N_14220);
and U15798 (N_15798,N_14748,N_14150);
nand U15799 (N_15799,N_14905,N_14456);
xnor U15800 (N_15800,N_14445,N_14769);
xor U15801 (N_15801,N_14783,N_14779);
and U15802 (N_15802,N_14142,N_14371);
nand U15803 (N_15803,N_14830,N_14191);
and U15804 (N_15804,N_14971,N_14533);
xor U15805 (N_15805,N_14840,N_14192);
nor U15806 (N_15806,N_14363,N_14866);
xnor U15807 (N_15807,N_14257,N_14082);
nand U15808 (N_15808,N_14797,N_14915);
xor U15809 (N_15809,N_14729,N_14114);
xor U15810 (N_15810,N_14507,N_14201);
nand U15811 (N_15811,N_14469,N_14218);
or U15812 (N_15812,N_14391,N_14568);
nor U15813 (N_15813,N_14615,N_14094);
or U15814 (N_15814,N_14437,N_14503);
and U15815 (N_15815,N_14114,N_14312);
and U15816 (N_15816,N_14424,N_14944);
xnor U15817 (N_15817,N_14143,N_14709);
xor U15818 (N_15818,N_14173,N_14159);
nand U15819 (N_15819,N_14164,N_14661);
and U15820 (N_15820,N_14321,N_14467);
or U15821 (N_15821,N_14710,N_14482);
xnor U15822 (N_15822,N_14586,N_14391);
and U15823 (N_15823,N_14260,N_14485);
and U15824 (N_15824,N_14256,N_14672);
or U15825 (N_15825,N_14007,N_14356);
xor U15826 (N_15826,N_14161,N_14383);
nand U15827 (N_15827,N_14260,N_14860);
and U15828 (N_15828,N_14663,N_14690);
and U15829 (N_15829,N_14219,N_14400);
and U15830 (N_15830,N_14369,N_14604);
and U15831 (N_15831,N_14827,N_14081);
nand U15832 (N_15832,N_14426,N_14880);
nand U15833 (N_15833,N_14176,N_14922);
nor U15834 (N_15834,N_14077,N_14911);
nand U15835 (N_15835,N_14690,N_14079);
or U15836 (N_15836,N_14541,N_14043);
nand U15837 (N_15837,N_14047,N_14758);
nand U15838 (N_15838,N_14501,N_14600);
xnor U15839 (N_15839,N_14875,N_14615);
nor U15840 (N_15840,N_14062,N_14292);
nand U15841 (N_15841,N_14789,N_14079);
xnor U15842 (N_15842,N_14752,N_14144);
nor U15843 (N_15843,N_14824,N_14785);
nand U15844 (N_15844,N_14317,N_14649);
xor U15845 (N_15845,N_14556,N_14897);
nand U15846 (N_15846,N_14155,N_14271);
xor U15847 (N_15847,N_14196,N_14677);
or U15848 (N_15848,N_14228,N_14545);
and U15849 (N_15849,N_14387,N_14853);
and U15850 (N_15850,N_14491,N_14249);
and U15851 (N_15851,N_14192,N_14356);
nand U15852 (N_15852,N_14179,N_14032);
nor U15853 (N_15853,N_14036,N_14926);
nand U15854 (N_15854,N_14844,N_14842);
and U15855 (N_15855,N_14176,N_14291);
and U15856 (N_15856,N_14541,N_14050);
nand U15857 (N_15857,N_14022,N_14754);
nor U15858 (N_15858,N_14162,N_14841);
nor U15859 (N_15859,N_14806,N_14701);
xor U15860 (N_15860,N_14825,N_14014);
nor U15861 (N_15861,N_14469,N_14456);
and U15862 (N_15862,N_14747,N_14384);
nor U15863 (N_15863,N_14142,N_14836);
nand U15864 (N_15864,N_14350,N_14605);
nand U15865 (N_15865,N_14092,N_14326);
or U15866 (N_15866,N_14460,N_14777);
nand U15867 (N_15867,N_14476,N_14813);
nor U15868 (N_15868,N_14343,N_14229);
xnor U15869 (N_15869,N_14320,N_14298);
and U15870 (N_15870,N_14166,N_14736);
nor U15871 (N_15871,N_14371,N_14261);
nor U15872 (N_15872,N_14109,N_14527);
or U15873 (N_15873,N_14305,N_14865);
or U15874 (N_15874,N_14766,N_14839);
and U15875 (N_15875,N_14836,N_14278);
nand U15876 (N_15876,N_14832,N_14305);
or U15877 (N_15877,N_14817,N_14041);
nand U15878 (N_15878,N_14512,N_14016);
and U15879 (N_15879,N_14243,N_14872);
nand U15880 (N_15880,N_14650,N_14530);
nor U15881 (N_15881,N_14425,N_14358);
nand U15882 (N_15882,N_14188,N_14002);
nand U15883 (N_15883,N_14874,N_14156);
nand U15884 (N_15884,N_14328,N_14128);
xnor U15885 (N_15885,N_14711,N_14792);
nor U15886 (N_15886,N_14067,N_14885);
nor U15887 (N_15887,N_14411,N_14075);
nor U15888 (N_15888,N_14807,N_14144);
nand U15889 (N_15889,N_14870,N_14754);
xor U15890 (N_15890,N_14305,N_14572);
nand U15891 (N_15891,N_14242,N_14481);
and U15892 (N_15892,N_14984,N_14296);
nand U15893 (N_15893,N_14475,N_14243);
or U15894 (N_15894,N_14957,N_14237);
or U15895 (N_15895,N_14130,N_14431);
and U15896 (N_15896,N_14006,N_14784);
or U15897 (N_15897,N_14122,N_14261);
nor U15898 (N_15898,N_14432,N_14020);
nand U15899 (N_15899,N_14514,N_14584);
nand U15900 (N_15900,N_14931,N_14216);
nor U15901 (N_15901,N_14304,N_14957);
nor U15902 (N_15902,N_14384,N_14109);
nor U15903 (N_15903,N_14659,N_14833);
nand U15904 (N_15904,N_14182,N_14687);
and U15905 (N_15905,N_14519,N_14246);
nand U15906 (N_15906,N_14815,N_14730);
nand U15907 (N_15907,N_14418,N_14621);
or U15908 (N_15908,N_14381,N_14235);
or U15909 (N_15909,N_14715,N_14335);
and U15910 (N_15910,N_14484,N_14333);
or U15911 (N_15911,N_14343,N_14161);
xor U15912 (N_15912,N_14747,N_14143);
or U15913 (N_15913,N_14893,N_14592);
nand U15914 (N_15914,N_14200,N_14304);
nand U15915 (N_15915,N_14570,N_14548);
or U15916 (N_15916,N_14194,N_14332);
or U15917 (N_15917,N_14857,N_14168);
and U15918 (N_15918,N_14117,N_14205);
or U15919 (N_15919,N_14807,N_14830);
xnor U15920 (N_15920,N_14356,N_14370);
and U15921 (N_15921,N_14758,N_14811);
nand U15922 (N_15922,N_14780,N_14009);
and U15923 (N_15923,N_14081,N_14508);
xor U15924 (N_15924,N_14625,N_14800);
nand U15925 (N_15925,N_14636,N_14506);
and U15926 (N_15926,N_14744,N_14499);
nand U15927 (N_15927,N_14735,N_14861);
nor U15928 (N_15928,N_14293,N_14929);
or U15929 (N_15929,N_14870,N_14703);
xor U15930 (N_15930,N_14426,N_14717);
or U15931 (N_15931,N_14385,N_14052);
nor U15932 (N_15932,N_14808,N_14120);
nor U15933 (N_15933,N_14113,N_14996);
nor U15934 (N_15934,N_14845,N_14716);
xnor U15935 (N_15935,N_14152,N_14998);
xnor U15936 (N_15936,N_14891,N_14881);
or U15937 (N_15937,N_14514,N_14286);
nand U15938 (N_15938,N_14734,N_14473);
nand U15939 (N_15939,N_14006,N_14647);
nand U15940 (N_15940,N_14716,N_14540);
nand U15941 (N_15941,N_14449,N_14493);
and U15942 (N_15942,N_14771,N_14174);
nand U15943 (N_15943,N_14662,N_14076);
nand U15944 (N_15944,N_14302,N_14656);
nand U15945 (N_15945,N_14409,N_14418);
and U15946 (N_15946,N_14382,N_14663);
nand U15947 (N_15947,N_14483,N_14659);
or U15948 (N_15948,N_14345,N_14597);
or U15949 (N_15949,N_14927,N_14536);
nor U15950 (N_15950,N_14319,N_14118);
nand U15951 (N_15951,N_14899,N_14785);
nor U15952 (N_15952,N_14135,N_14623);
or U15953 (N_15953,N_14361,N_14430);
nor U15954 (N_15954,N_14132,N_14424);
nand U15955 (N_15955,N_14309,N_14768);
nor U15956 (N_15956,N_14342,N_14252);
nor U15957 (N_15957,N_14325,N_14217);
or U15958 (N_15958,N_14461,N_14120);
or U15959 (N_15959,N_14140,N_14476);
nor U15960 (N_15960,N_14532,N_14125);
or U15961 (N_15961,N_14833,N_14308);
nand U15962 (N_15962,N_14185,N_14260);
and U15963 (N_15963,N_14621,N_14196);
xnor U15964 (N_15964,N_14803,N_14347);
nand U15965 (N_15965,N_14477,N_14379);
and U15966 (N_15966,N_14329,N_14131);
and U15967 (N_15967,N_14325,N_14398);
nand U15968 (N_15968,N_14842,N_14911);
nor U15969 (N_15969,N_14663,N_14524);
nand U15970 (N_15970,N_14719,N_14273);
nand U15971 (N_15971,N_14731,N_14313);
xor U15972 (N_15972,N_14847,N_14760);
and U15973 (N_15973,N_14210,N_14898);
and U15974 (N_15974,N_14477,N_14883);
and U15975 (N_15975,N_14774,N_14004);
or U15976 (N_15976,N_14471,N_14250);
nor U15977 (N_15977,N_14401,N_14187);
nor U15978 (N_15978,N_14748,N_14151);
or U15979 (N_15979,N_14893,N_14633);
nor U15980 (N_15980,N_14407,N_14993);
nor U15981 (N_15981,N_14747,N_14279);
nor U15982 (N_15982,N_14355,N_14025);
nor U15983 (N_15983,N_14722,N_14785);
nand U15984 (N_15984,N_14622,N_14270);
nor U15985 (N_15985,N_14171,N_14497);
nand U15986 (N_15986,N_14853,N_14596);
nand U15987 (N_15987,N_14625,N_14579);
nand U15988 (N_15988,N_14362,N_14617);
and U15989 (N_15989,N_14485,N_14279);
xnor U15990 (N_15990,N_14648,N_14061);
or U15991 (N_15991,N_14079,N_14387);
or U15992 (N_15992,N_14284,N_14940);
or U15993 (N_15993,N_14799,N_14589);
xnor U15994 (N_15994,N_14024,N_14537);
nor U15995 (N_15995,N_14101,N_14572);
nand U15996 (N_15996,N_14783,N_14049);
or U15997 (N_15997,N_14417,N_14152);
nor U15998 (N_15998,N_14719,N_14546);
or U15999 (N_15999,N_14673,N_14155);
nor U16000 (N_16000,N_15307,N_15376);
xnor U16001 (N_16001,N_15859,N_15914);
nor U16002 (N_16002,N_15576,N_15401);
and U16003 (N_16003,N_15662,N_15447);
nand U16004 (N_16004,N_15711,N_15897);
nand U16005 (N_16005,N_15125,N_15282);
or U16006 (N_16006,N_15552,N_15203);
nor U16007 (N_16007,N_15575,N_15237);
xnor U16008 (N_16008,N_15391,N_15500);
xnor U16009 (N_16009,N_15275,N_15337);
or U16010 (N_16010,N_15033,N_15315);
and U16011 (N_16011,N_15398,N_15143);
or U16012 (N_16012,N_15189,N_15541);
nand U16013 (N_16013,N_15122,N_15034);
xnor U16014 (N_16014,N_15329,N_15661);
xor U16015 (N_16015,N_15226,N_15073);
xor U16016 (N_16016,N_15865,N_15596);
and U16017 (N_16017,N_15412,N_15499);
or U16018 (N_16018,N_15011,N_15909);
or U16019 (N_16019,N_15736,N_15172);
nand U16020 (N_16020,N_15548,N_15845);
or U16021 (N_16021,N_15363,N_15180);
or U16022 (N_16022,N_15631,N_15165);
nand U16023 (N_16023,N_15389,N_15649);
or U16024 (N_16024,N_15557,N_15940);
nand U16025 (N_16025,N_15015,N_15078);
nor U16026 (N_16026,N_15217,N_15680);
nand U16027 (N_16027,N_15793,N_15258);
or U16028 (N_16028,N_15072,N_15799);
nand U16029 (N_16029,N_15096,N_15382);
xnor U16030 (N_16030,N_15050,N_15651);
xor U16031 (N_16031,N_15002,N_15469);
nor U16032 (N_16032,N_15092,N_15215);
nand U16033 (N_16033,N_15335,N_15403);
and U16034 (N_16034,N_15898,N_15147);
xor U16035 (N_16035,N_15957,N_15434);
nor U16036 (N_16036,N_15212,N_15229);
nand U16037 (N_16037,N_15842,N_15966);
nand U16038 (N_16038,N_15587,N_15350);
and U16039 (N_16039,N_15824,N_15027);
or U16040 (N_16040,N_15378,N_15234);
or U16041 (N_16041,N_15357,N_15452);
or U16042 (N_16042,N_15760,N_15747);
nand U16043 (N_16043,N_15303,N_15681);
or U16044 (N_16044,N_15106,N_15326);
nor U16045 (N_16045,N_15114,N_15042);
nor U16046 (N_16046,N_15394,N_15851);
nand U16047 (N_16047,N_15669,N_15145);
nor U16048 (N_16048,N_15956,N_15813);
or U16049 (N_16049,N_15100,N_15365);
nor U16050 (N_16050,N_15570,N_15495);
or U16051 (N_16051,N_15969,N_15513);
or U16052 (N_16052,N_15573,N_15103);
and U16053 (N_16053,N_15512,N_15444);
xnor U16054 (N_16054,N_15985,N_15392);
xor U16055 (N_16055,N_15302,N_15084);
nand U16056 (N_16056,N_15857,N_15617);
nand U16057 (N_16057,N_15435,N_15673);
and U16058 (N_16058,N_15525,N_15387);
xor U16059 (N_16059,N_15257,N_15546);
or U16060 (N_16060,N_15700,N_15150);
nand U16061 (N_16061,N_15724,N_15727);
or U16062 (N_16062,N_15827,N_15210);
nor U16063 (N_16063,N_15101,N_15655);
nor U16064 (N_16064,N_15549,N_15503);
or U16065 (N_16065,N_15584,N_15924);
and U16066 (N_16066,N_15031,N_15578);
nand U16067 (N_16067,N_15498,N_15107);
or U16068 (N_16068,N_15074,N_15944);
xnor U16069 (N_16069,N_15721,N_15798);
or U16070 (N_16070,N_15480,N_15136);
nor U16071 (N_16071,N_15884,N_15244);
xnor U16072 (N_16072,N_15064,N_15243);
xnor U16073 (N_16073,N_15225,N_15777);
or U16074 (N_16074,N_15466,N_15082);
and U16075 (N_16075,N_15019,N_15952);
nor U16076 (N_16076,N_15682,N_15818);
xnor U16077 (N_16077,N_15192,N_15671);
xnor U16078 (N_16078,N_15115,N_15975);
nand U16079 (N_16079,N_15872,N_15339);
or U16080 (N_16080,N_15611,N_15327);
and U16081 (N_16081,N_15691,N_15044);
xor U16082 (N_16082,N_15364,N_15685);
or U16083 (N_16083,N_15087,N_15920);
xnor U16084 (N_16084,N_15272,N_15762);
or U16085 (N_16085,N_15051,N_15245);
nand U16086 (N_16086,N_15756,N_15524);
nand U16087 (N_16087,N_15693,N_15585);
xor U16088 (N_16088,N_15062,N_15520);
nor U16089 (N_16089,N_15853,N_15869);
xnor U16090 (N_16090,N_15208,N_15195);
or U16091 (N_16091,N_15726,N_15953);
and U16092 (N_16092,N_15522,N_15336);
or U16093 (N_16093,N_15773,N_15406);
xnor U16094 (N_16094,N_15417,N_15252);
and U16095 (N_16095,N_15241,N_15105);
nand U16096 (N_16096,N_15852,N_15858);
nor U16097 (N_16097,N_15936,N_15769);
and U16098 (N_16098,N_15663,N_15407);
or U16099 (N_16099,N_15046,N_15181);
or U16100 (N_16100,N_15636,N_15856);
or U16101 (N_16101,N_15763,N_15986);
and U16102 (N_16102,N_15113,N_15193);
or U16103 (N_16103,N_15104,N_15487);
nand U16104 (N_16104,N_15345,N_15201);
xnor U16105 (N_16105,N_15477,N_15607);
xnor U16106 (N_16106,N_15875,N_15514);
or U16107 (N_16107,N_15534,N_15890);
nor U16108 (N_16108,N_15360,N_15259);
xor U16109 (N_16109,N_15112,N_15397);
and U16110 (N_16110,N_15701,N_15999);
xnor U16111 (N_16111,N_15830,N_15788);
or U16112 (N_16112,N_15964,N_15005);
nand U16113 (N_16113,N_15960,N_15137);
nor U16114 (N_16114,N_15504,N_15517);
or U16115 (N_16115,N_15348,N_15040);
nor U16116 (N_16116,N_15565,N_15039);
and U16117 (N_16117,N_15152,N_15057);
nor U16118 (N_16118,N_15874,N_15656);
and U16119 (N_16119,N_15288,N_15901);
nand U16120 (N_16120,N_15146,N_15566);
nand U16121 (N_16121,N_15831,N_15463);
or U16122 (N_16122,N_15130,N_15950);
xnor U16123 (N_16123,N_15413,N_15320);
xor U16124 (N_16124,N_15630,N_15714);
or U16125 (N_16125,N_15729,N_15010);
and U16126 (N_16126,N_15812,N_15863);
nand U16127 (N_16127,N_15294,N_15965);
nor U16128 (N_16128,N_15523,N_15984);
nand U16129 (N_16129,N_15732,N_15371);
nor U16130 (N_16130,N_15554,N_15695);
or U16131 (N_16131,N_15908,N_15070);
nand U16132 (N_16132,N_15943,N_15766);
and U16133 (N_16133,N_15892,N_15422);
xnor U16134 (N_16134,N_15713,N_15855);
nand U16135 (N_16135,N_15543,N_15870);
nor U16136 (N_16136,N_15755,N_15730);
or U16137 (N_16137,N_15608,N_15542);
or U16138 (N_16138,N_15415,N_15931);
and U16139 (N_16139,N_15474,N_15705);
and U16140 (N_16140,N_15481,N_15020);
or U16141 (N_16141,N_15707,N_15962);
or U16142 (N_16142,N_15638,N_15518);
nor U16143 (N_16143,N_15582,N_15988);
nand U16144 (N_16144,N_15399,N_15485);
and U16145 (N_16145,N_15922,N_15409);
and U16146 (N_16146,N_15102,N_15742);
nor U16147 (N_16147,N_15910,N_15323);
nand U16148 (N_16148,N_15928,N_15016);
or U16149 (N_16149,N_15774,N_15047);
and U16150 (N_16150,N_15614,N_15054);
and U16151 (N_16151,N_15262,N_15841);
and U16152 (N_16152,N_15359,N_15610);
or U16153 (N_16153,N_15847,N_15982);
or U16154 (N_16154,N_15176,N_15194);
nor U16155 (N_16155,N_15296,N_15531);
xor U16156 (N_16156,N_15540,N_15380);
xnor U16157 (N_16157,N_15483,N_15731);
nor U16158 (N_16158,N_15741,N_15438);
or U16159 (N_16159,N_15796,N_15697);
nand U16160 (N_16160,N_15672,N_15496);
nor U16161 (N_16161,N_15058,N_15589);
or U16162 (N_16162,N_15598,N_15489);
xor U16163 (N_16163,N_15306,N_15206);
nor U16164 (N_16164,N_15955,N_15224);
or U16165 (N_16165,N_15822,N_15634);
nor U16166 (N_16166,N_15604,N_15954);
and U16167 (N_16167,N_15390,N_15556);
nand U16168 (N_16168,N_15439,N_15289);
nor U16169 (N_16169,N_15699,N_15709);
nor U16170 (N_16170,N_15561,N_15008);
and U16171 (N_16171,N_15053,N_15287);
nor U16172 (N_16172,N_15923,N_15349);
or U16173 (N_16173,N_15222,N_15618);
and U16174 (N_16174,N_15751,N_15187);
nor U16175 (N_16175,N_15249,N_15242);
nand U16176 (N_16176,N_15024,N_15200);
xor U16177 (N_16177,N_15377,N_15746);
nand U16178 (N_16178,N_15416,N_15227);
nand U16179 (N_16179,N_15564,N_15128);
xor U16180 (N_16180,N_15052,N_15472);
or U16181 (N_16181,N_15911,N_15720);
nor U16182 (N_16182,N_15981,N_15285);
or U16183 (N_16183,N_15632,N_15299);
and U16184 (N_16184,N_15324,N_15828);
xor U16185 (N_16185,N_15595,N_15116);
xor U16186 (N_16186,N_15097,N_15490);
or U16187 (N_16187,N_15509,N_15133);
or U16188 (N_16188,N_15580,N_15939);
or U16189 (N_16189,N_15419,N_15846);
or U16190 (N_16190,N_15642,N_15160);
and U16191 (N_16191,N_15178,N_15085);
xor U16192 (N_16192,N_15148,N_15627);
xnor U16193 (N_16193,N_15161,N_15854);
nor U16194 (N_16194,N_15220,N_15980);
or U16195 (N_16195,N_15974,N_15805);
xnor U16196 (N_16196,N_15369,N_15740);
and U16197 (N_16197,N_15450,N_15779);
and U16198 (N_16198,N_15667,N_15384);
nand U16199 (N_16199,N_15712,N_15574);
or U16200 (N_16200,N_15135,N_15139);
or U16201 (N_16201,N_15658,N_15400);
nor U16202 (N_16202,N_15291,N_15759);
xor U16203 (N_16203,N_15300,N_15381);
and U16204 (N_16204,N_15433,N_15597);
and U16205 (N_16205,N_15319,N_15196);
or U16206 (N_16206,N_15022,N_15163);
or U16207 (N_16207,N_15159,N_15479);
and U16208 (N_16208,N_15037,N_15836);
xnor U16209 (N_16209,N_15312,N_15946);
nand U16210 (N_16210,N_15431,N_15571);
or U16211 (N_16211,N_15963,N_15265);
and U16212 (N_16212,N_15603,N_15421);
nand U16213 (N_16213,N_15794,N_15427);
or U16214 (N_16214,N_15674,N_15018);
nor U16215 (N_16215,N_15716,N_15157);
and U16216 (N_16216,N_15209,N_15676);
and U16217 (N_16217,N_15023,N_15079);
nor U16218 (N_16218,N_15095,N_15971);
nor U16219 (N_16219,N_15190,N_15000);
nand U16220 (N_16220,N_15448,N_15094);
nor U16221 (N_16221,N_15840,N_15132);
and U16222 (N_16222,N_15932,N_15801);
nand U16223 (N_16223,N_15167,N_15017);
nor U16224 (N_16224,N_15995,N_15248);
nor U16225 (N_16225,N_15886,N_15735);
nand U16226 (N_16226,N_15155,N_15366);
xor U16227 (N_16227,N_15110,N_15123);
xor U16228 (N_16228,N_15199,N_15213);
nor U16229 (N_16229,N_15835,N_15436);
nand U16230 (N_16230,N_15041,N_15532);
and U16231 (N_16231,N_15492,N_15907);
nand U16232 (N_16232,N_15346,N_15362);
xnor U16233 (N_16233,N_15071,N_15344);
nand U16234 (N_16234,N_15506,N_15205);
or U16235 (N_16235,N_15888,N_15792);
and U16236 (N_16236,N_15823,N_15887);
nand U16237 (N_16237,N_15588,N_15916);
nand U16238 (N_16238,N_15216,N_15470);
nor U16239 (N_16239,N_15972,N_15451);
xnor U16240 (N_16240,N_15098,N_15283);
and U16241 (N_16241,N_15592,N_15849);
and U16242 (N_16242,N_15606,N_15586);
xor U16243 (N_16243,N_15266,N_15816);
nor U16244 (N_16244,N_15202,N_15273);
or U16245 (N_16245,N_15725,N_15410);
nand U16246 (N_16246,N_15353,N_15544);
xor U16247 (N_16247,N_15679,N_15211);
or U16248 (N_16248,N_15219,N_15325);
xor U16249 (N_16249,N_15704,N_15441);
xor U16250 (N_16250,N_15622,N_15423);
nand U16251 (N_16251,N_15838,N_15906);
nand U16252 (N_16252,N_15083,N_15035);
nand U16253 (N_16253,N_15183,N_15281);
and U16254 (N_16254,N_15445,N_15060);
or U16255 (N_16255,N_15295,N_15065);
nand U16256 (N_16256,N_15625,N_15298);
and U16257 (N_16257,N_15577,N_15293);
nand U16258 (N_16258,N_15151,N_15328);
xnor U16259 (N_16259,N_15331,N_15129);
or U16260 (N_16260,N_15977,N_15066);
nor U16261 (N_16261,N_15921,N_15516);
and U16262 (N_16262,N_15119,N_15383);
nor U16263 (N_16263,N_15635,N_15987);
xor U16264 (N_16264,N_15260,N_15684);
nor U16265 (N_16265,N_15292,N_15269);
xor U16266 (N_16266,N_15510,N_15231);
nor U16267 (N_16267,N_15804,N_15169);
nor U16268 (N_16268,N_15026,N_15207);
or U16269 (N_16269,N_15765,N_15395);
nor U16270 (N_16270,N_15782,N_15028);
nand U16271 (N_16271,N_15996,N_15430);
and U16272 (N_16272,N_15743,N_15473);
or U16273 (N_16273,N_15068,N_15733);
and U16274 (N_16274,N_15748,N_15758);
xor U16275 (N_16275,N_15528,N_15917);
xnor U16276 (N_16276,N_15454,N_15710);
nor U16277 (N_16277,N_15218,N_15049);
and U16278 (N_16278,N_15059,N_15958);
nand U16279 (N_16279,N_15501,N_15278);
or U16280 (N_16280,N_15621,N_15305);
nor U16281 (N_16281,N_15505,N_15690);
nor U16282 (N_16282,N_15581,N_15829);
xor U16283 (N_16283,N_15388,N_15785);
nor U16284 (N_16284,N_15333,N_15223);
nand U16285 (N_16285,N_15553,N_15609);
nand U16286 (N_16286,N_15239,N_15286);
and U16287 (N_16287,N_15330,N_15791);
nand U16288 (N_16288,N_15453,N_15640);
and U16289 (N_16289,N_15264,N_15519);
xor U16290 (N_16290,N_15069,N_15012);
nand U16291 (N_16291,N_15770,N_15386);
or U16292 (N_16292,N_15004,N_15014);
nor U16293 (N_16293,N_15343,N_15781);
xor U16294 (N_16294,N_15032,N_15411);
and U16295 (N_16295,N_15698,N_15795);
nor U16296 (N_16296,N_15772,N_15692);
or U16297 (N_16297,N_15935,N_15476);
nor U16298 (N_16298,N_15455,N_15141);
xor U16299 (N_16299,N_15468,N_15990);
nor U16300 (N_16300,N_15738,N_15081);
nand U16301 (N_16301,N_15153,N_15089);
nand U16302 (N_16302,N_15170,N_15536);
nand U16303 (N_16303,N_15666,N_15899);
nor U16304 (N_16304,N_15228,N_15277);
xor U16305 (N_16305,N_15494,N_15332);
or U16306 (N_16306,N_15437,N_15605);
or U16307 (N_16307,N_15654,N_15356);
or U16308 (N_16308,N_15358,N_15652);
nor U16309 (N_16309,N_15379,N_15086);
nand U16310 (N_16310,N_15744,N_15117);
xnor U16311 (N_16311,N_15511,N_15091);
nand U16312 (N_16312,N_15030,N_15317);
xnor U16313 (N_16313,N_15374,N_15256);
xnor U16314 (N_16314,N_15013,N_15590);
and U16315 (N_16315,N_15650,N_15970);
nor U16316 (N_16316,N_15568,N_15061);
nor U16317 (N_16317,N_15547,N_15706);
xor U16318 (N_16318,N_15694,N_15983);
xnor U16319 (N_16319,N_15164,N_15367);
or U16320 (N_16320,N_15402,N_15373);
xnor U16321 (N_16321,N_15290,N_15967);
or U16322 (N_16322,N_15108,N_15310);
nand U16323 (N_16323,N_15904,N_15961);
nor U16324 (N_16324,N_15639,N_15230);
and U16325 (N_16325,N_15768,N_15168);
and U16326 (N_16326,N_15664,N_15342);
and U16327 (N_16327,N_15775,N_15815);
xnor U16328 (N_16328,N_15643,N_15121);
and U16329 (N_16329,N_15807,N_15530);
xnor U16330 (N_16330,N_15708,N_15602);
xor U16331 (N_16331,N_15533,N_15814);
and U16332 (N_16332,N_15029,N_15443);
xor U16333 (N_16333,N_15717,N_15653);
or U16334 (N_16334,N_15340,N_15959);
and U16335 (N_16335,N_15800,N_15526);
xor U16336 (N_16336,N_15308,N_15126);
xor U16337 (N_16337,N_15236,N_15545);
or U16338 (N_16338,N_15703,N_15926);
nand U16339 (N_16339,N_15626,N_15109);
and U16340 (N_16340,N_15594,N_15127);
or U16341 (N_16341,N_15043,N_15745);
xnor U16342 (N_16342,N_15396,N_15003);
xnor U16343 (N_16343,N_15214,N_15687);
or U16344 (N_16344,N_15997,N_15255);
or U16345 (N_16345,N_15826,N_15761);
xnor U16346 (N_16346,N_15502,N_15537);
nor U16347 (N_16347,N_15894,N_15280);
xnor U16348 (N_16348,N_15461,N_15560);
and U16349 (N_16349,N_15880,N_15825);
xor U16350 (N_16350,N_15124,N_15832);
or U16351 (N_16351,N_15036,N_15790);
nor U16352 (N_16352,N_15426,N_15877);
nand U16353 (N_16353,N_15462,N_15460);
nor U16354 (N_16354,N_15111,N_15171);
nor U16355 (N_16355,N_15428,N_15601);
nand U16356 (N_16356,N_15771,N_15787);
xor U16357 (N_16357,N_15456,N_15808);
or U16358 (N_16358,N_15633,N_15188);
or U16359 (N_16359,N_15620,N_15696);
nor U16360 (N_16360,N_15767,N_15254);
and U16361 (N_16361,N_15048,N_15271);
nand U16362 (N_16362,N_15757,N_15080);
nor U16363 (N_16363,N_15197,N_15878);
and U16364 (N_16364,N_15896,N_15951);
and U16365 (N_16365,N_15156,N_15821);
or U16366 (N_16366,N_15600,N_15871);
and U16367 (N_16367,N_15994,N_15860);
nand U16368 (N_16368,N_15361,N_15702);
nand U16369 (N_16369,N_15688,N_15240);
xor U16370 (N_16370,N_15613,N_15491);
nor U16371 (N_16371,N_15488,N_15616);
xor U16372 (N_16372,N_15629,N_15891);
and U16373 (N_16373,N_15583,N_15645);
and U16374 (N_16374,N_15021,N_15425);
xor U16375 (N_16375,N_15780,N_15442);
nand U16376 (N_16376,N_15045,N_15833);
and U16377 (N_16377,N_15677,N_15446);
xor U16378 (N_16378,N_15569,N_15998);
nand U16379 (N_16379,N_15868,N_15263);
nor U16380 (N_16380,N_15593,N_15558);
or U16381 (N_16381,N_15001,N_15885);
nand U16382 (N_16382,N_15976,N_15099);
nand U16383 (N_16383,N_15120,N_15862);
xnor U16384 (N_16384,N_15778,N_15251);
and U16385 (N_16385,N_15322,N_15551);
or U16386 (N_16386,N_15038,N_15819);
and U16387 (N_16387,N_15175,N_15486);
and U16388 (N_16388,N_15075,N_15134);
nand U16389 (N_16389,N_15311,N_15493);
xnor U16390 (N_16390,N_15246,N_15848);
or U16391 (N_16391,N_15783,N_15405);
nor U16392 (N_16392,N_15076,N_15198);
nor U16393 (N_16393,N_15478,N_15338);
nand U16394 (N_16394,N_15191,N_15689);
xor U16395 (N_16395,N_15131,N_15408);
xor U16396 (N_16396,N_15615,N_15683);
or U16397 (N_16397,N_15186,N_15056);
xor U16398 (N_16398,N_15508,N_15185);
nand U16399 (N_16399,N_15088,N_15660);
or U16400 (N_16400,N_15945,N_15458);
nand U16401 (N_16401,N_15806,N_15393);
nor U16402 (N_16402,N_15538,N_15728);
nand U16403 (N_16403,N_15929,N_15321);
and U16404 (N_16404,N_15686,N_15232);
nor U16405 (N_16405,N_15784,N_15723);
nor U16406 (N_16406,N_15883,N_15465);
nor U16407 (N_16407,N_15612,N_15449);
or U16408 (N_16408,N_15007,N_15341);
or U16409 (N_16409,N_15839,N_15949);
xor U16410 (N_16410,N_15077,N_15802);
or U16411 (N_16411,N_15253,N_15385);
nor U16412 (N_16412,N_15934,N_15475);
xor U16413 (N_16413,N_15515,N_15313);
xnor U16414 (N_16414,N_15314,N_15803);
nor U16415 (N_16415,N_15753,N_15347);
nand U16416 (N_16416,N_15093,N_15900);
or U16417 (N_16417,N_15250,N_15719);
or U16418 (N_16418,N_15641,N_15279);
and U16419 (N_16419,N_15989,N_15850);
xnor U16420 (N_16420,N_15429,N_15866);
or U16421 (N_16421,N_15734,N_15550);
or U16422 (N_16422,N_15591,N_15876);
or U16423 (N_16423,N_15567,N_15309);
nand U16424 (N_16424,N_15284,N_15267);
nand U16425 (N_16425,N_15370,N_15179);
and U16426 (N_16426,N_15467,N_15154);
nor U16427 (N_16427,N_15067,N_15233);
xor U16428 (N_16428,N_15810,N_15993);
or U16429 (N_16429,N_15118,N_15235);
or U16430 (N_16430,N_15572,N_15276);
or U16431 (N_16431,N_15665,N_15318);
nand U16432 (N_16432,N_15529,N_15912);
or U16433 (N_16433,N_15668,N_15268);
nand U16434 (N_16434,N_15375,N_15947);
xnor U16435 (N_16435,N_15140,N_15274);
nand U16436 (N_16436,N_15930,N_15301);
or U16437 (N_16437,N_15882,N_15174);
xnor U16438 (N_16438,N_15404,N_15352);
xnor U16439 (N_16439,N_15457,N_15881);
and U16440 (N_16440,N_15809,N_15166);
nand U16441 (N_16441,N_15913,N_15817);
and U16442 (N_16442,N_15937,N_15978);
nand U16443 (N_16443,N_15484,N_15424);
or U16444 (N_16444,N_15895,N_15162);
and U16445 (N_16445,N_15979,N_15905);
and U16446 (N_16446,N_15418,N_15142);
xor U16447 (N_16447,N_15628,N_15304);
or U16448 (N_16448,N_15414,N_15925);
nor U16449 (N_16449,N_15579,N_15138);
xnor U16450 (N_16450,N_15055,N_15948);
or U16451 (N_16451,N_15521,N_15739);
and U16452 (N_16452,N_15599,N_15973);
nand U16453 (N_16453,N_15555,N_15722);
and U16454 (N_16454,N_15659,N_15497);
xor U16455 (N_16455,N_15619,N_15090);
nand U16456 (N_16456,N_15843,N_15992);
and U16457 (N_16457,N_15471,N_15942);
xnor U16458 (N_16458,N_15919,N_15879);
nand U16459 (N_16459,N_15355,N_15440);
and U16460 (N_16460,N_15184,N_15811);
nand U16461 (N_16461,N_15368,N_15718);
nor U16462 (N_16462,N_15351,N_15025);
nand U16463 (N_16463,N_15623,N_15507);
and U16464 (N_16464,N_15991,N_15786);
nand U16465 (N_16465,N_15754,N_15789);
nand U16466 (N_16466,N_15776,N_15637);
and U16467 (N_16467,N_15837,N_15624);
or U16468 (N_16468,N_15562,N_15902);
or U16469 (N_16469,N_15354,N_15873);
and U16470 (N_16470,N_15563,N_15648);
nor U16471 (N_16471,N_15715,N_15535);
or U16472 (N_16472,N_15764,N_15432);
and U16473 (N_16473,N_15675,N_15158);
xnor U16474 (N_16474,N_15646,N_15903);
xor U16475 (N_16475,N_15861,N_15297);
and U16476 (N_16476,N_15539,N_15247);
nand U16477 (N_16477,N_15173,N_15559);
xor U16478 (N_16478,N_15657,N_15149);
and U16479 (N_16479,N_15316,N_15915);
and U16480 (N_16480,N_15270,N_15221);
xnor U16481 (N_16481,N_15238,N_15261);
nand U16482 (N_16482,N_15752,N_15006);
nor U16483 (N_16483,N_15464,N_15334);
nor U16484 (N_16484,N_15647,N_15527);
xor U16485 (N_16485,N_15177,N_15678);
nor U16486 (N_16486,N_15938,N_15737);
nor U16487 (N_16487,N_15893,N_15372);
or U16488 (N_16488,N_15144,N_15063);
nor U16489 (N_16489,N_15670,N_15844);
nand U16490 (N_16490,N_15927,N_15834);
or U16491 (N_16491,N_15968,N_15644);
or U16492 (N_16492,N_15820,N_15918);
and U16493 (N_16493,N_15749,N_15941);
xor U16494 (N_16494,N_15864,N_15889);
nor U16495 (N_16495,N_15182,N_15009);
xor U16496 (N_16496,N_15867,N_15750);
nand U16497 (N_16497,N_15933,N_15797);
xor U16498 (N_16498,N_15459,N_15204);
nor U16499 (N_16499,N_15420,N_15482);
xnor U16500 (N_16500,N_15343,N_15279);
and U16501 (N_16501,N_15213,N_15472);
xnor U16502 (N_16502,N_15185,N_15835);
xnor U16503 (N_16503,N_15641,N_15623);
or U16504 (N_16504,N_15270,N_15520);
and U16505 (N_16505,N_15028,N_15290);
xnor U16506 (N_16506,N_15169,N_15376);
xor U16507 (N_16507,N_15577,N_15689);
xnor U16508 (N_16508,N_15743,N_15249);
nor U16509 (N_16509,N_15525,N_15862);
or U16510 (N_16510,N_15728,N_15227);
and U16511 (N_16511,N_15475,N_15742);
nor U16512 (N_16512,N_15793,N_15581);
or U16513 (N_16513,N_15470,N_15921);
and U16514 (N_16514,N_15981,N_15379);
and U16515 (N_16515,N_15603,N_15988);
nor U16516 (N_16516,N_15667,N_15689);
nand U16517 (N_16517,N_15593,N_15391);
nand U16518 (N_16518,N_15052,N_15124);
xor U16519 (N_16519,N_15853,N_15283);
and U16520 (N_16520,N_15096,N_15421);
xor U16521 (N_16521,N_15041,N_15168);
and U16522 (N_16522,N_15647,N_15346);
and U16523 (N_16523,N_15579,N_15029);
or U16524 (N_16524,N_15131,N_15673);
or U16525 (N_16525,N_15249,N_15810);
or U16526 (N_16526,N_15137,N_15970);
xor U16527 (N_16527,N_15065,N_15474);
or U16528 (N_16528,N_15736,N_15392);
nor U16529 (N_16529,N_15170,N_15778);
nor U16530 (N_16530,N_15250,N_15228);
nor U16531 (N_16531,N_15659,N_15730);
nor U16532 (N_16532,N_15623,N_15214);
xnor U16533 (N_16533,N_15409,N_15632);
xor U16534 (N_16534,N_15081,N_15584);
or U16535 (N_16535,N_15938,N_15873);
nor U16536 (N_16536,N_15245,N_15003);
xnor U16537 (N_16537,N_15320,N_15466);
nand U16538 (N_16538,N_15349,N_15191);
nor U16539 (N_16539,N_15127,N_15192);
xnor U16540 (N_16540,N_15656,N_15075);
xor U16541 (N_16541,N_15747,N_15688);
nor U16542 (N_16542,N_15466,N_15628);
xnor U16543 (N_16543,N_15066,N_15898);
or U16544 (N_16544,N_15296,N_15056);
nor U16545 (N_16545,N_15037,N_15679);
and U16546 (N_16546,N_15693,N_15769);
nor U16547 (N_16547,N_15489,N_15102);
nor U16548 (N_16548,N_15835,N_15524);
nor U16549 (N_16549,N_15170,N_15811);
or U16550 (N_16550,N_15026,N_15456);
or U16551 (N_16551,N_15133,N_15349);
or U16552 (N_16552,N_15509,N_15046);
or U16553 (N_16553,N_15123,N_15023);
nand U16554 (N_16554,N_15126,N_15369);
xnor U16555 (N_16555,N_15719,N_15692);
or U16556 (N_16556,N_15541,N_15256);
and U16557 (N_16557,N_15303,N_15494);
nor U16558 (N_16558,N_15128,N_15568);
xor U16559 (N_16559,N_15511,N_15823);
or U16560 (N_16560,N_15398,N_15537);
nand U16561 (N_16561,N_15576,N_15743);
xnor U16562 (N_16562,N_15862,N_15647);
or U16563 (N_16563,N_15052,N_15992);
nand U16564 (N_16564,N_15228,N_15497);
nand U16565 (N_16565,N_15830,N_15317);
nand U16566 (N_16566,N_15390,N_15398);
and U16567 (N_16567,N_15155,N_15225);
and U16568 (N_16568,N_15161,N_15270);
or U16569 (N_16569,N_15396,N_15026);
nor U16570 (N_16570,N_15139,N_15307);
and U16571 (N_16571,N_15804,N_15845);
nor U16572 (N_16572,N_15690,N_15196);
nor U16573 (N_16573,N_15732,N_15143);
nand U16574 (N_16574,N_15599,N_15665);
or U16575 (N_16575,N_15768,N_15896);
nand U16576 (N_16576,N_15626,N_15879);
or U16577 (N_16577,N_15069,N_15769);
nor U16578 (N_16578,N_15946,N_15344);
xor U16579 (N_16579,N_15414,N_15865);
xnor U16580 (N_16580,N_15064,N_15728);
or U16581 (N_16581,N_15678,N_15416);
nor U16582 (N_16582,N_15623,N_15600);
nand U16583 (N_16583,N_15881,N_15199);
nor U16584 (N_16584,N_15652,N_15330);
xnor U16585 (N_16585,N_15149,N_15019);
xnor U16586 (N_16586,N_15175,N_15179);
nor U16587 (N_16587,N_15977,N_15292);
nor U16588 (N_16588,N_15607,N_15867);
nand U16589 (N_16589,N_15405,N_15917);
xor U16590 (N_16590,N_15297,N_15341);
and U16591 (N_16591,N_15778,N_15983);
or U16592 (N_16592,N_15015,N_15318);
xnor U16593 (N_16593,N_15050,N_15095);
and U16594 (N_16594,N_15294,N_15208);
nand U16595 (N_16595,N_15400,N_15179);
or U16596 (N_16596,N_15280,N_15686);
nor U16597 (N_16597,N_15685,N_15835);
or U16598 (N_16598,N_15025,N_15386);
and U16599 (N_16599,N_15592,N_15640);
xor U16600 (N_16600,N_15770,N_15304);
xnor U16601 (N_16601,N_15556,N_15778);
xnor U16602 (N_16602,N_15715,N_15079);
and U16603 (N_16603,N_15481,N_15910);
or U16604 (N_16604,N_15430,N_15231);
nor U16605 (N_16605,N_15686,N_15115);
and U16606 (N_16606,N_15460,N_15288);
xnor U16607 (N_16607,N_15589,N_15092);
xor U16608 (N_16608,N_15349,N_15155);
xnor U16609 (N_16609,N_15775,N_15187);
and U16610 (N_16610,N_15977,N_15072);
and U16611 (N_16611,N_15517,N_15934);
xor U16612 (N_16612,N_15556,N_15343);
and U16613 (N_16613,N_15157,N_15458);
nor U16614 (N_16614,N_15868,N_15430);
and U16615 (N_16615,N_15426,N_15003);
nor U16616 (N_16616,N_15578,N_15817);
nor U16617 (N_16617,N_15256,N_15817);
xor U16618 (N_16618,N_15293,N_15610);
or U16619 (N_16619,N_15017,N_15282);
and U16620 (N_16620,N_15307,N_15954);
nor U16621 (N_16621,N_15979,N_15946);
or U16622 (N_16622,N_15314,N_15128);
nor U16623 (N_16623,N_15943,N_15394);
nand U16624 (N_16624,N_15406,N_15942);
nand U16625 (N_16625,N_15282,N_15238);
nor U16626 (N_16626,N_15396,N_15185);
nor U16627 (N_16627,N_15815,N_15258);
and U16628 (N_16628,N_15894,N_15287);
and U16629 (N_16629,N_15022,N_15592);
nor U16630 (N_16630,N_15554,N_15887);
or U16631 (N_16631,N_15997,N_15850);
xnor U16632 (N_16632,N_15214,N_15225);
xor U16633 (N_16633,N_15717,N_15394);
nand U16634 (N_16634,N_15591,N_15139);
nand U16635 (N_16635,N_15362,N_15063);
nor U16636 (N_16636,N_15259,N_15857);
xnor U16637 (N_16637,N_15985,N_15562);
or U16638 (N_16638,N_15509,N_15468);
nor U16639 (N_16639,N_15783,N_15707);
xnor U16640 (N_16640,N_15384,N_15461);
nand U16641 (N_16641,N_15758,N_15674);
or U16642 (N_16642,N_15948,N_15783);
nor U16643 (N_16643,N_15248,N_15386);
nor U16644 (N_16644,N_15969,N_15082);
nor U16645 (N_16645,N_15074,N_15643);
xnor U16646 (N_16646,N_15290,N_15753);
nor U16647 (N_16647,N_15072,N_15318);
nand U16648 (N_16648,N_15408,N_15595);
nor U16649 (N_16649,N_15191,N_15572);
and U16650 (N_16650,N_15630,N_15380);
and U16651 (N_16651,N_15579,N_15434);
nand U16652 (N_16652,N_15330,N_15834);
and U16653 (N_16653,N_15473,N_15202);
xor U16654 (N_16654,N_15084,N_15852);
nor U16655 (N_16655,N_15333,N_15391);
or U16656 (N_16656,N_15249,N_15225);
or U16657 (N_16657,N_15974,N_15773);
nand U16658 (N_16658,N_15609,N_15733);
xor U16659 (N_16659,N_15173,N_15352);
nor U16660 (N_16660,N_15881,N_15900);
or U16661 (N_16661,N_15489,N_15336);
nand U16662 (N_16662,N_15361,N_15287);
or U16663 (N_16663,N_15067,N_15299);
nor U16664 (N_16664,N_15306,N_15381);
and U16665 (N_16665,N_15989,N_15157);
xnor U16666 (N_16666,N_15303,N_15782);
and U16667 (N_16667,N_15187,N_15051);
and U16668 (N_16668,N_15216,N_15663);
or U16669 (N_16669,N_15858,N_15546);
or U16670 (N_16670,N_15117,N_15373);
and U16671 (N_16671,N_15798,N_15628);
nand U16672 (N_16672,N_15955,N_15054);
xor U16673 (N_16673,N_15644,N_15005);
and U16674 (N_16674,N_15066,N_15841);
nor U16675 (N_16675,N_15661,N_15942);
or U16676 (N_16676,N_15488,N_15376);
nand U16677 (N_16677,N_15308,N_15962);
or U16678 (N_16678,N_15825,N_15434);
and U16679 (N_16679,N_15831,N_15307);
nor U16680 (N_16680,N_15024,N_15507);
nor U16681 (N_16681,N_15957,N_15853);
or U16682 (N_16682,N_15822,N_15490);
nor U16683 (N_16683,N_15060,N_15277);
and U16684 (N_16684,N_15559,N_15476);
nand U16685 (N_16685,N_15016,N_15326);
xnor U16686 (N_16686,N_15671,N_15496);
or U16687 (N_16687,N_15952,N_15535);
or U16688 (N_16688,N_15832,N_15033);
or U16689 (N_16689,N_15343,N_15336);
or U16690 (N_16690,N_15064,N_15120);
xnor U16691 (N_16691,N_15846,N_15111);
nor U16692 (N_16692,N_15472,N_15199);
or U16693 (N_16693,N_15587,N_15599);
or U16694 (N_16694,N_15504,N_15220);
and U16695 (N_16695,N_15858,N_15169);
xor U16696 (N_16696,N_15599,N_15629);
and U16697 (N_16697,N_15053,N_15798);
nor U16698 (N_16698,N_15093,N_15722);
or U16699 (N_16699,N_15863,N_15330);
nor U16700 (N_16700,N_15837,N_15657);
or U16701 (N_16701,N_15391,N_15052);
nand U16702 (N_16702,N_15600,N_15757);
or U16703 (N_16703,N_15285,N_15745);
and U16704 (N_16704,N_15611,N_15867);
nand U16705 (N_16705,N_15266,N_15776);
and U16706 (N_16706,N_15306,N_15911);
nand U16707 (N_16707,N_15411,N_15087);
or U16708 (N_16708,N_15510,N_15668);
nor U16709 (N_16709,N_15168,N_15642);
nor U16710 (N_16710,N_15082,N_15004);
xnor U16711 (N_16711,N_15256,N_15425);
nand U16712 (N_16712,N_15829,N_15236);
or U16713 (N_16713,N_15335,N_15972);
xor U16714 (N_16714,N_15691,N_15268);
and U16715 (N_16715,N_15416,N_15224);
or U16716 (N_16716,N_15984,N_15409);
and U16717 (N_16717,N_15846,N_15026);
or U16718 (N_16718,N_15557,N_15816);
xor U16719 (N_16719,N_15717,N_15797);
xnor U16720 (N_16720,N_15843,N_15367);
xnor U16721 (N_16721,N_15848,N_15795);
nor U16722 (N_16722,N_15691,N_15153);
or U16723 (N_16723,N_15166,N_15953);
and U16724 (N_16724,N_15308,N_15205);
and U16725 (N_16725,N_15451,N_15702);
or U16726 (N_16726,N_15227,N_15990);
and U16727 (N_16727,N_15664,N_15652);
nand U16728 (N_16728,N_15198,N_15703);
nor U16729 (N_16729,N_15782,N_15291);
or U16730 (N_16730,N_15177,N_15836);
or U16731 (N_16731,N_15383,N_15603);
and U16732 (N_16732,N_15277,N_15037);
xnor U16733 (N_16733,N_15152,N_15797);
or U16734 (N_16734,N_15555,N_15433);
and U16735 (N_16735,N_15906,N_15588);
nand U16736 (N_16736,N_15234,N_15843);
nand U16737 (N_16737,N_15538,N_15854);
and U16738 (N_16738,N_15706,N_15387);
nor U16739 (N_16739,N_15480,N_15756);
nor U16740 (N_16740,N_15709,N_15012);
nor U16741 (N_16741,N_15421,N_15163);
nor U16742 (N_16742,N_15734,N_15096);
nor U16743 (N_16743,N_15375,N_15713);
xor U16744 (N_16744,N_15530,N_15997);
nand U16745 (N_16745,N_15855,N_15501);
and U16746 (N_16746,N_15605,N_15502);
and U16747 (N_16747,N_15517,N_15349);
nand U16748 (N_16748,N_15459,N_15176);
nand U16749 (N_16749,N_15798,N_15152);
xnor U16750 (N_16750,N_15910,N_15819);
and U16751 (N_16751,N_15331,N_15252);
xnor U16752 (N_16752,N_15775,N_15064);
nor U16753 (N_16753,N_15915,N_15272);
or U16754 (N_16754,N_15238,N_15017);
and U16755 (N_16755,N_15387,N_15898);
xor U16756 (N_16756,N_15397,N_15217);
nor U16757 (N_16757,N_15101,N_15429);
nand U16758 (N_16758,N_15506,N_15881);
and U16759 (N_16759,N_15710,N_15181);
nand U16760 (N_16760,N_15418,N_15790);
and U16761 (N_16761,N_15705,N_15678);
nor U16762 (N_16762,N_15840,N_15540);
or U16763 (N_16763,N_15133,N_15614);
or U16764 (N_16764,N_15185,N_15980);
xnor U16765 (N_16765,N_15447,N_15406);
or U16766 (N_16766,N_15653,N_15832);
and U16767 (N_16767,N_15148,N_15333);
nor U16768 (N_16768,N_15072,N_15181);
and U16769 (N_16769,N_15184,N_15701);
or U16770 (N_16770,N_15524,N_15935);
or U16771 (N_16771,N_15939,N_15371);
nand U16772 (N_16772,N_15162,N_15595);
nor U16773 (N_16773,N_15932,N_15127);
xnor U16774 (N_16774,N_15827,N_15182);
xnor U16775 (N_16775,N_15257,N_15168);
xnor U16776 (N_16776,N_15973,N_15528);
nor U16777 (N_16777,N_15666,N_15654);
or U16778 (N_16778,N_15608,N_15910);
xor U16779 (N_16779,N_15034,N_15246);
or U16780 (N_16780,N_15733,N_15664);
and U16781 (N_16781,N_15011,N_15841);
nor U16782 (N_16782,N_15880,N_15518);
and U16783 (N_16783,N_15484,N_15251);
nand U16784 (N_16784,N_15626,N_15294);
or U16785 (N_16785,N_15658,N_15362);
xnor U16786 (N_16786,N_15976,N_15153);
nor U16787 (N_16787,N_15494,N_15421);
and U16788 (N_16788,N_15374,N_15429);
or U16789 (N_16789,N_15603,N_15770);
xor U16790 (N_16790,N_15914,N_15679);
xnor U16791 (N_16791,N_15484,N_15475);
or U16792 (N_16792,N_15776,N_15367);
and U16793 (N_16793,N_15080,N_15848);
nand U16794 (N_16794,N_15091,N_15999);
nand U16795 (N_16795,N_15709,N_15886);
nand U16796 (N_16796,N_15870,N_15469);
nand U16797 (N_16797,N_15766,N_15365);
xor U16798 (N_16798,N_15409,N_15055);
nand U16799 (N_16799,N_15677,N_15070);
nor U16800 (N_16800,N_15534,N_15057);
or U16801 (N_16801,N_15058,N_15684);
or U16802 (N_16802,N_15305,N_15394);
or U16803 (N_16803,N_15607,N_15344);
nor U16804 (N_16804,N_15958,N_15821);
or U16805 (N_16805,N_15562,N_15377);
or U16806 (N_16806,N_15698,N_15162);
nand U16807 (N_16807,N_15717,N_15038);
and U16808 (N_16808,N_15586,N_15252);
and U16809 (N_16809,N_15997,N_15018);
or U16810 (N_16810,N_15057,N_15287);
xnor U16811 (N_16811,N_15947,N_15419);
and U16812 (N_16812,N_15847,N_15978);
and U16813 (N_16813,N_15729,N_15307);
or U16814 (N_16814,N_15217,N_15083);
xnor U16815 (N_16815,N_15227,N_15785);
xor U16816 (N_16816,N_15434,N_15215);
xor U16817 (N_16817,N_15076,N_15284);
nand U16818 (N_16818,N_15965,N_15801);
nand U16819 (N_16819,N_15943,N_15200);
or U16820 (N_16820,N_15516,N_15049);
and U16821 (N_16821,N_15198,N_15206);
nand U16822 (N_16822,N_15440,N_15246);
xor U16823 (N_16823,N_15678,N_15399);
nor U16824 (N_16824,N_15517,N_15999);
xnor U16825 (N_16825,N_15130,N_15277);
and U16826 (N_16826,N_15563,N_15290);
xnor U16827 (N_16827,N_15617,N_15432);
and U16828 (N_16828,N_15255,N_15958);
nand U16829 (N_16829,N_15026,N_15434);
nor U16830 (N_16830,N_15325,N_15911);
and U16831 (N_16831,N_15092,N_15973);
nand U16832 (N_16832,N_15659,N_15574);
and U16833 (N_16833,N_15402,N_15197);
or U16834 (N_16834,N_15293,N_15148);
nor U16835 (N_16835,N_15036,N_15058);
or U16836 (N_16836,N_15782,N_15978);
xnor U16837 (N_16837,N_15249,N_15174);
xnor U16838 (N_16838,N_15302,N_15586);
nor U16839 (N_16839,N_15747,N_15903);
xor U16840 (N_16840,N_15128,N_15191);
xnor U16841 (N_16841,N_15409,N_15062);
xnor U16842 (N_16842,N_15416,N_15132);
nor U16843 (N_16843,N_15465,N_15599);
nand U16844 (N_16844,N_15567,N_15030);
xor U16845 (N_16845,N_15507,N_15222);
or U16846 (N_16846,N_15053,N_15348);
nor U16847 (N_16847,N_15848,N_15997);
or U16848 (N_16848,N_15644,N_15331);
xor U16849 (N_16849,N_15484,N_15209);
xnor U16850 (N_16850,N_15635,N_15243);
and U16851 (N_16851,N_15912,N_15407);
and U16852 (N_16852,N_15003,N_15399);
or U16853 (N_16853,N_15675,N_15514);
and U16854 (N_16854,N_15474,N_15331);
xnor U16855 (N_16855,N_15401,N_15695);
or U16856 (N_16856,N_15653,N_15624);
nor U16857 (N_16857,N_15225,N_15546);
xnor U16858 (N_16858,N_15331,N_15919);
nor U16859 (N_16859,N_15863,N_15760);
or U16860 (N_16860,N_15325,N_15765);
xnor U16861 (N_16861,N_15866,N_15518);
xor U16862 (N_16862,N_15020,N_15615);
or U16863 (N_16863,N_15473,N_15454);
xnor U16864 (N_16864,N_15901,N_15076);
and U16865 (N_16865,N_15797,N_15366);
or U16866 (N_16866,N_15325,N_15860);
and U16867 (N_16867,N_15216,N_15430);
or U16868 (N_16868,N_15924,N_15277);
and U16869 (N_16869,N_15292,N_15706);
nand U16870 (N_16870,N_15757,N_15255);
and U16871 (N_16871,N_15770,N_15180);
xor U16872 (N_16872,N_15085,N_15665);
xor U16873 (N_16873,N_15017,N_15184);
xnor U16874 (N_16874,N_15624,N_15672);
nand U16875 (N_16875,N_15125,N_15931);
nor U16876 (N_16876,N_15555,N_15564);
and U16877 (N_16877,N_15721,N_15771);
nor U16878 (N_16878,N_15902,N_15910);
nand U16879 (N_16879,N_15225,N_15375);
and U16880 (N_16880,N_15273,N_15234);
nand U16881 (N_16881,N_15162,N_15192);
or U16882 (N_16882,N_15700,N_15799);
xor U16883 (N_16883,N_15205,N_15021);
xor U16884 (N_16884,N_15181,N_15117);
nor U16885 (N_16885,N_15098,N_15865);
nor U16886 (N_16886,N_15144,N_15442);
nand U16887 (N_16887,N_15475,N_15848);
and U16888 (N_16888,N_15346,N_15090);
xor U16889 (N_16889,N_15728,N_15749);
nor U16890 (N_16890,N_15644,N_15627);
nor U16891 (N_16891,N_15579,N_15125);
xnor U16892 (N_16892,N_15907,N_15931);
or U16893 (N_16893,N_15832,N_15996);
nand U16894 (N_16894,N_15736,N_15224);
or U16895 (N_16895,N_15076,N_15170);
or U16896 (N_16896,N_15596,N_15792);
or U16897 (N_16897,N_15631,N_15460);
xor U16898 (N_16898,N_15383,N_15040);
and U16899 (N_16899,N_15137,N_15356);
or U16900 (N_16900,N_15943,N_15492);
xnor U16901 (N_16901,N_15556,N_15588);
and U16902 (N_16902,N_15422,N_15712);
xor U16903 (N_16903,N_15738,N_15361);
xor U16904 (N_16904,N_15734,N_15538);
and U16905 (N_16905,N_15813,N_15269);
xor U16906 (N_16906,N_15107,N_15563);
xnor U16907 (N_16907,N_15683,N_15717);
and U16908 (N_16908,N_15352,N_15533);
xor U16909 (N_16909,N_15637,N_15736);
and U16910 (N_16910,N_15704,N_15505);
xor U16911 (N_16911,N_15098,N_15353);
or U16912 (N_16912,N_15959,N_15703);
xor U16913 (N_16913,N_15158,N_15834);
nand U16914 (N_16914,N_15962,N_15737);
nor U16915 (N_16915,N_15056,N_15370);
and U16916 (N_16916,N_15538,N_15524);
or U16917 (N_16917,N_15641,N_15428);
xnor U16918 (N_16918,N_15210,N_15312);
or U16919 (N_16919,N_15024,N_15796);
xnor U16920 (N_16920,N_15127,N_15353);
nand U16921 (N_16921,N_15899,N_15667);
or U16922 (N_16922,N_15945,N_15025);
nor U16923 (N_16923,N_15994,N_15792);
xor U16924 (N_16924,N_15869,N_15504);
and U16925 (N_16925,N_15783,N_15202);
nor U16926 (N_16926,N_15208,N_15000);
or U16927 (N_16927,N_15835,N_15418);
nor U16928 (N_16928,N_15810,N_15297);
nor U16929 (N_16929,N_15215,N_15611);
nand U16930 (N_16930,N_15908,N_15548);
xor U16931 (N_16931,N_15414,N_15829);
nand U16932 (N_16932,N_15525,N_15435);
nor U16933 (N_16933,N_15080,N_15662);
xnor U16934 (N_16934,N_15731,N_15381);
nor U16935 (N_16935,N_15094,N_15821);
xnor U16936 (N_16936,N_15245,N_15637);
xor U16937 (N_16937,N_15060,N_15079);
or U16938 (N_16938,N_15834,N_15729);
and U16939 (N_16939,N_15682,N_15624);
and U16940 (N_16940,N_15930,N_15622);
nand U16941 (N_16941,N_15992,N_15078);
xnor U16942 (N_16942,N_15848,N_15455);
nand U16943 (N_16943,N_15519,N_15020);
xor U16944 (N_16944,N_15239,N_15887);
and U16945 (N_16945,N_15790,N_15369);
or U16946 (N_16946,N_15784,N_15086);
nand U16947 (N_16947,N_15729,N_15862);
and U16948 (N_16948,N_15312,N_15371);
xor U16949 (N_16949,N_15732,N_15240);
nand U16950 (N_16950,N_15514,N_15029);
or U16951 (N_16951,N_15499,N_15067);
or U16952 (N_16952,N_15022,N_15452);
or U16953 (N_16953,N_15524,N_15795);
nand U16954 (N_16954,N_15180,N_15134);
xnor U16955 (N_16955,N_15747,N_15929);
or U16956 (N_16956,N_15605,N_15479);
and U16957 (N_16957,N_15481,N_15416);
and U16958 (N_16958,N_15924,N_15545);
nand U16959 (N_16959,N_15659,N_15503);
and U16960 (N_16960,N_15018,N_15070);
or U16961 (N_16961,N_15803,N_15020);
and U16962 (N_16962,N_15714,N_15587);
xnor U16963 (N_16963,N_15950,N_15847);
or U16964 (N_16964,N_15473,N_15282);
nand U16965 (N_16965,N_15996,N_15525);
xnor U16966 (N_16966,N_15528,N_15844);
and U16967 (N_16967,N_15032,N_15283);
or U16968 (N_16968,N_15152,N_15836);
nor U16969 (N_16969,N_15511,N_15575);
nand U16970 (N_16970,N_15470,N_15610);
and U16971 (N_16971,N_15693,N_15258);
and U16972 (N_16972,N_15137,N_15200);
nor U16973 (N_16973,N_15290,N_15787);
or U16974 (N_16974,N_15567,N_15225);
nand U16975 (N_16975,N_15262,N_15968);
nor U16976 (N_16976,N_15991,N_15547);
or U16977 (N_16977,N_15119,N_15701);
nor U16978 (N_16978,N_15775,N_15765);
xor U16979 (N_16979,N_15550,N_15142);
nand U16980 (N_16980,N_15996,N_15726);
nor U16981 (N_16981,N_15338,N_15928);
nand U16982 (N_16982,N_15470,N_15607);
or U16983 (N_16983,N_15825,N_15012);
nand U16984 (N_16984,N_15849,N_15537);
nand U16985 (N_16985,N_15948,N_15452);
nand U16986 (N_16986,N_15778,N_15945);
and U16987 (N_16987,N_15359,N_15842);
nand U16988 (N_16988,N_15013,N_15029);
and U16989 (N_16989,N_15193,N_15320);
xor U16990 (N_16990,N_15058,N_15982);
xnor U16991 (N_16991,N_15252,N_15651);
xnor U16992 (N_16992,N_15267,N_15386);
and U16993 (N_16993,N_15052,N_15420);
and U16994 (N_16994,N_15999,N_15031);
nor U16995 (N_16995,N_15645,N_15854);
nand U16996 (N_16996,N_15084,N_15167);
and U16997 (N_16997,N_15937,N_15494);
nand U16998 (N_16998,N_15128,N_15343);
nor U16999 (N_16999,N_15541,N_15574);
xnor U17000 (N_17000,N_16920,N_16417);
xor U17001 (N_17001,N_16473,N_16895);
and U17002 (N_17002,N_16192,N_16114);
and U17003 (N_17003,N_16581,N_16050);
or U17004 (N_17004,N_16888,N_16152);
nor U17005 (N_17005,N_16383,N_16018);
and U17006 (N_17006,N_16489,N_16721);
and U17007 (N_17007,N_16154,N_16767);
xnor U17008 (N_17008,N_16651,N_16816);
xor U17009 (N_17009,N_16412,N_16270);
and U17010 (N_17010,N_16731,N_16670);
or U17011 (N_17011,N_16458,N_16355);
nor U17012 (N_17012,N_16541,N_16961);
or U17013 (N_17013,N_16750,N_16409);
or U17014 (N_17014,N_16638,N_16413);
and U17015 (N_17015,N_16785,N_16981);
nand U17016 (N_17016,N_16705,N_16525);
xnor U17017 (N_17017,N_16683,N_16499);
nor U17018 (N_17018,N_16319,N_16389);
nor U17019 (N_17019,N_16827,N_16034);
and U17020 (N_17020,N_16505,N_16357);
or U17021 (N_17021,N_16977,N_16886);
nand U17022 (N_17022,N_16483,N_16302);
nand U17023 (N_17023,N_16215,N_16928);
or U17024 (N_17024,N_16301,N_16444);
nor U17025 (N_17025,N_16599,N_16277);
nor U17026 (N_17026,N_16733,N_16632);
xnor U17027 (N_17027,N_16693,N_16808);
or U17028 (N_17028,N_16916,N_16479);
xor U17029 (N_17029,N_16268,N_16054);
or U17030 (N_17030,N_16751,N_16374);
or U17031 (N_17031,N_16972,N_16157);
xnor U17032 (N_17032,N_16156,N_16713);
and U17033 (N_17033,N_16452,N_16254);
xnor U17034 (N_17034,N_16144,N_16300);
or U17035 (N_17035,N_16818,N_16789);
or U17036 (N_17036,N_16837,N_16992);
or U17037 (N_17037,N_16607,N_16967);
or U17038 (N_17038,N_16704,N_16520);
nor U17039 (N_17039,N_16351,N_16968);
xor U17040 (N_17040,N_16454,N_16059);
nand U17041 (N_17041,N_16791,N_16347);
or U17042 (N_17042,N_16365,N_16882);
or U17043 (N_17043,N_16832,N_16681);
and U17044 (N_17044,N_16463,N_16392);
nand U17045 (N_17045,N_16080,N_16876);
nand U17046 (N_17046,N_16949,N_16570);
nor U17047 (N_17047,N_16899,N_16074);
and U17048 (N_17048,N_16963,N_16273);
xor U17049 (N_17049,N_16769,N_16376);
and U17050 (N_17050,N_16013,N_16253);
xnor U17051 (N_17051,N_16232,N_16137);
nor U17052 (N_17052,N_16561,N_16123);
and U17053 (N_17053,N_16461,N_16535);
or U17054 (N_17054,N_16323,N_16439);
nor U17055 (N_17055,N_16699,N_16025);
nand U17056 (N_17056,N_16709,N_16290);
or U17057 (N_17057,N_16288,N_16994);
nor U17058 (N_17058,N_16507,N_16143);
xor U17059 (N_17059,N_16966,N_16904);
and U17060 (N_17060,N_16142,N_16622);
nand U17061 (N_17061,N_16258,N_16026);
nand U17062 (N_17062,N_16732,N_16038);
xnor U17063 (N_17063,N_16612,N_16056);
nor U17064 (N_17064,N_16041,N_16504);
nand U17065 (N_17065,N_16222,N_16325);
nand U17066 (N_17066,N_16665,N_16883);
nor U17067 (N_17067,N_16000,N_16740);
or U17068 (N_17068,N_16574,N_16345);
nand U17069 (N_17069,N_16506,N_16102);
nand U17070 (N_17070,N_16335,N_16197);
or U17071 (N_17071,N_16231,N_16261);
or U17072 (N_17072,N_16905,N_16094);
or U17073 (N_17073,N_16488,N_16692);
nand U17074 (N_17074,N_16498,N_16263);
nor U17075 (N_17075,N_16195,N_16427);
nor U17076 (N_17076,N_16328,N_16324);
nor U17077 (N_17077,N_16341,N_16546);
nor U17078 (N_17078,N_16297,N_16111);
nor U17079 (N_17079,N_16957,N_16189);
nor U17080 (N_17080,N_16687,N_16202);
or U17081 (N_17081,N_16631,N_16039);
nand U17082 (N_17082,N_16012,N_16729);
xnor U17083 (N_17083,N_16861,N_16438);
or U17084 (N_17084,N_16746,N_16595);
nand U17085 (N_17085,N_16271,N_16233);
or U17086 (N_17086,N_16066,N_16022);
nor U17087 (N_17087,N_16199,N_16153);
nor U17088 (N_17088,N_16077,N_16947);
nand U17089 (N_17089,N_16698,N_16909);
and U17090 (N_17090,N_16216,N_16738);
xor U17091 (N_17091,N_16163,N_16696);
or U17092 (N_17092,N_16885,N_16623);
or U17093 (N_17093,N_16453,N_16762);
xnor U17094 (N_17094,N_16592,N_16641);
nand U17095 (N_17095,N_16255,N_16926);
or U17096 (N_17096,N_16008,N_16796);
xnor U17097 (N_17097,N_16027,N_16247);
nand U17098 (N_17098,N_16795,N_16941);
xor U17099 (N_17099,N_16537,N_16509);
xor U17100 (N_17100,N_16098,N_16471);
or U17101 (N_17101,N_16823,N_16423);
nor U17102 (N_17102,N_16933,N_16196);
and U17103 (N_17103,N_16125,N_16459);
nand U17104 (N_17104,N_16147,N_16118);
and U17105 (N_17105,N_16955,N_16431);
and U17106 (N_17106,N_16490,N_16180);
and U17107 (N_17107,N_16363,N_16855);
nand U17108 (N_17108,N_16893,N_16539);
nand U17109 (N_17109,N_16661,N_16478);
or U17110 (N_17110,N_16573,N_16062);
and U17111 (N_17111,N_16727,N_16419);
xnor U17112 (N_17112,N_16106,N_16690);
or U17113 (N_17113,N_16706,N_16274);
nor U17114 (N_17114,N_16129,N_16210);
nand U17115 (N_17115,N_16645,N_16282);
xnor U17116 (N_17116,N_16853,N_16628);
xnor U17117 (N_17117,N_16624,N_16408);
and U17118 (N_17118,N_16993,N_16446);
and U17119 (N_17119,N_16101,N_16029);
or U17120 (N_17120,N_16204,N_16477);
xnor U17121 (N_17121,N_16605,N_16394);
nand U17122 (N_17122,N_16646,N_16804);
or U17123 (N_17123,N_16894,N_16113);
and U17124 (N_17124,N_16810,N_16487);
nor U17125 (N_17125,N_16971,N_16688);
nor U17126 (N_17126,N_16549,N_16425);
nand U17127 (N_17127,N_16401,N_16572);
nor U17128 (N_17128,N_16346,N_16782);
nor U17129 (N_17129,N_16332,N_16133);
or U17130 (N_17130,N_16203,N_16829);
xor U17131 (N_17131,N_16072,N_16711);
and U17132 (N_17132,N_16975,N_16462);
or U17133 (N_17133,N_16672,N_16794);
xor U17134 (N_17134,N_16863,N_16435);
and U17135 (N_17135,N_16639,N_16495);
nand U17136 (N_17136,N_16226,N_16768);
and U17137 (N_17137,N_16787,N_16220);
nor U17138 (N_17138,N_16533,N_16775);
and U17139 (N_17139,N_16521,N_16660);
nand U17140 (N_17140,N_16181,N_16119);
nand U17141 (N_17141,N_16779,N_16173);
xnor U17142 (N_17142,N_16754,N_16650);
and U17143 (N_17143,N_16763,N_16124);
nand U17144 (N_17144,N_16793,N_16151);
or U17145 (N_17145,N_16707,N_16719);
and U17146 (N_17146,N_16964,N_16090);
xnor U17147 (N_17147,N_16285,N_16177);
nand U17148 (N_17148,N_16148,N_16329);
and U17149 (N_17149,N_16900,N_16340);
or U17150 (N_17150,N_16836,N_16988);
nor U17151 (N_17151,N_16860,N_16006);
and U17152 (N_17152,N_16428,N_16393);
and U17153 (N_17153,N_16112,N_16318);
and U17154 (N_17154,N_16141,N_16064);
and U17155 (N_17155,N_16480,N_16896);
or U17156 (N_17156,N_16398,N_16887);
and U17157 (N_17157,N_16803,N_16245);
nand U17158 (N_17158,N_16482,N_16206);
and U17159 (N_17159,N_16099,N_16815);
and U17160 (N_17160,N_16635,N_16958);
nand U17161 (N_17161,N_16223,N_16771);
xnor U17162 (N_17162,N_16096,N_16241);
or U17163 (N_17163,N_16500,N_16697);
and U17164 (N_17164,N_16606,N_16566);
nand U17165 (N_17165,N_16501,N_16472);
or U17166 (N_17166,N_16049,N_16040);
nor U17167 (N_17167,N_16044,N_16333);
nand U17168 (N_17168,N_16484,N_16674);
and U17169 (N_17169,N_16185,N_16221);
nand U17170 (N_17170,N_16265,N_16726);
and U17171 (N_17171,N_16184,N_16551);
or U17172 (N_17172,N_16851,N_16209);
nand U17173 (N_17173,N_16880,N_16822);
nand U17174 (N_17174,N_16280,N_16790);
or U17175 (N_17175,N_16873,N_16716);
xnor U17176 (N_17176,N_16379,N_16582);
nand U17177 (N_17177,N_16370,N_16455);
xnor U17178 (N_17178,N_16912,N_16310);
xnor U17179 (N_17179,N_16309,N_16655);
nor U17180 (N_17180,N_16432,N_16999);
and U17181 (N_17181,N_16200,N_16492);
or U17182 (N_17182,N_16313,N_16685);
or U17183 (N_17183,N_16361,N_16814);
or U17184 (N_17184,N_16294,N_16243);
and U17185 (N_17185,N_16367,N_16373);
nor U17186 (N_17186,N_16805,N_16677);
xor U17187 (N_17187,N_16009,N_16456);
and U17188 (N_17188,N_16703,N_16083);
xor U17189 (N_17189,N_16710,N_16756);
xor U17190 (N_17190,N_16925,N_16475);
and U17191 (N_17191,N_16491,N_16035);
nand U17192 (N_17192,N_16128,N_16673);
nand U17193 (N_17193,N_16517,N_16591);
nor U17194 (N_17194,N_16812,N_16036);
nand U17195 (N_17195,N_16922,N_16449);
nor U17196 (N_17196,N_16919,N_16293);
xnor U17197 (N_17197,N_16684,N_16720);
nor U17198 (N_17198,N_16846,N_16296);
xnor U17199 (N_17199,N_16217,N_16061);
xnor U17200 (N_17200,N_16979,N_16973);
xor U17201 (N_17201,N_16403,N_16969);
or U17202 (N_17202,N_16366,N_16020);
nand U17203 (N_17203,N_16053,N_16135);
and U17204 (N_17204,N_16918,N_16776);
nor U17205 (N_17205,N_16227,N_16902);
xor U17206 (N_17206,N_16759,N_16554);
and U17207 (N_17207,N_16126,N_16602);
and U17208 (N_17208,N_16436,N_16700);
nor U17209 (N_17209,N_16819,N_16802);
and U17210 (N_17210,N_16372,N_16866);
nor U17211 (N_17211,N_16278,N_16652);
or U17212 (N_17212,N_16609,N_16086);
nor U17213 (N_17213,N_16773,N_16741);
or U17214 (N_17214,N_16884,N_16758);
or U17215 (N_17215,N_16865,N_16174);
xnor U17216 (N_17216,N_16249,N_16275);
nand U17217 (N_17217,N_16630,N_16780);
nor U17218 (N_17218,N_16625,N_16619);
and U17219 (N_17219,N_16312,N_16248);
nor U17220 (N_17220,N_16381,N_16970);
xor U17221 (N_17221,N_16854,N_16171);
or U17222 (N_17222,N_16159,N_16161);
or U17223 (N_17223,N_16985,N_16214);
and U17224 (N_17224,N_16644,N_16911);
xnor U17225 (N_17225,N_16033,N_16877);
nand U17226 (N_17226,N_16559,N_16081);
xor U17227 (N_17227,N_16236,N_16540);
and U17228 (N_17228,N_16138,N_16809);
xor U17229 (N_17229,N_16104,N_16131);
and U17230 (N_17230,N_16228,N_16532);
xor U17231 (N_17231,N_16600,N_16075);
or U17232 (N_17232,N_16406,N_16330);
and U17233 (N_17233,N_16264,N_16543);
and U17234 (N_17234,N_16092,N_16334);
or U17235 (N_17235,N_16512,N_16991);
xnor U17236 (N_17236,N_16469,N_16648);
xnor U17237 (N_17237,N_16617,N_16744);
and U17238 (N_17238,N_16781,N_16434);
nor U17239 (N_17239,N_16353,N_16830);
xor U17240 (N_17240,N_16534,N_16753);
nor U17241 (N_17241,N_16465,N_16736);
nor U17242 (N_17242,N_16752,N_16948);
xor U17243 (N_17243,N_16160,N_16115);
xnor U17244 (N_17244,N_16003,N_16872);
or U17245 (N_17245,N_16359,N_16045);
or U17246 (N_17246,N_16450,N_16842);
xnor U17247 (N_17247,N_16337,N_16915);
nand U17248 (N_17248,N_16945,N_16664);
and U17249 (N_17249,N_16548,N_16695);
nor U17250 (N_17250,N_16354,N_16242);
and U17251 (N_17251,N_16874,N_16564);
or U17252 (N_17252,N_16005,N_16611);
nand U17253 (N_17253,N_16272,N_16134);
or U17254 (N_17254,N_16065,N_16937);
or U17255 (N_17255,N_16585,N_16850);
or U17256 (N_17256,N_16516,N_16722);
and U17257 (N_17257,N_16338,N_16420);
xor U17258 (N_17258,N_16244,N_16058);
nor U17259 (N_17259,N_16468,N_16680);
and U17260 (N_17260,N_16658,N_16788);
or U17261 (N_17261,N_16327,N_16042);
and U17262 (N_17262,N_16402,N_16682);
nor U17263 (N_17263,N_16982,N_16828);
nor U17264 (N_17264,N_16765,N_16730);
nor U17265 (N_17265,N_16831,N_16158);
nand U17266 (N_17266,N_16834,N_16870);
xnor U17267 (N_17267,N_16932,N_16095);
xnor U17268 (N_17268,N_16170,N_16770);
nor U17269 (N_17269,N_16636,N_16100);
and U17270 (N_17270,N_16878,N_16063);
and U17271 (N_17271,N_16194,N_16057);
or U17272 (N_17272,N_16046,N_16524);
and U17273 (N_17273,N_16784,N_16028);
nor U17274 (N_17274,N_16513,N_16048);
and U17275 (N_17275,N_16859,N_16717);
and U17276 (N_17276,N_16108,N_16826);
and U17277 (N_17277,N_16946,N_16596);
nand U17278 (N_17278,N_16120,N_16117);
or U17279 (N_17279,N_16457,N_16956);
or U17280 (N_17280,N_16903,N_16542);
nor U17281 (N_17281,N_16983,N_16901);
and U17282 (N_17282,N_16508,N_16924);
or U17283 (N_17283,N_16464,N_16519);
nand U17284 (N_17284,N_16890,N_16481);
or U17285 (N_17285,N_16089,N_16728);
nand U17286 (N_17286,N_16702,N_16503);
xnor U17287 (N_17287,N_16176,N_16360);
nor U17288 (N_17288,N_16974,N_16939);
nand U17289 (N_17289,N_16127,N_16284);
or U17290 (N_17290,N_16266,N_16349);
or U17291 (N_17291,N_16545,N_16218);
nor U17292 (N_17292,N_16667,N_16875);
xnor U17293 (N_17293,N_16743,N_16016);
or U17294 (N_17294,N_16356,N_16962);
nor U17295 (N_17295,N_16289,N_16544);
or U17296 (N_17296,N_16835,N_16640);
nor U17297 (N_17297,N_16723,N_16526);
nor U17298 (N_17298,N_16030,N_16906);
nor U17299 (N_17299,N_16426,N_16856);
and U17300 (N_17300,N_16257,N_16399);
nor U17301 (N_17301,N_16868,N_16165);
and U17302 (N_17302,N_16011,N_16343);
or U17303 (N_17303,N_16306,N_16430);
xor U17304 (N_17304,N_16493,N_16388);
or U17305 (N_17305,N_16068,N_16342);
nor U17306 (N_17306,N_16441,N_16317);
nand U17307 (N_17307,N_16395,N_16824);
nor U17308 (N_17308,N_16734,N_16188);
nor U17309 (N_17309,N_16350,N_16445);
or U17310 (N_17310,N_16862,N_16755);
xnor U17311 (N_17311,N_16421,N_16528);
or U17312 (N_17312,N_16183,N_16443);
nor U17313 (N_17313,N_16604,N_16518);
xnor U17314 (N_17314,N_16642,N_16764);
or U17315 (N_17315,N_16691,N_16577);
nand U17316 (N_17316,N_16397,N_16817);
nor U17317 (N_17317,N_16110,N_16286);
xnor U17318 (N_17318,N_16097,N_16198);
xnor U17319 (N_17319,N_16840,N_16140);
nand U17320 (N_17320,N_16400,N_16671);
nand U17321 (N_17321,N_16766,N_16010);
nor U17322 (N_17322,N_16615,N_16621);
nand U17323 (N_17323,N_16538,N_16881);
and U17324 (N_17324,N_16073,N_16235);
nor U17325 (N_17325,N_16792,N_16213);
nor U17326 (N_17326,N_16105,N_16742);
and U17327 (N_17327,N_16514,N_16485);
xnor U17328 (N_17328,N_16580,N_16307);
nand U17329 (N_17329,N_16201,N_16547);
nor U17330 (N_17330,N_16869,N_16069);
nand U17331 (N_17331,N_16989,N_16178);
nor U17332 (N_17332,N_16410,N_16908);
nor U17333 (N_17333,N_16339,N_16004);
nor U17334 (N_17334,N_16418,N_16404);
nor U17335 (N_17335,N_16515,N_16735);
and U17336 (N_17336,N_16291,N_16942);
nand U17337 (N_17337,N_16712,N_16078);
nor U17338 (N_17338,N_16191,N_16230);
xor U17339 (N_17339,N_16407,N_16913);
nand U17340 (N_17340,N_16259,N_16587);
nand U17341 (N_17341,N_16193,N_16739);
and U17342 (N_17342,N_16984,N_16914);
nor U17343 (N_17343,N_16643,N_16603);
nor U17344 (N_17344,N_16067,N_16558);
or U17345 (N_17345,N_16369,N_16447);
or U17346 (N_17346,N_16001,N_16806);
nor U17347 (N_17347,N_16364,N_16087);
nand U17348 (N_17348,N_16088,N_16380);
nand U17349 (N_17349,N_16694,N_16757);
nand U17350 (N_17350,N_16299,N_16557);
xnor U17351 (N_17351,N_16954,N_16959);
xor U17352 (N_17352,N_16237,N_16567);
xor U17353 (N_17353,N_16169,N_16225);
or U17354 (N_17354,N_16208,N_16637);
xor U17355 (N_17355,N_16931,N_16760);
nor U17356 (N_17356,N_16336,N_16470);
nor U17357 (N_17357,N_16749,N_16150);
or U17358 (N_17358,N_16960,N_16536);
xnor U17359 (N_17359,N_16283,N_16139);
or U17360 (N_17360,N_16416,N_16879);
nand U17361 (N_17361,N_16250,N_16316);
nor U17362 (N_17362,N_16082,N_16952);
nand U17363 (N_17363,N_16207,N_16889);
and U17364 (N_17364,N_16032,N_16167);
xnor U17365 (N_17365,N_16980,N_16303);
xor U17366 (N_17366,N_16689,N_16060);
and U17367 (N_17367,N_16362,N_16186);
nor U17368 (N_17368,N_16205,N_16633);
and U17369 (N_17369,N_16563,N_16593);
xnor U17370 (N_17370,N_16070,N_16023);
or U17371 (N_17371,N_16936,N_16718);
or U17372 (N_17372,N_16523,N_16530);
nor U17373 (N_17373,N_16986,N_16616);
nand U17374 (N_17374,N_16556,N_16320);
nor U17375 (N_17375,N_16260,N_16358);
nand U17376 (N_17376,N_16262,N_16848);
or U17377 (N_17377,N_16051,N_16579);
nor U17378 (N_17378,N_16076,N_16584);
nand U17379 (N_17379,N_16190,N_16411);
xnor U17380 (N_17380,N_16385,N_16384);
or U17381 (N_17381,N_16164,N_16747);
and U17382 (N_17382,N_16852,N_16943);
xnor U17383 (N_17383,N_16396,N_16725);
nor U17384 (N_17384,N_16838,N_16352);
or U17385 (N_17385,N_16898,N_16774);
nor U17386 (N_17386,N_16929,N_16252);
nor U17387 (N_17387,N_16847,N_16552);
nor U17388 (N_17388,N_16440,N_16414);
nand U17389 (N_17389,N_16390,N_16653);
or U17390 (N_17390,N_16675,N_16825);
or U17391 (N_17391,N_16976,N_16149);
nor U17392 (N_17392,N_16091,N_16575);
nand U17393 (N_17393,N_16162,N_16897);
and U17394 (N_17394,N_16304,N_16405);
nor U17395 (N_17395,N_16923,N_16620);
nor U17396 (N_17396,N_16024,N_16251);
nor U17397 (N_17397,N_16748,N_16571);
nand U17398 (N_17398,N_16424,N_16256);
or U17399 (N_17399,N_16927,N_16797);
xor U17400 (N_17400,N_16071,N_16669);
or U17401 (N_17401,N_16368,N_16531);
xnor U17402 (N_17402,N_16590,N_16839);
nor U17403 (N_17403,N_16807,N_16269);
and U17404 (N_17404,N_16662,N_16305);
nand U17405 (N_17405,N_16627,N_16281);
nor U17406 (N_17406,N_16820,N_16562);
nand U17407 (N_17407,N_16476,N_16344);
or U17408 (N_17408,N_16182,N_16084);
or U17409 (N_17409,N_16626,N_16331);
nand U17410 (N_17410,N_16858,N_16511);
xor U17411 (N_17411,N_16422,N_16657);
nand U17412 (N_17412,N_16234,N_16801);
nor U17413 (N_17413,N_16052,N_16938);
nor U17414 (N_17414,N_16017,N_16429);
xor U17415 (N_17415,N_16917,N_16569);
and U17416 (N_17416,N_16921,N_16867);
nor U17417 (N_17417,N_16085,N_16668);
xor U17418 (N_17418,N_16550,N_16935);
nor U17419 (N_17419,N_16136,N_16864);
nand U17420 (N_17420,N_16950,N_16654);
nand U17421 (N_17421,N_16841,N_16116);
nor U17422 (N_17422,N_16019,N_16745);
or U17423 (N_17423,N_16951,N_16714);
or U17424 (N_17424,N_16460,N_16871);
nor U17425 (N_17425,N_16560,N_16497);
nor U17426 (N_17426,N_16578,N_16415);
and U17427 (N_17427,N_16634,N_16267);
nand U17428 (N_17428,N_16629,N_16772);
or U17429 (N_17429,N_16348,N_16529);
nor U17430 (N_17430,N_16486,N_16555);
nor U17431 (N_17431,N_16015,N_16391);
or U17432 (N_17432,N_16647,N_16649);
or U17433 (N_17433,N_16998,N_16907);
nor U17434 (N_17434,N_16821,N_16813);
or U17435 (N_17435,N_16322,N_16007);
or U17436 (N_17436,N_16679,N_16522);
nand U17437 (N_17437,N_16002,N_16576);
or U17438 (N_17438,N_16502,N_16308);
xnor U17439 (N_17439,N_16783,N_16047);
nor U17440 (N_17440,N_16996,N_16724);
nor U17441 (N_17441,N_16833,N_16786);
or U17442 (N_17442,N_16168,N_16777);
nor U17443 (N_17443,N_16845,N_16997);
nand U17444 (N_17444,N_16451,N_16568);
xnor U17445 (N_17445,N_16103,N_16212);
or U17446 (N_17446,N_16844,N_16586);
nand U17447 (N_17447,N_16279,N_16708);
xnor U17448 (N_17448,N_16892,N_16211);
nor U17449 (N_17449,N_16145,N_16597);
nand U17450 (N_17450,N_16246,N_16676);
nor U17451 (N_17451,N_16467,N_16565);
nor U17452 (N_17452,N_16598,N_16109);
or U17453 (N_17453,N_16678,N_16799);
nand U17454 (N_17454,N_16953,N_16701);
xnor U17455 (N_17455,N_16442,N_16055);
or U17456 (N_17456,N_16166,N_16666);
and U17457 (N_17457,N_16849,N_16371);
and U17458 (N_17458,N_16295,N_16934);
xor U17459 (N_17459,N_16663,N_16172);
xor U17460 (N_17460,N_16229,N_16494);
and U17461 (N_17461,N_16239,N_16978);
nor U17462 (N_17462,N_16686,N_16079);
and U17463 (N_17463,N_16287,N_16107);
xor U17464 (N_17464,N_16179,N_16737);
and U17465 (N_17465,N_16122,N_16843);
xnor U17466 (N_17466,N_16175,N_16659);
nand U17467 (N_17467,N_16311,N_16037);
xor U17468 (N_17468,N_16146,N_16608);
xnor U17469 (N_17469,N_16382,N_16326);
nand U17470 (N_17470,N_16588,N_16377);
nand U17471 (N_17471,N_16474,N_16910);
or U17472 (N_17472,N_16130,N_16386);
and U17473 (N_17473,N_16238,N_16601);
and U17474 (N_17474,N_16553,N_16132);
xor U17475 (N_17475,N_16155,N_16292);
xor U17476 (N_17476,N_16656,N_16298);
and U17477 (N_17477,N_16995,N_16121);
or U17478 (N_17478,N_16448,N_16021);
xor U17479 (N_17479,N_16496,N_16891);
and U17480 (N_17480,N_16583,N_16987);
and U17481 (N_17481,N_16466,N_16375);
nand U17482 (N_17482,N_16761,N_16594);
or U17483 (N_17483,N_16314,N_16930);
nand U17484 (N_17484,N_16800,N_16315);
and U17485 (N_17485,N_16940,N_16527);
nand U17486 (N_17486,N_16857,N_16321);
nor U17487 (N_17487,N_16387,N_16014);
and U17488 (N_17488,N_16187,N_16798);
xor U17489 (N_17489,N_16589,N_16093);
or U17490 (N_17490,N_16811,N_16614);
and U17491 (N_17491,N_16043,N_16031);
or U17492 (N_17492,N_16219,N_16944);
nor U17493 (N_17493,N_16618,N_16276);
nor U17494 (N_17494,N_16990,N_16224);
or U17495 (N_17495,N_16378,N_16240);
nor U17496 (N_17496,N_16433,N_16610);
and U17497 (N_17497,N_16510,N_16778);
or U17498 (N_17498,N_16613,N_16715);
nor U17499 (N_17499,N_16965,N_16437);
nand U17500 (N_17500,N_16083,N_16007);
or U17501 (N_17501,N_16290,N_16278);
and U17502 (N_17502,N_16796,N_16914);
and U17503 (N_17503,N_16596,N_16050);
and U17504 (N_17504,N_16873,N_16856);
nor U17505 (N_17505,N_16012,N_16604);
or U17506 (N_17506,N_16436,N_16083);
nor U17507 (N_17507,N_16579,N_16455);
nor U17508 (N_17508,N_16229,N_16320);
nand U17509 (N_17509,N_16694,N_16364);
xor U17510 (N_17510,N_16434,N_16881);
xnor U17511 (N_17511,N_16779,N_16388);
nor U17512 (N_17512,N_16298,N_16282);
and U17513 (N_17513,N_16616,N_16507);
and U17514 (N_17514,N_16086,N_16706);
and U17515 (N_17515,N_16680,N_16376);
and U17516 (N_17516,N_16242,N_16741);
and U17517 (N_17517,N_16619,N_16848);
nor U17518 (N_17518,N_16254,N_16167);
nand U17519 (N_17519,N_16978,N_16564);
nor U17520 (N_17520,N_16397,N_16237);
nor U17521 (N_17521,N_16203,N_16564);
and U17522 (N_17522,N_16030,N_16000);
nand U17523 (N_17523,N_16165,N_16860);
nand U17524 (N_17524,N_16583,N_16339);
nand U17525 (N_17525,N_16572,N_16992);
nand U17526 (N_17526,N_16859,N_16371);
xor U17527 (N_17527,N_16772,N_16590);
nor U17528 (N_17528,N_16719,N_16260);
or U17529 (N_17529,N_16380,N_16875);
nand U17530 (N_17530,N_16204,N_16454);
and U17531 (N_17531,N_16853,N_16015);
nand U17532 (N_17532,N_16803,N_16852);
or U17533 (N_17533,N_16753,N_16987);
and U17534 (N_17534,N_16652,N_16427);
nand U17535 (N_17535,N_16546,N_16109);
xnor U17536 (N_17536,N_16582,N_16649);
xor U17537 (N_17537,N_16152,N_16797);
nor U17538 (N_17538,N_16234,N_16758);
and U17539 (N_17539,N_16288,N_16163);
or U17540 (N_17540,N_16681,N_16787);
nand U17541 (N_17541,N_16460,N_16539);
and U17542 (N_17542,N_16933,N_16024);
nor U17543 (N_17543,N_16790,N_16556);
nand U17544 (N_17544,N_16610,N_16056);
nand U17545 (N_17545,N_16743,N_16972);
nor U17546 (N_17546,N_16759,N_16329);
and U17547 (N_17547,N_16962,N_16172);
xor U17548 (N_17548,N_16776,N_16319);
and U17549 (N_17549,N_16959,N_16579);
xor U17550 (N_17550,N_16433,N_16904);
nor U17551 (N_17551,N_16796,N_16459);
and U17552 (N_17552,N_16297,N_16366);
and U17553 (N_17553,N_16332,N_16326);
nand U17554 (N_17554,N_16408,N_16308);
and U17555 (N_17555,N_16793,N_16953);
xnor U17556 (N_17556,N_16435,N_16994);
and U17557 (N_17557,N_16952,N_16698);
xnor U17558 (N_17558,N_16872,N_16115);
nor U17559 (N_17559,N_16029,N_16137);
xor U17560 (N_17560,N_16846,N_16092);
xor U17561 (N_17561,N_16772,N_16591);
nor U17562 (N_17562,N_16764,N_16540);
nor U17563 (N_17563,N_16855,N_16070);
nand U17564 (N_17564,N_16062,N_16749);
or U17565 (N_17565,N_16560,N_16301);
and U17566 (N_17566,N_16633,N_16848);
or U17567 (N_17567,N_16474,N_16792);
nand U17568 (N_17568,N_16186,N_16019);
xor U17569 (N_17569,N_16086,N_16663);
nand U17570 (N_17570,N_16171,N_16336);
and U17571 (N_17571,N_16390,N_16417);
and U17572 (N_17572,N_16574,N_16349);
xor U17573 (N_17573,N_16545,N_16081);
nor U17574 (N_17574,N_16226,N_16345);
and U17575 (N_17575,N_16353,N_16977);
or U17576 (N_17576,N_16771,N_16631);
and U17577 (N_17577,N_16048,N_16214);
and U17578 (N_17578,N_16500,N_16081);
nor U17579 (N_17579,N_16215,N_16717);
and U17580 (N_17580,N_16632,N_16835);
nand U17581 (N_17581,N_16397,N_16358);
or U17582 (N_17582,N_16635,N_16154);
nor U17583 (N_17583,N_16948,N_16458);
and U17584 (N_17584,N_16584,N_16312);
or U17585 (N_17585,N_16123,N_16718);
and U17586 (N_17586,N_16374,N_16803);
and U17587 (N_17587,N_16968,N_16411);
or U17588 (N_17588,N_16511,N_16003);
nand U17589 (N_17589,N_16192,N_16335);
nand U17590 (N_17590,N_16054,N_16633);
xor U17591 (N_17591,N_16332,N_16719);
xnor U17592 (N_17592,N_16594,N_16501);
nor U17593 (N_17593,N_16972,N_16055);
nand U17594 (N_17594,N_16232,N_16915);
or U17595 (N_17595,N_16500,N_16460);
or U17596 (N_17596,N_16929,N_16668);
and U17597 (N_17597,N_16227,N_16984);
nor U17598 (N_17598,N_16178,N_16189);
nand U17599 (N_17599,N_16774,N_16734);
nand U17600 (N_17600,N_16145,N_16179);
nor U17601 (N_17601,N_16296,N_16425);
xnor U17602 (N_17602,N_16444,N_16509);
xnor U17603 (N_17603,N_16195,N_16858);
nand U17604 (N_17604,N_16786,N_16944);
or U17605 (N_17605,N_16476,N_16024);
xor U17606 (N_17606,N_16031,N_16867);
nand U17607 (N_17607,N_16271,N_16982);
nor U17608 (N_17608,N_16654,N_16313);
xnor U17609 (N_17609,N_16885,N_16034);
and U17610 (N_17610,N_16055,N_16704);
and U17611 (N_17611,N_16234,N_16039);
xor U17612 (N_17612,N_16151,N_16851);
xnor U17613 (N_17613,N_16627,N_16826);
or U17614 (N_17614,N_16581,N_16983);
nor U17615 (N_17615,N_16265,N_16180);
or U17616 (N_17616,N_16366,N_16949);
nand U17617 (N_17617,N_16431,N_16831);
nand U17618 (N_17618,N_16830,N_16969);
xnor U17619 (N_17619,N_16557,N_16392);
and U17620 (N_17620,N_16522,N_16505);
nand U17621 (N_17621,N_16622,N_16211);
or U17622 (N_17622,N_16114,N_16005);
nor U17623 (N_17623,N_16421,N_16165);
xor U17624 (N_17624,N_16739,N_16317);
and U17625 (N_17625,N_16683,N_16658);
xor U17626 (N_17626,N_16456,N_16065);
and U17627 (N_17627,N_16170,N_16010);
and U17628 (N_17628,N_16434,N_16154);
and U17629 (N_17629,N_16496,N_16736);
nand U17630 (N_17630,N_16912,N_16127);
nand U17631 (N_17631,N_16196,N_16112);
xnor U17632 (N_17632,N_16694,N_16963);
and U17633 (N_17633,N_16155,N_16502);
nor U17634 (N_17634,N_16529,N_16470);
and U17635 (N_17635,N_16983,N_16290);
and U17636 (N_17636,N_16562,N_16278);
and U17637 (N_17637,N_16440,N_16193);
xor U17638 (N_17638,N_16195,N_16972);
xnor U17639 (N_17639,N_16358,N_16747);
nand U17640 (N_17640,N_16546,N_16161);
nor U17641 (N_17641,N_16232,N_16341);
nor U17642 (N_17642,N_16253,N_16043);
nor U17643 (N_17643,N_16788,N_16052);
nand U17644 (N_17644,N_16185,N_16933);
or U17645 (N_17645,N_16446,N_16243);
nand U17646 (N_17646,N_16160,N_16558);
nand U17647 (N_17647,N_16845,N_16651);
nand U17648 (N_17648,N_16847,N_16966);
nand U17649 (N_17649,N_16797,N_16251);
nand U17650 (N_17650,N_16931,N_16465);
nand U17651 (N_17651,N_16654,N_16749);
nand U17652 (N_17652,N_16413,N_16458);
nand U17653 (N_17653,N_16730,N_16470);
nand U17654 (N_17654,N_16427,N_16760);
and U17655 (N_17655,N_16739,N_16003);
nand U17656 (N_17656,N_16468,N_16704);
and U17657 (N_17657,N_16761,N_16729);
and U17658 (N_17658,N_16589,N_16675);
nor U17659 (N_17659,N_16869,N_16473);
xnor U17660 (N_17660,N_16932,N_16096);
or U17661 (N_17661,N_16832,N_16957);
or U17662 (N_17662,N_16255,N_16202);
nand U17663 (N_17663,N_16513,N_16646);
or U17664 (N_17664,N_16559,N_16532);
xor U17665 (N_17665,N_16148,N_16642);
and U17666 (N_17666,N_16272,N_16186);
nor U17667 (N_17667,N_16499,N_16122);
nand U17668 (N_17668,N_16678,N_16238);
or U17669 (N_17669,N_16522,N_16715);
or U17670 (N_17670,N_16165,N_16785);
nand U17671 (N_17671,N_16310,N_16109);
nor U17672 (N_17672,N_16895,N_16080);
xnor U17673 (N_17673,N_16181,N_16709);
nand U17674 (N_17674,N_16569,N_16040);
xnor U17675 (N_17675,N_16958,N_16986);
and U17676 (N_17676,N_16116,N_16624);
xnor U17677 (N_17677,N_16364,N_16737);
nor U17678 (N_17678,N_16076,N_16222);
or U17679 (N_17679,N_16740,N_16798);
nor U17680 (N_17680,N_16468,N_16008);
nand U17681 (N_17681,N_16926,N_16002);
nand U17682 (N_17682,N_16059,N_16927);
nand U17683 (N_17683,N_16024,N_16564);
nor U17684 (N_17684,N_16524,N_16931);
xor U17685 (N_17685,N_16722,N_16054);
nor U17686 (N_17686,N_16535,N_16401);
nand U17687 (N_17687,N_16979,N_16468);
nand U17688 (N_17688,N_16399,N_16500);
nand U17689 (N_17689,N_16975,N_16829);
xor U17690 (N_17690,N_16905,N_16769);
nand U17691 (N_17691,N_16398,N_16369);
nand U17692 (N_17692,N_16969,N_16476);
xor U17693 (N_17693,N_16442,N_16000);
xor U17694 (N_17694,N_16809,N_16992);
xor U17695 (N_17695,N_16390,N_16756);
xnor U17696 (N_17696,N_16165,N_16970);
xnor U17697 (N_17697,N_16533,N_16576);
or U17698 (N_17698,N_16308,N_16559);
nand U17699 (N_17699,N_16974,N_16856);
nand U17700 (N_17700,N_16747,N_16016);
nand U17701 (N_17701,N_16599,N_16349);
and U17702 (N_17702,N_16421,N_16496);
or U17703 (N_17703,N_16077,N_16592);
and U17704 (N_17704,N_16767,N_16388);
nand U17705 (N_17705,N_16801,N_16421);
nor U17706 (N_17706,N_16612,N_16450);
and U17707 (N_17707,N_16590,N_16357);
nor U17708 (N_17708,N_16099,N_16524);
xnor U17709 (N_17709,N_16676,N_16823);
nand U17710 (N_17710,N_16041,N_16660);
or U17711 (N_17711,N_16922,N_16499);
nand U17712 (N_17712,N_16724,N_16859);
nor U17713 (N_17713,N_16586,N_16408);
and U17714 (N_17714,N_16039,N_16233);
and U17715 (N_17715,N_16460,N_16338);
or U17716 (N_17716,N_16967,N_16786);
and U17717 (N_17717,N_16910,N_16513);
and U17718 (N_17718,N_16856,N_16331);
or U17719 (N_17719,N_16713,N_16925);
or U17720 (N_17720,N_16788,N_16457);
nand U17721 (N_17721,N_16906,N_16541);
nor U17722 (N_17722,N_16566,N_16887);
nor U17723 (N_17723,N_16703,N_16881);
nand U17724 (N_17724,N_16671,N_16014);
xnor U17725 (N_17725,N_16343,N_16178);
or U17726 (N_17726,N_16389,N_16778);
nand U17727 (N_17727,N_16556,N_16212);
xor U17728 (N_17728,N_16632,N_16964);
nand U17729 (N_17729,N_16025,N_16697);
xor U17730 (N_17730,N_16053,N_16824);
and U17731 (N_17731,N_16749,N_16975);
and U17732 (N_17732,N_16619,N_16144);
or U17733 (N_17733,N_16009,N_16785);
nor U17734 (N_17734,N_16115,N_16455);
nand U17735 (N_17735,N_16793,N_16121);
and U17736 (N_17736,N_16315,N_16101);
and U17737 (N_17737,N_16239,N_16158);
and U17738 (N_17738,N_16882,N_16593);
or U17739 (N_17739,N_16643,N_16507);
or U17740 (N_17740,N_16808,N_16480);
or U17741 (N_17741,N_16769,N_16733);
xor U17742 (N_17742,N_16994,N_16268);
nand U17743 (N_17743,N_16275,N_16515);
or U17744 (N_17744,N_16507,N_16529);
or U17745 (N_17745,N_16785,N_16746);
nor U17746 (N_17746,N_16093,N_16566);
nand U17747 (N_17747,N_16143,N_16604);
or U17748 (N_17748,N_16957,N_16005);
nand U17749 (N_17749,N_16038,N_16216);
xor U17750 (N_17750,N_16622,N_16276);
or U17751 (N_17751,N_16986,N_16143);
or U17752 (N_17752,N_16250,N_16679);
xor U17753 (N_17753,N_16342,N_16772);
or U17754 (N_17754,N_16743,N_16266);
or U17755 (N_17755,N_16377,N_16873);
xnor U17756 (N_17756,N_16903,N_16728);
xor U17757 (N_17757,N_16602,N_16337);
or U17758 (N_17758,N_16644,N_16723);
xnor U17759 (N_17759,N_16326,N_16351);
nor U17760 (N_17760,N_16411,N_16379);
or U17761 (N_17761,N_16551,N_16936);
xnor U17762 (N_17762,N_16025,N_16858);
and U17763 (N_17763,N_16284,N_16335);
nor U17764 (N_17764,N_16106,N_16316);
nand U17765 (N_17765,N_16299,N_16258);
xor U17766 (N_17766,N_16655,N_16274);
nand U17767 (N_17767,N_16956,N_16930);
and U17768 (N_17768,N_16173,N_16637);
xor U17769 (N_17769,N_16296,N_16464);
nand U17770 (N_17770,N_16304,N_16129);
and U17771 (N_17771,N_16848,N_16159);
and U17772 (N_17772,N_16659,N_16650);
nor U17773 (N_17773,N_16054,N_16946);
and U17774 (N_17774,N_16701,N_16154);
xor U17775 (N_17775,N_16305,N_16806);
and U17776 (N_17776,N_16285,N_16980);
nor U17777 (N_17777,N_16854,N_16148);
xnor U17778 (N_17778,N_16999,N_16530);
and U17779 (N_17779,N_16237,N_16885);
nor U17780 (N_17780,N_16883,N_16687);
xor U17781 (N_17781,N_16809,N_16662);
or U17782 (N_17782,N_16869,N_16432);
or U17783 (N_17783,N_16821,N_16464);
nor U17784 (N_17784,N_16806,N_16881);
nor U17785 (N_17785,N_16272,N_16225);
xor U17786 (N_17786,N_16587,N_16964);
or U17787 (N_17787,N_16478,N_16531);
nor U17788 (N_17788,N_16309,N_16100);
or U17789 (N_17789,N_16945,N_16874);
and U17790 (N_17790,N_16798,N_16022);
and U17791 (N_17791,N_16857,N_16520);
xor U17792 (N_17792,N_16076,N_16276);
and U17793 (N_17793,N_16820,N_16003);
and U17794 (N_17794,N_16789,N_16222);
nor U17795 (N_17795,N_16154,N_16763);
nand U17796 (N_17796,N_16454,N_16503);
nor U17797 (N_17797,N_16336,N_16756);
xor U17798 (N_17798,N_16053,N_16982);
xnor U17799 (N_17799,N_16098,N_16706);
and U17800 (N_17800,N_16349,N_16966);
xnor U17801 (N_17801,N_16140,N_16580);
nand U17802 (N_17802,N_16407,N_16931);
nor U17803 (N_17803,N_16258,N_16002);
nand U17804 (N_17804,N_16133,N_16984);
or U17805 (N_17805,N_16208,N_16270);
xnor U17806 (N_17806,N_16528,N_16475);
nand U17807 (N_17807,N_16880,N_16326);
xor U17808 (N_17808,N_16850,N_16502);
nor U17809 (N_17809,N_16627,N_16129);
xnor U17810 (N_17810,N_16064,N_16231);
and U17811 (N_17811,N_16369,N_16680);
and U17812 (N_17812,N_16597,N_16755);
or U17813 (N_17813,N_16051,N_16083);
nand U17814 (N_17814,N_16506,N_16141);
nor U17815 (N_17815,N_16324,N_16947);
xnor U17816 (N_17816,N_16176,N_16747);
or U17817 (N_17817,N_16961,N_16321);
or U17818 (N_17818,N_16750,N_16493);
or U17819 (N_17819,N_16271,N_16459);
nand U17820 (N_17820,N_16833,N_16789);
nand U17821 (N_17821,N_16886,N_16311);
and U17822 (N_17822,N_16568,N_16836);
or U17823 (N_17823,N_16590,N_16970);
nor U17824 (N_17824,N_16247,N_16581);
or U17825 (N_17825,N_16129,N_16482);
nor U17826 (N_17826,N_16638,N_16298);
xnor U17827 (N_17827,N_16434,N_16966);
xor U17828 (N_17828,N_16714,N_16133);
or U17829 (N_17829,N_16113,N_16371);
nand U17830 (N_17830,N_16454,N_16517);
and U17831 (N_17831,N_16797,N_16385);
or U17832 (N_17832,N_16422,N_16469);
xnor U17833 (N_17833,N_16592,N_16393);
or U17834 (N_17834,N_16512,N_16782);
nor U17835 (N_17835,N_16887,N_16649);
and U17836 (N_17836,N_16499,N_16776);
nand U17837 (N_17837,N_16921,N_16363);
and U17838 (N_17838,N_16447,N_16370);
nand U17839 (N_17839,N_16918,N_16546);
and U17840 (N_17840,N_16099,N_16148);
and U17841 (N_17841,N_16641,N_16621);
or U17842 (N_17842,N_16013,N_16970);
or U17843 (N_17843,N_16724,N_16157);
and U17844 (N_17844,N_16170,N_16468);
nand U17845 (N_17845,N_16965,N_16419);
or U17846 (N_17846,N_16403,N_16810);
nor U17847 (N_17847,N_16424,N_16335);
xnor U17848 (N_17848,N_16797,N_16780);
nand U17849 (N_17849,N_16535,N_16989);
and U17850 (N_17850,N_16974,N_16033);
and U17851 (N_17851,N_16535,N_16988);
or U17852 (N_17852,N_16549,N_16792);
nor U17853 (N_17853,N_16606,N_16546);
and U17854 (N_17854,N_16419,N_16820);
nand U17855 (N_17855,N_16625,N_16620);
or U17856 (N_17856,N_16284,N_16579);
or U17857 (N_17857,N_16381,N_16826);
and U17858 (N_17858,N_16104,N_16551);
xor U17859 (N_17859,N_16714,N_16487);
or U17860 (N_17860,N_16039,N_16593);
or U17861 (N_17861,N_16630,N_16860);
or U17862 (N_17862,N_16731,N_16119);
or U17863 (N_17863,N_16555,N_16863);
nand U17864 (N_17864,N_16214,N_16674);
or U17865 (N_17865,N_16386,N_16888);
xnor U17866 (N_17866,N_16755,N_16757);
or U17867 (N_17867,N_16037,N_16079);
nor U17868 (N_17868,N_16472,N_16239);
and U17869 (N_17869,N_16389,N_16727);
nand U17870 (N_17870,N_16595,N_16426);
or U17871 (N_17871,N_16413,N_16570);
or U17872 (N_17872,N_16746,N_16734);
nand U17873 (N_17873,N_16396,N_16371);
xnor U17874 (N_17874,N_16543,N_16194);
xor U17875 (N_17875,N_16248,N_16152);
xor U17876 (N_17876,N_16384,N_16696);
nand U17877 (N_17877,N_16656,N_16088);
or U17878 (N_17878,N_16411,N_16211);
nor U17879 (N_17879,N_16008,N_16927);
xor U17880 (N_17880,N_16875,N_16929);
or U17881 (N_17881,N_16125,N_16346);
xnor U17882 (N_17882,N_16967,N_16547);
nand U17883 (N_17883,N_16531,N_16441);
xor U17884 (N_17884,N_16359,N_16103);
or U17885 (N_17885,N_16956,N_16199);
and U17886 (N_17886,N_16306,N_16928);
nor U17887 (N_17887,N_16870,N_16534);
and U17888 (N_17888,N_16452,N_16739);
nor U17889 (N_17889,N_16403,N_16699);
or U17890 (N_17890,N_16587,N_16482);
and U17891 (N_17891,N_16177,N_16932);
xor U17892 (N_17892,N_16781,N_16449);
and U17893 (N_17893,N_16544,N_16402);
nor U17894 (N_17894,N_16475,N_16594);
xnor U17895 (N_17895,N_16786,N_16458);
and U17896 (N_17896,N_16917,N_16586);
nand U17897 (N_17897,N_16061,N_16841);
nor U17898 (N_17898,N_16832,N_16668);
xor U17899 (N_17899,N_16345,N_16922);
and U17900 (N_17900,N_16882,N_16533);
or U17901 (N_17901,N_16323,N_16733);
nor U17902 (N_17902,N_16272,N_16227);
and U17903 (N_17903,N_16812,N_16694);
and U17904 (N_17904,N_16919,N_16230);
xnor U17905 (N_17905,N_16750,N_16483);
or U17906 (N_17906,N_16500,N_16941);
and U17907 (N_17907,N_16733,N_16400);
nand U17908 (N_17908,N_16080,N_16976);
xnor U17909 (N_17909,N_16904,N_16964);
xnor U17910 (N_17910,N_16283,N_16700);
and U17911 (N_17911,N_16552,N_16013);
nor U17912 (N_17912,N_16944,N_16614);
nor U17913 (N_17913,N_16522,N_16589);
xor U17914 (N_17914,N_16003,N_16437);
xor U17915 (N_17915,N_16870,N_16484);
nand U17916 (N_17916,N_16615,N_16009);
xor U17917 (N_17917,N_16283,N_16424);
xor U17918 (N_17918,N_16906,N_16639);
nand U17919 (N_17919,N_16731,N_16148);
nor U17920 (N_17920,N_16253,N_16225);
nand U17921 (N_17921,N_16830,N_16920);
nand U17922 (N_17922,N_16395,N_16825);
and U17923 (N_17923,N_16644,N_16096);
or U17924 (N_17924,N_16204,N_16519);
xnor U17925 (N_17925,N_16225,N_16745);
nand U17926 (N_17926,N_16412,N_16647);
xor U17927 (N_17927,N_16289,N_16046);
nand U17928 (N_17928,N_16783,N_16922);
and U17929 (N_17929,N_16844,N_16785);
xnor U17930 (N_17930,N_16996,N_16207);
or U17931 (N_17931,N_16925,N_16221);
or U17932 (N_17932,N_16718,N_16747);
nor U17933 (N_17933,N_16700,N_16408);
and U17934 (N_17934,N_16187,N_16621);
or U17935 (N_17935,N_16552,N_16088);
nand U17936 (N_17936,N_16134,N_16794);
xor U17937 (N_17937,N_16842,N_16651);
xor U17938 (N_17938,N_16333,N_16744);
xor U17939 (N_17939,N_16893,N_16521);
nor U17940 (N_17940,N_16659,N_16463);
nor U17941 (N_17941,N_16639,N_16553);
nor U17942 (N_17942,N_16960,N_16036);
xor U17943 (N_17943,N_16157,N_16776);
nand U17944 (N_17944,N_16306,N_16592);
nand U17945 (N_17945,N_16266,N_16155);
nor U17946 (N_17946,N_16942,N_16846);
and U17947 (N_17947,N_16746,N_16469);
nand U17948 (N_17948,N_16756,N_16986);
and U17949 (N_17949,N_16397,N_16872);
xnor U17950 (N_17950,N_16464,N_16098);
and U17951 (N_17951,N_16471,N_16274);
and U17952 (N_17952,N_16912,N_16432);
nor U17953 (N_17953,N_16296,N_16827);
nand U17954 (N_17954,N_16286,N_16352);
and U17955 (N_17955,N_16170,N_16047);
or U17956 (N_17956,N_16626,N_16620);
xor U17957 (N_17957,N_16963,N_16889);
nand U17958 (N_17958,N_16549,N_16608);
nor U17959 (N_17959,N_16902,N_16662);
xor U17960 (N_17960,N_16358,N_16382);
xor U17961 (N_17961,N_16673,N_16721);
xnor U17962 (N_17962,N_16211,N_16753);
nor U17963 (N_17963,N_16358,N_16370);
nor U17964 (N_17964,N_16747,N_16741);
nand U17965 (N_17965,N_16292,N_16601);
xnor U17966 (N_17966,N_16153,N_16146);
or U17967 (N_17967,N_16236,N_16101);
xnor U17968 (N_17968,N_16530,N_16772);
or U17969 (N_17969,N_16924,N_16552);
xnor U17970 (N_17970,N_16188,N_16383);
nor U17971 (N_17971,N_16631,N_16808);
nand U17972 (N_17972,N_16935,N_16340);
xnor U17973 (N_17973,N_16047,N_16294);
nand U17974 (N_17974,N_16638,N_16407);
nor U17975 (N_17975,N_16787,N_16620);
and U17976 (N_17976,N_16397,N_16505);
xor U17977 (N_17977,N_16771,N_16025);
or U17978 (N_17978,N_16127,N_16887);
or U17979 (N_17979,N_16860,N_16992);
nor U17980 (N_17980,N_16576,N_16397);
xor U17981 (N_17981,N_16680,N_16508);
and U17982 (N_17982,N_16282,N_16861);
xnor U17983 (N_17983,N_16825,N_16396);
and U17984 (N_17984,N_16840,N_16483);
xnor U17985 (N_17985,N_16736,N_16005);
and U17986 (N_17986,N_16283,N_16094);
nor U17987 (N_17987,N_16319,N_16413);
nor U17988 (N_17988,N_16778,N_16240);
nand U17989 (N_17989,N_16404,N_16330);
nor U17990 (N_17990,N_16852,N_16678);
and U17991 (N_17991,N_16827,N_16055);
nand U17992 (N_17992,N_16301,N_16631);
nor U17993 (N_17993,N_16639,N_16813);
nand U17994 (N_17994,N_16438,N_16709);
nor U17995 (N_17995,N_16617,N_16585);
or U17996 (N_17996,N_16447,N_16023);
xor U17997 (N_17997,N_16652,N_16642);
nor U17998 (N_17998,N_16249,N_16326);
xnor U17999 (N_17999,N_16450,N_16084);
and U18000 (N_18000,N_17784,N_17605);
and U18001 (N_18001,N_17333,N_17819);
or U18002 (N_18002,N_17782,N_17561);
nand U18003 (N_18003,N_17789,N_17729);
or U18004 (N_18004,N_17715,N_17828);
xnor U18005 (N_18005,N_17946,N_17049);
or U18006 (N_18006,N_17877,N_17171);
and U18007 (N_18007,N_17960,N_17211);
xnor U18008 (N_18008,N_17385,N_17339);
or U18009 (N_18009,N_17697,N_17095);
nor U18010 (N_18010,N_17160,N_17735);
xor U18011 (N_18011,N_17806,N_17939);
xnor U18012 (N_18012,N_17815,N_17210);
and U18013 (N_18013,N_17928,N_17499);
nand U18014 (N_18014,N_17415,N_17080);
nand U18015 (N_18015,N_17014,N_17713);
or U18016 (N_18016,N_17324,N_17734);
xor U18017 (N_18017,N_17249,N_17243);
or U18018 (N_18018,N_17259,N_17525);
and U18019 (N_18019,N_17406,N_17477);
nor U18020 (N_18020,N_17889,N_17360);
and U18021 (N_18021,N_17368,N_17530);
or U18022 (N_18022,N_17706,N_17149);
xor U18023 (N_18023,N_17309,N_17809);
xor U18024 (N_18024,N_17232,N_17754);
nor U18025 (N_18025,N_17279,N_17817);
xor U18026 (N_18026,N_17076,N_17293);
nand U18027 (N_18027,N_17808,N_17265);
and U18028 (N_18028,N_17476,N_17051);
nand U18029 (N_18029,N_17114,N_17423);
nor U18030 (N_18030,N_17214,N_17518);
nand U18031 (N_18031,N_17134,N_17995);
and U18032 (N_18032,N_17804,N_17185);
xnor U18033 (N_18033,N_17359,N_17304);
nor U18034 (N_18034,N_17773,N_17927);
and U18035 (N_18035,N_17282,N_17341);
and U18036 (N_18036,N_17041,N_17987);
nand U18037 (N_18037,N_17197,N_17720);
xnor U18038 (N_18038,N_17418,N_17497);
and U18039 (N_18039,N_17913,N_17202);
or U18040 (N_18040,N_17492,N_17981);
nand U18041 (N_18041,N_17945,N_17598);
nor U18042 (N_18042,N_17200,N_17167);
and U18043 (N_18043,N_17206,N_17964);
or U18044 (N_18044,N_17609,N_17148);
nand U18045 (N_18045,N_17907,N_17740);
xnor U18046 (N_18046,N_17387,N_17066);
nand U18047 (N_18047,N_17331,N_17624);
xor U18048 (N_18048,N_17544,N_17676);
xnor U18049 (N_18049,N_17294,N_17412);
nand U18050 (N_18050,N_17348,N_17771);
nor U18051 (N_18051,N_17400,N_17498);
xnor U18052 (N_18052,N_17778,N_17527);
or U18053 (N_18053,N_17107,N_17025);
xor U18054 (N_18054,N_17108,N_17958);
xnor U18055 (N_18055,N_17356,N_17366);
or U18056 (N_18056,N_17422,N_17668);
xnor U18057 (N_18057,N_17541,N_17156);
xor U18058 (N_18058,N_17112,N_17702);
xor U18059 (N_18059,N_17984,N_17277);
and U18060 (N_18060,N_17959,N_17338);
or U18061 (N_18061,N_17435,N_17965);
nand U18062 (N_18062,N_17557,N_17452);
xnor U18063 (N_18063,N_17845,N_17005);
nor U18064 (N_18064,N_17260,N_17208);
xor U18065 (N_18065,N_17468,N_17161);
or U18066 (N_18066,N_17409,N_17831);
xor U18067 (N_18067,N_17736,N_17421);
nor U18068 (N_18068,N_17645,N_17336);
nor U18069 (N_18069,N_17128,N_17977);
xnor U18070 (N_18070,N_17417,N_17038);
xnor U18071 (N_18071,N_17508,N_17627);
xnor U18072 (N_18072,N_17425,N_17334);
nand U18073 (N_18073,N_17576,N_17162);
and U18074 (N_18074,N_17097,N_17432);
and U18075 (N_18075,N_17355,N_17876);
and U18076 (N_18076,N_17060,N_17071);
nand U18077 (N_18077,N_17219,N_17367);
nand U18078 (N_18078,N_17229,N_17626);
xor U18079 (N_18079,N_17257,N_17591);
nor U18080 (N_18080,N_17859,N_17788);
nor U18081 (N_18081,N_17374,N_17140);
xnor U18082 (N_18082,N_17398,N_17622);
and U18083 (N_18083,N_17079,N_17253);
nand U18084 (N_18084,N_17337,N_17892);
xor U18085 (N_18085,N_17388,N_17816);
and U18086 (N_18086,N_17436,N_17985);
xor U18087 (N_18087,N_17711,N_17667);
xor U18088 (N_18088,N_17188,N_17446);
nand U18089 (N_18089,N_17064,N_17004);
or U18090 (N_18090,N_17662,N_17558);
or U18091 (N_18091,N_17872,N_17708);
nand U18092 (N_18092,N_17777,N_17261);
xor U18093 (N_18093,N_17564,N_17144);
xor U18094 (N_18094,N_17491,N_17292);
nand U18095 (N_18095,N_17612,N_17517);
xor U18096 (N_18096,N_17187,N_17369);
or U18097 (N_18097,N_17587,N_17670);
and U18098 (N_18098,N_17967,N_17693);
or U18099 (N_18099,N_17472,N_17864);
and U18100 (N_18100,N_17552,N_17154);
nand U18101 (N_18101,N_17513,N_17424);
nor U18102 (N_18102,N_17048,N_17930);
nor U18103 (N_18103,N_17669,N_17785);
nor U18104 (N_18104,N_17094,N_17024);
and U18105 (N_18105,N_17482,N_17019);
and U18106 (N_18106,N_17999,N_17190);
nor U18107 (N_18107,N_17323,N_17286);
or U18108 (N_18108,N_17386,N_17506);
nor U18109 (N_18109,N_17177,N_17860);
nand U18110 (N_18110,N_17365,N_17798);
or U18111 (N_18111,N_17358,N_17245);
nor U18112 (N_18112,N_17057,N_17873);
xor U18113 (N_18113,N_17298,N_17616);
nor U18114 (N_18114,N_17281,N_17511);
and U18115 (N_18115,N_17794,N_17272);
nor U18116 (N_18116,N_17870,N_17878);
or U18117 (N_18117,N_17078,N_17081);
xnor U18118 (N_18118,N_17586,N_17610);
or U18119 (N_18119,N_17343,N_17940);
and U18120 (N_18120,N_17110,N_17638);
xor U18121 (N_18121,N_17002,N_17549);
or U18122 (N_18122,N_17833,N_17299);
and U18123 (N_18123,N_17650,N_17901);
nor U18124 (N_18124,N_17050,N_17838);
nand U18125 (N_18125,N_17373,N_17532);
xor U18126 (N_18126,N_17361,N_17514);
nor U18127 (N_18127,N_17931,N_17969);
nand U18128 (N_18128,N_17699,N_17628);
nand U18129 (N_18129,N_17893,N_17908);
nor U18130 (N_18130,N_17803,N_17534);
and U18131 (N_18131,N_17915,N_17755);
nand U18132 (N_18132,N_17199,N_17853);
or U18133 (N_18133,N_17462,N_17580);
or U18134 (N_18134,N_17251,N_17775);
xnor U18135 (N_18135,N_17102,N_17222);
xnor U18136 (N_18136,N_17133,N_17316);
xnor U18137 (N_18137,N_17320,N_17707);
nand U18138 (N_18138,N_17342,N_17768);
xnor U18139 (N_18139,N_17998,N_17625);
and U18140 (N_18140,N_17642,N_17207);
or U18141 (N_18141,N_17619,N_17973);
nand U18142 (N_18142,N_17158,N_17413);
nor U18143 (N_18143,N_17035,N_17994);
xor U18144 (N_18144,N_17218,N_17220);
nand U18145 (N_18145,N_17681,N_17377);
nor U18146 (N_18146,N_17380,N_17568);
and U18147 (N_18147,N_17692,N_17602);
or U18148 (N_18148,N_17463,N_17537);
and U18149 (N_18149,N_17685,N_17046);
or U18150 (N_18150,N_17906,N_17332);
xor U18151 (N_18151,N_17533,N_17440);
nor U18152 (N_18152,N_17879,N_17471);
or U18153 (N_18153,N_17826,N_17573);
nand U18154 (N_18154,N_17954,N_17791);
nand U18155 (N_18155,N_17405,N_17396);
xnor U18156 (N_18156,N_17478,N_17980);
nand U18157 (N_18157,N_17847,N_17466);
nor U18158 (N_18158,N_17957,N_17767);
and U18159 (N_18159,N_17712,N_17894);
nand U18160 (N_18160,N_17854,N_17291);
nor U18161 (N_18161,N_17666,N_17684);
xor U18162 (N_18162,N_17397,N_17834);
nand U18163 (N_18163,N_17869,N_17588);
and U18164 (N_18164,N_17234,N_17084);
nor U18165 (N_18165,N_17978,N_17454);
nor U18166 (N_18166,N_17792,N_17748);
and U18167 (N_18167,N_17636,N_17705);
xor U18168 (N_18168,N_17459,N_17383);
nor U18169 (N_18169,N_17473,N_17696);
or U18170 (N_18170,N_17236,N_17495);
and U18171 (N_18171,N_17820,N_17012);
nor U18172 (N_18172,N_17270,N_17678);
nand U18173 (N_18173,N_17848,N_17515);
xnor U18174 (N_18174,N_17934,N_17258);
and U18175 (N_18175,N_17614,N_17657);
or U18176 (N_18176,N_17083,N_17577);
nor U18177 (N_18177,N_17223,N_17011);
nand U18178 (N_18178,N_17918,N_17480);
xor U18179 (N_18179,N_17599,N_17151);
nor U18180 (N_18180,N_17111,N_17121);
nor U18181 (N_18181,N_17022,N_17240);
nor U18182 (N_18182,N_17840,N_17393);
nor U18183 (N_18183,N_17399,N_17392);
nand U18184 (N_18184,N_17929,N_17503);
or U18185 (N_18185,N_17823,N_17419);
or U18186 (N_18186,N_17867,N_17173);
xor U18187 (N_18187,N_17126,N_17528);
nand U18188 (N_18188,N_17841,N_17008);
nand U18189 (N_18189,N_17030,N_17013);
xnor U18190 (N_18190,N_17615,N_17956);
nand U18191 (N_18191,N_17664,N_17852);
or U18192 (N_18192,N_17802,N_17890);
nand U18193 (N_18193,N_17065,N_17920);
nand U18194 (N_18194,N_17724,N_17021);
nor U18195 (N_18195,N_17578,N_17150);
and U18196 (N_18196,N_17328,N_17354);
nand U18197 (N_18197,N_17861,N_17501);
and U18198 (N_18198,N_17225,N_17096);
or U18199 (N_18199,N_17824,N_17020);
and U18200 (N_18200,N_17944,N_17077);
or U18201 (N_18201,N_17512,N_17063);
or U18202 (N_18202,N_17592,N_17611);
or U18203 (N_18203,N_17988,N_17683);
xor U18204 (N_18204,N_17589,N_17040);
or U18205 (N_18205,N_17641,N_17091);
xnor U18206 (N_18206,N_17475,N_17175);
xor U18207 (N_18207,N_17490,N_17671);
or U18208 (N_18208,N_17857,N_17779);
and U18209 (N_18209,N_17655,N_17054);
xnor U18210 (N_18210,N_17204,N_17875);
nor U18211 (N_18211,N_17345,N_17898);
nor U18212 (N_18212,N_17523,N_17797);
nor U18213 (N_18213,N_17036,N_17474);
nand U18214 (N_18214,N_17590,N_17431);
xnor U18215 (N_18215,N_17215,N_17520);
nand U18216 (N_18216,N_17379,N_17357);
xnor U18217 (N_18217,N_17143,N_17271);
or U18218 (N_18218,N_17909,N_17353);
or U18219 (N_18219,N_17917,N_17184);
xor U18220 (N_18220,N_17248,N_17540);
and U18221 (N_18221,N_17163,N_17902);
xnor U18222 (N_18222,N_17437,N_17007);
xnor U18223 (N_18223,N_17903,N_17769);
xor U18224 (N_18224,N_17029,N_17453);
and U18225 (N_18225,N_17043,N_17009);
xnor U18226 (N_18226,N_17763,N_17562);
nor U18227 (N_18227,N_17716,N_17688);
xor U18228 (N_18228,N_17582,N_17147);
nand U18229 (N_18229,N_17526,N_17951);
nor U18230 (N_18230,N_17193,N_17070);
and U18231 (N_18231,N_17411,N_17465);
or U18232 (N_18232,N_17827,N_17179);
or U18233 (N_18233,N_17932,N_17686);
and U18234 (N_18234,N_17752,N_17855);
nand U18235 (N_18235,N_17765,N_17394);
and U18236 (N_18236,N_17275,N_17521);
nand U18237 (N_18237,N_17262,N_17774);
nand U18238 (N_18238,N_17201,N_17326);
nand U18239 (N_18239,N_17254,N_17566);
xor U18240 (N_18240,N_17382,N_17756);
and U18241 (N_18241,N_17829,N_17226);
and U18242 (N_18242,N_17743,N_17205);
nand U18243 (N_18243,N_17153,N_17087);
and U18244 (N_18244,N_17584,N_17289);
nor U18245 (N_18245,N_17677,N_17673);
or U18246 (N_18246,N_17255,N_17213);
nor U18247 (N_18247,N_17072,N_17180);
xor U18248 (N_18248,N_17347,N_17674);
and U18249 (N_18249,N_17821,N_17168);
nand U18250 (N_18250,N_17749,N_17547);
and U18251 (N_18251,N_17659,N_17123);
xor U18252 (N_18252,N_17737,N_17905);
xor U18253 (N_18253,N_17722,N_17125);
nand U18254 (N_18254,N_17037,N_17950);
xor U18255 (N_18255,N_17924,N_17658);
and U18256 (N_18256,N_17181,N_17027);
xnor U18257 (N_18257,N_17943,N_17648);
xnor U18258 (N_18258,N_17886,N_17799);
and U18259 (N_18259,N_17766,N_17224);
and U18260 (N_18260,N_17594,N_17186);
nor U18261 (N_18261,N_17451,N_17672);
xor U18262 (N_18262,N_17993,N_17138);
nand U18263 (N_18263,N_17241,N_17340);
xnor U18264 (N_18264,N_17941,N_17370);
nand U18265 (N_18265,N_17306,N_17493);
or U18266 (N_18266,N_17739,N_17704);
and U18267 (N_18267,N_17753,N_17433);
nor U18268 (N_18268,N_17026,N_17295);
or U18269 (N_18269,N_17308,N_17550);
xor U18270 (N_18270,N_17572,N_17384);
nand U18271 (N_18271,N_17656,N_17408);
xnor U18272 (N_18272,N_17703,N_17485);
nor U18273 (N_18273,N_17145,N_17962);
nand U18274 (N_18274,N_17073,N_17165);
and U18275 (N_18275,N_17885,N_17300);
nor U18276 (N_18276,N_17567,N_17970);
nand U18277 (N_18277,N_17313,N_17868);
nor U18278 (N_18278,N_17429,N_17975);
or U18279 (N_18279,N_17146,N_17483);
or U18280 (N_18280,N_17719,N_17100);
nand U18281 (N_18281,N_17912,N_17209);
and U18282 (N_18282,N_17212,N_17001);
and U18283 (N_18283,N_17710,N_17882);
nand U18284 (N_18284,N_17953,N_17727);
and U18285 (N_18285,N_17653,N_17067);
nor U18286 (N_18286,N_17757,N_17113);
nand U18287 (N_18287,N_17629,N_17644);
nand U18288 (N_18288,N_17319,N_17585);
nand U18289 (N_18289,N_17764,N_17844);
nand U18290 (N_18290,N_17937,N_17500);
xnor U18291 (N_18291,N_17176,N_17938);
xnor U18292 (N_18292,N_17575,N_17947);
or U18293 (N_18293,N_17198,N_17455);
nand U18294 (N_18294,N_17427,N_17839);
xor U18295 (N_18295,N_17709,N_17936);
and U18296 (N_18296,N_17781,N_17871);
xor U18297 (N_18297,N_17330,N_17438);
and U18298 (N_18298,N_17301,N_17690);
nand U18299 (N_18299,N_17082,N_17115);
xor U18300 (N_18300,N_17510,N_17730);
nand U18301 (N_18301,N_17652,N_17194);
nand U18302 (N_18302,N_17269,N_17595);
xor U18303 (N_18303,N_17296,N_17888);
nand U18304 (N_18304,N_17505,N_17256);
and U18305 (N_18305,N_17135,N_17329);
xnor U18306 (N_18306,N_17098,N_17276);
nand U18307 (N_18307,N_17793,N_17762);
and U18308 (N_18308,N_17812,N_17682);
nand U18309 (N_18309,N_17601,N_17312);
or U18310 (N_18310,N_17439,N_17085);
nor U18311 (N_18311,N_17911,N_17159);
and U18312 (N_18312,N_17621,N_17891);
or U18313 (N_18313,N_17571,N_17606);
and U18314 (N_18314,N_17059,N_17000);
and U18315 (N_18315,N_17430,N_17479);
nand U18316 (N_18316,N_17559,N_17310);
xnor U18317 (N_18317,N_17127,N_17910);
and U18318 (N_18318,N_17443,N_17221);
xor U18319 (N_18319,N_17287,N_17441);
nor U18320 (N_18320,N_17718,N_17372);
xor U18321 (N_18321,N_17700,N_17391);
xor U18322 (N_18322,N_17649,N_17402);
or U18323 (N_18323,N_17786,N_17244);
xnor U18324 (N_18324,N_17237,N_17457);
xor U18325 (N_18325,N_17783,N_17172);
xor U18326 (N_18326,N_17813,N_17280);
or U18327 (N_18327,N_17811,N_17543);
nor U18328 (N_18328,N_17874,N_17866);
or U18329 (N_18329,N_17851,N_17494);
and U18330 (N_18330,N_17132,N_17556);
or U18331 (N_18331,N_17613,N_17758);
and U18332 (N_18332,N_17721,N_17426);
and U18333 (N_18333,N_17105,N_17264);
nor U18334 (N_18334,N_17694,N_17850);
nor U18335 (N_18335,N_17631,N_17315);
nor U18336 (N_18336,N_17089,N_17991);
or U18337 (N_18337,N_17235,N_17502);
or U18338 (N_18338,N_17801,N_17887);
nand U18339 (N_18339,N_17344,N_17290);
xor U18340 (N_18340,N_17182,N_17434);
and U18341 (N_18341,N_17191,N_17058);
xor U18342 (N_18342,N_17003,N_17675);
nor U18343 (N_18343,N_17217,N_17742);
nand U18344 (N_18344,N_17461,N_17569);
and U18345 (N_18345,N_17522,N_17481);
or U18346 (N_18346,N_17551,N_17227);
nor U18347 (N_18347,N_17189,N_17583);
xnor U18348 (N_18348,N_17170,N_17283);
and U18349 (N_18349,N_17028,N_17099);
and U18350 (N_18350,N_17992,N_17375);
and U18351 (N_18351,N_17178,N_17689);
and U18352 (N_18352,N_17327,N_17103);
nand U18353 (N_18353,N_17196,N_17023);
nand U18354 (N_18354,N_17942,N_17088);
nand U18355 (N_18355,N_17725,N_17728);
xnor U18356 (N_18356,N_17321,N_17900);
and U18357 (N_18357,N_17104,N_17516);
nor U18358 (N_18358,N_17444,N_17553);
xor U18359 (N_18359,N_17899,N_17832);
nand U18360 (N_18360,N_17536,N_17835);
and U18361 (N_18361,N_17897,N_17266);
or U18362 (N_18362,N_17273,N_17056);
xor U18363 (N_18363,N_17531,N_17267);
nor U18364 (N_18364,N_17053,N_17968);
or U18365 (N_18365,N_17935,N_17796);
and U18366 (N_18366,N_17284,N_17318);
nand U18367 (N_18367,N_17810,N_17288);
nand U18368 (N_18368,N_17488,N_17130);
or U18369 (N_18369,N_17371,N_17731);
nor U18370 (N_18370,N_17252,N_17131);
nand U18371 (N_18371,N_17990,N_17116);
or U18372 (N_18372,N_17895,N_17574);
or U18373 (N_18373,N_17381,N_17842);
or U18374 (N_18374,N_17555,N_17971);
nand U18375 (N_18375,N_17747,N_17447);
or U18376 (N_18376,N_17546,N_17539);
nand U18377 (N_18377,N_17617,N_17033);
nor U18378 (N_18378,N_17118,N_17976);
or U18379 (N_18379,N_17790,N_17741);
or U18380 (N_18380,N_17389,N_17925);
xor U18381 (N_18381,N_17849,N_17603);
xor U18382 (N_18382,N_17579,N_17896);
and U18383 (N_18383,N_17955,N_17322);
or U18384 (N_18384,N_17701,N_17805);
xor U18385 (N_18385,N_17120,N_17018);
nand U18386 (N_18386,N_17166,N_17744);
nor U18387 (N_18387,N_17124,N_17966);
or U18388 (N_18388,N_17654,N_17129);
xnor U18389 (N_18389,N_17509,N_17407);
or U18390 (N_18390,N_17620,N_17157);
nor U18391 (N_18391,N_17442,N_17017);
and U18392 (N_18392,N_17274,N_17069);
or U18393 (N_18393,N_17750,N_17302);
nor U18394 (N_18394,N_17679,N_17448);
or U18395 (N_18395,N_17926,N_17307);
and U18396 (N_18396,N_17403,N_17632);
xor U18397 (N_18397,N_17618,N_17390);
or U18398 (N_18398,N_17643,N_17800);
and U18399 (N_18399,N_17242,N_17695);
xnor U18400 (N_18400,N_17231,N_17093);
xor U18401 (N_18401,N_17010,N_17404);
and U18402 (N_18402,N_17570,N_17152);
and U18403 (N_18403,N_17075,N_17691);
nor U18404 (N_18404,N_17351,N_17414);
and U18405 (N_18405,N_17814,N_17663);
and U18406 (N_18406,N_17548,N_17770);
xor U18407 (N_18407,N_17305,N_17445);
and U18408 (N_18408,N_17600,N_17881);
or U18409 (N_18409,N_17062,N_17487);
nor U18410 (N_18410,N_17880,N_17428);
or U18411 (N_18411,N_17136,N_17045);
nand U18412 (N_18412,N_17665,N_17660);
nand U18413 (N_18413,N_17714,N_17122);
nor U18414 (N_18414,N_17015,N_17883);
nand U18415 (N_18415,N_17637,N_17634);
and U18416 (N_18416,N_17865,N_17921);
or U18417 (N_18417,N_17593,N_17496);
or U18418 (N_18418,N_17504,N_17856);
nor U18419 (N_18419,N_17489,N_17216);
or U18420 (N_18420,N_17352,N_17738);
nor U18421 (N_18421,N_17787,N_17031);
and U18422 (N_18422,N_17006,N_17449);
nand U18423 (N_18423,N_17760,N_17646);
or U18424 (N_18424,N_17723,N_17119);
xor U18425 (N_18425,N_17914,N_17233);
or U18426 (N_18426,N_17807,N_17884);
nor U18427 (N_18427,N_17933,N_17680);
xor U18428 (N_18428,N_17607,N_17963);
and U18429 (N_18429,N_17979,N_17948);
and U18430 (N_18430,N_17349,N_17923);
or U18431 (N_18431,N_17862,N_17246);
or U18432 (N_18432,N_17106,N_17346);
nand U18433 (N_18433,N_17164,N_17142);
xnor U18434 (N_18434,N_17363,N_17263);
nand U18435 (N_18435,N_17239,N_17268);
nand U18436 (N_18436,N_17604,N_17410);
nand U18437 (N_18437,N_17795,N_17733);
nor U18438 (N_18438,N_17401,N_17238);
or U18439 (N_18439,N_17169,N_17846);
and U18440 (N_18440,N_17825,N_17623);
nand U18441 (N_18441,N_17044,N_17109);
nor U18442 (N_18442,N_17751,N_17032);
nand U18443 (N_18443,N_17362,N_17989);
nor U18444 (N_18444,N_17630,N_17836);
nand U18445 (N_18445,N_17545,N_17916);
nand U18446 (N_18446,N_17378,N_17818);
and U18447 (N_18447,N_17250,N_17780);
and U18448 (N_18448,N_17635,N_17843);
xnor U18449 (N_18449,N_17117,N_17155);
or U18450 (N_18450,N_17192,N_17470);
nand U18451 (N_18451,N_17542,N_17822);
nor U18452 (N_18452,N_17524,N_17230);
and U18453 (N_18453,N_17055,N_17858);
or U18454 (N_18454,N_17061,N_17174);
xnor U18455 (N_18455,N_17460,N_17139);
or U18456 (N_18456,N_17317,N_17297);
xnor U18457 (N_18457,N_17863,N_17376);
or U18458 (N_18458,N_17195,N_17464);
nor U18459 (N_18459,N_17074,N_17974);
and U18460 (N_18460,N_17687,N_17034);
or U18461 (N_18461,N_17467,N_17484);
or U18462 (N_18462,N_17228,N_17047);
or U18463 (N_18463,N_17554,N_17972);
nand U18464 (N_18464,N_17997,N_17904);
nor U18465 (N_18465,N_17647,N_17303);
xnor U18466 (N_18466,N_17952,N_17086);
nand U18467 (N_18467,N_17042,N_17746);
and U18468 (N_18468,N_17052,N_17639);
xnor U18469 (N_18469,N_17486,N_17519);
and U18470 (N_18470,N_17325,N_17581);
xnor U18471 (N_18471,N_17830,N_17450);
xor U18472 (N_18472,N_17597,N_17458);
xnor U18473 (N_18473,N_17068,N_17538);
xor U18474 (N_18474,N_17016,N_17247);
and U18475 (N_18475,N_17311,N_17772);
and U18476 (N_18476,N_17919,N_17092);
or U18477 (N_18477,N_17141,N_17314);
nand U18478 (N_18478,N_17633,N_17278);
nor U18479 (N_18479,N_17698,N_17745);
nand U18480 (N_18480,N_17469,N_17364);
nand U18481 (N_18481,N_17759,N_17651);
xnor U18482 (N_18482,N_17640,N_17285);
xor U18483 (N_18483,N_17732,N_17507);
xor U18484 (N_18484,N_17761,N_17456);
nor U18485 (N_18485,N_17395,N_17983);
and U18486 (N_18486,N_17726,N_17420);
and U18487 (N_18487,N_17986,N_17776);
xnor U18488 (N_18488,N_17560,N_17661);
xnor U18489 (N_18489,N_17608,N_17416);
and U18490 (N_18490,N_17535,N_17137);
or U18491 (N_18491,N_17717,N_17529);
xor U18492 (N_18492,N_17203,N_17350);
nor U18493 (N_18493,N_17596,N_17335);
and U18494 (N_18494,N_17949,N_17090);
xnor U18495 (N_18495,N_17563,N_17837);
nand U18496 (N_18496,N_17101,N_17961);
and U18497 (N_18497,N_17996,N_17922);
or U18498 (N_18498,N_17183,N_17565);
nor U18499 (N_18499,N_17039,N_17982);
nand U18500 (N_18500,N_17424,N_17123);
and U18501 (N_18501,N_17755,N_17609);
nor U18502 (N_18502,N_17222,N_17724);
or U18503 (N_18503,N_17746,N_17866);
or U18504 (N_18504,N_17801,N_17141);
nor U18505 (N_18505,N_17556,N_17736);
xnor U18506 (N_18506,N_17214,N_17683);
nor U18507 (N_18507,N_17607,N_17621);
nor U18508 (N_18508,N_17373,N_17648);
and U18509 (N_18509,N_17459,N_17607);
nor U18510 (N_18510,N_17123,N_17028);
xor U18511 (N_18511,N_17646,N_17966);
or U18512 (N_18512,N_17772,N_17237);
or U18513 (N_18513,N_17392,N_17150);
nand U18514 (N_18514,N_17697,N_17920);
or U18515 (N_18515,N_17665,N_17720);
nor U18516 (N_18516,N_17412,N_17039);
nand U18517 (N_18517,N_17504,N_17055);
and U18518 (N_18518,N_17578,N_17256);
nand U18519 (N_18519,N_17008,N_17077);
xor U18520 (N_18520,N_17982,N_17666);
nor U18521 (N_18521,N_17536,N_17192);
and U18522 (N_18522,N_17715,N_17980);
xnor U18523 (N_18523,N_17091,N_17862);
nor U18524 (N_18524,N_17609,N_17370);
or U18525 (N_18525,N_17519,N_17640);
and U18526 (N_18526,N_17224,N_17710);
and U18527 (N_18527,N_17931,N_17472);
nor U18528 (N_18528,N_17620,N_17524);
nand U18529 (N_18529,N_17604,N_17990);
nor U18530 (N_18530,N_17975,N_17377);
nor U18531 (N_18531,N_17343,N_17874);
and U18532 (N_18532,N_17455,N_17468);
or U18533 (N_18533,N_17773,N_17032);
nor U18534 (N_18534,N_17138,N_17939);
nand U18535 (N_18535,N_17540,N_17217);
or U18536 (N_18536,N_17215,N_17427);
and U18537 (N_18537,N_17469,N_17397);
or U18538 (N_18538,N_17785,N_17628);
nor U18539 (N_18539,N_17609,N_17904);
nor U18540 (N_18540,N_17029,N_17297);
or U18541 (N_18541,N_17341,N_17955);
nand U18542 (N_18542,N_17265,N_17693);
xnor U18543 (N_18543,N_17435,N_17977);
xor U18544 (N_18544,N_17714,N_17619);
xor U18545 (N_18545,N_17993,N_17089);
and U18546 (N_18546,N_17565,N_17058);
and U18547 (N_18547,N_17932,N_17127);
and U18548 (N_18548,N_17310,N_17421);
and U18549 (N_18549,N_17391,N_17712);
nand U18550 (N_18550,N_17695,N_17349);
or U18551 (N_18551,N_17446,N_17181);
xnor U18552 (N_18552,N_17316,N_17595);
nor U18553 (N_18553,N_17635,N_17201);
xnor U18554 (N_18554,N_17720,N_17590);
xnor U18555 (N_18555,N_17941,N_17076);
xnor U18556 (N_18556,N_17134,N_17885);
xnor U18557 (N_18557,N_17628,N_17517);
or U18558 (N_18558,N_17138,N_17558);
xor U18559 (N_18559,N_17245,N_17905);
nor U18560 (N_18560,N_17790,N_17056);
and U18561 (N_18561,N_17733,N_17764);
and U18562 (N_18562,N_17599,N_17962);
xnor U18563 (N_18563,N_17502,N_17651);
nor U18564 (N_18564,N_17614,N_17107);
nand U18565 (N_18565,N_17591,N_17058);
or U18566 (N_18566,N_17022,N_17087);
or U18567 (N_18567,N_17313,N_17104);
nor U18568 (N_18568,N_17273,N_17369);
or U18569 (N_18569,N_17513,N_17810);
xnor U18570 (N_18570,N_17908,N_17626);
and U18571 (N_18571,N_17198,N_17969);
xnor U18572 (N_18572,N_17120,N_17716);
xnor U18573 (N_18573,N_17746,N_17795);
and U18574 (N_18574,N_17840,N_17296);
or U18575 (N_18575,N_17759,N_17889);
nor U18576 (N_18576,N_17255,N_17025);
nor U18577 (N_18577,N_17541,N_17350);
nor U18578 (N_18578,N_17066,N_17285);
and U18579 (N_18579,N_17973,N_17652);
nor U18580 (N_18580,N_17103,N_17075);
nor U18581 (N_18581,N_17830,N_17530);
or U18582 (N_18582,N_17631,N_17526);
or U18583 (N_18583,N_17821,N_17917);
nor U18584 (N_18584,N_17036,N_17980);
or U18585 (N_18585,N_17008,N_17489);
nor U18586 (N_18586,N_17570,N_17980);
nand U18587 (N_18587,N_17852,N_17093);
or U18588 (N_18588,N_17968,N_17896);
and U18589 (N_18589,N_17748,N_17788);
nor U18590 (N_18590,N_17030,N_17057);
nand U18591 (N_18591,N_17823,N_17331);
or U18592 (N_18592,N_17360,N_17138);
xnor U18593 (N_18593,N_17791,N_17245);
nand U18594 (N_18594,N_17238,N_17064);
nor U18595 (N_18595,N_17719,N_17086);
or U18596 (N_18596,N_17247,N_17310);
and U18597 (N_18597,N_17257,N_17075);
xor U18598 (N_18598,N_17589,N_17088);
nor U18599 (N_18599,N_17172,N_17765);
or U18600 (N_18600,N_17096,N_17206);
and U18601 (N_18601,N_17249,N_17315);
nor U18602 (N_18602,N_17782,N_17437);
nand U18603 (N_18603,N_17626,N_17369);
nor U18604 (N_18604,N_17703,N_17973);
nor U18605 (N_18605,N_17094,N_17217);
nor U18606 (N_18606,N_17834,N_17330);
and U18607 (N_18607,N_17664,N_17962);
or U18608 (N_18608,N_17628,N_17542);
nor U18609 (N_18609,N_17921,N_17711);
nor U18610 (N_18610,N_17979,N_17134);
nor U18611 (N_18611,N_17702,N_17418);
xnor U18612 (N_18612,N_17360,N_17204);
and U18613 (N_18613,N_17125,N_17712);
nand U18614 (N_18614,N_17550,N_17069);
and U18615 (N_18615,N_17075,N_17280);
and U18616 (N_18616,N_17143,N_17281);
xnor U18617 (N_18617,N_17359,N_17155);
nor U18618 (N_18618,N_17335,N_17191);
xor U18619 (N_18619,N_17880,N_17506);
or U18620 (N_18620,N_17944,N_17935);
nor U18621 (N_18621,N_17896,N_17386);
xor U18622 (N_18622,N_17828,N_17258);
xnor U18623 (N_18623,N_17991,N_17204);
or U18624 (N_18624,N_17214,N_17779);
xor U18625 (N_18625,N_17261,N_17554);
and U18626 (N_18626,N_17533,N_17559);
and U18627 (N_18627,N_17477,N_17733);
xnor U18628 (N_18628,N_17959,N_17599);
nor U18629 (N_18629,N_17187,N_17491);
and U18630 (N_18630,N_17847,N_17916);
nand U18631 (N_18631,N_17038,N_17307);
nand U18632 (N_18632,N_17281,N_17039);
xnor U18633 (N_18633,N_17665,N_17621);
xnor U18634 (N_18634,N_17506,N_17505);
xnor U18635 (N_18635,N_17060,N_17545);
or U18636 (N_18636,N_17010,N_17225);
xnor U18637 (N_18637,N_17854,N_17932);
nand U18638 (N_18638,N_17496,N_17976);
xnor U18639 (N_18639,N_17679,N_17766);
nand U18640 (N_18640,N_17443,N_17829);
xnor U18641 (N_18641,N_17467,N_17679);
and U18642 (N_18642,N_17965,N_17106);
xnor U18643 (N_18643,N_17012,N_17488);
or U18644 (N_18644,N_17101,N_17914);
and U18645 (N_18645,N_17758,N_17544);
or U18646 (N_18646,N_17965,N_17095);
xor U18647 (N_18647,N_17171,N_17727);
xnor U18648 (N_18648,N_17596,N_17940);
xnor U18649 (N_18649,N_17103,N_17290);
xor U18650 (N_18650,N_17641,N_17103);
nor U18651 (N_18651,N_17821,N_17534);
nand U18652 (N_18652,N_17701,N_17079);
or U18653 (N_18653,N_17030,N_17570);
and U18654 (N_18654,N_17008,N_17472);
nand U18655 (N_18655,N_17635,N_17361);
nor U18656 (N_18656,N_17519,N_17615);
nand U18657 (N_18657,N_17275,N_17544);
nor U18658 (N_18658,N_17100,N_17539);
and U18659 (N_18659,N_17071,N_17329);
or U18660 (N_18660,N_17161,N_17513);
nor U18661 (N_18661,N_17561,N_17048);
nand U18662 (N_18662,N_17946,N_17854);
nor U18663 (N_18663,N_17936,N_17461);
nand U18664 (N_18664,N_17653,N_17563);
xor U18665 (N_18665,N_17056,N_17098);
xor U18666 (N_18666,N_17391,N_17925);
nor U18667 (N_18667,N_17523,N_17321);
and U18668 (N_18668,N_17136,N_17068);
or U18669 (N_18669,N_17187,N_17705);
or U18670 (N_18670,N_17960,N_17677);
or U18671 (N_18671,N_17631,N_17169);
or U18672 (N_18672,N_17613,N_17157);
nor U18673 (N_18673,N_17473,N_17354);
nand U18674 (N_18674,N_17128,N_17242);
or U18675 (N_18675,N_17512,N_17766);
xor U18676 (N_18676,N_17421,N_17262);
xnor U18677 (N_18677,N_17054,N_17429);
and U18678 (N_18678,N_17645,N_17260);
nand U18679 (N_18679,N_17852,N_17504);
or U18680 (N_18680,N_17149,N_17588);
or U18681 (N_18681,N_17195,N_17226);
xnor U18682 (N_18682,N_17882,N_17364);
nor U18683 (N_18683,N_17391,N_17663);
and U18684 (N_18684,N_17508,N_17327);
or U18685 (N_18685,N_17492,N_17252);
and U18686 (N_18686,N_17941,N_17837);
or U18687 (N_18687,N_17573,N_17474);
xnor U18688 (N_18688,N_17821,N_17467);
nand U18689 (N_18689,N_17759,N_17829);
nor U18690 (N_18690,N_17484,N_17047);
xor U18691 (N_18691,N_17930,N_17731);
nand U18692 (N_18692,N_17485,N_17959);
nand U18693 (N_18693,N_17563,N_17801);
nand U18694 (N_18694,N_17866,N_17547);
nor U18695 (N_18695,N_17193,N_17081);
nor U18696 (N_18696,N_17084,N_17297);
nand U18697 (N_18697,N_17920,N_17629);
and U18698 (N_18698,N_17196,N_17256);
xnor U18699 (N_18699,N_17460,N_17101);
and U18700 (N_18700,N_17045,N_17366);
nand U18701 (N_18701,N_17845,N_17474);
and U18702 (N_18702,N_17783,N_17975);
and U18703 (N_18703,N_17913,N_17410);
or U18704 (N_18704,N_17821,N_17721);
nand U18705 (N_18705,N_17765,N_17261);
nand U18706 (N_18706,N_17061,N_17820);
or U18707 (N_18707,N_17326,N_17874);
nand U18708 (N_18708,N_17475,N_17544);
nor U18709 (N_18709,N_17177,N_17838);
xnor U18710 (N_18710,N_17983,N_17883);
nor U18711 (N_18711,N_17041,N_17010);
nor U18712 (N_18712,N_17596,N_17179);
nor U18713 (N_18713,N_17636,N_17235);
nor U18714 (N_18714,N_17226,N_17559);
nand U18715 (N_18715,N_17992,N_17369);
xnor U18716 (N_18716,N_17208,N_17264);
xnor U18717 (N_18717,N_17958,N_17851);
nor U18718 (N_18718,N_17624,N_17830);
or U18719 (N_18719,N_17392,N_17202);
xnor U18720 (N_18720,N_17178,N_17047);
nor U18721 (N_18721,N_17584,N_17264);
or U18722 (N_18722,N_17538,N_17230);
nand U18723 (N_18723,N_17658,N_17551);
and U18724 (N_18724,N_17813,N_17534);
and U18725 (N_18725,N_17544,N_17185);
and U18726 (N_18726,N_17842,N_17481);
nand U18727 (N_18727,N_17678,N_17904);
and U18728 (N_18728,N_17967,N_17613);
nand U18729 (N_18729,N_17760,N_17719);
and U18730 (N_18730,N_17293,N_17623);
nor U18731 (N_18731,N_17270,N_17754);
xor U18732 (N_18732,N_17659,N_17428);
or U18733 (N_18733,N_17758,N_17984);
nand U18734 (N_18734,N_17634,N_17713);
or U18735 (N_18735,N_17450,N_17847);
nor U18736 (N_18736,N_17852,N_17265);
nor U18737 (N_18737,N_17014,N_17340);
and U18738 (N_18738,N_17937,N_17102);
nor U18739 (N_18739,N_17020,N_17665);
and U18740 (N_18740,N_17528,N_17920);
xor U18741 (N_18741,N_17146,N_17790);
and U18742 (N_18742,N_17011,N_17412);
and U18743 (N_18743,N_17797,N_17104);
nor U18744 (N_18744,N_17770,N_17877);
nand U18745 (N_18745,N_17789,N_17055);
xnor U18746 (N_18746,N_17008,N_17822);
or U18747 (N_18747,N_17998,N_17776);
nor U18748 (N_18748,N_17943,N_17662);
nor U18749 (N_18749,N_17224,N_17339);
and U18750 (N_18750,N_17104,N_17525);
xnor U18751 (N_18751,N_17550,N_17035);
and U18752 (N_18752,N_17519,N_17534);
nand U18753 (N_18753,N_17880,N_17720);
xor U18754 (N_18754,N_17972,N_17325);
or U18755 (N_18755,N_17385,N_17901);
and U18756 (N_18756,N_17363,N_17813);
or U18757 (N_18757,N_17948,N_17415);
or U18758 (N_18758,N_17045,N_17396);
xnor U18759 (N_18759,N_17969,N_17185);
nor U18760 (N_18760,N_17914,N_17872);
and U18761 (N_18761,N_17098,N_17496);
or U18762 (N_18762,N_17502,N_17655);
nand U18763 (N_18763,N_17761,N_17538);
nor U18764 (N_18764,N_17188,N_17101);
and U18765 (N_18765,N_17235,N_17001);
or U18766 (N_18766,N_17318,N_17253);
nand U18767 (N_18767,N_17018,N_17584);
and U18768 (N_18768,N_17645,N_17587);
nor U18769 (N_18769,N_17168,N_17600);
and U18770 (N_18770,N_17782,N_17460);
xor U18771 (N_18771,N_17121,N_17984);
or U18772 (N_18772,N_17654,N_17926);
nor U18773 (N_18773,N_17171,N_17542);
and U18774 (N_18774,N_17425,N_17492);
or U18775 (N_18775,N_17771,N_17549);
nor U18776 (N_18776,N_17048,N_17074);
and U18777 (N_18777,N_17121,N_17534);
xnor U18778 (N_18778,N_17911,N_17573);
and U18779 (N_18779,N_17272,N_17662);
nor U18780 (N_18780,N_17335,N_17673);
xnor U18781 (N_18781,N_17690,N_17529);
or U18782 (N_18782,N_17911,N_17305);
xor U18783 (N_18783,N_17934,N_17217);
nand U18784 (N_18784,N_17233,N_17623);
or U18785 (N_18785,N_17918,N_17380);
nand U18786 (N_18786,N_17996,N_17908);
nand U18787 (N_18787,N_17265,N_17510);
nor U18788 (N_18788,N_17234,N_17508);
nor U18789 (N_18789,N_17021,N_17396);
nor U18790 (N_18790,N_17540,N_17968);
and U18791 (N_18791,N_17445,N_17367);
nand U18792 (N_18792,N_17547,N_17452);
xor U18793 (N_18793,N_17858,N_17590);
nand U18794 (N_18794,N_17259,N_17752);
nor U18795 (N_18795,N_17391,N_17372);
or U18796 (N_18796,N_17984,N_17759);
nand U18797 (N_18797,N_17996,N_17825);
nand U18798 (N_18798,N_17812,N_17256);
or U18799 (N_18799,N_17225,N_17442);
nor U18800 (N_18800,N_17689,N_17073);
xnor U18801 (N_18801,N_17652,N_17793);
xor U18802 (N_18802,N_17433,N_17393);
xnor U18803 (N_18803,N_17574,N_17170);
xnor U18804 (N_18804,N_17824,N_17877);
nand U18805 (N_18805,N_17944,N_17249);
or U18806 (N_18806,N_17781,N_17510);
xnor U18807 (N_18807,N_17775,N_17636);
nor U18808 (N_18808,N_17468,N_17794);
xnor U18809 (N_18809,N_17683,N_17285);
nand U18810 (N_18810,N_17532,N_17321);
or U18811 (N_18811,N_17775,N_17960);
xor U18812 (N_18812,N_17121,N_17423);
nor U18813 (N_18813,N_17646,N_17677);
or U18814 (N_18814,N_17061,N_17912);
xnor U18815 (N_18815,N_17496,N_17790);
nand U18816 (N_18816,N_17984,N_17369);
nor U18817 (N_18817,N_17964,N_17646);
or U18818 (N_18818,N_17203,N_17176);
or U18819 (N_18819,N_17708,N_17881);
nand U18820 (N_18820,N_17631,N_17688);
nand U18821 (N_18821,N_17918,N_17542);
nor U18822 (N_18822,N_17484,N_17127);
xor U18823 (N_18823,N_17307,N_17249);
nand U18824 (N_18824,N_17895,N_17968);
nand U18825 (N_18825,N_17976,N_17464);
or U18826 (N_18826,N_17633,N_17797);
xor U18827 (N_18827,N_17287,N_17443);
nand U18828 (N_18828,N_17457,N_17796);
nor U18829 (N_18829,N_17996,N_17113);
nor U18830 (N_18830,N_17376,N_17307);
nor U18831 (N_18831,N_17224,N_17641);
and U18832 (N_18832,N_17491,N_17956);
xor U18833 (N_18833,N_17521,N_17698);
xor U18834 (N_18834,N_17296,N_17341);
or U18835 (N_18835,N_17069,N_17978);
xnor U18836 (N_18836,N_17207,N_17523);
xor U18837 (N_18837,N_17188,N_17005);
and U18838 (N_18838,N_17641,N_17884);
nor U18839 (N_18839,N_17758,N_17520);
or U18840 (N_18840,N_17788,N_17511);
and U18841 (N_18841,N_17314,N_17842);
xnor U18842 (N_18842,N_17654,N_17250);
xor U18843 (N_18843,N_17446,N_17911);
and U18844 (N_18844,N_17710,N_17919);
and U18845 (N_18845,N_17321,N_17850);
or U18846 (N_18846,N_17063,N_17385);
or U18847 (N_18847,N_17694,N_17722);
and U18848 (N_18848,N_17508,N_17966);
nor U18849 (N_18849,N_17548,N_17360);
or U18850 (N_18850,N_17538,N_17979);
xnor U18851 (N_18851,N_17073,N_17251);
and U18852 (N_18852,N_17767,N_17959);
and U18853 (N_18853,N_17542,N_17523);
and U18854 (N_18854,N_17735,N_17866);
and U18855 (N_18855,N_17378,N_17149);
or U18856 (N_18856,N_17598,N_17997);
and U18857 (N_18857,N_17689,N_17667);
nor U18858 (N_18858,N_17198,N_17822);
nand U18859 (N_18859,N_17907,N_17988);
and U18860 (N_18860,N_17760,N_17225);
and U18861 (N_18861,N_17368,N_17741);
nand U18862 (N_18862,N_17866,N_17929);
xor U18863 (N_18863,N_17186,N_17613);
or U18864 (N_18864,N_17374,N_17805);
nor U18865 (N_18865,N_17964,N_17575);
or U18866 (N_18866,N_17847,N_17954);
and U18867 (N_18867,N_17376,N_17270);
nand U18868 (N_18868,N_17388,N_17930);
nor U18869 (N_18869,N_17593,N_17039);
nor U18870 (N_18870,N_17814,N_17089);
nand U18871 (N_18871,N_17136,N_17307);
nand U18872 (N_18872,N_17597,N_17215);
or U18873 (N_18873,N_17088,N_17368);
or U18874 (N_18874,N_17645,N_17428);
xnor U18875 (N_18875,N_17607,N_17293);
and U18876 (N_18876,N_17090,N_17907);
or U18877 (N_18877,N_17990,N_17016);
and U18878 (N_18878,N_17815,N_17654);
and U18879 (N_18879,N_17637,N_17785);
nand U18880 (N_18880,N_17686,N_17554);
xnor U18881 (N_18881,N_17702,N_17826);
nand U18882 (N_18882,N_17044,N_17549);
or U18883 (N_18883,N_17061,N_17033);
or U18884 (N_18884,N_17081,N_17071);
or U18885 (N_18885,N_17444,N_17974);
nand U18886 (N_18886,N_17961,N_17040);
nor U18887 (N_18887,N_17994,N_17264);
xor U18888 (N_18888,N_17885,N_17363);
nor U18889 (N_18889,N_17738,N_17277);
nor U18890 (N_18890,N_17130,N_17930);
nand U18891 (N_18891,N_17102,N_17456);
and U18892 (N_18892,N_17194,N_17517);
or U18893 (N_18893,N_17132,N_17300);
or U18894 (N_18894,N_17411,N_17105);
and U18895 (N_18895,N_17081,N_17141);
nand U18896 (N_18896,N_17977,N_17664);
xnor U18897 (N_18897,N_17183,N_17588);
and U18898 (N_18898,N_17103,N_17956);
nor U18899 (N_18899,N_17915,N_17494);
nand U18900 (N_18900,N_17818,N_17148);
or U18901 (N_18901,N_17002,N_17773);
and U18902 (N_18902,N_17909,N_17580);
nor U18903 (N_18903,N_17707,N_17133);
and U18904 (N_18904,N_17154,N_17291);
nand U18905 (N_18905,N_17841,N_17048);
and U18906 (N_18906,N_17691,N_17785);
xnor U18907 (N_18907,N_17116,N_17863);
or U18908 (N_18908,N_17848,N_17223);
and U18909 (N_18909,N_17403,N_17418);
or U18910 (N_18910,N_17105,N_17833);
or U18911 (N_18911,N_17618,N_17417);
or U18912 (N_18912,N_17827,N_17577);
nand U18913 (N_18913,N_17003,N_17002);
nand U18914 (N_18914,N_17757,N_17372);
nor U18915 (N_18915,N_17588,N_17322);
and U18916 (N_18916,N_17999,N_17651);
nor U18917 (N_18917,N_17859,N_17341);
nor U18918 (N_18918,N_17154,N_17748);
nor U18919 (N_18919,N_17374,N_17796);
and U18920 (N_18920,N_17606,N_17728);
xnor U18921 (N_18921,N_17947,N_17245);
nand U18922 (N_18922,N_17338,N_17553);
xnor U18923 (N_18923,N_17144,N_17544);
and U18924 (N_18924,N_17348,N_17665);
and U18925 (N_18925,N_17977,N_17667);
or U18926 (N_18926,N_17298,N_17528);
and U18927 (N_18927,N_17568,N_17223);
nand U18928 (N_18928,N_17326,N_17672);
or U18929 (N_18929,N_17491,N_17384);
nand U18930 (N_18930,N_17379,N_17082);
and U18931 (N_18931,N_17442,N_17894);
xnor U18932 (N_18932,N_17463,N_17754);
nor U18933 (N_18933,N_17598,N_17041);
nor U18934 (N_18934,N_17679,N_17233);
xnor U18935 (N_18935,N_17672,N_17598);
nor U18936 (N_18936,N_17222,N_17737);
nor U18937 (N_18937,N_17457,N_17800);
xor U18938 (N_18938,N_17395,N_17174);
or U18939 (N_18939,N_17231,N_17027);
nand U18940 (N_18940,N_17007,N_17672);
nor U18941 (N_18941,N_17201,N_17626);
nor U18942 (N_18942,N_17059,N_17568);
nand U18943 (N_18943,N_17116,N_17738);
nand U18944 (N_18944,N_17973,N_17664);
xnor U18945 (N_18945,N_17281,N_17958);
and U18946 (N_18946,N_17446,N_17257);
xor U18947 (N_18947,N_17544,N_17695);
nand U18948 (N_18948,N_17429,N_17986);
nand U18949 (N_18949,N_17100,N_17948);
nand U18950 (N_18950,N_17958,N_17187);
xnor U18951 (N_18951,N_17368,N_17445);
nand U18952 (N_18952,N_17976,N_17963);
and U18953 (N_18953,N_17128,N_17501);
nand U18954 (N_18954,N_17358,N_17875);
nand U18955 (N_18955,N_17801,N_17562);
nor U18956 (N_18956,N_17515,N_17350);
or U18957 (N_18957,N_17640,N_17314);
and U18958 (N_18958,N_17687,N_17761);
nor U18959 (N_18959,N_17938,N_17540);
nor U18960 (N_18960,N_17526,N_17820);
nand U18961 (N_18961,N_17088,N_17837);
or U18962 (N_18962,N_17754,N_17863);
nor U18963 (N_18963,N_17971,N_17317);
or U18964 (N_18964,N_17003,N_17677);
and U18965 (N_18965,N_17645,N_17340);
and U18966 (N_18966,N_17212,N_17728);
or U18967 (N_18967,N_17781,N_17680);
xnor U18968 (N_18968,N_17696,N_17262);
nand U18969 (N_18969,N_17643,N_17386);
nor U18970 (N_18970,N_17024,N_17780);
and U18971 (N_18971,N_17827,N_17077);
nand U18972 (N_18972,N_17994,N_17900);
and U18973 (N_18973,N_17060,N_17852);
or U18974 (N_18974,N_17095,N_17368);
and U18975 (N_18975,N_17179,N_17225);
nand U18976 (N_18976,N_17099,N_17543);
xor U18977 (N_18977,N_17853,N_17661);
xor U18978 (N_18978,N_17399,N_17127);
or U18979 (N_18979,N_17581,N_17430);
and U18980 (N_18980,N_17207,N_17627);
nand U18981 (N_18981,N_17149,N_17324);
xnor U18982 (N_18982,N_17910,N_17297);
nand U18983 (N_18983,N_17807,N_17952);
nor U18984 (N_18984,N_17825,N_17576);
xor U18985 (N_18985,N_17340,N_17252);
nand U18986 (N_18986,N_17401,N_17650);
nand U18987 (N_18987,N_17978,N_17944);
nor U18988 (N_18988,N_17500,N_17098);
nand U18989 (N_18989,N_17140,N_17516);
xor U18990 (N_18990,N_17385,N_17190);
nand U18991 (N_18991,N_17347,N_17061);
and U18992 (N_18992,N_17453,N_17845);
and U18993 (N_18993,N_17824,N_17764);
nor U18994 (N_18994,N_17185,N_17639);
nand U18995 (N_18995,N_17661,N_17226);
and U18996 (N_18996,N_17071,N_17037);
xnor U18997 (N_18997,N_17078,N_17941);
nand U18998 (N_18998,N_17897,N_17173);
nand U18999 (N_18999,N_17057,N_17314);
xor U19000 (N_19000,N_18976,N_18582);
or U19001 (N_19001,N_18862,N_18206);
xor U19002 (N_19002,N_18097,N_18864);
nand U19003 (N_19003,N_18617,N_18535);
and U19004 (N_19004,N_18526,N_18095);
xnor U19005 (N_19005,N_18106,N_18392);
nor U19006 (N_19006,N_18844,N_18857);
nor U19007 (N_19007,N_18419,N_18974);
nand U19008 (N_19008,N_18902,N_18280);
nand U19009 (N_19009,N_18541,N_18145);
xor U19010 (N_19010,N_18602,N_18113);
and U19011 (N_19011,N_18321,N_18143);
nand U19012 (N_19012,N_18286,N_18613);
or U19013 (N_19013,N_18805,N_18637);
nor U19014 (N_19014,N_18929,N_18252);
and U19015 (N_19015,N_18247,N_18311);
nor U19016 (N_19016,N_18620,N_18749);
or U19017 (N_19017,N_18720,N_18624);
xnor U19018 (N_19018,N_18626,N_18779);
xnor U19019 (N_19019,N_18343,N_18552);
and U19020 (N_19020,N_18580,N_18411);
xnor U19021 (N_19021,N_18363,N_18813);
nand U19022 (N_19022,N_18258,N_18500);
xor U19023 (N_19023,N_18746,N_18763);
nor U19024 (N_19024,N_18506,N_18998);
nand U19025 (N_19025,N_18354,N_18731);
xnor U19026 (N_19026,N_18405,N_18319);
nand U19027 (N_19027,N_18249,N_18315);
or U19028 (N_19028,N_18532,N_18041);
nor U19029 (N_19029,N_18547,N_18255);
nor U19030 (N_19030,N_18140,N_18835);
and U19031 (N_19031,N_18949,N_18752);
xnor U19032 (N_19032,N_18911,N_18519);
nand U19033 (N_19033,N_18841,N_18825);
or U19034 (N_19034,N_18555,N_18717);
or U19035 (N_19035,N_18858,N_18655);
and U19036 (N_19036,N_18129,N_18478);
or U19037 (N_19037,N_18899,N_18110);
nor U19038 (N_19038,N_18175,N_18663);
nand U19039 (N_19039,N_18509,N_18855);
nand U19040 (N_19040,N_18473,N_18971);
or U19041 (N_19041,N_18156,N_18131);
nor U19042 (N_19042,N_18339,N_18525);
and U19043 (N_19043,N_18186,N_18107);
and U19044 (N_19044,N_18390,N_18067);
nor U19045 (N_19045,N_18462,N_18385);
or U19046 (N_19046,N_18963,N_18409);
or U19047 (N_19047,N_18927,N_18226);
and U19048 (N_19048,N_18705,N_18893);
and U19049 (N_19049,N_18061,N_18096);
nor U19050 (N_19050,N_18292,N_18799);
xnor U19051 (N_19051,N_18260,N_18290);
nand U19052 (N_19052,N_18202,N_18170);
nand U19053 (N_19053,N_18730,N_18220);
xnor U19054 (N_19054,N_18634,N_18843);
and U19055 (N_19055,N_18695,N_18660);
nor U19056 (N_19056,N_18433,N_18601);
or U19057 (N_19057,N_18570,N_18324);
nor U19058 (N_19058,N_18860,N_18036);
nand U19059 (N_19059,N_18137,N_18646);
or U19060 (N_19060,N_18169,N_18447);
nand U19061 (N_19061,N_18494,N_18584);
and U19062 (N_19062,N_18012,N_18573);
xor U19063 (N_19063,N_18149,N_18374);
nand U19064 (N_19064,N_18213,N_18699);
nor U19065 (N_19065,N_18788,N_18415);
xor U19066 (N_19066,N_18228,N_18874);
and U19067 (N_19067,N_18033,N_18125);
or U19068 (N_19068,N_18444,N_18314);
xnor U19069 (N_19069,N_18987,N_18100);
or U19070 (N_19070,N_18135,N_18649);
or U19071 (N_19071,N_18567,N_18109);
or U19072 (N_19072,N_18598,N_18372);
xor U19073 (N_19073,N_18597,N_18402);
nand U19074 (N_19074,N_18267,N_18901);
nand U19075 (N_19075,N_18189,N_18091);
nor U19076 (N_19076,N_18338,N_18043);
and U19077 (N_19077,N_18785,N_18001);
xnor U19078 (N_19078,N_18890,N_18839);
and U19079 (N_19079,N_18116,N_18854);
xor U19080 (N_19080,N_18394,N_18120);
xnor U19081 (N_19081,N_18913,N_18956);
and U19082 (N_19082,N_18069,N_18472);
nor U19083 (N_19083,N_18393,N_18397);
nor U19084 (N_19084,N_18968,N_18279);
or U19085 (N_19085,N_18115,N_18691);
nor U19086 (N_19086,N_18632,N_18052);
nor U19087 (N_19087,N_18177,N_18966);
or U19088 (N_19088,N_18119,N_18686);
xor U19089 (N_19089,N_18105,N_18128);
nand U19090 (N_19090,N_18797,N_18721);
nand U19091 (N_19091,N_18875,N_18905);
nand U19092 (N_19092,N_18004,N_18300);
and U19093 (N_19093,N_18511,N_18009);
nand U19094 (N_19094,N_18231,N_18693);
or U19095 (N_19095,N_18030,N_18370);
or U19096 (N_19096,N_18098,N_18235);
or U19097 (N_19097,N_18350,N_18992);
xnor U19098 (N_19098,N_18938,N_18867);
nor U19099 (N_19099,N_18356,N_18952);
and U19100 (N_19100,N_18062,N_18815);
or U19101 (N_19101,N_18625,N_18099);
xnor U19102 (N_19102,N_18700,N_18973);
nand U19103 (N_19103,N_18571,N_18709);
xnor U19104 (N_19104,N_18185,N_18631);
xor U19105 (N_19105,N_18895,N_18421);
xnor U19106 (N_19106,N_18248,N_18869);
nor U19107 (N_19107,N_18513,N_18310);
nor U19108 (N_19108,N_18190,N_18437);
nor U19109 (N_19109,N_18694,N_18171);
and U19110 (N_19110,N_18262,N_18092);
xor U19111 (N_19111,N_18124,N_18726);
nor U19112 (N_19112,N_18743,N_18126);
or U19113 (N_19113,N_18502,N_18521);
nand U19114 (N_19114,N_18104,N_18331);
nand U19115 (N_19115,N_18450,N_18272);
and U19116 (N_19116,N_18318,N_18484);
nor U19117 (N_19117,N_18636,N_18460);
nand U19118 (N_19118,N_18467,N_18810);
or U19119 (N_19119,N_18309,N_18147);
nor U19120 (N_19120,N_18764,N_18191);
nor U19121 (N_19121,N_18997,N_18496);
nand U19122 (N_19122,N_18876,N_18208);
and U19123 (N_19123,N_18819,N_18919);
or U19124 (N_19124,N_18470,N_18600);
xor U19125 (N_19125,N_18389,N_18751);
nor U19126 (N_19126,N_18789,N_18492);
nor U19127 (N_19127,N_18403,N_18776);
or U19128 (N_19128,N_18616,N_18572);
or U19129 (N_19129,N_18714,N_18712);
nand U19130 (N_19130,N_18281,N_18887);
or U19131 (N_19131,N_18475,N_18682);
or U19132 (N_19132,N_18975,N_18576);
xnor U19133 (N_19133,N_18837,N_18935);
or U19134 (N_19134,N_18622,N_18355);
nor U19135 (N_19135,N_18423,N_18607);
nand U19136 (N_19136,N_18044,N_18882);
or U19137 (N_19137,N_18594,N_18733);
nand U19138 (N_19138,N_18505,N_18930);
xor U19139 (N_19139,N_18988,N_18545);
nor U19140 (N_19140,N_18851,N_18692);
xor U19141 (N_19141,N_18736,N_18045);
xor U19142 (N_19142,N_18474,N_18289);
and U19143 (N_19143,N_18690,N_18954);
or U19144 (N_19144,N_18561,N_18564);
nand U19145 (N_19145,N_18828,N_18793);
xnor U19146 (N_19146,N_18359,N_18674);
nand U19147 (N_19147,N_18653,N_18102);
or U19148 (N_19148,N_18408,N_18948);
xnor U19149 (N_19149,N_18083,N_18273);
xor U19150 (N_19150,N_18641,N_18336);
xor U19151 (N_19151,N_18227,N_18603);
nor U19152 (N_19152,N_18643,N_18141);
or U19153 (N_19153,N_18656,N_18784);
and U19154 (N_19154,N_18464,N_18765);
nor U19155 (N_19155,N_18728,N_18836);
nor U19156 (N_19156,N_18215,N_18969);
nand U19157 (N_19157,N_18063,N_18961);
nor U19158 (N_19158,N_18775,N_18629);
and U19159 (N_19159,N_18565,N_18586);
nor U19160 (N_19160,N_18546,N_18017);
nand U19161 (N_19161,N_18885,N_18676);
nand U19162 (N_19162,N_18136,N_18387);
xnor U19163 (N_19163,N_18592,N_18880);
nor U19164 (N_19164,N_18823,N_18933);
xnor U19165 (N_19165,N_18516,N_18926);
and U19166 (N_19166,N_18027,N_18884);
nor U19167 (N_19167,N_18970,N_18678);
or U19168 (N_19168,N_18647,N_18853);
and U19169 (N_19169,N_18654,N_18243);
xor U19170 (N_19170,N_18605,N_18293);
or U19171 (N_19171,N_18153,N_18003);
nor U19172 (N_19172,N_18233,N_18924);
nor U19173 (N_19173,N_18361,N_18900);
and U19174 (N_19174,N_18307,N_18439);
or U19175 (N_19175,N_18589,N_18777);
nor U19176 (N_19176,N_18955,N_18544);
nand U19177 (N_19177,N_18639,N_18368);
nor U19178 (N_19178,N_18889,N_18781);
nand U19179 (N_19179,N_18298,N_18416);
nor U19180 (N_19180,N_18357,N_18740);
nand U19181 (N_19181,N_18005,N_18630);
xnor U19182 (N_19182,N_18168,N_18514);
xor U19183 (N_19183,N_18266,N_18121);
nor U19184 (N_19184,N_18652,N_18308);
nor U19185 (N_19185,N_18209,N_18224);
or U19186 (N_19186,N_18058,N_18000);
or U19187 (N_19187,N_18146,N_18367);
or U19188 (N_19188,N_18928,N_18078);
and U19189 (N_19189,N_18093,N_18945);
or U19190 (N_19190,N_18379,N_18008);
nor U19191 (N_19191,N_18218,N_18082);
xnor U19192 (N_19192,N_18342,N_18047);
and U19193 (N_19193,N_18123,N_18039);
nand U19194 (N_19194,N_18959,N_18211);
xnor U19195 (N_19195,N_18380,N_18440);
nand U19196 (N_19196,N_18822,N_18879);
or U19197 (N_19197,N_18477,N_18804);
or U19198 (N_19198,N_18811,N_18877);
or U19199 (N_19199,N_18406,N_18790);
nor U19200 (N_19200,N_18801,N_18967);
nand U19201 (N_19201,N_18050,N_18701);
nor U19202 (N_19202,N_18878,N_18989);
nor U19203 (N_19203,N_18865,N_18329);
and U19204 (N_19204,N_18127,N_18520);
xor U19205 (N_19205,N_18739,N_18303);
xor U19206 (N_19206,N_18486,N_18794);
or U19207 (N_19207,N_18084,N_18427);
nand U19208 (N_19208,N_18378,N_18197);
xor U19209 (N_19209,N_18590,N_18627);
or U19210 (N_19210,N_18537,N_18246);
nand U19211 (N_19211,N_18184,N_18196);
nor U19212 (N_19212,N_18724,N_18138);
xor U19213 (N_19213,N_18734,N_18671);
nor U19214 (N_19214,N_18432,N_18452);
xor U19215 (N_19215,N_18435,N_18103);
or U19216 (N_19216,N_18783,N_18090);
or U19217 (N_19217,N_18426,N_18194);
nand U19218 (N_19218,N_18480,N_18362);
nand U19219 (N_19219,N_18217,N_18471);
xor U19220 (N_19220,N_18337,N_18834);
nor U19221 (N_19221,N_18562,N_18294);
nor U19222 (N_19222,N_18604,N_18375);
and U19223 (N_19223,N_18264,N_18278);
nand U19224 (N_19224,N_18330,N_18181);
nor U19225 (N_19225,N_18263,N_18301);
xnor U19226 (N_19226,N_18302,N_18530);
nor U19227 (N_19227,N_18787,N_18838);
and U19228 (N_19228,N_18468,N_18942);
or U19229 (N_19229,N_18953,N_18325);
or U19230 (N_19230,N_18863,N_18936);
xor U19231 (N_19231,N_18587,N_18167);
xnor U19232 (N_19232,N_18048,N_18088);
and U19233 (N_19233,N_18850,N_18680);
nor U19234 (N_19234,N_18434,N_18774);
xnor U19235 (N_19235,N_18398,N_18487);
or U19236 (N_19236,N_18495,N_18019);
nand U19237 (N_19237,N_18883,N_18606);
xnor U19238 (N_19238,N_18072,N_18698);
nor U19239 (N_19239,N_18897,N_18556);
nand U19240 (N_19240,N_18188,N_18738);
nor U19241 (N_19241,N_18316,N_18931);
or U19242 (N_19242,N_18922,N_18595);
nand U19243 (N_19243,N_18812,N_18888);
nand U19244 (N_19244,N_18445,N_18619);
and U19245 (N_19245,N_18577,N_18304);
nor U19246 (N_19246,N_18575,N_18507);
and U19247 (N_19247,N_18010,N_18234);
nand U19248 (N_19248,N_18485,N_18917);
and U19249 (N_19249,N_18960,N_18055);
nor U19250 (N_19250,N_18896,N_18972);
xnor U19251 (N_19251,N_18287,N_18327);
nand U19252 (N_19252,N_18192,N_18847);
or U19253 (N_19253,N_18497,N_18079);
and U19254 (N_19254,N_18569,N_18754);
nand U19255 (N_19255,N_18621,N_18579);
nand U19256 (N_19256,N_18087,N_18707);
and U19257 (N_19257,N_18463,N_18642);
and U19258 (N_19258,N_18396,N_18716);
or U19259 (N_19259,N_18111,N_18727);
or U19260 (N_19260,N_18182,N_18101);
nor U19261 (N_19261,N_18094,N_18907);
nand U19262 (N_19262,N_18710,N_18157);
or U19263 (N_19263,N_18207,N_18759);
nand U19264 (N_19264,N_18683,N_18456);
or U19265 (N_19265,N_18829,N_18719);
and U19266 (N_19266,N_18664,N_18032);
and U19267 (N_19267,N_18689,N_18257);
nor U19268 (N_19268,N_18984,N_18348);
xnor U19269 (N_19269,N_18221,N_18915);
nor U19270 (N_19270,N_18214,N_18501);
nor U19271 (N_19271,N_18852,N_18941);
nor U19272 (N_19272,N_18773,N_18762);
nor U19273 (N_19273,N_18122,N_18152);
or U19274 (N_19274,N_18065,N_18977);
and U19275 (N_19275,N_18200,N_18155);
nor U19276 (N_19276,N_18769,N_18995);
nand U19277 (N_19277,N_18623,N_18659);
xor U19278 (N_19278,N_18291,N_18665);
nor U19279 (N_19279,N_18566,N_18791);
nor U19280 (N_19280,N_18198,N_18628);
and U19281 (N_19281,N_18934,N_18112);
or U19282 (N_19282,N_18585,N_18947);
nand U19283 (N_19283,N_18524,N_18022);
xor U19284 (N_19284,N_18780,N_18269);
and U19285 (N_19285,N_18792,N_18557);
xnor U19286 (N_19286,N_18183,N_18282);
nor U19287 (N_19287,N_18018,N_18908);
xnor U19288 (N_19288,N_18817,N_18089);
xor U19289 (N_19289,N_18178,N_18503);
and U19290 (N_19290,N_18295,N_18640);
and U19291 (N_19291,N_18904,N_18542);
xnor U19292 (N_19292,N_18508,N_18981);
nor U19293 (N_19293,N_18076,N_18075);
or U19294 (N_19294,N_18238,N_18469);
nor U19295 (N_19295,N_18158,N_18334);
nor U19296 (N_19296,N_18846,N_18187);
and U19297 (N_19297,N_18558,N_18428);
or U19298 (N_19298,N_18024,N_18236);
nand U19299 (N_19299,N_18015,N_18554);
nor U19300 (N_19300,N_18457,N_18230);
nand U19301 (N_19301,N_18453,N_18476);
nor U19302 (N_19302,N_18800,N_18870);
nand U19303 (N_19303,N_18560,N_18268);
and U19304 (N_19304,N_18943,N_18725);
xor U19305 (N_19305,N_18245,N_18451);
or U19306 (N_19306,N_18056,N_18299);
or U19307 (N_19307,N_18199,N_18261);
nand U19308 (N_19308,N_18679,N_18028);
nand U19309 (N_19309,N_18222,N_18772);
or U19310 (N_19310,N_18459,N_18735);
or U19311 (N_19311,N_18814,N_18771);
xor U19312 (N_19312,N_18872,N_18068);
and U19313 (N_19313,N_18894,N_18162);
xnor U19314 (N_19314,N_18991,N_18400);
nand U19315 (N_19315,N_18054,N_18768);
or U19316 (N_19316,N_18333,N_18448);
nor U19317 (N_19317,N_18824,N_18986);
and U19318 (N_19318,N_18553,N_18254);
or U19319 (N_19319,N_18244,N_18993);
and U19320 (N_19320,N_18618,N_18395);
nand U19321 (N_19321,N_18670,N_18490);
or U19322 (N_19322,N_18430,N_18358);
nand U19323 (N_19323,N_18596,N_18909);
nor U19324 (N_19324,N_18353,N_18212);
and U19325 (N_19325,N_18650,N_18609);
xor U19326 (N_19326,N_18133,N_18668);
nand U19327 (N_19327,N_18550,N_18482);
or U19328 (N_19328,N_18729,N_18528);
or U19329 (N_19329,N_18704,N_18351);
nand U19330 (N_19330,N_18081,N_18431);
xor U19331 (N_19331,N_18479,N_18070);
or U19332 (N_19332,N_18842,N_18615);
nand U19333 (N_19333,N_18944,N_18349);
nand U19334 (N_19334,N_18667,N_18386);
nand U19335 (N_19335,N_18366,N_18504);
nand U19336 (N_19336,N_18536,N_18071);
nand U19337 (N_19337,N_18270,N_18982);
nor U19338 (N_19338,N_18345,N_18795);
and U19339 (N_19339,N_18910,N_18438);
and U19340 (N_19340,N_18436,N_18612);
nand U19341 (N_19341,N_18023,N_18407);
and U19342 (N_19342,N_18687,N_18173);
and U19343 (N_19343,N_18770,N_18950);
or U19344 (N_19344,N_18742,N_18335);
and U19345 (N_19345,N_18250,N_18745);
nand U19346 (N_19346,N_18086,N_18161);
or U19347 (N_19347,N_18831,N_18648);
or U19348 (N_19348,N_18006,N_18306);
nor U19349 (N_19349,N_18049,N_18253);
nor U19350 (N_19350,N_18996,N_18946);
nor U19351 (N_19351,N_18886,N_18697);
nand U19352 (N_19352,N_18757,N_18821);
xor U19353 (N_19353,N_18713,N_18688);
or U19354 (N_19354,N_18593,N_18673);
nand U19355 (N_19355,N_18527,N_18417);
nor U19356 (N_19356,N_18978,N_18046);
xor U19357 (N_19357,N_18059,N_18251);
nor U19358 (N_19358,N_18684,N_18174);
nand U19359 (N_19359,N_18446,N_18538);
nand U19360 (N_19360,N_18401,N_18994);
xor U19361 (N_19361,N_18715,N_18237);
nor U19362 (N_19362,N_18515,N_18702);
nor U19363 (N_19363,N_18591,N_18581);
xnor U19364 (N_19364,N_18165,N_18499);
nor U19365 (N_19365,N_18332,N_18510);
nand U19366 (N_19366,N_18718,N_18798);
xnor U19367 (N_19367,N_18493,N_18574);
xnor U19368 (N_19368,N_18965,N_18549);
or U19369 (N_19369,N_18455,N_18611);
or U19370 (N_19370,N_18999,N_18951);
or U19371 (N_19371,N_18563,N_18533);
or U19372 (N_19372,N_18203,N_18830);
nor U19373 (N_19373,N_18035,N_18013);
or U19374 (N_19374,N_18703,N_18489);
and U19375 (N_19375,N_18465,N_18412);
and U19376 (N_19376,N_18259,N_18559);
or U19377 (N_19377,N_18816,N_18285);
nor U19378 (N_19378,N_18920,N_18675);
xnor U19379 (N_19379,N_18179,N_18661);
nor U19380 (N_19380,N_18551,N_18866);
or U19381 (N_19381,N_18283,N_18364);
nor U19382 (N_19382,N_18413,N_18381);
or U19383 (N_19383,N_18371,N_18229);
nor U19384 (N_19384,N_18645,N_18741);
nor U19385 (N_19385,N_18818,N_18180);
or U19386 (N_19386,N_18488,N_18614);
xor U19387 (N_19387,N_18352,N_18539);
nand U19388 (N_19388,N_18205,N_18962);
nor U19389 (N_19389,N_18808,N_18420);
and U19390 (N_19390,N_18414,N_18384);
or U19391 (N_19391,N_18025,N_18681);
nor U19392 (N_19392,N_18132,N_18038);
nand U19393 (N_19393,N_18782,N_18377);
nor U19394 (N_19394,N_18014,N_18861);
or U19395 (N_19395,N_18114,N_18164);
or U19396 (N_19396,N_18980,N_18964);
or U19397 (N_19397,N_18912,N_18376);
xnor U19398 (N_19398,N_18424,N_18449);
nor U19399 (N_19399,N_18937,N_18983);
or U19400 (N_19400,N_18166,N_18297);
xnor U19401 (N_19401,N_18873,N_18906);
or U19402 (N_19402,N_18365,N_18466);
nor U19403 (N_19403,N_18066,N_18442);
nand U19404 (N_19404,N_18328,N_18429);
nand U19405 (N_19405,N_18060,N_18568);
nor U19406 (N_19406,N_18176,N_18708);
or U19407 (N_19407,N_18940,N_18341);
nor U19408 (N_19408,N_18748,N_18296);
nand U19409 (N_19409,N_18903,N_18921);
and U19410 (N_19410,N_18031,N_18523);
xor U19411 (N_19411,N_18677,N_18802);
nor U19412 (N_19412,N_18323,N_18118);
nand U19413 (N_19413,N_18806,N_18662);
or U19414 (N_19414,N_18150,N_18284);
nor U19415 (N_19415,N_18441,N_18848);
nor U19416 (N_19416,N_18481,N_18305);
and U19417 (N_19417,N_18633,N_18193);
xor U19418 (N_19418,N_18312,N_18277);
nor U19419 (N_19419,N_18756,N_18638);
nor U19420 (N_19420,N_18871,N_18347);
nand U19421 (N_19421,N_18074,N_18275);
xnor U19422 (N_19422,N_18422,N_18753);
xnor U19423 (N_19423,N_18957,N_18021);
nor U19424 (N_19424,N_18077,N_18522);
and U19425 (N_19425,N_18159,N_18340);
and U19426 (N_19426,N_18750,N_18239);
nor U19427 (N_19427,N_18760,N_18914);
or U19428 (N_19428,N_18242,N_18932);
nor U19429 (N_19429,N_18142,N_18425);
xor U19430 (N_19430,N_18744,N_18651);
nor U19431 (N_19431,N_18461,N_18761);
xnor U19432 (N_19432,N_18820,N_18256);
and U19433 (N_19433,N_18531,N_18344);
and U19434 (N_19434,N_18240,N_18073);
nand U19435 (N_19435,N_18918,N_18383);
and U19436 (N_19436,N_18672,N_18360);
nor U19437 (N_19437,N_18807,N_18758);
or U19438 (N_19438,N_18737,N_18037);
or U19439 (N_19439,N_18599,N_18322);
nor U19440 (N_19440,N_18856,N_18985);
xor U19441 (N_19441,N_18410,N_18160);
nand U19442 (N_19442,N_18543,N_18454);
and U19443 (N_19443,N_18723,N_18517);
or U19444 (N_19444,N_18979,N_18276);
xnor U19445 (N_19445,N_18418,N_18534);
and U19446 (N_19446,N_18134,N_18313);
xor U19447 (N_19447,N_18232,N_18064);
xnor U19448 (N_19448,N_18382,N_18766);
xnor U19449 (N_19449,N_18404,N_18053);
nand U19450 (N_19450,N_18939,N_18809);
nor U19451 (N_19451,N_18271,N_18139);
or U19452 (N_19452,N_18388,N_18151);
and U19453 (N_19453,N_18840,N_18990);
and U19454 (N_19454,N_18498,N_18320);
nor U19455 (N_19455,N_18706,N_18610);
nor U19456 (N_19456,N_18891,N_18029);
nor U19457 (N_19457,N_18210,N_18826);
or U19458 (N_19458,N_18223,N_18925);
xor U19459 (N_19459,N_18608,N_18849);
or U19460 (N_19460,N_18042,N_18767);
xor U19461 (N_19461,N_18051,N_18898);
xor U19462 (N_19462,N_18747,N_18148);
or U19463 (N_19463,N_18443,N_18172);
xnor U19464 (N_19464,N_18881,N_18108);
nand U19465 (N_19465,N_18786,N_18512);
or U19466 (N_19466,N_18666,N_18644);
nor U19467 (N_19467,N_18007,N_18016);
nand U19468 (N_19468,N_18635,N_18732);
and U19469 (N_19469,N_18669,N_18483);
nor U19470 (N_19470,N_18578,N_18288);
or U19471 (N_19471,N_18326,N_18274);
or U19472 (N_19472,N_18588,N_18225);
xor U19473 (N_19473,N_18216,N_18892);
xnor U19474 (N_19474,N_18696,N_18369);
xor U19475 (N_19475,N_18399,N_18057);
xor U19476 (N_19476,N_18144,N_18845);
nand U19477 (N_19477,N_18391,N_18832);
nand U19478 (N_19478,N_18491,N_18657);
and U19479 (N_19479,N_18011,N_18346);
xor U19480 (N_19480,N_18540,N_18458);
nor U19481 (N_19481,N_18026,N_18833);
nand U19482 (N_19482,N_18548,N_18916);
nor U19483 (N_19483,N_18529,N_18265);
nand U19484 (N_19484,N_18085,N_18117);
or U19485 (N_19485,N_18923,N_18317);
nand U19486 (N_19486,N_18020,N_18827);
nor U19487 (N_19487,N_18868,N_18201);
xor U19488 (N_19488,N_18711,N_18778);
nand U19489 (N_19489,N_18219,N_18130);
nor U19490 (N_19490,N_18080,N_18034);
or U19491 (N_19491,N_18958,N_18373);
nor U19492 (N_19492,N_18002,N_18040);
nor U19493 (N_19493,N_18685,N_18154);
and U19494 (N_19494,N_18583,N_18195);
xnor U19495 (N_19495,N_18796,N_18859);
and U19496 (N_19496,N_18755,N_18204);
xor U19497 (N_19497,N_18241,N_18803);
or U19498 (N_19498,N_18722,N_18163);
nand U19499 (N_19499,N_18518,N_18658);
xor U19500 (N_19500,N_18970,N_18554);
and U19501 (N_19501,N_18490,N_18351);
nor U19502 (N_19502,N_18088,N_18008);
or U19503 (N_19503,N_18716,N_18585);
nor U19504 (N_19504,N_18715,N_18393);
or U19505 (N_19505,N_18399,N_18241);
and U19506 (N_19506,N_18468,N_18465);
or U19507 (N_19507,N_18247,N_18315);
or U19508 (N_19508,N_18772,N_18630);
and U19509 (N_19509,N_18183,N_18109);
nor U19510 (N_19510,N_18262,N_18727);
or U19511 (N_19511,N_18803,N_18009);
xnor U19512 (N_19512,N_18681,N_18805);
or U19513 (N_19513,N_18075,N_18352);
nand U19514 (N_19514,N_18179,N_18247);
nand U19515 (N_19515,N_18784,N_18866);
xnor U19516 (N_19516,N_18203,N_18994);
or U19517 (N_19517,N_18927,N_18934);
and U19518 (N_19518,N_18140,N_18453);
and U19519 (N_19519,N_18382,N_18779);
and U19520 (N_19520,N_18340,N_18945);
xor U19521 (N_19521,N_18915,N_18689);
nor U19522 (N_19522,N_18363,N_18140);
nand U19523 (N_19523,N_18294,N_18305);
or U19524 (N_19524,N_18737,N_18203);
and U19525 (N_19525,N_18298,N_18181);
xnor U19526 (N_19526,N_18939,N_18309);
nand U19527 (N_19527,N_18368,N_18464);
nand U19528 (N_19528,N_18659,N_18206);
and U19529 (N_19529,N_18110,N_18054);
xor U19530 (N_19530,N_18539,N_18712);
nand U19531 (N_19531,N_18928,N_18948);
nor U19532 (N_19532,N_18121,N_18206);
nor U19533 (N_19533,N_18950,N_18689);
and U19534 (N_19534,N_18911,N_18350);
and U19535 (N_19535,N_18625,N_18008);
nor U19536 (N_19536,N_18953,N_18893);
and U19537 (N_19537,N_18448,N_18681);
nand U19538 (N_19538,N_18536,N_18949);
and U19539 (N_19539,N_18244,N_18895);
nor U19540 (N_19540,N_18809,N_18081);
nand U19541 (N_19541,N_18825,N_18250);
nand U19542 (N_19542,N_18702,N_18888);
and U19543 (N_19543,N_18514,N_18255);
nand U19544 (N_19544,N_18919,N_18021);
xor U19545 (N_19545,N_18732,N_18331);
nand U19546 (N_19546,N_18664,N_18669);
and U19547 (N_19547,N_18447,N_18962);
and U19548 (N_19548,N_18523,N_18560);
or U19549 (N_19549,N_18440,N_18564);
and U19550 (N_19550,N_18641,N_18076);
xor U19551 (N_19551,N_18675,N_18049);
or U19552 (N_19552,N_18472,N_18434);
nor U19553 (N_19553,N_18973,N_18626);
nor U19554 (N_19554,N_18335,N_18437);
xor U19555 (N_19555,N_18312,N_18454);
xor U19556 (N_19556,N_18249,N_18062);
nor U19557 (N_19557,N_18565,N_18292);
nand U19558 (N_19558,N_18700,N_18782);
or U19559 (N_19559,N_18275,N_18764);
nor U19560 (N_19560,N_18706,N_18296);
xor U19561 (N_19561,N_18466,N_18456);
xor U19562 (N_19562,N_18988,N_18367);
nor U19563 (N_19563,N_18232,N_18271);
xnor U19564 (N_19564,N_18334,N_18728);
or U19565 (N_19565,N_18053,N_18418);
xor U19566 (N_19566,N_18942,N_18085);
or U19567 (N_19567,N_18823,N_18244);
xor U19568 (N_19568,N_18256,N_18127);
nor U19569 (N_19569,N_18294,N_18479);
nand U19570 (N_19570,N_18599,N_18392);
and U19571 (N_19571,N_18553,N_18126);
nor U19572 (N_19572,N_18165,N_18779);
and U19573 (N_19573,N_18866,N_18215);
nand U19574 (N_19574,N_18023,N_18245);
or U19575 (N_19575,N_18463,N_18364);
and U19576 (N_19576,N_18912,N_18672);
or U19577 (N_19577,N_18714,N_18819);
or U19578 (N_19578,N_18112,N_18114);
nor U19579 (N_19579,N_18037,N_18914);
xor U19580 (N_19580,N_18146,N_18192);
xnor U19581 (N_19581,N_18179,N_18737);
xor U19582 (N_19582,N_18047,N_18473);
nor U19583 (N_19583,N_18843,N_18698);
and U19584 (N_19584,N_18073,N_18428);
xnor U19585 (N_19585,N_18067,N_18336);
nor U19586 (N_19586,N_18993,N_18442);
nor U19587 (N_19587,N_18842,N_18476);
xor U19588 (N_19588,N_18030,N_18420);
xnor U19589 (N_19589,N_18168,N_18225);
or U19590 (N_19590,N_18215,N_18155);
nand U19591 (N_19591,N_18356,N_18255);
xnor U19592 (N_19592,N_18124,N_18595);
xnor U19593 (N_19593,N_18509,N_18499);
and U19594 (N_19594,N_18124,N_18712);
nand U19595 (N_19595,N_18609,N_18565);
xnor U19596 (N_19596,N_18442,N_18390);
nand U19597 (N_19597,N_18542,N_18039);
xnor U19598 (N_19598,N_18226,N_18174);
nor U19599 (N_19599,N_18293,N_18024);
nor U19600 (N_19600,N_18307,N_18395);
and U19601 (N_19601,N_18864,N_18678);
xor U19602 (N_19602,N_18366,N_18264);
or U19603 (N_19603,N_18476,N_18064);
nand U19604 (N_19604,N_18523,N_18042);
nand U19605 (N_19605,N_18569,N_18301);
xnor U19606 (N_19606,N_18704,N_18047);
nand U19607 (N_19607,N_18530,N_18463);
nor U19608 (N_19608,N_18140,N_18174);
and U19609 (N_19609,N_18217,N_18687);
or U19610 (N_19610,N_18139,N_18671);
and U19611 (N_19611,N_18176,N_18562);
xnor U19612 (N_19612,N_18480,N_18868);
nand U19613 (N_19613,N_18220,N_18867);
xnor U19614 (N_19614,N_18179,N_18628);
nand U19615 (N_19615,N_18534,N_18196);
nand U19616 (N_19616,N_18994,N_18519);
xor U19617 (N_19617,N_18824,N_18826);
or U19618 (N_19618,N_18300,N_18864);
xnor U19619 (N_19619,N_18458,N_18494);
nor U19620 (N_19620,N_18584,N_18553);
nor U19621 (N_19621,N_18332,N_18925);
or U19622 (N_19622,N_18820,N_18245);
and U19623 (N_19623,N_18072,N_18544);
and U19624 (N_19624,N_18609,N_18042);
nand U19625 (N_19625,N_18578,N_18577);
or U19626 (N_19626,N_18543,N_18760);
nand U19627 (N_19627,N_18700,N_18816);
and U19628 (N_19628,N_18683,N_18973);
or U19629 (N_19629,N_18130,N_18434);
nand U19630 (N_19630,N_18991,N_18831);
or U19631 (N_19631,N_18315,N_18715);
nor U19632 (N_19632,N_18946,N_18614);
nor U19633 (N_19633,N_18021,N_18572);
or U19634 (N_19634,N_18949,N_18559);
xnor U19635 (N_19635,N_18275,N_18894);
and U19636 (N_19636,N_18399,N_18761);
and U19637 (N_19637,N_18384,N_18906);
and U19638 (N_19638,N_18244,N_18505);
or U19639 (N_19639,N_18593,N_18335);
nand U19640 (N_19640,N_18650,N_18548);
and U19641 (N_19641,N_18511,N_18791);
nand U19642 (N_19642,N_18986,N_18286);
and U19643 (N_19643,N_18011,N_18523);
xnor U19644 (N_19644,N_18435,N_18030);
nand U19645 (N_19645,N_18139,N_18730);
xor U19646 (N_19646,N_18668,N_18466);
xor U19647 (N_19647,N_18116,N_18566);
nand U19648 (N_19648,N_18858,N_18747);
nor U19649 (N_19649,N_18909,N_18464);
and U19650 (N_19650,N_18336,N_18551);
nand U19651 (N_19651,N_18341,N_18253);
or U19652 (N_19652,N_18873,N_18623);
xor U19653 (N_19653,N_18349,N_18310);
nor U19654 (N_19654,N_18380,N_18447);
and U19655 (N_19655,N_18474,N_18322);
xnor U19656 (N_19656,N_18415,N_18621);
or U19657 (N_19657,N_18962,N_18531);
xor U19658 (N_19658,N_18563,N_18867);
and U19659 (N_19659,N_18327,N_18444);
nand U19660 (N_19660,N_18556,N_18944);
and U19661 (N_19661,N_18023,N_18597);
nor U19662 (N_19662,N_18272,N_18278);
and U19663 (N_19663,N_18801,N_18679);
xor U19664 (N_19664,N_18049,N_18942);
xor U19665 (N_19665,N_18609,N_18400);
nand U19666 (N_19666,N_18189,N_18631);
xor U19667 (N_19667,N_18143,N_18440);
and U19668 (N_19668,N_18184,N_18512);
and U19669 (N_19669,N_18341,N_18090);
or U19670 (N_19670,N_18370,N_18284);
or U19671 (N_19671,N_18328,N_18017);
nand U19672 (N_19672,N_18680,N_18329);
or U19673 (N_19673,N_18844,N_18048);
nand U19674 (N_19674,N_18203,N_18092);
xnor U19675 (N_19675,N_18251,N_18161);
nor U19676 (N_19676,N_18685,N_18567);
nor U19677 (N_19677,N_18841,N_18591);
xnor U19678 (N_19678,N_18127,N_18326);
nand U19679 (N_19679,N_18417,N_18216);
and U19680 (N_19680,N_18860,N_18712);
nor U19681 (N_19681,N_18937,N_18224);
or U19682 (N_19682,N_18865,N_18134);
or U19683 (N_19683,N_18003,N_18822);
xnor U19684 (N_19684,N_18621,N_18717);
xnor U19685 (N_19685,N_18723,N_18685);
or U19686 (N_19686,N_18177,N_18431);
xor U19687 (N_19687,N_18554,N_18204);
xnor U19688 (N_19688,N_18104,N_18857);
and U19689 (N_19689,N_18972,N_18779);
nor U19690 (N_19690,N_18944,N_18601);
xnor U19691 (N_19691,N_18155,N_18887);
or U19692 (N_19692,N_18667,N_18250);
xor U19693 (N_19693,N_18327,N_18007);
and U19694 (N_19694,N_18426,N_18196);
and U19695 (N_19695,N_18600,N_18794);
or U19696 (N_19696,N_18568,N_18198);
or U19697 (N_19697,N_18990,N_18852);
and U19698 (N_19698,N_18084,N_18960);
nand U19699 (N_19699,N_18321,N_18512);
nand U19700 (N_19700,N_18144,N_18493);
nand U19701 (N_19701,N_18188,N_18895);
nand U19702 (N_19702,N_18032,N_18568);
nor U19703 (N_19703,N_18516,N_18256);
nand U19704 (N_19704,N_18747,N_18857);
and U19705 (N_19705,N_18985,N_18146);
or U19706 (N_19706,N_18325,N_18863);
xor U19707 (N_19707,N_18186,N_18572);
nor U19708 (N_19708,N_18107,N_18342);
xor U19709 (N_19709,N_18623,N_18216);
or U19710 (N_19710,N_18276,N_18700);
and U19711 (N_19711,N_18619,N_18921);
nand U19712 (N_19712,N_18460,N_18374);
nand U19713 (N_19713,N_18331,N_18272);
nand U19714 (N_19714,N_18134,N_18946);
nor U19715 (N_19715,N_18033,N_18002);
nand U19716 (N_19716,N_18378,N_18517);
or U19717 (N_19717,N_18727,N_18583);
nor U19718 (N_19718,N_18504,N_18257);
or U19719 (N_19719,N_18849,N_18603);
or U19720 (N_19720,N_18824,N_18361);
and U19721 (N_19721,N_18535,N_18673);
nor U19722 (N_19722,N_18939,N_18758);
nor U19723 (N_19723,N_18642,N_18550);
xor U19724 (N_19724,N_18375,N_18883);
and U19725 (N_19725,N_18551,N_18703);
or U19726 (N_19726,N_18325,N_18363);
xor U19727 (N_19727,N_18673,N_18666);
nor U19728 (N_19728,N_18485,N_18570);
and U19729 (N_19729,N_18021,N_18350);
or U19730 (N_19730,N_18480,N_18739);
or U19731 (N_19731,N_18215,N_18122);
nor U19732 (N_19732,N_18551,N_18111);
or U19733 (N_19733,N_18555,N_18431);
or U19734 (N_19734,N_18727,N_18718);
nor U19735 (N_19735,N_18769,N_18511);
nor U19736 (N_19736,N_18507,N_18856);
nor U19737 (N_19737,N_18970,N_18508);
xor U19738 (N_19738,N_18344,N_18411);
and U19739 (N_19739,N_18516,N_18628);
and U19740 (N_19740,N_18750,N_18333);
and U19741 (N_19741,N_18914,N_18039);
nand U19742 (N_19742,N_18827,N_18960);
or U19743 (N_19743,N_18306,N_18061);
and U19744 (N_19744,N_18302,N_18906);
and U19745 (N_19745,N_18330,N_18127);
nor U19746 (N_19746,N_18443,N_18704);
or U19747 (N_19747,N_18574,N_18337);
or U19748 (N_19748,N_18792,N_18982);
and U19749 (N_19749,N_18541,N_18802);
xor U19750 (N_19750,N_18207,N_18194);
and U19751 (N_19751,N_18590,N_18403);
nand U19752 (N_19752,N_18835,N_18547);
nor U19753 (N_19753,N_18357,N_18030);
or U19754 (N_19754,N_18960,N_18297);
and U19755 (N_19755,N_18206,N_18692);
or U19756 (N_19756,N_18926,N_18641);
nor U19757 (N_19757,N_18607,N_18971);
or U19758 (N_19758,N_18090,N_18981);
nor U19759 (N_19759,N_18630,N_18694);
or U19760 (N_19760,N_18415,N_18206);
nor U19761 (N_19761,N_18703,N_18701);
nand U19762 (N_19762,N_18671,N_18288);
xor U19763 (N_19763,N_18973,N_18415);
nor U19764 (N_19764,N_18921,N_18017);
nand U19765 (N_19765,N_18816,N_18053);
xor U19766 (N_19766,N_18854,N_18746);
and U19767 (N_19767,N_18629,N_18778);
nand U19768 (N_19768,N_18746,N_18058);
or U19769 (N_19769,N_18465,N_18023);
nand U19770 (N_19770,N_18312,N_18707);
nand U19771 (N_19771,N_18558,N_18387);
xor U19772 (N_19772,N_18127,N_18880);
nand U19773 (N_19773,N_18402,N_18051);
xnor U19774 (N_19774,N_18712,N_18865);
or U19775 (N_19775,N_18968,N_18110);
nor U19776 (N_19776,N_18867,N_18266);
nand U19777 (N_19777,N_18919,N_18487);
or U19778 (N_19778,N_18631,N_18232);
nand U19779 (N_19779,N_18724,N_18945);
xnor U19780 (N_19780,N_18905,N_18298);
nand U19781 (N_19781,N_18086,N_18393);
and U19782 (N_19782,N_18509,N_18622);
xor U19783 (N_19783,N_18844,N_18770);
or U19784 (N_19784,N_18410,N_18329);
xor U19785 (N_19785,N_18619,N_18793);
or U19786 (N_19786,N_18882,N_18847);
xnor U19787 (N_19787,N_18913,N_18751);
or U19788 (N_19788,N_18111,N_18570);
and U19789 (N_19789,N_18577,N_18094);
xor U19790 (N_19790,N_18191,N_18621);
or U19791 (N_19791,N_18334,N_18753);
nand U19792 (N_19792,N_18981,N_18241);
xnor U19793 (N_19793,N_18414,N_18732);
or U19794 (N_19794,N_18457,N_18033);
and U19795 (N_19795,N_18696,N_18031);
nand U19796 (N_19796,N_18245,N_18757);
xor U19797 (N_19797,N_18014,N_18125);
nand U19798 (N_19798,N_18129,N_18356);
nand U19799 (N_19799,N_18729,N_18360);
nand U19800 (N_19800,N_18852,N_18420);
and U19801 (N_19801,N_18323,N_18387);
or U19802 (N_19802,N_18647,N_18248);
nand U19803 (N_19803,N_18023,N_18707);
xor U19804 (N_19804,N_18814,N_18268);
and U19805 (N_19805,N_18965,N_18487);
xor U19806 (N_19806,N_18826,N_18471);
nand U19807 (N_19807,N_18702,N_18576);
and U19808 (N_19808,N_18674,N_18217);
or U19809 (N_19809,N_18699,N_18436);
and U19810 (N_19810,N_18513,N_18318);
or U19811 (N_19811,N_18069,N_18982);
or U19812 (N_19812,N_18056,N_18597);
or U19813 (N_19813,N_18653,N_18716);
and U19814 (N_19814,N_18386,N_18909);
and U19815 (N_19815,N_18119,N_18812);
and U19816 (N_19816,N_18919,N_18721);
xnor U19817 (N_19817,N_18925,N_18243);
xnor U19818 (N_19818,N_18638,N_18889);
xor U19819 (N_19819,N_18496,N_18948);
or U19820 (N_19820,N_18299,N_18956);
nand U19821 (N_19821,N_18486,N_18979);
or U19822 (N_19822,N_18026,N_18928);
xnor U19823 (N_19823,N_18996,N_18908);
nand U19824 (N_19824,N_18138,N_18718);
xnor U19825 (N_19825,N_18460,N_18540);
or U19826 (N_19826,N_18691,N_18580);
nand U19827 (N_19827,N_18274,N_18975);
nand U19828 (N_19828,N_18342,N_18088);
xnor U19829 (N_19829,N_18852,N_18049);
xor U19830 (N_19830,N_18464,N_18545);
or U19831 (N_19831,N_18116,N_18663);
and U19832 (N_19832,N_18246,N_18982);
nor U19833 (N_19833,N_18810,N_18730);
nor U19834 (N_19834,N_18238,N_18569);
nand U19835 (N_19835,N_18801,N_18767);
xor U19836 (N_19836,N_18323,N_18096);
xnor U19837 (N_19837,N_18034,N_18918);
or U19838 (N_19838,N_18288,N_18012);
xor U19839 (N_19839,N_18407,N_18269);
or U19840 (N_19840,N_18342,N_18548);
nand U19841 (N_19841,N_18140,N_18446);
or U19842 (N_19842,N_18016,N_18721);
xor U19843 (N_19843,N_18627,N_18209);
xor U19844 (N_19844,N_18034,N_18942);
and U19845 (N_19845,N_18581,N_18947);
or U19846 (N_19846,N_18321,N_18932);
xnor U19847 (N_19847,N_18408,N_18438);
nand U19848 (N_19848,N_18947,N_18029);
or U19849 (N_19849,N_18882,N_18998);
xor U19850 (N_19850,N_18625,N_18569);
or U19851 (N_19851,N_18329,N_18772);
nand U19852 (N_19852,N_18662,N_18680);
xor U19853 (N_19853,N_18983,N_18158);
xnor U19854 (N_19854,N_18788,N_18399);
xnor U19855 (N_19855,N_18030,N_18964);
or U19856 (N_19856,N_18064,N_18104);
nor U19857 (N_19857,N_18846,N_18520);
and U19858 (N_19858,N_18460,N_18378);
nand U19859 (N_19859,N_18163,N_18318);
nor U19860 (N_19860,N_18617,N_18899);
xor U19861 (N_19861,N_18866,N_18390);
nand U19862 (N_19862,N_18280,N_18227);
and U19863 (N_19863,N_18637,N_18813);
nor U19864 (N_19864,N_18000,N_18755);
nand U19865 (N_19865,N_18755,N_18581);
nand U19866 (N_19866,N_18537,N_18257);
or U19867 (N_19867,N_18530,N_18787);
or U19868 (N_19868,N_18146,N_18467);
nand U19869 (N_19869,N_18855,N_18219);
and U19870 (N_19870,N_18347,N_18570);
xor U19871 (N_19871,N_18884,N_18311);
or U19872 (N_19872,N_18899,N_18437);
nor U19873 (N_19873,N_18604,N_18584);
xor U19874 (N_19874,N_18435,N_18734);
nand U19875 (N_19875,N_18117,N_18269);
nand U19876 (N_19876,N_18315,N_18327);
nand U19877 (N_19877,N_18719,N_18534);
nand U19878 (N_19878,N_18998,N_18363);
or U19879 (N_19879,N_18748,N_18548);
xor U19880 (N_19880,N_18765,N_18186);
xnor U19881 (N_19881,N_18387,N_18097);
xor U19882 (N_19882,N_18338,N_18336);
xor U19883 (N_19883,N_18813,N_18721);
nor U19884 (N_19884,N_18237,N_18342);
or U19885 (N_19885,N_18231,N_18335);
nand U19886 (N_19886,N_18332,N_18805);
xnor U19887 (N_19887,N_18197,N_18470);
or U19888 (N_19888,N_18251,N_18680);
nand U19889 (N_19889,N_18307,N_18593);
nor U19890 (N_19890,N_18546,N_18236);
or U19891 (N_19891,N_18534,N_18446);
and U19892 (N_19892,N_18425,N_18537);
nand U19893 (N_19893,N_18651,N_18080);
xnor U19894 (N_19894,N_18918,N_18579);
or U19895 (N_19895,N_18556,N_18007);
nand U19896 (N_19896,N_18290,N_18616);
and U19897 (N_19897,N_18754,N_18306);
nand U19898 (N_19898,N_18544,N_18479);
or U19899 (N_19899,N_18943,N_18195);
nand U19900 (N_19900,N_18427,N_18659);
xnor U19901 (N_19901,N_18582,N_18187);
or U19902 (N_19902,N_18740,N_18618);
and U19903 (N_19903,N_18012,N_18658);
and U19904 (N_19904,N_18514,N_18782);
xor U19905 (N_19905,N_18309,N_18779);
and U19906 (N_19906,N_18343,N_18280);
nand U19907 (N_19907,N_18158,N_18628);
and U19908 (N_19908,N_18972,N_18127);
or U19909 (N_19909,N_18546,N_18298);
nor U19910 (N_19910,N_18522,N_18266);
xor U19911 (N_19911,N_18094,N_18488);
and U19912 (N_19912,N_18860,N_18665);
and U19913 (N_19913,N_18471,N_18504);
and U19914 (N_19914,N_18312,N_18636);
nand U19915 (N_19915,N_18382,N_18195);
or U19916 (N_19916,N_18815,N_18793);
or U19917 (N_19917,N_18871,N_18131);
and U19918 (N_19918,N_18251,N_18409);
and U19919 (N_19919,N_18679,N_18100);
xor U19920 (N_19920,N_18111,N_18804);
and U19921 (N_19921,N_18086,N_18078);
xor U19922 (N_19922,N_18086,N_18254);
and U19923 (N_19923,N_18362,N_18326);
or U19924 (N_19924,N_18829,N_18113);
nor U19925 (N_19925,N_18264,N_18590);
nand U19926 (N_19926,N_18312,N_18367);
nor U19927 (N_19927,N_18986,N_18681);
nor U19928 (N_19928,N_18440,N_18451);
or U19929 (N_19929,N_18661,N_18276);
nand U19930 (N_19930,N_18978,N_18557);
nor U19931 (N_19931,N_18991,N_18686);
or U19932 (N_19932,N_18033,N_18679);
xor U19933 (N_19933,N_18657,N_18202);
or U19934 (N_19934,N_18568,N_18668);
nand U19935 (N_19935,N_18236,N_18751);
nand U19936 (N_19936,N_18284,N_18176);
xnor U19937 (N_19937,N_18805,N_18580);
and U19938 (N_19938,N_18609,N_18646);
or U19939 (N_19939,N_18105,N_18501);
nor U19940 (N_19940,N_18046,N_18909);
nand U19941 (N_19941,N_18742,N_18081);
nand U19942 (N_19942,N_18010,N_18139);
nor U19943 (N_19943,N_18834,N_18599);
nor U19944 (N_19944,N_18789,N_18683);
nor U19945 (N_19945,N_18575,N_18722);
and U19946 (N_19946,N_18166,N_18019);
or U19947 (N_19947,N_18742,N_18108);
or U19948 (N_19948,N_18890,N_18583);
nor U19949 (N_19949,N_18666,N_18906);
nor U19950 (N_19950,N_18419,N_18647);
and U19951 (N_19951,N_18098,N_18688);
and U19952 (N_19952,N_18277,N_18895);
nor U19953 (N_19953,N_18363,N_18003);
and U19954 (N_19954,N_18444,N_18729);
and U19955 (N_19955,N_18247,N_18357);
nand U19956 (N_19956,N_18554,N_18107);
nand U19957 (N_19957,N_18629,N_18564);
nor U19958 (N_19958,N_18415,N_18756);
or U19959 (N_19959,N_18494,N_18003);
or U19960 (N_19960,N_18640,N_18876);
nand U19961 (N_19961,N_18886,N_18210);
nand U19962 (N_19962,N_18366,N_18712);
nand U19963 (N_19963,N_18024,N_18875);
or U19964 (N_19964,N_18169,N_18581);
nand U19965 (N_19965,N_18553,N_18742);
or U19966 (N_19966,N_18159,N_18697);
nand U19967 (N_19967,N_18817,N_18981);
nor U19968 (N_19968,N_18368,N_18154);
and U19969 (N_19969,N_18799,N_18262);
or U19970 (N_19970,N_18669,N_18947);
nor U19971 (N_19971,N_18486,N_18621);
nand U19972 (N_19972,N_18579,N_18493);
or U19973 (N_19973,N_18883,N_18318);
and U19974 (N_19974,N_18746,N_18868);
xnor U19975 (N_19975,N_18032,N_18475);
nand U19976 (N_19976,N_18031,N_18573);
nor U19977 (N_19977,N_18087,N_18816);
or U19978 (N_19978,N_18174,N_18152);
xnor U19979 (N_19979,N_18703,N_18493);
and U19980 (N_19980,N_18119,N_18141);
xor U19981 (N_19981,N_18908,N_18437);
and U19982 (N_19982,N_18644,N_18359);
and U19983 (N_19983,N_18920,N_18996);
nor U19984 (N_19984,N_18728,N_18866);
and U19985 (N_19985,N_18744,N_18023);
nor U19986 (N_19986,N_18848,N_18994);
nor U19987 (N_19987,N_18919,N_18839);
nor U19988 (N_19988,N_18827,N_18695);
and U19989 (N_19989,N_18152,N_18979);
nand U19990 (N_19990,N_18353,N_18196);
or U19991 (N_19991,N_18027,N_18175);
xor U19992 (N_19992,N_18012,N_18324);
or U19993 (N_19993,N_18669,N_18440);
nand U19994 (N_19994,N_18599,N_18480);
nor U19995 (N_19995,N_18290,N_18653);
and U19996 (N_19996,N_18031,N_18839);
nor U19997 (N_19997,N_18529,N_18112);
or U19998 (N_19998,N_18624,N_18549);
or U19999 (N_19999,N_18062,N_18155);
nor U20000 (N_20000,N_19444,N_19561);
and U20001 (N_20001,N_19057,N_19259);
and U20002 (N_20002,N_19384,N_19182);
nand U20003 (N_20003,N_19228,N_19572);
and U20004 (N_20004,N_19526,N_19743);
nor U20005 (N_20005,N_19287,N_19310);
and U20006 (N_20006,N_19091,N_19293);
or U20007 (N_20007,N_19985,N_19318);
and U20008 (N_20008,N_19665,N_19388);
and U20009 (N_20009,N_19632,N_19816);
xnor U20010 (N_20010,N_19161,N_19063);
xor U20011 (N_20011,N_19194,N_19564);
nand U20012 (N_20012,N_19284,N_19213);
or U20013 (N_20013,N_19181,N_19753);
xnor U20014 (N_20014,N_19639,N_19558);
nand U20015 (N_20015,N_19716,N_19476);
nand U20016 (N_20016,N_19676,N_19389);
and U20017 (N_20017,N_19175,N_19799);
nor U20018 (N_20018,N_19528,N_19608);
nand U20019 (N_20019,N_19510,N_19423);
nand U20020 (N_20020,N_19226,N_19280);
or U20021 (N_20021,N_19415,N_19711);
nand U20022 (N_20022,N_19603,N_19512);
and U20023 (N_20023,N_19801,N_19539);
nor U20024 (N_20024,N_19039,N_19611);
xor U20025 (N_20025,N_19080,N_19852);
nand U20026 (N_20026,N_19068,N_19715);
or U20027 (N_20027,N_19366,N_19469);
and U20028 (N_20028,N_19976,N_19565);
nand U20029 (N_20029,N_19073,N_19505);
or U20030 (N_20030,N_19000,N_19867);
nand U20031 (N_20031,N_19997,N_19036);
or U20032 (N_20032,N_19133,N_19405);
and U20033 (N_20033,N_19911,N_19829);
nor U20034 (N_20034,N_19798,N_19647);
nor U20035 (N_20035,N_19028,N_19687);
or U20036 (N_20036,N_19104,N_19783);
or U20037 (N_20037,N_19762,N_19788);
and U20038 (N_20038,N_19099,N_19842);
or U20039 (N_20039,N_19873,N_19595);
nand U20040 (N_20040,N_19920,N_19996);
and U20041 (N_20041,N_19999,N_19645);
or U20042 (N_20042,N_19882,N_19365);
xor U20043 (N_20043,N_19797,N_19907);
xor U20044 (N_20044,N_19767,N_19468);
and U20045 (N_20045,N_19236,N_19464);
and U20046 (N_20046,N_19584,N_19966);
and U20047 (N_20047,N_19978,N_19901);
or U20048 (N_20048,N_19625,N_19338);
nor U20049 (N_20049,N_19532,N_19321);
and U20050 (N_20050,N_19195,N_19106);
and U20051 (N_20051,N_19936,N_19176);
and U20052 (N_20052,N_19125,N_19832);
xnor U20053 (N_20053,N_19589,N_19810);
nand U20054 (N_20054,N_19067,N_19433);
and U20055 (N_20055,N_19878,N_19261);
nor U20056 (N_20056,N_19568,N_19764);
xnor U20057 (N_20057,N_19846,N_19504);
or U20058 (N_20058,N_19225,N_19605);
nand U20059 (N_20059,N_19171,N_19369);
nor U20060 (N_20060,N_19138,N_19734);
and U20061 (N_20061,N_19332,N_19484);
nor U20062 (N_20062,N_19136,N_19507);
and U20063 (N_20063,N_19214,N_19038);
or U20064 (N_20064,N_19071,N_19898);
nor U20065 (N_20065,N_19344,N_19818);
or U20066 (N_20066,N_19612,N_19706);
or U20067 (N_20067,N_19056,N_19269);
or U20068 (N_20068,N_19440,N_19436);
and U20069 (N_20069,N_19904,N_19992);
xor U20070 (N_20070,N_19302,N_19574);
nor U20071 (N_20071,N_19265,N_19411);
xor U20072 (N_20072,N_19995,N_19243);
nand U20073 (N_20073,N_19749,N_19520);
xor U20074 (N_20074,N_19570,N_19777);
nor U20075 (N_20075,N_19342,N_19858);
and U20076 (N_20076,N_19972,N_19640);
or U20077 (N_20077,N_19193,N_19130);
nor U20078 (N_20078,N_19679,N_19566);
or U20079 (N_20079,N_19399,N_19703);
xnor U20080 (N_20080,N_19353,N_19820);
nor U20081 (N_20081,N_19202,N_19337);
nor U20082 (N_20082,N_19147,N_19299);
xor U20083 (N_20083,N_19724,N_19208);
and U20084 (N_20084,N_19308,N_19917);
xor U20085 (N_20085,N_19438,N_19981);
nand U20086 (N_20086,N_19560,N_19479);
and U20087 (N_20087,N_19790,N_19025);
and U20088 (N_20088,N_19628,N_19103);
and U20089 (N_20089,N_19970,N_19094);
and U20090 (N_20090,N_19060,N_19721);
and U20091 (N_20091,N_19222,N_19641);
nand U20092 (N_20092,N_19069,N_19467);
xnor U20093 (N_20093,N_19412,N_19159);
nand U20094 (N_20094,N_19210,N_19049);
or U20095 (N_20095,N_19102,N_19553);
or U20096 (N_20096,N_19821,N_19227);
nor U20097 (N_20097,N_19922,N_19478);
nand U20098 (N_20098,N_19508,N_19591);
and U20099 (N_20099,N_19569,N_19352);
and U20100 (N_20100,N_19634,N_19708);
or U20101 (N_20101,N_19778,N_19160);
nor U20102 (N_20102,N_19989,N_19607);
xnor U20103 (N_20103,N_19908,N_19295);
xor U20104 (N_20104,N_19270,N_19495);
or U20105 (N_20105,N_19417,N_19154);
and U20106 (N_20106,N_19745,N_19223);
and U20107 (N_20107,N_19522,N_19865);
nor U20108 (N_20108,N_19646,N_19670);
or U20109 (N_20109,N_19152,N_19343);
or U20110 (N_20110,N_19918,N_19340);
nor U20111 (N_20111,N_19017,N_19533);
nor U20112 (N_20112,N_19671,N_19610);
nand U20113 (N_20113,N_19792,N_19040);
and U20114 (N_20114,N_19705,N_19179);
or U20115 (N_20115,N_19163,N_19298);
nand U20116 (N_20116,N_19112,N_19317);
nor U20117 (N_20117,N_19198,N_19902);
and U20118 (N_20118,N_19822,N_19597);
xor U20119 (N_20119,N_19551,N_19747);
nand U20120 (N_20120,N_19111,N_19237);
nor U20121 (N_20121,N_19325,N_19364);
or U20122 (N_20122,N_19011,N_19961);
or U20123 (N_20123,N_19741,N_19001);
nand U20124 (N_20124,N_19126,N_19370);
and U20125 (N_20125,N_19482,N_19492);
nand U20126 (N_20126,N_19037,N_19662);
nor U20127 (N_20127,N_19914,N_19095);
or U20128 (N_20128,N_19473,N_19431);
and U20129 (N_20129,N_19475,N_19066);
xor U20130 (N_20130,N_19916,N_19523);
and U20131 (N_20131,N_19241,N_19189);
or U20132 (N_20132,N_19165,N_19075);
or U20133 (N_20133,N_19651,N_19132);
and U20134 (N_20134,N_19022,N_19768);
xor U20135 (N_20135,N_19348,N_19502);
nand U20136 (N_20136,N_19041,N_19268);
and U20137 (N_20137,N_19454,N_19733);
nand U20138 (N_20138,N_19315,N_19903);
nor U20139 (N_20139,N_19391,N_19928);
nor U20140 (N_20140,N_19546,N_19013);
xor U20141 (N_20141,N_19371,N_19659);
nor U20142 (N_20142,N_19969,N_19868);
or U20143 (N_20143,N_19187,N_19896);
nor U20144 (N_20144,N_19872,N_19117);
nand U20145 (N_20145,N_19627,N_19447);
nor U20146 (N_20146,N_19998,N_19082);
xnor U20147 (N_20147,N_19979,N_19601);
nand U20148 (N_20148,N_19459,N_19373);
and U20149 (N_20149,N_19116,N_19127);
xor U20150 (N_20150,N_19205,N_19453);
nand U20151 (N_20151,N_19004,N_19847);
and U20152 (N_20152,N_19256,N_19139);
xnor U20153 (N_20153,N_19919,N_19363);
or U20154 (N_20154,N_19772,N_19808);
nor U20155 (N_20155,N_19756,N_19575);
nor U20156 (N_20156,N_19292,N_19623);
nand U20157 (N_20157,N_19650,N_19758);
and U20158 (N_20158,N_19658,N_19812);
nor U20159 (N_20159,N_19582,N_19064);
or U20160 (N_20160,N_19644,N_19486);
and U20161 (N_20161,N_19421,N_19264);
or U20162 (N_20162,N_19588,N_19947);
or U20163 (N_20163,N_19185,N_19912);
xor U20164 (N_20164,N_19613,N_19831);
xnor U20165 (N_20165,N_19144,N_19124);
or U20166 (N_20166,N_19910,N_19660);
xor U20167 (N_20167,N_19844,N_19752);
and U20168 (N_20168,N_19290,N_19948);
nor U20169 (N_20169,N_19047,N_19407);
and U20170 (N_20170,N_19974,N_19984);
or U20171 (N_20171,N_19500,N_19673);
or U20172 (N_20172,N_19770,N_19032);
or U20173 (N_20173,N_19090,N_19334);
and U20174 (N_20174,N_19240,N_19326);
nand U20175 (N_20175,N_19414,N_19455);
and U20176 (N_20176,N_19465,N_19531);
nor U20177 (N_20177,N_19314,N_19804);
xor U20178 (N_20178,N_19341,N_19172);
xnor U20179 (N_20179,N_19699,N_19380);
nand U20180 (N_20180,N_19020,N_19294);
nor U20181 (N_20181,N_19814,N_19760);
and U20182 (N_20182,N_19953,N_19986);
and U20183 (N_20183,N_19143,N_19113);
nor U20184 (N_20184,N_19007,N_19184);
xnor U20185 (N_20185,N_19305,N_19925);
nor U20186 (N_20186,N_19381,N_19451);
nand U20187 (N_20187,N_19696,N_19602);
nor U20188 (N_20188,N_19875,N_19689);
xor U20189 (N_20189,N_19681,N_19796);
or U20190 (N_20190,N_19445,N_19636);
or U20191 (N_20191,N_19296,N_19174);
or U20192 (N_20192,N_19690,N_19471);
xor U20193 (N_20193,N_19629,N_19887);
xor U20194 (N_20194,N_19016,N_19496);
nand U20195 (N_20195,N_19221,N_19516);
nor U20196 (N_20196,N_19537,N_19803);
or U20197 (N_20197,N_19311,N_19076);
or U20198 (N_20198,N_19331,N_19990);
and U20199 (N_20199,N_19404,N_19450);
or U20200 (N_20200,N_19664,N_19012);
xor U20201 (N_20201,N_19432,N_19894);
or U20202 (N_20202,N_19286,N_19950);
xor U20203 (N_20203,N_19489,N_19400);
nor U20204 (N_20204,N_19915,N_19178);
or U20205 (N_20205,N_19534,N_19114);
and U20206 (N_20206,N_19149,N_19230);
nor U20207 (N_20207,N_19669,N_19006);
xnor U20208 (N_20208,N_19281,N_19245);
and U20209 (N_20209,N_19973,N_19283);
or U20210 (N_20210,N_19834,N_19677);
or U20211 (N_20211,N_19258,N_19637);
nor U20212 (N_20212,N_19249,N_19750);
and U20213 (N_20213,N_19253,N_19543);
nor U20214 (N_20214,N_19631,N_19385);
nor U20215 (N_20215,N_19759,N_19050);
and U20216 (N_20216,N_19470,N_19190);
or U20217 (N_20217,N_19170,N_19320);
and U20218 (N_20218,N_19098,N_19672);
xnor U20219 (N_20219,N_19379,N_19871);
xnor U20220 (N_20220,N_19604,N_19443);
and U20221 (N_20221,N_19648,N_19666);
nand U20222 (N_20222,N_19525,N_19786);
and U20223 (N_20223,N_19577,N_19954);
nand U20224 (N_20224,N_19813,N_19110);
nand U20225 (N_20225,N_19840,N_19769);
xnor U20226 (N_20226,N_19324,N_19924);
nand U20227 (N_20227,N_19550,N_19586);
nor U20228 (N_20228,N_19958,N_19065);
and U20229 (N_20229,N_19555,N_19218);
xnor U20230 (N_20230,N_19619,N_19649);
xor U20231 (N_20231,N_19053,N_19698);
and U20232 (N_20232,N_19590,N_19336);
nand U20233 (N_20233,N_19861,N_19598);
and U20234 (N_20234,N_19773,N_19817);
or U20235 (N_20235,N_19939,N_19600);
and U20236 (N_20236,N_19335,N_19105);
and U20237 (N_20237,N_19626,N_19559);
nor U20238 (N_20238,N_19420,N_19633);
or U20239 (N_20239,N_19782,N_19115);
or U20240 (N_20240,N_19250,N_19735);
nor U20241 (N_20241,N_19988,N_19192);
nor U20242 (N_20242,N_19277,N_19885);
nand U20243 (N_20243,N_19694,N_19488);
and U20244 (N_20244,N_19146,N_19680);
nor U20245 (N_20245,N_19029,N_19313);
and U20246 (N_20246,N_19397,N_19862);
or U20247 (N_20247,N_19833,N_19643);
xnor U20248 (N_20248,N_19806,N_19491);
and U20249 (N_20249,N_19956,N_19191);
and U20250 (N_20250,N_19889,N_19460);
and U20251 (N_20251,N_19275,N_19009);
nand U20252 (N_20252,N_19642,N_19282);
nor U20253 (N_20253,N_19562,N_19072);
and U20254 (N_20254,N_19350,N_19955);
xnor U20255 (N_20255,N_19054,N_19118);
or U20256 (N_20256,N_19592,N_19088);
nor U20257 (N_20257,N_19480,N_19573);
and U20258 (N_20258,N_19893,N_19481);
nor U20259 (N_20259,N_19203,N_19257);
nor U20260 (N_20260,N_19635,N_19309);
or U20261 (N_20261,N_19538,N_19630);
or U20262 (N_20262,N_19678,N_19890);
nor U20263 (N_20263,N_19425,N_19289);
nand U20264 (N_20264,N_19312,N_19390);
or U20265 (N_20265,N_19836,N_19031);
xor U20266 (N_20266,N_19406,N_19005);
and U20267 (N_20267,N_19120,N_19233);
xor U20268 (N_20268,N_19501,N_19437);
and U20269 (N_20269,N_19946,N_19197);
nor U20270 (N_20270,N_19055,N_19622);
xor U20271 (N_20271,N_19167,N_19514);
nand U20272 (N_20272,N_19361,N_19306);
and U20273 (N_20273,N_19078,N_19606);
or U20274 (N_20274,N_19328,N_19485);
nor U20275 (N_20275,N_19209,N_19866);
nor U20276 (N_20276,N_19567,N_19392);
nand U20277 (N_20277,N_19329,N_19018);
or U20278 (N_20278,N_19864,N_19129);
nor U20279 (N_20279,N_19509,N_19244);
nand U20280 (N_20280,N_19211,N_19863);
nor U20281 (N_20281,N_19059,N_19273);
nand U20282 (N_20282,N_19616,N_19316);
nor U20283 (N_20283,N_19354,N_19376);
xnor U20284 (N_20284,N_19661,N_19323);
nor U20285 (N_20285,N_19932,N_19717);
nand U20286 (N_20286,N_19372,N_19702);
nand U20287 (N_20287,N_19186,N_19707);
or U20288 (N_20288,N_19419,N_19201);
or U20289 (N_20289,N_19122,N_19942);
xnor U20290 (N_20290,N_19008,N_19135);
xor U20291 (N_20291,N_19692,N_19688);
nand U20292 (N_20292,N_19895,N_19736);
and U20293 (N_20293,N_19929,N_19021);
nor U20294 (N_20294,N_19434,N_19271);
nor U20295 (N_20295,N_19754,N_19527);
or U20296 (N_20296,N_19541,N_19940);
and U20297 (N_20297,N_19980,N_19728);
xor U20298 (N_20298,N_19474,N_19837);
and U20299 (N_20299,N_19819,N_19087);
or U20300 (N_20300,N_19712,N_19401);
xor U20301 (N_20301,N_19805,N_19246);
xnor U20302 (N_20302,N_19010,N_19251);
xor U20303 (N_20303,N_19857,N_19079);
and U20304 (N_20304,N_19360,N_19499);
and U20305 (N_20305,N_19701,N_19300);
nand U20306 (N_20306,N_19351,N_19971);
and U20307 (N_20307,N_19150,N_19785);
or U20308 (N_20308,N_19853,N_19652);
nand U20309 (N_20309,N_19377,N_19835);
and U20310 (N_20310,N_19382,N_19780);
nor U20311 (N_20311,N_19166,N_19276);
nand U20312 (N_20312,N_19155,N_19386);
or U20313 (N_20313,N_19905,N_19272);
or U20314 (N_20314,N_19145,N_19183);
or U20315 (N_20315,N_19860,N_19358);
and U20316 (N_20316,N_19933,N_19472);
nand U20317 (N_20317,N_19375,N_19594);
xor U20318 (N_20318,N_19206,N_19685);
nand U20319 (N_20319,N_19503,N_19930);
nor U20320 (N_20320,N_19886,N_19739);
xor U20321 (N_20321,N_19164,N_19188);
xor U20322 (N_20322,N_19618,N_19148);
nor U20323 (N_20323,N_19457,N_19074);
nor U20324 (N_20324,N_19695,N_19725);
or U20325 (N_20325,N_19859,N_19880);
nor U20326 (N_20326,N_19897,N_19108);
xnor U20327 (N_20327,N_19439,N_19044);
and U20328 (N_20328,N_19034,N_19535);
nand U20329 (N_20329,N_19959,N_19416);
nor U20330 (N_20330,N_19937,N_19097);
or U20331 (N_20331,N_19374,N_19156);
xnor U20332 (N_20332,N_19547,N_19356);
nor U20333 (N_20333,N_19435,N_19121);
nand U20334 (N_20334,N_19429,N_19494);
nor U20335 (N_20335,N_19693,N_19809);
nor U20336 (N_20336,N_19349,N_19949);
nand U20337 (N_20337,N_19262,N_19052);
and U20338 (N_20338,N_19548,N_19675);
xnor U20339 (N_20339,N_19229,N_19802);
and U20340 (N_20340,N_19771,N_19609);
xor U20341 (N_20341,N_19709,N_19003);
and U20342 (N_20342,N_19545,N_19587);
nand U20343 (N_20343,N_19668,N_19906);
or U20344 (N_20344,N_19718,N_19913);
xor U20345 (N_20345,N_19517,N_19248);
nand U20346 (N_20346,N_19683,N_19900);
or U20347 (N_20347,N_19849,N_19430);
nor U20348 (N_20348,N_19775,N_19700);
xor U20349 (N_20349,N_19731,N_19422);
nand U20350 (N_20350,N_19874,N_19199);
xnor U20351 (N_20351,N_19585,N_19583);
nand U20352 (N_20352,N_19058,N_19506);
xor U20353 (N_20353,N_19424,N_19498);
xnor U20354 (N_20354,N_19322,N_19288);
and U20355 (N_20355,N_19217,N_19935);
nor U20356 (N_20356,N_19413,N_19776);
xnor U20357 (N_20357,N_19719,N_19409);
nor U20358 (N_20358,N_19839,N_19563);
nand U20359 (N_20359,N_19291,N_19765);
or U20360 (N_20360,N_19466,N_19303);
and U20361 (N_20361,N_19657,N_19109);
nand U20362 (N_20362,N_19119,N_19720);
and U20363 (N_20363,N_19513,N_19845);
xor U20364 (N_20364,N_19200,N_19791);
and U20365 (N_20365,N_19304,N_19779);
and U20366 (N_20366,N_19938,N_19571);
nor U20367 (N_20367,N_19394,N_19811);
and U20368 (N_20368,N_19751,N_19727);
or U20369 (N_20369,N_19869,N_19061);
or U20370 (N_20370,N_19656,N_19945);
xnor U20371 (N_20371,N_19931,N_19162);
and U20372 (N_20372,N_19378,N_19339);
nor U20373 (N_20373,N_19823,N_19267);
nand U20374 (N_20374,N_19043,N_19461);
or U20375 (N_20375,N_19691,N_19704);
or U20376 (N_20376,N_19511,N_19141);
or U20377 (N_20377,N_19697,N_19231);
or U20378 (N_20378,N_19398,N_19870);
nor U20379 (N_20379,N_19173,N_19795);
nor U20380 (N_20380,N_19019,N_19396);
nand U20381 (N_20381,N_19204,N_19987);
nand U20382 (N_20382,N_19442,N_19554);
and U20383 (N_20383,N_19621,N_19827);
xnor U20384 (N_20384,N_19487,N_19710);
nor U20385 (N_20385,N_19964,N_19083);
xor U20386 (N_20386,N_19158,N_19944);
xor U20387 (N_20387,N_19524,N_19740);
nor U20388 (N_20388,N_19219,N_19387);
nand U20389 (N_20389,N_19084,N_19046);
nor U20390 (N_20390,N_19383,N_19252);
or U20391 (N_20391,N_19123,N_19825);
xnor U20392 (N_20392,N_19714,N_19667);
nand U20393 (N_20393,N_19952,N_19794);
or U20394 (N_20394,N_19140,N_19448);
nand U20395 (N_20395,N_19216,N_19347);
and U20396 (N_20396,N_19254,N_19620);
or U20397 (N_20397,N_19909,N_19926);
xnor U20398 (N_20398,N_19490,N_19892);
nand U20399 (N_20399,N_19235,N_19856);
nand U20400 (N_20400,N_19774,N_19529);
and U20401 (N_20401,N_19826,N_19168);
nand U20402 (N_20402,N_19991,N_19763);
nor U20403 (N_20403,N_19848,N_19196);
and U20404 (N_20404,N_19757,N_19131);
xnor U20405 (N_20405,N_19838,N_19232);
or U20406 (N_20406,N_19993,N_19483);
and U20407 (N_20407,N_19030,N_19142);
nand U20408 (N_20408,N_19255,N_19975);
or U20409 (N_20409,N_19519,N_19319);
nand U20410 (N_20410,N_19549,N_19960);
or U20411 (N_20411,N_19092,N_19247);
and U20412 (N_20412,N_19238,N_19841);
xor U20413 (N_20413,N_19536,N_19544);
and U20414 (N_20414,N_19212,N_19737);
xnor U20415 (N_20415,N_19883,N_19614);
or U20416 (N_20416,N_19393,N_19345);
nor U20417 (N_20417,N_19048,N_19368);
xnor U20418 (N_20418,N_19515,N_19968);
nand U20419 (N_20419,N_19449,N_19081);
xor U20420 (N_20420,N_19748,N_19042);
nand U20421 (N_20421,N_19279,N_19815);
nor U20422 (N_20422,N_19403,N_19830);
nor U20423 (N_20423,N_19713,N_19497);
xnor U20424 (N_20424,N_19051,N_19002);
xnor U20425 (N_20425,N_19234,N_19285);
and U20426 (N_20426,N_19107,N_19965);
nor U20427 (N_20427,N_19367,N_19941);
or U20428 (N_20428,N_19026,N_19014);
nor U20429 (N_20429,N_19761,N_19408);
nand U20430 (N_20430,N_19977,N_19578);
nand U20431 (N_20431,N_19220,N_19428);
nand U20432 (N_20432,N_19521,N_19157);
nor U20433 (N_20433,N_19327,N_19301);
xnor U20434 (N_20434,N_19800,N_19557);
nand U20435 (N_20435,N_19355,N_19101);
nand U20436 (N_20436,N_19426,N_19879);
or U20437 (N_20437,N_19540,N_19684);
or U20438 (N_20438,N_19876,N_19096);
xor U20439 (N_20439,N_19333,N_19807);
or U20440 (N_20440,N_19742,N_19746);
or U20441 (N_20441,N_19884,N_19477);
xor U20442 (N_20442,N_19726,N_19024);
or U20443 (N_20443,N_19686,N_19452);
nand U20444 (N_20444,N_19274,N_19086);
nand U20445 (N_20445,N_19242,N_19653);
and U20446 (N_20446,N_19732,N_19177);
and U20447 (N_20447,N_19169,N_19446);
and U20448 (N_20448,N_19153,N_19100);
xor U20449 (N_20449,N_19580,N_19957);
xnor U20450 (N_20450,N_19346,N_19793);
or U20451 (N_20451,N_19239,N_19617);
or U20452 (N_20452,N_19784,N_19410);
or U20453 (N_20453,N_19093,N_19266);
xnor U20454 (N_20454,N_19828,N_19462);
xnor U20455 (N_20455,N_19730,N_19755);
nand U20456 (N_20456,N_19089,N_19855);
xnor U20457 (N_20457,N_19441,N_19891);
nand U20458 (N_20458,N_19663,N_19458);
or U20459 (N_20459,N_19556,N_19682);
nand U20460 (N_20460,N_19888,N_19729);
or U20461 (N_20461,N_19260,N_19654);
nand U20462 (N_20462,N_19923,N_19579);
and U20463 (N_20463,N_19151,N_19297);
nand U20464 (N_20464,N_19463,N_19615);
or U20465 (N_20465,N_19027,N_19023);
or U20466 (N_20466,N_19357,N_19134);
and U20467 (N_20467,N_19982,N_19542);
xnor U20468 (N_20468,N_19877,N_19359);
nand U20469 (N_20469,N_19552,N_19951);
and U20470 (N_20470,N_19077,N_19362);
nor U20471 (N_20471,N_19263,N_19738);
xor U20472 (N_20472,N_19850,N_19638);
or U20473 (N_20473,N_19851,N_19456);
xor U20474 (N_20474,N_19418,N_19674);
and U20475 (N_20475,N_19307,N_19085);
xor U20476 (N_20476,N_19207,N_19843);
and U20477 (N_20477,N_19789,N_19070);
and U20478 (N_20478,N_19035,N_19927);
or U20479 (N_20479,N_19599,N_19330);
xor U20480 (N_20480,N_19781,N_19596);
nor U20481 (N_20481,N_19062,N_19593);
nor U20482 (N_20482,N_19899,N_19824);
xnor U20483 (N_20483,N_19787,N_19395);
or U20484 (N_20484,N_19137,N_19128);
and U20485 (N_20485,N_19983,N_19722);
xor U20486 (N_20486,N_19723,N_19881);
and U20487 (N_20487,N_19921,N_19224);
or U20488 (N_20488,N_19427,N_19576);
nor U20489 (N_20489,N_19943,N_19994);
nand U20490 (N_20490,N_19744,N_19581);
xor U20491 (N_20491,N_19766,N_19402);
and U20492 (N_20492,N_19493,N_19045);
nor U20493 (N_20493,N_19854,N_19962);
and U20494 (N_20494,N_19180,N_19530);
xnor U20495 (N_20495,N_19518,N_19934);
nand U20496 (N_20496,N_19215,N_19278);
nand U20497 (N_20497,N_19655,N_19963);
and U20498 (N_20498,N_19967,N_19015);
and U20499 (N_20499,N_19033,N_19624);
xnor U20500 (N_20500,N_19809,N_19878);
nor U20501 (N_20501,N_19198,N_19532);
and U20502 (N_20502,N_19983,N_19054);
or U20503 (N_20503,N_19884,N_19235);
xnor U20504 (N_20504,N_19849,N_19816);
nand U20505 (N_20505,N_19321,N_19311);
nor U20506 (N_20506,N_19891,N_19694);
xor U20507 (N_20507,N_19611,N_19320);
and U20508 (N_20508,N_19109,N_19979);
xor U20509 (N_20509,N_19276,N_19799);
and U20510 (N_20510,N_19231,N_19102);
or U20511 (N_20511,N_19094,N_19649);
nand U20512 (N_20512,N_19223,N_19644);
or U20513 (N_20513,N_19889,N_19298);
nand U20514 (N_20514,N_19974,N_19885);
nor U20515 (N_20515,N_19398,N_19257);
xor U20516 (N_20516,N_19809,N_19364);
xnor U20517 (N_20517,N_19020,N_19870);
or U20518 (N_20518,N_19465,N_19524);
nand U20519 (N_20519,N_19517,N_19199);
or U20520 (N_20520,N_19413,N_19090);
or U20521 (N_20521,N_19385,N_19770);
nand U20522 (N_20522,N_19105,N_19782);
and U20523 (N_20523,N_19519,N_19618);
xor U20524 (N_20524,N_19770,N_19642);
and U20525 (N_20525,N_19130,N_19823);
xor U20526 (N_20526,N_19678,N_19742);
nand U20527 (N_20527,N_19189,N_19717);
or U20528 (N_20528,N_19230,N_19815);
xnor U20529 (N_20529,N_19392,N_19266);
nor U20530 (N_20530,N_19980,N_19247);
and U20531 (N_20531,N_19301,N_19263);
xor U20532 (N_20532,N_19579,N_19777);
nor U20533 (N_20533,N_19086,N_19358);
nor U20534 (N_20534,N_19522,N_19691);
and U20535 (N_20535,N_19522,N_19999);
nand U20536 (N_20536,N_19196,N_19722);
xor U20537 (N_20537,N_19839,N_19737);
nand U20538 (N_20538,N_19683,N_19403);
and U20539 (N_20539,N_19990,N_19246);
and U20540 (N_20540,N_19646,N_19426);
xor U20541 (N_20541,N_19651,N_19549);
or U20542 (N_20542,N_19803,N_19277);
xor U20543 (N_20543,N_19586,N_19445);
nor U20544 (N_20544,N_19578,N_19190);
or U20545 (N_20545,N_19971,N_19013);
xnor U20546 (N_20546,N_19857,N_19777);
nor U20547 (N_20547,N_19302,N_19314);
and U20548 (N_20548,N_19139,N_19202);
and U20549 (N_20549,N_19954,N_19463);
and U20550 (N_20550,N_19044,N_19658);
nor U20551 (N_20551,N_19767,N_19466);
or U20552 (N_20552,N_19037,N_19571);
nor U20553 (N_20553,N_19904,N_19146);
or U20554 (N_20554,N_19598,N_19889);
and U20555 (N_20555,N_19510,N_19598);
and U20556 (N_20556,N_19656,N_19443);
xor U20557 (N_20557,N_19340,N_19428);
nand U20558 (N_20558,N_19095,N_19617);
and U20559 (N_20559,N_19225,N_19382);
nand U20560 (N_20560,N_19324,N_19285);
xor U20561 (N_20561,N_19368,N_19531);
and U20562 (N_20562,N_19731,N_19805);
and U20563 (N_20563,N_19313,N_19209);
xnor U20564 (N_20564,N_19910,N_19109);
nand U20565 (N_20565,N_19260,N_19114);
xnor U20566 (N_20566,N_19620,N_19976);
xnor U20567 (N_20567,N_19213,N_19680);
nand U20568 (N_20568,N_19521,N_19538);
and U20569 (N_20569,N_19209,N_19686);
nor U20570 (N_20570,N_19798,N_19894);
xor U20571 (N_20571,N_19868,N_19508);
nand U20572 (N_20572,N_19439,N_19758);
nand U20573 (N_20573,N_19364,N_19763);
and U20574 (N_20574,N_19660,N_19460);
or U20575 (N_20575,N_19445,N_19634);
xnor U20576 (N_20576,N_19477,N_19320);
or U20577 (N_20577,N_19303,N_19359);
nor U20578 (N_20578,N_19636,N_19194);
or U20579 (N_20579,N_19048,N_19230);
or U20580 (N_20580,N_19735,N_19715);
nor U20581 (N_20581,N_19712,N_19835);
nand U20582 (N_20582,N_19195,N_19124);
and U20583 (N_20583,N_19129,N_19943);
xnor U20584 (N_20584,N_19452,N_19715);
nor U20585 (N_20585,N_19736,N_19002);
and U20586 (N_20586,N_19696,N_19112);
and U20587 (N_20587,N_19007,N_19094);
nand U20588 (N_20588,N_19433,N_19952);
nand U20589 (N_20589,N_19865,N_19102);
nand U20590 (N_20590,N_19323,N_19001);
nand U20591 (N_20591,N_19817,N_19961);
nor U20592 (N_20592,N_19258,N_19156);
and U20593 (N_20593,N_19927,N_19240);
nand U20594 (N_20594,N_19529,N_19698);
and U20595 (N_20595,N_19491,N_19139);
or U20596 (N_20596,N_19533,N_19641);
nor U20597 (N_20597,N_19493,N_19376);
nand U20598 (N_20598,N_19225,N_19525);
nor U20599 (N_20599,N_19756,N_19103);
or U20600 (N_20600,N_19298,N_19455);
and U20601 (N_20601,N_19308,N_19650);
or U20602 (N_20602,N_19365,N_19640);
nand U20603 (N_20603,N_19192,N_19954);
nor U20604 (N_20604,N_19648,N_19435);
and U20605 (N_20605,N_19509,N_19367);
nand U20606 (N_20606,N_19765,N_19979);
or U20607 (N_20607,N_19650,N_19490);
or U20608 (N_20608,N_19657,N_19709);
xnor U20609 (N_20609,N_19068,N_19943);
nor U20610 (N_20610,N_19315,N_19066);
nor U20611 (N_20611,N_19308,N_19679);
xor U20612 (N_20612,N_19912,N_19368);
nand U20613 (N_20613,N_19995,N_19119);
nor U20614 (N_20614,N_19855,N_19853);
xnor U20615 (N_20615,N_19504,N_19880);
nor U20616 (N_20616,N_19508,N_19281);
and U20617 (N_20617,N_19099,N_19660);
or U20618 (N_20618,N_19142,N_19572);
or U20619 (N_20619,N_19295,N_19829);
or U20620 (N_20620,N_19405,N_19622);
and U20621 (N_20621,N_19322,N_19815);
and U20622 (N_20622,N_19466,N_19440);
and U20623 (N_20623,N_19282,N_19591);
or U20624 (N_20624,N_19074,N_19266);
xor U20625 (N_20625,N_19066,N_19877);
nor U20626 (N_20626,N_19019,N_19898);
or U20627 (N_20627,N_19920,N_19139);
and U20628 (N_20628,N_19336,N_19079);
nor U20629 (N_20629,N_19519,N_19632);
nand U20630 (N_20630,N_19874,N_19284);
nand U20631 (N_20631,N_19245,N_19023);
nand U20632 (N_20632,N_19014,N_19831);
xnor U20633 (N_20633,N_19234,N_19937);
or U20634 (N_20634,N_19506,N_19322);
and U20635 (N_20635,N_19435,N_19977);
nand U20636 (N_20636,N_19790,N_19429);
xnor U20637 (N_20637,N_19465,N_19512);
and U20638 (N_20638,N_19711,N_19401);
xor U20639 (N_20639,N_19810,N_19947);
nand U20640 (N_20640,N_19768,N_19998);
xnor U20641 (N_20641,N_19049,N_19721);
nor U20642 (N_20642,N_19518,N_19646);
or U20643 (N_20643,N_19633,N_19681);
nand U20644 (N_20644,N_19477,N_19003);
nor U20645 (N_20645,N_19492,N_19854);
nand U20646 (N_20646,N_19752,N_19587);
nor U20647 (N_20647,N_19938,N_19245);
xnor U20648 (N_20648,N_19651,N_19975);
nand U20649 (N_20649,N_19389,N_19416);
and U20650 (N_20650,N_19716,N_19226);
xnor U20651 (N_20651,N_19037,N_19641);
or U20652 (N_20652,N_19524,N_19822);
nand U20653 (N_20653,N_19602,N_19399);
nand U20654 (N_20654,N_19235,N_19152);
and U20655 (N_20655,N_19442,N_19049);
or U20656 (N_20656,N_19018,N_19127);
nor U20657 (N_20657,N_19236,N_19251);
xnor U20658 (N_20658,N_19044,N_19598);
nor U20659 (N_20659,N_19363,N_19639);
or U20660 (N_20660,N_19847,N_19299);
nor U20661 (N_20661,N_19768,N_19302);
and U20662 (N_20662,N_19416,N_19901);
and U20663 (N_20663,N_19884,N_19343);
nor U20664 (N_20664,N_19372,N_19778);
and U20665 (N_20665,N_19898,N_19968);
nand U20666 (N_20666,N_19081,N_19391);
nand U20667 (N_20667,N_19265,N_19165);
or U20668 (N_20668,N_19432,N_19706);
nor U20669 (N_20669,N_19176,N_19160);
xnor U20670 (N_20670,N_19210,N_19278);
nand U20671 (N_20671,N_19705,N_19413);
and U20672 (N_20672,N_19226,N_19742);
or U20673 (N_20673,N_19271,N_19957);
or U20674 (N_20674,N_19215,N_19635);
xor U20675 (N_20675,N_19487,N_19307);
xnor U20676 (N_20676,N_19182,N_19838);
xor U20677 (N_20677,N_19949,N_19298);
xor U20678 (N_20678,N_19424,N_19510);
xor U20679 (N_20679,N_19706,N_19536);
xnor U20680 (N_20680,N_19909,N_19772);
xor U20681 (N_20681,N_19196,N_19432);
xnor U20682 (N_20682,N_19647,N_19192);
or U20683 (N_20683,N_19940,N_19178);
nor U20684 (N_20684,N_19709,N_19865);
xor U20685 (N_20685,N_19172,N_19037);
nand U20686 (N_20686,N_19195,N_19779);
xor U20687 (N_20687,N_19636,N_19490);
nand U20688 (N_20688,N_19525,N_19075);
nand U20689 (N_20689,N_19171,N_19056);
xnor U20690 (N_20690,N_19668,N_19099);
or U20691 (N_20691,N_19349,N_19287);
or U20692 (N_20692,N_19058,N_19476);
nand U20693 (N_20693,N_19571,N_19149);
nor U20694 (N_20694,N_19660,N_19820);
nor U20695 (N_20695,N_19714,N_19872);
or U20696 (N_20696,N_19775,N_19450);
or U20697 (N_20697,N_19703,N_19642);
and U20698 (N_20698,N_19293,N_19329);
nor U20699 (N_20699,N_19000,N_19728);
and U20700 (N_20700,N_19541,N_19335);
xnor U20701 (N_20701,N_19256,N_19868);
nor U20702 (N_20702,N_19817,N_19545);
nand U20703 (N_20703,N_19030,N_19184);
and U20704 (N_20704,N_19290,N_19633);
xor U20705 (N_20705,N_19595,N_19185);
xnor U20706 (N_20706,N_19553,N_19889);
nand U20707 (N_20707,N_19012,N_19252);
or U20708 (N_20708,N_19675,N_19537);
xor U20709 (N_20709,N_19037,N_19907);
nand U20710 (N_20710,N_19850,N_19780);
nand U20711 (N_20711,N_19820,N_19316);
nor U20712 (N_20712,N_19354,N_19056);
nor U20713 (N_20713,N_19578,N_19335);
xor U20714 (N_20714,N_19599,N_19551);
or U20715 (N_20715,N_19428,N_19016);
or U20716 (N_20716,N_19643,N_19650);
and U20717 (N_20717,N_19624,N_19865);
and U20718 (N_20718,N_19304,N_19780);
or U20719 (N_20719,N_19748,N_19356);
nand U20720 (N_20720,N_19905,N_19095);
nand U20721 (N_20721,N_19090,N_19232);
nand U20722 (N_20722,N_19291,N_19041);
or U20723 (N_20723,N_19381,N_19654);
or U20724 (N_20724,N_19010,N_19135);
or U20725 (N_20725,N_19555,N_19560);
or U20726 (N_20726,N_19147,N_19201);
nor U20727 (N_20727,N_19406,N_19311);
xnor U20728 (N_20728,N_19139,N_19338);
nand U20729 (N_20729,N_19302,N_19738);
nand U20730 (N_20730,N_19865,N_19901);
xnor U20731 (N_20731,N_19427,N_19575);
nor U20732 (N_20732,N_19118,N_19655);
and U20733 (N_20733,N_19918,N_19310);
nand U20734 (N_20734,N_19265,N_19458);
and U20735 (N_20735,N_19394,N_19557);
xor U20736 (N_20736,N_19981,N_19725);
or U20737 (N_20737,N_19386,N_19271);
or U20738 (N_20738,N_19683,N_19092);
xnor U20739 (N_20739,N_19837,N_19692);
nand U20740 (N_20740,N_19577,N_19407);
and U20741 (N_20741,N_19422,N_19404);
xnor U20742 (N_20742,N_19430,N_19086);
nor U20743 (N_20743,N_19997,N_19389);
xnor U20744 (N_20744,N_19552,N_19741);
or U20745 (N_20745,N_19708,N_19153);
nand U20746 (N_20746,N_19351,N_19360);
nand U20747 (N_20747,N_19934,N_19886);
or U20748 (N_20748,N_19978,N_19472);
xor U20749 (N_20749,N_19616,N_19819);
or U20750 (N_20750,N_19182,N_19696);
xnor U20751 (N_20751,N_19301,N_19190);
or U20752 (N_20752,N_19473,N_19580);
xor U20753 (N_20753,N_19536,N_19926);
and U20754 (N_20754,N_19419,N_19849);
nor U20755 (N_20755,N_19930,N_19360);
nor U20756 (N_20756,N_19279,N_19696);
or U20757 (N_20757,N_19313,N_19595);
or U20758 (N_20758,N_19656,N_19652);
nand U20759 (N_20759,N_19713,N_19019);
nand U20760 (N_20760,N_19662,N_19765);
nor U20761 (N_20761,N_19053,N_19543);
nand U20762 (N_20762,N_19274,N_19431);
xnor U20763 (N_20763,N_19154,N_19068);
nand U20764 (N_20764,N_19942,N_19873);
or U20765 (N_20765,N_19551,N_19920);
nor U20766 (N_20766,N_19675,N_19575);
and U20767 (N_20767,N_19819,N_19768);
nor U20768 (N_20768,N_19025,N_19987);
nand U20769 (N_20769,N_19261,N_19320);
or U20770 (N_20770,N_19802,N_19523);
or U20771 (N_20771,N_19462,N_19458);
and U20772 (N_20772,N_19979,N_19668);
nand U20773 (N_20773,N_19922,N_19811);
nor U20774 (N_20774,N_19430,N_19555);
nand U20775 (N_20775,N_19576,N_19736);
and U20776 (N_20776,N_19854,N_19878);
xor U20777 (N_20777,N_19815,N_19617);
xor U20778 (N_20778,N_19721,N_19477);
and U20779 (N_20779,N_19149,N_19772);
or U20780 (N_20780,N_19482,N_19899);
xnor U20781 (N_20781,N_19540,N_19017);
nor U20782 (N_20782,N_19180,N_19377);
or U20783 (N_20783,N_19927,N_19339);
and U20784 (N_20784,N_19020,N_19793);
or U20785 (N_20785,N_19881,N_19708);
or U20786 (N_20786,N_19622,N_19447);
and U20787 (N_20787,N_19717,N_19028);
nor U20788 (N_20788,N_19727,N_19375);
nor U20789 (N_20789,N_19783,N_19725);
nand U20790 (N_20790,N_19425,N_19537);
xor U20791 (N_20791,N_19884,N_19586);
nand U20792 (N_20792,N_19759,N_19464);
nor U20793 (N_20793,N_19947,N_19194);
or U20794 (N_20794,N_19304,N_19876);
or U20795 (N_20795,N_19674,N_19970);
and U20796 (N_20796,N_19209,N_19288);
or U20797 (N_20797,N_19027,N_19329);
or U20798 (N_20798,N_19368,N_19618);
and U20799 (N_20799,N_19456,N_19030);
or U20800 (N_20800,N_19704,N_19534);
nor U20801 (N_20801,N_19398,N_19801);
or U20802 (N_20802,N_19200,N_19683);
nor U20803 (N_20803,N_19455,N_19040);
xor U20804 (N_20804,N_19814,N_19397);
xnor U20805 (N_20805,N_19665,N_19486);
and U20806 (N_20806,N_19433,N_19370);
and U20807 (N_20807,N_19629,N_19154);
and U20808 (N_20808,N_19337,N_19562);
nand U20809 (N_20809,N_19649,N_19090);
or U20810 (N_20810,N_19846,N_19247);
xor U20811 (N_20811,N_19323,N_19176);
nand U20812 (N_20812,N_19298,N_19796);
nand U20813 (N_20813,N_19460,N_19972);
and U20814 (N_20814,N_19282,N_19361);
nor U20815 (N_20815,N_19337,N_19388);
nor U20816 (N_20816,N_19237,N_19956);
and U20817 (N_20817,N_19088,N_19737);
and U20818 (N_20818,N_19443,N_19823);
nor U20819 (N_20819,N_19235,N_19354);
nor U20820 (N_20820,N_19419,N_19956);
xor U20821 (N_20821,N_19887,N_19306);
xor U20822 (N_20822,N_19061,N_19854);
xnor U20823 (N_20823,N_19135,N_19308);
xnor U20824 (N_20824,N_19086,N_19524);
and U20825 (N_20825,N_19657,N_19853);
nor U20826 (N_20826,N_19614,N_19503);
or U20827 (N_20827,N_19079,N_19903);
nor U20828 (N_20828,N_19063,N_19433);
nand U20829 (N_20829,N_19833,N_19335);
and U20830 (N_20830,N_19708,N_19336);
and U20831 (N_20831,N_19606,N_19865);
or U20832 (N_20832,N_19618,N_19041);
nand U20833 (N_20833,N_19062,N_19186);
and U20834 (N_20834,N_19070,N_19096);
nand U20835 (N_20835,N_19918,N_19382);
xnor U20836 (N_20836,N_19860,N_19732);
nor U20837 (N_20837,N_19190,N_19511);
xor U20838 (N_20838,N_19180,N_19304);
and U20839 (N_20839,N_19666,N_19927);
or U20840 (N_20840,N_19114,N_19224);
and U20841 (N_20841,N_19788,N_19901);
nor U20842 (N_20842,N_19706,N_19832);
and U20843 (N_20843,N_19246,N_19076);
nor U20844 (N_20844,N_19516,N_19433);
xnor U20845 (N_20845,N_19058,N_19192);
nand U20846 (N_20846,N_19724,N_19090);
nor U20847 (N_20847,N_19142,N_19586);
or U20848 (N_20848,N_19289,N_19865);
xnor U20849 (N_20849,N_19351,N_19753);
xnor U20850 (N_20850,N_19699,N_19470);
xnor U20851 (N_20851,N_19027,N_19442);
or U20852 (N_20852,N_19717,N_19930);
xor U20853 (N_20853,N_19875,N_19860);
nand U20854 (N_20854,N_19636,N_19145);
nor U20855 (N_20855,N_19118,N_19791);
xor U20856 (N_20856,N_19084,N_19087);
or U20857 (N_20857,N_19763,N_19745);
xnor U20858 (N_20858,N_19946,N_19511);
or U20859 (N_20859,N_19825,N_19972);
xnor U20860 (N_20860,N_19579,N_19506);
or U20861 (N_20861,N_19717,N_19938);
nor U20862 (N_20862,N_19397,N_19301);
nor U20863 (N_20863,N_19513,N_19502);
and U20864 (N_20864,N_19097,N_19417);
nor U20865 (N_20865,N_19719,N_19697);
and U20866 (N_20866,N_19965,N_19633);
and U20867 (N_20867,N_19988,N_19864);
nor U20868 (N_20868,N_19650,N_19818);
nor U20869 (N_20869,N_19167,N_19328);
xnor U20870 (N_20870,N_19690,N_19199);
xnor U20871 (N_20871,N_19977,N_19233);
xor U20872 (N_20872,N_19368,N_19432);
nand U20873 (N_20873,N_19633,N_19687);
nand U20874 (N_20874,N_19902,N_19917);
or U20875 (N_20875,N_19379,N_19020);
and U20876 (N_20876,N_19456,N_19025);
and U20877 (N_20877,N_19473,N_19954);
or U20878 (N_20878,N_19316,N_19182);
xor U20879 (N_20879,N_19188,N_19602);
xnor U20880 (N_20880,N_19111,N_19607);
xor U20881 (N_20881,N_19562,N_19850);
nor U20882 (N_20882,N_19947,N_19236);
and U20883 (N_20883,N_19109,N_19331);
nand U20884 (N_20884,N_19379,N_19745);
nand U20885 (N_20885,N_19139,N_19553);
xor U20886 (N_20886,N_19276,N_19290);
or U20887 (N_20887,N_19644,N_19047);
nor U20888 (N_20888,N_19524,N_19607);
and U20889 (N_20889,N_19478,N_19068);
or U20890 (N_20890,N_19271,N_19330);
xnor U20891 (N_20891,N_19443,N_19769);
nor U20892 (N_20892,N_19036,N_19424);
or U20893 (N_20893,N_19631,N_19512);
nand U20894 (N_20894,N_19907,N_19134);
and U20895 (N_20895,N_19184,N_19975);
and U20896 (N_20896,N_19119,N_19306);
and U20897 (N_20897,N_19658,N_19097);
nor U20898 (N_20898,N_19113,N_19472);
xor U20899 (N_20899,N_19872,N_19442);
xnor U20900 (N_20900,N_19555,N_19978);
xor U20901 (N_20901,N_19902,N_19840);
xnor U20902 (N_20902,N_19294,N_19534);
nand U20903 (N_20903,N_19581,N_19133);
xor U20904 (N_20904,N_19935,N_19008);
nor U20905 (N_20905,N_19787,N_19797);
or U20906 (N_20906,N_19635,N_19801);
nor U20907 (N_20907,N_19225,N_19582);
and U20908 (N_20908,N_19112,N_19999);
nand U20909 (N_20909,N_19499,N_19514);
nor U20910 (N_20910,N_19192,N_19681);
nand U20911 (N_20911,N_19251,N_19399);
nand U20912 (N_20912,N_19671,N_19524);
or U20913 (N_20913,N_19166,N_19131);
or U20914 (N_20914,N_19951,N_19223);
or U20915 (N_20915,N_19738,N_19650);
or U20916 (N_20916,N_19846,N_19723);
xnor U20917 (N_20917,N_19642,N_19434);
nor U20918 (N_20918,N_19206,N_19912);
nor U20919 (N_20919,N_19298,N_19592);
and U20920 (N_20920,N_19327,N_19381);
xor U20921 (N_20921,N_19714,N_19823);
nand U20922 (N_20922,N_19817,N_19605);
nand U20923 (N_20923,N_19742,N_19597);
nor U20924 (N_20924,N_19338,N_19782);
nor U20925 (N_20925,N_19164,N_19651);
nand U20926 (N_20926,N_19285,N_19960);
xor U20927 (N_20927,N_19425,N_19928);
or U20928 (N_20928,N_19097,N_19319);
nor U20929 (N_20929,N_19669,N_19588);
nor U20930 (N_20930,N_19988,N_19285);
and U20931 (N_20931,N_19690,N_19980);
nand U20932 (N_20932,N_19887,N_19355);
and U20933 (N_20933,N_19626,N_19127);
or U20934 (N_20934,N_19102,N_19501);
nor U20935 (N_20935,N_19419,N_19137);
nor U20936 (N_20936,N_19263,N_19350);
nand U20937 (N_20937,N_19448,N_19359);
nand U20938 (N_20938,N_19309,N_19920);
xnor U20939 (N_20939,N_19529,N_19418);
nor U20940 (N_20940,N_19319,N_19804);
xnor U20941 (N_20941,N_19401,N_19850);
xnor U20942 (N_20942,N_19374,N_19320);
nand U20943 (N_20943,N_19644,N_19871);
or U20944 (N_20944,N_19763,N_19411);
nor U20945 (N_20945,N_19039,N_19646);
xor U20946 (N_20946,N_19460,N_19973);
xnor U20947 (N_20947,N_19490,N_19718);
and U20948 (N_20948,N_19636,N_19724);
and U20949 (N_20949,N_19692,N_19694);
nand U20950 (N_20950,N_19906,N_19590);
nand U20951 (N_20951,N_19867,N_19612);
xnor U20952 (N_20952,N_19704,N_19093);
nand U20953 (N_20953,N_19696,N_19145);
nand U20954 (N_20954,N_19088,N_19643);
nor U20955 (N_20955,N_19712,N_19753);
and U20956 (N_20956,N_19902,N_19963);
xor U20957 (N_20957,N_19877,N_19869);
nor U20958 (N_20958,N_19450,N_19680);
and U20959 (N_20959,N_19070,N_19630);
or U20960 (N_20960,N_19433,N_19870);
xnor U20961 (N_20961,N_19815,N_19611);
or U20962 (N_20962,N_19736,N_19849);
and U20963 (N_20963,N_19690,N_19681);
or U20964 (N_20964,N_19759,N_19085);
xor U20965 (N_20965,N_19575,N_19691);
nand U20966 (N_20966,N_19264,N_19056);
nor U20967 (N_20967,N_19055,N_19375);
or U20968 (N_20968,N_19610,N_19268);
or U20969 (N_20969,N_19889,N_19961);
nand U20970 (N_20970,N_19643,N_19281);
nand U20971 (N_20971,N_19336,N_19662);
or U20972 (N_20972,N_19230,N_19122);
or U20973 (N_20973,N_19485,N_19114);
nand U20974 (N_20974,N_19447,N_19124);
nor U20975 (N_20975,N_19897,N_19417);
nor U20976 (N_20976,N_19443,N_19009);
xnor U20977 (N_20977,N_19942,N_19120);
xnor U20978 (N_20978,N_19187,N_19864);
nor U20979 (N_20979,N_19690,N_19817);
and U20980 (N_20980,N_19726,N_19137);
nor U20981 (N_20981,N_19032,N_19377);
nor U20982 (N_20982,N_19630,N_19269);
or U20983 (N_20983,N_19547,N_19185);
or U20984 (N_20984,N_19623,N_19639);
and U20985 (N_20985,N_19298,N_19625);
nand U20986 (N_20986,N_19631,N_19496);
nor U20987 (N_20987,N_19650,N_19829);
and U20988 (N_20988,N_19043,N_19333);
nor U20989 (N_20989,N_19490,N_19443);
xor U20990 (N_20990,N_19694,N_19102);
nor U20991 (N_20991,N_19770,N_19283);
xor U20992 (N_20992,N_19267,N_19668);
nand U20993 (N_20993,N_19370,N_19344);
nand U20994 (N_20994,N_19902,N_19266);
nand U20995 (N_20995,N_19798,N_19242);
xnor U20996 (N_20996,N_19262,N_19939);
nor U20997 (N_20997,N_19524,N_19761);
or U20998 (N_20998,N_19619,N_19511);
nor U20999 (N_20999,N_19829,N_19016);
and U21000 (N_21000,N_20542,N_20718);
nor U21001 (N_21001,N_20702,N_20637);
nand U21002 (N_21002,N_20316,N_20011);
nor U21003 (N_21003,N_20684,N_20783);
nor U21004 (N_21004,N_20974,N_20601);
xnor U21005 (N_21005,N_20680,N_20977);
or U21006 (N_21006,N_20227,N_20144);
and U21007 (N_21007,N_20916,N_20234);
or U21008 (N_21008,N_20930,N_20108);
or U21009 (N_21009,N_20388,N_20228);
nand U21010 (N_21010,N_20931,N_20806);
or U21011 (N_21011,N_20247,N_20477);
xor U21012 (N_21012,N_20310,N_20107);
nor U21013 (N_21013,N_20958,N_20179);
nor U21014 (N_21014,N_20088,N_20696);
or U21015 (N_21015,N_20733,N_20431);
nor U21016 (N_21016,N_20466,N_20889);
and U21017 (N_21017,N_20219,N_20877);
xnor U21018 (N_21018,N_20404,N_20315);
xor U21019 (N_21019,N_20762,N_20985);
nor U21020 (N_21020,N_20638,N_20997);
and U21021 (N_21021,N_20043,N_20933);
xnor U21022 (N_21022,N_20541,N_20288);
or U21023 (N_21023,N_20087,N_20306);
or U21024 (N_21024,N_20355,N_20722);
or U21025 (N_21025,N_20941,N_20617);
xor U21026 (N_21026,N_20505,N_20325);
xor U21027 (N_21027,N_20176,N_20128);
or U21028 (N_21028,N_20482,N_20990);
or U21029 (N_21029,N_20553,N_20622);
xnor U21030 (N_21030,N_20309,N_20821);
xnor U21031 (N_21031,N_20459,N_20465);
nand U21032 (N_21032,N_20546,N_20585);
and U21033 (N_21033,N_20472,N_20221);
xor U21034 (N_21034,N_20236,N_20999);
and U21035 (N_21035,N_20616,N_20868);
nor U21036 (N_21036,N_20249,N_20803);
and U21037 (N_21037,N_20788,N_20293);
and U21038 (N_21038,N_20470,N_20863);
and U21039 (N_21039,N_20526,N_20818);
xnor U21040 (N_21040,N_20345,N_20023);
nand U21041 (N_21041,N_20858,N_20017);
nand U21042 (N_21042,N_20403,N_20887);
xor U21043 (N_21043,N_20343,N_20149);
xnor U21044 (N_21044,N_20346,N_20327);
nor U21045 (N_21045,N_20586,N_20436);
or U21046 (N_21046,N_20678,N_20137);
and U21047 (N_21047,N_20556,N_20486);
nor U21048 (N_21048,N_20802,N_20516);
nand U21049 (N_21049,N_20847,N_20708);
and U21050 (N_21050,N_20199,N_20256);
xnor U21051 (N_21051,N_20218,N_20625);
or U21052 (N_21052,N_20611,N_20357);
and U21053 (N_21053,N_20194,N_20822);
xnor U21054 (N_21054,N_20870,N_20648);
nand U21055 (N_21055,N_20152,N_20523);
nor U21056 (N_21056,N_20569,N_20753);
nor U21057 (N_21057,N_20304,N_20740);
xnor U21058 (N_21058,N_20575,N_20039);
nand U21059 (N_21059,N_20591,N_20350);
and U21060 (N_21060,N_20214,N_20857);
and U21061 (N_21061,N_20848,N_20447);
nand U21062 (N_21062,N_20905,N_20947);
xnor U21063 (N_21063,N_20410,N_20675);
xor U21064 (N_21064,N_20850,N_20534);
nor U21065 (N_21065,N_20353,N_20914);
xnor U21066 (N_21066,N_20281,N_20764);
nor U21067 (N_21067,N_20506,N_20994);
nor U21068 (N_21068,N_20370,N_20484);
nor U21069 (N_21069,N_20051,N_20628);
or U21070 (N_21070,N_20499,N_20792);
nand U21071 (N_21071,N_20957,N_20864);
nand U21072 (N_21072,N_20965,N_20473);
or U21073 (N_21073,N_20102,N_20837);
nor U21074 (N_21074,N_20250,N_20824);
nand U21075 (N_21075,N_20169,N_20763);
xor U21076 (N_21076,N_20339,N_20492);
nand U21077 (N_21077,N_20070,N_20125);
xor U21078 (N_21078,N_20369,N_20799);
xor U21079 (N_21079,N_20001,N_20418);
xor U21080 (N_21080,N_20592,N_20709);
and U21081 (N_21081,N_20642,N_20462);
xor U21082 (N_21082,N_20026,N_20552);
or U21083 (N_21083,N_20437,N_20226);
nand U21084 (N_21084,N_20254,N_20147);
nor U21085 (N_21085,N_20402,N_20082);
nor U21086 (N_21086,N_20421,N_20823);
or U21087 (N_21087,N_20768,N_20291);
xor U21088 (N_21088,N_20987,N_20098);
and U21089 (N_21089,N_20111,N_20307);
xnor U21090 (N_21090,N_20399,N_20121);
and U21091 (N_21091,N_20422,N_20992);
nor U21092 (N_21092,N_20498,N_20723);
nor U21093 (N_21093,N_20564,N_20903);
and U21094 (N_21094,N_20779,N_20649);
nor U21095 (N_21095,N_20430,N_20314);
xor U21096 (N_21096,N_20123,N_20861);
or U21097 (N_21097,N_20183,N_20319);
xnor U21098 (N_21098,N_20576,N_20652);
xnor U21099 (N_21099,N_20804,N_20699);
and U21100 (N_21100,N_20342,N_20513);
or U21101 (N_21101,N_20973,N_20311);
and U21102 (N_21102,N_20298,N_20452);
nor U21103 (N_21103,N_20873,N_20368);
and U21104 (N_21104,N_20392,N_20561);
nor U21105 (N_21105,N_20756,N_20908);
nor U21106 (N_21106,N_20106,N_20366);
or U21107 (N_21107,N_20519,N_20248);
nor U21108 (N_21108,N_20720,N_20529);
nand U21109 (N_21109,N_20295,N_20998);
or U21110 (N_21110,N_20690,N_20805);
nor U21111 (N_21111,N_20025,N_20324);
nand U21112 (N_21112,N_20002,N_20225);
nor U21113 (N_21113,N_20165,N_20765);
or U21114 (N_21114,N_20501,N_20798);
and U21115 (N_21115,N_20911,N_20487);
xnor U21116 (N_21116,N_20015,N_20196);
and U21117 (N_21117,N_20009,N_20099);
nand U21118 (N_21118,N_20193,N_20323);
nor U21119 (N_21119,N_20464,N_20520);
nor U21120 (N_21120,N_20286,N_20886);
or U21121 (N_21121,N_20174,N_20010);
nand U21122 (N_21122,N_20361,N_20441);
nand U21123 (N_21123,N_20728,N_20476);
or U21124 (N_21124,N_20621,N_20145);
xnor U21125 (N_21125,N_20782,N_20915);
or U21126 (N_21126,N_20683,N_20831);
nor U21127 (N_21127,N_20273,N_20047);
or U21128 (N_21128,N_20049,N_20117);
xor U21129 (N_21129,N_20660,N_20597);
and U21130 (N_21130,N_20712,N_20351);
or U21131 (N_21131,N_20817,N_20830);
or U21132 (N_21132,N_20742,N_20540);
nor U21133 (N_21133,N_20984,N_20434);
nor U21134 (N_21134,N_20217,N_20953);
nand U21135 (N_21135,N_20521,N_20747);
nand U21136 (N_21136,N_20587,N_20890);
or U21137 (N_21137,N_20500,N_20262);
or U21138 (N_21138,N_20277,N_20632);
or U21139 (N_21139,N_20926,N_20938);
xor U21140 (N_21140,N_20725,N_20394);
and U21141 (N_21141,N_20003,N_20919);
xnor U21142 (N_21142,N_20548,N_20135);
nor U21143 (N_21143,N_20420,N_20963);
nand U21144 (N_21144,N_20906,N_20185);
xor U21145 (N_21145,N_20734,N_20608);
nor U21146 (N_21146,N_20489,N_20882);
nor U21147 (N_21147,N_20807,N_20643);
nor U21148 (N_21148,N_20239,N_20400);
xnor U21149 (N_21149,N_20016,N_20153);
or U21150 (N_21150,N_20703,N_20260);
and U21151 (N_21151,N_20669,N_20457);
nor U21152 (N_21152,N_20800,N_20922);
xnor U21153 (N_21153,N_20860,N_20014);
nand U21154 (N_21154,N_20533,N_20000);
or U21155 (N_21155,N_20253,N_20257);
nor U21156 (N_21156,N_20382,N_20697);
nor U21157 (N_21157,N_20766,N_20606);
and U21158 (N_21158,N_20920,N_20859);
nand U21159 (N_21159,N_20639,N_20425);
and U21160 (N_21160,N_20503,N_20545);
nor U21161 (N_21161,N_20381,N_20896);
or U21162 (N_21162,N_20651,N_20579);
nand U21163 (N_21163,N_20409,N_20220);
and U21164 (N_21164,N_20810,N_20613);
or U21165 (N_21165,N_20849,N_20899);
nand U21166 (N_21166,N_20633,N_20666);
and U21167 (N_21167,N_20707,N_20738);
or U21168 (N_21168,N_20655,N_20808);
nand U21169 (N_21169,N_20897,N_20384);
nor U21170 (N_21170,N_20417,N_20727);
nand U21171 (N_21171,N_20761,N_20892);
nor U21172 (N_21172,N_20093,N_20146);
nor U21173 (N_21173,N_20395,N_20950);
or U21174 (N_21174,N_20875,N_20955);
and U21175 (N_21175,N_20332,N_20274);
and U21176 (N_21176,N_20757,N_20695);
and U21177 (N_21177,N_20423,N_20432);
xnor U21178 (N_21178,N_20453,N_20658);
nor U21179 (N_21179,N_20184,N_20245);
nand U21180 (N_21180,N_20936,N_20347);
xnor U21181 (N_21181,N_20175,N_20211);
nor U21182 (N_21182,N_20558,N_20318);
xor U21183 (N_21183,N_20944,N_20203);
nor U21184 (N_21184,N_20018,N_20834);
xnor U21185 (N_21185,N_20312,N_20913);
xnor U21186 (N_21186,N_20191,N_20960);
and U21187 (N_21187,N_20907,N_20044);
nand U21188 (N_21188,N_20110,N_20134);
and U21189 (N_21189,N_20485,N_20940);
xor U21190 (N_21190,N_20893,N_20888);
or U21191 (N_21191,N_20789,N_20054);
or U21192 (N_21192,N_20004,N_20910);
nand U21193 (N_21193,N_20571,N_20209);
xor U21194 (N_21194,N_20598,N_20854);
xor U21195 (N_21195,N_20636,N_20538);
and U21196 (N_21196,N_20746,N_20917);
nand U21197 (N_21197,N_20580,N_20966);
nor U21198 (N_21198,N_20356,N_20901);
xnor U21199 (N_21199,N_20630,N_20334);
xnor U21200 (N_21200,N_20451,N_20775);
nand U21201 (N_21201,N_20590,N_20924);
xnor U21202 (N_21202,N_20689,N_20692);
and U21203 (N_21203,N_20150,N_20737);
nand U21204 (N_21204,N_20401,N_20237);
and U21205 (N_21205,N_20034,N_20371);
nor U21206 (N_21206,N_20701,N_20216);
nor U21207 (N_21207,N_20641,N_20988);
or U21208 (N_21208,N_20204,N_20059);
nand U21209 (N_21209,N_20035,N_20020);
and U21210 (N_21210,N_20839,N_20036);
nand U21211 (N_21211,N_20340,N_20898);
or U21212 (N_21212,N_20657,N_20101);
nand U21213 (N_21213,N_20488,N_20030);
xor U21214 (N_21214,N_20233,N_20584);
nand U21215 (N_21215,N_20092,N_20359);
or U21216 (N_21216,N_20405,N_20267);
nor U21217 (N_21217,N_20943,N_20467);
nand U21218 (N_21218,N_20749,N_20284);
nand U21219 (N_21219,N_20066,N_20397);
nor U21220 (N_21220,N_20507,N_20682);
nand U21221 (N_21221,N_20141,N_20089);
nor U21222 (N_21222,N_20952,N_20038);
nor U21223 (N_21223,N_20058,N_20856);
nand U21224 (N_21224,N_20544,N_20222);
or U21225 (N_21225,N_20158,N_20653);
nand U21226 (N_21226,N_20212,N_20321);
or U21227 (N_21227,N_20168,N_20445);
nor U21228 (N_21228,N_20385,N_20440);
nor U21229 (N_21229,N_20365,N_20378);
or U21230 (N_21230,N_20661,N_20724);
or U21231 (N_21231,N_20177,N_20739);
nor U21232 (N_21232,N_20674,N_20069);
and U21233 (N_21233,N_20570,N_20627);
nor U21234 (N_21234,N_20681,N_20713);
and U21235 (N_21235,N_20308,N_20180);
and U21236 (N_21236,N_20978,N_20448);
and U21237 (N_21237,N_20894,N_20959);
nand U21238 (N_21238,N_20603,N_20372);
xor U21239 (N_21239,N_20995,N_20045);
xor U21240 (N_21240,N_20289,N_20776);
and U21241 (N_21241,N_20354,N_20640);
and U21242 (N_21242,N_20474,N_20543);
and U21243 (N_21243,N_20527,N_20600);
xor U21244 (N_21244,N_20008,N_20454);
or U21245 (N_21245,N_20170,N_20055);
xor U21246 (N_21246,N_20964,N_20155);
nand U21247 (N_21247,N_20969,N_20411);
xor U21248 (N_21248,N_20406,N_20925);
xnor U21249 (N_21249,N_20968,N_20238);
and U21250 (N_21250,N_20232,N_20280);
and U21251 (N_21251,N_20126,N_20075);
nor U21252 (N_21252,N_20942,N_20700);
nand U21253 (N_21253,N_20444,N_20171);
nand U21254 (N_21254,N_20634,N_20563);
or U21255 (N_21255,N_20255,N_20412);
nand U21256 (N_21256,N_20829,N_20103);
xor U21257 (N_21257,N_20794,N_20872);
xnor U21258 (N_21258,N_20945,N_20079);
nand U21259 (N_21259,N_20261,N_20362);
nor U21260 (N_21260,N_20131,N_20647);
nand U21261 (N_21261,N_20605,N_20843);
and U21262 (N_21262,N_20483,N_20080);
xnor U21263 (N_21263,N_20027,N_20113);
nand U21264 (N_21264,N_20883,N_20084);
or U21265 (N_21265,N_20980,N_20156);
and U21266 (N_21266,N_20827,N_20816);
nand U21267 (N_21267,N_20317,N_20244);
xnor U21268 (N_21268,N_20844,N_20105);
xor U21269 (N_21269,N_20604,N_20754);
xor U21270 (N_21270,N_20292,N_20373);
and U21271 (N_21271,N_20567,N_20268);
xnor U21272 (N_21272,N_20909,N_20951);
nor U21273 (N_21273,N_20846,N_20918);
xor U21274 (N_21274,N_20793,N_20852);
nor U21275 (N_21275,N_20972,N_20932);
or U21276 (N_21276,N_20549,N_20554);
and U21277 (N_21277,N_20819,N_20900);
nand U21278 (N_21278,N_20706,N_20672);
and U21279 (N_21279,N_20522,N_20525);
and U21280 (N_21280,N_20568,N_20599);
nand U21281 (N_21281,N_20407,N_20202);
nand U21282 (N_21282,N_20299,N_20508);
xnor U21283 (N_21283,N_20230,N_20891);
and U21284 (N_21284,N_20364,N_20928);
nand U21285 (N_21285,N_20866,N_20352);
or U21286 (N_21286,N_20979,N_20996);
xnor U21287 (N_21287,N_20867,N_20537);
nand U21288 (N_21288,N_20455,N_20029);
nand U21289 (N_21289,N_20815,N_20282);
or U21290 (N_21290,N_20614,N_20704);
or U21291 (N_21291,N_20731,N_20668);
or U21292 (N_21292,N_20624,N_20265);
xor U21293 (N_21293,N_20842,N_20294);
or U21294 (N_21294,N_20266,N_20490);
xor U21295 (N_21295,N_20391,N_20333);
and U21296 (N_21296,N_20518,N_20743);
xor U21297 (N_21297,N_20021,N_20383);
or U21298 (N_21298,N_20832,N_20934);
and U21299 (N_21299,N_20715,N_20389);
nand U21300 (N_21300,N_20205,N_20290);
nor U21301 (N_21301,N_20297,N_20132);
or U21302 (N_21302,N_20428,N_20547);
xor U21303 (N_21303,N_20471,N_20456);
nand U21304 (N_21304,N_20278,N_20094);
or U21305 (N_21305,N_20338,N_20114);
and U21306 (N_21306,N_20885,N_20264);
and U21307 (N_21307,N_20744,N_20118);
nor U21308 (N_21308,N_20825,N_20755);
nand U21309 (N_21309,N_20083,N_20673);
and U21310 (N_21310,N_20157,N_20033);
or U21311 (N_21311,N_20659,N_20687);
nand U21312 (N_21312,N_20791,N_20670);
xor U21313 (N_21313,N_20797,N_20531);
or U21314 (N_21314,N_20677,N_20902);
nand U21315 (N_21315,N_20654,N_20935);
nor U21316 (N_21316,N_20005,N_20595);
or U21317 (N_21317,N_20172,N_20122);
nor U21318 (N_21318,N_20693,N_20646);
nor U21319 (N_21319,N_20296,N_20949);
nand U21320 (N_21320,N_20064,N_20574);
or U21321 (N_21321,N_20539,N_20679);
nor U21322 (N_21322,N_20215,N_20024);
or U21323 (N_21323,N_20182,N_20013);
and U21324 (N_21324,N_20735,N_20853);
nand U21325 (N_21325,N_20989,N_20811);
nor U21326 (N_21326,N_20050,N_20535);
xnor U21327 (N_21327,N_20186,N_20838);
or U21328 (N_21328,N_20429,N_20139);
nor U21329 (N_21329,N_20780,N_20777);
xor U21330 (N_21330,N_20062,N_20074);
nor U21331 (N_21331,N_20065,N_20159);
nor U21332 (N_21332,N_20190,N_20581);
and U21333 (N_21333,N_20491,N_20691);
nor U21334 (N_21334,N_20326,N_20077);
and U21335 (N_21335,N_20469,N_20986);
and U21336 (N_21336,N_20751,N_20833);
and U21337 (N_21337,N_20303,N_20167);
xnor U21338 (N_21338,N_20481,N_20192);
or U21339 (N_21339,N_20285,N_20588);
or U21340 (N_21340,N_20458,N_20210);
nor U21341 (N_21341,N_20865,N_20786);
or U21342 (N_21342,N_20698,N_20187);
nand U21343 (N_21343,N_20478,N_20337);
nor U21344 (N_21344,N_20130,N_20201);
nor U21345 (N_21345,N_20258,N_20688);
nor U21346 (N_21346,N_20726,N_20813);
nor U21347 (N_21347,N_20671,N_20609);
nand U21348 (N_21348,N_20981,N_20040);
nand U21349 (N_21349,N_20375,N_20729);
nand U21350 (N_21350,N_20551,N_20787);
nor U21351 (N_21351,N_20300,N_20479);
or U21352 (N_21352,N_20663,N_20577);
and U21353 (N_21353,N_20615,N_20302);
or U21354 (N_21354,N_20665,N_20716);
and U21355 (N_21355,N_20583,N_20927);
and U21356 (N_21356,N_20229,N_20136);
and U21357 (N_21357,N_20895,N_20970);
xor U21358 (N_21358,N_20714,N_20619);
or U21359 (N_21359,N_20532,N_20127);
nor U21360 (N_21360,N_20840,N_20120);
nand U21361 (N_21361,N_20468,N_20769);
or U21362 (N_21362,N_20450,N_20504);
or U21363 (N_21363,N_20904,N_20224);
nand U21364 (N_21364,N_20784,N_20251);
nor U21365 (N_21365,N_20097,N_20390);
or U21366 (N_21366,N_20862,N_20770);
or U21367 (N_21367,N_20667,N_20560);
or U21368 (N_21368,N_20785,N_20252);
and U21369 (N_21369,N_20528,N_20536);
xor U21370 (N_21370,N_20078,N_20962);
nand U21371 (N_21371,N_20085,N_20349);
or U21372 (N_21372,N_20869,N_20320);
nor U21373 (N_21373,N_20305,N_20090);
or U21374 (N_21374,N_20063,N_20975);
or U21375 (N_21375,N_20594,N_20279);
nor U21376 (N_21376,N_20645,N_20119);
nand U21377 (N_21377,N_20138,N_20424);
and U21378 (N_21378,N_20801,N_20387);
xor U21379 (N_21379,N_20644,N_20795);
nand U21380 (N_21380,N_20573,N_20610);
and U21381 (N_21381,N_20884,N_20376);
and U21382 (N_21382,N_20937,N_20496);
or U21383 (N_21383,N_20719,N_20662);
xor U21384 (N_21384,N_20511,N_20650);
xnor U21385 (N_21385,N_20578,N_20143);
nor U21386 (N_21386,N_20686,N_20160);
nand U21387 (N_21387,N_20773,N_20037);
nand U21388 (N_21388,N_20771,N_20912);
and U21389 (N_21389,N_20923,N_20475);
nand U21390 (N_21390,N_20096,N_20269);
nand U21391 (N_21391,N_20752,N_20328);
and U21392 (N_21392,N_20971,N_20426);
or U21393 (N_21393,N_20042,N_20348);
and U21394 (N_21394,N_20976,N_20946);
nand U21395 (N_21395,N_20263,N_20198);
xnor U21396 (N_21396,N_20480,N_20929);
xnor U21397 (N_21397,N_20961,N_20415);
and U21398 (N_21398,N_20393,N_20748);
nor U21399 (N_21399,N_20416,N_20855);
and U21400 (N_21400,N_20993,N_20438);
nand U21401 (N_21401,N_20335,N_20322);
nand U21402 (N_21402,N_20596,N_20517);
xnor U21403 (N_21403,N_20530,N_20344);
and U21404 (N_21404,N_20774,N_20705);
nor U21405 (N_21405,N_20112,N_20197);
xor U21406 (N_21406,N_20772,N_20732);
nor U21407 (N_21407,N_20367,N_20100);
nor U21408 (N_21408,N_20967,N_20664);
xnor U21409 (N_21409,N_20283,N_20515);
and U21410 (N_21410,N_20502,N_20271);
nand U21411 (N_21411,N_20052,N_20007);
nand U21412 (N_21412,N_20778,N_20874);
and U21413 (N_21413,N_20745,N_20142);
or U21414 (N_21414,N_20493,N_20151);
xnor U21415 (N_21415,N_20876,N_20276);
and U21416 (N_21416,N_20956,N_20259);
or U21417 (N_21417,N_20443,N_20717);
nand U21418 (N_21418,N_20685,N_20760);
or U21419 (N_21419,N_20566,N_20140);
nor U21420 (N_21420,N_20991,N_20240);
xor U21421 (N_21421,N_20494,N_20046);
and U21422 (N_21422,N_20270,N_20067);
nand U21423 (N_21423,N_20954,N_20759);
xnor U21424 (N_21424,N_20461,N_20386);
xnor U21425 (N_21425,N_20019,N_20061);
or U21426 (N_21426,N_20880,N_20790);
or U21427 (N_21427,N_20162,N_20828);
or U21428 (N_21428,N_20076,N_20374);
and U21429 (N_21429,N_20439,N_20329);
and U21430 (N_21430,N_20736,N_20056);
or U21431 (N_21431,N_20071,N_20730);
nand U21432 (N_21432,N_20331,N_20572);
or U21433 (N_21433,N_20178,N_20767);
nor U21434 (N_21434,N_20750,N_20032);
nand U21435 (N_21435,N_20053,N_20148);
xnor U21436 (N_21436,N_20208,N_20012);
and U21437 (N_21437,N_20781,N_20629);
and U21438 (N_21438,N_20091,N_20358);
and U21439 (N_21439,N_20243,N_20006);
or U21440 (N_21440,N_20095,N_20948);
nor U21441 (N_21441,N_20559,N_20495);
or U21442 (N_21442,N_20982,N_20509);
or U21443 (N_21443,N_20398,N_20656);
or U21444 (N_21444,N_20272,N_20275);
nand U21445 (N_21445,N_20195,N_20116);
nand U21446 (N_21446,N_20189,N_20433);
or U21447 (N_21447,N_20983,N_20301);
xnor U21448 (N_21448,N_20231,N_20631);
xor U21449 (N_21449,N_20435,N_20836);
or U21450 (N_21450,N_20360,N_20086);
or U21451 (N_21451,N_20820,N_20129);
and U21452 (N_21452,N_20620,N_20618);
or U21453 (N_21453,N_20826,N_20235);
and U21454 (N_21454,N_20626,N_20073);
xor U21455 (N_21455,N_20341,N_20427);
xnor U21456 (N_21456,N_20133,N_20741);
and U21457 (N_21457,N_20607,N_20022);
nor U21458 (N_21458,N_20242,N_20419);
nand U21459 (N_21459,N_20166,N_20593);
xor U21460 (N_21460,N_20081,N_20164);
nor U21461 (N_21461,N_20814,N_20602);
nand U21462 (N_21462,N_20057,N_20845);
or U21463 (N_21463,N_20060,N_20206);
nor U21464 (N_21464,N_20173,N_20188);
nor U21465 (N_21465,N_20246,N_20104);
or U21466 (N_21466,N_20835,N_20694);
nand U21467 (N_21467,N_20623,N_20200);
nand U21468 (N_21468,N_20881,N_20363);
or U21469 (N_21469,N_20414,N_20068);
xor U21470 (N_21470,N_20512,N_20565);
nand U21471 (N_21471,N_20161,N_20557);
and U21472 (N_21472,N_20241,N_20413);
nor U21473 (N_21473,N_20758,N_20207);
xor U21474 (N_21474,N_20871,N_20449);
nor U21475 (N_21475,N_20721,N_20676);
xnor U21476 (N_21476,N_20442,N_20446);
nor U21477 (N_21477,N_20796,N_20028);
or U21478 (N_21478,N_20379,N_20851);
xnor U21479 (N_21479,N_20048,N_20396);
or U21480 (N_21480,N_20287,N_20710);
and U21481 (N_21481,N_20181,N_20711);
xor U21482 (N_21482,N_20377,N_20812);
or U21483 (N_21483,N_20330,N_20510);
nand U21484 (N_21484,N_20313,N_20879);
or U21485 (N_21485,N_20115,N_20921);
nand U21486 (N_21486,N_20336,N_20072);
nor U21487 (N_21487,N_20109,N_20497);
or U21488 (N_21488,N_20939,N_20408);
and U21489 (N_21489,N_20809,N_20582);
xor U21490 (N_21490,N_20213,N_20562);
nor U21491 (N_21491,N_20154,N_20878);
nor U21492 (N_21492,N_20514,N_20524);
nand U21493 (N_21493,N_20124,N_20555);
nand U21494 (N_21494,N_20031,N_20589);
or U21495 (N_21495,N_20380,N_20041);
nand U21496 (N_21496,N_20550,N_20460);
nor U21497 (N_21497,N_20841,N_20635);
nand U21498 (N_21498,N_20612,N_20463);
and U21499 (N_21499,N_20163,N_20223);
xnor U21500 (N_21500,N_20662,N_20813);
nand U21501 (N_21501,N_20893,N_20936);
and U21502 (N_21502,N_20684,N_20313);
nand U21503 (N_21503,N_20035,N_20572);
and U21504 (N_21504,N_20383,N_20302);
or U21505 (N_21505,N_20090,N_20008);
and U21506 (N_21506,N_20216,N_20124);
and U21507 (N_21507,N_20583,N_20065);
or U21508 (N_21508,N_20594,N_20140);
nand U21509 (N_21509,N_20952,N_20071);
or U21510 (N_21510,N_20884,N_20971);
nand U21511 (N_21511,N_20380,N_20440);
nor U21512 (N_21512,N_20667,N_20013);
or U21513 (N_21513,N_20000,N_20179);
or U21514 (N_21514,N_20067,N_20424);
and U21515 (N_21515,N_20168,N_20899);
and U21516 (N_21516,N_20071,N_20691);
nand U21517 (N_21517,N_20705,N_20411);
nand U21518 (N_21518,N_20031,N_20179);
nor U21519 (N_21519,N_20543,N_20576);
nor U21520 (N_21520,N_20366,N_20150);
nor U21521 (N_21521,N_20217,N_20849);
nor U21522 (N_21522,N_20634,N_20740);
nand U21523 (N_21523,N_20104,N_20313);
nand U21524 (N_21524,N_20207,N_20579);
and U21525 (N_21525,N_20829,N_20216);
nand U21526 (N_21526,N_20790,N_20168);
and U21527 (N_21527,N_20302,N_20065);
xnor U21528 (N_21528,N_20697,N_20511);
xnor U21529 (N_21529,N_20509,N_20662);
nand U21530 (N_21530,N_20158,N_20360);
nand U21531 (N_21531,N_20804,N_20582);
xnor U21532 (N_21532,N_20295,N_20025);
and U21533 (N_21533,N_20003,N_20031);
nor U21534 (N_21534,N_20371,N_20536);
nor U21535 (N_21535,N_20399,N_20195);
or U21536 (N_21536,N_20526,N_20518);
or U21537 (N_21537,N_20677,N_20083);
or U21538 (N_21538,N_20379,N_20333);
nor U21539 (N_21539,N_20473,N_20339);
or U21540 (N_21540,N_20633,N_20548);
nor U21541 (N_21541,N_20837,N_20559);
nor U21542 (N_21542,N_20828,N_20569);
xnor U21543 (N_21543,N_20370,N_20973);
xor U21544 (N_21544,N_20777,N_20767);
nand U21545 (N_21545,N_20060,N_20104);
or U21546 (N_21546,N_20778,N_20098);
nand U21547 (N_21547,N_20861,N_20798);
xnor U21548 (N_21548,N_20551,N_20414);
nand U21549 (N_21549,N_20534,N_20551);
nor U21550 (N_21550,N_20158,N_20312);
and U21551 (N_21551,N_20092,N_20707);
nand U21552 (N_21552,N_20554,N_20699);
and U21553 (N_21553,N_20000,N_20444);
xnor U21554 (N_21554,N_20049,N_20827);
nor U21555 (N_21555,N_20353,N_20940);
xor U21556 (N_21556,N_20577,N_20169);
nor U21557 (N_21557,N_20600,N_20871);
nand U21558 (N_21558,N_20477,N_20600);
nand U21559 (N_21559,N_20837,N_20677);
xnor U21560 (N_21560,N_20912,N_20365);
or U21561 (N_21561,N_20133,N_20338);
xnor U21562 (N_21562,N_20890,N_20690);
nor U21563 (N_21563,N_20064,N_20079);
and U21564 (N_21564,N_20122,N_20283);
xnor U21565 (N_21565,N_20047,N_20568);
nor U21566 (N_21566,N_20636,N_20203);
or U21567 (N_21567,N_20171,N_20497);
nand U21568 (N_21568,N_20343,N_20232);
and U21569 (N_21569,N_20340,N_20102);
and U21570 (N_21570,N_20751,N_20412);
and U21571 (N_21571,N_20556,N_20541);
nor U21572 (N_21572,N_20084,N_20683);
nand U21573 (N_21573,N_20767,N_20947);
xnor U21574 (N_21574,N_20127,N_20594);
and U21575 (N_21575,N_20952,N_20878);
and U21576 (N_21576,N_20564,N_20221);
and U21577 (N_21577,N_20037,N_20252);
nand U21578 (N_21578,N_20764,N_20569);
and U21579 (N_21579,N_20586,N_20055);
and U21580 (N_21580,N_20156,N_20515);
and U21581 (N_21581,N_20816,N_20441);
and U21582 (N_21582,N_20768,N_20677);
or U21583 (N_21583,N_20936,N_20837);
or U21584 (N_21584,N_20318,N_20177);
xor U21585 (N_21585,N_20687,N_20260);
nand U21586 (N_21586,N_20599,N_20059);
and U21587 (N_21587,N_20493,N_20126);
nor U21588 (N_21588,N_20920,N_20074);
nor U21589 (N_21589,N_20155,N_20007);
nor U21590 (N_21590,N_20087,N_20021);
nand U21591 (N_21591,N_20973,N_20836);
nor U21592 (N_21592,N_20716,N_20538);
nand U21593 (N_21593,N_20545,N_20163);
nand U21594 (N_21594,N_20313,N_20100);
xor U21595 (N_21595,N_20480,N_20761);
and U21596 (N_21596,N_20197,N_20867);
and U21597 (N_21597,N_20323,N_20670);
or U21598 (N_21598,N_20579,N_20317);
and U21599 (N_21599,N_20841,N_20118);
xnor U21600 (N_21600,N_20826,N_20013);
nand U21601 (N_21601,N_20439,N_20929);
and U21602 (N_21602,N_20333,N_20273);
nor U21603 (N_21603,N_20549,N_20274);
or U21604 (N_21604,N_20088,N_20469);
or U21605 (N_21605,N_20831,N_20553);
nand U21606 (N_21606,N_20519,N_20337);
xnor U21607 (N_21607,N_20169,N_20259);
nand U21608 (N_21608,N_20637,N_20978);
or U21609 (N_21609,N_20634,N_20385);
and U21610 (N_21610,N_20835,N_20821);
nand U21611 (N_21611,N_20680,N_20359);
nor U21612 (N_21612,N_20080,N_20104);
or U21613 (N_21613,N_20002,N_20031);
nor U21614 (N_21614,N_20325,N_20843);
xor U21615 (N_21615,N_20411,N_20649);
nand U21616 (N_21616,N_20886,N_20855);
and U21617 (N_21617,N_20437,N_20578);
nor U21618 (N_21618,N_20214,N_20626);
and U21619 (N_21619,N_20894,N_20758);
xnor U21620 (N_21620,N_20171,N_20374);
nand U21621 (N_21621,N_20763,N_20039);
or U21622 (N_21622,N_20782,N_20554);
nand U21623 (N_21623,N_20391,N_20386);
and U21624 (N_21624,N_20773,N_20368);
xor U21625 (N_21625,N_20012,N_20265);
nand U21626 (N_21626,N_20047,N_20942);
xnor U21627 (N_21627,N_20790,N_20592);
and U21628 (N_21628,N_20614,N_20669);
nor U21629 (N_21629,N_20432,N_20820);
or U21630 (N_21630,N_20744,N_20912);
and U21631 (N_21631,N_20181,N_20228);
nor U21632 (N_21632,N_20675,N_20215);
or U21633 (N_21633,N_20265,N_20681);
nand U21634 (N_21634,N_20428,N_20064);
xnor U21635 (N_21635,N_20646,N_20895);
nand U21636 (N_21636,N_20436,N_20476);
and U21637 (N_21637,N_20033,N_20218);
xnor U21638 (N_21638,N_20803,N_20084);
or U21639 (N_21639,N_20351,N_20292);
nand U21640 (N_21640,N_20672,N_20054);
and U21641 (N_21641,N_20536,N_20387);
nand U21642 (N_21642,N_20455,N_20787);
nor U21643 (N_21643,N_20721,N_20404);
nor U21644 (N_21644,N_20290,N_20320);
nor U21645 (N_21645,N_20660,N_20529);
nor U21646 (N_21646,N_20322,N_20153);
and U21647 (N_21647,N_20560,N_20871);
xor U21648 (N_21648,N_20165,N_20529);
nand U21649 (N_21649,N_20094,N_20914);
nand U21650 (N_21650,N_20548,N_20394);
or U21651 (N_21651,N_20223,N_20641);
and U21652 (N_21652,N_20386,N_20912);
nor U21653 (N_21653,N_20226,N_20609);
nor U21654 (N_21654,N_20099,N_20113);
nand U21655 (N_21655,N_20288,N_20863);
and U21656 (N_21656,N_20198,N_20015);
nand U21657 (N_21657,N_20853,N_20305);
nand U21658 (N_21658,N_20082,N_20083);
xnor U21659 (N_21659,N_20632,N_20844);
nor U21660 (N_21660,N_20989,N_20426);
xnor U21661 (N_21661,N_20131,N_20097);
xnor U21662 (N_21662,N_20496,N_20208);
and U21663 (N_21663,N_20182,N_20778);
nor U21664 (N_21664,N_20473,N_20021);
nand U21665 (N_21665,N_20475,N_20169);
xor U21666 (N_21666,N_20648,N_20375);
xnor U21667 (N_21667,N_20981,N_20047);
nor U21668 (N_21668,N_20059,N_20164);
and U21669 (N_21669,N_20908,N_20197);
xor U21670 (N_21670,N_20720,N_20819);
or U21671 (N_21671,N_20318,N_20958);
nor U21672 (N_21672,N_20201,N_20823);
nor U21673 (N_21673,N_20860,N_20867);
nand U21674 (N_21674,N_20290,N_20250);
or U21675 (N_21675,N_20130,N_20572);
xor U21676 (N_21676,N_20085,N_20685);
nor U21677 (N_21677,N_20512,N_20343);
nand U21678 (N_21678,N_20988,N_20338);
and U21679 (N_21679,N_20453,N_20047);
nor U21680 (N_21680,N_20756,N_20401);
nor U21681 (N_21681,N_20830,N_20391);
xor U21682 (N_21682,N_20771,N_20227);
or U21683 (N_21683,N_20721,N_20827);
and U21684 (N_21684,N_20456,N_20692);
and U21685 (N_21685,N_20730,N_20979);
and U21686 (N_21686,N_20978,N_20379);
and U21687 (N_21687,N_20438,N_20175);
nor U21688 (N_21688,N_20773,N_20509);
and U21689 (N_21689,N_20559,N_20140);
nand U21690 (N_21690,N_20842,N_20441);
nor U21691 (N_21691,N_20103,N_20312);
nand U21692 (N_21692,N_20374,N_20959);
nor U21693 (N_21693,N_20005,N_20617);
or U21694 (N_21694,N_20472,N_20571);
and U21695 (N_21695,N_20096,N_20362);
or U21696 (N_21696,N_20726,N_20056);
nand U21697 (N_21697,N_20789,N_20343);
nor U21698 (N_21698,N_20276,N_20436);
and U21699 (N_21699,N_20668,N_20745);
or U21700 (N_21700,N_20748,N_20088);
or U21701 (N_21701,N_20582,N_20371);
nand U21702 (N_21702,N_20500,N_20016);
nor U21703 (N_21703,N_20228,N_20280);
nand U21704 (N_21704,N_20050,N_20195);
nand U21705 (N_21705,N_20964,N_20992);
nor U21706 (N_21706,N_20846,N_20437);
and U21707 (N_21707,N_20582,N_20004);
nand U21708 (N_21708,N_20702,N_20705);
nand U21709 (N_21709,N_20199,N_20410);
and U21710 (N_21710,N_20628,N_20444);
xor U21711 (N_21711,N_20276,N_20132);
or U21712 (N_21712,N_20662,N_20629);
and U21713 (N_21713,N_20940,N_20084);
nand U21714 (N_21714,N_20647,N_20418);
nand U21715 (N_21715,N_20155,N_20328);
xnor U21716 (N_21716,N_20662,N_20253);
xor U21717 (N_21717,N_20205,N_20287);
or U21718 (N_21718,N_20767,N_20419);
xor U21719 (N_21719,N_20936,N_20690);
nor U21720 (N_21720,N_20109,N_20743);
nor U21721 (N_21721,N_20162,N_20223);
xnor U21722 (N_21722,N_20878,N_20279);
xnor U21723 (N_21723,N_20102,N_20651);
nand U21724 (N_21724,N_20191,N_20280);
and U21725 (N_21725,N_20830,N_20596);
and U21726 (N_21726,N_20437,N_20171);
or U21727 (N_21727,N_20873,N_20662);
nor U21728 (N_21728,N_20217,N_20552);
nand U21729 (N_21729,N_20166,N_20819);
nor U21730 (N_21730,N_20310,N_20501);
xnor U21731 (N_21731,N_20498,N_20530);
and U21732 (N_21732,N_20032,N_20257);
or U21733 (N_21733,N_20183,N_20066);
and U21734 (N_21734,N_20412,N_20746);
and U21735 (N_21735,N_20151,N_20561);
and U21736 (N_21736,N_20577,N_20590);
xnor U21737 (N_21737,N_20334,N_20609);
and U21738 (N_21738,N_20579,N_20296);
nand U21739 (N_21739,N_20218,N_20043);
and U21740 (N_21740,N_20783,N_20092);
or U21741 (N_21741,N_20196,N_20055);
or U21742 (N_21742,N_20077,N_20155);
and U21743 (N_21743,N_20476,N_20209);
and U21744 (N_21744,N_20100,N_20533);
and U21745 (N_21745,N_20438,N_20525);
xor U21746 (N_21746,N_20938,N_20743);
xor U21747 (N_21747,N_20981,N_20329);
xnor U21748 (N_21748,N_20755,N_20791);
and U21749 (N_21749,N_20275,N_20911);
or U21750 (N_21750,N_20088,N_20092);
or U21751 (N_21751,N_20770,N_20157);
xor U21752 (N_21752,N_20392,N_20954);
nand U21753 (N_21753,N_20237,N_20329);
nand U21754 (N_21754,N_20395,N_20044);
xor U21755 (N_21755,N_20261,N_20360);
xnor U21756 (N_21756,N_20762,N_20081);
and U21757 (N_21757,N_20254,N_20462);
and U21758 (N_21758,N_20890,N_20415);
nor U21759 (N_21759,N_20929,N_20839);
nor U21760 (N_21760,N_20966,N_20623);
nor U21761 (N_21761,N_20553,N_20647);
xor U21762 (N_21762,N_20212,N_20480);
xnor U21763 (N_21763,N_20393,N_20269);
and U21764 (N_21764,N_20706,N_20686);
and U21765 (N_21765,N_20557,N_20149);
nand U21766 (N_21766,N_20165,N_20550);
xnor U21767 (N_21767,N_20815,N_20943);
nand U21768 (N_21768,N_20925,N_20984);
nand U21769 (N_21769,N_20140,N_20270);
xor U21770 (N_21770,N_20392,N_20253);
xnor U21771 (N_21771,N_20094,N_20653);
xor U21772 (N_21772,N_20389,N_20992);
nand U21773 (N_21773,N_20130,N_20941);
or U21774 (N_21774,N_20497,N_20946);
and U21775 (N_21775,N_20025,N_20336);
or U21776 (N_21776,N_20054,N_20057);
or U21777 (N_21777,N_20986,N_20332);
or U21778 (N_21778,N_20165,N_20392);
nor U21779 (N_21779,N_20657,N_20331);
nand U21780 (N_21780,N_20189,N_20208);
nor U21781 (N_21781,N_20160,N_20880);
xnor U21782 (N_21782,N_20976,N_20537);
xnor U21783 (N_21783,N_20679,N_20342);
and U21784 (N_21784,N_20268,N_20094);
nand U21785 (N_21785,N_20026,N_20295);
nor U21786 (N_21786,N_20290,N_20292);
and U21787 (N_21787,N_20642,N_20511);
or U21788 (N_21788,N_20676,N_20593);
xor U21789 (N_21789,N_20659,N_20008);
nand U21790 (N_21790,N_20927,N_20097);
or U21791 (N_21791,N_20891,N_20622);
or U21792 (N_21792,N_20074,N_20008);
xor U21793 (N_21793,N_20510,N_20839);
xnor U21794 (N_21794,N_20940,N_20149);
or U21795 (N_21795,N_20130,N_20287);
or U21796 (N_21796,N_20794,N_20406);
and U21797 (N_21797,N_20877,N_20870);
nor U21798 (N_21798,N_20272,N_20243);
nand U21799 (N_21799,N_20831,N_20707);
xnor U21800 (N_21800,N_20795,N_20257);
nor U21801 (N_21801,N_20065,N_20845);
xnor U21802 (N_21802,N_20084,N_20934);
or U21803 (N_21803,N_20864,N_20302);
nand U21804 (N_21804,N_20957,N_20004);
xor U21805 (N_21805,N_20399,N_20900);
nand U21806 (N_21806,N_20578,N_20313);
xnor U21807 (N_21807,N_20208,N_20153);
xor U21808 (N_21808,N_20475,N_20680);
and U21809 (N_21809,N_20470,N_20949);
and U21810 (N_21810,N_20909,N_20985);
and U21811 (N_21811,N_20122,N_20895);
or U21812 (N_21812,N_20115,N_20305);
nand U21813 (N_21813,N_20076,N_20603);
nor U21814 (N_21814,N_20195,N_20363);
xor U21815 (N_21815,N_20181,N_20464);
and U21816 (N_21816,N_20150,N_20899);
or U21817 (N_21817,N_20564,N_20399);
nand U21818 (N_21818,N_20684,N_20511);
xnor U21819 (N_21819,N_20285,N_20451);
xnor U21820 (N_21820,N_20611,N_20469);
nand U21821 (N_21821,N_20517,N_20052);
or U21822 (N_21822,N_20003,N_20196);
nand U21823 (N_21823,N_20725,N_20544);
nor U21824 (N_21824,N_20777,N_20940);
xor U21825 (N_21825,N_20847,N_20532);
and U21826 (N_21826,N_20290,N_20869);
and U21827 (N_21827,N_20733,N_20205);
or U21828 (N_21828,N_20900,N_20542);
nand U21829 (N_21829,N_20331,N_20632);
nand U21830 (N_21830,N_20451,N_20453);
and U21831 (N_21831,N_20961,N_20681);
xor U21832 (N_21832,N_20013,N_20829);
nor U21833 (N_21833,N_20270,N_20660);
and U21834 (N_21834,N_20771,N_20899);
nand U21835 (N_21835,N_20265,N_20873);
nand U21836 (N_21836,N_20280,N_20753);
nand U21837 (N_21837,N_20438,N_20292);
nor U21838 (N_21838,N_20349,N_20855);
nor U21839 (N_21839,N_20701,N_20980);
nand U21840 (N_21840,N_20033,N_20141);
and U21841 (N_21841,N_20822,N_20283);
nand U21842 (N_21842,N_20030,N_20145);
nor U21843 (N_21843,N_20403,N_20804);
xnor U21844 (N_21844,N_20612,N_20530);
or U21845 (N_21845,N_20250,N_20483);
or U21846 (N_21846,N_20499,N_20704);
nor U21847 (N_21847,N_20109,N_20114);
xnor U21848 (N_21848,N_20651,N_20766);
xor U21849 (N_21849,N_20940,N_20551);
or U21850 (N_21850,N_20463,N_20002);
nand U21851 (N_21851,N_20837,N_20276);
and U21852 (N_21852,N_20890,N_20172);
and U21853 (N_21853,N_20015,N_20938);
or U21854 (N_21854,N_20638,N_20255);
and U21855 (N_21855,N_20024,N_20160);
xor U21856 (N_21856,N_20409,N_20085);
or U21857 (N_21857,N_20166,N_20255);
and U21858 (N_21858,N_20040,N_20871);
and U21859 (N_21859,N_20604,N_20293);
nand U21860 (N_21860,N_20914,N_20701);
or U21861 (N_21861,N_20171,N_20645);
xor U21862 (N_21862,N_20400,N_20916);
xor U21863 (N_21863,N_20114,N_20268);
nor U21864 (N_21864,N_20961,N_20947);
and U21865 (N_21865,N_20194,N_20157);
and U21866 (N_21866,N_20787,N_20608);
and U21867 (N_21867,N_20333,N_20244);
nor U21868 (N_21868,N_20586,N_20214);
nor U21869 (N_21869,N_20979,N_20119);
and U21870 (N_21870,N_20053,N_20516);
or U21871 (N_21871,N_20930,N_20584);
or U21872 (N_21872,N_20833,N_20178);
and U21873 (N_21873,N_20448,N_20346);
nand U21874 (N_21874,N_20568,N_20725);
nor U21875 (N_21875,N_20889,N_20973);
and U21876 (N_21876,N_20790,N_20310);
or U21877 (N_21877,N_20833,N_20524);
nand U21878 (N_21878,N_20095,N_20174);
or U21879 (N_21879,N_20405,N_20894);
nand U21880 (N_21880,N_20307,N_20663);
or U21881 (N_21881,N_20068,N_20129);
xnor U21882 (N_21882,N_20994,N_20844);
and U21883 (N_21883,N_20740,N_20657);
and U21884 (N_21884,N_20490,N_20868);
xor U21885 (N_21885,N_20016,N_20873);
xnor U21886 (N_21886,N_20636,N_20389);
nand U21887 (N_21887,N_20532,N_20659);
nor U21888 (N_21888,N_20606,N_20961);
xor U21889 (N_21889,N_20303,N_20118);
xnor U21890 (N_21890,N_20484,N_20924);
nor U21891 (N_21891,N_20290,N_20104);
or U21892 (N_21892,N_20667,N_20961);
xor U21893 (N_21893,N_20792,N_20384);
or U21894 (N_21894,N_20494,N_20910);
nor U21895 (N_21895,N_20916,N_20107);
xor U21896 (N_21896,N_20034,N_20893);
xnor U21897 (N_21897,N_20445,N_20360);
nor U21898 (N_21898,N_20132,N_20353);
nor U21899 (N_21899,N_20564,N_20487);
nor U21900 (N_21900,N_20035,N_20190);
nor U21901 (N_21901,N_20558,N_20030);
or U21902 (N_21902,N_20196,N_20281);
nand U21903 (N_21903,N_20210,N_20419);
and U21904 (N_21904,N_20861,N_20158);
or U21905 (N_21905,N_20044,N_20099);
nor U21906 (N_21906,N_20054,N_20039);
or U21907 (N_21907,N_20858,N_20203);
xor U21908 (N_21908,N_20115,N_20974);
nor U21909 (N_21909,N_20346,N_20948);
nand U21910 (N_21910,N_20147,N_20888);
xor U21911 (N_21911,N_20298,N_20771);
nor U21912 (N_21912,N_20939,N_20208);
nand U21913 (N_21913,N_20111,N_20560);
or U21914 (N_21914,N_20926,N_20568);
or U21915 (N_21915,N_20053,N_20764);
or U21916 (N_21916,N_20105,N_20265);
or U21917 (N_21917,N_20814,N_20813);
and U21918 (N_21918,N_20694,N_20015);
and U21919 (N_21919,N_20023,N_20575);
and U21920 (N_21920,N_20567,N_20622);
or U21921 (N_21921,N_20298,N_20729);
nor U21922 (N_21922,N_20221,N_20513);
nor U21923 (N_21923,N_20478,N_20876);
xor U21924 (N_21924,N_20768,N_20085);
xnor U21925 (N_21925,N_20049,N_20915);
xor U21926 (N_21926,N_20536,N_20889);
nor U21927 (N_21927,N_20436,N_20446);
and U21928 (N_21928,N_20821,N_20427);
or U21929 (N_21929,N_20792,N_20784);
nor U21930 (N_21930,N_20340,N_20434);
or U21931 (N_21931,N_20010,N_20851);
nand U21932 (N_21932,N_20494,N_20035);
xnor U21933 (N_21933,N_20948,N_20110);
nand U21934 (N_21934,N_20607,N_20372);
nand U21935 (N_21935,N_20544,N_20248);
or U21936 (N_21936,N_20330,N_20557);
nor U21937 (N_21937,N_20795,N_20955);
or U21938 (N_21938,N_20760,N_20717);
and U21939 (N_21939,N_20548,N_20267);
and U21940 (N_21940,N_20605,N_20593);
nor U21941 (N_21941,N_20679,N_20888);
nand U21942 (N_21942,N_20465,N_20509);
xnor U21943 (N_21943,N_20916,N_20951);
and U21944 (N_21944,N_20139,N_20622);
or U21945 (N_21945,N_20378,N_20898);
nand U21946 (N_21946,N_20130,N_20428);
nor U21947 (N_21947,N_20596,N_20422);
nand U21948 (N_21948,N_20745,N_20726);
nand U21949 (N_21949,N_20420,N_20191);
or U21950 (N_21950,N_20982,N_20301);
or U21951 (N_21951,N_20374,N_20907);
xnor U21952 (N_21952,N_20702,N_20172);
nand U21953 (N_21953,N_20472,N_20941);
and U21954 (N_21954,N_20597,N_20242);
or U21955 (N_21955,N_20568,N_20394);
xor U21956 (N_21956,N_20165,N_20907);
xnor U21957 (N_21957,N_20627,N_20959);
and U21958 (N_21958,N_20807,N_20891);
nor U21959 (N_21959,N_20043,N_20193);
and U21960 (N_21960,N_20203,N_20435);
nor U21961 (N_21961,N_20777,N_20583);
and U21962 (N_21962,N_20502,N_20872);
nand U21963 (N_21963,N_20835,N_20722);
nor U21964 (N_21964,N_20481,N_20773);
or U21965 (N_21965,N_20517,N_20617);
nor U21966 (N_21966,N_20204,N_20837);
or U21967 (N_21967,N_20448,N_20285);
nor U21968 (N_21968,N_20336,N_20972);
nor U21969 (N_21969,N_20213,N_20427);
or U21970 (N_21970,N_20764,N_20800);
xnor U21971 (N_21971,N_20252,N_20184);
xnor U21972 (N_21972,N_20308,N_20630);
or U21973 (N_21973,N_20595,N_20437);
or U21974 (N_21974,N_20935,N_20520);
or U21975 (N_21975,N_20585,N_20414);
and U21976 (N_21976,N_20857,N_20445);
nor U21977 (N_21977,N_20005,N_20379);
xor U21978 (N_21978,N_20901,N_20656);
xor U21979 (N_21979,N_20216,N_20274);
and U21980 (N_21980,N_20682,N_20195);
nor U21981 (N_21981,N_20095,N_20546);
nor U21982 (N_21982,N_20622,N_20389);
or U21983 (N_21983,N_20169,N_20521);
nand U21984 (N_21984,N_20587,N_20974);
and U21985 (N_21985,N_20926,N_20251);
xnor U21986 (N_21986,N_20767,N_20349);
nand U21987 (N_21987,N_20600,N_20722);
or U21988 (N_21988,N_20112,N_20224);
xor U21989 (N_21989,N_20980,N_20981);
nor U21990 (N_21990,N_20421,N_20738);
and U21991 (N_21991,N_20255,N_20551);
xor U21992 (N_21992,N_20646,N_20893);
nand U21993 (N_21993,N_20982,N_20721);
xnor U21994 (N_21994,N_20937,N_20311);
nor U21995 (N_21995,N_20178,N_20933);
nor U21996 (N_21996,N_20456,N_20306);
and U21997 (N_21997,N_20729,N_20800);
nor U21998 (N_21998,N_20681,N_20272);
nand U21999 (N_21999,N_20145,N_20597);
or U22000 (N_22000,N_21354,N_21716);
or U22001 (N_22001,N_21203,N_21845);
or U22002 (N_22002,N_21705,N_21639);
nand U22003 (N_22003,N_21435,N_21282);
nand U22004 (N_22004,N_21137,N_21686);
nor U22005 (N_22005,N_21249,N_21221);
and U22006 (N_22006,N_21696,N_21576);
or U22007 (N_22007,N_21041,N_21365);
xor U22008 (N_22008,N_21059,N_21875);
and U22009 (N_22009,N_21232,N_21720);
xnor U22010 (N_22010,N_21955,N_21828);
or U22011 (N_22011,N_21426,N_21063);
and U22012 (N_22012,N_21322,N_21323);
nand U22013 (N_22013,N_21465,N_21445);
xor U22014 (N_22014,N_21771,N_21848);
nand U22015 (N_22015,N_21053,N_21056);
nor U22016 (N_22016,N_21958,N_21613);
nor U22017 (N_22017,N_21795,N_21064);
nor U22018 (N_22018,N_21935,N_21852);
and U22019 (N_22019,N_21976,N_21805);
xor U22020 (N_22020,N_21938,N_21051);
nand U22021 (N_22021,N_21261,N_21395);
xor U22022 (N_22022,N_21178,N_21279);
nand U22023 (N_22023,N_21708,N_21346);
nor U22024 (N_22024,N_21554,N_21572);
xor U22025 (N_22025,N_21623,N_21113);
nand U22026 (N_22026,N_21819,N_21460);
or U22027 (N_22027,N_21177,N_21704);
nor U22028 (N_22028,N_21683,N_21306);
and U22029 (N_22029,N_21389,N_21454);
or U22030 (N_22030,N_21746,N_21422);
and U22031 (N_22031,N_21072,N_21563);
xor U22032 (N_22032,N_21277,N_21187);
xor U22033 (N_22033,N_21268,N_21122);
nand U22034 (N_22034,N_21448,N_21790);
xor U22035 (N_22035,N_21786,N_21728);
and U22036 (N_22036,N_21183,N_21995);
nand U22037 (N_22037,N_21710,N_21689);
nand U22038 (N_22038,N_21257,N_21224);
and U22039 (N_22039,N_21396,N_21974);
nor U22040 (N_22040,N_21707,N_21991);
nand U22041 (N_22041,N_21698,N_21896);
xor U22042 (N_22042,N_21255,N_21632);
nor U22043 (N_22043,N_21289,N_21333);
and U22044 (N_22044,N_21114,N_21909);
or U22045 (N_22045,N_21436,N_21250);
nand U22046 (N_22046,N_21595,N_21592);
nor U22047 (N_22047,N_21823,N_21315);
or U22048 (N_22048,N_21060,N_21309);
xor U22049 (N_22049,N_21350,N_21058);
or U22050 (N_22050,N_21248,N_21959);
or U22051 (N_22051,N_21622,N_21159);
xnor U22052 (N_22052,N_21917,N_21530);
xnor U22053 (N_22053,N_21412,N_21128);
xor U22054 (N_22054,N_21711,N_21195);
or U22055 (N_22055,N_21544,N_21290);
or U22056 (N_22056,N_21300,N_21320);
and U22057 (N_22057,N_21830,N_21768);
xor U22058 (N_22058,N_21584,N_21497);
nand U22059 (N_22059,N_21449,N_21491);
xnor U22060 (N_22060,N_21509,N_21985);
and U22061 (N_22061,N_21406,N_21370);
xnor U22062 (N_22062,N_21831,N_21408);
nor U22063 (N_22063,N_21011,N_21314);
or U22064 (N_22064,N_21732,N_21508);
and U22065 (N_22065,N_21087,N_21597);
or U22066 (N_22066,N_21241,N_21007);
and U22067 (N_22067,N_21285,N_21086);
nand U22068 (N_22068,N_21299,N_21463);
or U22069 (N_22069,N_21336,N_21905);
xor U22070 (N_22070,N_21880,N_21681);
xor U22071 (N_22071,N_21235,N_21656);
or U22072 (N_22072,N_21380,N_21772);
and U22073 (N_22073,N_21504,N_21402);
or U22074 (N_22074,N_21853,N_21915);
and U22075 (N_22075,N_21457,N_21062);
xnor U22076 (N_22076,N_21994,N_21170);
or U22077 (N_22077,N_21349,N_21145);
or U22078 (N_22078,N_21283,N_21218);
nand U22079 (N_22079,N_21001,N_21256);
or U22080 (N_22080,N_21580,N_21479);
or U22081 (N_22081,N_21398,N_21245);
nand U22082 (N_22082,N_21782,N_21134);
nor U22083 (N_22083,N_21238,N_21547);
or U22084 (N_22084,N_21152,N_21918);
xor U22085 (N_22085,N_21319,N_21367);
and U22086 (N_22086,N_21943,N_21219);
or U22087 (N_22087,N_21269,N_21045);
or U22088 (N_22088,N_21032,N_21179);
xor U22089 (N_22089,N_21847,N_21736);
or U22090 (N_22090,N_21793,N_21230);
or U22091 (N_22091,N_21171,N_21416);
xnor U22092 (N_22092,N_21920,N_21749);
nand U22093 (N_22093,N_21528,N_21898);
nor U22094 (N_22094,N_21131,N_21461);
or U22095 (N_22095,N_21097,N_21127);
or U22096 (N_22096,N_21616,N_21886);
xor U22097 (N_22097,N_21796,N_21548);
nand U22098 (N_22098,N_21048,N_21857);
nand U22099 (N_22099,N_21685,N_21557);
xnor U22100 (N_22100,N_21537,N_21375);
nand U22101 (N_22101,N_21215,N_21302);
or U22102 (N_22102,N_21574,N_21964);
xnor U22103 (N_22103,N_21259,N_21526);
or U22104 (N_22104,N_21769,N_21017);
or U22105 (N_22105,N_21669,N_21270);
or U22106 (N_22106,N_21027,N_21956);
nand U22107 (N_22107,N_21675,N_21678);
or U22108 (N_22108,N_21579,N_21641);
or U22109 (N_22109,N_21676,N_21751);
or U22110 (N_22110,N_21680,N_21957);
xnor U22111 (N_22111,N_21442,N_21263);
or U22112 (N_22112,N_21721,N_21693);
nor U22113 (N_22113,N_21013,N_21397);
nor U22114 (N_22114,N_21541,N_21872);
nor U22115 (N_22115,N_21950,N_21111);
or U22116 (N_22116,N_21316,N_21654);
or U22117 (N_22117,N_21840,N_21779);
and U22118 (N_22118,N_21409,N_21419);
xor U22119 (N_22119,N_21907,N_21390);
or U22120 (N_22120,N_21106,N_21858);
nand U22121 (N_22121,N_21369,N_21602);
nand U22122 (N_22122,N_21026,N_21386);
and U22123 (N_22123,N_21405,N_21891);
or U22124 (N_22124,N_21201,N_21031);
or U22125 (N_22125,N_21975,N_21094);
and U22126 (N_22126,N_21077,N_21288);
xor U22127 (N_22127,N_21176,N_21908);
and U22128 (N_22128,N_21940,N_21627);
and U22129 (N_22129,N_21427,N_21564);
xor U22130 (N_22130,N_21560,N_21144);
nand U22131 (N_22131,N_21214,N_21157);
xnor U22132 (N_22132,N_21738,N_21212);
or U22133 (N_22133,N_21029,N_21861);
nand U22134 (N_22134,N_21362,N_21495);
or U22135 (N_22135,N_21521,N_21462);
and U22136 (N_22136,N_21892,N_21534);
and U22137 (N_22137,N_21832,N_21281);
or U22138 (N_22138,N_21879,N_21867);
xor U22139 (N_22139,N_21722,N_21266);
xor U22140 (N_22140,N_21699,N_21525);
nand U22141 (N_22141,N_21050,N_21643);
and U22142 (N_22142,N_21192,N_21142);
or U22143 (N_22143,N_21934,N_21765);
xnor U22144 (N_22144,N_21931,N_21120);
or U22145 (N_22145,N_21992,N_21717);
and U22146 (N_22146,N_21837,N_21735);
nor U22147 (N_22147,N_21480,N_21399);
and U22148 (N_22148,N_21359,N_21624);
nor U22149 (N_22149,N_21432,N_21229);
or U22150 (N_22150,N_21684,N_21864);
nor U22151 (N_22151,N_21260,N_21274);
nand U22152 (N_22152,N_21589,N_21997);
or U22153 (N_22153,N_21865,N_21207);
nand U22154 (N_22154,N_21527,N_21726);
or U22155 (N_22155,N_21523,N_21822);
or U22156 (N_22156,N_21014,N_21360);
nand U22157 (N_22157,N_21690,N_21640);
nand U22158 (N_22158,N_21567,N_21433);
xor U22159 (N_22159,N_21493,N_21724);
nand U22160 (N_22160,N_21753,N_21816);
and U22161 (N_22161,N_21827,N_21582);
xor U22162 (N_22162,N_21522,N_21265);
nand U22163 (N_22163,N_21904,N_21671);
nor U22164 (N_22164,N_21668,N_21503);
xor U22165 (N_22165,N_21102,N_21164);
xnor U22166 (N_22166,N_21307,N_21980);
xnor U22167 (N_22167,N_21090,N_21379);
nor U22168 (N_22168,N_21634,N_21264);
xnor U22169 (N_22169,N_21903,N_21093);
nor U22170 (N_22170,N_21666,N_21325);
and U22171 (N_22171,N_21791,N_21967);
xnor U22172 (N_22172,N_21468,N_21130);
and U22173 (N_22173,N_21701,N_21762);
or U22174 (N_22174,N_21351,N_21443);
or U22175 (N_22175,N_21107,N_21520);
and U22176 (N_22176,N_21621,N_21844);
xnor U22177 (N_22177,N_21785,N_21437);
and U22178 (N_22178,N_21910,N_21108);
xor U22179 (N_22179,N_21251,N_21930);
nand U22180 (N_22180,N_21650,N_21709);
nor U22181 (N_22181,N_21376,N_21764);
and U22182 (N_22182,N_21737,N_21970);
or U22183 (N_22183,N_21303,N_21665);
or U22184 (N_22184,N_21440,N_21658);
or U22185 (N_22185,N_21781,N_21514);
xor U22186 (N_22186,N_21916,N_21278);
or U22187 (N_22187,N_21963,N_21510);
xor U22188 (N_22188,N_21885,N_21894);
nand U22189 (N_22189,N_21899,N_21545);
xnor U22190 (N_22190,N_21425,N_21809);
or U22191 (N_22191,N_21944,N_21513);
and U22192 (N_22192,N_21789,N_21340);
and U22193 (N_22193,N_21850,N_21774);
or U22194 (N_22194,N_21186,N_21984);
and U22195 (N_22195,N_21338,N_21546);
nor U22196 (N_22196,N_21401,N_21608);
or U22197 (N_22197,N_21876,N_21648);
nor U22198 (N_22198,N_21755,N_21040);
or U22199 (N_22199,N_21743,N_21010);
or U22200 (N_22200,N_21391,N_21926);
nand U22201 (N_22201,N_21986,N_21517);
or U22202 (N_22202,N_21005,N_21893);
or U22203 (N_22203,N_21092,N_21889);
or U22204 (N_22204,N_21382,N_21039);
or U22205 (N_22205,N_21752,N_21361);
or U22206 (N_22206,N_21198,N_21500);
nor U22207 (N_22207,N_21364,N_21190);
nor U22208 (N_22208,N_21467,N_21777);
nand U22209 (N_22209,N_21953,N_21378);
xor U22210 (N_22210,N_21015,N_21182);
and U22211 (N_22211,N_21038,N_21759);
xor U22212 (N_22212,N_21125,N_21133);
xnor U22213 (N_22213,N_21512,N_21150);
xor U22214 (N_22214,N_21439,N_21078);
xor U22215 (N_22215,N_21043,N_21609);
nand U22216 (N_22216,N_21598,N_21363);
xor U22217 (N_22217,N_21109,N_21573);
nor U22218 (N_22218,N_21124,N_21585);
or U22219 (N_22219,N_21863,N_21611);
nor U22220 (N_22220,N_21838,N_21403);
or U22221 (N_22221,N_21551,N_21859);
nand U22222 (N_22222,N_21651,N_21477);
xor U22223 (N_22223,N_21836,N_21697);
nor U22224 (N_22224,N_21817,N_21223);
or U22225 (N_22225,N_21118,N_21210);
xor U22226 (N_22226,N_21856,N_21301);
or U22227 (N_22227,N_21653,N_21156);
nand U22228 (N_22228,N_21244,N_21679);
xor U22229 (N_22229,N_21694,N_21066);
nand U22230 (N_22230,N_21415,N_21162);
nor U22231 (N_22231,N_21494,N_21091);
xor U22232 (N_22232,N_21052,N_21146);
or U22233 (N_22233,N_21163,N_21536);
nand U22234 (N_22234,N_21583,N_21246);
or U22235 (N_22235,N_21550,N_21549);
or U22236 (N_22236,N_21115,N_21441);
nand U22237 (N_22237,N_21571,N_21947);
or U22238 (N_22238,N_21447,N_21706);
nand U22239 (N_22239,N_21960,N_21911);
xor U22240 (N_22240,N_21098,N_21371);
or U22241 (N_22241,N_21326,N_21253);
nand U22242 (N_22242,N_21730,N_21021);
or U22243 (N_22243,N_21141,N_21169);
xor U22244 (N_22244,N_21870,N_21797);
nand U22245 (N_22245,N_21343,N_21175);
nand U22246 (N_22246,N_21151,N_21339);
and U22247 (N_22247,N_21132,N_21160);
xor U22248 (N_22248,N_21312,N_21418);
nand U22249 (N_22249,N_21996,N_21407);
nor U22250 (N_22250,N_21474,N_21095);
and U22251 (N_22251,N_21217,N_21070);
and U22252 (N_22252,N_21939,N_21538);
and U22253 (N_22253,N_21516,N_21507);
or U22254 (N_22254,N_21023,N_21682);
or U22255 (N_22255,N_21153,N_21625);
nand U22256 (N_22256,N_21100,N_21922);
nand U22257 (N_22257,N_21455,N_21272);
xnor U22258 (N_22258,N_21154,N_21105);
and U22259 (N_22259,N_21096,N_21287);
or U22260 (N_22260,N_21515,N_21296);
and U22261 (N_22261,N_21842,N_21877);
xor U22262 (N_22262,N_21049,N_21660);
and U22263 (N_22263,N_21044,N_21475);
nor U22264 (N_22264,N_21388,N_21297);
nand U22265 (N_22265,N_21293,N_21887);
and U22266 (N_22266,N_21237,N_21900);
and U22267 (N_22267,N_21035,N_21925);
nand U22268 (N_22268,N_21065,N_21047);
and U22269 (N_22269,N_21496,N_21080);
or U22270 (N_22270,N_21635,N_21804);
nand U22271 (N_22271,N_21321,N_21148);
nand U22272 (N_22272,N_21057,N_21729);
or U22273 (N_22273,N_21135,N_21139);
nor U22274 (N_22274,N_21687,N_21610);
xnor U22275 (N_22275,N_21883,N_21155);
nand U22276 (N_22276,N_21890,N_21199);
or U22277 (N_22277,N_21982,N_21929);
or U22278 (N_22278,N_21394,N_21647);
nand U22279 (N_22279,N_21633,N_21628);
nor U22280 (N_22280,N_21869,N_21846);
and U22281 (N_22281,N_21194,N_21138);
nand U22282 (N_22282,N_21642,N_21763);
nand U22283 (N_22283,N_21173,N_21562);
nor U22284 (N_22284,N_21637,N_21191);
nand U22285 (N_22285,N_21747,N_21353);
and U22286 (N_22286,N_21941,N_21998);
xor U22287 (N_22287,N_21028,N_21381);
nor U22288 (N_22288,N_21030,N_21291);
and U22289 (N_22289,N_21404,N_21076);
and U22290 (N_22290,N_21631,N_21531);
nor U22291 (N_22291,N_21978,N_21488);
nand U22292 (N_22292,N_21143,N_21607);
xor U22293 (N_22293,N_21489,N_21638);
nand U22294 (N_22294,N_21271,N_21233);
nand U22295 (N_22295,N_21220,N_21239);
and U22296 (N_22296,N_21824,N_21101);
nand U22297 (N_22297,N_21902,N_21225);
xor U22298 (N_22298,N_21811,N_21775);
nor U22299 (N_22299,N_21841,N_21629);
nand U22300 (N_22300,N_21295,N_21843);
or U22301 (N_22301,N_21254,N_21670);
nor U22302 (N_22302,N_21766,N_21068);
nor U22303 (N_22303,N_21973,N_21599);
xnor U22304 (N_22304,N_21464,N_21617);
nand U22305 (N_22305,N_21601,N_21006);
nand U22306 (N_22306,N_21073,N_21161);
or U22307 (N_22307,N_21833,N_21189);
nand U22308 (N_22308,N_21486,N_21788);
nand U22309 (N_22309,N_21410,N_21444);
nand U22310 (N_22310,N_21104,N_21802);
xor U22311 (N_22311,N_21117,N_21636);
nand U22312 (N_22312,N_21818,N_21037);
nor U22313 (N_22313,N_21262,N_21919);
nand U22314 (N_22314,N_21387,N_21498);
or U22315 (N_22315,N_21061,N_21815);
and U22316 (N_22316,N_21429,N_21414);
xor U22317 (N_22317,N_21074,N_21335);
or U22318 (N_22318,N_21862,N_21147);
nand U22319 (N_22319,N_21228,N_21662);
xnor U22320 (N_22320,N_21897,N_21556);
nor U22321 (N_22321,N_21542,N_21025);
or U22322 (N_22322,N_21969,N_21334);
and U22323 (N_22323,N_21099,N_21569);
xor U22324 (N_22324,N_21649,N_21482);
and U22325 (N_22325,N_21661,N_21174);
nand U22326 (N_22326,N_21116,N_21317);
and U22327 (N_22327,N_21874,N_21966);
or U22328 (N_22328,N_21332,N_21924);
xor U22329 (N_22329,N_21088,N_21566);
nor U22330 (N_22330,N_21987,N_21206);
and U22331 (N_22331,N_21756,N_21373);
or U22332 (N_22332,N_21715,N_21196);
xor U22333 (N_22333,N_21760,N_21712);
xor U22334 (N_22334,N_21761,N_21347);
or U22335 (N_22335,N_21112,N_21591);
nor U22336 (N_22336,N_21055,N_21280);
and U22337 (N_22337,N_21646,N_21434);
nand U22338 (N_22338,N_21672,N_21803);
nor U22339 (N_22339,N_21552,N_21331);
nand U22340 (N_22340,N_21718,N_21558);
nor U22341 (N_22341,N_21559,N_21745);
nor U22342 (N_22342,N_21868,N_21368);
nor U22343 (N_22343,N_21612,N_21377);
xor U22344 (N_22344,N_21276,N_21129);
nor U22345 (N_22345,N_21519,N_21423);
or U22346 (N_22346,N_21532,N_21851);
xnor U22347 (N_22347,N_21501,N_21773);
and U22348 (N_22348,N_21505,N_21481);
nor U22349 (N_22349,N_21860,N_21535);
nand U22350 (N_22350,N_21392,N_21231);
or U22351 (N_22351,N_21324,N_21358);
and U22352 (N_22352,N_21744,N_21921);
or U22353 (N_22353,N_21723,N_21492);
xnor U22354 (N_22354,N_21511,N_21677);
and U22355 (N_22355,N_21881,N_21476);
nor U22356 (N_22356,N_21329,N_21968);
and U22357 (N_22357,N_21075,N_21172);
nor U22358 (N_22358,N_21878,N_21471);
and U22359 (N_22359,N_21620,N_21748);
nand U22360 (N_22360,N_21085,N_21298);
and U22361 (N_22361,N_21692,N_21424);
nor U22362 (N_22362,N_21575,N_21993);
nor U22363 (N_22363,N_21949,N_21603);
nor U22364 (N_22364,N_21374,N_21518);
nor U22365 (N_22365,N_21020,N_21733);
nor U22366 (N_22366,N_21691,N_21932);
xnor U22367 (N_22367,N_21002,N_21181);
nor U22368 (N_22368,N_21807,N_21197);
nand U22369 (N_22369,N_21742,N_21553);
nand U22370 (N_22370,N_21588,N_21470);
xnor U22371 (N_22371,N_21180,N_21543);
and U22372 (N_22372,N_21384,N_21741);
nor U22373 (N_22373,N_21529,N_21798);
and U22374 (N_22374,N_21204,N_21466);
or U22375 (N_22375,N_21411,N_21357);
or U22376 (N_22376,N_21213,N_21999);
nor U22377 (N_22377,N_21778,N_21019);
xnor U22378 (N_22378,N_21149,N_21784);
and U22379 (N_22379,N_21003,N_21615);
xor U22380 (N_22380,N_21311,N_21600);
or U22381 (N_22381,N_21590,N_21450);
nand U22382 (N_22382,N_21344,N_21024);
nand U22383 (N_22383,N_21792,N_21242);
xnor U22384 (N_22384,N_21740,N_21702);
nor U22385 (N_22385,N_21438,N_21839);
nand U22386 (N_22386,N_21989,N_21016);
xnor U22387 (N_22387,N_21451,N_21855);
xor U22388 (N_22388,N_21168,N_21914);
and U22389 (N_22389,N_21808,N_21485);
and U22390 (N_22390,N_21866,N_21829);
xnor U22391 (N_22391,N_21913,N_21258);
nor U22392 (N_22392,N_21252,N_21417);
nand U22393 (N_22393,N_21659,N_21000);
and U22394 (N_22394,N_21946,N_21446);
nand U22395 (N_22395,N_21933,N_21036);
and U22396 (N_22396,N_21727,N_21216);
nor U22397 (N_22397,N_21645,N_21568);
nand U22398 (N_22398,N_21854,N_21188);
xor U22399 (N_22399,N_21393,N_21069);
nand U22400 (N_22400,N_21121,N_21452);
nand U22401 (N_22401,N_21754,N_21923);
nand U22402 (N_22402,N_21304,N_21565);
xor U22403 (N_22403,N_21988,N_21103);
and U22404 (N_22404,N_21385,N_21945);
or U22405 (N_22405,N_21972,N_21459);
and U22406 (N_22406,N_21472,N_21337);
nor U22407 (N_22407,N_21082,N_21356);
nor U22408 (N_22408,N_21570,N_21873);
nand U22409 (N_22409,N_21713,N_21012);
nand U22410 (N_22410,N_21688,N_21596);
or U22411 (N_22411,N_21604,N_21383);
xor U22412 (N_22412,N_21205,N_21555);
xor U22413 (N_22413,N_21421,N_21342);
nand U22414 (N_22414,N_21912,N_21952);
xnor U22415 (N_22415,N_21499,N_21355);
xnor U22416 (N_22416,N_21979,N_21054);
or U22417 (N_22417,N_21165,N_21825);
xor U22418 (N_22418,N_21725,N_21273);
nor U22419 (N_22419,N_21067,N_21961);
nand U22420 (N_22420,N_21895,N_21185);
xor U22421 (N_22421,N_21084,N_21524);
or U22422 (N_22422,N_21420,N_21757);
nand U22423 (N_22423,N_21731,N_21313);
nand U22424 (N_22424,N_21714,N_21954);
nor U22425 (N_22425,N_21126,N_21734);
nor U22426 (N_22426,N_21906,N_21664);
and U22427 (N_22427,N_21540,N_21936);
or U22428 (N_22428,N_21750,N_21348);
and U22429 (N_22429,N_21123,N_21208);
or U22430 (N_22430,N_21275,N_21593);
and U22431 (N_22431,N_21430,N_21308);
nor U22432 (N_22432,N_21267,N_21366);
and U22433 (N_22433,N_21539,N_21081);
or U22434 (N_22434,N_21783,N_21614);
nand U22435 (N_22435,N_21089,N_21810);
or U22436 (N_22436,N_21110,N_21674);
nor U22437 (N_22437,N_21801,N_21473);
nor U22438 (N_22438,N_21990,N_21136);
and U22439 (N_22439,N_21884,N_21700);
nand U22440 (N_22440,N_21243,N_21226);
xor U22441 (N_22441,N_21587,N_21882);
nand U22442 (N_22442,N_21456,N_21849);
xnor U22443 (N_22443,N_21502,N_21167);
nor U22444 (N_22444,N_21719,N_21234);
nand U22445 (N_22445,N_21937,N_21506);
xor U22446 (N_22446,N_21806,N_21200);
nand U22447 (N_22447,N_21780,N_21901);
or U22448 (N_22448,N_21928,N_21305);
or U22449 (N_22449,N_21594,N_21372);
nor U22450 (N_22450,N_21657,N_21453);
and U22451 (N_22451,N_21079,N_21166);
xnor U22452 (N_22452,N_21618,N_21981);
and U22453 (N_22453,N_21431,N_21799);
and U22454 (N_22454,N_21428,N_21951);
xor U22455 (N_22455,N_21222,N_21812);
xnor U22456 (N_22456,N_21655,N_21813);
xor U22457 (N_22457,N_21652,N_21484);
xnor U22458 (N_22458,N_21942,N_21758);
nor U22459 (N_22459,N_21834,N_21965);
and U22460 (N_22460,N_21619,N_21794);
nor U22461 (N_22461,N_21983,N_21770);
or U22462 (N_22462,N_21240,N_21581);
nand U22463 (N_22463,N_21577,N_21478);
xor U22464 (N_22464,N_21022,N_21871);
nand U22465 (N_22465,N_21345,N_21948);
xnor U22466 (N_22466,N_21328,N_21458);
nor U22467 (N_22467,N_21490,N_21630);
or U22468 (N_22468,N_21211,N_21413);
nand U22469 (N_22469,N_21318,N_21483);
nand U22470 (N_22470,N_21046,N_21352);
nor U22471 (N_22471,N_21814,N_21835);
or U22472 (N_22472,N_21193,N_21247);
nor U22473 (N_22473,N_21008,N_21606);
nor U22474 (N_22474,N_21071,N_21158);
and U22475 (N_22475,N_21971,N_21561);
or U22476 (N_22476,N_21977,N_21695);
xor U22477 (N_22477,N_21578,N_21626);
xnor U22478 (N_22478,N_21202,N_21605);
nor U22479 (N_22479,N_21294,N_21888);
and U22480 (N_22480,N_21800,N_21292);
nor U22481 (N_22481,N_21739,N_21469);
xor U22482 (N_22482,N_21140,N_21310);
xnor U22483 (N_22483,N_21826,N_21487);
nor U22484 (N_22484,N_21184,N_21962);
or U22485 (N_22485,N_21663,N_21776);
xnor U22486 (N_22486,N_21644,N_21400);
and U22487 (N_22487,N_21236,N_21004);
nor U22488 (N_22488,N_21341,N_21083);
nor U22489 (N_22489,N_21821,N_21533);
nor U22490 (N_22490,N_21018,N_21586);
or U22491 (N_22491,N_21033,N_21284);
nand U22492 (N_22492,N_21327,N_21703);
nor U22493 (N_22493,N_21673,N_21820);
and U22494 (N_22494,N_21927,N_21767);
or U22495 (N_22495,N_21667,N_21787);
nand U22496 (N_22496,N_21119,N_21227);
nand U22497 (N_22497,N_21330,N_21034);
nor U22498 (N_22498,N_21042,N_21209);
nand U22499 (N_22499,N_21286,N_21009);
nor U22500 (N_22500,N_21101,N_21713);
or U22501 (N_22501,N_21543,N_21708);
nor U22502 (N_22502,N_21367,N_21201);
nor U22503 (N_22503,N_21806,N_21203);
nand U22504 (N_22504,N_21444,N_21771);
nor U22505 (N_22505,N_21760,N_21312);
and U22506 (N_22506,N_21986,N_21155);
or U22507 (N_22507,N_21835,N_21385);
xnor U22508 (N_22508,N_21015,N_21188);
and U22509 (N_22509,N_21453,N_21509);
or U22510 (N_22510,N_21314,N_21068);
nor U22511 (N_22511,N_21073,N_21038);
and U22512 (N_22512,N_21271,N_21189);
or U22513 (N_22513,N_21000,N_21151);
xor U22514 (N_22514,N_21593,N_21980);
or U22515 (N_22515,N_21692,N_21192);
and U22516 (N_22516,N_21983,N_21124);
or U22517 (N_22517,N_21743,N_21070);
xnor U22518 (N_22518,N_21004,N_21186);
nor U22519 (N_22519,N_21633,N_21982);
and U22520 (N_22520,N_21406,N_21455);
xnor U22521 (N_22521,N_21039,N_21486);
or U22522 (N_22522,N_21557,N_21376);
and U22523 (N_22523,N_21149,N_21232);
and U22524 (N_22524,N_21229,N_21577);
nand U22525 (N_22525,N_21441,N_21209);
xor U22526 (N_22526,N_21830,N_21165);
xnor U22527 (N_22527,N_21243,N_21500);
xnor U22528 (N_22528,N_21225,N_21726);
xnor U22529 (N_22529,N_21247,N_21072);
xor U22530 (N_22530,N_21136,N_21174);
nand U22531 (N_22531,N_21268,N_21466);
nand U22532 (N_22532,N_21978,N_21990);
and U22533 (N_22533,N_21956,N_21207);
nor U22534 (N_22534,N_21412,N_21859);
and U22535 (N_22535,N_21381,N_21886);
or U22536 (N_22536,N_21643,N_21571);
nor U22537 (N_22537,N_21032,N_21328);
nor U22538 (N_22538,N_21965,N_21317);
nor U22539 (N_22539,N_21716,N_21037);
and U22540 (N_22540,N_21137,N_21539);
nor U22541 (N_22541,N_21074,N_21259);
nand U22542 (N_22542,N_21086,N_21432);
or U22543 (N_22543,N_21763,N_21369);
or U22544 (N_22544,N_21410,N_21066);
or U22545 (N_22545,N_21208,N_21122);
and U22546 (N_22546,N_21506,N_21081);
nor U22547 (N_22547,N_21015,N_21480);
nor U22548 (N_22548,N_21286,N_21882);
xnor U22549 (N_22549,N_21128,N_21825);
or U22550 (N_22550,N_21496,N_21797);
nand U22551 (N_22551,N_21794,N_21189);
nor U22552 (N_22552,N_21999,N_21030);
and U22553 (N_22553,N_21914,N_21634);
nand U22554 (N_22554,N_21677,N_21649);
nor U22555 (N_22555,N_21641,N_21068);
or U22556 (N_22556,N_21672,N_21058);
or U22557 (N_22557,N_21178,N_21906);
nand U22558 (N_22558,N_21348,N_21101);
or U22559 (N_22559,N_21917,N_21100);
nand U22560 (N_22560,N_21891,N_21227);
xor U22561 (N_22561,N_21832,N_21793);
xnor U22562 (N_22562,N_21570,N_21512);
and U22563 (N_22563,N_21230,N_21279);
xor U22564 (N_22564,N_21691,N_21272);
and U22565 (N_22565,N_21079,N_21386);
nand U22566 (N_22566,N_21227,N_21453);
nor U22567 (N_22567,N_21044,N_21634);
nand U22568 (N_22568,N_21446,N_21860);
xnor U22569 (N_22569,N_21060,N_21163);
nand U22570 (N_22570,N_21229,N_21188);
nor U22571 (N_22571,N_21636,N_21323);
or U22572 (N_22572,N_21714,N_21753);
nor U22573 (N_22573,N_21685,N_21378);
nor U22574 (N_22574,N_21198,N_21362);
nand U22575 (N_22575,N_21654,N_21411);
xor U22576 (N_22576,N_21722,N_21242);
nand U22577 (N_22577,N_21227,N_21671);
nand U22578 (N_22578,N_21316,N_21142);
xnor U22579 (N_22579,N_21365,N_21093);
or U22580 (N_22580,N_21209,N_21974);
or U22581 (N_22581,N_21746,N_21489);
xor U22582 (N_22582,N_21081,N_21608);
nand U22583 (N_22583,N_21163,N_21607);
and U22584 (N_22584,N_21628,N_21989);
and U22585 (N_22585,N_21523,N_21672);
xnor U22586 (N_22586,N_21619,N_21482);
nor U22587 (N_22587,N_21543,N_21627);
or U22588 (N_22588,N_21199,N_21871);
xnor U22589 (N_22589,N_21443,N_21183);
nor U22590 (N_22590,N_21924,N_21171);
nand U22591 (N_22591,N_21925,N_21716);
xor U22592 (N_22592,N_21533,N_21835);
nand U22593 (N_22593,N_21886,N_21017);
or U22594 (N_22594,N_21126,N_21678);
nor U22595 (N_22595,N_21516,N_21769);
and U22596 (N_22596,N_21284,N_21296);
xnor U22597 (N_22597,N_21515,N_21069);
xnor U22598 (N_22598,N_21643,N_21949);
xnor U22599 (N_22599,N_21142,N_21319);
nand U22600 (N_22600,N_21946,N_21988);
xnor U22601 (N_22601,N_21690,N_21735);
xnor U22602 (N_22602,N_21955,N_21198);
and U22603 (N_22603,N_21855,N_21046);
nand U22604 (N_22604,N_21032,N_21475);
or U22605 (N_22605,N_21831,N_21929);
or U22606 (N_22606,N_21259,N_21549);
nand U22607 (N_22607,N_21551,N_21603);
nor U22608 (N_22608,N_21618,N_21929);
nand U22609 (N_22609,N_21512,N_21748);
xnor U22610 (N_22610,N_21217,N_21304);
nand U22611 (N_22611,N_21214,N_21013);
nand U22612 (N_22612,N_21728,N_21213);
nand U22613 (N_22613,N_21314,N_21530);
nand U22614 (N_22614,N_21523,N_21882);
and U22615 (N_22615,N_21707,N_21814);
nor U22616 (N_22616,N_21941,N_21353);
xnor U22617 (N_22617,N_21963,N_21188);
xor U22618 (N_22618,N_21385,N_21211);
nor U22619 (N_22619,N_21833,N_21759);
nand U22620 (N_22620,N_21574,N_21873);
nor U22621 (N_22621,N_21640,N_21369);
nor U22622 (N_22622,N_21637,N_21087);
xnor U22623 (N_22623,N_21682,N_21622);
nor U22624 (N_22624,N_21842,N_21123);
nor U22625 (N_22625,N_21070,N_21839);
xor U22626 (N_22626,N_21579,N_21970);
and U22627 (N_22627,N_21738,N_21168);
xnor U22628 (N_22628,N_21319,N_21524);
xor U22629 (N_22629,N_21771,N_21431);
nor U22630 (N_22630,N_21933,N_21443);
xor U22631 (N_22631,N_21155,N_21871);
nand U22632 (N_22632,N_21374,N_21338);
nand U22633 (N_22633,N_21795,N_21025);
xnor U22634 (N_22634,N_21533,N_21730);
xnor U22635 (N_22635,N_21577,N_21179);
nand U22636 (N_22636,N_21150,N_21433);
nor U22637 (N_22637,N_21920,N_21383);
or U22638 (N_22638,N_21742,N_21976);
or U22639 (N_22639,N_21422,N_21998);
and U22640 (N_22640,N_21438,N_21869);
xor U22641 (N_22641,N_21577,N_21630);
nand U22642 (N_22642,N_21617,N_21408);
and U22643 (N_22643,N_21806,N_21079);
and U22644 (N_22644,N_21870,N_21919);
nand U22645 (N_22645,N_21367,N_21748);
or U22646 (N_22646,N_21598,N_21682);
nor U22647 (N_22647,N_21804,N_21875);
nand U22648 (N_22648,N_21968,N_21525);
nand U22649 (N_22649,N_21698,N_21094);
and U22650 (N_22650,N_21279,N_21305);
nor U22651 (N_22651,N_21154,N_21085);
xor U22652 (N_22652,N_21136,N_21518);
or U22653 (N_22653,N_21310,N_21881);
xnor U22654 (N_22654,N_21682,N_21689);
and U22655 (N_22655,N_21686,N_21905);
nand U22656 (N_22656,N_21856,N_21326);
or U22657 (N_22657,N_21057,N_21841);
xnor U22658 (N_22658,N_21512,N_21946);
or U22659 (N_22659,N_21060,N_21429);
and U22660 (N_22660,N_21720,N_21320);
nand U22661 (N_22661,N_21936,N_21293);
and U22662 (N_22662,N_21939,N_21366);
nor U22663 (N_22663,N_21223,N_21094);
or U22664 (N_22664,N_21610,N_21928);
xnor U22665 (N_22665,N_21311,N_21340);
and U22666 (N_22666,N_21438,N_21197);
nor U22667 (N_22667,N_21823,N_21127);
and U22668 (N_22668,N_21825,N_21367);
nor U22669 (N_22669,N_21194,N_21304);
xor U22670 (N_22670,N_21651,N_21363);
and U22671 (N_22671,N_21569,N_21934);
or U22672 (N_22672,N_21626,N_21553);
xnor U22673 (N_22673,N_21155,N_21705);
nor U22674 (N_22674,N_21112,N_21204);
xnor U22675 (N_22675,N_21068,N_21047);
or U22676 (N_22676,N_21969,N_21751);
nor U22677 (N_22677,N_21600,N_21911);
nor U22678 (N_22678,N_21764,N_21683);
nor U22679 (N_22679,N_21278,N_21291);
and U22680 (N_22680,N_21932,N_21826);
and U22681 (N_22681,N_21818,N_21279);
xor U22682 (N_22682,N_21575,N_21635);
nand U22683 (N_22683,N_21686,N_21363);
or U22684 (N_22684,N_21284,N_21340);
or U22685 (N_22685,N_21888,N_21234);
nor U22686 (N_22686,N_21900,N_21189);
nor U22687 (N_22687,N_21180,N_21630);
nor U22688 (N_22688,N_21700,N_21265);
or U22689 (N_22689,N_21346,N_21076);
nand U22690 (N_22690,N_21335,N_21969);
and U22691 (N_22691,N_21378,N_21159);
nand U22692 (N_22692,N_21361,N_21907);
or U22693 (N_22693,N_21975,N_21253);
or U22694 (N_22694,N_21674,N_21760);
and U22695 (N_22695,N_21158,N_21559);
and U22696 (N_22696,N_21847,N_21226);
and U22697 (N_22697,N_21613,N_21278);
xor U22698 (N_22698,N_21795,N_21415);
nand U22699 (N_22699,N_21839,N_21627);
or U22700 (N_22700,N_21073,N_21678);
nand U22701 (N_22701,N_21729,N_21754);
xnor U22702 (N_22702,N_21162,N_21123);
nor U22703 (N_22703,N_21599,N_21988);
xnor U22704 (N_22704,N_21381,N_21885);
nor U22705 (N_22705,N_21740,N_21183);
nand U22706 (N_22706,N_21518,N_21860);
nor U22707 (N_22707,N_21403,N_21607);
or U22708 (N_22708,N_21059,N_21990);
nand U22709 (N_22709,N_21729,N_21104);
or U22710 (N_22710,N_21638,N_21309);
and U22711 (N_22711,N_21891,N_21783);
nand U22712 (N_22712,N_21637,N_21208);
nand U22713 (N_22713,N_21706,N_21099);
xnor U22714 (N_22714,N_21437,N_21663);
nand U22715 (N_22715,N_21720,N_21297);
or U22716 (N_22716,N_21403,N_21957);
xnor U22717 (N_22717,N_21178,N_21717);
nor U22718 (N_22718,N_21758,N_21505);
xor U22719 (N_22719,N_21655,N_21551);
xor U22720 (N_22720,N_21102,N_21697);
and U22721 (N_22721,N_21736,N_21770);
nand U22722 (N_22722,N_21383,N_21334);
or U22723 (N_22723,N_21396,N_21140);
nor U22724 (N_22724,N_21469,N_21701);
and U22725 (N_22725,N_21309,N_21377);
xor U22726 (N_22726,N_21368,N_21346);
xnor U22727 (N_22727,N_21578,N_21364);
nand U22728 (N_22728,N_21890,N_21605);
xnor U22729 (N_22729,N_21636,N_21255);
nand U22730 (N_22730,N_21827,N_21210);
nor U22731 (N_22731,N_21808,N_21703);
or U22732 (N_22732,N_21621,N_21334);
nor U22733 (N_22733,N_21286,N_21529);
xnor U22734 (N_22734,N_21423,N_21609);
nand U22735 (N_22735,N_21134,N_21862);
nor U22736 (N_22736,N_21662,N_21546);
xor U22737 (N_22737,N_21451,N_21129);
nand U22738 (N_22738,N_21807,N_21791);
xor U22739 (N_22739,N_21078,N_21742);
nor U22740 (N_22740,N_21256,N_21386);
xor U22741 (N_22741,N_21691,N_21372);
nand U22742 (N_22742,N_21731,N_21213);
nor U22743 (N_22743,N_21917,N_21741);
or U22744 (N_22744,N_21697,N_21216);
xnor U22745 (N_22745,N_21576,N_21900);
and U22746 (N_22746,N_21995,N_21096);
nor U22747 (N_22747,N_21573,N_21634);
xor U22748 (N_22748,N_21874,N_21608);
xor U22749 (N_22749,N_21022,N_21147);
and U22750 (N_22750,N_21001,N_21642);
nor U22751 (N_22751,N_21782,N_21875);
xnor U22752 (N_22752,N_21616,N_21767);
and U22753 (N_22753,N_21850,N_21438);
xnor U22754 (N_22754,N_21211,N_21597);
nor U22755 (N_22755,N_21929,N_21567);
nor U22756 (N_22756,N_21656,N_21748);
xnor U22757 (N_22757,N_21211,N_21843);
and U22758 (N_22758,N_21658,N_21278);
and U22759 (N_22759,N_21568,N_21922);
and U22760 (N_22760,N_21188,N_21710);
nor U22761 (N_22761,N_21211,N_21826);
nand U22762 (N_22762,N_21048,N_21101);
and U22763 (N_22763,N_21739,N_21369);
nand U22764 (N_22764,N_21352,N_21377);
xnor U22765 (N_22765,N_21144,N_21174);
xnor U22766 (N_22766,N_21829,N_21297);
nand U22767 (N_22767,N_21378,N_21773);
and U22768 (N_22768,N_21735,N_21742);
nor U22769 (N_22769,N_21680,N_21230);
nor U22770 (N_22770,N_21694,N_21809);
nand U22771 (N_22771,N_21510,N_21294);
and U22772 (N_22772,N_21906,N_21888);
xnor U22773 (N_22773,N_21983,N_21612);
and U22774 (N_22774,N_21478,N_21323);
nand U22775 (N_22775,N_21416,N_21787);
or U22776 (N_22776,N_21888,N_21985);
nand U22777 (N_22777,N_21998,N_21893);
or U22778 (N_22778,N_21323,N_21277);
nor U22779 (N_22779,N_21809,N_21263);
or U22780 (N_22780,N_21843,N_21937);
xnor U22781 (N_22781,N_21040,N_21638);
nor U22782 (N_22782,N_21958,N_21013);
xnor U22783 (N_22783,N_21189,N_21116);
or U22784 (N_22784,N_21473,N_21298);
and U22785 (N_22785,N_21990,N_21492);
nand U22786 (N_22786,N_21000,N_21195);
nand U22787 (N_22787,N_21155,N_21649);
nor U22788 (N_22788,N_21161,N_21165);
nor U22789 (N_22789,N_21649,N_21461);
nand U22790 (N_22790,N_21808,N_21085);
nor U22791 (N_22791,N_21479,N_21892);
or U22792 (N_22792,N_21553,N_21397);
nand U22793 (N_22793,N_21297,N_21431);
nand U22794 (N_22794,N_21773,N_21914);
nor U22795 (N_22795,N_21702,N_21026);
xnor U22796 (N_22796,N_21410,N_21838);
xnor U22797 (N_22797,N_21764,N_21470);
xor U22798 (N_22798,N_21827,N_21738);
or U22799 (N_22799,N_21375,N_21695);
xor U22800 (N_22800,N_21635,N_21253);
and U22801 (N_22801,N_21152,N_21123);
xnor U22802 (N_22802,N_21838,N_21927);
nor U22803 (N_22803,N_21944,N_21277);
or U22804 (N_22804,N_21685,N_21570);
and U22805 (N_22805,N_21971,N_21468);
and U22806 (N_22806,N_21179,N_21852);
and U22807 (N_22807,N_21277,N_21761);
nor U22808 (N_22808,N_21494,N_21737);
or U22809 (N_22809,N_21634,N_21941);
or U22810 (N_22810,N_21136,N_21319);
xor U22811 (N_22811,N_21888,N_21231);
and U22812 (N_22812,N_21427,N_21826);
and U22813 (N_22813,N_21203,N_21196);
nor U22814 (N_22814,N_21290,N_21610);
nor U22815 (N_22815,N_21004,N_21393);
and U22816 (N_22816,N_21373,N_21963);
or U22817 (N_22817,N_21866,N_21494);
nand U22818 (N_22818,N_21168,N_21712);
or U22819 (N_22819,N_21504,N_21540);
nor U22820 (N_22820,N_21000,N_21039);
nor U22821 (N_22821,N_21662,N_21443);
nor U22822 (N_22822,N_21172,N_21310);
xor U22823 (N_22823,N_21442,N_21235);
or U22824 (N_22824,N_21837,N_21454);
or U22825 (N_22825,N_21914,N_21883);
xnor U22826 (N_22826,N_21506,N_21935);
xnor U22827 (N_22827,N_21740,N_21298);
and U22828 (N_22828,N_21236,N_21143);
and U22829 (N_22829,N_21894,N_21730);
and U22830 (N_22830,N_21873,N_21875);
or U22831 (N_22831,N_21098,N_21528);
and U22832 (N_22832,N_21767,N_21806);
or U22833 (N_22833,N_21092,N_21928);
xor U22834 (N_22834,N_21102,N_21655);
xor U22835 (N_22835,N_21490,N_21749);
nor U22836 (N_22836,N_21154,N_21604);
or U22837 (N_22837,N_21801,N_21834);
and U22838 (N_22838,N_21650,N_21864);
xnor U22839 (N_22839,N_21929,N_21720);
nand U22840 (N_22840,N_21030,N_21935);
nand U22841 (N_22841,N_21666,N_21118);
and U22842 (N_22842,N_21989,N_21221);
nand U22843 (N_22843,N_21160,N_21474);
xor U22844 (N_22844,N_21052,N_21921);
xor U22845 (N_22845,N_21358,N_21523);
xnor U22846 (N_22846,N_21986,N_21288);
xnor U22847 (N_22847,N_21125,N_21380);
nor U22848 (N_22848,N_21447,N_21404);
and U22849 (N_22849,N_21345,N_21266);
xnor U22850 (N_22850,N_21198,N_21732);
or U22851 (N_22851,N_21393,N_21780);
nor U22852 (N_22852,N_21146,N_21891);
or U22853 (N_22853,N_21785,N_21185);
nand U22854 (N_22854,N_21930,N_21119);
and U22855 (N_22855,N_21143,N_21944);
or U22856 (N_22856,N_21576,N_21367);
nor U22857 (N_22857,N_21843,N_21364);
and U22858 (N_22858,N_21181,N_21283);
and U22859 (N_22859,N_21376,N_21827);
and U22860 (N_22860,N_21559,N_21598);
nand U22861 (N_22861,N_21901,N_21702);
nor U22862 (N_22862,N_21451,N_21881);
or U22863 (N_22863,N_21716,N_21307);
nand U22864 (N_22864,N_21229,N_21146);
xor U22865 (N_22865,N_21498,N_21112);
and U22866 (N_22866,N_21408,N_21124);
nand U22867 (N_22867,N_21541,N_21641);
nor U22868 (N_22868,N_21833,N_21701);
xnor U22869 (N_22869,N_21370,N_21849);
and U22870 (N_22870,N_21146,N_21707);
xnor U22871 (N_22871,N_21061,N_21573);
or U22872 (N_22872,N_21376,N_21494);
or U22873 (N_22873,N_21214,N_21366);
nand U22874 (N_22874,N_21687,N_21632);
nor U22875 (N_22875,N_21094,N_21555);
and U22876 (N_22876,N_21406,N_21194);
xnor U22877 (N_22877,N_21700,N_21837);
nand U22878 (N_22878,N_21954,N_21488);
nor U22879 (N_22879,N_21354,N_21345);
and U22880 (N_22880,N_21701,N_21662);
or U22881 (N_22881,N_21776,N_21388);
nand U22882 (N_22882,N_21238,N_21981);
xnor U22883 (N_22883,N_21795,N_21746);
and U22884 (N_22884,N_21331,N_21163);
xor U22885 (N_22885,N_21887,N_21732);
nor U22886 (N_22886,N_21092,N_21832);
nand U22887 (N_22887,N_21528,N_21669);
and U22888 (N_22888,N_21625,N_21949);
nand U22889 (N_22889,N_21400,N_21548);
xor U22890 (N_22890,N_21607,N_21310);
and U22891 (N_22891,N_21001,N_21924);
nand U22892 (N_22892,N_21300,N_21343);
xnor U22893 (N_22893,N_21760,N_21743);
xnor U22894 (N_22894,N_21147,N_21748);
nor U22895 (N_22895,N_21807,N_21858);
and U22896 (N_22896,N_21373,N_21231);
nand U22897 (N_22897,N_21561,N_21394);
or U22898 (N_22898,N_21473,N_21422);
nand U22899 (N_22899,N_21273,N_21224);
xor U22900 (N_22900,N_21576,N_21365);
nor U22901 (N_22901,N_21417,N_21408);
and U22902 (N_22902,N_21172,N_21230);
and U22903 (N_22903,N_21515,N_21612);
nor U22904 (N_22904,N_21739,N_21744);
nor U22905 (N_22905,N_21170,N_21295);
or U22906 (N_22906,N_21254,N_21850);
or U22907 (N_22907,N_21197,N_21882);
nor U22908 (N_22908,N_21372,N_21360);
nand U22909 (N_22909,N_21168,N_21164);
or U22910 (N_22910,N_21871,N_21329);
xor U22911 (N_22911,N_21273,N_21766);
or U22912 (N_22912,N_21290,N_21125);
xor U22913 (N_22913,N_21380,N_21721);
and U22914 (N_22914,N_21289,N_21046);
and U22915 (N_22915,N_21250,N_21607);
nor U22916 (N_22916,N_21711,N_21444);
or U22917 (N_22917,N_21693,N_21507);
and U22918 (N_22918,N_21433,N_21174);
and U22919 (N_22919,N_21830,N_21762);
nor U22920 (N_22920,N_21071,N_21082);
nor U22921 (N_22921,N_21069,N_21492);
nand U22922 (N_22922,N_21728,N_21637);
nor U22923 (N_22923,N_21154,N_21932);
and U22924 (N_22924,N_21053,N_21402);
nor U22925 (N_22925,N_21866,N_21048);
or U22926 (N_22926,N_21378,N_21137);
and U22927 (N_22927,N_21419,N_21595);
nand U22928 (N_22928,N_21297,N_21796);
or U22929 (N_22929,N_21565,N_21507);
nand U22930 (N_22930,N_21018,N_21986);
xor U22931 (N_22931,N_21748,N_21984);
and U22932 (N_22932,N_21020,N_21075);
xnor U22933 (N_22933,N_21367,N_21945);
xnor U22934 (N_22934,N_21599,N_21629);
and U22935 (N_22935,N_21453,N_21892);
nand U22936 (N_22936,N_21938,N_21114);
nor U22937 (N_22937,N_21183,N_21032);
or U22938 (N_22938,N_21176,N_21055);
xor U22939 (N_22939,N_21816,N_21695);
or U22940 (N_22940,N_21009,N_21331);
nor U22941 (N_22941,N_21199,N_21015);
xnor U22942 (N_22942,N_21567,N_21554);
nand U22943 (N_22943,N_21954,N_21331);
xor U22944 (N_22944,N_21527,N_21292);
nor U22945 (N_22945,N_21134,N_21198);
and U22946 (N_22946,N_21315,N_21276);
and U22947 (N_22947,N_21373,N_21055);
and U22948 (N_22948,N_21757,N_21167);
xnor U22949 (N_22949,N_21803,N_21886);
and U22950 (N_22950,N_21283,N_21895);
xor U22951 (N_22951,N_21596,N_21012);
nor U22952 (N_22952,N_21889,N_21378);
nor U22953 (N_22953,N_21086,N_21257);
and U22954 (N_22954,N_21353,N_21070);
or U22955 (N_22955,N_21843,N_21504);
and U22956 (N_22956,N_21783,N_21426);
nor U22957 (N_22957,N_21240,N_21858);
and U22958 (N_22958,N_21093,N_21435);
and U22959 (N_22959,N_21413,N_21018);
xor U22960 (N_22960,N_21783,N_21647);
xor U22961 (N_22961,N_21642,N_21203);
xnor U22962 (N_22962,N_21530,N_21372);
xnor U22963 (N_22963,N_21694,N_21370);
nand U22964 (N_22964,N_21228,N_21408);
nor U22965 (N_22965,N_21640,N_21731);
nor U22966 (N_22966,N_21557,N_21426);
nor U22967 (N_22967,N_21975,N_21499);
nor U22968 (N_22968,N_21544,N_21363);
nor U22969 (N_22969,N_21091,N_21618);
nand U22970 (N_22970,N_21972,N_21684);
or U22971 (N_22971,N_21307,N_21308);
nand U22972 (N_22972,N_21755,N_21134);
or U22973 (N_22973,N_21514,N_21952);
nand U22974 (N_22974,N_21184,N_21071);
nand U22975 (N_22975,N_21851,N_21793);
nor U22976 (N_22976,N_21202,N_21864);
or U22977 (N_22977,N_21768,N_21944);
and U22978 (N_22978,N_21089,N_21369);
or U22979 (N_22979,N_21565,N_21222);
or U22980 (N_22980,N_21586,N_21045);
nand U22981 (N_22981,N_21838,N_21509);
xor U22982 (N_22982,N_21193,N_21093);
nor U22983 (N_22983,N_21618,N_21259);
and U22984 (N_22984,N_21931,N_21576);
nand U22985 (N_22985,N_21259,N_21658);
or U22986 (N_22986,N_21767,N_21796);
or U22987 (N_22987,N_21925,N_21658);
nor U22988 (N_22988,N_21013,N_21515);
nand U22989 (N_22989,N_21367,N_21896);
or U22990 (N_22990,N_21388,N_21068);
nand U22991 (N_22991,N_21160,N_21001);
nor U22992 (N_22992,N_21525,N_21230);
nor U22993 (N_22993,N_21721,N_21065);
and U22994 (N_22994,N_21642,N_21215);
and U22995 (N_22995,N_21871,N_21130);
nand U22996 (N_22996,N_21283,N_21844);
or U22997 (N_22997,N_21173,N_21503);
nor U22998 (N_22998,N_21519,N_21232);
nand U22999 (N_22999,N_21496,N_21851);
nand U23000 (N_23000,N_22331,N_22879);
or U23001 (N_23001,N_22136,N_22281);
or U23002 (N_23002,N_22716,N_22585);
or U23003 (N_23003,N_22721,N_22480);
nor U23004 (N_23004,N_22330,N_22777);
or U23005 (N_23005,N_22884,N_22176);
and U23006 (N_23006,N_22822,N_22905);
and U23007 (N_23007,N_22040,N_22044);
nand U23008 (N_23008,N_22260,N_22515);
nand U23009 (N_23009,N_22823,N_22850);
nor U23010 (N_23010,N_22987,N_22558);
nand U23011 (N_23011,N_22456,N_22144);
and U23012 (N_23012,N_22030,N_22848);
xnor U23013 (N_23013,N_22572,N_22403);
nor U23014 (N_23014,N_22396,N_22242);
nor U23015 (N_23015,N_22561,N_22781);
xnor U23016 (N_23016,N_22744,N_22697);
nand U23017 (N_23017,N_22195,N_22100);
xor U23018 (N_23018,N_22160,N_22730);
or U23019 (N_23019,N_22227,N_22996);
and U23020 (N_23020,N_22683,N_22601);
and U23021 (N_23021,N_22257,N_22593);
or U23022 (N_23022,N_22372,N_22285);
or U23023 (N_23023,N_22825,N_22941);
nor U23024 (N_23024,N_22115,N_22284);
and U23025 (N_23025,N_22663,N_22179);
and U23026 (N_23026,N_22741,N_22387);
nand U23027 (N_23027,N_22604,N_22971);
or U23028 (N_23028,N_22214,N_22643);
nand U23029 (N_23029,N_22117,N_22449);
nor U23030 (N_23030,N_22221,N_22889);
or U23031 (N_23031,N_22826,N_22321);
or U23032 (N_23032,N_22805,N_22090);
or U23033 (N_23033,N_22333,N_22288);
xor U23034 (N_23034,N_22525,N_22123);
xor U23035 (N_23035,N_22246,N_22279);
nand U23036 (N_23036,N_22578,N_22358);
nor U23037 (N_23037,N_22802,N_22484);
or U23038 (N_23038,N_22225,N_22896);
or U23039 (N_23039,N_22510,N_22014);
or U23040 (N_23040,N_22588,N_22171);
and U23041 (N_23041,N_22340,N_22230);
nand U23042 (N_23042,N_22064,N_22217);
xor U23043 (N_23043,N_22058,N_22363);
and U23044 (N_23044,N_22459,N_22674);
and U23045 (N_23045,N_22618,N_22133);
or U23046 (N_23046,N_22570,N_22218);
and U23047 (N_23047,N_22914,N_22019);
nor U23048 (N_23048,N_22175,N_22555);
nand U23049 (N_23049,N_22609,N_22569);
and U23050 (N_23050,N_22606,N_22617);
nand U23051 (N_23051,N_22845,N_22289);
or U23052 (N_23052,N_22745,N_22507);
nor U23053 (N_23053,N_22628,N_22912);
nand U23054 (N_23054,N_22297,N_22282);
or U23055 (N_23055,N_22167,N_22771);
nand U23056 (N_23056,N_22423,N_22792);
or U23057 (N_23057,N_22788,N_22046);
xnor U23058 (N_23058,N_22184,N_22587);
xor U23059 (N_23059,N_22471,N_22979);
nor U23060 (N_23060,N_22186,N_22296);
xor U23061 (N_23061,N_22003,N_22327);
nand U23062 (N_23062,N_22513,N_22390);
xor U23063 (N_23063,N_22549,N_22583);
nand U23064 (N_23064,N_22276,N_22371);
nand U23065 (N_23065,N_22215,N_22675);
nand U23066 (N_23066,N_22765,N_22841);
nand U23067 (N_23067,N_22840,N_22707);
nand U23068 (N_23068,N_22931,N_22473);
nor U23069 (N_23069,N_22520,N_22148);
and U23070 (N_23070,N_22667,N_22008);
nor U23071 (N_23071,N_22436,N_22581);
xor U23072 (N_23072,N_22997,N_22529);
nor U23073 (N_23073,N_22240,N_22020);
and U23074 (N_23074,N_22737,N_22669);
nand U23075 (N_23075,N_22178,N_22223);
nor U23076 (N_23076,N_22143,N_22145);
or U23077 (N_23077,N_22362,N_22075);
xor U23078 (N_23078,N_22277,N_22576);
nor U23079 (N_23079,N_22222,N_22047);
xnor U23080 (N_23080,N_22205,N_22154);
nor U23081 (N_23081,N_22901,N_22194);
nor U23082 (N_23082,N_22642,N_22665);
nand U23083 (N_23083,N_22259,N_22485);
nand U23084 (N_23084,N_22861,N_22092);
and U23085 (N_23085,N_22081,N_22342);
nor U23086 (N_23086,N_22174,N_22180);
xnor U23087 (N_23087,N_22334,N_22655);
xor U23088 (N_23088,N_22651,N_22932);
xor U23089 (N_23089,N_22798,N_22084);
or U23090 (N_23090,N_22873,N_22393);
xnor U23091 (N_23091,N_22349,N_22364);
nor U23092 (N_23092,N_22536,N_22063);
nand U23093 (N_23093,N_22943,N_22089);
nand U23094 (N_23094,N_22165,N_22768);
xnor U23095 (N_23095,N_22129,N_22368);
nor U23096 (N_23096,N_22374,N_22793);
nor U23097 (N_23097,N_22530,N_22164);
or U23098 (N_23098,N_22553,N_22658);
nand U23099 (N_23099,N_22468,N_22703);
or U23100 (N_23100,N_22859,N_22440);
nand U23101 (N_23101,N_22603,N_22018);
and U23102 (N_23102,N_22037,N_22237);
and U23103 (N_23103,N_22073,N_22649);
nor U23104 (N_23104,N_22815,N_22220);
nand U23105 (N_23105,N_22800,N_22016);
nor U23106 (N_23106,N_22489,N_22060);
or U23107 (N_23107,N_22447,N_22968);
or U23108 (N_23108,N_22827,N_22646);
and U23109 (N_23109,N_22397,N_22494);
and U23110 (N_23110,N_22162,N_22476);
nand U23111 (N_23111,N_22361,N_22672);
and U23112 (N_23112,N_22157,N_22776);
xnor U23113 (N_23113,N_22072,N_22865);
and U23114 (N_23114,N_22566,N_22543);
nor U23115 (N_23115,N_22954,N_22634);
nor U23116 (N_23116,N_22866,N_22808);
nand U23117 (N_23117,N_22273,N_22382);
xor U23118 (N_23118,N_22161,N_22487);
nand U23119 (N_23119,N_22657,N_22500);
or U23120 (N_23120,N_22355,N_22395);
nor U23121 (N_23121,N_22977,N_22066);
nor U23122 (N_23122,N_22211,N_22557);
nor U23123 (N_23123,N_22448,N_22424);
and U23124 (N_23124,N_22369,N_22614);
or U23125 (N_23125,N_22079,N_22263);
xor U23126 (N_23126,N_22883,N_22753);
nor U23127 (N_23127,N_22385,N_22109);
xnor U23128 (N_23128,N_22457,N_22735);
xor U23129 (N_23129,N_22252,N_22727);
nand U23130 (N_23130,N_22055,N_22465);
nand U23131 (N_23131,N_22376,N_22346);
nor U23132 (N_23132,N_22538,N_22758);
nor U23133 (N_23133,N_22034,N_22085);
nand U23134 (N_23134,N_22711,N_22812);
and U23135 (N_23135,N_22661,N_22907);
and U23136 (N_23136,N_22626,N_22314);
nand U23137 (N_23137,N_22036,N_22106);
and U23138 (N_23138,N_22300,N_22219);
xnor U23139 (N_23139,N_22769,N_22105);
or U23140 (N_23140,N_22107,N_22247);
nand U23141 (N_23141,N_22024,N_22291);
or U23142 (N_23142,N_22140,N_22904);
and U23143 (N_23143,N_22728,N_22560);
or U23144 (N_23144,N_22152,N_22607);
nor U23145 (N_23145,N_22233,N_22791);
nand U23146 (N_23146,N_22445,N_22173);
nand U23147 (N_23147,N_22130,N_22888);
xnor U23148 (N_23148,N_22622,N_22344);
and U23149 (N_23149,N_22189,N_22498);
nor U23150 (N_23150,N_22341,N_22691);
or U23151 (N_23151,N_22267,N_22653);
xnor U23152 (N_23152,N_22057,N_22128);
nor U23153 (N_23153,N_22563,N_22980);
nand U23154 (N_23154,N_22755,N_22097);
nand U23155 (N_23155,N_22989,N_22871);
xor U23156 (N_23156,N_22299,N_22415);
nor U23157 (N_23157,N_22295,N_22461);
nand U23158 (N_23158,N_22504,N_22261);
xor U23159 (N_23159,N_22935,N_22898);
nor U23160 (N_23160,N_22310,N_22354);
or U23161 (N_23161,N_22025,N_22293);
nand U23162 (N_23162,N_22837,N_22528);
nand U23163 (N_23163,N_22596,N_22146);
nand U23164 (N_23164,N_22937,N_22497);
nor U23165 (N_23165,N_22951,N_22973);
nand U23166 (N_23166,N_22113,N_22985);
xnor U23167 (N_23167,N_22431,N_22239);
nor U23168 (N_23168,N_22235,N_22104);
xnor U23169 (N_23169,N_22479,N_22481);
nor U23170 (N_23170,N_22645,N_22541);
xor U23171 (N_23171,N_22794,N_22615);
nor U23172 (N_23172,N_22894,N_22589);
or U23173 (N_23173,N_22212,N_22890);
and U23174 (N_23174,N_22590,N_22630);
xor U23175 (N_23175,N_22399,N_22947);
or U23176 (N_23176,N_22762,N_22686);
xnor U23177 (N_23177,N_22303,N_22469);
xor U23178 (N_23178,N_22417,N_22710);
nand U23179 (N_23179,N_22969,N_22595);
or U23180 (N_23180,N_22455,N_22023);
nand U23181 (N_23181,N_22842,N_22552);
xnor U23182 (N_23182,N_22118,N_22564);
or U23183 (N_23183,N_22992,N_22425);
nor U23184 (N_23184,N_22191,N_22013);
and U23185 (N_23185,N_22780,N_22704);
nand U23186 (N_23186,N_22982,N_22198);
and U23187 (N_23187,N_22656,N_22360);
nand U23188 (N_23188,N_22502,N_22574);
and U23189 (N_23189,N_22945,N_22681);
xnor U23190 (N_23190,N_22210,N_22463);
nand U23191 (N_23191,N_22389,N_22108);
nand U23192 (N_23192,N_22384,N_22268);
and U23193 (N_23193,N_22526,N_22648);
or U23194 (N_23194,N_22886,N_22168);
and U23195 (N_23195,N_22241,N_22501);
or U23196 (N_23196,N_22867,N_22957);
nand U23197 (N_23197,N_22633,N_22414);
nand U23198 (N_23198,N_22809,N_22814);
nor U23199 (N_23199,N_22472,N_22801);
and U23200 (N_23200,N_22357,N_22839);
nand U23201 (N_23201,N_22684,N_22482);
nor U23202 (N_23202,N_22673,N_22206);
and U23203 (N_23203,N_22994,N_22253);
and U23204 (N_23204,N_22880,N_22467);
nor U23205 (N_23205,N_22856,N_22820);
xor U23206 (N_23206,N_22203,N_22356);
and U23207 (N_23207,N_22616,N_22126);
and U23208 (N_23208,N_22742,N_22006);
and U23209 (N_23209,N_22610,N_22519);
nand U23210 (N_23210,N_22659,N_22668);
nand U23211 (N_23211,N_22045,N_22153);
or U23212 (N_23212,N_22627,N_22757);
nand U23213 (N_23213,N_22065,N_22620);
nor U23214 (N_23214,N_22517,N_22787);
or U23215 (N_23215,N_22591,N_22600);
xor U23216 (N_23216,N_22197,N_22111);
and U23217 (N_23217,N_22110,N_22038);
nor U23218 (N_23218,N_22015,N_22803);
xor U23219 (N_23219,N_22836,N_22895);
nand U23220 (N_23220,N_22682,N_22923);
nand U23221 (N_23221,N_22772,N_22920);
nor U23222 (N_23222,N_22554,N_22548);
or U23223 (N_23223,N_22725,N_22156);
or U23224 (N_23224,N_22204,N_22124);
nand U23225 (N_23225,N_22335,N_22244);
and U23226 (N_23226,N_22413,N_22767);
nand U23227 (N_23227,N_22302,N_22860);
and U23228 (N_23228,N_22408,N_22052);
or U23229 (N_23229,N_22470,N_22568);
xnor U23230 (N_23230,N_22067,N_22450);
or U23231 (N_23231,N_22187,N_22488);
nand U23232 (N_23232,N_22086,N_22854);
or U23233 (N_23233,N_22613,N_22720);
or U23234 (N_23234,N_22199,N_22407);
or U23235 (N_23235,N_22756,N_22512);
xor U23236 (N_23236,N_22005,N_22091);
nor U23237 (N_23237,N_22438,N_22849);
xor U23238 (N_23238,N_22714,N_22950);
nand U23239 (N_23239,N_22754,N_22995);
or U23240 (N_23240,N_22017,N_22311);
nand U23241 (N_23241,N_22934,N_22592);
nand U23242 (N_23242,N_22352,N_22773);
nand U23243 (N_23243,N_22275,N_22933);
and U23244 (N_23244,N_22004,N_22386);
or U23245 (N_23245,N_22690,N_22208);
xor U23246 (N_23246,N_22926,N_22453);
nand U23247 (N_23247,N_22200,N_22747);
nand U23248 (N_23248,N_22088,N_22676);
xnor U23249 (N_23249,N_22294,N_22007);
xnor U23250 (N_23250,N_22050,N_22598);
nor U23251 (N_23251,N_22158,N_22039);
nor U23252 (N_23252,N_22550,N_22444);
and U23253 (N_23253,N_22251,N_22292);
nand U23254 (N_23254,N_22694,N_22033);
nor U23255 (N_23255,N_22544,N_22492);
nor U23256 (N_23256,N_22817,N_22639);
xnor U23257 (N_23257,N_22636,N_22185);
and U23258 (N_23258,N_22192,N_22172);
xnor U23259 (N_23259,N_22427,N_22594);
nand U23260 (N_23260,N_22687,N_22435);
xor U23261 (N_23261,N_22775,N_22010);
nand U23262 (N_23262,N_22051,N_22011);
nor U23263 (N_23263,N_22567,N_22743);
xnor U23264 (N_23264,N_22316,N_22782);
nor U23265 (N_23265,N_22611,N_22764);
and U23266 (N_23266,N_22207,N_22759);
xor U23267 (N_23267,N_22324,N_22274);
nand U23268 (N_23268,N_22308,N_22692);
nand U23269 (N_23269,N_22723,N_22338);
and U23270 (N_23270,N_22083,N_22132);
nor U23271 (N_23271,N_22127,N_22584);
xnor U23272 (N_23272,N_22698,N_22786);
and U23273 (N_23273,N_22958,N_22232);
nor U23274 (N_23274,N_22851,N_22952);
nand U23275 (N_23275,N_22032,N_22542);
nor U23276 (N_23276,N_22307,N_22991);
or U23277 (N_23277,N_22437,N_22049);
xnor U23278 (N_23278,N_22422,N_22042);
nand U23279 (N_23279,N_22893,N_22751);
nor U23280 (N_23280,N_22434,N_22844);
and U23281 (N_23281,N_22093,N_22819);
and U23282 (N_23282,N_22795,N_22102);
and U23283 (N_23283,N_22891,N_22027);
nand U23284 (N_23284,N_22623,N_22832);
nand U23285 (N_23285,N_22406,N_22881);
xor U23286 (N_23286,N_22940,N_22428);
xnor U23287 (N_23287,N_22378,N_22163);
or U23288 (N_23288,N_22899,N_22121);
nor U23289 (N_23289,N_22999,N_22678);
and U23290 (N_23290,N_22970,N_22875);
or U23291 (N_23291,N_22579,N_22359);
xor U23292 (N_23292,N_22929,N_22580);
xnor U23293 (N_23293,N_22332,N_22347);
xnor U23294 (N_23294,N_22466,N_22551);
nand U23295 (N_23295,N_22712,N_22000);
nand U23296 (N_23296,N_22188,N_22892);
and U23297 (N_23297,N_22540,N_22224);
nor U23298 (N_23298,N_22229,N_22717);
nor U23299 (N_23299,N_22640,N_22068);
and U23300 (N_23300,N_22226,N_22821);
xor U23301 (N_23301,N_22625,N_22234);
or U23302 (N_23302,N_22608,N_22028);
nand U23303 (N_23303,N_22631,N_22421);
nand U23304 (N_23304,N_22029,N_22602);
xnor U23305 (N_23305,N_22831,N_22441);
nor U23306 (N_23306,N_22258,N_22975);
nand U23307 (N_23307,N_22026,N_22829);
and U23308 (N_23308,N_22597,N_22458);
xnor U23309 (N_23309,N_22779,N_22265);
and U23310 (N_23310,N_22443,N_22715);
nor U23311 (N_23311,N_22978,N_22412);
or U23312 (N_23312,N_22269,N_22546);
xnor U23313 (N_23313,N_22984,N_22002);
and U23314 (N_23314,N_22624,N_22924);
xor U23315 (N_23315,N_22706,N_22411);
nor U23316 (N_23316,N_22155,N_22981);
nor U23317 (N_23317,N_22280,N_22365);
xor U23318 (N_23318,N_22960,N_22953);
nand U23319 (N_23319,N_22695,N_22922);
or U23320 (N_23320,N_22909,N_22582);
or U23321 (N_23321,N_22320,N_22993);
nor U23322 (N_23322,N_22149,N_22317);
xor U23323 (N_23323,N_22719,N_22599);
and U23324 (N_23324,N_22547,N_22329);
or U23325 (N_23325,N_22370,N_22571);
xnor U23326 (N_23326,N_22539,N_22278);
xor U23327 (N_23327,N_22936,N_22043);
or U23328 (N_23328,N_22381,N_22699);
nor U23329 (N_23329,N_22054,N_22847);
xnor U23330 (N_23330,N_22664,N_22182);
xnor U23331 (N_23331,N_22159,N_22677);
xor U23332 (N_23332,N_22243,N_22974);
xor U23333 (N_23333,N_22972,N_22784);
nand U23334 (N_23334,N_22420,N_22323);
xnor U23335 (N_23335,N_22789,N_22141);
xor U23336 (N_23336,N_22731,N_22913);
nand U23337 (N_23337,N_22647,N_22442);
and U23338 (N_23338,N_22287,N_22071);
nor U23339 (N_23339,N_22729,N_22496);
nand U23340 (N_23340,N_22967,N_22897);
or U23341 (N_23341,N_22760,N_22309);
nand U23342 (N_23342,N_22418,N_22919);
and U23343 (N_23343,N_22505,N_22722);
or U23344 (N_23344,N_22948,N_22652);
nor U23345 (N_23345,N_22988,N_22116);
or U23346 (N_23346,N_22521,N_22125);
or U23347 (N_23347,N_22120,N_22961);
nor U23348 (N_23348,N_22325,N_22048);
nand U23349 (N_23349,N_22245,N_22486);
and U23350 (N_23350,N_22946,N_22377);
or U23351 (N_23351,N_22343,N_22870);
and U23352 (N_23352,N_22353,N_22575);
nand U23353 (N_23353,N_22499,N_22433);
nor U23354 (N_23354,N_22070,N_22404);
and U23355 (N_23355,N_22766,N_22254);
and U23356 (N_23356,N_22740,N_22119);
xor U23357 (N_23357,N_22925,N_22761);
and U23358 (N_23358,N_22493,N_22375);
nor U23359 (N_23359,N_22074,N_22490);
nand U23360 (N_23360,N_22451,N_22545);
and U23361 (N_23361,N_22900,N_22533);
or U23362 (N_23362,N_22351,N_22949);
nand U23363 (N_23363,N_22348,N_22078);
nor U23364 (N_23364,N_22990,N_22394);
xor U23365 (N_23365,N_22477,N_22059);
or U23366 (N_23366,N_22738,N_22270);
nand U23367 (N_23367,N_22565,N_22495);
xnor U23368 (N_23368,N_22965,N_22213);
and U23369 (N_23369,N_22885,N_22882);
xor U23370 (N_23370,N_22855,N_22400);
or U23371 (N_23371,N_22577,N_22910);
nor U23372 (N_23372,N_22290,N_22514);
and U23373 (N_23373,N_22852,N_22619);
and U23374 (N_23374,N_22231,N_22650);
and U23375 (N_23375,N_22662,N_22264);
nor U23376 (N_23376,N_22373,N_22306);
nand U23377 (N_23377,N_22138,N_22432);
nor U23378 (N_23378,N_22518,N_22644);
or U23379 (N_23379,N_22887,N_22478);
nor U23380 (N_23380,N_22464,N_22535);
or U23381 (N_23381,N_22062,N_22452);
or U23382 (N_23382,N_22266,N_22419);
xor U23383 (N_23383,N_22405,N_22137);
nand U23384 (N_23384,N_22638,N_22559);
nor U23385 (N_23385,N_22022,N_22916);
or U23386 (N_23386,N_22315,N_22304);
or U23387 (N_23387,N_22098,N_22439);
or U23388 (N_23388,N_22878,N_22483);
xnor U23389 (N_23389,N_22903,N_22379);
or U23390 (N_23390,N_22928,N_22056);
nand U23391 (N_23391,N_22523,N_22053);
xnor U23392 (N_23392,N_22401,N_22632);
xor U23393 (N_23393,N_22862,N_22688);
and U23394 (N_23394,N_22021,N_22209);
or U23395 (N_23395,N_22001,N_22818);
nor U23396 (N_23396,N_22193,N_22956);
nor U23397 (N_23397,N_22702,N_22524);
nand U23398 (N_23398,N_22748,N_22562);
xor U23399 (N_23399,N_22475,N_22286);
xor U23400 (N_23400,N_22828,N_22305);
nand U23401 (N_23401,N_22312,N_22183);
xnor U23402 (N_23402,N_22135,N_22696);
and U23403 (N_23403,N_22012,N_22076);
and U23404 (N_23404,N_22508,N_22170);
xnor U23405 (N_23405,N_22637,N_22701);
and U23406 (N_23406,N_22537,N_22556);
and U23407 (N_23407,N_22942,N_22778);
nor U23408 (N_23408,N_22713,N_22868);
xnor U23409 (N_23409,N_22087,N_22061);
nor U23410 (N_23410,N_22454,N_22586);
nor U23411 (N_23411,N_22804,N_22734);
nand U23412 (N_23412,N_22750,N_22122);
nand U23413 (N_23413,N_22446,N_22196);
xor U23414 (N_23414,N_22749,N_22770);
or U23415 (N_23415,N_22383,N_22095);
and U23416 (N_23416,N_22635,N_22460);
nand U23417 (N_23417,N_22705,N_22816);
xor U23418 (N_23418,N_22534,N_22392);
nor U23419 (N_23419,N_22660,N_22917);
or U23420 (N_23420,N_22732,N_22918);
xor U23421 (N_23421,N_22236,N_22746);
nand U23422 (N_23422,N_22838,N_22774);
and U23423 (N_23423,N_22983,N_22339);
xnor U23424 (N_23424,N_22248,N_22228);
nor U23425 (N_23425,N_22906,N_22272);
nand U23426 (N_23426,N_22255,N_22326);
or U23427 (N_23427,N_22134,N_22872);
and U23428 (N_23428,N_22201,N_22491);
and U23429 (N_23429,N_22573,N_22966);
nand U23430 (N_23430,N_22921,N_22939);
nor U23431 (N_23431,N_22398,N_22319);
and U23432 (N_23432,N_22077,N_22874);
or U23433 (N_23433,N_22824,N_22938);
xnor U23434 (N_23434,N_22430,N_22689);
or U23435 (N_23435,N_22009,N_22834);
and U23436 (N_23436,N_22959,N_22930);
xnor U23437 (N_23437,N_22797,N_22301);
nor U23438 (N_23438,N_22151,N_22869);
or U23439 (N_23439,N_22944,N_22752);
xor U23440 (N_23440,N_22336,N_22328);
or U23441 (N_23441,N_22709,N_22641);
xor U23442 (N_23442,N_22503,N_22096);
and U23443 (N_23443,N_22718,N_22216);
and U23444 (N_23444,N_22511,N_22806);
xor U23445 (N_23445,N_22256,N_22864);
or U23446 (N_23446,N_22531,N_22671);
and U23447 (N_23447,N_22366,N_22739);
nand U23448 (N_23448,N_22283,N_22736);
and U23449 (N_23449,N_22666,N_22114);
and U23450 (N_23450,N_22955,N_22846);
and U23451 (N_23451,N_22041,N_22629);
nor U23452 (N_23452,N_22835,N_22733);
nand U23453 (N_23453,N_22103,N_22313);
nor U23454 (N_23454,N_22876,N_22612);
nor U23455 (N_23455,N_22250,N_22262);
nand U23456 (N_23456,N_22853,N_22506);
nor U23457 (N_23457,N_22345,N_22877);
nand U23458 (N_23458,N_22147,N_22131);
nor U23459 (N_23459,N_22976,N_22318);
or U23460 (N_23460,N_22799,N_22783);
and U23461 (N_23461,N_22142,N_22388);
xnor U23462 (N_23462,N_22190,N_22249);
or U23463 (N_23463,N_22679,N_22810);
or U23464 (N_23464,N_22426,N_22962);
or U23465 (N_23465,N_22911,N_22915);
or U23466 (N_23466,N_22685,N_22654);
xor U23467 (N_23467,N_22509,N_22708);
nand U23468 (N_23468,N_22522,N_22830);
or U23469 (N_23469,N_22474,N_22350);
and U23470 (N_23470,N_22169,N_22843);
and U23471 (N_23471,N_22516,N_22409);
xor U23472 (N_23472,N_22857,N_22670);
or U23473 (N_23473,N_22532,N_22693);
xnor U23474 (N_23474,N_22271,N_22202);
xor U23475 (N_23475,N_22700,N_22367);
xnor U23476 (N_23476,N_22166,N_22031);
nor U23477 (N_23477,N_22462,N_22402);
and U23478 (N_23478,N_22391,N_22380);
nand U23479 (N_23479,N_22927,N_22527);
nand U23480 (N_23480,N_22986,N_22908);
or U23481 (N_23481,N_22069,N_22101);
nor U23482 (N_23482,N_22790,N_22082);
and U23483 (N_23483,N_22998,N_22785);
nand U23484 (N_23484,N_22902,N_22337);
xnor U23485 (N_23485,N_22035,N_22833);
nor U23486 (N_23486,N_22099,N_22680);
nor U23487 (N_23487,N_22863,N_22080);
nor U23488 (N_23488,N_22322,N_22763);
and U23489 (N_23489,N_22605,N_22858);
nor U23490 (N_23490,N_22181,N_22811);
or U23491 (N_23491,N_22724,N_22429);
or U23492 (N_23492,N_22410,N_22726);
xnor U23493 (N_23493,N_22094,N_22416);
or U23494 (N_23494,N_22964,N_22139);
nor U23495 (N_23495,N_22177,N_22807);
or U23496 (N_23496,N_22112,N_22238);
nand U23497 (N_23497,N_22150,N_22298);
nand U23498 (N_23498,N_22621,N_22796);
nand U23499 (N_23499,N_22963,N_22813);
or U23500 (N_23500,N_22832,N_22145);
or U23501 (N_23501,N_22267,N_22610);
and U23502 (N_23502,N_22604,N_22780);
nand U23503 (N_23503,N_22650,N_22540);
xor U23504 (N_23504,N_22130,N_22067);
xnor U23505 (N_23505,N_22631,N_22923);
xnor U23506 (N_23506,N_22482,N_22237);
and U23507 (N_23507,N_22952,N_22602);
xor U23508 (N_23508,N_22401,N_22898);
xnor U23509 (N_23509,N_22613,N_22893);
xnor U23510 (N_23510,N_22750,N_22446);
or U23511 (N_23511,N_22141,N_22030);
nor U23512 (N_23512,N_22625,N_22779);
nand U23513 (N_23513,N_22419,N_22248);
nand U23514 (N_23514,N_22053,N_22347);
and U23515 (N_23515,N_22343,N_22462);
or U23516 (N_23516,N_22693,N_22880);
or U23517 (N_23517,N_22951,N_22485);
nor U23518 (N_23518,N_22284,N_22931);
and U23519 (N_23519,N_22888,N_22640);
xnor U23520 (N_23520,N_22285,N_22241);
or U23521 (N_23521,N_22234,N_22934);
or U23522 (N_23522,N_22146,N_22000);
or U23523 (N_23523,N_22820,N_22374);
xnor U23524 (N_23524,N_22595,N_22258);
nor U23525 (N_23525,N_22134,N_22292);
and U23526 (N_23526,N_22808,N_22450);
nand U23527 (N_23527,N_22736,N_22730);
and U23528 (N_23528,N_22211,N_22309);
and U23529 (N_23529,N_22744,N_22438);
nand U23530 (N_23530,N_22231,N_22969);
and U23531 (N_23531,N_22122,N_22431);
and U23532 (N_23532,N_22758,N_22477);
nor U23533 (N_23533,N_22430,N_22518);
nand U23534 (N_23534,N_22533,N_22686);
or U23535 (N_23535,N_22950,N_22615);
nand U23536 (N_23536,N_22302,N_22720);
or U23537 (N_23537,N_22344,N_22764);
xor U23538 (N_23538,N_22964,N_22755);
or U23539 (N_23539,N_22074,N_22540);
nor U23540 (N_23540,N_22285,N_22478);
or U23541 (N_23541,N_22591,N_22300);
or U23542 (N_23542,N_22339,N_22151);
xnor U23543 (N_23543,N_22575,N_22070);
and U23544 (N_23544,N_22974,N_22318);
xor U23545 (N_23545,N_22897,N_22453);
nor U23546 (N_23546,N_22236,N_22277);
and U23547 (N_23547,N_22944,N_22339);
nor U23548 (N_23548,N_22976,N_22325);
or U23549 (N_23549,N_22029,N_22662);
nor U23550 (N_23550,N_22717,N_22259);
or U23551 (N_23551,N_22986,N_22542);
or U23552 (N_23552,N_22591,N_22744);
nand U23553 (N_23553,N_22292,N_22937);
or U23554 (N_23554,N_22079,N_22250);
xnor U23555 (N_23555,N_22649,N_22663);
nor U23556 (N_23556,N_22202,N_22150);
nand U23557 (N_23557,N_22338,N_22266);
or U23558 (N_23558,N_22205,N_22513);
or U23559 (N_23559,N_22943,N_22808);
nand U23560 (N_23560,N_22332,N_22044);
nand U23561 (N_23561,N_22116,N_22813);
or U23562 (N_23562,N_22524,N_22256);
or U23563 (N_23563,N_22012,N_22272);
xnor U23564 (N_23564,N_22811,N_22159);
nor U23565 (N_23565,N_22703,N_22171);
xnor U23566 (N_23566,N_22794,N_22798);
nand U23567 (N_23567,N_22648,N_22973);
and U23568 (N_23568,N_22398,N_22942);
or U23569 (N_23569,N_22515,N_22354);
xor U23570 (N_23570,N_22492,N_22836);
xnor U23571 (N_23571,N_22821,N_22918);
nand U23572 (N_23572,N_22245,N_22297);
or U23573 (N_23573,N_22357,N_22181);
nor U23574 (N_23574,N_22385,N_22127);
nand U23575 (N_23575,N_22711,N_22082);
or U23576 (N_23576,N_22330,N_22493);
and U23577 (N_23577,N_22572,N_22173);
nor U23578 (N_23578,N_22884,N_22064);
nand U23579 (N_23579,N_22212,N_22456);
or U23580 (N_23580,N_22422,N_22598);
nand U23581 (N_23581,N_22468,N_22455);
nand U23582 (N_23582,N_22497,N_22736);
xor U23583 (N_23583,N_22545,N_22165);
nor U23584 (N_23584,N_22942,N_22277);
or U23585 (N_23585,N_22841,N_22322);
and U23586 (N_23586,N_22853,N_22190);
and U23587 (N_23587,N_22323,N_22942);
nand U23588 (N_23588,N_22829,N_22837);
or U23589 (N_23589,N_22520,N_22001);
or U23590 (N_23590,N_22647,N_22863);
or U23591 (N_23591,N_22032,N_22949);
nand U23592 (N_23592,N_22631,N_22256);
xor U23593 (N_23593,N_22197,N_22350);
nor U23594 (N_23594,N_22094,N_22404);
nor U23595 (N_23595,N_22165,N_22229);
and U23596 (N_23596,N_22512,N_22129);
nor U23597 (N_23597,N_22143,N_22674);
xnor U23598 (N_23598,N_22755,N_22159);
and U23599 (N_23599,N_22356,N_22596);
nand U23600 (N_23600,N_22052,N_22527);
and U23601 (N_23601,N_22396,N_22025);
or U23602 (N_23602,N_22301,N_22142);
or U23603 (N_23603,N_22027,N_22160);
xnor U23604 (N_23604,N_22404,N_22313);
nor U23605 (N_23605,N_22955,N_22055);
or U23606 (N_23606,N_22534,N_22985);
or U23607 (N_23607,N_22210,N_22620);
and U23608 (N_23608,N_22121,N_22209);
xnor U23609 (N_23609,N_22273,N_22099);
nand U23610 (N_23610,N_22282,N_22166);
or U23611 (N_23611,N_22937,N_22059);
or U23612 (N_23612,N_22628,N_22354);
or U23613 (N_23613,N_22256,N_22068);
and U23614 (N_23614,N_22789,N_22928);
xnor U23615 (N_23615,N_22578,N_22075);
and U23616 (N_23616,N_22311,N_22104);
nor U23617 (N_23617,N_22968,N_22573);
nand U23618 (N_23618,N_22494,N_22523);
or U23619 (N_23619,N_22231,N_22265);
nor U23620 (N_23620,N_22056,N_22696);
nor U23621 (N_23621,N_22067,N_22147);
nand U23622 (N_23622,N_22978,N_22608);
nand U23623 (N_23623,N_22814,N_22745);
xnor U23624 (N_23624,N_22765,N_22348);
nor U23625 (N_23625,N_22983,N_22009);
xnor U23626 (N_23626,N_22111,N_22488);
and U23627 (N_23627,N_22489,N_22042);
nor U23628 (N_23628,N_22259,N_22316);
nand U23629 (N_23629,N_22002,N_22532);
nand U23630 (N_23630,N_22666,N_22130);
nand U23631 (N_23631,N_22292,N_22651);
xor U23632 (N_23632,N_22965,N_22756);
nor U23633 (N_23633,N_22870,N_22527);
and U23634 (N_23634,N_22819,N_22169);
or U23635 (N_23635,N_22851,N_22752);
and U23636 (N_23636,N_22255,N_22482);
or U23637 (N_23637,N_22043,N_22161);
nand U23638 (N_23638,N_22140,N_22022);
nand U23639 (N_23639,N_22457,N_22822);
or U23640 (N_23640,N_22515,N_22330);
and U23641 (N_23641,N_22976,N_22143);
nor U23642 (N_23642,N_22641,N_22204);
nor U23643 (N_23643,N_22848,N_22988);
nand U23644 (N_23644,N_22759,N_22637);
and U23645 (N_23645,N_22686,N_22830);
and U23646 (N_23646,N_22726,N_22821);
xnor U23647 (N_23647,N_22635,N_22809);
nor U23648 (N_23648,N_22734,N_22256);
xor U23649 (N_23649,N_22355,N_22068);
nor U23650 (N_23650,N_22440,N_22155);
xor U23651 (N_23651,N_22940,N_22033);
nor U23652 (N_23652,N_22433,N_22556);
or U23653 (N_23653,N_22022,N_22002);
and U23654 (N_23654,N_22671,N_22185);
or U23655 (N_23655,N_22634,N_22829);
or U23656 (N_23656,N_22872,N_22393);
or U23657 (N_23657,N_22538,N_22484);
xnor U23658 (N_23658,N_22003,N_22035);
or U23659 (N_23659,N_22591,N_22692);
or U23660 (N_23660,N_22778,N_22704);
xnor U23661 (N_23661,N_22654,N_22676);
nor U23662 (N_23662,N_22626,N_22107);
or U23663 (N_23663,N_22284,N_22775);
nand U23664 (N_23664,N_22140,N_22669);
xnor U23665 (N_23665,N_22289,N_22081);
nand U23666 (N_23666,N_22388,N_22888);
or U23667 (N_23667,N_22246,N_22133);
and U23668 (N_23668,N_22053,N_22604);
or U23669 (N_23669,N_22484,N_22955);
nand U23670 (N_23670,N_22135,N_22927);
xor U23671 (N_23671,N_22260,N_22616);
and U23672 (N_23672,N_22754,N_22188);
xnor U23673 (N_23673,N_22149,N_22949);
nand U23674 (N_23674,N_22461,N_22456);
and U23675 (N_23675,N_22058,N_22696);
xnor U23676 (N_23676,N_22269,N_22909);
xnor U23677 (N_23677,N_22735,N_22529);
nor U23678 (N_23678,N_22454,N_22913);
xor U23679 (N_23679,N_22015,N_22044);
nor U23680 (N_23680,N_22643,N_22650);
or U23681 (N_23681,N_22734,N_22541);
xnor U23682 (N_23682,N_22936,N_22108);
or U23683 (N_23683,N_22378,N_22570);
nand U23684 (N_23684,N_22894,N_22397);
nand U23685 (N_23685,N_22684,N_22008);
and U23686 (N_23686,N_22025,N_22674);
and U23687 (N_23687,N_22821,N_22086);
xnor U23688 (N_23688,N_22265,N_22961);
nor U23689 (N_23689,N_22292,N_22505);
xor U23690 (N_23690,N_22716,N_22120);
nor U23691 (N_23691,N_22810,N_22441);
or U23692 (N_23692,N_22141,N_22398);
and U23693 (N_23693,N_22143,N_22857);
nand U23694 (N_23694,N_22209,N_22840);
and U23695 (N_23695,N_22228,N_22059);
or U23696 (N_23696,N_22149,N_22988);
or U23697 (N_23697,N_22953,N_22435);
and U23698 (N_23698,N_22321,N_22432);
and U23699 (N_23699,N_22625,N_22810);
xor U23700 (N_23700,N_22636,N_22127);
nand U23701 (N_23701,N_22680,N_22916);
xor U23702 (N_23702,N_22079,N_22038);
xnor U23703 (N_23703,N_22756,N_22197);
or U23704 (N_23704,N_22883,N_22060);
nand U23705 (N_23705,N_22636,N_22364);
nand U23706 (N_23706,N_22630,N_22107);
and U23707 (N_23707,N_22340,N_22629);
xnor U23708 (N_23708,N_22664,N_22772);
nor U23709 (N_23709,N_22408,N_22794);
nor U23710 (N_23710,N_22056,N_22149);
nand U23711 (N_23711,N_22578,N_22194);
xnor U23712 (N_23712,N_22932,N_22428);
or U23713 (N_23713,N_22918,N_22942);
nor U23714 (N_23714,N_22905,N_22602);
and U23715 (N_23715,N_22953,N_22782);
and U23716 (N_23716,N_22265,N_22987);
nand U23717 (N_23717,N_22655,N_22868);
nor U23718 (N_23718,N_22323,N_22724);
nand U23719 (N_23719,N_22389,N_22924);
or U23720 (N_23720,N_22769,N_22775);
or U23721 (N_23721,N_22967,N_22015);
xnor U23722 (N_23722,N_22403,N_22158);
xnor U23723 (N_23723,N_22223,N_22037);
nand U23724 (N_23724,N_22115,N_22100);
and U23725 (N_23725,N_22693,N_22612);
or U23726 (N_23726,N_22206,N_22371);
and U23727 (N_23727,N_22254,N_22560);
nor U23728 (N_23728,N_22967,N_22697);
nand U23729 (N_23729,N_22698,N_22249);
nand U23730 (N_23730,N_22942,N_22051);
or U23731 (N_23731,N_22719,N_22860);
and U23732 (N_23732,N_22398,N_22278);
nand U23733 (N_23733,N_22800,N_22351);
and U23734 (N_23734,N_22281,N_22622);
nand U23735 (N_23735,N_22888,N_22817);
or U23736 (N_23736,N_22223,N_22224);
nor U23737 (N_23737,N_22486,N_22693);
nand U23738 (N_23738,N_22606,N_22812);
nand U23739 (N_23739,N_22521,N_22946);
nand U23740 (N_23740,N_22630,N_22103);
or U23741 (N_23741,N_22302,N_22509);
xor U23742 (N_23742,N_22277,N_22979);
or U23743 (N_23743,N_22306,N_22201);
nor U23744 (N_23744,N_22488,N_22224);
or U23745 (N_23745,N_22291,N_22479);
xnor U23746 (N_23746,N_22410,N_22678);
xnor U23747 (N_23747,N_22575,N_22727);
or U23748 (N_23748,N_22775,N_22715);
nor U23749 (N_23749,N_22034,N_22376);
nor U23750 (N_23750,N_22712,N_22123);
nand U23751 (N_23751,N_22385,N_22827);
nor U23752 (N_23752,N_22202,N_22074);
nor U23753 (N_23753,N_22747,N_22673);
and U23754 (N_23754,N_22279,N_22996);
and U23755 (N_23755,N_22944,N_22891);
nand U23756 (N_23756,N_22795,N_22620);
xnor U23757 (N_23757,N_22394,N_22724);
xor U23758 (N_23758,N_22057,N_22385);
nor U23759 (N_23759,N_22753,N_22074);
and U23760 (N_23760,N_22075,N_22147);
or U23761 (N_23761,N_22433,N_22015);
xor U23762 (N_23762,N_22005,N_22269);
nand U23763 (N_23763,N_22439,N_22976);
nor U23764 (N_23764,N_22832,N_22541);
and U23765 (N_23765,N_22569,N_22671);
and U23766 (N_23766,N_22012,N_22058);
nand U23767 (N_23767,N_22198,N_22156);
nor U23768 (N_23768,N_22070,N_22178);
nor U23769 (N_23769,N_22742,N_22398);
and U23770 (N_23770,N_22642,N_22745);
xnor U23771 (N_23771,N_22134,N_22679);
nand U23772 (N_23772,N_22195,N_22557);
xnor U23773 (N_23773,N_22646,N_22582);
xnor U23774 (N_23774,N_22521,N_22559);
xnor U23775 (N_23775,N_22084,N_22495);
or U23776 (N_23776,N_22893,N_22172);
nand U23777 (N_23777,N_22268,N_22206);
xor U23778 (N_23778,N_22606,N_22409);
and U23779 (N_23779,N_22761,N_22876);
xor U23780 (N_23780,N_22621,N_22204);
xnor U23781 (N_23781,N_22182,N_22794);
nand U23782 (N_23782,N_22785,N_22514);
nand U23783 (N_23783,N_22785,N_22240);
or U23784 (N_23784,N_22749,N_22454);
nor U23785 (N_23785,N_22148,N_22555);
nor U23786 (N_23786,N_22265,N_22781);
xor U23787 (N_23787,N_22931,N_22125);
or U23788 (N_23788,N_22061,N_22191);
nor U23789 (N_23789,N_22001,N_22891);
and U23790 (N_23790,N_22150,N_22426);
and U23791 (N_23791,N_22442,N_22554);
xnor U23792 (N_23792,N_22832,N_22173);
nand U23793 (N_23793,N_22776,N_22650);
or U23794 (N_23794,N_22346,N_22747);
nand U23795 (N_23795,N_22447,N_22379);
nand U23796 (N_23796,N_22110,N_22321);
and U23797 (N_23797,N_22001,N_22281);
nand U23798 (N_23798,N_22791,N_22686);
nor U23799 (N_23799,N_22599,N_22986);
nor U23800 (N_23800,N_22103,N_22141);
nor U23801 (N_23801,N_22325,N_22161);
or U23802 (N_23802,N_22110,N_22285);
and U23803 (N_23803,N_22273,N_22416);
or U23804 (N_23804,N_22562,N_22821);
or U23805 (N_23805,N_22451,N_22671);
nor U23806 (N_23806,N_22160,N_22896);
or U23807 (N_23807,N_22897,N_22425);
and U23808 (N_23808,N_22297,N_22368);
nand U23809 (N_23809,N_22257,N_22470);
and U23810 (N_23810,N_22155,N_22381);
nand U23811 (N_23811,N_22571,N_22655);
nor U23812 (N_23812,N_22570,N_22512);
or U23813 (N_23813,N_22730,N_22912);
nor U23814 (N_23814,N_22693,N_22116);
xnor U23815 (N_23815,N_22381,N_22886);
or U23816 (N_23816,N_22018,N_22132);
nor U23817 (N_23817,N_22287,N_22674);
nand U23818 (N_23818,N_22718,N_22277);
xnor U23819 (N_23819,N_22814,N_22833);
and U23820 (N_23820,N_22975,N_22972);
or U23821 (N_23821,N_22066,N_22001);
nand U23822 (N_23822,N_22258,N_22908);
nor U23823 (N_23823,N_22563,N_22405);
nor U23824 (N_23824,N_22527,N_22592);
nand U23825 (N_23825,N_22208,N_22862);
nand U23826 (N_23826,N_22476,N_22406);
or U23827 (N_23827,N_22230,N_22809);
or U23828 (N_23828,N_22127,N_22329);
or U23829 (N_23829,N_22764,N_22453);
nor U23830 (N_23830,N_22661,N_22571);
xnor U23831 (N_23831,N_22831,N_22478);
and U23832 (N_23832,N_22863,N_22758);
and U23833 (N_23833,N_22523,N_22273);
nand U23834 (N_23834,N_22712,N_22449);
and U23835 (N_23835,N_22540,N_22257);
or U23836 (N_23836,N_22248,N_22986);
nor U23837 (N_23837,N_22042,N_22591);
and U23838 (N_23838,N_22224,N_22744);
and U23839 (N_23839,N_22280,N_22319);
nand U23840 (N_23840,N_22383,N_22099);
nand U23841 (N_23841,N_22139,N_22865);
nor U23842 (N_23842,N_22629,N_22852);
nor U23843 (N_23843,N_22738,N_22700);
xor U23844 (N_23844,N_22928,N_22073);
or U23845 (N_23845,N_22458,N_22194);
nor U23846 (N_23846,N_22318,N_22046);
nor U23847 (N_23847,N_22563,N_22041);
and U23848 (N_23848,N_22253,N_22478);
nor U23849 (N_23849,N_22708,N_22294);
or U23850 (N_23850,N_22003,N_22959);
nor U23851 (N_23851,N_22917,N_22725);
xnor U23852 (N_23852,N_22308,N_22543);
nor U23853 (N_23853,N_22134,N_22628);
and U23854 (N_23854,N_22923,N_22403);
or U23855 (N_23855,N_22673,N_22146);
or U23856 (N_23856,N_22515,N_22894);
xnor U23857 (N_23857,N_22939,N_22882);
nand U23858 (N_23858,N_22793,N_22265);
nor U23859 (N_23859,N_22924,N_22043);
and U23860 (N_23860,N_22885,N_22298);
and U23861 (N_23861,N_22572,N_22507);
nand U23862 (N_23862,N_22966,N_22619);
and U23863 (N_23863,N_22956,N_22109);
xnor U23864 (N_23864,N_22358,N_22223);
nor U23865 (N_23865,N_22416,N_22380);
nand U23866 (N_23866,N_22873,N_22510);
xor U23867 (N_23867,N_22492,N_22049);
xor U23868 (N_23868,N_22841,N_22948);
and U23869 (N_23869,N_22303,N_22791);
nand U23870 (N_23870,N_22653,N_22743);
xor U23871 (N_23871,N_22814,N_22491);
or U23872 (N_23872,N_22508,N_22415);
or U23873 (N_23873,N_22823,N_22520);
xor U23874 (N_23874,N_22972,N_22608);
or U23875 (N_23875,N_22556,N_22895);
nor U23876 (N_23876,N_22509,N_22498);
xor U23877 (N_23877,N_22295,N_22763);
nor U23878 (N_23878,N_22773,N_22454);
nand U23879 (N_23879,N_22192,N_22769);
and U23880 (N_23880,N_22067,N_22292);
xnor U23881 (N_23881,N_22838,N_22594);
or U23882 (N_23882,N_22010,N_22278);
nand U23883 (N_23883,N_22670,N_22902);
and U23884 (N_23884,N_22606,N_22058);
nor U23885 (N_23885,N_22035,N_22555);
nor U23886 (N_23886,N_22411,N_22944);
nand U23887 (N_23887,N_22136,N_22530);
nand U23888 (N_23888,N_22431,N_22924);
nand U23889 (N_23889,N_22344,N_22298);
and U23890 (N_23890,N_22817,N_22942);
xnor U23891 (N_23891,N_22772,N_22016);
xor U23892 (N_23892,N_22350,N_22475);
nor U23893 (N_23893,N_22559,N_22577);
and U23894 (N_23894,N_22247,N_22044);
and U23895 (N_23895,N_22189,N_22737);
xor U23896 (N_23896,N_22480,N_22147);
or U23897 (N_23897,N_22526,N_22680);
nor U23898 (N_23898,N_22377,N_22236);
xnor U23899 (N_23899,N_22280,N_22044);
xnor U23900 (N_23900,N_22305,N_22621);
or U23901 (N_23901,N_22550,N_22710);
nor U23902 (N_23902,N_22293,N_22839);
xnor U23903 (N_23903,N_22968,N_22719);
nand U23904 (N_23904,N_22410,N_22943);
or U23905 (N_23905,N_22164,N_22446);
and U23906 (N_23906,N_22823,N_22233);
or U23907 (N_23907,N_22756,N_22277);
and U23908 (N_23908,N_22279,N_22694);
or U23909 (N_23909,N_22876,N_22686);
and U23910 (N_23910,N_22994,N_22949);
nand U23911 (N_23911,N_22696,N_22744);
nor U23912 (N_23912,N_22871,N_22190);
nand U23913 (N_23913,N_22050,N_22365);
nand U23914 (N_23914,N_22812,N_22867);
and U23915 (N_23915,N_22422,N_22738);
nor U23916 (N_23916,N_22201,N_22627);
xor U23917 (N_23917,N_22654,N_22168);
or U23918 (N_23918,N_22034,N_22073);
nand U23919 (N_23919,N_22038,N_22434);
or U23920 (N_23920,N_22939,N_22191);
or U23921 (N_23921,N_22487,N_22734);
or U23922 (N_23922,N_22011,N_22479);
nand U23923 (N_23923,N_22640,N_22037);
xnor U23924 (N_23924,N_22996,N_22806);
and U23925 (N_23925,N_22270,N_22790);
or U23926 (N_23926,N_22627,N_22637);
xor U23927 (N_23927,N_22100,N_22417);
or U23928 (N_23928,N_22010,N_22151);
or U23929 (N_23929,N_22473,N_22559);
or U23930 (N_23930,N_22951,N_22757);
or U23931 (N_23931,N_22389,N_22853);
nand U23932 (N_23932,N_22938,N_22391);
or U23933 (N_23933,N_22507,N_22578);
and U23934 (N_23934,N_22797,N_22083);
or U23935 (N_23935,N_22306,N_22063);
nand U23936 (N_23936,N_22444,N_22334);
or U23937 (N_23937,N_22713,N_22087);
nand U23938 (N_23938,N_22013,N_22216);
xor U23939 (N_23939,N_22299,N_22424);
or U23940 (N_23940,N_22783,N_22789);
nand U23941 (N_23941,N_22705,N_22749);
nor U23942 (N_23942,N_22250,N_22401);
or U23943 (N_23943,N_22969,N_22746);
or U23944 (N_23944,N_22041,N_22667);
or U23945 (N_23945,N_22776,N_22689);
and U23946 (N_23946,N_22977,N_22430);
or U23947 (N_23947,N_22511,N_22264);
nand U23948 (N_23948,N_22477,N_22522);
or U23949 (N_23949,N_22861,N_22091);
nor U23950 (N_23950,N_22372,N_22295);
or U23951 (N_23951,N_22079,N_22457);
and U23952 (N_23952,N_22959,N_22312);
or U23953 (N_23953,N_22206,N_22178);
or U23954 (N_23954,N_22032,N_22735);
or U23955 (N_23955,N_22532,N_22032);
or U23956 (N_23956,N_22357,N_22101);
and U23957 (N_23957,N_22197,N_22121);
nor U23958 (N_23958,N_22885,N_22917);
xnor U23959 (N_23959,N_22186,N_22109);
nand U23960 (N_23960,N_22933,N_22839);
nor U23961 (N_23961,N_22083,N_22278);
or U23962 (N_23962,N_22098,N_22305);
xnor U23963 (N_23963,N_22767,N_22463);
xnor U23964 (N_23964,N_22176,N_22064);
nand U23965 (N_23965,N_22568,N_22913);
or U23966 (N_23966,N_22794,N_22650);
nor U23967 (N_23967,N_22838,N_22983);
nand U23968 (N_23968,N_22969,N_22469);
or U23969 (N_23969,N_22471,N_22007);
nand U23970 (N_23970,N_22005,N_22965);
xnor U23971 (N_23971,N_22876,N_22517);
and U23972 (N_23972,N_22939,N_22443);
and U23973 (N_23973,N_22450,N_22161);
nor U23974 (N_23974,N_22175,N_22500);
nor U23975 (N_23975,N_22420,N_22788);
and U23976 (N_23976,N_22686,N_22596);
and U23977 (N_23977,N_22009,N_22452);
or U23978 (N_23978,N_22583,N_22704);
nor U23979 (N_23979,N_22114,N_22850);
or U23980 (N_23980,N_22648,N_22452);
xor U23981 (N_23981,N_22420,N_22587);
or U23982 (N_23982,N_22257,N_22976);
nand U23983 (N_23983,N_22062,N_22338);
nand U23984 (N_23984,N_22385,N_22786);
nor U23985 (N_23985,N_22190,N_22824);
nor U23986 (N_23986,N_22560,N_22854);
nand U23987 (N_23987,N_22302,N_22044);
nand U23988 (N_23988,N_22682,N_22456);
and U23989 (N_23989,N_22094,N_22245);
nor U23990 (N_23990,N_22695,N_22894);
and U23991 (N_23991,N_22066,N_22693);
nand U23992 (N_23992,N_22376,N_22899);
nand U23993 (N_23993,N_22010,N_22063);
or U23994 (N_23994,N_22081,N_22110);
xnor U23995 (N_23995,N_22482,N_22803);
or U23996 (N_23996,N_22930,N_22320);
nand U23997 (N_23997,N_22411,N_22580);
nor U23998 (N_23998,N_22481,N_22306);
nor U23999 (N_23999,N_22641,N_22004);
xnor U24000 (N_24000,N_23536,N_23833);
xnor U24001 (N_24001,N_23651,N_23842);
xnor U24002 (N_24002,N_23747,N_23425);
or U24003 (N_24003,N_23931,N_23848);
nor U24004 (N_24004,N_23904,N_23976);
nand U24005 (N_24005,N_23789,N_23790);
xnor U24006 (N_24006,N_23450,N_23600);
or U24007 (N_24007,N_23427,N_23123);
nor U24008 (N_24008,N_23712,N_23434);
and U24009 (N_24009,N_23535,N_23922);
nand U24010 (N_24010,N_23203,N_23834);
nand U24011 (N_24011,N_23346,N_23301);
or U24012 (N_24012,N_23460,N_23540);
xnor U24013 (N_24013,N_23787,N_23571);
or U24014 (N_24014,N_23523,N_23576);
nand U24015 (N_24015,N_23205,N_23312);
nand U24016 (N_24016,N_23101,N_23290);
or U24017 (N_24017,N_23366,N_23652);
xnor U24018 (N_24018,N_23007,N_23257);
and U24019 (N_24019,N_23231,N_23826);
nand U24020 (N_24020,N_23748,N_23449);
or U24021 (N_24021,N_23376,N_23024);
and U24022 (N_24022,N_23067,N_23823);
nor U24023 (N_24023,N_23059,N_23248);
nor U24024 (N_24024,N_23733,N_23810);
or U24025 (N_24025,N_23817,N_23136);
nand U24026 (N_24026,N_23813,N_23282);
nand U24027 (N_24027,N_23031,N_23738);
or U24028 (N_24028,N_23554,N_23721);
and U24029 (N_24029,N_23951,N_23035);
xnor U24030 (N_24030,N_23029,N_23681);
xnor U24031 (N_24031,N_23084,N_23529);
and U24032 (N_24032,N_23377,N_23378);
and U24033 (N_24033,N_23947,N_23300);
nand U24034 (N_24034,N_23279,N_23461);
nand U24035 (N_24035,N_23433,N_23843);
or U24036 (N_24036,N_23133,N_23187);
nand U24037 (N_24037,N_23556,N_23723);
or U24038 (N_24038,N_23821,N_23752);
and U24039 (N_24039,N_23184,N_23422);
nand U24040 (N_24040,N_23125,N_23226);
nor U24041 (N_24041,N_23470,N_23354);
nand U24042 (N_24042,N_23982,N_23224);
nor U24043 (N_24043,N_23400,N_23132);
nor U24044 (N_24044,N_23838,N_23581);
or U24045 (N_24045,N_23418,N_23528);
and U24046 (N_24046,N_23241,N_23961);
nand U24047 (N_24047,N_23754,N_23941);
or U24048 (N_24048,N_23739,N_23795);
xnor U24049 (N_24049,N_23771,N_23977);
or U24050 (N_24050,N_23166,N_23619);
xnor U24051 (N_24051,N_23895,N_23153);
nand U24052 (N_24052,N_23611,N_23917);
xnor U24053 (N_24053,N_23714,N_23592);
xor U24054 (N_24054,N_23113,N_23948);
nand U24055 (N_24055,N_23837,N_23785);
nor U24056 (N_24056,N_23486,N_23524);
or U24057 (N_24057,N_23437,N_23359);
or U24058 (N_24058,N_23962,N_23860);
xor U24059 (N_24059,N_23511,N_23987);
nand U24060 (N_24060,N_23866,N_23896);
or U24061 (N_24061,N_23942,N_23381);
or U24062 (N_24062,N_23273,N_23678);
or U24063 (N_24063,N_23902,N_23385);
nand U24064 (N_24064,N_23401,N_23316);
and U24065 (N_24065,N_23189,N_23872);
xnor U24066 (N_24066,N_23626,N_23575);
or U24067 (N_24067,N_23713,N_23799);
nand U24068 (N_24068,N_23637,N_23076);
nand U24069 (N_24069,N_23516,N_23918);
and U24070 (N_24070,N_23394,N_23676);
nor U24071 (N_24071,N_23371,N_23983);
or U24072 (N_24072,N_23036,N_23933);
nor U24073 (N_24073,N_23151,N_23130);
nor U24074 (N_24074,N_23037,N_23436);
xnor U24075 (N_24075,N_23538,N_23882);
or U24076 (N_24076,N_23938,N_23343);
nand U24077 (N_24077,N_23202,N_23768);
xnor U24078 (N_24078,N_23491,N_23507);
nor U24079 (N_24079,N_23155,N_23469);
or U24080 (N_24080,N_23050,N_23215);
or U24081 (N_24081,N_23986,N_23596);
xnor U24082 (N_24082,N_23278,N_23981);
nor U24083 (N_24083,N_23158,N_23077);
xor U24084 (N_24084,N_23495,N_23275);
or U24085 (N_24085,N_23318,N_23426);
and U24086 (N_24086,N_23665,N_23533);
xnor U24087 (N_24087,N_23479,N_23310);
nand U24088 (N_24088,N_23672,N_23539);
xnor U24089 (N_24089,N_23852,N_23169);
nor U24090 (N_24090,N_23906,N_23749);
and U24091 (N_24091,N_23091,N_23143);
xnor U24092 (N_24092,N_23692,N_23492);
xnor U24093 (N_24093,N_23392,N_23573);
nor U24094 (N_24094,N_23658,N_23361);
nand U24095 (N_24095,N_23116,N_23435);
nor U24096 (N_24096,N_23660,N_23574);
nand U24097 (N_24097,N_23766,N_23175);
nor U24098 (N_24098,N_23518,N_23191);
nor U24099 (N_24099,N_23625,N_23264);
and U24100 (N_24100,N_23876,N_23193);
or U24101 (N_24101,N_23796,N_23409);
and U24102 (N_24102,N_23375,N_23402);
xnor U24103 (N_24103,N_23332,N_23729);
nor U24104 (N_24104,N_23763,N_23062);
and U24105 (N_24105,N_23246,N_23788);
or U24106 (N_24106,N_23056,N_23499);
xnor U24107 (N_24107,N_23086,N_23643);
nor U24108 (N_24108,N_23755,N_23949);
nor U24109 (N_24109,N_23281,N_23373);
nor U24110 (N_24110,N_23496,N_23840);
and U24111 (N_24111,N_23502,N_23558);
and U24112 (N_24112,N_23888,N_23635);
and U24113 (N_24113,N_23334,N_23302);
nand U24114 (N_24114,N_23033,N_23365);
nor U24115 (N_24115,N_23707,N_23487);
and U24116 (N_24116,N_23548,N_23867);
or U24117 (N_24117,N_23068,N_23628);
or U24118 (N_24118,N_23288,N_23182);
or U24119 (N_24119,N_23965,N_23432);
and U24120 (N_24120,N_23034,N_23777);
and U24121 (N_24121,N_23363,N_23659);
nor U24122 (N_24122,N_23464,N_23701);
and U24123 (N_24123,N_23657,N_23251);
xor U24124 (N_24124,N_23724,N_23131);
nand U24125 (N_24125,N_23975,N_23892);
xnor U24126 (N_24126,N_23974,N_23229);
and U24127 (N_24127,N_23268,N_23283);
or U24128 (N_24128,N_23504,N_23720);
xor U24129 (N_24129,N_23806,N_23990);
or U24130 (N_24130,N_23579,N_23075);
xnor U24131 (N_24131,N_23805,N_23853);
xnor U24132 (N_24132,N_23772,N_23862);
xnor U24133 (N_24133,N_23884,N_23715);
nor U24134 (N_24134,N_23519,N_23515);
and U24135 (N_24135,N_23471,N_23505);
xnor U24136 (N_24136,N_23526,N_23463);
nand U24137 (N_24137,N_23773,N_23988);
nand U24138 (N_24138,N_23330,N_23686);
xor U24139 (N_24139,N_23956,N_23991);
xnor U24140 (N_24140,N_23280,N_23815);
nor U24141 (N_24141,N_23362,N_23909);
and U24142 (N_24142,N_23655,N_23380);
nand U24143 (N_24143,N_23177,N_23305);
and U24144 (N_24144,N_23306,N_23412);
nand U24145 (N_24145,N_23157,N_23198);
nand U24146 (N_24146,N_23924,N_23117);
and U24147 (N_24147,N_23857,N_23874);
and U24148 (N_24148,N_23820,N_23667);
or U24149 (N_24149,N_23928,N_23040);
or U24150 (N_24150,N_23683,N_23816);
nor U24151 (N_24151,N_23172,N_23083);
or U24152 (N_24152,N_23159,N_23213);
nand U24153 (N_24153,N_23134,N_23616);
nor U24154 (N_24154,N_23446,N_23939);
xor U24155 (N_24155,N_23295,N_23138);
or U24156 (N_24156,N_23465,N_23360);
nand U24157 (N_24157,N_23064,N_23026);
nand U24158 (N_24158,N_23480,N_23908);
or U24159 (N_24159,N_23483,N_23049);
nand U24160 (N_24160,N_23699,N_23258);
nor U24161 (N_24161,N_23110,N_23398);
and U24162 (N_24162,N_23836,N_23052);
nand U24163 (N_24163,N_23054,N_23079);
xnor U24164 (N_24164,N_23121,N_23237);
or U24165 (N_24165,N_23244,N_23845);
nor U24166 (N_24166,N_23889,N_23081);
xor U24167 (N_24167,N_23970,N_23442);
or U24168 (N_24168,N_23038,N_23139);
or U24169 (N_24169,N_23679,N_23913);
nor U24170 (N_24170,N_23124,N_23071);
and U24171 (N_24171,N_23717,N_23630);
or U24172 (N_24172,N_23980,N_23569);
xnor U24173 (N_24173,N_23580,N_23760);
nor U24174 (N_24174,N_23314,N_23127);
xor U24175 (N_24175,N_23522,N_23710);
nand U24176 (N_24176,N_23186,N_23243);
nor U24177 (N_24177,N_23448,N_23666);
nand U24178 (N_24178,N_23291,N_23870);
or U24179 (N_24179,N_23217,N_23620);
or U24180 (N_24180,N_23277,N_23741);
nor U24181 (N_24181,N_23794,N_23122);
nor U24182 (N_24182,N_23093,N_23145);
nand U24183 (N_24183,N_23180,N_23832);
nor U24184 (N_24184,N_23368,N_23053);
or U24185 (N_24185,N_23232,N_23353);
xor U24186 (N_24186,N_23689,N_23430);
and U24187 (N_24187,N_23957,N_23473);
nor U24188 (N_24188,N_23897,N_23905);
nor U24189 (N_24189,N_23379,N_23930);
nand U24190 (N_24190,N_23051,N_23100);
nand U24191 (N_24191,N_23259,N_23791);
nand U24192 (N_24192,N_23682,N_23188);
and U24193 (N_24193,N_23728,N_23043);
xor U24194 (N_24194,N_23570,N_23800);
nor U24195 (N_24195,N_23252,N_23058);
nand U24196 (N_24196,N_23673,N_23255);
and U24197 (N_24197,N_23099,N_23021);
and U24198 (N_24198,N_23160,N_23750);
xor U24199 (N_24199,N_23530,N_23740);
xnor U24200 (N_24200,N_23684,N_23289);
xor U24201 (N_24201,N_23105,N_23644);
and U24202 (N_24202,N_23944,N_23937);
nand U24203 (N_24203,N_23731,N_23200);
nand U24204 (N_24204,N_23339,N_23841);
xnor U24205 (N_24205,N_23964,N_23674);
or U24206 (N_24206,N_23225,N_23612);
nor U24207 (N_24207,N_23835,N_23214);
nor U24208 (N_24208,N_23410,N_23112);
nor U24209 (N_24209,N_23615,N_23025);
nor U24210 (N_24210,N_23146,N_23656);
xor U24211 (N_24211,N_23745,N_23164);
nand U24212 (N_24212,N_23935,N_23703);
nor U24213 (N_24213,N_23584,N_23256);
nor U24214 (N_24214,N_23421,N_23424);
or U24215 (N_24215,N_23253,N_23156);
and U24216 (N_24216,N_23591,N_23195);
xnor U24217 (N_24217,N_23585,N_23456);
nand U24218 (N_24218,N_23716,N_23690);
and U24219 (N_24219,N_23671,N_23565);
nor U24220 (N_24220,N_23774,N_23769);
or U24221 (N_24221,N_23984,N_23779);
nor U24222 (N_24222,N_23120,N_23639);
nand U24223 (N_24223,N_23736,N_23002);
nand U24224 (N_24224,N_23793,N_23563);
nor U24225 (N_24225,N_23221,N_23708);
nor U24226 (N_24226,N_23893,N_23072);
nand U24227 (N_24227,N_23209,N_23685);
or U24228 (N_24228,N_23618,N_23627);
or U24229 (N_24229,N_23631,N_23452);
and U24230 (N_24230,N_23017,N_23654);
nor U24231 (N_24231,N_23307,N_23313);
xnor U24232 (N_24232,N_23770,N_23525);
xor U24233 (N_24233,N_23780,N_23814);
xor U24234 (N_24234,N_23020,N_23445);
and U24235 (N_24235,N_23397,N_23910);
or U24236 (N_24236,N_23331,N_23923);
or U24237 (N_24237,N_23521,N_23677);
xnor U24238 (N_24238,N_23952,N_23783);
nor U24239 (N_24239,N_23722,N_23107);
nor U24240 (N_24240,N_23531,N_23932);
or U24241 (N_24241,N_23080,N_23044);
nor U24242 (N_24242,N_23967,N_23664);
xor U24243 (N_24243,N_23199,N_23621);
nor U24244 (N_24244,N_23216,N_23073);
nand U24245 (N_24245,N_23998,N_23792);
nand U24246 (N_24246,N_23008,N_23096);
nor U24247 (N_24247,N_23403,N_23147);
xor U24248 (N_24248,N_23871,N_23687);
nor U24249 (N_24249,N_23012,N_23019);
and U24250 (N_24250,N_23417,N_23388);
and U24251 (N_24251,N_23856,N_23711);
and U24252 (N_24252,N_23901,N_23284);
or U24253 (N_24253,N_23594,N_23734);
nor U24254 (N_24254,N_23048,N_23326);
nand U24255 (N_24255,N_23233,N_23605);
or U24256 (N_24256,N_23358,N_23894);
or U24257 (N_24257,N_23624,N_23118);
or U24258 (N_24258,N_23276,N_23744);
nor U24259 (N_24259,N_23144,N_23577);
or U24260 (N_24260,N_23955,N_23765);
or U24261 (N_24261,N_23509,N_23597);
xnor U24262 (N_24262,N_23356,N_23490);
and U24263 (N_24263,N_23439,N_23335);
nor U24264 (N_24264,N_23802,N_23775);
nand U24265 (N_24265,N_23472,N_23608);
nand U24266 (N_24266,N_23061,N_23041);
or U24267 (N_24267,N_23527,N_23174);
xor U24268 (N_24268,N_23484,N_23467);
nand U24269 (N_24269,N_23270,N_23219);
nand U24270 (N_24270,N_23545,N_23693);
nand U24271 (N_24271,N_23803,N_23859);
or U24272 (N_24272,N_23494,N_23688);
and U24273 (N_24273,N_23032,N_23269);
and U24274 (N_24274,N_23730,N_23055);
xor U24275 (N_24275,N_23443,N_23329);
xnor U24276 (N_24276,N_23582,N_23344);
nor U24277 (N_24277,N_23593,N_23396);
nor U24278 (N_24278,N_23613,N_23261);
nand U24279 (N_24279,N_23801,N_23886);
or U24280 (N_24280,N_23778,N_23285);
nor U24281 (N_24281,N_23969,N_23603);
or U24282 (N_24282,N_23348,N_23271);
nand U24283 (N_24283,N_23920,N_23082);
nor U24284 (N_24284,N_23929,N_23323);
xnor U24285 (N_24285,N_23165,N_23304);
xnor U24286 (N_24286,N_23898,N_23868);
and U24287 (N_24287,N_23847,N_23098);
nand U24288 (N_24288,N_23459,N_23634);
or U24289 (N_24289,N_23234,N_23351);
nor U24290 (N_24290,N_23680,N_23042);
or U24291 (N_24291,N_23812,N_23382);
xor U24292 (N_24292,N_23726,N_23431);
xnor U24293 (N_24293,N_23764,N_23649);
or U24294 (N_24294,N_23719,N_23781);
nand U24295 (N_24295,N_23230,N_23784);
nand U24296 (N_24296,N_23732,N_23762);
and U24297 (N_24297,N_23236,N_23455);
xnor U24298 (N_24298,N_23477,N_23089);
nor U24299 (N_24299,N_23196,N_23709);
or U24300 (N_24300,N_23485,N_23534);
nand U24301 (N_24301,N_23458,N_23429);
xnor U24302 (N_24302,N_23364,N_23263);
nand U24303 (N_24303,N_23336,N_23950);
nor U24304 (N_24304,N_23891,N_23212);
and U24305 (N_24305,N_23228,N_23474);
or U24306 (N_24306,N_23617,N_23451);
nor U24307 (N_24307,N_23702,N_23475);
nor U24308 (N_24308,N_23757,N_23863);
nand U24309 (N_24309,N_23065,N_23009);
nor U24310 (N_24310,N_23150,N_23357);
or U24311 (N_24311,N_23190,N_23598);
xor U24312 (N_24312,N_23415,N_23846);
and U24313 (N_24313,N_23537,N_23869);
xor U24314 (N_24314,N_23387,N_23405);
or U24315 (N_24315,N_23109,N_23006);
or U24316 (N_24316,N_23245,N_23014);
or U24317 (N_24317,N_23997,N_23296);
or U24318 (N_24318,N_23811,N_23010);
and U24319 (N_24319,N_23183,N_23171);
and U24320 (N_24320,N_23807,N_23958);
nor U24321 (N_24321,N_23129,N_23108);
or U24322 (N_24322,N_23883,N_23004);
or U24323 (N_24323,N_23670,N_23207);
nand U24324 (N_24324,N_23865,N_23423);
or U24325 (N_24325,N_23066,N_23406);
and U24326 (N_24326,N_23561,N_23994);
xnor U24327 (N_24327,N_23238,N_23759);
nor U24328 (N_24328,N_23877,N_23168);
and U24329 (N_24329,N_23650,N_23566);
and U24330 (N_24330,N_23743,N_23555);
nand U24331 (N_24331,N_23367,N_23963);
xnor U24332 (N_24332,N_23640,N_23727);
and U24333 (N_24333,N_23444,N_23322);
xor U24334 (N_24334,N_23642,N_23559);
or U24335 (N_24335,N_23602,N_23549);
nand U24336 (N_24336,N_23900,N_23500);
or U24337 (N_24337,N_23979,N_23510);
nor U24338 (N_24338,N_23972,N_23399);
nand U24339 (N_24339,N_23532,N_23114);
nand U24340 (N_24340,N_23247,N_23493);
nor U24341 (N_24341,N_23309,N_23804);
xor U24342 (N_24342,N_23185,N_23718);
and U24343 (N_24343,N_23973,N_23355);
or U24344 (N_24344,N_23704,N_23641);
and U24345 (N_24345,N_23992,N_23223);
nand U24346 (N_24346,N_23604,N_23645);
nand U24347 (N_24347,N_23552,N_23440);
xor U24348 (N_24348,N_23315,N_23022);
xnor U24349 (N_24349,N_23696,N_23661);
and U24350 (N_24350,N_23560,N_23317);
nor U24351 (N_24351,N_23320,N_23911);
nand U24352 (N_24352,N_23137,N_23758);
nor U24353 (N_24353,N_23646,N_23861);
xnor U24354 (N_24354,N_23636,N_23384);
nor U24355 (N_24355,N_23520,N_23737);
nor U24356 (N_24356,N_23498,N_23782);
or U24357 (N_24357,N_23797,N_23849);
or U24358 (N_24358,N_23553,N_23338);
nand U24359 (N_24359,N_23013,N_23167);
xor U24360 (N_24360,N_23586,N_23926);
or U24361 (N_24361,N_23106,N_23063);
nand U24362 (N_24362,N_23092,N_23030);
or U24363 (N_24363,N_23342,N_23181);
nand U24364 (N_24364,N_23419,N_23001);
or U24365 (N_24365,N_23003,N_23027);
nand U24366 (N_24366,N_23220,N_23943);
xnor U24367 (N_24367,N_23925,N_23550);
or U24368 (N_24368,N_23208,N_23919);
or U24369 (N_24369,N_23851,N_23327);
nand U24370 (N_24370,N_23016,N_23135);
nor U24371 (N_24371,N_23267,N_23966);
or U24372 (N_24372,N_23936,N_23163);
and U24373 (N_24373,N_23391,N_23887);
nor U24374 (N_24374,N_23457,N_23023);
xor U24375 (N_24375,N_23864,N_23927);
nor U24376 (N_24376,N_23000,N_23292);
nor U24377 (N_24377,N_23822,N_23201);
or U24378 (N_24378,N_23568,N_23878);
and U24379 (N_24379,N_23638,N_23324);
nand U24380 (N_24380,N_23506,N_23249);
nor U24381 (N_24381,N_23503,N_23829);
xnor U24382 (N_24382,N_23162,N_23178);
or U24383 (N_24383,N_23087,N_23149);
and U24384 (N_24384,N_23194,N_23395);
nor U24385 (N_24385,N_23880,N_23078);
nor U24386 (N_24386,N_23045,N_23543);
or U24387 (N_24387,N_23648,N_23697);
and U24388 (N_24388,N_23633,N_23416);
or U24389 (N_24389,N_23668,N_23468);
nor U24390 (N_24390,N_23954,N_23173);
xor U24391 (N_24391,N_23321,N_23154);
and U24392 (N_24392,N_23272,N_23614);
nand U24393 (N_24393,N_23546,N_23308);
nor U24394 (N_24394,N_23945,N_23753);
or U24395 (N_24395,N_23047,N_23476);
and U24396 (N_24396,N_23197,N_23809);
xnor U24397 (N_24397,N_23547,N_23915);
xor U24398 (N_24398,N_23319,N_23294);
nor U24399 (N_24399,N_23140,N_23890);
xor U24400 (N_24400,N_23386,N_23227);
and U24401 (N_24401,N_23240,N_23907);
nor U24402 (N_24402,N_23239,N_23501);
nor U24403 (N_24403,N_23662,N_23383);
or U24404 (N_24404,N_23695,N_23767);
nand U24405 (N_24405,N_23374,N_23632);
nand U24406 (N_24406,N_23069,N_23609);
nor U24407 (N_24407,N_23148,N_23462);
nor U24408 (N_24408,N_23345,N_23333);
xor U24409 (N_24409,N_23818,N_23606);
or U24410 (N_24410,N_23705,N_23428);
nor U24411 (N_24411,N_23588,N_23875);
or U24412 (N_24412,N_23015,N_23254);
and U24413 (N_24413,N_23946,N_23912);
and U24414 (N_24414,N_23497,N_23482);
and U24415 (N_24415,N_23018,N_23512);
nand U24416 (N_24416,N_23960,N_23706);
xnor U24417 (N_24417,N_23453,N_23663);
or U24418 (N_24418,N_23204,N_23297);
and U24419 (N_24419,N_23206,N_23095);
and U24420 (N_24420,N_23337,N_23347);
or U24421 (N_24421,N_23057,N_23831);
nand U24422 (N_24422,N_23746,N_23250);
or U24423 (N_24423,N_23088,N_23070);
nand U24424 (N_24424,N_23141,N_23060);
and U24425 (N_24425,N_23447,N_23265);
or U24426 (N_24426,N_23102,N_23590);
nor U24427 (N_24427,N_23372,N_23589);
nand U24428 (N_24428,N_23039,N_23786);
and U24429 (N_24429,N_23104,N_23179);
or U24430 (N_24430,N_23959,N_23293);
xnor U24431 (N_24431,N_23481,N_23404);
xnor U24432 (N_24432,N_23514,N_23567);
xnor U24433 (N_24433,N_23756,N_23735);
xor U24434 (N_24434,N_23466,N_23587);
and U24435 (N_24435,N_23694,N_23260);
xnor U24436 (N_24436,N_23873,N_23274);
nand U24437 (N_24437,N_23855,N_23578);
nor U24438 (N_24438,N_23517,N_23218);
and U24439 (N_24439,N_23210,N_23622);
nor U24440 (N_24440,N_23629,N_23170);
or U24441 (N_24441,N_23222,N_23299);
nor U24442 (N_24442,N_23341,N_23085);
and U24443 (N_24443,N_23325,N_23542);
xor U24444 (N_24444,N_23389,N_23830);
nor U24445 (N_24445,N_23700,N_23407);
nor U24446 (N_24446,N_23489,N_23819);
nand U24447 (N_24447,N_23557,N_23242);
nand U24448 (N_24448,N_23126,N_23414);
xor U24449 (N_24449,N_23393,N_23827);
xnor U24450 (N_24450,N_23311,N_23090);
nor U24451 (N_24451,N_23097,N_23508);
or U24452 (N_24452,N_23903,N_23751);
nand U24453 (N_24453,N_23562,N_23369);
nor U24454 (N_24454,N_23303,N_23441);
or U24455 (N_24455,N_23572,N_23599);
nand U24456 (N_24456,N_23776,N_23370);
or U24457 (N_24457,N_23742,N_23940);
xor U24458 (N_24458,N_23328,N_23691);
and U24459 (N_24459,N_23028,N_23235);
and U24460 (N_24460,N_23899,N_23824);
and U24461 (N_24461,N_23858,N_23287);
nand U24462 (N_24462,N_23879,N_23881);
nand U24463 (N_24463,N_23211,N_23996);
nand U24464 (N_24464,N_23349,N_23390);
xnor U24465 (N_24465,N_23011,N_23103);
xor U24466 (N_24466,N_23005,N_23286);
xor U24467 (N_24467,N_23916,N_23607);
nand U24468 (N_24468,N_23340,N_23623);
and U24469 (N_24469,N_23454,N_23989);
xor U24470 (N_24470,N_23595,N_23698);
xor U24471 (N_24471,N_23142,N_23262);
nor U24472 (N_24472,N_23413,N_23583);
xnor U24473 (N_24473,N_23854,N_23046);
or U24474 (N_24474,N_23978,N_23094);
nand U24475 (N_24475,N_23993,N_23921);
nand U24476 (N_24476,N_23828,N_23914);
and U24477 (N_24477,N_23411,N_23352);
nor U24478 (N_24478,N_23298,N_23808);
nor U24479 (N_24479,N_23478,N_23408);
xnor U24480 (N_24480,N_23885,N_23761);
xnor U24481 (N_24481,N_23610,N_23839);
nand U24482 (N_24482,N_23192,N_23115);
and U24483 (N_24483,N_23420,N_23968);
nand U24484 (N_24484,N_23551,N_23176);
nand U24485 (N_24485,N_23488,N_23669);
nor U24486 (N_24486,N_23161,N_23119);
or U24487 (N_24487,N_23971,N_23074);
nand U24488 (N_24488,N_23999,N_23350);
and U24489 (N_24489,N_23152,N_23541);
and U24490 (N_24490,N_23128,N_23844);
nor U24491 (N_24491,N_23953,N_23647);
xor U24492 (N_24492,N_23111,N_23798);
and U24493 (N_24493,N_23653,N_23995);
or U24494 (N_24494,N_23675,N_23513);
and U24495 (N_24495,N_23725,N_23266);
nand U24496 (N_24496,N_23825,N_23934);
nor U24497 (N_24497,N_23544,N_23601);
nand U24498 (N_24498,N_23438,N_23985);
xnor U24499 (N_24499,N_23850,N_23564);
or U24500 (N_24500,N_23321,N_23002);
or U24501 (N_24501,N_23455,N_23963);
and U24502 (N_24502,N_23044,N_23027);
nand U24503 (N_24503,N_23102,N_23761);
and U24504 (N_24504,N_23025,N_23555);
nor U24505 (N_24505,N_23313,N_23408);
nand U24506 (N_24506,N_23007,N_23265);
xor U24507 (N_24507,N_23332,N_23696);
or U24508 (N_24508,N_23899,N_23700);
nand U24509 (N_24509,N_23836,N_23458);
xnor U24510 (N_24510,N_23440,N_23150);
and U24511 (N_24511,N_23508,N_23046);
nand U24512 (N_24512,N_23484,N_23088);
nand U24513 (N_24513,N_23258,N_23904);
or U24514 (N_24514,N_23972,N_23842);
nor U24515 (N_24515,N_23822,N_23350);
xnor U24516 (N_24516,N_23543,N_23696);
nor U24517 (N_24517,N_23945,N_23031);
and U24518 (N_24518,N_23306,N_23216);
and U24519 (N_24519,N_23425,N_23945);
nand U24520 (N_24520,N_23114,N_23298);
nor U24521 (N_24521,N_23076,N_23523);
and U24522 (N_24522,N_23235,N_23054);
xnor U24523 (N_24523,N_23064,N_23629);
nor U24524 (N_24524,N_23544,N_23504);
nand U24525 (N_24525,N_23877,N_23404);
xnor U24526 (N_24526,N_23350,N_23272);
nand U24527 (N_24527,N_23174,N_23178);
and U24528 (N_24528,N_23960,N_23052);
and U24529 (N_24529,N_23063,N_23621);
xnor U24530 (N_24530,N_23771,N_23933);
nor U24531 (N_24531,N_23868,N_23786);
and U24532 (N_24532,N_23869,N_23555);
nor U24533 (N_24533,N_23341,N_23255);
nand U24534 (N_24534,N_23782,N_23631);
nand U24535 (N_24535,N_23007,N_23636);
or U24536 (N_24536,N_23599,N_23253);
xnor U24537 (N_24537,N_23417,N_23999);
nor U24538 (N_24538,N_23961,N_23963);
or U24539 (N_24539,N_23172,N_23407);
and U24540 (N_24540,N_23403,N_23827);
and U24541 (N_24541,N_23924,N_23435);
nand U24542 (N_24542,N_23466,N_23273);
and U24543 (N_24543,N_23284,N_23604);
and U24544 (N_24544,N_23301,N_23203);
nand U24545 (N_24545,N_23724,N_23168);
or U24546 (N_24546,N_23232,N_23452);
nor U24547 (N_24547,N_23600,N_23551);
and U24548 (N_24548,N_23572,N_23047);
and U24549 (N_24549,N_23341,N_23198);
nor U24550 (N_24550,N_23800,N_23904);
and U24551 (N_24551,N_23548,N_23978);
nand U24552 (N_24552,N_23493,N_23080);
nor U24553 (N_24553,N_23753,N_23151);
or U24554 (N_24554,N_23430,N_23490);
xnor U24555 (N_24555,N_23466,N_23435);
xnor U24556 (N_24556,N_23199,N_23422);
xnor U24557 (N_24557,N_23766,N_23892);
xor U24558 (N_24558,N_23988,N_23256);
nor U24559 (N_24559,N_23519,N_23468);
or U24560 (N_24560,N_23493,N_23535);
nor U24561 (N_24561,N_23599,N_23850);
xor U24562 (N_24562,N_23312,N_23578);
nand U24563 (N_24563,N_23630,N_23425);
nand U24564 (N_24564,N_23067,N_23005);
or U24565 (N_24565,N_23376,N_23884);
nand U24566 (N_24566,N_23867,N_23864);
nor U24567 (N_24567,N_23091,N_23406);
nand U24568 (N_24568,N_23547,N_23653);
or U24569 (N_24569,N_23671,N_23258);
or U24570 (N_24570,N_23715,N_23213);
and U24571 (N_24571,N_23334,N_23907);
nand U24572 (N_24572,N_23506,N_23166);
nor U24573 (N_24573,N_23168,N_23213);
and U24574 (N_24574,N_23059,N_23041);
nand U24575 (N_24575,N_23576,N_23137);
nand U24576 (N_24576,N_23678,N_23119);
nand U24577 (N_24577,N_23819,N_23892);
nand U24578 (N_24578,N_23966,N_23133);
nand U24579 (N_24579,N_23728,N_23730);
or U24580 (N_24580,N_23193,N_23329);
nand U24581 (N_24581,N_23575,N_23525);
nor U24582 (N_24582,N_23440,N_23509);
nand U24583 (N_24583,N_23032,N_23722);
or U24584 (N_24584,N_23205,N_23632);
or U24585 (N_24585,N_23414,N_23174);
nor U24586 (N_24586,N_23903,N_23669);
nor U24587 (N_24587,N_23179,N_23332);
xor U24588 (N_24588,N_23369,N_23387);
nand U24589 (N_24589,N_23784,N_23386);
nand U24590 (N_24590,N_23602,N_23360);
xnor U24591 (N_24591,N_23012,N_23366);
nor U24592 (N_24592,N_23743,N_23853);
xnor U24593 (N_24593,N_23853,N_23060);
xnor U24594 (N_24594,N_23740,N_23665);
xnor U24595 (N_24595,N_23096,N_23137);
and U24596 (N_24596,N_23544,N_23262);
nand U24597 (N_24597,N_23248,N_23432);
nand U24598 (N_24598,N_23104,N_23470);
nor U24599 (N_24599,N_23160,N_23197);
nor U24600 (N_24600,N_23083,N_23864);
nor U24601 (N_24601,N_23599,N_23346);
nand U24602 (N_24602,N_23678,N_23577);
xnor U24603 (N_24603,N_23034,N_23002);
nand U24604 (N_24604,N_23435,N_23373);
nand U24605 (N_24605,N_23812,N_23195);
and U24606 (N_24606,N_23350,N_23897);
nand U24607 (N_24607,N_23205,N_23943);
nand U24608 (N_24608,N_23910,N_23446);
nor U24609 (N_24609,N_23148,N_23539);
nor U24610 (N_24610,N_23138,N_23804);
xnor U24611 (N_24611,N_23472,N_23176);
or U24612 (N_24612,N_23111,N_23947);
nand U24613 (N_24613,N_23991,N_23556);
nand U24614 (N_24614,N_23103,N_23541);
nor U24615 (N_24615,N_23643,N_23138);
and U24616 (N_24616,N_23693,N_23946);
or U24617 (N_24617,N_23556,N_23582);
nor U24618 (N_24618,N_23109,N_23018);
or U24619 (N_24619,N_23034,N_23948);
and U24620 (N_24620,N_23850,N_23364);
nand U24621 (N_24621,N_23656,N_23030);
and U24622 (N_24622,N_23436,N_23122);
or U24623 (N_24623,N_23147,N_23714);
nor U24624 (N_24624,N_23276,N_23278);
or U24625 (N_24625,N_23939,N_23653);
or U24626 (N_24626,N_23786,N_23114);
or U24627 (N_24627,N_23268,N_23295);
and U24628 (N_24628,N_23925,N_23759);
xnor U24629 (N_24629,N_23175,N_23802);
nand U24630 (N_24630,N_23618,N_23426);
nand U24631 (N_24631,N_23119,N_23748);
or U24632 (N_24632,N_23382,N_23389);
and U24633 (N_24633,N_23867,N_23569);
nor U24634 (N_24634,N_23367,N_23137);
xor U24635 (N_24635,N_23733,N_23788);
or U24636 (N_24636,N_23650,N_23112);
xor U24637 (N_24637,N_23353,N_23712);
nand U24638 (N_24638,N_23933,N_23475);
or U24639 (N_24639,N_23423,N_23026);
nor U24640 (N_24640,N_23251,N_23707);
and U24641 (N_24641,N_23947,N_23920);
xnor U24642 (N_24642,N_23665,N_23952);
xnor U24643 (N_24643,N_23048,N_23535);
or U24644 (N_24644,N_23447,N_23564);
nand U24645 (N_24645,N_23632,N_23068);
or U24646 (N_24646,N_23363,N_23284);
xnor U24647 (N_24647,N_23274,N_23746);
nand U24648 (N_24648,N_23690,N_23669);
xnor U24649 (N_24649,N_23026,N_23752);
xnor U24650 (N_24650,N_23963,N_23682);
xor U24651 (N_24651,N_23160,N_23215);
or U24652 (N_24652,N_23317,N_23660);
and U24653 (N_24653,N_23333,N_23129);
and U24654 (N_24654,N_23131,N_23443);
xor U24655 (N_24655,N_23921,N_23991);
xnor U24656 (N_24656,N_23892,N_23271);
xnor U24657 (N_24657,N_23607,N_23210);
nor U24658 (N_24658,N_23431,N_23927);
nor U24659 (N_24659,N_23686,N_23948);
nor U24660 (N_24660,N_23875,N_23110);
nor U24661 (N_24661,N_23334,N_23491);
or U24662 (N_24662,N_23992,N_23178);
xnor U24663 (N_24663,N_23726,N_23621);
and U24664 (N_24664,N_23964,N_23478);
or U24665 (N_24665,N_23931,N_23807);
and U24666 (N_24666,N_23379,N_23817);
nor U24667 (N_24667,N_23200,N_23757);
nand U24668 (N_24668,N_23683,N_23140);
and U24669 (N_24669,N_23043,N_23347);
and U24670 (N_24670,N_23412,N_23646);
nand U24671 (N_24671,N_23832,N_23260);
nand U24672 (N_24672,N_23282,N_23657);
or U24673 (N_24673,N_23380,N_23327);
nand U24674 (N_24674,N_23428,N_23666);
and U24675 (N_24675,N_23825,N_23313);
nand U24676 (N_24676,N_23867,N_23287);
nand U24677 (N_24677,N_23507,N_23557);
nor U24678 (N_24678,N_23244,N_23379);
nand U24679 (N_24679,N_23471,N_23141);
nand U24680 (N_24680,N_23204,N_23308);
and U24681 (N_24681,N_23230,N_23634);
or U24682 (N_24682,N_23076,N_23377);
nor U24683 (N_24683,N_23849,N_23814);
xor U24684 (N_24684,N_23457,N_23732);
xnor U24685 (N_24685,N_23540,N_23679);
xnor U24686 (N_24686,N_23321,N_23860);
nor U24687 (N_24687,N_23936,N_23034);
nor U24688 (N_24688,N_23178,N_23117);
xnor U24689 (N_24689,N_23623,N_23332);
and U24690 (N_24690,N_23936,N_23377);
xnor U24691 (N_24691,N_23626,N_23548);
xnor U24692 (N_24692,N_23735,N_23684);
nor U24693 (N_24693,N_23334,N_23775);
and U24694 (N_24694,N_23828,N_23568);
nor U24695 (N_24695,N_23319,N_23602);
xor U24696 (N_24696,N_23206,N_23901);
nand U24697 (N_24697,N_23646,N_23726);
nor U24698 (N_24698,N_23309,N_23191);
or U24699 (N_24699,N_23109,N_23293);
xnor U24700 (N_24700,N_23164,N_23027);
and U24701 (N_24701,N_23225,N_23576);
and U24702 (N_24702,N_23046,N_23295);
nand U24703 (N_24703,N_23281,N_23695);
nand U24704 (N_24704,N_23401,N_23547);
and U24705 (N_24705,N_23382,N_23354);
xnor U24706 (N_24706,N_23448,N_23358);
nand U24707 (N_24707,N_23190,N_23307);
or U24708 (N_24708,N_23474,N_23494);
xnor U24709 (N_24709,N_23343,N_23266);
nor U24710 (N_24710,N_23302,N_23271);
nor U24711 (N_24711,N_23761,N_23849);
nand U24712 (N_24712,N_23049,N_23885);
xnor U24713 (N_24713,N_23273,N_23557);
xnor U24714 (N_24714,N_23506,N_23852);
and U24715 (N_24715,N_23769,N_23349);
xnor U24716 (N_24716,N_23184,N_23147);
or U24717 (N_24717,N_23785,N_23344);
nor U24718 (N_24718,N_23039,N_23872);
nor U24719 (N_24719,N_23460,N_23543);
nand U24720 (N_24720,N_23156,N_23869);
nor U24721 (N_24721,N_23507,N_23593);
and U24722 (N_24722,N_23935,N_23249);
xor U24723 (N_24723,N_23220,N_23981);
nand U24724 (N_24724,N_23133,N_23581);
nor U24725 (N_24725,N_23262,N_23631);
and U24726 (N_24726,N_23760,N_23658);
nor U24727 (N_24727,N_23269,N_23239);
or U24728 (N_24728,N_23708,N_23044);
xor U24729 (N_24729,N_23245,N_23203);
nor U24730 (N_24730,N_23661,N_23832);
nand U24731 (N_24731,N_23923,N_23166);
nand U24732 (N_24732,N_23002,N_23325);
or U24733 (N_24733,N_23518,N_23156);
nand U24734 (N_24734,N_23043,N_23611);
or U24735 (N_24735,N_23944,N_23873);
or U24736 (N_24736,N_23100,N_23005);
xnor U24737 (N_24737,N_23852,N_23328);
nand U24738 (N_24738,N_23530,N_23919);
and U24739 (N_24739,N_23683,N_23907);
xor U24740 (N_24740,N_23517,N_23229);
xor U24741 (N_24741,N_23028,N_23064);
nand U24742 (N_24742,N_23827,N_23160);
nand U24743 (N_24743,N_23203,N_23548);
nor U24744 (N_24744,N_23532,N_23093);
or U24745 (N_24745,N_23751,N_23128);
nand U24746 (N_24746,N_23733,N_23883);
and U24747 (N_24747,N_23638,N_23960);
nand U24748 (N_24748,N_23473,N_23163);
nand U24749 (N_24749,N_23734,N_23884);
and U24750 (N_24750,N_23721,N_23100);
nor U24751 (N_24751,N_23979,N_23581);
nand U24752 (N_24752,N_23103,N_23705);
nand U24753 (N_24753,N_23023,N_23608);
nor U24754 (N_24754,N_23367,N_23016);
xor U24755 (N_24755,N_23014,N_23534);
nor U24756 (N_24756,N_23595,N_23790);
xnor U24757 (N_24757,N_23767,N_23448);
nor U24758 (N_24758,N_23560,N_23336);
and U24759 (N_24759,N_23436,N_23228);
and U24760 (N_24760,N_23422,N_23441);
nand U24761 (N_24761,N_23847,N_23164);
nor U24762 (N_24762,N_23810,N_23957);
nand U24763 (N_24763,N_23491,N_23128);
or U24764 (N_24764,N_23613,N_23272);
xnor U24765 (N_24765,N_23264,N_23578);
nor U24766 (N_24766,N_23759,N_23334);
and U24767 (N_24767,N_23873,N_23562);
and U24768 (N_24768,N_23782,N_23442);
or U24769 (N_24769,N_23989,N_23387);
nor U24770 (N_24770,N_23574,N_23061);
xnor U24771 (N_24771,N_23201,N_23369);
and U24772 (N_24772,N_23862,N_23785);
and U24773 (N_24773,N_23365,N_23088);
and U24774 (N_24774,N_23717,N_23993);
or U24775 (N_24775,N_23851,N_23666);
or U24776 (N_24776,N_23788,N_23896);
or U24777 (N_24777,N_23225,N_23328);
and U24778 (N_24778,N_23410,N_23599);
or U24779 (N_24779,N_23104,N_23958);
nor U24780 (N_24780,N_23660,N_23801);
and U24781 (N_24781,N_23238,N_23435);
and U24782 (N_24782,N_23323,N_23654);
nor U24783 (N_24783,N_23016,N_23930);
nor U24784 (N_24784,N_23070,N_23652);
nand U24785 (N_24785,N_23125,N_23515);
nor U24786 (N_24786,N_23101,N_23298);
nand U24787 (N_24787,N_23102,N_23400);
xor U24788 (N_24788,N_23924,N_23685);
nand U24789 (N_24789,N_23713,N_23137);
xnor U24790 (N_24790,N_23333,N_23580);
and U24791 (N_24791,N_23512,N_23698);
or U24792 (N_24792,N_23796,N_23413);
or U24793 (N_24793,N_23674,N_23746);
nor U24794 (N_24794,N_23066,N_23769);
nand U24795 (N_24795,N_23158,N_23806);
xor U24796 (N_24796,N_23676,N_23389);
and U24797 (N_24797,N_23450,N_23280);
nand U24798 (N_24798,N_23577,N_23161);
and U24799 (N_24799,N_23137,N_23216);
or U24800 (N_24800,N_23387,N_23236);
nand U24801 (N_24801,N_23759,N_23921);
and U24802 (N_24802,N_23568,N_23870);
or U24803 (N_24803,N_23271,N_23588);
xnor U24804 (N_24804,N_23147,N_23103);
nor U24805 (N_24805,N_23495,N_23066);
nand U24806 (N_24806,N_23081,N_23615);
or U24807 (N_24807,N_23654,N_23480);
nor U24808 (N_24808,N_23402,N_23384);
xor U24809 (N_24809,N_23067,N_23965);
or U24810 (N_24810,N_23607,N_23896);
and U24811 (N_24811,N_23687,N_23002);
and U24812 (N_24812,N_23158,N_23595);
or U24813 (N_24813,N_23210,N_23330);
nor U24814 (N_24814,N_23158,N_23476);
nand U24815 (N_24815,N_23482,N_23472);
nand U24816 (N_24816,N_23589,N_23032);
xor U24817 (N_24817,N_23693,N_23810);
xnor U24818 (N_24818,N_23602,N_23884);
or U24819 (N_24819,N_23161,N_23208);
xor U24820 (N_24820,N_23650,N_23519);
xor U24821 (N_24821,N_23445,N_23215);
xor U24822 (N_24822,N_23688,N_23861);
nor U24823 (N_24823,N_23427,N_23568);
and U24824 (N_24824,N_23030,N_23340);
nor U24825 (N_24825,N_23704,N_23409);
nor U24826 (N_24826,N_23700,N_23421);
and U24827 (N_24827,N_23010,N_23150);
nand U24828 (N_24828,N_23429,N_23011);
and U24829 (N_24829,N_23456,N_23829);
nand U24830 (N_24830,N_23490,N_23184);
xor U24831 (N_24831,N_23404,N_23478);
nor U24832 (N_24832,N_23446,N_23743);
or U24833 (N_24833,N_23222,N_23754);
nand U24834 (N_24834,N_23616,N_23988);
xor U24835 (N_24835,N_23058,N_23598);
nand U24836 (N_24836,N_23045,N_23150);
or U24837 (N_24837,N_23186,N_23882);
or U24838 (N_24838,N_23320,N_23879);
and U24839 (N_24839,N_23062,N_23930);
or U24840 (N_24840,N_23486,N_23442);
or U24841 (N_24841,N_23293,N_23019);
or U24842 (N_24842,N_23523,N_23032);
xor U24843 (N_24843,N_23863,N_23455);
nand U24844 (N_24844,N_23809,N_23187);
or U24845 (N_24845,N_23708,N_23302);
or U24846 (N_24846,N_23393,N_23286);
or U24847 (N_24847,N_23530,N_23606);
or U24848 (N_24848,N_23052,N_23049);
and U24849 (N_24849,N_23992,N_23135);
and U24850 (N_24850,N_23394,N_23097);
nor U24851 (N_24851,N_23059,N_23476);
nor U24852 (N_24852,N_23834,N_23625);
nand U24853 (N_24853,N_23196,N_23612);
and U24854 (N_24854,N_23645,N_23018);
nor U24855 (N_24855,N_23447,N_23137);
and U24856 (N_24856,N_23046,N_23612);
xnor U24857 (N_24857,N_23612,N_23255);
nand U24858 (N_24858,N_23650,N_23311);
and U24859 (N_24859,N_23522,N_23821);
nand U24860 (N_24860,N_23704,N_23209);
nand U24861 (N_24861,N_23503,N_23083);
xnor U24862 (N_24862,N_23554,N_23980);
nand U24863 (N_24863,N_23366,N_23018);
nor U24864 (N_24864,N_23428,N_23517);
or U24865 (N_24865,N_23946,N_23599);
xnor U24866 (N_24866,N_23086,N_23760);
or U24867 (N_24867,N_23277,N_23606);
nand U24868 (N_24868,N_23602,N_23241);
and U24869 (N_24869,N_23119,N_23860);
or U24870 (N_24870,N_23777,N_23091);
or U24871 (N_24871,N_23514,N_23480);
nor U24872 (N_24872,N_23315,N_23934);
nor U24873 (N_24873,N_23036,N_23506);
nor U24874 (N_24874,N_23171,N_23425);
xnor U24875 (N_24875,N_23061,N_23939);
or U24876 (N_24876,N_23931,N_23219);
xor U24877 (N_24877,N_23031,N_23413);
xor U24878 (N_24878,N_23969,N_23677);
or U24879 (N_24879,N_23770,N_23559);
or U24880 (N_24880,N_23047,N_23065);
nor U24881 (N_24881,N_23350,N_23866);
or U24882 (N_24882,N_23413,N_23072);
or U24883 (N_24883,N_23706,N_23642);
nand U24884 (N_24884,N_23454,N_23537);
xor U24885 (N_24885,N_23545,N_23304);
nor U24886 (N_24886,N_23374,N_23765);
xnor U24887 (N_24887,N_23018,N_23196);
nand U24888 (N_24888,N_23346,N_23690);
or U24889 (N_24889,N_23054,N_23383);
xnor U24890 (N_24890,N_23827,N_23025);
and U24891 (N_24891,N_23651,N_23309);
or U24892 (N_24892,N_23776,N_23433);
nand U24893 (N_24893,N_23583,N_23696);
and U24894 (N_24894,N_23351,N_23149);
nor U24895 (N_24895,N_23700,N_23687);
or U24896 (N_24896,N_23507,N_23898);
xor U24897 (N_24897,N_23311,N_23391);
xnor U24898 (N_24898,N_23023,N_23115);
and U24899 (N_24899,N_23163,N_23087);
and U24900 (N_24900,N_23238,N_23773);
nor U24901 (N_24901,N_23186,N_23589);
and U24902 (N_24902,N_23653,N_23803);
or U24903 (N_24903,N_23661,N_23922);
and U24904 (N_24904,N_23574,N_23105);
and U24905 (N_24905,N_23431,N_23788);
xnor U24906 (N_24906,N_23011,N_23540);
or U24907 (N_24907,N_23370,N_23899);
nor U24908 (N_24908,N_23249,N_23529);
xnor U24909 (N_24909,N_23430,N_23957);
or U24910 (N_24910,N_23386,N_23234);
or U24911 (N_24911,N_23364,N_23189);
xnor U24912 (N_24912,N_23461,N_23382);
or U24913 (N_24913,N_23847,N_23981);
nor U24914 (N_24914,N_23866,N_23527);
xnor U24915 (N_24915,N_23637,N_23798);
nor U24916 (N_24916,N_23300,N_23149);
xor U24917 (N_24917,N_23149,N_23937);
nand U24918 (N_24918,N_23805,N_23460);
nand U24919 (N_24919,N_23285,N_23784);
or U24920 (N_24920,N_23813,N_23723);
nand U24921 (N_24921,N_23002,N_23199);
and U24922 (N_24922,N_23792,N_23669);
nand U24923 (N_24923,N_23014,N_23083);
nand U24924 (N_24924,N_23379,N_23310);
xnor U24925 (N_24925,N_23007,N_23824);
nor U24926 (N_24926,N_23354,N_23398);
or U24927 (N_24927,N_23184,N_23728);
nor U24928 (N_24928,N_23017,N_23933);
nand U24929 (N_24929,N_23722,N_23304);
or U24930 (N_24930,N_23810,N_23212);
nand U24931 (N_24931,N_23483,N_23244);
nand U24932 (N_24932,N_23600,N_23069);
xnor U24933 (N_24933,N_23996,N_23229);
nor U24934 (N_24934,N_23681,N_23253);
nor U24935 (N_24935,N_23375,N_23267);
xnor U24936 (N_24936,N_23694,N_23760);
xnor U24937 (N_24937,N_23610,N_23636);
and U24938 (N_24938,N_23842,N_23693);
xor U24939 (N_24939,N_23092,N_23790);
nor U24940 (N_24940,N_23217,N_23249);
nand U24941 (N_24941,N_23469,N_23285);
or U24942 (N_24942,N_23633,N_23173);
xor U24943 (N_24943,N_23782,N_23132);
xor U24944 (N_24944,N_23205,N_23088);
nor U24945 (N_24945,N_23762,N_23305);
and U24946 (N_24946,N_23171,N_23348);
and U24947 (N_24947,N_23320,N_23680);
nand U24948 (N_24948,N_23468,N_23034);
nand U24949 (N_24949,N_23205,N_23049);
and U24950 (N_24950,N_23982,N_23704);
or U24951 (N_24951,N_23279,N_23711);
or U24952 (N_24952,N_23109,N_23831);
and U24953 (N_24953,N_23377,N_23842);
xnor U24954 (N_24954,N_23465,N_23906);
or U24955 (N_24955,N_23574,N_23804);
xor U24956 (N_24956,N_23279,N_23401);
and U24957 (N_24957,N_23209,N_23444);
xor U24958 (N_24958,N_23286,N_23159);
and U24959 (N_24959,N_23754,N_23271);
nor U24960 (N_24960,N_23058,N_23172);
or U24961 (N_24961,N_23673,N_23700);
nor U24962 (N_24962,N_23533,N_23154);
xnor U24963 (N_24963,N_23276,N_23382);
and U24964 (N_24964,N_23883,N_23521);
or U24965 (N_24965,N_23427,N_23589);
xor U24966 (N_24966,N_23392,N_23938);
nand U24967 (N_24967,N_23843,N_23081);
and U24968 (N_24968,N_23762,N_23127);
nand U24969 (N_24969,N_23725,N_23061);
and U24970 (N_24970,N_23060,N_23386);
nand U24971 (N_24971,N_23843,N_23122);
nand U24972 (N_24972,N_23264,N_23731);
xnor U24973 (N_24973,N_23713,N_23349);
xnor U24974 (N_24974,N_23591,N_23292);
or U24975 (N_24975,N_23580,N_23500);
or U24976 (N_24976,N_23922,N_23478);
nor U24977 (N_24977,N_23293,N_23925);
nor U24978 (N_24978,N_23605,N_23704);
and U24979 (N_24979,N_23544,N_23720);
nor U24980 (N_24980,N_23995,N_23678);
and U24981 (N_24981,N_23622,N_23004);
nor U24982 (N_24982,N_23029,N_23395);
or U24983 (N_24983,N_23759,N_23605);
and U24984 (N_24984,N_23184,N_23267);
xor U24985 (N_24985,N_23133,N_23329);
and U24986 (N_24986,N_23114,N_23422);
nor U24987 (N_24987,N_23078,N_23524);
or U24988 (N_24988,N_23016,N_23887);
nand U24989 (N_24989,N_23983,N_23780);
and U24990 (N_24990,N_23888,N_23771);
nand U24991 (N_24991,N_23209,N_23158);
and U24992 (N_24992,N_23582,N_23447);
nor U24993 (N_24993,N_23633,N_23884);
and U24994 (N_24994,N_23817,N_23413);
or U24995 (N_24995,N_23925,N_23257);
and U24996 (N_24996,N_23626,N_23419);
xor U24997 (N_24997,N_23169,N_23305);
and U24998 (N_24998,N_23595,N_23952);
xnor U24999 (N_24999,N_23703,N_23207);
or U25000 (N_25000,N_24134,N_24962);
xor U25001 (N_25001,N_24720,N_24291);
nor U25002 (N_25002,N_24673,N_24709);
or U25003 (N_25003,N_24512,N_24542);
nor U25004 (N_25004,N_24901,N_24548);
nand U25005 (N_25005,N_24399,N_24359);
nand U25006 (N_25006,N_24922,N_24212);
xor U25007 (N_25007,N_24747,N_24917);
xor U25008 (N_25008,N_24361,N_24337);
nor U25009 (N_25009,N_24480,N_24386);
and U25010 (N_25010,N_24382,N_24025);
nand U25011 (N_25011,N_24681,N_24330);
and U25012 (N_25012,N_24978,N_24558);
or U25013 (N_25013,N_24357,N_24507);
and U25014 (N_25014,N_24077,N_24501);
and U25015 (N_25015,N_24995,N_24105);
and U25016 (N_25016,N_24260,N_24145);
xor U25017 (N_25017,N_24178,N_24336);
nor U25018 (N_25018,N_24969,N_24071);
or U25019 (N_25019,N_24426,N_24907);
or U25020 (N_25020,N_24109,N_24283);
xnor U25021 (N_25021,N_24365,N_24470);
or U25022 (N_25022,N_24515,N_24717);
nand U25023 (N_25023,N_24831,N_24510);
nor U25024 (N_25024,N_24887,N_24492);
or U25025 (N_25025,N_24862,N_24708);
or U25026 (N_25026,N_24166,N_24618);
or U25027 (N_25027,N_24724,N_24885);
xor U25028 (N_25028,N_24646,N_24697);
xnor U25029 (N_25029,N_24019,N_24443);
xor U25030 (N_25030,N_24861,N_24826);
nor U25031 (N_25031,N_24063,N_24363);
nor U25032 (N_25032,N_24857,N_24240);
or U25033 (N_25033,N_24564,N_24088);
and U25034 (N_25034,N_24214,N_24913);
and U25035 (N_25035,N_24853,N_24349);
or U25036 (N_25036,N_24035,N_24529);
xnor U25037 (N_25037,N_24964,N_24433);
nor U25038 (N_25038,N_24199,N_24074);
nand U25039 (N_25039,N_24723,N_24645);
xor U25040 (N_25040,N_24085,N_24356);
xor U25041 (N_25041,N_24476,N_24555);
or U25042 (N_25042,N_24008,N_24301);
and U25043 (N_25043,N_24094,N_24251);
xor U25044 (N_25044,N_24338,N_24345);
and U25045 (N_25045,N_24486,N_24845);
nand U25046 (N_25046,N_24671,N_24783);
nor U25047 (N_25047,N_24284,N_24554);
nand U25048 (N_25048,N_24712,N_24144);
nor U25049 (N_25049,N_24619,N_24463);
xor U25050 (N_25050,N_24224,N_24967);
and U25051 (N_25051,N_24730,N_24482);
nand U25052 (N_25052,N_24523,N_24597);
and U25053 (N_25053,N_24466,N_24891);
or U25054 (N_25054,N_24531,N_24689);
nand U25055 (N_25055,N_24381,N_24435);
nand U25056 (N_25056,N_24606,N_24687);
nor U25057 (N_25057,N_24763,N_24659);
or U25058 (N_25058,N_24136,N_24150);
and U25059 (N_25059,N_24794,N_24699);
or U25060 (N_25060,N_24582,N_24966);
and U25061 (N_25061,N_24131,N_24350);
nand U25062 (N_25062,N_24308,N_24781);
or U25063 (N_25063,N_24117,N_24755);
and U25064 (N_25064,N_24552,N_24469);
nand U25065 (N_25065,N_24812,N_24406);
xor U25066 (N_25066,N_24255,N_24248);
and U25067 (N_25067,N_24648,N_24431);
nor U25068 (N_25068,N_24825,N_24231);
or U25069 (N_25069,N_24366,N_24209);
xor U25070 (N_25070,N_24402,N_24745);
xor U25071 (N_25071,N_24153,N_24066);
xnor U25072 (N_25072,N_24961,N_24353);
or U25073 (N_25073,N_24772,N_24344);
xor U25074 (N_25074,N_24220,N_24587);
or U25075 (N_25075,N_24654,N_24513);
or U25076 (N_25076,N_24686,N_24398);
nand U25077 (N_25077,N_24737,N_24722);
and U25078 (N_25078,N_24270,N_24418);
or U25079 (N_25079,N_24522,N_24617);
and U25080 (N_25080,N_24777,N_24296);
nor U25081 (N_25081,N_24932,N_24824);
xnor U25082 (N_25082,N_24930,N_24976);
or U25083 (N_25083,N_24154,N_24124);
xor U25084 (N_25084,N_24293,N_24414);
or U25085 (N_25085,N_24233,N_24559);
nand U25086 (N_25086,N_24385,N_24565);
nand U25087 (N_25087,N_24729,N_24459);
nand U25088 (N_25088,N_24351,N_24180);
nor U25089 (N_25089,N_24493,N_24550);
nand U25090 (N_25090,N_24206,N_24354);
or U25091 (N_25091,N_24685,N_24910);
or U25092 (N_25092,N_24079,N_24888);
or U25093 (N_25093,N_24388,N_24241);
nor U25094 (N_25094,N_24836,N_24900);
or U25095 (N_25095,N_24649,N_24412);
or U25096 (N_25096,N_24946,N_24848);
nor U25097 (N_25097,N_24537,N_24702);
nand U25098 (N_25098,N_24111,N_24926);
and U25099 (N_25099,N_24101,N_24139);
or U25100 (N_25100,N_24860,N_24416);
xor U25101 (N_25101,N_24315,N_24496);
xnor U25102 (N_25102,N_24477,N_24525);
and U25103 (N_25103,N_24249,N_24440);
xor U25104 (N_25104,N_24949,N_24622);
nor U25105 (N_25105,N_24464,N_24731);
and U25106 (N_25106,N_24140,N_24918);
or U25107 (N_25107,N_24786,N_24122);
nor U25108 (N_25108,N_24034,N_24504);
and U25109 (N_25109,N_24458,N_24688);
or U25110 (N_25110,N_24302,N_24149);
and U25111 (N_25111,N_24563,N_24938);
and U25112 (N_25112,N_24757,N_24256);
or U25113 (N_25113,N_24438,N_24695);
and U25114 (N_25114,N_24895,N_24514);
xor U25115 (N_25115,N_24779,N_24666);
nor U25116 (N_25116,N_24157,N_24893);
nand U25117 (N_25117,N_24636,N_24959);
nor U25118 (N_25118,N_24445,N_24185);
or U25119 (N_25119,N_24289,N_24583);
nand U25120 (N_25120,N_24838,N_24767);
nor U25121 (N_25121,N_24939,N_24096);
nand U25122 (N_25122,N_24674,N_24164);
xor U25123 (N_25123,N_24653,N_24190);
or U25124 (N_25124,N_24741,N_24100);
and U25125 (N_25125,N_24234,N_24881);
nand U25126 (N_25126,N_24298,N_24277);
nor U25127 (N_25127,N_24883,N_24539);
or U25128 (N_25128,N_24295,N_24115);
nand U25129 (N_25129,N_24791,N_24183);
nand U25130 (N_25130,N_24765,N_24271);
nor U25131 (N_25131,N_24454,N_24257);
or U25132 (N_25132,N_24629,N_24084);
xor U25133 (N_25133,N_24801,N_24427);
xnor U25134 (N_25134,N_24128,N_24549);
and U25135 (N_25135,N_24230,N_24667);
xnor U25136 (N_25136,N_24508,N_24753);
and U25137 (N_25137,N_24165,N_24846);
xnor U25138 (N_25138,N_24871,N_24093);
xnor U25139 (N_25139,N_24607,N_24647);
and U25140 (N_25140,N_24303,N_24914);
nor U25141 (N_25141,N_24170,N_24006);
nand U25142 (N_25142,N_24682,N_24087);
or U25143 (N_25143,N_24809,N_24215);
nand U25144 (N_25144,N_24865,N_24625);
nor U25145 (N_25145,N_24442,N_24343);
xor U25146 (N_25146,N_24080,N_24994);
nand U25147 (N_25147,N_24162,N_24076);
or U25148 (N_25148,N_24275,N_24404);
nand U25149 (N_25149,N_24841,N_24670);
nor U25150 (N_25150,N_24112,N_24187);
xnor U25151 (N_25151,N_24141,N_24143);
and U25152 (N_25152,N_24596,N_24272);
or U25153 (N_25153,N_24713,N_24668);
xor U25154 (N_25154,N_24310,N_24941);
xor U25155 (N_25155,N_24108,N_24339);
nand U25156 (N_25156,N_24567,N_24665);
and U25157 (N_25157,N_24370,N_24817);
nand U25158 (N_25158,N_24444,N_24325);
nand U25159 (N_25159,N_24274,N_24952);
xor U25160 (N_25160,N_24894,N_24616);
nor U25161 (N_25161,N_24389,N_24519);
or U25162 (N_25162,N_24201,N_24304);
nor U25163 (N_25163,N_24656,N_24499);
and U25164 (N_25164,N_24973,N_24589);
and U25165 (N_25165,N_24182,N_24547);
nor U25166 (N_25166,N_24725,N_24527);
and U25167 (N_25167,N_24059,N_24528);
or U25168 (N_25168,N_24262,N_24278);
or U25169 (N_25169,N_24908,N_24061);
or U25170 (N_25170,N_24120,N_24749);
nand U25171 (N_25171,N_24912,N_24375);
nand U25172 (N_25172,N_24759,N_24005);
and U25173 (N_25173,N_24488,N_24655);
and U25174 (N_25174,N_24481,N_24658);
xor U25175 (N_25175,N_24998,N_24615);
nand U25176 (N_25176,N_24761,N_24516);
xor U25177 (N_25177,N_24732,N_24855);
nand U25178 (N_25178,N_24965,N_24152);
and U25179 (N_25179,N_24208,N_24229);
nand U25180 (N_25180,N_24015,N_24147);
xor U25181 (N_25181,N_24568,N_24191);
nand U25182 (N_25182,N_24696,N_24859);
nor U25183 (N_25183,N_24854,N_24879);
nor U25184 (N_25184,N_24569,N_24027);
nor U25185 (N_25185,N_24632,N_24038);
xnor U25186 (N_25186,N_24158,N_24391);
or U25187 (N_25187,N_24748,N_24690);
nand U25188 (N_25188,N_24750,N_24614);
and U25189 (N_25189,N_24953,N_24039);
and U25190 (N_25190,N_24378,N_24506);
or U25191 (N_25191,N_24680,N_24288);
xor U25192 (N_25192,N_24543,N_24221);
and U25193 (N_25193,N_24736,N_24313);
and U25194 (N_25194,N_24553,N_24798);
xor U25195 (N_25195,N_24011,N_24802);
nand U25196 (N_25196,N_24882,N_24012);
xor U25197 (N_25197,N_24950,N_24205);
nand U25198 (N_25198,N_24827,N_24979);
and U25199 (N_25199,N_24328,N_24931);
xnor U25200 (N_25200,N_24362,N_24613);
xnor U25201 (N_25201,N_24905,N_24788);
nand U25202 (N_25202,N_24580,N_24460);
and U25203 (N_25203,N_24306,N_24526);
and U25204 (N_25204,N_24662,N_24021);
nor U25205 (N_25205,N_24721,N_24919);
and U25206 (N_25206,N_24273,N_24776);
and U25207 (N_25207,N_24218,N_24520);
or U25208 (N_25208,N_24876,N_24806);
xor U25209 (N_25209,N_24963,N_24148);
and U25210 (N_25210,N_24573,N_24322);
nor U25211 (N_25211,N_24425,N_24623);
nor U25212 (N_25212,N_24287,N_24054);
nand U25213 (N_25213,N_24408,N_24728);
nand U25214 (N_25214,N_24127,N_24678);
nor U25215 (N_25215,N_24174,N_24804);
nor U25216 (N_25216,N_24727,N_24906);
and U25217 (N_25217,N_24052,N_24631);
xnor U25218 (N_25218,N_24001,N_24576);
nand U25219 (N_25219,N_24204,N_24316);
xor U25220 (N_25220,N_24498,N_24415);
nor U25221 (N_25221,N_24473,N_24243);
xor U25222 (N_25222,N_24822,N_24851);
nor U25223 (N_25223,N_24013,N_24207);
or U25224 (N_25224,N_24123,N_24534);
xnor U25225 (N_25225,N_24676,N_24714);
xnor U25226 (N_25226,N_24333,N_24099);
and U25227 (N_25227,N_24790,N_24297);
nor U25228 (N_25228,N_24915,N_24238);
nor U25229 (N_25229,N_24660,N_24171);
xor U25230 (N_25230,N_24037,N_24245);
or U25231 (N_25231,N_24999,N_24210);
xor U25232 (N_25232,N_24742,N_24196);
or U25233 (N_25233,N_24811,N_24002);
or U25234 (N_25234,N_24975,N_24432);
xor U25235 (N_25235,N_24113,N_24672);
xnor U25236 (N_25236,N_24311,N_24637);
nor U25237 (N_25237,N_24624,N_24816);
nand U25238 (N_25238,N_24449,N_24186);
xnor U25239 (N_25239,N_24320,N_24067);
nor U25240 (N_25240,N_24715,N_24216);
nor U25241 (N_25241,N_24177,N_24223);
nand U25242 (N_25242,N_24500,N_24146);
or U25243 (N_25243,N_24269,N_24225);
and U25244 (N_25244,N_24675,N_24650);
nor U25245 (N_25245,N_24371,N_24467);
and U25246 (N_25246,N_24490,N_24996);
nor U25247 (N_25247,N_24593,N_24064);
or U25248 (N_25248,N_24423,N_24397);
and U25249 (N_25249,N_24828,N_24775);
nand U25250 (N_25250,N_24261,N_24484);
nand U25251 (N_25251,N_24943,N_24497);
xnor U25252 (N_25252,N_24348,N_24661);
and U25253 (N_25253,N_24595,N_24869);
nand U25254 (N_25254,N_24051,N_24835);
and U25255 (N_25255,N_24807,N_24521);
xnor U25256 (N_25256,N_24192,N_24487);
and U25257 (N_25257,N_24003,N_24103);
nor U25258 (N_25258,N_24307,N_24424);
nor U25259 (N_25259,N_24055,N_24368);
nand U25260 (N_25260,N_24247,N_24692);
nor U25261 (N_25261,N_24073,N_24927);
xnor U25262 (N_25262,N_24991,N_24319);
xor U25263 (N_25263,N_24384,N_24823);
and U25264 (N_25264,N_24898,N_24125);
and U25265 (N_25265,N_24160,N_24834);
nor U25266 (N_25266,N_24299,N_24119);
nand U25267 (N_25267,N_24639,N_24340);
nor U25268 (N_25268,N_24902,N_24010);
nor U25269 (N_25269,N_24078,N_24403);
or U25270 (N_25270,N_24448,N_24474);
nor U25271 (N_25271,N_24292,N_24993);
nor U25272 (N_25272,N_24980,N_24852);
xnor U25273 (N_25273,N_24453,N_24899);
or U25274 (N_25274,N_24142,N_24451);
and U25275 (N_25275,N_24172,N_24441);
nor U25276 (N_25276,N_24644,N_24844);
xnor U25277 (N_25277,N_24461,N_24417);
xnor U25278 (N_25278,N_24837,N_24377);
and U25279 (N_25279,N_24818,N_24787);
nand U25280 (N_25280,N_24664,N_24264);
xor U25281 (N_25281,N_24754,N_24267);
or U25282 (N_25282,N_24584,N_24020);
nand U25283 (N_25283,N_24360,N_24669);
nand U25284 (N_25284,N_24222,N_24955);
nor U25285 (N_25285,N_24849,N_24535);
nor U25286 (N_25286,N_24990,N_24380);
xor U25287 (N_25287,N_24988,N_24740);
and U25288 (N_25288,N_24098,N_24739);
nor U25289 (N_25289,N_24227,N_24634);
xor U25290 (N_25290,N_24060,N_24226);
and U25291 (N_25291,N_24574,N_24188);
xnor U25292 (N_25292,N_24305,N_24341);
nand U25293 (N_25293,N_24133,N_24813);
nand U25294 (N_25294,N_24570,N_24556);
nand U25295 (N_25295,N_24770,N_24491);
or U25296 (N_25296,N_24452,N_24373);
or U25297 (N_25297,N_24766,N_24300);
or U25298 (N_25298,N_24974,N_24923);
xor U25299 (N_25299,N_24024,N_24904);
xor U25300 (N_25300,N_24735,N_24411);
or U25301 (N_25301,N_24419,N_24312);
xor U25302 (N_25302,N_24603,N_24815);
or U25303 (N_25303,N_24203,N_24110);
and U25304 (N_25304,N_24586,N_24450);
nor U25305 (N_25305,N_24422,N_24874);
or U25306 (N_25306,N_24407,N_24546);
and U25307 (N_25307,N_24410,N_24246);
and U25308 (N_25308,N_24358,N_24651);
or U25309 (N_25309,N_24601,N_24258);
or U25310 (N_25310,N_24983,N_24045);
and U25311 (N_25311,N_24698,N_24718);
or U25312 (N_25312,N_24608,N_24850);
xnor U25313 (N_25313,N_24733,N_24156);
xnor U25314 (N_25314,N_24058,N_24706);
and U25315 (N_25315,N_24000,N_24872);
xor U25316 (N_25316,N_24236,N_24585);
xnor U25317 (N_25317,N_24956,N_24374);
nor U25318 (N_25318,N_24774,N_24232);
xnor U25319 (N_25319,N_24752,N_24475);
xnor U25320 (N_25320,N_24916,N_24518);
nand U25321 (N_25321,N_24560,N_24046);
nand U25322 (N_25322,N_24805,N_24532);
or U25323 (N_25323,N_24591,N_24960);
xor U25324 (N_25324,N_24609,N_24266);
xor U25325 (N_25325,N_24799,N_24065);
and U25326 (N_25326,N_24372,N_24856);
xnor U25327 (N_25327,N_24383,N_24892);
and U25328 (N_25328,N_24942,N_24981);
nor U25329 (N_25329,N_24116,N_24705);
and U25330 (N_25330,N_24421,N_24842);
nand U25331 (N_25331,N_24800,N_24579);
nor U25332 (N_25332,N_24700,N_24168);
nand U25333 (N_25333,N_24935,N_24909);
nand U25334 (N_25334,N_24434,N_24756);
xor U25335 (N_25335,N_24771,N_24877);
or U25336 (N_25336,N_24462,N_24029);
nor U25337 (N_25337,N_24551,N_24161);
xor U25338 (N_25338,N_24977,N_24968);
or U25339 (N_25339,N_24092,N_24880);
and U25340 (N_25340,N_24179,N_24286);
and U25341 (N_25341,N_24982,N_24184);
xnor U25342 (N_25342,N_24875,N_24782);
nand U25343 (N_25343,N_24957,N_24040);
xor U25344 (N_25344,N_24683,N_24326);
and U25345 (N_25345,N_24472,N_24934);
or U25346 (N_25346,N_24413,N_24870);
and U25347 (N_25347,N_24132,N_24387);
and U25348 (N_25348,N_24323,N_24768);
nor U25349 (N_25349,N_24332,N_24810);
nand U25350 (N_25350,N_24590,N_24604);
nor U25351 (N_25351,N_24920,N_24561);
nand U25352 (N_25352,N_24984,N_24478);
nor U25353 (N_25353,N_24562,N_24620);
or U25354 (N_25354,N_24173,N_24014);
and U25355 (N_25355,N_24566,N_24511);
xnor U25356 (N_25356,N_24509,N_24602);
and U25357 (N_25357,N_24279,N_24704);
or U25358 (N_25358,N_24137,N_24971);
and U25359 (N_25359,N_24195,N_24420);
or U25360 (N_25360,N_24367,N_24376);
and U25361 (N_25361,N_24711,N_24118);
or U25362 (N_25362,N_24181,N_24536);
or U25363 (N_25363,N_24219,N_24228);
xnor U25364 (N_25364,N_24503,N_24540);
or U25365 (N_25365,N_24897,N_24954);
nor U25366 (N_25366,N_24886,N_24198);
nand U25367 (N_25367,N_24471,N_24889);
nor U25368 (N_25368,N_24072,N_24086);
and U25369 (N_25369,N_24679,N_24707);
or U25370 (N_25370,N_24578,N_24793);
and U25371 (N_25371,N_24839,N_24327);
nor U25372 (N_25372,N_24290,N_24863);
nor U25373 (N_25373,N_24483,N_24250);
xor U25374 (N_25374,N_24868,N_24611);
nor U25375 (N_25375,N_24594,N_24138);
nand U25376 (N_25376,N_24126,N_24840);
xnor U25377 (N_25377,N_24612,N_24719);
and U25378 (N_25378,N_24533,N_24400);
xnor U25379 (N_25379,N_24948,N_24884);
or U25380 (N_25380,N_24684,N_24347);
xor U25381 (N_25381,N_24265,N_24254);
xnor U25382 (N_25382,N_24044,N_24989);
nor U25383 (N_25383,N_24524,N_24769);
and U25384 (N_25384,N_24334,N_24987);
xnor U25385 (N_25385,N_24778,N_24517);
nor U25386 (N_25386,N_24022,N_24764);
xor U25387 (N_25387,N_24947,N_24992);
and U25388 (N_25388,N_24053,N_24502);
nand U25389 (N_25389,N_24057,N_24627);
and U25390 (N_25390,N_24821,N_24703);
or U25391 (N_25391,N_24792,N_24056);
and U25392 (N_25392,N_24866,N_24318);
xnor U25393 (N_25393,N_24691,N_24716);
or U25394 (N_25394,N_24036,N_24068);
or U25395 (N_25395,N_24744,N_24933);
or U25396 (N_25396,N_24239,N_24762);
nand U25397 (N_25397,N_24263,N_24189);
or U25398 (N_25398,N_24494,N_24575);
or U25399 (N_25399,N_24097,N_24630);
xnor U25400 (N_25400,N_24430,N_24331);
nor U25401 (N_25401,N_24924,N_24577);
nor U25402 (N_25402,N_24041,N_24048);
nand U25403 (N_25403,N_24652,N_24944);
xor U25404 (N_25404,N_24075,N_24069);
and U25405 (N_25405,N_24864,N_24396);
or U25406 (N_25406,N_24446,N_24049);
and U25407 (N_25407,N_24925,N_24890);
or U25408 (N_25408,N_24091,N_24176);
or U25409 (N_25409,N_24710,N_24495);
nor U25410 (N_25410,N_24004,N_24610);
xor U25411 (N_25411,N_24104,N_24878);
xnor U25412 (N_25412,N_24642,N_24734);
xnor U25413 (N_25413,N_24541,N_24217);
or U25414 (N_25414,N_24163,N_24043);
or U25415 (N_25415,N_24090,N_24592);
and U25416 (N_25416,N_24095,N_24276);
and U25417 (N_25417,N_24390,N_24701);
nand U25418 (N_25418,N_24070,N_24106);
xor U25419 (N_25419,N_24833,N_24640);
or U25420 (N_25420,N_24167,N_24082);
nor U25421 (N_25421,N_24751,N_24940);
nor U25422 (N_25422,N_24819,N_24159);
nand U25423 (N_25423,N_24785,N_24259);
nand U25424 (N_25424,N_24429,N_24588);
nor U25425 (N_25425,N_24242,N_24694);
nor U25426 (N_25426,N_24628,N_24253);
nor U25427 (N_25427,N_24530,N_24572);
and U25428 (N_25428,N_24832,N_24197);
or U25429 (N_25429,N_24773,N_24867);
xor U25430 (N_25430,N_24814,N_24028);
nor U25431 (N_25431,N_24937,N_24169);
or U25432 (N_25432,N_24784,N_24042);
or U25433 (N_25433,N_24843,N_24758);
and U25434 (N_25434,N_24026,N_24829);
xor U25435 (N_25435,N_24468,N_24281);
xnor U25436 (N_25436,N_24439,N_24581);
and U25437 (N_25437,N_24803,N_24455);
nand U25438 (N_25438,N_24294,N_24928);
nand U25439 (N_25439,N_24401,N_24329);
nor U25440 (N_25440,N_24285,N_24135);
and U25441 (N_25441,N_24738,N_24465);
nand U25442 (N_25442,N_24379,N_24050);
nand U25443 (N_25443,N_24235,N_24268);
nor U25444 (N_25444,N_24324,N_24795);
xor U25445 (N_25445,N_24081,N_24395);
xor U25446 (N_25446,N_24921,N_24342);
nand U25447 (N_25447,N_24936,N_24820);
nor U25448 (N_25448,N_24621,N_24194);
nor U25449 (N_25449,N_24200,N_24023);
or U25450 (N_25450,N_24626,N_24945);
nand U25451 (N_25451,N_24309,N_24352);
nor U25452 (N_25452,N_24896,N_24911);
and U25453 (N_25453,N_24130,N_24605);
or U25454 (N_25454,N_24317,N_24155);
xnor U25455 (N_25455,N_24107,N_24405);
nor U25456 (N_25456,N_24693,N_24393);
and U25457 (N_25457,N_24780,N_24544);
nand U25458 (N_25458,N_24986,N_24789);
and U25459 (N_25459,N_24797,N_24958);
and U25460 (N_25460,N_24903,N_24129);
or U25461 (N_25461,N_24016,N_24252);
nand U25462 (N_25462,N_24972,N_24456);
or U25463 (N_25463,N_24858,N_24033);
nor U25464 (N_25464,N_24571,N_24102);
and U25465 (N_25465,N_24663,N_24437);
xnor U25466 (N_25466,N_24505,N_24951);
xor U25467 (N_25467,N_24280,N_24677);
and U25468 (N_25468,N_24031,N_24346);
or U25469 (N_25469,N_24538,N_24089);
nand U25470 (N_25470,N_24746,N_24314);
or U25471 (N_25471,N_24175,N_24083);
nand U25472 (N_25472,N_24743,N_24355);
xor U25473 (N_25473,N_24657,N_24830);
or U25474 (N_25474,N_24321,N_24436);
xnor U25475 (N_25475,N_24489,N_24760);
and U25476 (N_25476,N_24643,N_24047);
and U25477 (N_25477,N_24847,N_24335);
or U25478 (N_25478,N_24545,N_24062);
or U25479 (N_25479,N_24485,N_24017);
or U25480 (N_25480,N_24114,N_24213);
or U25481 (N_25481,N_24457,N_24244);
and U25482 (N_25482,N_24970,N_24428);
and U25483 (N_25483,N_24018,N_24641);
nor U25484 (N_25484,N_24726,N_24985);
nor U25485 (N_25485,N_24873,N_24599);
nand U25486 (N_25486,N_24600,N_24409);
or U25487 (N_25487,N_24635,N_24364);
xnor U25488 (N_25488,N_24638,N_24557);
or U25489 (N_25489,N_24447,N_24007);
nor U25490 (N_25490,N_24202,N_24479);
and U25491 (N_25491,N_24030,N_24282);
or U25492 (N_25492,N_24369,N_24796);
and U25493 (N_25493,N_24633,N_24997);
nor U25494 (N_25494,N_24598,N_24808);
xnor U25495 (N_25495,N_24394,N_24032);
nand U25496 (N_25496,N_24009,N_24193);
nor U25497 (N_25497,N_24392,N_24929);
xnor U25498 (N_25498,N_24151,N_24237);
nor U25499 (N_25499,N_24121,N_24211);
xnor U25500 (N_25500,N_24496,N_24411);
xor U25501 (N_25501,N_24650,N_24821);
xor U25502 (N_25502,N_24818,N_24378);
nor U25503 (N_25503,N_24769,N_24836);
xor U25504 (N_25504,N_24631,N_24428);
xor U25505 (N_25505,N_24085,N_24046);
xor U25506 (N_25506,N_24379,N_24732);
nor U25507 (N_25507,N_24438,N_24483);
xnor U25508 (N_25508,N_24603,N_24951);
nor U25509 (N_25509,N_24828,N_24467);
or U25510 (N_25510,N_24892,N_24446);
xnor U25511 (N_25511,N_24737,N_24741);
nor U25512 (N_25512,N_24585,N_24829);
nor U25513 (N_25513,N_24746,N_24286);
nand U25514 (N_25514,N_24945,N_24622);
and U25515 (N_25515,N_24211,N_24132);
or U25516 (N_25516,N_24561,N_24257);
xor U25517 (N_25517,N_24424,N_24760);
or U25518 (N_25518,N_24889,N_24682);
nor U25519 (N_25519,N_24317,N_24811);
nand U25520 (N_25520,N_24538,N_24471);
nand U25521 (N_25521,N_24151,N_24461);
nand U25522 (N_25522,N_24519,N_24411);
nor U25523 (N_25523,N_24172,N_24314);
and U25524 (N_25524,N_24715,N_24134);
nor U25525 (N_25525,N_24004,N_24892);
xnor U25526 (N_25526,N_24532,N_24987);
or U25527 (N_25527,N_24533,N_24476);
or U25528 (N_25528,N_24931,N_24003);
xor U25529 (N_25529,N_24113,N_24784);
and U25530 (N_25530,N_24116,N_24039);
nand U25531 (N_25531,N_24501,N_24298);
xnor U25532 (N_25532,N_24844,N_24462);
xor U25533 (N_25533,N_24577,N_24667);
nand U25534 (N_25534,N_24605,N_24340);
or U25535 (N_25535,N_24658,N_24386);
and U25536 (N_25536,N_24024,N_24911);
nor U25537 (N_25537,N_24324,N_24765);
and U25538 (N_25538,N_24741,N_24706);
and U25539 (N_25539,N_24116,N_24805);
or U25540 (N_25540,N_24244,N_24064);
or U25541 (N_25541,N_24924,N_24399);
nor U25542 (N_25542,N_24909,N_24137);
and U25543 (N_25543,N_24485,N_24786);
xor U25544 (N_25544,N_24176,N_24485);
xnor U25545 (N_25545,N_24173,N_24845);
nor U25546 (N_25546,N_24139,N_24023);
nand U25547 (N_25547,N_24821,N_24556);
or U25548 (N_25548,N_24368,N_24821);
and U25549 (N_25549,N_24240,N_24811);
nand U25550 (N_25550,N_24912,N_24224);
or U25551 (N_25551,N_24668,N_24395);
nor U25552 (N_25552,N_24268,N_24140);
xor U25553 (N_25553,N_24730,N_24270);
nand U25554 (N_25554,N_24519,N_24400);
nor U25555 (N_25555,N_24977,N_24511);
nor U25556 (N_25556,N_24211,N_24709);
nor U25557 (N_25557,N_24279,N_24074);
nand U25558 (N_25558,N_24059,N_24333);
nand U25559 (N_25559,N_24528,N_24436);
or U25560 (N_25560,N_24986,N_24278);
xor U25561 (N_25561,N_24221,N_24998);
or U25562 (N_25562,N_24984,N_24300);
nand U25563 (N_25563,N_24998,N_24560);
or U25564 (N_25564,N_24946,N_24150);
and U25565 (N_25565,N_24877,N_24698);
nand U25566 (N_25566,N_24684,N_24972);
or U25567 (N_25567,N_24702,N_24129);
nand U25568 (N_25568,N_24123,N_24733);
nor U25569 (N_25569,N_24550,N_24889);
xnor U25570 (N_25570,N_24952,N_24298);
and U25571 (N_25571,N_24321,N_24722);
nand U25572 (N_25572,N_24344,N_24302);
nor U25573 (N_25573,N_24442,N_24703);
xnor U25574 (N_25574,N_24472,N_24593);
xor U25575 (N_25575,N_24104,N_24245);
nor U25576 (N_25576,N_24695,N_24089);
nor U25577 (N_25577,N_24152,N_24681);
and U25578 (N_25578,N_24270,N_24626);
nand U25579 (N_25579,N_24116,N_24642);
and U25580 (N_25580,N_24582,N_24873);
nand U25581 (N_25581,N_24874,N_24121);
or U25582 (N_25582,N_24458,N_24988);
or U25583 (N_25583,N_24699,N_24752);
xor U25584 (N_25584,N_24644,N_24544);
xnor U25585 (N_25585,N_24371,N_24174);
xnor U25586 (N_25586,N_24749,N_24882);
xnor U25587 (N_25587,N_24607,N_24845);
and U25588 (N_25588,N_24419,N_24036);
nand U25589 (N_25589,N_24339,N_24218);
nor U25590 (N_25590,N_24173,N_24239);
nand U25591 (N_25591,N_24661,N_24953);
and U25592 (N_25592,N_24915,N_24699);
nor U25593 (N_25593,N_24935,N_24373);
xor U25594 (N_25594,N_24233,N_24296);
xor U25595 (N_25595,N_24444,N_24606);
and U25596 (N_25596,N_24891,N_24378);
or U25597 (N_25597,N_24526,N_24961);
xnor U25598 (N_25598,N_24914,N_24335);
nor U25599 (N_25599,N_24272,N_24023);
nand U25600 (N_25600,N_24856,N_24708);
xor U25601 (N_25601,N_24790,N_24440);
or U25602 (N_25602,N_24679,N_24825);
xor U25603 (N_25603,N_24528,N_24176);
nand U25604 (N_25604,N_24691,N_24442);
or U25605 (N_25605,N_24688,N_24218);
or U25606 (N_25606,N_24789,N_24377);
nand U25607 (N_25607,N_24530,N_24928);
and U25608 (N_25608,N_24847,N_24936);
and U25609 (N_25609,N_24458,N_24387);
or U25610 (N_25610,N_24413,N_24453);
xnor U25611 (N_25611,N_24264,N_24774);
xnor U25612 (N_25612,N_24040,N_24562);
nor U25613 (N_25613,N_24281,N_24736);
nand U25614 (N_25614,N_24958,N_24183);
xnor U25615 (N_25615,N_24282,N_24816);
or U25616 (N_25616,N_24461,N_24081);
nand U25617 (N_25617,N_24118,N_24372);
nor U25618 (N_25618,N_24689,N_24558);
nand U25619 (N_25619,N_24434,N_24068);
xnor U25620 (N_25620,N_24955,N_24933);
xnor U25621 (N_25621,N_24926,N_24958);
xnor U25622 (N_25622,N_24388,N_24724);
and U25623 (N_25623,N_24802,N_24455);
nand U25624 (N_25624,N_24586,N_24231);
xnor U25625 (N_25625,N_24247,N_24290);
nand U25626 (N_25626,N_24176,N_24992);
nand U25627 (N_25627,N_24622,N_24736);
or U25628 (N_25628,N_24379,N_24511);
nand U25629 (N_25629,N_24841,N_24402);
xor U25630 (N_25630,N_24751,N_24373);
nand U25631 (N_25631,N_24735,N_24009);
nor U25632 (N_25632,N_24597,N_24483);
and U25633 (N_25633,N_24818,N_24089);
nor U25634 (N_25634,N_24249,N_24923);
nor U25635 (N_25635,N_24586,N_24750);
xnor U25636 (N_25636,N_24417,N_24241);
and U25637 (N_25637,N_24630,N_24285);
or U25638 (N_25638,N_24287,N_24384);
and U25639 (N_25639,N_24189,N_24118);
or U25640 (N_25640,N_24861,N_24513);
and U25641 (N_25641,N_24317,N_24567);
nor U25642 (N_25642,N_24186,N_24831);
or U25643 (N_25643,N_24174,N_24146);
and U25644 (N_25644,N_24191,N_24774);
nor U25645 (N_25645,N_24258,N_24205);
nor U25646 (N_25646,N_24839,N_24107);
nand U25647 (N_25647,N_24384,N_24418);
xor U25648 (N_25648,N_24134,N_24086);
or U25649 (N_25649,N_24213,N_24482);
or U25650 (N_25650,N_24094,N_24455);
and U25651 (N_25651,N_24259,N_24961);
xnor U25652 (N_25652,N_24843,N_24397);
and U25653 (N_25653,N_24001,N_24111);
xnor U25654 (N_25654,N_24574,N_24259);
nand U25655 (N_25655,N_24337,N_24956);
nand U25656 (N_25656,N_24776,N_24634);
or U25657 (N_25657,N_24873,N_24551);
and U25658 (N_25658,N_24569,N_24733);
nor U25659 (N_25659,N_24052,N_24302);
nand U25660 (N_25660,N_24895,N_24867);
and U25661 (N_25661,N_24142,N_24973);
nand U25662 (N_25662,N_24918,N_24851);
or U25663 (N_25663,N_24875,N_24184);
or U25664 (N_25664,N_24734,N_24567);
or U25665 (N_25665,N_24246,N_24775);
and U25666 (N_25666,N_24806,N_24386);
and U25667 (N_25667,N_24147,N_24726);
nor U25668 (N_25668,N_24418,N_24238);
or U25669 (N_25669,N_24529,N_24616);
nand U25670 (N_25670,N_24589,N_24742);
and U25671 (N_25671,N_24258,N_24093);
nand U25672 (N_25672,N_24651,N_24640);
xnor U25673 (N_25673,N_24676,N_24991);
or U25674 (N_25674,N_24356,N_24315);
nand U25675 (N_25675,N_24904,N_24705);
xor U25676 (N_25676,N_24485,N_24742);
xor U25677 (N_25677,N_24801,N_24516);
nor U25678 (N_25678,N_24500,N_24074);
and U25679 (N_25679,N_24387,N_24938);
xor U25680 (N_25680,N_24699,N_24019);
nand U25681 (N_25681,N_24339,N_24402);
or U25682 (N_25682,N_24007,N_24621);
nor U25683 (N_25683,N_24779,N_24157);
and U25684 (N_25684,N_24771,N_24026);
nand U25685 (N_25685,N_24403,N_24387);
nor U25686 (N_25686,N_24757,N_24249);
and U25687 (N_25687,N_24740,N_24248);
nand U25688 (N_25688,N_24053,N_24224);
or U25689 (N_25689,N_24171,N_24261);
nand U25690 (N_25690,N_24188,N_24458);
nand U25691 (N_25691,N_24844,N_24271);
and U25692 (N_25692,N_24233,N_24137);
nand U25693 (N_25693,N_24401,N_24151);
nand U25694 (N_25694,N_24557,N_24282);
nor U25695 (N_25695,N_24674,N_24619);
or U25696 (N_25696,N_24871,N_24279);
and U25697 (N_25697,N_24418,N_24803);
and U25698 (N_25698,N_24531,N_24276);
or U25699 (N_25699,N_24360,N_24276);
or U25700 (N_25700,N_24281,N_24011);
nor U25701 (N_25701,N_24130,N_24949);
nand U25702 (N_25702,N_24316,N_24837);
nor U25703 (N_25703,N_24125,N_24960);
or U25704 (N_25704,N_24751,N_24057);
or U25705 (N_25705,N_24915,N_24419);
and U25706 (N_25706,N_24011,N_24755);
xor U25707 (N_25707,N_24953,N_24453);
and U25708 (N_25708,N_24954,N_24652);
xor U25709 (N_25709,N_24526,N_24104);
nand U25710 (N_25710,N_24309,N_24394);
xnor U25711 (N_25711,N_24151,N_24994);
and U25712 (N_25712,N_24523,N_24164);
and U25713 (N_25713,N_24917,N_24674);
nor U25714 (N_25714,N_24220,N_24410);
and U25715 (N_25715,N_24508,N_24425);
xnor U25716 (N_25716,N_24930,N_24730);
and U25717 (N_25717,N_24267,N_24191);
nand U25718 (N_25718,N_24061,N_24172);
nand U25719 (N_25719,N_24577,N_24412);
nor U25720 (N_25720,N_24999,N_24373);
xor U25721 (N_25721,N_24559,N_24783);
nor U25722 (N_25722,N_24374,N_24501);
nand U25723 (N_25723,N_24072,N_24348);
xnor U25724 (N_25724,N_24560,N_24210);
or U25725 (N_25725,N_24997,N_24049);
and U25726 (N_25726,N_24205,N_24953);
nand U25727 (N_25727,N_24796,N_24351);
and U25728 (N_25728,N_24982,N_24269);
or U25729 (N_25729,N_24884,N_24840);
nor U25730 (N_25730,N_24262,N_24153);
or U25731 (N_25731,N_24245,N_24027);
or U25732 (N_25732,N_24380,N_24224);
nand U25733 (N_25733,N_24774,N_24158);
xnor U25734 (N_25734,N_24503,N_24329);
xnor U25735 (N_25735,N_24130,N_24391);
xnor U25736 (N_25736,N_24828,N_24038);
nor U25737 (N_25737,N_24996,N_24416);
nand U25738 (N_25738,N_24051,N_24752);
or U25739 (N_25739,N_24180,N_24333);
nor U25740 (N_25740,N_24463,N_24090);
nand U25741 (N_25741,N_24173,N_24548);
or U25742 (N_25742,N_24007,N_24954);
nor U25743 (N_25743,N_24165,N_24659);
nand U25744 (N_25744,N_24109,N_24372);
or U25745 (N_25745,N_24677,N_24661);
or U25746 (N_25746,N_24012,N_24420);
nand U25747 (N_25747,N_24957,N_24650);
or U25748 (N_25748,N_24098,N_24205);
and U25749 (N_25749,N_24846,N_24004);
xnor U25750 (N_25750,N_24765,N_24148);
and U25751 (N_25751,N_24147,N_24548);
or U25752 (N_25752,N_24299,N_24357);
nor U25753 (N_25753,N_24340,N_24076);
and U25754 (N_25754,N_24495,N_24380);
nor U25755 (N_25755,N_24118,N_24634);
nor U25756 (N_25756,N_24971,N_24253);
and U25757 (N_25757,N_24708,N_24547);
nor U25758 (N_25758,N_24028,N_24877);
or U25759 (N_25759,N_24940,N_24723);
nand U25760 (N_25760,N_24900,N_24201);
nor U25761 (N_25761,N_24975,N_24830);
nor U25762 (N_25762,N_24203,N_24059);
nand U25763 (N_25763,N_24158,N_24279);
xor U25764 (N_25764,N_24784,N_24819);
xnor U25765 (N_25765,N_24063,N_24425);
xnor U25766 (N_25766,N_24665,N_24109);
and U25767 (N_25767,N_24246,N_24085);
or U25768 (N_25768,N_24257,N_24141);
xor U25769 (N_25769,N_24076,N_24937);
nand U25770 (N_25770,N_24406,N_24551);
or U25771 (N_25771,N_24143,N_24510);
nor U25772 (N_25772,N_24540,N_24939);
xor U25773 (N_25773,N_24990,N_24743);
xor U25774 (N_25774,N_24410,N_24023);
or U25775 (N_25775,N_24718,N_24571);
xnor U25776 (N_25776,N_24446,N_24674);
nand U25777 (N_25777,N_24248,N_24886);
or U25778 (N_25778,N_24602,N_24370);
or U25779 (N_25779,N_24064,N_24197);
and U25780 (N_25780,N_24002,N_24052);
nor U25781 (N_25781,N_24225,N_24455);
nor U25782 (N_25782,N_24953,N_24779);
xor U25783 (N_25783,N_24288,N_24730);
nand U25784 (N_25784,N_24036,N_24019);
or U25785 (N_25785,N_24450,N_24264);
xnor U25786 (N_25786,N_24917,N_24033);
and U25787 (N_25787,N_24859,N_24955);
and U25788 (N_25788,N_24511,N_24010);
and U25789 (N_25789,N_24802,N_24970);
and U25790 (N_25790,N_24682,N_24841);
or U25791 (N_25791,N_24436,N_24774);
or U25792 (N_25792,N_24440,N_24815);
nor U25793 (N_25793,N_24750,N_24456);
or U25794 (N_25794,N_24739,N_24668);
nor U25795 (N_25795,N_24563,N_24484);
nand U25796 (N_25796,N_24160,N_24503);
and U25797 (N_25797,N_24675,N_24844);
xnor U25798 (N_25798,N_24885,N_24966);
and U25799 (N_25799,N_24378,N_24200);
xor U25800 (N_25800,N_24069,N_24121);
xnor U25801 (N_25801,N_24322,N_24907);
nand U25802 (N_25802,N_24653,N_24083);
and U25803 (N_25803,N_24868,N_24018);
xnor U25804 (N_25804,N_24742,N_24054);
nor U25805 (N_25805,N_24548,N_24550);
and U25806 (N_25806,N_24934,N_24911);
xnor U25807 (N_25807,N_24284,N_24059);
or U25808 (N_25808,N_24868,N_24102);
nand U25809 (N_25809,N_24747,N_24240);
or U25810 (N_25810,N_24780,N_24853);
or U25811 (N_25811,N_24995,N_24202);
nor U25812 (N_25812,N_24119,N_24141);
nor U25813 (N_25813,N_24877,N_24842);
nor U25814 (N_25814,N_24264,N_24218);
and U25815 (N_25815,N_24316,N_24968);
nand U25816 (N_25816,N_24805,N_24332);
or U25817 (N_25817,N_24756,N_24388);
xnor U25818 (N_25818,N_24525,N_24875);
xor U25819 (N_25819,N_24300,N_24641);
or U25820 (N_25820,N_24118,N_24046);
xnor U25821 (N_25821,N_24959,N_24288);
nor U25822 (N_25822,N_24858,N_24126);
or U25823 (N_25823,N_24573,N_24832);
nand U25824 (N_25824,N_24774,N_24248);
nor U25825 (N_25825,N_24313,N_24368);
xnor U25826 (N_25826,N_24382,N_24601);
nor U25827 (N_25827,N_24180,N_24733);
and U25828 (N_25828,N_24900,N_24709);
xnor U25829 (N_25829,N_24150,N_24399);
xnor U25830 (N_25830,N_24644,N_24782);
nand U25831 (N_25831,N_24011,N_24259);
and U25832 (N_25832,N_24432,N_24859);
nor U25833 (N_25833,N_24794,N_24891);
nand U25834 (N_25834,N_24949,N_24679);
xor U25835 (N_25835,N_24481,N_24978);
nor U25836 (N_25836,N_24460,N_24115);
xnor U25837 (N_25837,N_24304,N_24696);
and U25838 (N_25838,N_24919,N_24872);
or U25839 (N_25839,N_24579,N_24768);
xor U25840 (N_25840,N_24508,N_24021);
xnor U25841 (N_25841,N_24525,N_24561);
nand U25842 (N_25842,N_24405,N_24983);
nor U25843 (N_25843,N_24300,N_24344);
or U25844 (N_25844,N_24627,N_24511);
xnor U25845 (N_25845,N_24682,N_24927);
nor U25846 (N_25846,N_24889,N_24314);
nand U25847 (N_25847,N_24635,N_24251);
nor U25848 (N_25848,N_24705,N_24304);
or U25849 (N_25849,N_24170,N_24251);
or U25850 (N_25850,N_24620,N_24437);
nand U25851 (N_25851,N_24268,N_24665);
or U25852 (N_25852,N_24740,N_24391);
and U25853 (N_25853,N_24965,N_24797);
and U25854 (N_25854,N_24097,N_24170);
nand U25855 (N_25855,N_24173,N_24780);
or U25856 (N_25856,N_24866,N_24653);
and U25857 (N_25857,N_24285,N_24751);
or U25858 (N_25858,N_24875,N_24667);
and U25859 (N_25859,N_24611,N_24896);
and U25860 (N_25860,N_24924,N_24532);
or U25861 (N_25861,N_24683,N_24110);
xor U25862 (N_25862,N_24121,N_24313);
nand U25863 (N_25863,N_24254,N_24631);
nand U25864 (N_25864,N_24715,N_24410);
xnor U25865 (N_25865,N_24654,N_24469);
nand U25866 (N_25866,N_24629,N_24466);
and U25867 (N_25867,N_24773,N_24462);
and U25868 (N_25868,N_24898,N_24059);
nand U25869 (N_25869,N_24064,N_24272);
nor U25870 (N_25870,N_24343,N_24054);
and U25871 (N_25871,N_24189,N_24549);
nand U25872 (N_25872,N_24165,N_24782);
or U25873 (N_25873,N_24452,N_24445);
xor U25874 (N_25874,N_24397,N_24427);
or U25875 (N_25875,N_24524,N_24442);
and U25876 (N_25876,N_24717,N_24590);
nand U25877 (N_25877,N_24658,N_24119);
and U25878 (N_25878,N_24747,N_24460);
and U25879 (N_25879,N_24599,N_24790);
xor U25880 (N_25880,N_24842,N_24060);
nor U25881 (N_25881,N_24353,N_24462);
or U25882 (N_25882,N_24404,N_24538);
xnor U25883 (N_25883,N_24024,N_24743);
nor U25884 (N_25884,N_24028,N_24793);
nor U25885 (N_25885,N_24642,N_24026);
nand U25886 (N_25886,N_24081,N_24078);
nor U25887 (N_25887,N_24757,N_24970);
or U25888 (N_25888,N_24558,N_24009);
and U25889 (N_25889,N_24489,N_24632);
and U25890 (N_25890,N_24989,N_24792);
xor U25891 (N_25891,N_24258,N_24353);
nand U25892 (N_25892,N_24282,N_24880);
nand U25893 (N_25893,N_24866,N_24076);
xnor U25894 (N_25894,N_24880,N_24536);
nand U25895 (N_25895,N_24114,N_24419);
nor U25896 (N_25896,N_24446,N_24790);
nor U25897 (N_25897,N_24684,N_24134);
nand U25898 (N_25898,N_24080,N_24467);
and U25899 (N_25899,N_24649,N_24972);
nor U25900 (N_25900,N_24066,N_24775);
or U25901 (N_25901,N_24080,N_24908);
nand U25902 (N_25902,N_24745,N_24711);
nor U25903 (N_25903,N_24377,N_24730);
nor U25904 (N_25904,N_24330,N_24176);
and U25905 (N_25905,N_24797,N_24002);
or U25906 (N_25906,N_24041,N_24338);
nand U25907 (N_25907,N_24418,N_24118);
and U25908 (N_25908,N_24631,N_24352);
or U25909 (N_25909,N_24690,N_24087);
and U25910 (N_25910,N_24418,N_24676);
or U25911 (N_25911,N_24374,N_24478);
nand U25912 (N_25912,N_24006,N_24005);
or U25913 (N_25913,N_24909,N_24176);
and U25914 (N_25914,N_24371,N_24095);
and U25915 (N_25915,N_24860,N_24724);
nor U25916 (N_25916,N_24788,N_24962);
nor U25917 (N_25917,N_24076,N_24705);
or U25918 (N_25918,N_24793,N_24321);
nor U25919 (N_25919,N_24168,N_24754);
nand U25920 (N_25920,N_24854,N_24007);
nor U25921 (N_25921,N_24630,N_24497);
or U25922 (N_25922,N_24689,N_24792);
xnor U25923 (N_25923,N_24112,N_24369);
nor U25924 (N_25924,N_24736,N_24855);
nand U25925 (N_25925,N_24881,N_24103);
nor U25926 (N_25926,N_24973,N_24372);
and U25927 (N_25927,N_24399,N_24231);
nand U25928 (N_25928,N_24615,N_24059);
nor U25929 (N_25929,N_24027,N_24213);
and U25930 (N_25930,N_24596,N_24576);
or U25931 (N_25931,N_24427,N_24274);
xor U25932 (N_25932,N_24317,N_24070);
and U25933 (N_25933,N_24122,N_24378);
nor U25934 (N_25934,N_24720,N_24965);
nor U25935 (N_25935,N_24691,N_24778);
xor U25936 (N_25936,N_24106,N_24105);
nand U25937 (N_25937,N_24915,N_24295);
or U25938 (N_25938,N_24568,N_24700);
nand U25939 (N_25939,N_24595,N_24241);
nand U25940 (N_25940,N_24249,N_24364);
and U25941 (N_25941,N_24675,N_24411);
nand U25942 (N_25942,N_24064,N_24994);
xor U25943 (N_25943,N_24909,N_24076);
nor U25944 (N_25944,N_24370,N_24321);
or U25945 (N_25945,N_24595,N_24246);
and U25946 (N_25946,N_24626,N_24941);
nor U25947 (N_25947,N_24133,N_24505);
xnor U25948 (N_25948,N_24018,N_24390);
or U25949 (N_25949,N_24224,N_24961);
nor U25950 (N_25950,N_24641,N_24841);
nand U25951 (N_25951,N_24272,N_24855);
nor U25952 (N_25952,N_24924,N_24569);
nand U25953 (N_25953,N_24218,N_24864);
xor U25954 (N_25954,N_24705,N_24216);
nand U25955 (N_25955,N_24402,N_24768);
nand U25956 (N_25956,N_24152,N_24370);
xnor U25957 (N_25957,N_24139,N_24066);
xor U25958 (N_25958,N_24004,N_24954);
xor U25959 (N_25959,N_24681,N_24293);
nand U25960 (N_25960,N_24134,N_24554);
nor U25961 (N_25961,N_24406,N_24164);
xnor U25962 (N_25962,N_24774,N_24360);
and U25963 (N_25963,N_24914,N_24871);
and U25964 (N_25964,N_24176,N_24823);
xnor U25965 (N_25965,N_24131,N_24618);
xor U25966 (N_25966,N_24129,N_24194);
nor U25967 (N_25967,N_24844,N_24119);
and U25968 (N_25968,N_24455,N_24471);
and U25969 (N_25969,N_24686,N_24272);
and U25970 (N_25970,N_24023,N_24322);
xnor U25971 (N_25971,N_24664,N_24484);
nor U25972 (N_25972,N_24815,N_24613);
or U25973 (N_25973,N_24401,N_24356);
and U25974 (N_25974,N_24489,N_24782);
xor U25975 (N_25975,N_24100,N_24744);
and U25976 (N_25976,N_24201,N_24175);
xnor U25977 (N_25977,N_24394,N_24253);
nor U25978 (N_25978,N_24602,N_24549);
and U25979 (N_25979,N_24781,N_24588);
nand U25980 (N_25980,N_24496,N_24152);
xnor U25981 (N_25981,N_24661,N_24713);
nor U25982 (N_25982,N_24195,N_24137);
and U25983 (N_25983,N_24955,N_24273);
nor U25984 (N_25984,N_24321,N_24358);
and U25985 (N_25985,N_24209,N_24843);
or U25986 (N_25986,N_24257,N_24071);
and U25987 (N_25987,N_24355,N_24226);
xor U25988 (N_25988,N_24612,N_24508);
nand U25989 (N_25989,N_24023,N_24470);
and U25990 (N_25990,N_24768,N_24276);
nand U25991 (N_25991,N_24415,N_24111);
xor U25992 (N_25992,N_24787,N_24111);
nor U25993 (N_25993,N_24406,N_24400);
nand U25994 (N_25994,N_24708,N_24641);
nor U25995 (N_25995,N_24236,N_24013);
xnor U25996 (N_25996,N_24169,N_24891);
and U25997 (N_25997,N_24236,N_24168);
or U25998 (N_25998,N_24262,N_24041);
nor U25999 (N_25999,N_24268,N_24833);
nor U26000 (N_26000,N_25520,N_25624);
nor U26001 (N_26001,N_25631,N_25017);
xor U26002 (N_26002,N_25111,N_25584);
or U26003 (N_26003,N_25806,N_25916);
or U26004 (N_26004,N_25507,N_25989);
xor U26005 (N_26005,N_25807,N_25918);
and U26006 (N_26006,N_25604,N_25677);
or U26007 (N_26007,N_25510,N_25766);
or U26008 (N_26008,N_25881,N_25575);
nand U26009 (N_26009,N_25342,N_25725);
and U26010 (N_26010,N_25194,N_25121);
nor U26011 (N_26011,N_25034,N_25508);
nor U26012 (N_26012,N_25910,N_25407);
or U26013 (N_26013,N_25669,N_25934);
and U26014 (N_26014,N_25386,N_25158);
xnor U26015 (N_26015,N_25739,N_25556);
or U26016 (N_26016,N_25526,N_25994);
or U26017 (N_26017,N_25229,N_25853);
or U26018 (N_26018,N_25496,N_25021);
and U26019 (N_26019,N_25044,N_25244);
nand U26020 (N_26020,N_25478,N_25441);
xor U26021 (N_26021,N_25691,N_25950);
or U26022 (N_26022,N_25007,N_25845);
nand U26023 (N_26023,N_25912,N_25268);
or U26024 (N_26024,N_25660,N_25415);
and U26025 (N_26025,N_25540,N_25605);
or U26026 (N_26026,N_25247,N_25871);
or U26027 (N_26027,N_25923,N_25969);
nor U26028 (N_26028,N_25266,N_25642);
nor U26029 (N_26029,N_25444,N_25582);
and U26030 (N_26030,N_25330,N_25637);
nor U26031 (N_26031,N_25080,N_25799);
xnor U26032 (N_26032,N_25919,N_25543);
and U26033 (N_26033,N_25824,N_25302);
and U26034 (N_26034,N_25908,N_25672);
nor U26035 (N_26035,N_25051,N_25841);
nand U26036 (N_26036,N_25494,N_25993);
or U26037 (N_26037,N_25214,N_25428);
and U26038 (N_26038,N_25114,N_25329);
xnor U26039 (N_26039,N_25535,N_25569);
xnor U26040 (N_26040,N_25468,N_25749);
or U26041 (N_26041,N_25418,N_25636);
or U26042 (N_26042,N_25294,N_25399);
and U26043 (N_26043,N_25944,N_25177);
and U26044 (N_26044,N_25692,N_25814);
nor U26045 (N_26045,N_25180,N_25346);
nand U26046 (N_26046,N_25589,N_25829);
xor U26047 (N_26047,N_25992,N_25457);
nand U26048 (N_26048,N_25400,N_25168);
and U26049 (N_26049,N_25967,N_25727);
nor U26050 (N_26050,N_25859,N_25706);
and U26051 (N_26051,N_25865,N_25423);
nor U26052 (N_26052,N_25913,N_25959);
xor U26053 (N_26053,N_25377,N_25723);
nor U26054 (N_26054,N_25708,N_25961);
xnor U26055 (N_26055,N_25554,N_25277);
nand U26056 (N_26056,N_25075,N_25395);
nor U26057 (N_26057,N_25254,N_25664);
nand U26058 (N_26058,N_25225,N_25843);
xnor U26059 (N_26059,N_25008,N_25394);
nand U26060 (N_26060,N_25109,N_25553);
or U26061 (N_26061,N_25092,N_25499);
xnor U26062 (N_26062,N_25138,N_25975);
or U26063 (N_26063,N_25747,N_25634);
nand U26064 (N_26064,N_25403,N_25523);
xnor U26065 (N_26065,N_25943,N_25787);
xor U26066 (N_26066,N_25301,N_25956);
nor U26067 (N_26067,N_25370,N_25223);
and U26068 (N_26068,N_25501,N_25700);
nand U26069 (N_26069,N_25753,N_25729);
and U26070 (N_26070,N_25601,N_25931);
nor U26071 (N_26071,N_25383,N_25470);
or U26072 (N_26072,N_25065,N_25350);
nor U26073 (N_26073,N_25968,N_25057);
xnor U26074 (N_26074,N_25699,N_25161);
or U26075 (N_26075,N_25459,N_25550);
xor U26076 (N_26076,N_25996,N_25612);
xor U26077 (N_26077,N_25037,N_25820);
xnor U26078 (N_26078,N_25658,N_25782);
or U26079 (N_26079,N_25868,N_25489);
or U26080 (N_26080,N_25061,N_25963);
or U26081 (N_26081,N_25292,N_25670);
nand U26082 (N_26082,N_25680,N_25957);
nand U26083 (N_26083,N_25883,N_25497);
xor U26084 (N_26084,N_25711,N_25724);
nand U26085 (N_26085,N_25909,N_25185);
xnor U26086 (N_26086,N_25282,N_25079);
and U26087 (N_26087,N_25863,N_25886);
xnor U26088 (N_26088,N_25907,N_25143);
or U26089 (N_26089,N_25887,N_25182);
nor U26090 (N_26090,N_25434,N_25512);
nor U26091 (N_26091,N_25581,N_25867);
or U26092 (N_26092,N_25381,N_25305);
and U26093 (N_26093,N_25447,N_25222);
xor U26094 (N_26094,N_25189,N_25487);
xor U26095 (N_26095,N_25667,N_25651);
nand U26096 (N_26096,N_25655,N_25014);
xor U26097 (N_26097,N_25564,N_25382);
or U26098 (N_26098,N_25673,N_25524);
xnor U26099 (N_26099,N_25084,N_25378);
or U26100 (N_26100,N_25933,N_25498);
or U26101 (N_26101,N_25476,N_25480);
nand U26102 (N_26102,N_25755,N_25164);
nor U26103 (N_26103,N_25165,N_25684);
xnor U26104 (N_26104,N_25210,N_25942);
and U26105 (N_26105,N_25442,N_25769);
xor U26106 (N_26106,N_25840,N_25774);
xor U26107 (N_26107,N_25253,N_25693);
xnor U26108 (N_26108,N_25484,N_25573);
xor U26109 (N_26109,N_25761,N_25740);
nor U26110 (N_26110,N_25032,N_25701);
nor U26111 (N_26111,N_25215,N_25081);
nor U26112 (N_26112,N_25259,N_25445);
nand U26113 (N_26113,N_25786,N_25615);
xnor U26114 (N_26114,N_25816,N_25297);
and U26115 (N_26115,N_25027,N_25473);
xor U26116 (N_26116,N_25183,N_25107);
nand U26117 (N_26117,N_25152,N_25062);
and U26118 (N_26118,N_25924,N_25241);
or U26119 (N_26119,N_25530,N_25662);
and U26120 (N_26120,N_25326,N_25228);
or U26121 (N_26121,N_25561,N_25101);
nor U26122 (N_26122,N_25074,N_25522);
or U26123 (N_26123,N_25973,N_25439);
nor U26124 (N_26124,N_25393,N_25200);
nor U26125 (N_26125,N_25320,N_25619);
or U26126 (N_26126,N_25683,N_25714);
or U26127 (N_26127,N_25965,N_25617);
nor U26128 (N_26128,N_25201,N_25647);
and U26129 (N_26129,N_25851,N_25610);
nor U26130 (N_26130,N_25469,N_25713);
nand U26131 (N_26131,N_25679,N_25492);
nor U26132 (N_26132,N_25771,N_25269);
and U26133 (N_26133,N_25668,N_25758);
nand U26134 (N_26134,N_25145,N_25698);
nand U26135 (N_26135,N_25308,N_25538);
xnor U26136 (N_26136,N_25426,N_25060);
nand U26137 (N_26137,N_25935,N_25261);
nand U26138 (N_26138,N_25040,N_25646);
nor U26139 (N_26139,N_25757,N_25951);
nand U26140 (N_26140,N_25327,N_25118);
and U26141 (N_26141,N_25379,N_25020);
and U26142 (N_26142,N_25641,N_25456);
or U26143 (N_26143,N_25744,N_25003);
nor U26144 (N_26144,N_25629,N_25517);
and U26145 (N_26145,N_25202,N_25140);
nor U26146 (N_26146,N_25325,N_25271);
and U26147 (N_26147,N_25345,N_25306);
or U26148 (N_26148,N_25056,N_25359);
xnor U26149 (N_26149,N_25162,N_25134);
nor U26150 (N_26150,N_25406,N_25337);
xor U26151 (N_26151,N_25891,N_25255);
or U26152 (N_26152,N_25640,N_25614);
or U26153 (N_26153,N_25167,N_25455);
or U26154 (N_26154,N_25542,N_25050);
nand U26155 (N_26155,N_25022,N_25844);
nor U26156 (N_26156,N_25129,N_25477);
nor U26157 (N_26157,N_25654,N_25388);
and U26158 (N_26158,N_25870,N_25785);
xnor U26159 (N_26159,N_25095,N_25351);
xor U26160 (N_26160,N_25312,N_25800);
and U26161 (N_26161,N_25644,N_25984);
nor U26162 (N_26162,N_25153,N_25733);
nand U26163 (N_26163,N_25756,N_25310);
or U26164 (N_26164,N_25846,N_25450);
nor U26165 (N_26165,N_25882,N_25068);
nor U26166 (N_26166,N_25026,N_25142);
nor U26167 (N_26167,N_25243,N_25300);
nor U26168 (N_26168,N_25879,N_25106);
nand U26169 (N_26169,N_25174,N_25098);
nor U26170 (N_26170,N_25119,N_25097);
nor U26171 (N_26171,N_25227,N_25112);
nor U26172 (N_26172,N_25211,N_25117);
nand U26173 (N_26173,N_25436,N_25169);
nor U26174 (N_26174,N_25380,N_25519);
and U26175 (N_26175,N_25532,N_25921);
nand U26176 (N_26176,N_25052,N_25869);
nand U26177 (N_26177,N_25568,N_25557);
nand U26178 (N_26178,N_25876,N_25071);
nand U26179 (N_26179,N_25043,N_25115);
or U26180 (N_26180,N_25953,N_25001);
or U26181 (N_26181,N_25533,N_25064);
xnor U26182 (N_26182,N_25028,N_25322);
nand U26183 (N_26183,N_25110,N_25465);
nor U26184 (N_26184,N_25945,N_25549);
and U26185 (N_26185,N_25888,N_25331);
or U26186 (N_26186,N_25528,N_25285);
nand U26187 (N_26187,N_25073,N_25938);
and U26188 (N_26188,N_25046,N_25810);
nor U26189 (N_26189,N_25630,N_25263);
nand U26190 (N_26190,N_25541,N_25628);
or U26191 (N_26191,N_25854,N_25726);
xor U26192 (N_26192,N_25276,N_25408);
or U26193 (N_26193,N_25190,N_25390);
nor U26194 (N_26194,N_25884,N_25414);
nand U26195 (N_26195,N_25131,N_25937);
xnor U26196 (N_26196,N_25735,N_25525);
nand U26197 (N_26197,N_25606,N_25094);
or U26198 (N_26198,N_25103,N_25411);
and U26199 (N_26199,N_25077,N_25332);
nand U26200 (N_26200,N_25838,N_25592);
nor U26201 (N_26201,N_25750,N_25796);
or U26202 (N_26202,N_25954,N_25374);
or U26203 (N_26203,N_25917,N_25448);
or U26204 (N_26204,N_25925,N_25777);
nor U26205 (N_26205,N_25939,N_25552);
or U26206 (N_26206,N_25602,N_25260);
xor U26207 (N_26207,N_25705,N_25878);
nand U26208 (N_26208,N_25929,N_25986);
nor U26209 (N_26209,N_25421,N_25754);
nor U26210 (N_26210,N_25410,N_25387);
nor U26211 (N_26211,N_25503,N_25148);
or U26212 (N_26212,N_25175,N_25852);
and U26213 (N_26213,N_25462,N_25633);
xnor U26214 (N_26214,N_25096,N_25621);
or U26215 (N_26215,N_25000,N_25252);
nor U26216 (N_26216,N_25089,N_25318);
and U26217 (N_26217,N_25425,N_25430);
or U26218 (N_26218,N_25139,N_25836);
or U26219 (N_26219,N_25127,N_25941);
nand U26220 (N_26220,N_25927,N_25719);
xnor U26221 (N_26221,N_25220,N_25539);
and U26222 (N_26222,N_25355,N_25193);
or U26223 (N_26223,N_25746,N_25273);
or U26224 (N_26224,N_25828,N_25665);
xnor U26225 (N_26225,N_25588,N_25563);
and U26226 (N_26226,N_25309,N_25005);
nand U26227 (N_26227,N_25690,N_25659);
nor U26228 (N_26228,N_25159,N_25995);
or U26229 (N_26229,N_25289,N_25135);
or U26230 (N_26230,N_25334,N_25583);
nand U26231 (N_26231,N_25548,N_25352);
nand U26232 (N_26232,N_25555,N_25249);
or U26233 (N_26233,N_25120,N_25250);
xor U26234 (N_26234,N_25197,N_25696);
nand U26235 (N_26235,N_25960,N_25695);
xor U26236 (N_26236,N_25980,N_25608);
xnor U26237 (N_26237,N_25454,N_25897);
nand U26238 (N_26238,N_25544,N_25591);
nor U26239 (N_26239,N_25023,N_25343);
xnor U26240 (N_26240,N_25186,N_25398);
nand U26241 (N_26241,N_25347,N_25587);
and U26242 (N_26242,N_25048,N_25815);
xnor U26243 (N_26243,N_25645,N_25835);
or U26244 (N_26244,N_25926,N_25874);
and U26245 (N_26245,N_25805,N_25099);
nor U26246 (N_26246,N_25570,N_25427);
xnor U26247 (N_26247,N_25483,N_25262);
nor U26248 (N_26248,N_25217,N_25781);
or U26249 (N_26249,N_25072,N_25505);
xor U26250 (N_26250,N_25002,N_25504);
nor U26251 (N_26251,N_25546,N_25248);
or U26252 (N_26252,N_25536,N_25904);
xnor U26253 (N_26253,N_25404,N_25371);
or U26254 (N_26254,N_25176,N_25966);
nor U26255 (N_26255,N_25751,N_25237);
or U26256 (N_26256,N_25819,N_25857);
and U26257 (N_26257,N_25146,N_25979);
xor U26258 (N_26258,N_25594,N_25104);
and U26259 (N_26259,N_25981,N_25181);
xnor U26260 (N_26260,N_25978,N_25803);
nor U26261 (N_26261,N_25491,N_25204);
nand U26262 (N_26262,N_25559,N_25206);
and U26263 (N_26263,N_25596,N_25137);
nor U26264 (N_26264,N_25811,N_25607);
and U26265 (N_26265,N_25609,N_25593);
and U26266 (N_26266,N_25316,N_25136);
nand U26267 (N_26267,N_25246,N_25281);
and U26268 (N_26268,N_25042,N_25962);
or U26269 (N_26269,N_25191,N_25715);
and U26270 (N_26270,N_25900,N_25759);
xor U26271 (N_26271,N_25431,N_25336);
nand U26272 (N_26272,N_25770,N_25808);
nor U26273 (N_26273,N_25283,N_25236);
nor U26274 (N_26274,N_25576,N_25652);
nand U26275 (N_26275,N_25147,N_25367);
nand U26276 (N_26276,N_25230,N_25784);
and U26277 (N_26277,N_25982,N_25936);
xor U26278 (N_26278,N_25620,N_25375);
nor U26279 (N_26279,N_25486,N_25817);
or U26280 (N_26280,N_25760,N_25716);
and U26281 (N_26281,N_25417,N_25270);
and U26282 (N_26282,N_25160,N_25710);
and U26283 (N_26283,N_25433,N_25338);
or U26284 (N_26284,N_25625,N_25502);
or U26285 (N_26285,N_25251,N_25313);
xnor U26286 (N_26286,N_25232,N_25558);
nand U26287 (N_26287,N_25964,N_25391);
and U26288 (N_26288,N_25265,N_25412);
nand U26289 (N_26289,N_25616,N_25123);
nor U26290 (N_26290,N_25362,N_25850);
xnor U26291 (N_26291,N_25833,N_25720);
xor U26292 (N_26292,N_25877,N_25173);
nor U26293 (N_26293,N_25264,N_25892);
xor U26294 (N_26294,N_25813,N_25529);
or U26295 (N_26295,N_25019,N_25413);
nor U26296 (N_26296,N_25045,N_25440);
or U26297 (N_26297,N_25323,N_25511);
and U26298 (N_26298,N_25090,N_25901);
or U26299 (N_26299,N_25474,N_25156);
nor U26300 (N_26300,N_25335,N_25358);
nor U26301 (N_26301,N_25049,N_25035);
nand U26302 (N_26302,N_25622,N_25472);
and U26303 (N_26303,N_25847,N_25363);
xor U26304 (N_26304,N_25272,N_25626);
nand U26305 (N_26305,N_25238,N_25578);
nor U26306 (N_26306,N_25066,N_25409);
nor U26307 (N_26307,N_25721,N_25764);
or U26308 (N_26308,N_25794,N_25639);
nand U26309 (N_26309,N_25792,N_25574);
nor U26310 (N_26310,N_25392,N_25566);
nand U26311 (N_26311,N_25765,N_25737);
nor U26312 (N_26312,N_25788,N_25067);
xor U26313 (N_26313,N_25856,N_25464);
nor U26314 (N_26314,N_25718,N_25830);
nand U26315 (N_26315,N_25855,N_25862);
nand U26316 (N_26316,N_25213,N_25467);
xor U26317 (N_26317,N_25036,N_25990);
xnor U26318 (N_26318,N_25366,N_25955);
nand U26319 (N_26319,N_25278,N_25424);
nor U26320 (N_26320,N_25632,N_25722);
and U26321 (N_26321,N_25443,N_25172);
or U26322 (N_26322,N_25087,N_25102);
and U26323 (N_26323,N_25207,N_25743);
and U26324 (N_26324,N_25738,N_25873);
xor U26325 (N_26325,N_25116,N_25258);
or U26326 (N_26326,N_25531,N_25745);
nand U26327 (N_26327,N_25972,N_25493);
and U26328 (N_26328,N_25638,N_25930);
xnor U26329 (N_26329,N_25880,N_25033);
xor U26330 (N_26330,N_25063,N_25130);
xnor U26331 (N_26331,N_25618,N_25623);
or U26332 (N_26332,N_25778,N_25132);
and U26333 (N_26333,N_25681,N_25999);
xnor U26334 (N_26334,N_25889,N_25694);
or U26335 (N_26335,N_25298,N_25154);
xnor U26336 (N_26336,N_25914,N_25178);
nand U26337 (N_26337,N_25653,N_25742);
xnor U26338 (N_26338,N_25333,N_25603);
and U26339 (N_26339,N_25429,N_25970);
nand U26340 (N_26340,N_25795,N_25905);
nor U26341 (N_26341,N_25070,N_25171);
nand U26342 (N_26342,N_25015,N_25082);
nor U26343 (N_26343,N_25842,N_25293);
nand U26344 (N_26344,N_25170,N_25661);
nand U26345 (N_26345,N_25686,N_25196);
and U26346 (N_26346,N_25915,N_25422);
and U26347 (N_26347,N_25419,N_25697);
and U26348 (N_26348,N_25240,N_25288);
nand U26349 (N_26349,N_25012,N_25702);
and U26350 (N_26350,N_25341,N_25985);
nor U26351 (N_26351,N_25775,N_25242);
and U26352 (N_26352,N_25179,N_25416);
nor U26353 (N_26353,N_25898,N_25041);
xor U26354 (N_26354,N_25086,N_25224);
xnor U26355 (N_26355,N_25233,N_25357);
nand U26356 (N_26356,N_25689,N_25038);
nor U26357 (N_26357,N_25078,N_25348);
or U26358 (N_26358,N_25006,N_25976);
nor U26359 (N_26359,N_25577,N_25150);
nand U26360 (N_26360,N_25849,N_25821);
nor U26361 (N_26361,N_25004,N_25198);
nor U26362 (N_26362,N_25812,N_25896);
nor U26363 (N_26363,N_25314,N_25537);
nor U26364 (N_26364,N_25011,N_25703);
nand U26365 (N_26365,N_25598,N_25024);
xnor U26366 (N_26366,N_25518,N_25940);
nand U26367 (N_26367,N_25894,N_25998);
or U26368 (N_26368,N_25091,N_25280);
and U26369 (N_26369,N_25054,N_25364);
or U26370 (N_26370,N_25479,N_25495);
and U26371 (N_26371,N_25946,N_25643);
or U26372 (N_26372,N_25047,N_25991);
xnor U26373 (N_26373,N_25365,N_25802);
and U26374 (N_26374,N_25321,N_25971);
nor U26375 (N_26375,N_25353,N_25789);
and U26376 (N_26376,N_25100,N_25125);
and U26377 (N_26377,N_25122,N_25834);
nor U26378 (N_26378,N_25674,N_25438);
nand U26379 (N_26379,N_25650,N_25069);
and U26380 (N_26380,N_25199,N_25356);
nor U26381 (N_26381,N_25151,N_25219);
and U26382 (N_26382,N_25983,N_25157);
or U26383 (N_26383,N_25590,N_25488);
xnor U26384 (N_26384,N_25205,N_25858);
xnor U26385 (N_26385,N_25823,N_25216);
nor U26386 (N_26386,N_25373,N_25039);
and U26387 (N_26387,N_25822,N_25435);
nand U26388 (N_26388,N_25595,N_25952);
or U26389 (N_26389,N_25466,N_25031);
nor U26390 (N_26390,N_25053,N_25906);
or U26391 (N_26391,N_25932,N_25328);
nand U26392 (N_26392,N_25284,N_25728);
xor U26393 (N_26393,N_25825,N_25762);
and U26394 (N_26394,N_25149,N_25958);
and U26395 (N_26395,N_25565,N_25385);
nand U26396 (N_26396,N_25303,N_25797);
and U26397 (N_26397,N_25837,N_25195);
or U26398 (N_26398,N_25752,N_25093);
or U26399 (N_26399,N_25126,N_25911);
nor U26400 (N_26400,N_25580,N_25687);
nand U26401 (N_26401,N_25453,N_25704);
xnor U26402 (N_26402,N_25029,N_25656);
xor U26403 (N_26403,N_25184,N_25613);
or U26404 (N_26404,N_25389,N_25826);
xnor U26405 (N_26405,N_25267,N_25239);
nand U26406 (N_26406,N_25490,N_25221);
nand U26407 (N_26407,N_25013,N_25562);
nand U26408 (N_26408,N_25304,N_25226);
xnor U26409 (N_26409,N_25083,N_25730);
or U26410 (N_26410,N_25920,N_25475);
nor U26411 (N_26411,N_25988,N_25571);
xor U26412 (N_26412,N_25663,N_25256);
or U26413 (N_26413,N_25875,N_25513);
nand U26414 (N_26414,N_25451,N_25514);
nand U26415 (N_26415,N_25586,N_25809);
and U26416 (N_26416,N_25275,N_25832);
nor U26417 (N_26417,N_25291,N_25369);
nor U26418 (N_26418,N_25903,N_25482);
nand U26419 (N_26419,N_25506,N_25128);
nand U26420 (N_26420,N_25212,N_25257);
nand U26421 (N_26421,N_25009,N_25864);
nand U26422 (N_26422,N_25449,N_25368);
and U26423 (N_26423,N_25567,N_25560);
or U26424 (N_26424,N_25627,N_25360);
xor U26425 (N_26425,N_25839,N_25376);
xnor U26426 (N_26426,N_25748,N_25678);
and U26427 (N_26427,N_25675,N_25349);
xnor U26428 (N_26428,N_25405,N_25732);
and U26429 (N_26429,N_25585,N_25471);
nand U26430 (N_26430,N_25827,N_25773);
nor U26431 (N_26431,N_25245,N_25113);
and U26432 (N_26432,N_25279,N_25798);
and U26433 (N_26433,N_25657,N_25712);
nand U26434 (N_26434,N_25311,N_25287);
nor U26435 (N_26435,N_25676,N_25780);
nand U26436 (N_26436,N_25768,N_25779);
nand U26437 (N_26437,N_25790,N_25763);
nor U26438 (N_26438,N_25804,N_25515);
and U26439 (N_26439,N_25058,N_25319);
or U26440 (N_26440,N_25521,N_25861);
nand U26441 (N_26441,N_25709,N_25974);
or U26442 (N_26442,N_25299,N_25124);
nor U26443 (N_26443,N_25402,N_25648);
xor U26444 (N_26444,N_25509,N_25192);
nand U26445 (N_26445,N_25688,N_25446);
nand U26446 (N_26446,N_25635,N_25384);
and U26447 (N_26447,N_25579,N_25361);
or U26448 (N_26448,N_25317,N_25599);
nor U26449 (N_26449,N_25707,N_25286);
nor U26450 (N_26450,N_25296,N_25324);
nand U26451 (N_26451,N_25059,N_25734);
nor U26452 (N_26452,N_25372,N_25018);
and U26453 (N_26453,N_25500,N_25893);
and U26454 (N_26454,N_25947,N_25534);
nor U26455 (N_26455,N_25307,N_25485);
nor U26456 (N_26456,N_25030,N_25890);
and U26457 (N_26457,N_25987,N_25885);
nor U26458 (N_26458,N_25597,N_25741);
xor U26459 (N_26459,N_25231,N_25866);
and U26460 (N_26460,N_25088,N_25776);
or U26461 (N_26461,N_25831,N_25234);
nand U26462 (N_26462,N_25397,N_25611);
and U26463 (N_26463,N_25600,N_25848);
and U26464 (N_26464,N_25801,N_25458);
xor U26465 (N_26465,N_25108,N_25401);
nor U26466 (N_26466,N_25209,N_25452);
nand U26467 (N_26467,N_25203,N_25977);
nor U26468 (N_26468,N_25463,N_25922);
xor U26469 (N_26469,N_25339,N_25315);
xnor U26470 (N_26470,N_25649,N_25527);
or U26471 (N_26471,N_25144,N_25344);
nand U26472 (N_26472,N_25547,N_25997);
nor U26473 (N_26473,N_25902,N_25791);
nand U26474 (N_26474,N_25895,N_25717);
nor U26475 (N_26475,N_25860,N_25685);
or U26476 (N_26476,N_25460,N_25731);
nor U26477 (N_26477,N_25188,N_25793);
nor U26478 (N_26478,N_25105,N_25572);
nand U26479 (N_26479,N_25461,N_25155);
nor U26480 (N_26480,N_25899,N_25166);
nor U26481 (N_26481,N_25235,N_25736);
nand U26482 (N_26482,N_25290,N_25218);
nand U26483 (N_26483,N_25010,N_25682);
nand U26484 (N_26484,N_25025,N_25948);
nor U26485 (N_26485,N_25872,N_25545);
and U26486 (N_26486,N_25928,N_25671);
nand U26487 (N_26487,N_25772,N_25274);
and U26488 (N_26488,N_25767,N_25340);
and U26489 (N_26489,N_25516,N_25141);
nor U26490 (N_26490,N_25437,N_25949);
xnor U26491 (N_26491,N_25076,N_25666);
and U26492 (N_26492,N_25396,N_25163);
or U26493 (N_26493,N_25783,N_25085);
xor U26494 (N_26494,N_25187,N_25551);
and U26495 (N_26495,N_25295,N_25420);
and U26496 (N_26496,N_25208,N_25055);
and U26497 (N_26497,N_25481,N_25133);
nor U26498 (N_26498,N_25818,N_25016);
or U26499 (N_26499,N_25432,N_25354);
and U26500 (N_26500,N_25151,N_25477);
nand U26501 (N_26501,N_25716,N_25118);
nor U26502 (N_26502,N_25784,N_25736);
or U26503 (N_26503,N_25121,N_25908);
nand U26504 (N_26504,N_25249,N_25673);
or U26505 (N_26505,N_25225,N_25441);
nand U26506 (N_26506,N_25691,N_25086);
or U26507 (N_26507,N_25990,N_25254);
and U26508 (N_26508,N_25123,N_25148);
xor U26509 (N_26509,N_25060,N_25441);
nand U26510 (N_26510,N_25376,N_25503);
xnor U26511 (N_26511,N_25136,N_25841);
xor U26512 (N_26512,N_25872,N_25510);
and U26513 (N_26513,N_25226,N_25845);
or U26514 (N_26514,N_25993,N_25343);
or U26515 (N_26515,N_25646,N_25699);
nand U26516 (N_26516,N_25586,N_25365);
nor U26517 (N_26517,N_25853,N_25962);
xnor U26518 (N_26518,N_25730,N_25637);
or U26519 (N_26519,N_25325,N_25121);
xor U26520 (N_26520,N_25292,N_25069);
nand U26521 (N_26521,N_25919,N_25511);
nor U26522 (N_26522,N_25742,N_25366);
and U26523 (N_26523,N_25401,N_25571);
or U26524 (N_26524,N_25542,N_25658);
nor U26525 (N_26525,N_25799,N_25281);
and U26526 (N_26526,N_25141,N_25558);
xor U26527 (N_26527,N_25395,N_25301);
or U26528 (N_26528,N_25306,N_25617);
xnor U26529 (N_26529,N_25852,N_25919);
xor U26530 (N_26530,N_25541,N_25286);
xor U26531 (N_26531,N_25300,N_25389);
nor U26532 (N_26532,N_25093,N_25646);
and U26533 (N_26533,N_25380,N_25536);
nand U26534 (N_26534,N_25052,N_25925);
nand U26535 (N_26535,N_25264,N_25767);
nor U26536 (N_26536,N_25333,N_25267);
or U26537 (N_26537,N_25009,N_25166);
and U26538 (N_26538,N_25186,N_25739);
and U26539 (N_26539,N_25639,N_25461);
xor U26540 (N_26540,N_25888,N_25459);
xor U26541 (N_26541,N_25118,N_25427);
or U26542 (N_26542,N_25711,N_25371);
nor U26543 (N_26543,N_25102,N_25770);
or U26544 (N_26544,N_25384,N_25948);
xor U26545 (N_26545,N_25553,N_25688);
xor U26546 (N_26546,N_25751,N_25766);
nor U26547 (N_26547,N_25923,N_25094);
xnor U26548 (N_26548,N_25438,N_25503);
or U26549 (N_26549,N_25034,N_25625);
nor U26550 (N_26550,N_25110,N_25995);
and U26551 (N_26551,N_25899,N_25195);
nor U26552 (N_26552,N_25965,N_25019);
and U26553 (N_26553,N_25683,N_25362);
or U26554 (N_26554,N_25828,N_25783);
nand U26555 (N_26555,N_25725,N_25330);
nand U26556 (N_26556,N_25608,N_25574);
and U26557 (N_26557,N_25566,N_25218);
xnor U26558 (N_26558,N_25316,N_25178);
nor U26559 (N_26559,N_25142,N_25350);
or U26560 (N_26560,N_25540,N_25422);
nor U26561 (N_26561,N_25350,N_25770);
xnor U26562 (N_26562,N_25228,N_25405);
xnor U26563 (N_26563,N_25268,N_25644);
nor U26564 (N_26564,N_25069,N_25671);
and U26565 (N_26565,N_25773,N_25297);
nor U26566 (N_26566,N_25164,N_25395);
nor U26567 (N_26567,N_25549,N_25791);
or U26568 (N_26568,N_25284,N_25534);
or U26569 (N_26569,N_25284,N_25410);
nor U26570 (N_26570,N_25109,N_25089);
nand U26571 (N_26571,N_25063,N_25918);
nor U26572 (N_26572,N_25935,N_25780);
nor U26573 (N_26573,N_25075,N_25994);
and U26574 (N_26574,N_25423,N_25275);
or U26575 (N_26575,N_25920,N_25616);
xnor U26576 (N_26576,N_25386,N_25469);
or U26577 (N_26577,N_25073,N_25962);
xor U26578 (N_26578,N_25360,N_25510);
xnor U26579 (N_26579,N_25421,N_25215);
and U26580 (N_26580,N_25161,N_25004);
xor U26581 (N_26581,N_25912,N_25228);
and U26582 (N_26582,N_25411,N_25299);
and U26583 (N_26583,N_25635,N_25097);
or U26584 (N_26584,N_25359,N_25667);
xnor U26585 (N_26585,N_25288,N_25555);
nor U26586 (N_26586,N_25815,N_25143);
and U26587 (N_26587,N_25435,N_25292);
xor U26588 (N_26588,N_25233,N_25579);
or U26589 (N_26589,N_25117,N_25574);
nor U26590 (N_26590,N_25046,N_25383);
xnor U26591 (N_26591,N_25248,N_25227);
nand U26592 (N_26592,N_25876,N_25902);
nand U26593 (N_26593,N_25098,N_25236);
and U26594 (N_26594,N_25661,N_25757);
nand U26595 (N_26595,N_25814,N_25421);
xor U26596 (N_26596,N_25597,N_25212);
nand U26597 (N_26597,N_25334,N_25239);
nand U26598 (N_26598,N_25795,N_25569);
nand U26599 (N_26599,N_25054,N_25959);
nand U26600 (N_26600,N_25735,N_25126);
and U26601 (N_26601,N_25131,N_25126);
nor U26602 (N_26602,N_25617,N_25735);
and U26603 (N_26603,N_25289,N_25130);
xor U26604 (N_26604,N_25156,N_25120);
xor U26605 (N_26605,N_25733,N_25649);
xnor U26606 (N_26606,N_25622,N_25731);
or U26607 (N_26607,N_25783,N_25588);
or U26608 (N_26608,N_25265,N_25507);
nor U26609 (N_26609,N_25757,N_25119);
nor U26610 (N_26610,N_25747,N_25005);
or U26611 (N_26611,N_25974,N_25012);
xor U26612 (N_26612,N_25457,N_25740);
and U26613 (N_26613,N_25253,N_25512);
nor U26614 (N_26614,N_25858,N_25377);
xor U26615 (N_26615,N_25616,N_25188);
nor U26616 (N_26616,N_25139,N_25883);
nand U26617 (N_26617,N_25876,N_25176);
xor U26618 (N_26618,N_25176,N_25688);
xnor U26619 (N_26619,N_25812,N_25874);
xor U26620 (N_26620,N_25230,N_25990);
nor U26621 (N_26621,N_25722,N_25317);
nand U26622 (N_26622,N_25453,N_25139);
xnor U26623 (N_26623,N_25232,N_25113);
nand U26624 (N_26624,N_25601,N_25901);
nor U26625 (N_26625,N_25719,N_25405);
xnor U26626 (N_26626,N_25562,N_25768);
nand U26627 (N_26627,N_25818,N_25634);
and U26628 (N_26628,N_25804,N_25305);
nand U26629 (N_26629,N_25737,N_25263);
nand U26630 (N_26630,N_25431,N_25542);
or U26631 (N_26631,N_25100,N_25987);
nor U26632 (N_26632,N_25216,N_25708);
nand U26633 (N_26633,N_25443,N_25112);
and U26634 (N_26634,N_25326,N_25913);
and U26635 (N_26635,N_25465,N_25488);
and U26636 (N_26636,N_25295,N_25356);
xnor U26637 (N_26637,N_25300,N_25982);
or U26638 (N_26638,N_25042,N_25060);
and U26639 (N_26639,N_25590,N_25752);
and U26640 (N_26640,N_25043,N_25207);
or U26641 (N_26641,N_25355,N_25174);
or U26642 (N_26642,N_25949,N_25166);
xor U26643 (N_26643,N_25641,N_25531);
nand U26644 (N_26644,N_25090,N_25038);
or U26645 (N_26645,N_25120,N_25649);
nor U26646 (N_26646,N_25948,N_25230);
nor U26647 (N_26647,N_25688,N_25674);
and U26648 (N_26648,N_25684,N_25687);
xor U26649 (N_26649,N_25804,N_25546);
and U26650 (N_26650,N_25814,N_25064);
and U26651 (N_26651,N_25990,N_25971);
nor U26652 (N_26652,N_25838,N_25497);
nor U26653 (N_26653,N_25277,N_25952);
nand U26654 (N_26654,N_25754,N_25939);
xnor U26655 (N_26655,N_25752,N_25944);
and U26656 (N_26656,N_25875,N_25015);
nand U26657 (N_26657,N_25575,N_25259);
or U26658 (N_26658,N_25282,N_25872);
nor U26659 (N_26659,N_25157,N_25188);
nor U26660 (N_26660,N_25528,N_25286);
nor U26661 (N_26661,N_25143,N_25635);
and U26662 (N_26662,N_25168,N_25802);
nor U26663 (N_26663,N_25124,N_25506);
or U26664 (N_26664,N_25153,N_25761);
xor U26665 (N_26665,N_25529,N_25631);
nor U26666 (N_26666,N_25638,N_25286);
nor U26667 (N_26667,N_25118,N_25178);
xor U26668 (N_26668,N_25118,N_25171);
nor U26669 (N_26669,N_25600,N_25220);
nand U26670 (N_26670,N_25973,N_25834);
and U26671 (N_26671,N_25027,N_25510);
nand U26672 (N_26672,N_25235,N_25392);
xor U26673 (N_26673,N_25695,N_25739);
xor U26674 (N_26674,N_25291,N_25379);
nor U26675 (N_26675,N_25861,N_25175);
or U26676 (N_26676,N_25593,N_25416);
or U26677 (N_26677,N_25763,N_25499);
xnor U26678 (N_26678,N_25904,N_25446);
or U26679 (N_26679,N_25507,N_25750);
nand U26680 (N_26680,N_25879,N_25375);
xor U26681 (N_26681,N_25558,N_25828);
or U26682 (N_26682,N_25772,N_25365);
nor U26683 (N_26683,N_25454,N_25457);
nand U26684 (N_26684,N_25029,N_25495);
nand U26685 (N_26685,N_25337,N_25209);
and U26686 (N_26686,N_25085,N_25428);
nand U26687 (N_26687,N_25948,N_25177);
or U26688 (N_26688,N_25553,N_25477);
or U26689 (N_26689,N_25657,N_25634);
nand U26690 (N_26690,N_25494,N_25830);
and U26691 (N_26691,N_25270,N_25372);
or U26692 (N_26692,N_25804,N_25234);
nand U26693 (N_26693,N_25657,N_25757);
and U26694 (N_26694,N_25826,N_25374);
xor U26695 (N_26695,N_25599,N_25617);
or U26696 (N_26696,N_25018,N_25404);
or U26697 (N_26697,N_25712,N_25606);
xor U26698 (N_26698,N_25187,N_25295);
or U26699 (N_26699,N_25749,N_25313);
and U26700 (N_26700,N_25188,N_25663);
or U26701 (N_26701,N_25603,N_25141);
nor U26702 (N_26702,N_25173,N_25178);
xor U26703 (N_26703,N_25283,N_25017);
nand U26704 (N_26704,N_25729,N_25329);
nand U26705 (N_26705,N_25324,N_25699);
or U26706 (N_26706,N_25868,N_25124);
or U26707 (N_26707,N_25822,N_25973);
nand U26708 (N_26708,N_25085,N_25616);
and U26709 (N_26709,N_25987,N_25228);
and U26710 (N_26710,N_25924,N_25046);
nand U26711 (N_26711,N_25421,N_25055);
nor U26712 (N_26712,N_25794,N_25121);
or U26713 (N_26713,N_25961,N_25954);
or U26714 (N_26714,N_25425,N_25040);
xnor U26715 (N_26715,N_25022,N_25705);
and U26716 (N_26716,N_25418,N_25802);
nand U26717 (N_26717,N_25159,N_25638);
or U26718 (N_26718,N_25023,N_25342);
xor U26719 (N_26719,N_25802,N_25750);
and U26720 (N_26720,N_25002,N_25578);
xnor U26721 (N_26721,N_25369,N_25822);
or U26722 (N_26722,N_25582,N_25431);
or U26723 (N_26723,N_25372,N_25476);
nor U26724 (N_26724,N_25792,N_25937);
xor U26725 (N_26725,N_25641,N_25848);
or U26726 (N_26726,N_25656,N_25406);
xnor U26727 (N_26727,N_25561,N_25145);
or U26728 (N_26728,N_25154,N_25766);
and U26729 (N_26729,N_25306,N_25007);
nor U26730 (N_26730,N_25597,N_25556);
or U26731 (N_26731,N_25319,N_25881);
or U26732 (N_26732,N_25623,N_25903);
and U26733 (N_26733,N_25922,N_25899);
nor U26734 (N_26734,N_25059,N_25854);
nor U26735 (N_26735,N_25581,N_25520);
or U26736 (N_26736,N_25350,N_25388);
or U26737 (N_26737,N_25707,N_25864);
or U26738 (N_26738,N_25988,N_25684);
nand U26739 (N_26739,N_25135,N_25630);
nor U26740 (N_26740,N_25620,N_25445);
nand U26741 (N_26741,N_25569,N_25589);
and U26742 (N_26742,N_25281,N_25625);
and U26743 (N_26743,N_25938,N_25894);
nor U26744 (N_26744,N_25138,N_25026);
xnor U26745 (N_26745,N_25144,N_25952);
xnor U26746 (N_26746,N_25181,N_25692);
and U26747 (N_26747,N_25342,N_25449);
or U26748 (N_26748,N_25293,N_25434);
nor U26749 (N_26749,N_25455,N_25973);
nor U26750 (N_26750,N_25192,N_25929);
xnor U26751 (N_26751,N_25955,N_25034);
nand U26752 (N_26752,N_25237,N_25732);
nand U26753 (N_26753,N_25924,N_25129);
nand U26754 (N_26754,N_25742,N_25508);
xor U26755 (N_26755,N_25685,N_25927);
nand U26756 (N_26756,N_25672,N_25736);
nand U26757 (N_26757,N_25693,N_25925);
nand U26758 (N_26758,N_25559,N_25476);
and U26759 (N_26759,N_25568,N_25562);
xnor U26760 (N_26760,N_25007,N_25675);
or U26761 (N_26761,N_25129,N_25940);
xor U26762 (N_26762,N_25929,N_25767);
or U26763 (N_26763,N_25807,N_25101);
or U26764 (N_26764,N_25172,N_25771);
or U26765 (N_26765,N_25079,N_25094);
nor U26766 (N_26766,N_25424,N_25515);
xor U26767 (N_26767,N_25059,N_25189);
nand U26768 (N_26768,N_25140,N_25066);
nand U26769 (N_26769,N_25177,N_25212);
xnor U26770 (N_26770,N_25916,N_25121);
nand U26771 (N_26771,N_25833,N_25574);
xor U26772 (N_26772,N_25515,N_25134);
xnor U26773 (N_26773,N_25977,N_25391);
nor U26774 (N_26774,N_25715,N_25799);
or U26775 (N_26775,N_25618,N_25516);
xor U26776 (N_26776,N_25515,N_25429);
and U26777 (N_26777,N_25919,N_25474);
or U26778 (N_26778,N_25327,N_25234);
nor U26779 (N_26779,N_25971,N_25322);
nor U26780 (N_26780,N_25428,N_25952);
or U26781 (N_26781,N_25205,N_25674);
or U26782 (N_26782,N_25827,N_25633);
or U26783 (N_26783,N_25589,N_25877);
nand U26784 (N_26784,N_25857,N_25184);
and U26785 (N_26785,N_25626,N_25729);
nand U26786 (N_26786,N_25201,N_25030);
or U26787 (N_26787,N_25274,N_25333);
and U26788 (N_26788,N_25189,N_25985);
and U26789 (N_26789,N_25405,N_25632);
and U26790 (N_26790,N_25638,N_25062);
xor U26791 (N_26791,N_25488,N_25079);
or U26792 (N_26792,N_25344,N_25059);
or U26793 (N_26793,N_25560,N_25956);
and U26794 (N_26794,N_25377,N_25005);
or U26795 (N_26795,N_25586,N_25372);
and U26796 (N_26796,N_25610,N_25540);
or U26797 (N_26797,N_25125,N_25753);
nand U26798 (N_26798,N_25996,N_25390);
xor U26799 (N_26799,N_25417,N_25723);
xnor U26800 (N_26800,N_25499,N_25108);
or U26801 (N_26801,N_25423,N_25610);
nand U26802 (N_26802,N_25791,N_25686);
or U26803 (N_26803,N_25059,N_25375);
nand U26804 (N_26804,N_25241,N_25739);
xnor U26805 (N_26805,N_25052,N_25098);
and U26806 (N_26806,N_25819,N_25612);
xor U26807 (N_26807,N_25053,N_25904);
xor U26808 (N_26808,N_25566,N_25158);
and U26809 (N_26809,N_25912,N_25201);
or U26810 (N_26810,N_25048,N_25019);
nand U26811 (N_26811,N_25402,N_25484);
nor U26812 (N_26812,N_25970,N_25559);
and U26813 (N_26813,N_25507,N_25446);
or U26814 (N_26814,N_25294,N_25957);
nor U26815 (N_26815,N_25545,N_25975);
and U26816 (N_26816,N_25150,N_25075);
or U26817 (N_26817,N_25264,N_25633);
nand U26818 (N_26818,N_25689,N_25324);
or U26819 (N_26819,N_25231,N_25057);
and U26820 (N_26820,N_25984,N_25254);
and U26821 (N_26821,N_25476,N_25659);
nand U26822 (N_26822,N_25067,N_25156);
nand U26823 (N_26823,N_25069,N_25888);
nand U26824 (N_26824,N_25914,N_25445);
nand U26825 (N_26825,N_25106,N_25417);
nand U26826 (N_26826,N_25946,N_25344);
or U26827 (N_26827,N_25484,N_25013);
xor U26828 (N_26828,N_25007,N_25712);
xor U26829 (N_26829,N_25251,N_25799);
or U26830 (N_26830,N_25051,N_25755);
or U26831 (N_26831,N_25368,N_25289);
xnor U26832 (N_26832,N_25174,N_25520);
nand U26833 (N_26833,N_25139,N_25549);
and U26834 (N_26834,N_25429,N_25731);
nor U26835 (N_26835,N_25533,N_25476);
nand U26836 (N_26836,N_25749,N_25907);
xnor U26837 (N_26837,N_25636,N_25751);
nand U26838 (N_26838,N_25035,N_25067);
or U26839 (N_26839,N_25125,N_25252);
nand U26840 (N_26840,N_25949,N_25001);
xnor U26841 (N_26841,N_25770,N_25233);
xor U26842 (N_26842,N_25356,N_25898);
and U26843 (N_26843,N_25828,N_25943);
nor U26844 (N_26844,N_25456,N_25285);
and U26845 (N_26845,N_25476,N_25812);
xor U26846 (N_26846,N_25400,N_25971);
and U26847 (N_26847,N_25145,N_25183);
nand U26848 (N_26848,N_25195,N_25512);
xnor U26849 (N_26849,N_25888,N_25355);
or U26850 (N_26850,N_25757,N_25522);
and U26851 (N_26851,N_25649,N_25192);
nor U26852 (N_26852,N_25774,N_25161);
and U26853 (N_26853,N_25362,N_25746);
and U26854 (N_26854,N_25008,N_25662);
xnor U26855 (N_26855,N_25181,N_25328);
or U26856 (N_26856,N_25078,N_25977);
or U26857 (N_26857,N_25708,N_25267);
nand U26858 (N_26858,N_25405,N_25291);
xor U26859 (N_26859,N_25473,N_25853);
and U26860 (N_26860,N_25611,N_25362);
or U26861 (N_26861,N_25826,N_25678);
or U26862 (N_26862,N_25374,N_25143);
nand U26863 (N_26863,N_25739,N_25679);
nor U26864 (N_26864,N_25422,N_25995);
nor U26865 (N_26865,N_25742,N_25035);
nor U26866 (N_26866,N_25404,N_25375);
or U26867 (N_26867,N_25006,N_25821);
nor U26868 (N_26868,N_25085,N_25559);
or U26869 (N_26869,N_25177,N_25183);
nand U26870 (N_26870,N_25605,N_25323);
and U26871 (N_26871,N_25397,N_25027);
or U26872 (N_26872,N_25336,N_25914);
or U26873 (N_26873,N_25085,N_25916);
nand U26874 (N_26874,N_25419,N_25676);
and U26875 (N_26875,N_25836,N_25304);
or U26876 (N_26876,N_25761,N_25690);
nor U26877 (N_26877,N_25814,N_25914);
and U26878 (N_26878,N_25846,N_25978);
or U26879 (N_26879,N_25912,N_25348);
and U26880 (N_26880,N_25672,N_25599);
xor U26881 (N_26881,N_25979,N_25753);
nand U26882 (N_26882,N_25135,N_25087);
and U26883 (N_26883,N_25994,N_25638);
and U26884 (N_26884,N_25709,N_25282);
nand U26885 (N_26885,N_25086,N_25562);
xnor U26886 (N_26886,N_25111,N_25460);
xor U26887 (N_26887,N_25117,N_25553);
xor U26888 (N_26888,N_25245,N_25877);
nor U26889 (N_26889,N_25188,N_25382);
or U26890 (N_26890,N_25050,N_25867);
nor U26891 (N_26891,N_25374,N_25872);
nor U26892 (N_26892,N_25150,N_25782);
nor U26893 (N_26893,N_25644,N_25699);
and U26894 (N_26894,N_25298,N_25165);
and U26895 (N_26895,N_25130,N_25284);
and U26896 (N_26896,N_25908,N_25730);
nand U26897 (N_26897,N_25239,N_25773);
or U26898 (N_26898,N_25225,N_25795);
nor U26899 (N_26899,N_25490,N_25774);
and U26900 (N_26900,N_25988,N_25010);
and U26901 (N_26901,N_25164,N_25330);
nand U26902 (N_26902,N_25038,N_25107);
nor U26903 (N_26903,N_25630,N_25002);
nor U26904 (N_26904,N_25561,N_25514);
or U26905 (N_26905,N_25062,N_25004);
xor U26906 (N_26906,N_25432,N_25355);
xor U26907 (N_26907,N_25489,N_25978);
and U26908 (N_26908,N_25959,N_25292);
nand U26909 (N_26909,N_25527,N_25178);
or U26910 (N_26910,N_25537,N_25429);
xor U26911 (N_26911,N_25607,N_25900);
nor U26912 (N_26912,N_25650,N_25693);
nor U26913 (N_26913,N_25964,N_25350);
nor U26914 (N_26914,N_25607,N_25586);
nor U26915 (N_26915,N_25760,N_25182);
nor U26916 (N_26916,N_25061,N_25564);
and U26917 (N_26917,N_25389,N_25904);
nand U26918 (N_26918,N_25505,N_25546);
nand U26919 (N_26919,N_25759,N_25393);
xnor U26920 (N_26920,N_25160,N_25358);
nand U26921 (N_26921,N_25782,N_25052);
and U26922 (N_26922,N_25314,N_25518);
xnor U26923 (N_26923,N_25436,N_25211);
nand U26924 (N_26924,N_25086,N_25823);
nand U26925 (N_26925,N_25428,N_25386);
or U26926 (N_26926,N_25477,N_25542);
nor U26927 (N_26927,N_25225,N_25584);
or U26928 (N_26928,N_25655,N_25567);
nand U26929 (N_26929,N_25820,N_25985);
and U26930 (N_26930,N_25907,N_25978);
nor U26931 (N_26931,N_25499,N_25232);
xor U26932 (N_26932,N_25647,N_25374);
or U26933 (N_26933,N_25004,N_25504);
nor U26934 (N_26934,N_25837,N_25566);
nand U26935 (N_26935,N_25429,N_25392);
nand U26936 (N_26936,N_25699,N_25187);
or U26937 (N_26937,N_25135,N_25440);
xnor U26938 (N_26938,N_25189,N_25407);
or U26939 (N_26939,N_25681,N_25374);
and U26940 (N_26940,N_25053,N_25892);
and U26941 (N_26941,N_25998,N_25370);
or U26942 (N_26942,N_25550,N_25712);
or U26943 (N_26943,N_25865,N_25712);
or U26944 (N_26944,N_25972,N_25118);
and U26945 (N_26945,N_25846,N_25541);
nand U26946 (N_26946,N_25025,N_25606);
nor U26947 (N_26947,N_25701,N_25130);
and U26948 (N_26948,N_25165,N_25755);
xnor U26949 (N_26949,N_25767,N_25119);
nor U26950 (N_26950,N_25065,N_25640);
or U26951 (N_26951,N_25364,N_25351);
xnor U26952 (N_26952,N_25701,N_25915);
nand U26953 (N_26953,N_25152,N_25656);
or U26954 (N_26954,N_25381,N_25349);
or U26955 (N_26955,N_25024,N_25950);
or U26956 (N_26956,N_25955,N_25838);
nor U26957 (N_26957,N_25700,N_25945);
xnor U26958 (N_26958,N_25113,N_25590);
or U26959 (N_26959,N_25007,N_25366);
and U26960 (N_26960,N_25725,N_25466);
and U26961 (N_26961,N_25699,N_25475);
xnor U26962 (N_26962,N_25726,N_25394);
xnor U26963 (N_26963,N_25440,N_25976);
xor U26964 (N_26964,N_25435,N_25007);
and U26965 (N_26965,N_25422,N_25453);
nor U26966 (N_26966,N_25253,N_25110);
and U26967 (N_26967,N_25296,N_25325);
nand U26968 (N_26968,N_25813,N_25500);
nand U26969 (N_26969,N_25181,N_25188);
and U26970 (N_26970,N_25395,N_25104);
and U26971 (N_26971,N_25203,N_25599);
xnor U26972 (N_26972,N_25297,N_25621);
or U26973 (N_26973,N_25448,N_25440);
and U26974 (N_26974,N_25299,N_25321);
and U26975 (N_26975,N_25675,N_25580);
nand U26976 (N_26976,N_25235,N_25410);
and U26977 (N_26977,N_25052,N_25787);
xnor U26978 (N_26978,N_25398,N_25295);
nand U26979 (N_26979,N_25214,N_25345);
nand U26980 (N_26980,N_25142,N_25448);
or U26981 (N_26981,N_25432,N_25701);
or U26982 (N_26982,N_25162,N_25852);
xor U26983 (N_26983,N_25060,N_25094);
nand U26984 (N_26984,N_25764,N_25889);
and U26985 (N_26985,N_25364,N_25013);
and U26986 (N_26986,N_25666,N_25540);
xor U26987 (N_26987,N_25368,N_25187);
nand U26988 (N_26988,N_25588,N_25513);
or U26989 (N_26989,N_25242,N_25927);
xnor U26990 (N_26990,N_25384,N_25017);
xnor U26991 (N_26991,N_25582,N_25191);
nand U26992 (N_26992,N_25708,N_25530);
nor U26993 (N_26993,N_25496,N_25282);
or U26994 (N_26994,N_25522,N_25157);
or U26995 (N_26995,N_25455,N_25650);
or U26996 (N_26996,N_25685,N_25455);
nand U26997 (N_26997,N_25627,N_25327);
nand U26998 (N_26998,N_25316,N_25674);
and U26999 (N_26999,N_25364,N_25790);
or U27000 (N_27000,N_26761,N_26569);
nor U27001 (N_27001,N_26530,N_26263);
nor U27002 (N_27002,N_26164,N_26995);
xor U27003 (N_27003,N_26946,N_26933);
or U27004 (N_27004,N_26275,N_26089);
nor U27005 (N_27005,N_26235,N_26757);
and U27006 (N_27006,N_26481,N_26850);
nor U27007 (N_27007,N_26607,N_26445);
or U27008 (N_27008,N_26811,N_26448);
xnor U27009 (N_27009,N_26870,N_26450);
and U27010 (N_27010,N_26921,N_26495);
and U27011 (N_27011,N_26456,N_26666);
nor U27012 (N_27012,N_26286,N_26825);
nand U27013 (N_27013,N_26401,N_26985);
and U27014 (N_27014,N_26233,N_26515);
or U27015 (N_27015,N_26041,N_26628);
or U27016 (N_27016,N_26693,N_26932);
xnor U27017 (N_27017,N_26767,N_26517);
xnor U27018 (N_27018,N_26649,N_26028);
xnor U27019 (N_27019,N_26637,N_26103);
nand U27020 (N_27020,N_26679,N_26443);
nor U27021 (N_27021,N_26846,N_26192);
and U27022 (N_27022,N_26625,N_26620);
nand U27023 (N_27023,N_26437,N_26650);
xor U27024 (N_27024,N_26913,N_26380);
xnor U27025 (N_27025,N_26480,N_26189);
nor U27026 (N_27026,N_26409,N_26144);
nor U27027 (N_27027,N_26796,N_26229);
nand U27028 (N_27028,N_26542,N_26922);
nand U27029 (N_27029,N_26467,N_26877);
xor U27030 (N_27030,N_26728,N_26357);
or U27031 (N_27031,N_26312,N_26708);
xnor U27032 (N_27032,N_26266,N_26543);
and U27033 (N_27033,N_26347,N_26828);
nand U27034 (N_27034,N_26786,N_26826);
nor U27035 (N_27035,N_26176,N_26115);
nand U27036 (N_27036,N_26213,N_26011);
or U27037 (N_27037,N_26285,N_26865);
xnor U27038 (N_27038,N_26948,N_26411);
nor U27039 (N_27039,N_26433,N_26474);
nand U27040 (N_27040,N_26020,N_26158);
nor U27041 (N_27041,N_26425,N_26241);
nand U27042 (N_27042,N_26676,N_26686);
or U27043 (N_27043,N_26001,N_26440);
nor U27044 (N_27044,N_26141,N_26402);
nand U27045 (N_27045,N_26238,N_26697);
or U27046 (N_27046,N_26912,N_26598);
nor U27047 (N_27047,N_26048,N_26505);
and U27048 (N_27048,N_26050,N_26071);
nor U27049 (N_27049,N_26717,N_26981);
xnor U27050 (N_27050,N_26799,N_26122);
nand U27051 (N_27051,N_26837,N_26379);
xor U27052 (N_27052,N_26352,N_26499);
xnor U27053 (N_27053,N_26582,N_26430);
nand U27054 (N_27054,N_26835,N_26484);
nor U27055 (N_27055,N_26138,N_26733);
and U27056 (N_27056,N_26868,N_26952);
xnor U27057 (N_27057,N_26120,N_26814);
xnor U27058 (N_27058,N_26427,N_26310);
nor U27059 (N_27059,N_26876,N_26389);
or U27060 (N_27060,N_26586,N_26337);
nand U27061 (N_27061,N_26565,N_26217);
xnor U27062 (N_27062,N_26082,N_26604);
nor U27063 (N_27063,N_26738,N_26461);
nand U27064 (N_27064,N_26602,N_26810);
and U27065 (N_27065,N_26252,N_26834);
nand U27066 (N_27066,N_26118,N_26124);
nand U27067 (N_27067,N_26688,N_26070);
or U27068 (N_27068,N_26507,N_26764);
nand U27069 (N_27069,N_26655,N_26462);
and U27070 (N_27070,N_26299,N_26571);
and U27071 (N_27071,N_26540,N_26851);
nor U27072 (N_27072,N_26955,N_26648);
nand U27073 (N_27073,N_26642,N_26917);
or U27074 (N_27074,N_26501,N_26829);
xnor U27075 (N_27075,N_26559,N_26858);
or U27076 (N_27076,N_26174,N_26493);
nand U27077 (N_27077,N_26359,N_26691);
nand U27078 (N_27078,N_26790,N_26705);
nand U27079 (N_27079,N_26202,N_26095);
nor U27080 (N_27080,N_26532,N_26351);
nor U27081 (N_27081,N_26477,N_26662);
or U27082 (N_27082,N_26135,N_26794);
or U27083 (N_27083,N_26998,N_26378);
xor U27084 (N_27084,N_26335,N_26634);
nand U27085 (N_27085,N_26110,N_26168);
nand U27086 (N_27086,N_26342,N_26781);
nor U27087 (N_27087,N_26550,N_26004);
or U27088 (N_27088,N_26316,N_26538);
nand U27089 (N_27089,N_26191,N_26570);
and U27090 (N_27090,N_26581,N_26249);
and U27091 (N_27091,N_26804,N_26240);
xor U27092 (N_27092,N_26894,N_26371);
or U27093 (N_27093,N_26326,N_26419);
or U27094 (N_27094,N_26911,N_26633);
nor U27095 (N_27095,N_26300,N_26105);
or U27096 (N_27096,N_26372,N_26257);
nor U27097 (N_27097,N_26522,N_26606);
and U27098 (N_27098,N_26857,N_26377);
xnor U27099 (N_27099,N_26546,N_26303);
and U27100 (N_27100,N_26151,N_26157);
nor U27101 (N_27101,N_26088,N_26974);
xnor U27102 (N_27102,N_26340,N_26483);
xnor U27103 (N_27103,N_26646,N_26621);
nand U27104 (N_27104,N_26801,N_26265);
nand U27105 (N_27105,N_26816,N_26127);
nand U27106 (N_27106,N_26111,N_26042);
nor U27107 (N_27107,N_26701,N_26924);
and U27108 (N_27108,N_26227,N_26119);
and U27109 (N_27109,N_26594,N_26769);
nor U27110 (N_27110,N_26306,N_26329);
xor U27111 (N_27111,N_26636,N_26962);
and U27112 (N_27112,N_26798,N_26317);
xor U27113 (N_27113,N_26668,N_26319);
nand U27114 (N_27114,N_26595,N_26830);
and U27115 (N_27115,N_26023,N_26181);
and U27116 (N_27116,N_26086,N_26866);
or U27117 (N_27117,N_26274,N_26803);
nand U27118 (N_27118,N_26114,N_26576);
and U27119 (N_27119,N_26725,N_26381);
nand U27120 (N_27120,N_26096,N_26920);
or U27121 (N_27121,N_26729,N_26490);
nor U27122 (N_27122,N_26018,N_26087);
and U27123 (N_27123,N_26287,N_26321);
nor U27124 (N_27124,N_26514,N_26072);
nand U27125 (N_27125,N_26815,N_26945);
nor U27126 (N_27126,N_26328,N_26188);
nor U27127 (N_27127,N_26787,N_26314);
nor U27128 (N_27128,N_26556,N_26972);
nand U27129 (N_27129,N_26752,N_26564);
nand U27130 (N_27130,N_26510,N_26612);
nor U27131 (N_27131,N_26553,N_26195);
xnor U27132 (N_27132,N_26979,N_26671);
xor U27133 (N_27133,N_26605,N_26073);
nor U27134 (N_27134,N_26751,N_26957);
or U27135 (N_27135,N_26627,N_26619);
nand U27136 (N_27136,N_26583,N_26529);
nand U27137 (N_27137,N_26234,N_26388);
and U27138 (N_27138,N_26785,N_26364);
nor U27139 (N_27139,N_26873,N_26898);
and U27140 (N_27140,N_26879,N_26054);
nand U27141 (N_27141,N_26267,N_26052);
xor U27142 (N_27142,N_26682,N_26953);
nand U27143 (N_27143,N_26147,N_26035);
and U27144 (N_27144,N_26201,N_26549);
or U27145 (N_27145,N_26083,N_26079);
xor U27146 (N_27146,N_26236,N_26534);
or U27147 (N_27147,N_26899,N_26021);
nand U27148 (N_27148,N_26256,N_26003);
xor U27149 (N_27149,N_26369,N_26029);
nand U27150 (N_27150,N_26470,N_26283);
nand U27151 (N_27151,N_26040,N_26533);
or U27152 (N_27152,N_26843,N_26797);
xnor U27153 (N_27153,N_26117,N_26768);
nor U27154 (N_27154,N_26373,N_26131);
or U27155 (N_27155,N_26297,N_26719);
and U27156 (N_27156,N_26163,N_26006);
and U27157 (N_27157,N_26750,N_26696);
and U27158 (N_27158,N_26745,N_26394);
nor U27159 (N_27159,N_26491,N_26415);
and U27160 (N_27160,N_26931,N_26155);
or U27161 (N_27161,N_26434,N_26929);
xnor U27162 (N_27162,N_26338,N_26390);
and U27163 (N_27163,N_26414,N_26116);
or U27164 (N_27164,N_26432,N_26665);
and U27165 (N_27165,N_26882,N_26961);
and U27166 (N_27166,N_26944,N_26245);
and U27167 (N_27167,N_26090,N_26988);
nor U27168 (N_27168,N_26022,N_26853);
and U27169 (N_27169,N_26396,N_26459);
and U27170 (N_27170,N_26254,N_26413);
xnor U27171 (N_27171,N_26458,N_26383);
xnor U27172 (N_27172,N_26792,N_26673);
nand U27173 (N_27173,N_26685,N_26647);
nor U27174 (N_27174,N_26889,N_26775);
nand U27175 (N_27175,N_26061,N_26271);
xor U27176 (N_27176,N_26892,N_26473);
nand U27177 (N_27177,N_26171,N_26183);
or U27178 (N_27178,N_26503,N_26942);
nand U27179 (N_27179,N_26108,N_26428);
or U27180 (N_27180,N_26143,N_26154);
and U27181 (N_27181,N_26034,N_26126);
or U27182 (N_27182,N_26991,N_26575);
or U27183 (N_27183,N_26353,N_26017);
nand U27184 (N_27184,N_26856,N_26968);
nand U27185 (N_27185,N_26938,N_26327);
nand U27186 (N_27186,N_26551,N_26601);
nor U27187 (N_27187,N_26259,N_26626);
xnor U27188 (N_27188,N_26807,N_26983);
and U27189 (N_27189,N_26743,N_26165);
xor U27190 (N_27190,N_26354,N_26291);
nor U27191 (N_27191,N_26282,N_26502);
nand U27192 (N_27192,N_26949,N_26078);
and U27193 (N_27193,N_26162,N_26094);
and U27194 (N_27194,N_26221,N_26793);
or U27195 (N_27195,N_26439,N_26186);
nor U27196 (N_27196,N_26196,N_26320);
xnor U27197 (N_27197,N_26718,N_26289);
xor U27198 (N_27198,N_26260,N_26992);
nand U27199 (N_27199,N_26404,N_26466);
nand U27200 (N_27200,N_26180,N_26926);
or U27201 (N_27201,N_26080,N_26224);
or U27202 (N_27202,N_26230,N_26005);
xor U27203 (N_27203,N_26486,N_26527);
nand U27204 (N_27204,N_26426,N_26129);
xnor U27205 (N_27205,N_26896,N_26277);
or U27206 (N_27206,N_26914,N_26190);
xor U27207 (N_27207,N_26216,N_26406);
or U27208 (N_27208,N_26927,N_26805);
nor U27209 (N_27209,N_26101,N_26706);
nor U27210 (N_27210,N_26600,N_26410);
or U27211 (N_27211,N_26045,N_26008);
nor U27212 (N_27212,N_26167,N_26204);
or U27213 (N_27213,N_26239,N_26698);
or U27214 (N_27214,N_26778,N_26641);
and U27215 (N_27215,N_26208,N_26547);
xnor U27216 (N_27216,N_26468,N_26187);
or U27217 (N_27217,N_26199,N_26077);
nand U27218 (N_27218,N_26024,N_26496);
and U27219 (N_27219,N_26791,N_26178);
or U27220 (N_27220,N_26109,N_26137);
and U27221 (N_27221,N_26272,N_26941);
nand U27222 (N_27222,N_26513,N_26046);
and U27223 (N_27223,N_26893,N_26971);
nand U27224 (N_27224,N_26152,N_26362);
nor U27225 (N_27225,N_26611,N_26871);
xor U27226 (N_27226,N_26471,N_26446);
or U27227 (N_27227,N_26910,N_26007);
and U27228 (N_27228,N_26614,N_26984);
and U27229 (N_27229,N_26997,N_26656);
and U27230 (N_27230,N_26016,N_26153);
nor U27231 (N_27231,N_26408,N_26169);
and U27232 (N_27232,N_26521,N_26457);
nand U27233 (N_27233,N_26897,N_26242);
or U27234 (N_27234,N_26497,N_26156);
or U27235 (N_27235,N_26640,N_26066);
and U27236 (N_27236,N_26301,N_26715);
and U27237 (N_27237,N_26305,N_26387);
and U27238 (N_27238,N_26469,N_26964);
nor U27239 (N_27239,N_26043,N_26742);
nor U27240 (N_27240,N_26777,N_26906);
xor U27241 (N_27241,N_26068,N_26731);
and U27242 (N_27242,N_26032,N_26250);
nand U27243 (N_27243,N_26085,N_26753);
or U27244 (N_27244,N_26215,N_26436);
and U27245 (N_27245,N_26667,N_26093);
and U27246 (N_27246,N_26142,N_26528);
nor U27247 (N_27247,N_26999,N_26059);
or U27248 (N_27248,N_26392,N_26782);
and U27249 (N_27249,N_26711,N_26345);
xnor U27250 (N_27250,N_26652,N_26121);
or U27251 (N_27251,N_26883,N_26772);
and U27252 (N_27252,N_26919,N_26677);
xnor U27253 (N_27253,N_26504,N_26603);
and U27254 (N_27254,N_26617,N_26632);
and U27255 (N_27255,N_26887,N_26276);
or U27256 (N_27256,N_26511,N_26759);
or U27257 (N_27257,N_26726,N_26592);
and U27258 (N_27258,N_26322,N_26076);
and U27259 (N_27259,N_26700,N_26488);
nor U27260 (N_27260,N_26566,N_26916);
nand U27261 (N_27261,N_26280,N_26128);
or U27262 (N_27262,N_26736,N_26537);
nor U27263 (N_27263,N_26780,N_26248);
xor U27264 (N_27264,N_26523,N_26884);
and U27265 (N_27265,N_26855,N_26506);
and U27266 (N_27266,N_26279,N_26500);
and U27267 (N_27267,N_26139,N_26047);
and U27268 (N_27268,N_26175,N_26293);
nand U27269 (N_27269,N_26989,N_26049);
nand U27270 (N_27270,N_26261,N_26675);
nor U27271 (N_27271,N_26935,N_26026);
nor U27272 (N_27272,N_26722,N_26455);
and U27273 (N_27273,N_26584,N_26019);
and U27274 (N_27274,N_26993,N_26395);
xnor U27275 (N_27275,N_26994,N_26770);
and U27276 (N_27276,N_26758,N_26444);
xor U27277 (N_27277,N_26747,N_26374);
and U27278 (N_27278,N_26901,N_26037);
nor U27279 (N_27279,N_26431,N_26000);
nand U27280 (N_27280,N_26453,N_26194);
or U27281 (N_27281,N_26177,N_26756);
or U27282 (N_27282,N_26292,N_26464);
nand U27283 (N_27283,N_26862,N_26908);
xor U27284 (N_27284,N_26541,N_26773);
nor U27285 (N_27285,N_26653,N_26909);
or U27286 (N_27286,N_26694,N_26051);
xnor U27287 (N_27287,N_26343,N_26845);
or U27288 (N_27288,N_26552,N_26572);
or U27289 (N_27289,N_26025,N_26623);
or U27290 (N_27290,N_26064,N_26476);
and U27291 (N_27291,N_26687,N_26881);
or U27292 (N_27292,N_26568,N_26067);
nor U27293 (N_27293,N_26978,N_26746);
nand U27294 (N_27294,N_26014,N_26664);
and U27295 (N_27295,N_26727,N_26358);
and U27296 (N_27296,N_26635,N_26324);
xor U27297 (N_27297,N_26900,N_26813);
or U27298 (N_27298,N_26661,N_26442);
nand U27299 (N_27299,N_26982,N_26721);
or U27300 (N_27300,N_26423,N_26062);
and U27301 (N_27301,N_26819,N_26251);
or U27302 (N_27302,N_26593,N_26193);
xor U27303 (N_27303,N_26692,N_26934);
xor U27304 (N_27304,N_26098,N_26332);
or U27305 (N_27305,N_26384,N_26382);
xnor U27306 (N_27306,N_26561,N_26222);
nand U27307 (N_27307,N_26678,N_26060);
nor U27308 (N_27308,N_26860,N_26295);
or U27309 (N_27309,N_26789,N_26822);
nor U27310 (N_27310,N_26184,N_26112);
xnor U27311 (N_27311,N_26107,N_26424);
xnor U27312 (N_27312,N_26220,N_26516);
nand U27313 (N_27313,N_26330,N_26363);
and U27314 (N_27314,N_26478,N_26015);
xnor U27315 (N_27315,N_26106,N_26832);
nand U27316 (N_27316,N_26563,N_26827);
and U27317 (N_27317,N_26928,N_26346);
and U27318 (N_27318,N_26859,N_26278);
xor U27319 (N_27319,N_26302,N_26148);
and U27320 (N_27320,N_26247,N_26589);
and U27321 (N_27321,N_26925,N_26638);
or U27322 (N_27322,N_26441,N_26760);
xnor U27323 (N_27323,N_26038,N_26902);
and U27324 (N_27324,N_26056,N_26714);
nand U27325 (N_27325,N_26954,N_26097);
and U27326 (N_27326,N_26730,N_26878);
nor U27327 (N_27327,N_26710,N_26657);
and U27328 (N_27328,N_26965,N_26318);
and U27329 (N_27329,N_26036,N_26699);
or U27330 (N_27330,N_26132,N_26783);
xor U27331 (N_27331,N_26735,N_26573);
nor U27332 (N_27332,N_26539,N_26818);
nand U27333 (N_27333,N_26861,N_26724);
nor U27334 (N_27334,N_26134,N_26416);
or U27335 (N_27335,N_26027,N_26058);
xor U27336 (N_27336,N_26203,N_26092);
and U27337 (N_27337,N_26872,N_26947);
and U27338 (N_27338,N_26099,N_26739);
nor U27339 (N_27339,N_26460,N_26209);
and U27340 (N_27340,N_26986,N_26885);
xor U27341 (N_27341,N_26683,N_26226);
nand U27342 (N_27342,N_26223,N_26231);
xor U27343 (N_27343,N_26802,N_26960);
nand U27344 (N_27344,N_26421,N_26702);
xnor U27345 (N_27345,N_26307,N_26173);
nand U27346 (N_27346,N_26405,N_26323);
and U27347 (N_27347,N_26225,N_26065);
and U27348 (N_27348,N_26831,N_26057);
nor U27349 (N_27349,N_26429,N_26562);
xor U27350 (N_27350,N_26304,N_26309);
nand U27351 (N_27351,N_26741,N_26639);
or U27352 (N_27352,N_26918,N_26366);
nand U27353 (N_27353,N_26578,N_26557);
nand U27354 (N_27354,N_26074,N_26334);
nor U27355 (N_27355,N_26723,N_26774);
and U27356 (N_27356,N_26800,N_26417);
nand U27357 (N_27357,N_26704,N_26170);
or U27358 (N_27358,N_26766,N_26498);
or U27359 (N_27359,N_26585,N_26763);
nor U27360 (N_27360,N_26211,N_26084);
nand U27361 (N_27361,N_26579,N_26244);
nor U27362 (N_27362,N_26264,N_26400);
xor U27363 (N_27363,N_26618,N_26608);
or U27364 (N_27364,N_26849,N_26689);
or U27365 (N_27365,N_26494,N_26597);
or U27366 (N_27366,N_26133,N_26841);
nor U27367 (N_27367,N_26670,N_26232);
xor U27368 (N_27368,N_26273,N_26755);
or U27369 (N_27369,N_26355,N_26438);
or U27370 (N_27370,N_26643,N_26385);
nor U27371 (N_27371,N_26654,N_26361);
or U27372 (N_27372,N_26875,N_26218);
nand U27373 (N_27373,N_26149,N_26482);
nand U27374 (N_27374,N_26590,N_26923);
or U27375 (N_27375,N_26588,N_26397);
or U27376 (N_27376,N_26709,N_26281);
xnor U27377 (N_27377,N_26560,N_26969);
and U27378 (N_27378,N_26681,N_26644);
xnor U27379 (N_27379,N_26610,N_26904);
nand U27380 (N_27380,N_26658,N_26130);
xnor U27381 (N_27381,N_26616,N_26869);
nor U27382 (N_27382,N_26418,N_26145);
nand U27383 (N_27383,N_26210,N_26350);
nor U27384 (N_27384,N_26903,N_26852);
xor U27385 (N_27385,N_26663,N_26412);
nor U27386 (N_27386,N_26890,N_26707);
nand U27387 (N_27387,N_26548,N_26713);
and U27388 (N_27388,N_26959,N_26847);
xnor U27389 (N_27389,N_26631,N_26228);
nor U27390 (N_27390,N_26246,N_26262);
nor U27391 (N_27391,N_26940,N_26449);
nand U27392 (N_27392,N_26740,N_26895);
or U27393 (N_27393,N_26368,N_26255);
or U27394 (N_27394,N_26207,N_26874);
and U27395 (N_27395,N_26863,N_26013);
nor U27396 (N_27396,N_26009,N_26905);
and U27397 (N_27397,N_26967,N_26508);
nor U27398 (N_27398,N_26950,N_26339);
nand U27399 (N_27399,N_26545,N_26298);
or U27400 (N_27400,N_26206,N_26422);
nor U27401 (N_27401,N_26996,N_26720);
nand U27402 (N_27402,N_26356,N_26844);
or U27403 (N_27403,N_26613,N_26958);
and U27404 (N_27404,N_26447,N_26839);
nor U27405 (N_27405,N_26288,N_26712);
nor U27406 (N_27406,N_26732,N_26672);
or U27407 (N_27407,N_26182,N_26587);
xor U27408 (N_27408,N_26348,N_26010);
nor U27409 (N_27409,N_26771,N_26341);
or U27410 (N_27410,N_26669,N_26465);
xnor U27411 (N_27411,N_26596,N_26659);
nor U27412 (N_27412,N_26817,N_26290);
nand U27413 (N_27413,N_26536,N_26237);
or U27414 (N_27414,N_26012,N_26102);
and U27415 (N_27415,N_26867,N_26651);
nand U27416 (N_27416,N_26970,N_26526);
nor U27417 (N_27417,N_26930,N_26313);
xor U27418 (N_27418,N_26939,N_26308);
and U27419 (N_27419,N_26113,N_26990);
and U27420 (N_27420,N_26053,N_26146);
xnor U27421 (N_27421,N_26376,N_26716);
nand U27422 (N_27422,N_26956,N_26044);
nand U27423 (N_27423,N_26033,N_26809);
or U27424 (N_27424,N_26331,N_26104);
nor U27425 (N_27425,N_26973,N_26531);
nand U27426 (N_27426,N_26762,N_26645);
nand U27427 (N_27427,N_26512,N_26848);
or U27428 (N_27428,N_26684,N_26269);
or U27429 (N_27429,N_26936,N_26479);
nand U27430 (N_27430,N_26943,N_26407);
or U27431 (N_27431,N_26695,N_26375);
or U27432 (N_27432,N_26140,N_26391);
nand U27433 (N_27433,N_26325,N_26591);
and U27434 (N_27434,N_26349,N_26172);
and U27435 (N_27435,N_26823,N_26365);
nand U27436 (N_27436,N_26489,N_26567);
nand U27437 (N_27437,N_26420,N_26580);
nor U27438 (N_27438,N_26854,N_26069);
or U27439 (N_27439,N_26951,N_26891);
xnor U27440 (N_27440,N_26100,N_26836);
or U27441 (N_27441,N_26205,N_26744);
nor U27442 (N_27442,N_26975,N_26002);
nor U27443 (N_27443,N_26136,N_26393);
xor U27444 (N_27444,N_26398,N_26386);
nand U27445 (N_27445,N_26179,N_26734);
nand U27446 (N_27446,N_26435,N_26344);
xnor U27447 (N_27447,N_26161,N_26840);
nand U27448 (N_27448,N_26197,N_26629);
xor U27449 (N_27449,N_26824,N_26243);
and U27450 (N_27450,N_26452,N_26150);
and U27451 (N_27451,N_26976,N_26185);
and U27452 (N_27452,N_26808,N_26518);
or U27453 (N_27453,N_26660,N_26091);
xnor U27454 (N_27454,N_26748,N_26031);
or U27455 (N_27455,N_26125,N_26599);
nor U27456 (N_27456,N_26160,N_26544);
xor U27457 (N_27457,N_26367,N_26333);
or U27458 (N_27458,N_26915,N_26524);
nor U27459 (N_27459,N_26788,N_26485);
and U27460 (N_27460,N_26399,N_26888);
and U27461 (N_27461,N_26680,N_26159);
or U27462 (N_27462,N_26055,N_26907);
nor U27463 (N_27463,N_26624,N_26370);
and U27464 (N_27464,N_26838,N_26284);
xnor U27465 (N_27465,N_26558,N_26520);
xnor U27466 (N_27466,N_26219,N_26880);
and U27467 (N_27467,N_26615,N_26030);
nand U27468 (N_27468,N_26765,N_26475);
and U27469 (N_27469,N_26784,N_26296);
and U27470 (N_27470,N_26535,N_26166);
nand U27471 (N_27471,N_26268,N_26463);
and U27472 (N_27472,N_26754,N_26574);
nor U27473 (N_27473,N_26270,N_26776);
xor U27474 (N_27474,N_26703,N_26311);
and U27475 (N_27475,N_26609,N_26821);
xnor U27476 (N_27476,N_26360,N_26779);
nand U27477 (N_27477,N_26253,N_26749);
or U27478 (N_27478,N_26198,N_26336);
or U27479 (N_27479,N_26081,N_26622);
xnor U27480 (N_27480,N_26812,N_26977);
nand U27481 (N_27481,N_26472,N_26980);
nor U27482 (N_27482,N_26039,N_26737);
nand U27483 (N_27483,N_26123,N_26842);
and U27484 (N_27484,N_26454,N_26690);
nand U27485 (N_27485,N_26200,N_26833);
or U27486 (N_27486,N_26630,N_26525);
nor U27487 (N_27487,N_26509,N_26487);
and U27488 (N_27488,N_26820,N_26492);
or U27489 (N_27489,N_26519,N_26864);
and U27490 (N_27490,N_26258,N_26795);
and U27491 (N_27491,N_26806,N_26886);
nand U27492 (N_27492,N_26214,N_26403);
xor U27493 (N_27493,N_26294,N_26937);
or U27494 (N_27494,N_26966,N_26555);
nor U27495 (N_27495,N_26212,N_26063);
or U27496 (N_27496,N_26987,N_26577);
nand U27497 (N_27497,N_26963,N_26554);
or U27498 (N_27498,N_26674,N_26315);
or U27499 (N_27499,N_26075,N_26451);
or U27500 (N_27500,N_26341,N_26204);
xor U27501 (N_27501,N_26662,N_26523);
or U27502 (N_27502,N_26747,N_26991);
xnor U27503 (N_27503,N_26016,N_26020);
and U27504 (N_27504,N_26375,N_26120);
nand U27505 (N_27505,N_26628,N_26904);
nand U27506 (N_27506,N_26727,N_26391);
nand U27507 (N_27507,N_26516,N_26953);
nand U27508 (N_27508,N_26471,N_26454);
and U27509 (N_27509,N_26523,N_26845);
xnor U27510 (N_27510,N_26749,N_26491);
nand U27511 (N_27511,N_26799,N_26549);
or U27512 (N_27512,N_26772,N_26153);
nor U27513 (N_27513,N_26825,N_26561);
and U27514 (N_27514,N_26489,N_26562);
nor U27515 (N_27515,N_26097,N_26030);
nor U27516 (N_27516,N_26863,N_26884);
and U27517 (N_27517,N_26930,N_26900);
xnor U27518 (N_27518,N_26437,N_26422);
nor U27519 (N_27519,N_26503,N_26289);
and U27520 (N_27520,N_26482,N_26703);
or U27521 (N_27521,N_26034,N_26913);
nand U27522 (N_27522,N_26473,N_26802);
nor U27523 (N_27523,N_26538,N_26254);
or U27524 (N_27524,N_26274,N_26912);
nor U27525 (N_27525,N_26288,N_26444);
xor U27526 (N_27526,N_26787,N_26884);
nor U27527 (N_27527,N_26503,N_26535);
nor U27528 (N_27528,N_26997,N_26723);
nor U27529 (N_27529,N_26927,N_26707);
and U27530 (N_27530,N_26937,N_26276);
nand U27531 (N_27531,N_26017,N_26990);
and U27532 (N_27532,N_26479,N_26485);
xnor U27533 (N_27533,N_26038,N_26780);
or U27534 (N_27534,N_26223,N_26193);
and U27535 (N_27535,N_26103,N_26998);
and U27536 (N_27536,N_26422,N_26994);
and U27537 (N_27537,N_26314,N_26944);
nand U27538 (N_27538,N_26744,N_26048);
xnor U27539 (N_27539,N_26914,N_26893);
and U27540 (N_27540,N_26977,N_26352);
nor U27541 (N_27541,N_26859,N_26874);
xnor U27542 (N_27542,N_26642,N_26238);
nor U27543 (N_27543,N_26203,N_26171);
xnor U27544 (N_27544,N_26967,N_26850);
nand U27545 (N_27545,N_26165,N_26989);
nor U27546 (N_27546,N_26382,N_26723);
nor U27547 (N_27547,N_26710,N_26716);
xnor U27548 (N_27548,N_26628,N_26587);
xnor U27549 (N_27549,N_26177,N_26204);
or U27550 (N_27550,N_26716,N_26330);
and U27551 (N_27551,N_26320,N_26818);
or U27552 (N_27552,N_26099,N_26087);
or U27553 (N_27553,N_26578,N_26887);
xor U27554 (N_27554,N_26463,N_26110);
xnor U27555 (N_27555,N_26219,N_26862);
nand U27556 (N_27556,N_26092,N_26276);
nand U27557 (N_27557,N_26105,N_26597);
nor U27558 (N_27558,N_26256,N_26322);
xor U27559 (N_27559,N_26399,N_26840);
and U27560 (N_27560,N_26634,N_26991);
nand U27561 (N_27561,N_26598,N_26850);
nor U27562 (N_27562,N_26403,N_26184);
or U27563 (N_27563,N_26866,N_26041);
and U27564 (N_27564,N_26392,N_26419);
nor U27565 (N_27565,N_26461,N_26507);
nor U27566 (N_27566,N_26819,N_26479);
xor U27567 (N_27567,N_26252,N_26302);
or U27568 (N_27568,N_26404,N_26931);
or U27569 (N_27569,N_26617,N_26707);
nor U27570 (N_27570,N_26800,N_26160);
xor U27571 (N_27571,N_26824,N_26084);
or U27572 (N_27572,N_26318,N_26510);
nor U27573 (N_27573,N_26972,N_26407);
and U27574 (N_27574,N_26290,N_26112);
nor U27575 (N_27575,N_26649,N_26419);
xor U27576 (N_27576,N_26121,N_26018);
xnor U27577 (N_27577,N_26210,N_26503);
nor U27578 (N_27578,N_26332,N_26845);
nand U27579 (N_27579,N_26084,N_26189);
nand U27580 (N_27580,N_26451,N_26219);
xor U27581 (N_27581,N_26680,N_26118);
nand U27582 (N_27582,N_26979,N_26684);
or U27583 (N_27583,N_26978,N_26081);
xnor U27584 (N_27584,N_26849,N_26824);
or U27585 (N_27585,N_26707,N_26684);
or U27586 (N_27586,N_26726,N_26406);
nand U27587 (N_27587,N_26419,N_26986);
or U27588 (N_27588,N_26914,N_26609);
and U27589 (N_27589,N_26551,N_26250);
or U27590 (N_27590,N_26637,N_26162);
nor U27591 (N_27591,N_26863,N_26223);
and U27592 (N_27592,N_26195,N_26763);
and U27593 (N_27593,N_26393,N_26281);
nand U27594 (N_27594,N_26671,N_26778);
nand U27595 (N_27595,N_26179,N_26649);
and U27596 (N_27596,N_26984,N_26598);
or U27597 (N_27597,N_26292,N_26932);
xnor U27598 (N_27598,N_26693,N_26537);
nor U27599 (N_27599,N_26421,N_26404);
and U27600 (N_27600,N_26670,N_26290);
nor U27601 (N_27601,N_26617,N_26790);
nor U27602 (N_27602,N_26472,N_26863);
and U27603 (N_27603,N_26038,N_26022);
nor U27604 (N_27604,N_26290,N_26923);
nor U27605 (N_27605,N_26503,N_26053);
or U27606 (N_27606,N_26766,N_26348);
xor U27607 (N_27607,N_26668,N_26716);
nor U27608 (N_27608,N_26332,N_26497);
or U27609 (N_27609,N_26493,N_26116);
nor U27610 (N_27610,N_26092,N_26932);
nor U27611 (N_27611,N_26578,N_26766);
and U27612 (N_27612,N_26019,N_26200);
or U27613 (N_27613,N_26675,N_26708);
nand U27614 (N_27614,N_26273,N_26594);
or U27615 (N_27615,N_26705,N_26132);
or U27616 (N_27616,N_26620,N_26697);
xor U27617 (N_27617,N_26484,N_26409);
xnor U27618 (N_27618,N_26367,N_26713);
nand U27619 (N_27619,N_26103,N_26958);
nor U27620 (N_27620,N_26423,N_26747);
xor U27621 (N_27621,N_26152,N_26930);
xnor U27622 (N_27622,N_26588,N_26229);
nand U27623 (N_27623,N_26842,N_26413);
and U27624 (N_27624,N_26331,N_26498);
and U27625 (N_27625,N_26098,N_26474);
xnor U27626 (N_27626,N_26214,N_26650);
and U27627 (N_27627,N_26732,N_26378);
or U27628 (N_27628,N_26739,N_26298);
nor U27629 (N_27629,N_26723,N_26480);
xnor U27630 (N_27630,N_26174,N_26286);
and U27631 (N_27631,N_26862,N_26331);
or U27632 (N_27632,N_26584,N_26038);
and U27633 (N_27633,N_26394,N_26194);
nor U27634 (N_27634,N_26592,N_26303);
nand U27635 (N_27635,N_26847,N_26929);
and U27636 (N_27636,N_26137,N_26290);
nor U27637 (N_27637,N_26191,N_26726);
nand U27638 (N_27638,N_26709,N_26429);
xnor U27639 (N_27639,N_26048,N_26017);
or U27640 (N_27640,N_26764,N_26668);
xnor U27641 (N_27641,N_26956,N_26978);
nor U27642 (N_27642,N_26573,N_26841);
or U27643 (N_27643,N_26205,N_26616);
xor U27644 (N_27644,N_26716,N_26784);
and U27645 (N_27645,N_26830,N_26372);
nor U27646 (N_27646,N_26905,N_26664);
nor U27647 (N_27647,N_26664,N_26150);
and U27648 (N_27648,N_26289,N_26426);
xor U27649 (N_27649,N_26591,N_26516);
nand U27650 (N_27650,N_26899,N_26911);
xor U27651 (N_27651,N_26154,N_26376);
nor U27652 (N_27652,N_26099,N_26906);
nor U27653 (N_27653,N_26134,N_26517);
xor U27654 (N_27654,N_26634,N_26454);
and U27655 (N_27655,N_26352,N_26512);
xor U27656 (N_27656,N_26124,N_26573);
or U27657 (N_27657,N_26851,N_26165);
xnor U27658 (N_27658,N_26509,N_26765);
and U27659 (N_27659,N_26669,N_26360);
nor U27660 (N_27660,N_26923,N_26659);
xnor U27661 (N_27661,N_26784,N_26361);
and U27662 (N_27662,N_26380,N_26673);
nor U27663 (N_27663,N_26156,N_26807);
nor U27664 (N_27664,N_26534,N_26671);
nor U27665 (N_27665,N_26386,N_26161);
nand U27666 (N_27666,N_26798,N_26944);
and U27667 (N_27667,N_26416,N_26538);
or U27668 (N_27668,N_26205,N_26561);
xor U27669 (N_27669,N_26843,N_26820);
nor U27670 (N_27670,N_26564,N_26096);
or U27671 (N_27671,N_26764,N_26694);
nor U27672 (N_27672,N_26193,N_26462);
nor U27673 (N_27673,N_26058,N_26708);
nand U27674 (N_27674,N_26780,N_26325);
nand U27675 (N_27675,N_26665,N_26289);
and U27676 (N_27676,N_26620,N_26484);
nor U27677 (N_27677,N_26556,N_26739);
or U27678 (N_27678,N_26967,N_26102);
and U27679 (N_27679,N_26280,N_26426);
and U27680 (N_27680,N_26343,N_26794);
nand U27681 (N_27681,N_26179,N_26841);
nand U27682 (N_27682,N_26981,N_26588);
and U27683 (N_27683,N_26985,N_26811);
xor U27684 (N_27684,N_26003,N_26011);
and U27685 (N_27685,N_26229,N_26002);
xnor U27686 (N_27686,N_26017,N_26642);
nand U27687 (N_27687,N_26378,N_26950);
nand U27688 (N_27688,N_26914,N_26005);
or U27689 (N_27689,N_26481,N_26812);
or U27690 (N_27690,N_26299,N_26892);
nand U27691 (N_27691,N_26610,N_26420);
or U27692 (N_27692,N_26699,N_26196);
nand U27693 (N_27693,N_26666,N_26315);
nand U27694 (N_27694,N_26393,N_26005);
nor U27695 (N_27695,N_26114,N_26607);
or U27696 (N_27696,N_26016,N_26579);
or U27697 (N_27697,N_26417,N_26595);
nor U27698 (N_27698,N_26839,N_26713);
xor U27699 (N_27699,N_26721,N_26529);
nor U27700 (N_27700,N_26423,N_26663);
xor U27701 (N_27701,N_26884,N_26874);
and U27702 (N_27702,N_26421,N_26247);
nor U27703 (N_27703,N_26382,N_26059);
nand U27704 (N_27704,N_26448,N_26204);
or U27705 (N_27705,N_26597,N_26688);
and U27706 (N_27706,N_26436,N_26746);
or U27707 (N_27707,N_26044,N_26603);
and U27708 (N_27708,N_26860,N_26792);
nand U27709 (N_27709,N_26480,N_26652);
nor U27710 (N_27710,N_26496,N_26401);
nor U27711 (N_27711,N_26043,N_26688);
nand U27712 (N_27712,N_26060,N_26047);
or U27713 (N_27713,N_26708,N_26874);
nand U27714 (N_27714,N_26173,N_26255);
nor U27715 (N_27715,N_26371,N_26507);
nor U27716 (N_27716,N_26933,N_26318);
or U27717 (N_27717,N_26935,N_26926);
or U27718 (N_27718,N_26568,N_26375);
nor U27719 (N_27719,N_26278,N_26544);
and U27720 (N_27720,N_26904,N_26878);
and U27721 (N_27721,N_26053,N_26673);
or U27722 (N_27722,N_26206,N_26020);
xor U27723 (N_27723,N_26784,N_26481);
xnor U27724 (N_27724,N_26133,N_26636);
or U27725 (N_27725,N_26924,N_26448);
nand U27726 (N_27726,N_26370,N_26413);
nand U27727 (N_27727,N_26222,N_26152);
xor U27728 (N_27728,N_26982,N_26409);
or U27729 (N_27729,N_26883,N_26915);
or U27730 (N_27730,N_26359,N_26167);
nor U27731 (N_27731,N_26843,N_26099);
nor U27732 (N_27732,N_26762,N_26279);
nand U27733 (N_27733,N_26730,N_26868);
and U27734 (N_27734,N_26062,N_26618);
or U27735 (N_27735,N_26008,N_26548);
nor U27736 (N_27736,N_26428,N_26007);
and U27737 (N_27737,N_26181,N_26528);
nor U27738 (N_27738,N_26276,N_26899);
xnor U27739 (N_27739,N_26664,N_26041);
or U27740 (N_27740,N_26672,N_26729);
and U27741 (N_27741,N_26493,N_26499);
and U27742 (N_27742,N_26177,N_26757);
and U27743 (N_27743,N_26865,N_26792);
nand U27744 (N_27744,N_26143,N_26453);
or U27745 (N_27745,N_26463,N_26964);
or U27746 (N_27746,N_26951,N_26483);
and U27747 (N_27747,N_26215,N_26672);
or U27748 (N_27748,N_26081,N_26599);
nor U27749 (N_27749,N_26840,N_26260);
nor U27750 (N_27750,N_26000,N_26264);
and U27751 (N_27751,N_26614,N_26139);
and U27752 (N_27752,N_26836,N_26204);
and U27753 (N_27753,N_26227,N_26096);
and U27754 (N_27754,N_26540,N_26646);
and U27755 (N_27755,N_26643,N_26411);
xnor U27756 (N_27756,N_26851,N_26805);
nor U27757 (N_27757,N_26712,N_26229);
or U27758 (N_27758,N_26138,N_26101);
and U27759 (N_27759,N_26754,N_26372);
or U27760 (N_27760,N_26721,N_26025);
nand U27761 (N_27761,N_26945,N_26039);
nand U27762 (N_27762,N_26443,N_26111);
xnor U27763 (N_27763,N_26140,N_26673);
nor U27764 (N_27764,N_26761,N_26996);
xor U27765 (N_27765,N_26160,N_26589);
xor U27766 (N_27766,N_26449,N_26160);
nand U27767 (N_27767,N_26666,N_26631);
or U27768 (N_27768,N_26075,N_26465);
nand U27769 (N_27769,N_26175,N_26396);
and U27770 (N_27770,N_26560,N_26383);
xor U27771 (N_27771,N_26878,N_26133);
nand U27772 (N_27772,N_26707,N_26776);
and U27773 (N_27773,N_26918,N_26467);
nor U27774 (N_27774,N_26358,N_26448);
or U27775 (N_27775,N_26346,N_26157);
and U27776 (N_27776,N_26140,N_26823);
xor U27777 (N_27777,N_26525,N_26227);
xnor U27778 (N_27778,N_26498,N_26232);
nor U27779 (N_27779,N_26315,N_26837);
nor U27780 (N_27780,N_26558,N_26099);
or U27781 (N_27781,N_26700,N_26036);
nor U27782 (N_27782,N_26724,N_26552);
or U27783 (N_27783,N_26279,N_26400);
nor U27784 (N_27784,N_26107,N_26206);
or U27785 (N_27785,N_26456,N_26990);
nor U27786 (N_27786,N_26349,N_26770);
xor U27787 (N_27787,N_26449,N_26926);
nand U27788 (N_27788,N_26958,N_26833);
nor U27789 (N_27789,N_26132,N_26611);
nand U27790 (N_27790,N_26225,N_26358);
or U27791 (N_27791,N_26488,N_26820);
nor U27792 (N_27792,N_26144,N_26956);
and U27793 (N_27793,N_26236,N_26868);
nor U27794 (N_27794,N_26081,N_26284);
nor U27795 (N_27795,N_26994,N_26851);
nand U27796 (N_27796,N_26310,N_26200);
xor U27797 (N_27797,N_26823,N_26062);
and U27798 (N_27798,N_26311,N_26194);
or U27799 (N_27799,N_26276,N_26708);
or U27800 (N_27800,N_26620,N_26040);
and U27801 (N_27801,N_26810,N_26428);
or U27802 (N_27802,N_26244,N_26894);
and U27803 (N_27803,N_26056,N_26837);
nand U27804 (N_27804,N_26064,N_26721);
nand U27805 (N_27805,N_26394,N_26461);
xor U27806 (N_27806,N_26577,N_26633);
or U27807 (N_27807,N_26513,N_26537);
or U27808 (N_27808,N_26489,N_26808);
and U27809 (N_27809,N_26123,N_26809);
xor U27810 (N_27810,N_26050,N_26006);
xnor U27811 (N_27811,N_26931,N_26336);
nor U27812 (N_27812,N_26062,N_26425);
xor U27813 (N_27813,N_26223,N_26771);
nand U27814 (N_27814,N_26634,N_26586);
nand U27815 (N_27815,N_26640,N_26909);
and U27816 (N_27816,N_26392,N_26493);
or U27817 (N_27817,N_26358,N_26656);
or U27818 (N_27818,N_26542,N_26709);
or U27819 (N_27819,N_26542,N_26855);
and U27820 (N_27820,N_26708,N_26801);
xnor U27821 (N_27821,N_26231,N_26982);
xnor U27822 (N_27822,N_26269,N_26498);
nand U27823 (N_27823,N_26596,N_26993);
nor U27824 (N_27824,N_26846,N_26514);
or U27825 (N_27825,N_26725,N_26117);
xnor U27826 (N_27826,N_26194,N_26156);
or U27827 (N_27827,N_26015,N_26056);
or U27828 (N_27828,N_26268,N_26185);
nand U27829 (N_27829,N_26255,N_26004);
nand U27830 (N_27830,N_26522,N_26582);
or U27831 (N_27831,N_26600,N_26561);
nor U27832 (N_27832,N_26478,N_26050);
nor U27833 (N_27833,N_26620,N_26265);
or U27834 (N_27834,N_26906,N_26781);
nor U27835 (N_27835,N_26798,N_26141);
or U27836 (N_27836,N_26640,N_26447);
or U27837 (N_27837,N_26235,N_26577);
nor U27838 (N_27838,N_26029,N_26700);
nand U27839 (N_27839,N_26178,N_26540);
nor U27840 (N_27840,N_26896,N_26460);
xnor U27841 (N_27841,N_26302,N_26744);
nor U27842 (N_27842,N_26940,N_26820);
and U27843 (N_27843,N_26668,N_26548);
nor U27844 (N_27844,N_26054,N_26701);
xor U27845 (N_27845,N_26873,N_26848);
nor U27846 (N_27846,N_26402,N_26900);
nand U27847 (N_27847,N_26206,N_26682);
and U27848 (N_27848,N_26896,N_26110);
xor U27849 (N_27849,N_26240,N_26864);
xor U27850 (N_27850,N_26073,N_26880);
and U27851 (N_27851,N_26735,N_26627);
nand U27852 (N_27852,N_26156,N_26365);
or U27853 (N_27853,N_26480,N_26459);
nor U27854 (N_27854,N_26124,N_26647);
nor U27855 (N_27855,N_26386,N_26186);
and U27856 (N_27856,N_26591,N_26781);
nand U27857 (N_27857,N_26048,N_26103);
nand U27858 (N_27858,N_26754,N_26681);
or U27859 (N_27859,N_26895,N_26580);
or U27860 (N_27860,N_26475,N_26341);
and U27861 (N_27861,N_26913,N_26822);
nor U27862 (N_27862,N_26097,N_26761);
and U27863 (N_27863,N_26012,N_26413);
xnor U27864 (N_27864,N_26880,N_26550);
and U27865 (N_27865,N_26340,N_26438);
or U27866 (N_27866,N_26206,N_26405);
xor U27867 (N_27867,N_26166,N_26494);
or U27868 (N_27868,N_26728,N_26939);
or U27869 (N_27869,N_26684,N_26374);
nor U27870 (N_27870,N_26694,N_26306);
nand U27871 (N_27871,N_26570,N_26636);
nor U27872 (N_27872,N_26876,N_26034);
and U27873 (N_27873,N_26266,N_26472);
nand U27874 (N_27874,N_26683,N_26147);
nand U27875 (N_27875,N_26710,N_26863);
xor U27876 (N_27876,N_26831,N_26531);
nand U27877 (N_27877,N_26876,N_26831);
or U27878 (N_27878,N_26896,N_26942);
or U27879 (N_27879,N_26372,N_26442);
nor U27880 (N_27880,N_26487,N_26072);
and U27881 (N_27881,N_26598,N_26741);
xnor U27882 (N_27882,N_26540,N_26286);
or U27883 (N_27883,N_26110,N_26478);
nor U27884 (N_27884,N_26797,N_26327);
nor U27885 (N_27885,N_26035,N_26391);
and U27886 (N_27886,N_26963,N_26458);
and U27887 (N_27887,N_26543,N_26288);
xnor U27888 (N_27888,N_26053,N_26371);
nand U27889 (N_27889,N_26774,N_26771);
and U27890 (N_27890,N_26001,N_26326);
and U27891 (N_27891,N_26632,N_26712);
nand U27892 (N_27892,N_26664,N_26400);
or U27893 (N_27893,N_26968,N_26724);
or U27894 (N_27894,N_26595,N_26165);
nand U27895 (N_27895,N_26269,N_26759);
and U27896 (N_27896,N_26279,N_26336);
and U27897 (N_27897,N_26379,N_26701);
xnor U27898 (N_27898,N_26204,N_26572);
or U27899 (N_27899,N_26769,N_26010);
xnor U27900 (N_27900,N_26097,N_26072);
or U27901 (N_27901,N_26496,N_26588);
nor U27902 (N_27902,N_26062,N_26019);
nor U27903 (N_27903,N_26305,N_26178);
xor U27904 (N_27904,N_26889,N_26824);
nand U27905 (N_27905,N_26843,N_26929);
nand U27906 (N_27906,N_26255,N_26027);
xor U27907 (N_27907,N_26041,N_26647);
nor U27908 (N_27908,N_26708,N_26660);
and U27909 (N_27909,N_26093,N_26242);
nor U27910 (N_27910,N_26304,N_26045);
nor U27911 (N_27911,N_26725,N_26384);
and U27912 (N_27912,N_26022,N_26206);
and U27913 (N_27913,N_26663,N_26081);
or U27914 (N_27914,N_26767,N_26727);
nor U27915 (N_27915,N_26842,N_26128);
xnor U27916 (N_27916,N_26397,N_26573);
nor U27917 (N_27917,N_26056,N_26621);
nor U27918 (N_27918,N_26519,N_26436);
nor U27919 (N_27919,N_26386,N_26635);
nand U27920 (N_27920,N_26791,N_26961);
nand U27921 (N_27921,N_26327,N_26740);
nor U27922 (N_27922,N_26675,N_26360);
nor U27923 (N_27923,N_26904,N_26648);
and U27924 (N_27924,N_26021,N_26679);
nor U27925 (N_27925,N_26991,N_26459);
nand U27926 (N_27926,N_26427,N_26268);
or U27927 (N_27927,N_26338,N_26679);
nor U27928 (N_27928,N_26186,N_26925);
or U27929 (N_27929,N_26419,N_26807);
or U27930 (N_27930,N_26100,N_26950);
nor U27931 (N_27931,N_26141,N_26241);
nor U27932 (N_27932,N_26832,N_26693);
nand U27933 (N_27933,N_26992,N_26301);
xor U27934 (N_27934,N_26167,N_26112);
or U27935 (N_27935,N_26388,N_26941);
nor U27936 (N_27936,N_26445,N_26323);
xnor U27937 (N_27937,N_26089,N_26826);
xor U27938 (N_27938,N_26200,N_26937);
and U27939 (N_27939,N_26970,N_26127);
nand U27940 (N_27940,N_26833,N_26141);
nor U27941 (N_27941,N_26853,N_26815);
or U27942 (N_27942,N_26503,N_26058);
or U27943 (N_27943,N_26395,N_26465);
xor U27944 (N_27944,N_26688,N_26999);
and U27945 (N_27945,N_26498,N_26501);
or U27946 (N_27946,N_26400,N_26602);
xor U27947 (N_27947,N_26081,N_26390);
and U27948 (N_27948,N_26780,N_26705);
or U27949 (N_27949,N_26827,N_26165);
nand U27950 (N_27950,N_26380,N_26403);
nor U27951 (N_27951,N_26144,N_26788);
nor U27952 (N_27952,N_26510,N_26687);
nor U27953 (N_27953,N_26301,N_26948);
nand U27954 (N_27954,N_26032,N_26297);
and U27955 (N_27955,N_26015,N_26691);
and U27956 (N_27956,N_26272,N_26355);
xor U27957 (N_27957,N_26064,N_26359);
or U27958 (N_27958,N_26124,N_26170);
nor U27959 (N_27959,N_26493,N_26766);
and U27960 (N_27960,N_26090,N_26412);
nand U27961 (N_27961,N_26162,N_26197);
and U27962 (N_27962,N_26907,N_26476);
nand U27963 (N_27963,N_26855,N_26473);
nand U27964 (N_27964,N_26295,N_26248);
and U27965 (N_27965,N_26884,N_26304);
nand U27966 (N_27966,N_26605,N_26867);
nand U27967 (N_27967,N_26436,N_26438);
xor U27968 (N_27968,N_26319,N_26911);
and U27969 (N_27969,N_26928,N_26257);
nand U27970 (N_27970,N_26778,N_26977);
or U27971 (N_27971,N_26793,N_26964);
or U27972 (N_27972,N_26668,N_26675);
and U27973 (N_27973,N_26834,N_26925);
nand U27974 (N_27974,N_26607,N_26504);
nand U27975 (N_27975,N_26415,N_26296);
nor U27976 (N_27976,N_26153,N_26278);
xor U27977 (N_27977,N_26205,N_26181);
nand U27978 (N_27978,N_26352,N_26160);
or U27979 (N_27979,N_26756,N_26217);
xnor U27980 (N_27980,N_26132,N_26764);
or U27981 (N_27981,N_26046,N_26162);
or U27982 (N_27982,N_26822,N_26647);
or U27983 (N_27983,N_26557,N_26817);
nor U27984 (N_27984,N_26788,N_26467);
nand U27985 (N_27985,N_26386,N_26169);
nor U27986 (N_27986,N_26882,N_26907);
xor U27987 (N_27987,N_26458,N_26979);
nor U27988 (N_27988,N_26723,N_26246);
xnor U27989 (N_27989,N_26157,N_26816);
nor U27990 (N_27990,N_26652,N_26593);
xor U27991 (N_27991,N_26921,N_26408);
nor U27992 (N_27992,N_26709,N_26568);
nor U27993 (N_27993,N_26608,N_26054);
and U27994 (N_27994,N_26717,N_26585);
and U27995 (N_27995,N_26782,N_26804);
nand U27996 (N_27996,N_26607,N_26000);
or U27997 (N_27997,N_26684,N_26349);
or U27998 (N_27998,N_26978,N_26357);
or U27999 (N_27999,N_26715,N_26562);
nor U28000 (N_28000,N_27665,N_27449);
or U28001 (N_28001,N_27161,N_27589);
or U28002 (N_28002,N_27671,N_27151);
xor U28003 (N_28003,N_27374,N_27229);
and U28004 (N_28004,N_27350,N_27525);
nor U28005 (N_28005,N_27450,N_27501);
and U28006 (N_28006,N_27647,N_27339);
and U28007 (N_28007,N_27578,N_27454);
xor U28008 (N_28008,N_27199,N_27863);
xnor U28009 (N_28009,N_27539,N_27176);
nor U28010 (N_28010,N_27220,N_27907);
xor U28011 (N_28011,N_27856,N_27858);
or U28012 (N_28012,N_27834,N_27222);
nand U28013 (N_28013,N_27184,N_27235);
and U28014 (N_28014,N_27205,N_27861);
and U28015 (N_28015,N_27346,N_27909);
and U28016 (N_28016,N_27568,N_27328);
and U28017 (N_28017,N_27860,N_27726);
nor U28018 (N_28018,N_27756,N_27285);
or U28019 (N_28019,N_27778,N_27215);
and U28020 (N_28020,N_27893,N_27982);
nor U28021 (N_28021,N_27470,N_27761);
nand U28022 (N_28022,N_27476,N_27195);
nand U28023 (N_28023,N_27791,N_27074);
nor U28024 (N_28024,N_27685,N_27786);
nand U28025 (N_28025,N_27518,N_27737);
nand U28026 (N_28026,N_27773,N_27129);
and U28027 (N_28027,N_27931,N_27182);
or U28028 (N_28028,N_27849,N_27748);
or U28029 (N_28029,N_27755,N_27677);
or U28030 (N_28030,N_27028,N_27260);
nand U28031 (N_28031,N_27356,N_27419);
xor U28032 (N_28032,N_27366,N_27230);
xnor U28033 (N_28033,N_27088,N_27968);
nand U28034 (N_28034,N_27134,N_27365);
nor U28035 (N_28035,N_27186,N_27768);
xnor U28036 (N_28036,N_27289,N_27401);
nor U28037 (N_28037,N_27337,N_27936);
and U28038 (N_28038,N_27293,N_27505);
nor U28039 (N_28039,N_27969,N_27524);
and U28040 (N_28040,N_27190,N_27654);
nor U28041 (N_28041,N_27790,N_27455);
nor U28042 (N_28042,N_27261,N_27713);
and U28043 (N_28043,N_27206,N_27057);
nor U28044 (N_28044,N_27036,N_27140);
and U28045 (N_28045,N_27110,N_27800);
nor U28046 (N_28046,N_27839,N_27574);
xnor U28047 (N_28047,N_27692,N_27885);
nor U28048 (N_28048,N_27546,N_27271);
nand U28049 (N_28049,N_27663,N_27711);
or U28050 (N_28050,N_27444,N_27447);
nor U28051 (N_28051,N_27407,N_27270);
or U28052 (N_28052,N_27256,N_27548);
xnor U28053 (N_28053,N_27996,N_27650);
nand U28054 (N_28054,N_27845,N_27104);
nor U28055 (N_28055,N_27462,N_27352);
nor U28056 (N_28056,N_27978,N_27515);
nor U28057 (N_28057,N_27794,N_27379);
nor U28058 (N_28058,N_27167,N_27509);
nand U28059 (N_28059,N_27141,N_27932);
or U28060 (N_28060,N_27133,N_27810);
xnor U28061 (N_28061,N_27779,N_27880);
nand U28062 (N_28062,N_27322,N_27171);
xor U28063 (N_28063,N_27188,N_27543);
nor U28064 (N_28064,N_27914,N_27891);
nand U28065 (N_28065,N_27106,N_27306);
or U28066 (N_28066,N_27537,N_27632);
xnor U28067 (N_28067,N_27646,N_27488);
xor U28068 (N_28068,N_27612,N_27248);
nand U28069 (N_28069,N_27662,N_27701);
and U28070 (N_28070,N_27915,N_27466);
nand U28071 (N_28071,N_27441,N_27682);
nor U28072 (N_28072,N_27926,N_27198);
or U28073 (N_28073,N_27942,N_27999);
nor U28074 (N_28074,N_27239,N_27850);
or U28075 (N_28075,N_27517,N_27338);
nor U28076 (N_28076,N_27014,N_27812);
and U28077 (N_28077,N_27103,N_27012);
and U28078 (N_28078,N_27687,N_27838);
nand U28079 (N_28079,N_27808,N_27175);
nand U28080 (N_28080,N_27181,N_27570);
nor U28081 (N_28081,N_27991,N_27189);
xnor U28082 (N_28082,N_27183,N_27118);
or U28083 (N_28083,N_27301,N_27935);
or U28084 (N_28084,N_27376,N_27920);
and U28085 (N_28085,N_27272,N_27811);
nor U28086 (N_28086,N_27866,N_27976);
nor U28087 (N_28087,N_27855,N_27562);
nand U28088 (N_28088,N_27819,N_27253);
nand U28089 (N_28089,N_27180,N_27435);
and U28090 (N_28090,N_27255,N_27284);
xor U28091 (N_28091,N_27010,N_27776);
or U28092 (N_28092,N_27705,N_27157);
xor U28093 (N_28093,N_27656,N_27152);
or U28094 (N_28094,N_27298,N_27381);
nor U28095 (N_28095,N_27130,N_27623);
nor U28096 (N_28096,N_27442,N_27314);
xor U28097 (N_28097,N_27373,N_27496);
nand U28098 (N_28098,N_27963,N_27251);
or U28099 (N_28099,N_27032,N_27565);
and U28100 (N_28100,N_27307,N_27681);
nor U28101 (N_28101,N_27056,N_27415);
xnor U28102 (N_28102,N_27109,N_27030);
or U28103 (N_28103,N_27257,N_27053);
nand U28104 (N_28104,N_27712,N_27445);
or U28105 (N_28105,N_27008,N_27164);
nand U28106 (N_28106,N_27234,N_27813);
or U28107 (N_28107,N_27689,N_27657);
nor U28108 (N_28108,N_27390,N_27026);
and U28109 (N_28109,N_27925,N_27486);
nand U28110 (N_28110,N_27410,N_27785);
or U28111 (N_28111,N_27459,N_27604);
nand U28112 (N_28112,N_27553,N_27400);
nor U28113 (N_28113,N_27990,N_27413);
and U28114 (N_28114,N_27055,N_27916);
or U28115 (N_28115,N_27516,N_27734);
nand U28116 (N_28116,N_27159,N_27512);
and U28117 (N_28117,N_27347,N_27933);
or U28118 (N_28118,N_27949,N_27383);
and U28119 (N_28119,N_27923,N_27414);
and U28120 (N_28120,N_27440,N_27579);
and U28121 (N_28121,N_27448,N_27841);
or U28122 (N_28122,N_27331,N_27136);
nor U28123 (N_28123,N_27047,N_27492);
or U28124 (N_28124,N_27142,N_27070);
nor U28125 (N_28125,N_27258,N_27250);
nor U28126 (N_28126,N_27762,N_27870);
nand U28127 (N_28127,N_27487,N_27924);
nor U28128 (N_28128,N_27054,N_27002);
and U28129 (N_28129,N_27985,N_27150);
xnor U28130 (N_28130,N_27479,N_27912);
nand U28131 (N_28131,N_27829,N_27236);
xnor U28132 (N_28132,N_27581,N_27867);
nor U28133 (N_28133,N_27040,N_27742);
xor U28134 (N_28134,N_27947,N_27636);
nand U28135 (N_28135,N_27817,N_27340);
nor U28136 (N_28136,N_27956,N_27502);
and U28137 (N_28137,N_27994,N_27266);
nor U28138 (N_28138,N_27704,N_27830);
nor U28139 (N_28139,N_27017,N_27769);
xnor U28140 (N_28140,N_27310,N_27661);
nor U28141 (N_28141,N_27523,N_27918);
or U28142 (N_28142,N_27992,N_27904);
and U28143 (N_28143,N_27315,N_27464);
or U28144 (N_28144,N_27264,N_27023);
and U28145 (N_28145,N_27165,N_27600);
or U28146 (N_28146,N_27732,N_27637);
nand U28147 (N_28147,N_27007,N_27280);
nand U28148 (N_28148,N_27513,N_27369);
nor U28149 (N_28149,N_27249,N_27308);
nand U28150 (N_28150,N_27938,N_27836);
nor U28151 (N_28151,N_27719,N_27342);
xor U28152 (N_28152,N_27588,N_27320);
or U28153 (N_28153,N_27491,N_27847);
nor U28154 (N_28154,N_27541,N_27670);
and U28155 (N_28155,N_27006,N_27622);
xor U28156 (N_28156,N_27898,N_27997);
or U28157 (N_28157,N_27137,N_27745);
or U28158 (N_28158,N_27408,N_27341);
or U28159 (N_28159,N_27065,N_27886);
nor U28160 (N_28160,N_27254,N_27783);
nor U28161 (N_28161,N_27608,N_27864);
xor U28162 (N_28162,N_27451,N_27333);
xnor U28163 (N_28163,N_27433,N_27883);
nand U28164 (N_28164,N_27169,N_27981);
xor U28165 (N_28165,N_27927,N_27378);
nand U28166 (N_28166,N_27594,N_27094);
nor U28167 (N_28167,N_27717,N_27563);
nand U28168 (N_28168,N_27843,N_27031);
nand U28169 (N_28169,N_27766,N_27672);
and U28170 (N_28170,N_27018,N_27245);
and U28171 (N_28171,N_27640,N_27716);
xnor U28172 (N_28172,N_27090,N_27598);
nand U28173 (N_28173,N_27591,N_27542);
or U28174 (N_28174,N_27831,N_27889);
and U28175 (N_28175,N_27382,N_27452);
nand U28176 (N_28176,N_27075,N_27709);
xnor U28177 (N_28177,N_27399,N_27240);
nor U28178 (N_28178,N_27765,N_27678);
nor U28179 (N_28179,N_27823,N_27360);
or U28180 (N_28180,N_27232,N_27416);
or U28181 (N_28181,N_27204,N_27219);
xnor U28182 (N_28182,N_27368,N_27559);
nor U28183 (N_28183,N_27013,N_27805);
nor U28184 (N_28184,N_27004,N_27406);
nand U28185 (N_28185,N_27039,N_27780);
xor U28186 (N_28186,N_27560,N_27443);
nand U28187 (N_28187,N_27900,N_27770);
xnor U28188 (N_28188,N_27101,N_27434);
and U28189 (N_28189,N_27621,N_27021);
nand U28190 (N_28190,N_27336,N_27585);
or U28191 (N_28191,N_27547,N_27531);
nor U28192 (N_28192,N_27475,N_27166);
nor U28193 (N_28193,N_27644,N_27071);
nand U28194 (N_28194,N_27353,N_27639);
nor U28195 (N_28195,N_27292,N_27767);
and U28196 (N_28196,N_27457,N_27624);
xor U28197 (N_28197,N_27837,N_27821);
xor U28198 (N_28198,N_27193,N_27828);
and U28199 (N_28199,N_27172,N_27357);
nand U28200 (N_28200,N_27659,N_27951);
nand U28201 (N_28201,N_27312,N_27558);
nor U28202 (N_28202,N_27877,N_27741);
nand U28203 (N_28203,N_27510,N_27059);
xor U28204 (N_28204,N_27939,N_27263);
xor U28205 (N_28205,N_27730,N_27080);
xnor U28206 (N_28206,N_27595,N_27422);
and U28207 (N_28207,N_27634,N_27268);
nand U28208 (N_28208,N_27185,N_27179);
xnor U28209 (N_28209,N_27439,N_27987);
nand U28210 (N_28210,N_27241,N_27122);
and U28211 (N_28211,N_27123,N_27706);
xor U28212 (N_28212,N_27526,N_27297);
and U28213 (N_28213,N_27156,N_27262);
xnor U28214 (N_28214,N_27428,N_27989);
and U28215 (N_28215,N_27750,N_27566);
nand U28216 (N_28216,N_27603,N_27868);
nand U28217 (N_28217,N_27710,N_27265);
nor U28218 (N_28218,N_27477,N_27417);
and U28219 (N_28219,N_27691,N_27120);
nand U28220 (N_28220,N_27522,N_27027);
xnor U28221 (N_28221,N_27132,N_27899);
nand U28222 (N_28222,N_27102,N_27158);
nor U28223 (N_28223,N_27873,N_27354);
xor U28224 (N_28224,N_27698,N_27163);
nor U28225 (N_28225,N_27100,N_27051);
and U28226 (N_28226,N_27597,N_27645);
nand U28227 (N_28227,N_27798,N_27820);
or U28228 (N_28228,N_27816,N_27749);
and U28229 (N_28229,N_27393,N_27940);
or U28230 (N_28230,N_27325,N_27286);
xnor U28231 (N_28231,N_27370,N_27740);
nor U28232 (N_28232,N_27695,N_27784);
or U28233 (N_28233,N_27038,N_27019);
nand U28234 (N_28234,N_27041,N_27641);
xor U28235 (N_28235,N_27529,N_27403);
nor U28236 (N_28236,N_27962,N_27601);
nor U28237 (N_28237,N_27246,N_27398);
nand U28238 (N_28238,N_27775,N_27064);
nand U28239 (N_28239,N_27627,N_27826);
nand U28240 (N_28240,N_27972,N_27429);
xnor U28241 (N_28241,N_27571,N_27679);
or U28242 (N_28242,N_27299,N_27950);
xnor U28243 (N_28243,N_27804,N_27888);
xor U28244 (N_28244,N_27114,N_27467);
nor U28245 (N_28245,N_27922,N_27580);
and U28246 (N_28246,N_27535,N_27807);
nand U28247 (N_28247,N_27676,N_27209);
xor U28248 (N_28248,N_27386,N_27469);
xnor U28249 (N_28249,N_27105,N_27733);
and U28250 (N_28250,N_27519,N_27126);
xor U28251 (N_28251,N_27009,N_27960);
nand U28252 (N_28252,N_27721,N_27921);
xor U28253 (N_28253,N_27049,N_27890);
nand U28254 (N_28254,N_27735,N_27564);
xnor U28255 (N_28255,N_27667,N_27037);
or U28256 (N_28256,N_27093,N_27952);
xor U28257 (N_28257,N_27375,N_27660);
nand U28258 (N_28258,N_27001,N_27000);
nor U28259 (N_28259,N_27979,N_27503);
nand U28260 (N_28260,N_27842,N_27569);
nand U28261 (N_28261,N_27143,N_27533);
and U28262 (N_28262,N_27832,N_27202);
or U28263 (N_28263,N_27789,N_27033);
nor U28264 (N_28264,N_27084,N_27896);
or U28265 (N_28265,N_27882,N_27556);
and U28266 (N_28266,N_27696,N_27584);
xor U28267 (N_28267,N_27472,N_27471);
xor U28268 (N_28268,N_27605,N_27048);
or U28269 (N_28269,N_27117,N_27988);
nor U28270 (N_28270,N_27984,N_27729);
nor U28271 (N_28271,N_27977,N_27046);
nor U28272 (N_28272,N_27674,N_27825);
and U28273 (N_28273,N_27290,N_27231);
xnor U28274 (N_28274,N_27154,N_27803);
and U28275 (N_28275,N_27324,N_27957);
and U28276 (N_28276,N_27304,N_27527);
nor U28277 (N_28277,N_27361,N_27629);
nor U28278 (N_28278,N_27108,N_27971);
nand U28279 (N_28279,N_27772,N_27015);
nand U28280 (N_28280,N_27911,N_27799);
xor U28281 (N_28281,N_27430,N_27224);
or U28282 (N_28282,N_27576,N_27680);
nand U28283 (N_28283,N_27693,N_27210);
or U28284 (N_28284,N_27908,N_27690);
xor U28285 (N_28285,N_27617,N_27943);
nand U28286 (N_28286,N_27252,N_27635);
nor U28287 (N_28287,N_27752,N_27282);
and U28288 (N_28288,N_27930,N_27178);
nor U28289 (N_28289,N_27625,N_27489);
and U28290 (N_28290,N_27887,N_27387);
xnor U28291 (N_28291,N_27587,N_27633);
and U28292 (N_28292,N_27731,N_27355);
or U28293 (N_28293,N_27853,N_27349);
nand U28294 (N_28294,N_27801,N_27555);
and U28295 (N_28295,N_27431,N_27045);
or U28296 (N_28296,N_27481,N_27411);
or U28297 (N_28297,N_27953,N_27929);
xnor U28298 (N_28298,N_27494,N_27020);
or U28299 (N_28299,N_27484,N_27388);
xor U28300 (N_28300,N_27302,N_27112);
xor U28301 (N_28301,N_27424,N_27371);
nand U28302 (N_28302,N_27066,N_27099);
xnor U28303 (N_28303,N_27363,N_27316);
and U28304 (N_28304,N_27022,N_27233);
or U28305 (N_28305,N_27139,N_27396);
and U28306 (N_28306,N_27421,N_27975);
nor U28307 (N_28307,N_27335,N_27892);
xnor U28308 (N_28308,N_27458,N_27964);
nand U28309 (N_28309,N_27217,N_27707);
or U28310 (N_28310,N_27086,N_27664);
xor U28311 (N_28311,N_27788,N_27247);
and U28312 (N_28312,N_27702,N_27872);
or U28313 (N_28313,N_27753,N_27278);
or U28314 (N_28314,N_27196,N_27500);
xnor U28315 (N_28315,N_27177,N_27277);
nand U28316 (N_28316,N_27980,N_27763);
or U28317 (N_28317,N_27242,N_27092);
nand U28318 (N_28318,N_27714,N_27683);
nand U28319 (N_28319,N_27514,N_27694);
nand U28320 (N_28320,N_27050,N_27534);
xnor U28321 (N_28321,N_27747,N_27283);
and U28322 (N_28322,N_27586,N_27067);
or U28323 (N_28323,N_27961,N_27743);
nor U28324 (N_28324,N_27493,N_27311);
nand U28325 (N_28325,N_27934,N_27998);
or U28326 (N_28326,N_27453,N_27986);
or U28327 (N_28327,N_27317,N_27876);
and U28328 (N_28328,N_27857,N_27402);
xor U28329 (N_28329,N_27536,N_27613);
xor U28330 (N_28330,N_27135,N_27699);
nand U28331 (N_28331,N_27508,N_27119);
nor U28332 (N_28332,N_27881,N_27226);
and U28333 (N_28333,N_27759,N_27630);
nand U28334 (N_28334,N_27967,N_27865);
xor U28335 (N_28335,N_27029,N_27824);
xor U28336 (N_28336,N_27862,N_27060);
nand U28337 (N_28337,N_27582,N_27993);
nand U28338 (N_28338,N_27498,N_27906);
nand U28339 (N_28339,N_27362,N_27276);
xnor U28340 (N_28340,N_27507,N_27116);
or U28341 (N_28341,N_27025,N_27194);
xor U28342 (N_28342,N_27395,N_27557);
nor U28343 (N_28343,N_27330,N_27802);
and U28344 (N_28344,N_27173,N_27974);
and U28345 (N_28345,N_27225,N_27153);
and U28346 (N_28346,N_27572,N_27653);
nand U28347 (N_28347,N_27295,N_27684);
and U28348 (N_28348,N_27746,N_27955);
or U28349 (N_28349,N_27567,N_27473);
nand U28350 (N_28350,N_27288,N_27024);
nand U28351 (N_28351,N_27851,N_27544);
and U28352 (N_28352,N_27884,N_27609);
or U28353 (N_28353,N_27358,N_27296);
and U28354 (N_28354,N_27063,N_27874);
and U28355 (N_28355,N_27372,N_27468);
or U28356 (N_28356,N_27532,N_27300);
nor U28357 (N_28357,N_27835,N_27545);
or U28358 (N_28358,N_27797,N_27787);
and U28359 (N_28359,N_27208,N_27364);
nor U28360 (N_28360,N_27593,N_27607);
and U28361 (N_28361,N_27111,N_27287);
nand U28362 (N_28362,N_27655,N_27425);
or U28363 (N_28363,N_27554,N_27561);
nand U28364 (N_28364,N_27069,N_27970);
or U28365 (N_28365,N_27162,N_27432);
xnor U28366 (N_28366,N_27506,N_27385);
and U28367 (N_28367,N_27076,N_27854);
nand U28368 (N_28368,N_27903,N_27638);
or U28369 (N_28369,N_27959,N_27078);
or U28370 (N_28370,N_27966,N_27200);
and U28371 (N_28371,N_27329,N_27344);
and U28372 (N_28372,N_27207,N_27483);
or U28373 (N_28373,N_27723,N_27902);
nand U28374 (N_28374,N_27648,N_27016);
and U28375 (N_28375,N_27958,N_27274);
nand U28376 (N_28376,N_27323,N_27897);
xor U28377 (N_28377,N_27042,N_27818);
and U28378 (N_28378,N_27697,N_27115);
nor U28379 (N_28379,N_27079,N_27197);
xnor U28380 (N_28380,N_27774,N_27146);
nand U28381 (N_28381,N_27223,N_27614);
or U28382 (N_28382,N_27313,N_27575);
and U28383 (N_28383,N_27326,N_27279);
xor U28384 (N_28384,N_27538,N_27058);
or U28385 (N_28385,N_27550,N_27822);
and U28386 (N_28386,N_27616,N_27795);
nor U28387 (N_28387,N_27035,N_27305);
and U28388 (N_28388,N_27218,N_27945);
nand U28389 (N_28389,N_27214,N_27666);
and U28390 (N_28390,N_27781,N_27504);
nor U28391 (N_28391,N_27520,N_27669);
nor U28392 (N_28392,N_27573,N_27148);
or U28393 (N_28393,N_27725,N_27715);
xnor U28394 (N_28394,N_27490,N_27334);
xnor U28395 (N_28395,N_27549,N_27269);
xnor U28396 (N_28396,N_27995,N_27793);
nand U28397 (N_28397,N_27227,N_27160);
or U28398 (N_28398,N_27348,N_27082);
and U28399 (N_28399,N_27642,N_27777);
nand U28400 (N_28400,N_27380,N_27894);
and U28401 (N_28401,N_27626,N_27131);
or U28402 (N_28402,N_27673,N_27782);
and U28403 (N_28403,N_27044,N_27409);
or U28404 (N_28404,N_27688,N_27062);
or U28405 (N_28405,N_27618,N_27436);
or U28406 (N_28406,N_27391,N_27700);
nand U28407 (N_28407,N_27446,N_27461);
xor U28408 (N_28408,N_27703,N_27081);
and U28409 (N_28409,N_27155,N_27244);
and U28410 (N_28410,N_27345,N_27658);
xnor U28411 (N_28411,N_27061,N_27003);
nor U28412 (N_28412,N_27211,N_27221);
nand U28413 (N_28413,N_27760,N_27879);
xnor U28414 (N_28414,N_27846,N_27460);
nor U28415 (N_28415,N_27610,N_27125);
or U28416 (N_28416,N_27815,N_27203);
xnor U28417 (N_28417,N_27259,N_27083);
or U28418 (N_28418,N_27187,N_27583);
nor U28419 (N_28419,N_27552,N_27859);
nor U28420 (N_28420,N_27771,N_27919);
and U28421 (N_28421,N_27191,N_27599);
nor U28422 (N_28422,N_27343,N_27392);
xnor U28423 (N_28423,N_27649,N_27170);
or U28424 (N_28424,N_27944,N_27764);
nand U28425 (N_28425,N_27954,N_27814);
xor U28426 (N_28426,N_27073,N_27412);
or U28427 (N_28427,N_27420,N_27739);
nor U28428 (N_28428,N_27928,N_27708);
or U28429 (N_28429,N_27332,N_27384);
nor U28430 (N_28430,N_27577,N_27631);
nor U28431 (N_28431,N_27121,N_27973);
or U28432 (N_28432,N_27351,N_27095);
xnor U28433 (N_28433,N_27474,N_27281);
or U28434 (N_28434,N_27511,N_27147);
nor U28435 (N_28435,N_27827,N_27497);
nand U28436 (N_28436,N_27495,N_27068);
nor U28437 (N_28437,N_27878,N_27377);
or U28438 (N_28438,N_27418,N_27871);
xnor U28439 (N_28439,N_27098,N_27144);
and U28440 (N_28440,N_27423,N_27174);
nand U28441 (N_28441,N_27318,N_27675);
nand U28442 (N_28442,N_27611,N_27852);
or U28443 (N_28443,N_27192,N_27736);
or U28444 (N_28444,N_27465,N_27913);
nand U28445 (N_28445,N_27905,N_27606);
or U28446 (N_28446,N_27275,N_27615);
xnor U28447 (N_28447,N_27686,N_27480);
xnor U28448 (N_28448,N_27359,N_27273);
nor U28449 (N_28449,N_27405,N_27869);
nor U28450 (N_28450,N_27456,N_27720);
and U28451 (N_28451,N_27528,N_27895);
xnor U28452 (N_28452,N_27397,N_27796);
nand U28453 (N_28453,N_27309,N_27946);
nor U28454 (N_28454,N_27727,N_27722);
nand U28455 (N_28455,N_27394,N_27201);
or U28456 (N_28456,N_27485,N_27321);
nand U28457 (N_28457,N_27651,N_27643);
and U28458 (N_28458,N_27034,N_27319);
xor U28459 (N_28459,N_27728,N_27238);
xor U28460 (N_28460,N_27724,N_27937);
nand U28461 (N_28461,N_27602,N_27901);
nand U28462 (N_28462,N_27228,N_27809);
nor U28463 (N_28463,N_27011,N_27941);
nor U28464 (N_28464,N_27540,N_27875);
xor U28465 (N_28465,N_27404,N_27620);
xnor U28466 (N_28466,N_27438,N_27792);
nor U28467 (N_28467,N_27628,N_27149);
xor U28468 (N_28468,N_27043,N_27463);
nor U28469 (N_28469,N_27530,N_27389);
or U28470 (N_28470,N_27668,N_27551);
and U28471 (N_28471,N_27757,N_27303);
or U28472 (N_28472,N_27427,N_27243);
nor U28473 (N_28473,N_27077,N_27596);
nor U28474 (N_28474,N_27138,N_27127);
and U28475 (N_28475,N_27948,N_27367);
nor U28476 (N_28476,N_27107,N_27212);
nand U28477 (N_28477,N_27124,N_27085);
nand U28478 (N_28478,N_27965,N_27833);
nand U28479 (N_28479,N_27145,N_27294);
xnor U28480 (N_28480,N_27267,N_27213);
or U28481 (N_28481,N_27751,N_27237);
or U28482 (N_28482,N_27478,N_27128);
nor U28483 (N_28483,N_27590,N_27738);
and U28484 (N_28484,N_27005,N_27096);
or U28485 (N_28485,N_27758,N_27844);
nor U28486 (N_28486,N_27426,N_27840);
xnor U28487 (N_28487,N_27917,N_27592);
and U28488 (N_28488,N_27482,N_27619);
and U28489 (N_28489,N_27744,N_27113);
and U28490 (N_28490,N_27216,N_27910);
and U28491 (N_28491,N_27652,N_27848);
or U28492 (N_28492,N_27499,N_27806);
or U28493 (N_28493,N_27087,N_27052);
xor U28494 (N_28494,N_27437,N_27327);
and U28495 (N_28495,N_27718,N_27089);
xnor U28496 (N_28496,N_27291,N_27521);
xor U28497 (N_28497,N_27168,N_27097);
or U28498 (N_28498,N_27983,N_27754);
and U28499 (N_28499,N_27072,N_27091);
nand U28500 (N_28500,N_27484,N_27175);
or U28501 (N_28501,N_27345,N_27627);
xor U28502 (N_28502,N_27411,N_27064);
nor U28503 (N_28503,N_27781,N_27101);
and U28504 (N_28504,N_27261,N_27353);
xnor U28505 (N_28505,N_27647,N_27588);
xnor U28506 (N_28506,N_27378,N_27359);
or U28507 (N_28507,N_27729,N_27088);
nor U28508 (N_28508,N_27237,N_27995);
or U28509 (N_28509,N_27694,N_27624);
nand U28510 (N_28510,N_27751,N_27415);
and U28511 (N_28511,N_27082,N_27661);
and U28512 (N_28512,N_27042,N_27493);
nand U28513 (N_28513,N_27549,N_27314);
nor U28514 (N_28514,N_27260,N_27411);
and U28515 (N_28515,N_27029,N_27707);
or U28516 (N_28516,N_27952,N_27860);
or U28517 (N_28517,N_27534,N_27084);
nor U28518 (N_28518,N_27991,N_27121);
nor U28519 (N_28519,N_27412,N_27134);
and U28520 (N_28520,N_27100,N_27946);
or U28521 (N_28521,N_27718,N_27920);
nor U28522 (N_28522,N_27908,N_27885);
and U28523 (N_28523,N_27477,N_27493);
and U28524 (N_28524,N_27549,N_27815);
nand U28525 (N_28525,N_27433,N_27784);
nand U28526 (N_28526,N_27629,N_27488);
xor U28527 (N_28527,N_27878,N_27271);
xnor U28528 (N_28528,N_27575,N_27168);
or U28529 (N_28529,N_27795,N_27385);
and U28530 (N_28530,N_27189,N_27996);
nor U28531 (N_28531,N_27521,N_27078);
nor U28532 (N_28532,N_27854,N_27137);
nand U28533 (N_28533,N_27615,N_27957);
nor U28534 (N_28534,N_27210,N_27245);
and U28535 (N_28535,N_27481,N_27600);
xor U28536 (N_28536,N_27073,N_27576);
xnor U28537 (N_28537,N_27550,N_27218);
nand U28538 (N_28538,N_27631,N_27090);
nor U28539 (N_28539,N_27166,N_27602);
or U28540 (N_28540,N_27829,N_27352);
xor U28541 (N_28541,N_27601,N_27976);
and U28542 (N_28542,N_27983,N_27664);
and U28543 (N_28543,N_27970,N_27801);
and U28544 (N_28544,N_27651,N_27183);
and U28545 (N_28545,N_27185,N_27832);
nand U28546 (N_28546,N_27812,N_27567);
nor U28547 (N_28547,N_27147,N_27024);
xnor U28548 (N_28548,N_27698,N_27645);
and U28549 (N_28549,N_27792,N_27767);
nand U28550 (N_28550,N_27807,N_27542);
nor U28551 (N_28551,N_27584,N_27775);
xnor U28552 (N_28552,N_27346,N_27420);
xor U28553 (N_28553,N_27463,N_27487);
nand U28554 (N_28554,N_27087,N_27836);
and U28555 (N_28555,N_27554,N_27792);
nor U28556 (N_28556,N_27935,N_27065);
nand U28557 (N_28557,N_27584,N_27656);
xor U28558 (N_28558,N_27845,N_27244);
xor U28559 (N_28559,N_27763,N_27773);
nor U28560 (N_28560,N_27259,N_27903);
xnor U28561 (N_28561,N_27137,N_27142);
xor U28562 (N_28562,N_27020,N_27676);
and U28563 (N_28563,N_27002,N_27121);
and U28564 (N_28564,N_27486,N_27733);
nand U28565 (N_28565,N_27626,N_27933);
nand U28566 (N_28566,N_27502,N_27467);
or U28567 (N_28567,N_27163,N_27323);
nor U28568 (N_28568,N_27641,N_27104);
xor U28569 (N_28569,N_27546,N_27115);
or U28570 (N_28570,N_27440,N_27014);
xor U28571 (N_28571,N_27134,N_27919);
nor U28572 (N_28572,N_27747,N_27204);
and U28573 (N_28573,N_27090,N_27528);
or U28574 (N_28574,N_27089,N_27598);
or U28575 (N_28575,N_27354,N_27957);
or U28576 (N_28576,N_27576,N_27773);
and U28577 (N_28577,N_27102,N_27407);
or U28578 (N_28578,N_27047,N_27243);
nor U28579 (N_28579,N_27284,N_27094);
and U28580 (N_28580,N_27565,N_27881);
or U28581 (N_28581,N_27461,N_27811);
xnor U28582 (N_28582,N_27425,N_27320);
and U28583 (N_28583,N_27953,N_27576);
or U28584 (N_28584,N_27121,N_27131);
and U28585 (N_28585,N_27129,N_27501);
xor U28586 (N_28586,N_27138,N_27424);
xnor U28587 (N_28587,N_27780,N_27078);
nor U28588 (N_28588,N_27840,N_27702);
nand U28589 (N_28589,N_27208,N_27035);
nor U28590 (N_28590,N_27372,N_27892);
and U28591 (N_28591,N_27538,N_27371);
nand U28592 (N_28592,N_27743,N_27452);
nand U28593 (N_28593,N_27931,N_27793);
nand U28594 (N_28594,N_27636,N_27736);
nor U28595 (N_28595,N_27336,N_27697);
xnor U28596 (N_28596,N_27591,N_27120);
nor U28597 (N_28597,N_27263,N_27240);
xor U28598 (N_28598,N_27061,N_27980);
nand U28599 (N_28599,N_27234,N_27046);
or U28600 (N_28600,N_27383,N_27432);
or U28601 (N_28601,N_27730,N_27440);
and U28602 (N_28602,N_27017,N_27884);
nor U28603 (N_28603,N_27114,N_27248);
and U28604 (N_28604,N_27317,N_27887);
and U28605 (N_28605,N_27105,N_27150);
nor U28606 (N_28606,N_27802,N_27764);
or U28607 (N_28607,N_27315,N_27165);
or U28608 (N_28608,N_27228,N_27579);
nand U28609 (N_28609,N_27769,N_27715);
and U28610 (N_28610,N_27672,N_27994);
nor U28611 (N_28611,N_27825,N_27093);
nor U28612 (N_28612,N_27731,N_27757);
or U28613 (N_28613,N_27691,N_27996);
or U28614 (N_28614,N_27979,N_27966);
and U28615 (N_28615,N_27738,N_27628);
or U28616 (N_28616,N_27435,N_27471);
or U28617 (N_28617,N_27195,N_27571);
and U28618 (N_28618,N_27839,N_27046);
and U28619 (N_28619,N_27418,N_27394);
nand U28620 (N_28620,N_27824,N_27698);
and U28621 (N_28621,N_27435,N_27206);
or U28622 (N_28622,N_27693,N_27769);
xor U28623 (N_28623,N_27589,N_27588);
or U28624 (N_28624,N_27805,N_27045);
nand U28625 (N_28625,N_27863,N_27672);
or U28626 (N_28626,N_27617,N_27177);
xnor U28627 (N_28627,N_27017,N_27261);
or U28628 (N_28628,N_27417,N_27878);
nand U28629 (N_28629,N_27637,N_27282);
nand U28630 (N_28630,N_27745,N_27849);
nor U28631 (N_28631,N_27591,N_27140);
nand U28632 (N_28632,N_27251,N_27567);
nand U28633 (N_28633,N_27828,N_27848);
nand U28634 (N_28634,N_27497,N_27312);
or U28635 (N_28635,N_27927,N_27021);
xor U28636 (N_28636,N_27835,N_27544);
nor U28637 (N_28637,N_27949,N_27834);
nand U28638 (N_28638,N_27152,N_27682);
or U28639 (N_28639,N_27425,N_27532);
and U28640 (N_28640,N_27698,N_27756);
nand U28641 (N_28641,N_27857,N_27416);
or U28642 (N_28642,N_27400,N_27125);
nor U28643 (N_28643,N_27214,N_27101);
xnor U28644 (N_28644,N_27352,N_27037);
nand U28645 (N_28645,N_27309,N_27335);
nand U28646 (N_28646,N_27930,N_27554);
xor U28647 (N_28647,N_27479,N_27805);
nand U28648 (N_28648,N_27667,N_27399);
and U28649 (N_28649,N_27120,N_27704);
or U28650 (N_28650,N_27066,N_27132);
or U28651 (N_28651,N_27458,N_27457);
nor U28652 (N_28652,N_27407,N_27254);
nand U28653 (N_28653,N_27493,N_27081);
xor U28654 (N_28654,N_27238,N_27891);
and U28655 (N_28655,N_27571,N_27438);
and U28656 (N_28656,N_27705,N_27669);
xor U28657 (N_28657,N_27433,N_27214);
xnor U28658 (N_28658,N_27629,N_27158);
xor U28659 (N_28659,N_27355,N_27514);
nor U28660 (N_28660,N_27967,N_27425);
nand U28661 (N_28661,N_27279,N_27876);
nor U28662 (N_28662,N_27585,N_27459);
and U28663 (N_28663,N_27077,N_27727);
xor U28664 (N_28664,N_27237,N_27469);
xor U28665 (N_28665,N_27255,N_27109);
and U28666 (N_28666,N_27490,N_27281);
nor U28667 (N_28667,N_27792,N_27779);
xnor U28668 (N_28668,N_27837,N_27381);
or U28669 (N_28669,N_27519,N_27342);
xnor U28670 (N_28670,N_27966,N_27249);
nand U28671 (N_28671,N_27431,N_27768);
nand U28672 (N_28672,N_27791,N_27357);
or U28673 (N_28673,N_27066,N_27903);
or U28674 (N_28674,N_27903,N_27979);
nand U28675 (N_28675,N_27204,N_27517);
or U28676 (N_28676,N_27533,N_27550);
and U28677 (N_28677,N_27115,N_27388);
or U28678 (N_28678,N_27772,N_27456);
and U28679 (N_28679,N_27610,N_27513);
nand U28680 (N_28680,N_27900,N_27453);
or U28681 (N_28681,N_27239,N_27487);
nand U28682 (N_28682,N_27938,N_27990);
and U28683 (N_28683,N_27906,N_27108);
xnor U28684 (N_28684,N_27122,N_27132);
nor U28685 (N_28685,N_27105,N_27129);
nor U28686 (N_28686,N_27206,N_27306);
and U28687 (N_28687,N_27013,N_27537);
or U28688 (N_28688,N_27473,N_27972);
or U28689 (N_28689,N_27483,N_27477);
and U28690 (N_28690,N_27498,N_27191);
xor U28691 (N_28691,N_27910,N_27115);
nand U28692 (N_28692,N_27534,N_27100);
nor U28693 (N_28693,N_27781,N_27435);
xnor U28694 (N_28694,N_27581,N_27465);
xnor U28695 (N_28695,N_27217,N_27708);
and U28696 (N_28696,N_27723,N_27704);
and U28697 (N_28697,N_27526,N_27966);
and U28698 (N_28698,N_27425,N_27406);
nor U28699 (N_28699,N_27068,N_27735);
xnor U28700 (N_28700,N_27047,N_27476);
or U28701 (N_28701,N_27279,N_27154);
xor U28702 (N_28702,N_27064,N_27740);
xnor U28703 (N_28703,N_27519,N_27128);
nor U28704 (N_28704,N_27032,N_27931);
nand U28705 (N_28705,N_27466,N_27778);
nand U28706 (N_28706,N_27542,N_27361);
xnor U28707 (N_28707,N_27090,N_27987);
or U28708 (N_28708,N_27693,N_27723);
nand U28709 (N_28709,N_27827,N_27728);
xor U28710 (N_28710,N_27245,N_27979);
and U28711 (N_28711,N_27639,N_27490);
and U28712 (N_28712,N_27544,N_27565);
nor U28713 (N_28713,N_27392,N_27182);
nand U28714 (N_28714,N_27876,N_27570);
nor U28715 (N_28715,N_27789,N_27768);
or U28716 (N_28716,N_27033,N_27591);
nand U28717 (N_28717,N_27921,N_27417);
and U28718 (N_28718,N_27719,N_27635);
and U28719 (N_28719,N_27124,N_27262);
nor U28720 (N_28720,N_27264,N_27412);
and U28721 (N_28721,N_27692,N_27559);
and U28722 (N_28722,N_27744,N_27536);
and U28723 (N_28723,N_27843,N_27813);
or U28724 (N_28724,N_27430,N_27613);
and U28725 (N_28725,N_27004,N_27935);
nor U28726 (N_28726,N_27893,N_27082);
nor U28727 (N_28727,N_27848,N_27479);
or U28728 (N_28728,N_27617,N_27259);
xor U28729 (N_28729,N_27104,N_27000);
xor U28730 (N_28730,N_27066,N_27740);
nand U28731 (N_28731,N_27415,N_27563);
and U28732 (N_28732,N_27497,N_27125);
nor U28733 (N_28733,N_27332,N_27007);
xnor U28734 (N_28734,N_27829,N_27102);
and U28735 (N_28735,N_27059,N_27477);
and U28736 (N_28736,N_27093,N_27648);
xor U28737 (N_28737,N_27436,N_27680);
nand U28738 (N_28738,N_27414,N_27246);
or U28739 (N_28739,N_27742,N_27927);
and U28740 (N_28740,N_27673,N_27788);
and U28741 (N_28741,N_27659,N_27643);
nand U28742 (N_28742,N_27230,N_27822);
and U28743 (N_28743,N_27138,N_27246);
or U28744 (N_28744,N_27590,N_27803);
nor U28745 (N_28745,N_27332,N_27708);
or U28746 (N_28746,N_27699,N_27682);
nand U28747 (N_28747,N_27995,N_27062);
nor U28748 (N_28748,N_27959,N_27787);
nand U28749 (N_28749,N_27642,N_27007);
nand U28750 (N_28750,N_27016,N_27134);
and U28751 (N_28751,N_27385,N_27332);
nand U28752 (N_28752,N_27249,N_27744);
nor U28753 (N_28753,N_27210,N_27783);
or U28754 (N_28754,N_27560,N_27436);
nand U28755 (N_28755,N_27531,N_27294);
xnor U28756 (N_28756,N_27165,N_27119);
xnor U28757 (N_28757,N_27023,N_27942);
and U28758 (N_28758,N_27744,N_27118);
nand U28759 (N_28759,N_27155,N_27308);
nor U28760 (N_28760,N_27895,N_27976);
nand U28761 (N_28761,N_27311,N_27806);
xnor U28762 (N_28762,N_27578,N_27652);
xor U28763 (N_28763,N_27741,N_27956);
or U28764 (N_28764,N_27385,N_27645);
nor U28765 (N_28765,N_27706,N_27956);
nand U28766 (N_28766,N_27362,N_27704);
nor U28767 (N_28767,N_27836,N_27196);
nand U28768 (N_28768,N_27780,N_27566);
nand U28769 (N_28769,N_27284,N_27147);
or U28770 (N_28770,N_27542,N_27674);
nand U28771 (N_28771,N_27763,N_27957);
and U28772 (N_28772,N_27717,N_27032);
xnor U28773 (N_28773,N_27965,N_27666);
nand U28774 (N_28774,N_27972,N_27127);
nor U28775 (N_28775,N_27627,N_27252);
xor U28776 (N_28776,N_27049,N_27247);
nand U28777 (N_28777,N_27515,N_27669);
or U28778 (N_28778,N_27617,N_27857);
nor U28779 (N_28779,N_27186,N_27696);
nor U28780 (N_28780,N_27592,N_27879);
xnor U28781 (N_28781,N_27506,N_27796);
and U28782 (N_28782,N_27449,N_27507);
xor U28783 (N_28783,N_27574,N_27887);
nand U28784 (N_28784,N_27759,N_27281);
nor U28785 (N_28785,N_27563,N_27970);
and U28786 (N_28786,N_27163,N_27609);
nand U28787 (N_28787,N_27308,N_27853);
and U28788 (N_28788,N_27123,N_27413);
or U28789 (N_28789,N_27991,N_27704);
and U28790 (N_28790,N_27666,N_27664);
nor U28791 (N_28791,N_27676,N_27224);
nor U28792 (N_28792,N_27929,N_27865);
and U28793 (N_28793,N_27900,N_27791);
xor U28794 (N_28794,N_27905,N_27951);
and U28795 (N_28795,N_27942,N_27821);
nor U28796 (N_28796,N_27284,N_27919);
xnor U28797 (N_28797,N_27689,N_27400);
nand U28798 (N_28798,N_27248,N_27358);
nand U28799 (N_28799,N_27870,N_27631);
xor U28800 (N_28800,N_27450,N_27911);
nor U28801 (N_28801,N_27282,N_27387);
xnor U28802 (N_28802,N_27630,N_27296);
nor U28803 (N_28803,N_27046,N_27490);
nor U28804 (N_28804,N_27515,N_27183);
xnor U28805 (N_28805,N_27429,N_27342);
and U28806 (N_28806,N_27610,N_27643);
nand U28807 (N_28807,N_27495,N_27281);
nand U28808 (N_28808,N_27361,N_27992);
nand U28809 (N_28809,N_27742,N_27576);
xnor U28810 (N_28810,N_27345,N_27311);
or U28811 (N_28811,N_27065,N_27652);
xor U28812 (N_28812,N_27728,N_27546);
or U28813 (N_28813,N_27205,N_27963);
nor U28814 (N_28814,N_27889,N_27817);
nor U28815 (N_28815,N_27497,N_27169);
nor U28816 (N_28816,N_27946,N_27902);
or U28817 (N_28817,N_27657,N_27762);
or U28818 (N_28818,N_27333,N_27297);
nand U28819 (N_28819,N_27544,N_27993);
or U28820 (N_28820,N_27589,N_27437);
and U28821 (N_28821,N_27707,N_27692);
and U28822 (N_28822,N_27160,N_27180);
xor U28823 (N_28823,N_27993,N_27659);
nand U28824 (N_28824,N_27862,N_27066);
nor U28825 (N_28825,N_27752,N_27487);
or U28826 (N_28826,N_27651,N_27764);
nand U28827 (N_28827,N_27828,N_27586);
xor U28828 (N_28828,N_27599,N_27537);
and U28829 (N_28829,N_27437,N_27307);
xor U28830 (N_28830,N_27664,N_27692);
and U28831 (N_28831,N_27859,N_27681);
xor U28832 (N_28832,N_27934,N_27246);
xor U28833 (N_28833,N_27409,N_27228);
xor U28834 (N_28834,N_27198,N_27331);
nor U28835 (N_28835,N_27717,N_27183);
and U28836 (N_28836,N_27732,N_27818);
and U28837 (N_28837,N_27752,N_27500);
nand U28838 (N_28838,N_27918,N_27823);
nand U28839 (N_28839,N_27385,N_27915);
nand U28840 (N_28840,N_27694,N_27060);
and U28841 (N_28841,N_27472,N_27860);
xnor U28842 (N_28842,N_27480,N_27872);
xnor U28843 (N_28843,N_27648,N_27213);
nor U28844 (N_28844,N_27094,N_27080);
and U28845 (N_28845,N_27471,N_27461);
and U28846 (N_28846,N_27393,N_27657);
or U28847 (N_28847,N_27067,N_27453);
and U28848 (N_28848,N_27380,N_27170);
nand U28849 (N_28849,N_27257,N_27293);
nand U28850 (N_28850,N_27038,N_27338);
nor U28851 (N_28851,N_27514,N_27311);
and U28852 (N_28852,N_27983,N_27049);
nor U28853 (N_28853,N_27640,N_27032);
xor U28854 (N_28854,N_27277,N_27593);
and U28855 (N_28855,N_27771,N_27423);
nor U28856 (N_28856,N_27407,N_27670);
xor U28857 (N_28857,N_27956,N_27459);
xnor U28858 (N_28858,N_27485,N_27314);
or U28859 (N_28859,N_27015,N_27705);
xor U28860 (N_28860,N_27917,N_27948);
nand U28861 (N_28861,N_27486,N_27658);
and U28862 (N_28862,N_27093,N_27718);
and U28863 (N_28863,N_27908,N_27662);
xor U28864 (N_28864,N_27747,N_27408);
or U28865 (N_28865,N_27323,N_27905);
or U28866 (N_28866,N_27975,N_27022);
or U28867 (N_28867,N_27854,N_27729);
or U28868 (N_28868,N_27994,N_27037);
and U28869 (N_28869,N_27102,N_27139);
and U28870 (N_28870,N_27891,N_27225);
or U28871 (N_28871,N_27330,N_27145);
nor U28872 (N_28872,N_27912,N_27590);
xor U28873 (N_28873,N_27668,N_27270);
or U28874 (N_28874,N_27865,N_27302);
xnor U28875 (N_28875,N_27136,N_27957);
nor U28876 (N_28876,N_27125,N_27666);
or U28877 (N_28877,N_27327,N_27723);
nor U28878 (N_28878,N_27747,N_27017);
or U28879 (N_28879,N_27874,N_27887);
and U28880 (N_28880,N_27034,N_27148);
nand U28881 (N_28881,N_27780,N_27933);
and U28882 (N_28882,N_27211,N_27959);
xor U28883 (N_28883,N_27498,N_27647);
and U28884 (N_28884,N_27596,N_27221);
nor U28885 (N_28885,N_27729,N_27565);
and U28886 (N_28886,N_27487,N_27210);
xor U28887 (N_28887,N_27932,N_27173);
nand U28888 (N_28888,N_27731,N_27162);
xnor U28889 (N_28889,N_27796,N_27724);
xnor U28890 (N_28890,N_27508,N_27680);
nor U28891 (N_28891,N_27405,N_27004);
nand U28892 (N_28892,N_27814,N_27539);
and U28893 (N_28893,N_27637,N_27145);
xnor U28894 (N_28894,N_27804,N_27900);
nor U28895 (N_28895,N_27329,N_27536);
and U28896 (N_28896,N_27529,N_27837);
nor U28897 (N_28897,N_27199,N_27422);
or U28898 (N_28898,N_27950,N_27616);
or U28899 (N_28899,N_27799,N_27275);
nor U28900 (N_28900,N_27332,N_27548);
or U28901 (N_28901,N_27666,N_27917);
or U28902 (N_28902,N_27898,N_27175);
or U28903 (N_28903,N_27262,N_27641);
xnor U28904 (N_28904,N_27222,N_27822);
nor U28905 (N_28905,N_27997,N_27804);
or U28906 (N_28906,N_27808,N_27501);
nand U28907 (N_28907,N_27064,N_27159);
and U28908 (N_28908,N_27715,N_27706);
and U28909 (N_28909,N_27207,N_27301);
nor U28910 (N_28910,N_27251,N_27171);
and U28911 (N_28911,N_27632,N_27411);
xnor U28912 (N_28912,N_27421,N_27933);
xnor U28913 (N_28913,N_27950,N_27977);
xnor U28914 (N_28914,N_27277,N_27721);
and U28915 (N_28915,N_27316,N_27151);
nor U28916 (N_28916,N_27666,N_27629);
nand U28917 (N_28917,N_27327,N_27876);
and U28918 (N_28918,N_27103,N_27059);
nand U28919 (N_28919,N_27330,N_27636);
or U28920 (N_28920,N_27294,N_27669);
xor U28921 (N_28921,N_27785,N_27037);
xor U28922 (N_28922,N_27984,N_27138);
and U28923 (N_28923,N_27868,N_27844);
nor U28924 (N_28924,N_27459,N_27544);
and U28925 (N_28925,N_27990,N_27107);
or U28926 (N_28926,N_27313,N_27132);
or U28927 (N_28927,N_27441,N_27828);
and U28928 (N_28928,N_27062,N_27163);
nand U28929 (N_28929,N_27992,N_27531);
nor U28930 (N_28930,N_27509,N_27021);
xnor U28931 (N_28931,N_27546,N_27859);
nor U28932 (N_28932,N_27173,N_27885);
nand U28933 (N_28933,N_27574,N_27900);
nand U28934 (N_28934,N_27454,N_27125);
and U28935 (N_28935,N_27562,N_27865);
or U28936 (N_28936,N_27888,N_27677);
nor U28937 (N_28937,N_27304,N_27846);
xor U28938 (N_28938,N_27900,N_27273);
and U28939 (N_28939,N_27908,N_27111);
and U28940 (N_28940,N_27999,N_27292);
or U28941 (N_28941,N_27389,N_27317);
or U28942 (N_28942,N_27556,N_27718);
xor U28943 (N_28943,N_27047,N_27262);
nand U28944 (N_28944,N_27248,N_27557);
and U28945 (N_28945,N_27739,N_27535);
nand U28946 (N_28946,N_27294,N_27419);
nor U28947 (N_28947,N_27001,N_27857);
nor U28948 (N_28948,N_27998,N_27006);
or U28949 (N_28949,N_27453,N_27106);
or U28950 (N_28950,N_27190,N_27959);
and U28951 (N_28951,N_27929,N_27357);
nor U28952 (N_28952,N_27336,N_27532);
nor U28953 (N_28953,N_27667,N_27646);
or U28954 (N_28954,N_27828,N_27220);
or U28955 (N_28955,N_27846,N_27400);
nand U28956 (N_28956,N_27932,N_27748);
nor U28957 (N_28957,N_27340,N_27518);
xor U28958 (N_28958,N_27755,N_27398);
or U28959 (N_28959,N_27733,N_27242);
nand U28960 (N_28960,N_27908,N_27824);
nand U28961 (N_28961,N_27626,N_27904);
nand U28962 (N_28962,N_27491,N_27461);
or U28963 (N_28963,N_27695,N_27303);
nand U28964 (N_28964,N_27898,N_27591);
and U28965 (N_28965,N_27079,N_27236);
nor U28966 (N_28966,N_27626,N_27201);
nor U28967 (N_28967,N_27964,N_27674);
or U28968 (N_28968,N_27109,N_27620);
xnor U28969 (N_28969,N_27714,N_27274);
nand U28970 (N_28970,N_27132,N_27451);
nand U28971 (N_28971,N_27960,N_27674);
nand U28972 (N_28972,N_27056,N_27956);
xor U28973 (N_28973,N_27440,N_27967);
and U28974 (N_28974,N_27783,N_27740);
nor U28975 (N_28975,N_27800,N_27996);
xor U28976 (N_28976,N_27033,N_27602);
nand U28977 (N_28977,N_27017,N_27684);
nor U28978 (N_28978,N_27586,N_27018);
or U28979 (N_28979,N_27644,N_27241);
nand U28980 (N_28980,N_27280,N_27394);
nor U28981 (N_28981,N_27025,N_27993);
nand U28982 (N_28982,N_27862,N_27642);
nand U28983 (N_28983,N_27136,N_27162);
xor U28984 (N_28984,N_27127,N_27242);
or U28985 (N_28985,N_27935,N_27999);
xnor U28986 (N_28986,N_27085,N_27416);
nor U28987 (N_28987,N_27833,N_27452);
nand U28988 (N_28988,N_27595,N_27558);
nor U28989 (N_28989,N_27063,N_27833);
nand U28990 (N_28990,N_27969,N_27875);
nand U28991 (N_28991,N_27740,N_27302);
nor U28992 (N_28992,N_27061,N_27568);
nor U28993 (N_28993,N_27867,N_27763);
and U28994 (N_28994,N_27460,N_27759);
and U28995 (N_28995,N_27948,N_27128);
nor U28996 (N_28996,N_27609,N_27839);
xor U28997 (N_28997,N_27079,N_27128);
nand U28998 (N_28998,N_27916,N_27228);
and U28999 (N_28999,N_27964,N_27396);
xor U29000 (N_29000,N_28017,N_28456);
nor U29001 (N_29001,N_28149,N_28040);
or U29002 (N_29002,N_28649,N_28144);
nor U29003 (N_29003,N_28642,N_28795);
nor U29004 (N_29004,N_28091,N_28305);
xor U29005 (N_29005,N_28001,N_28662);
and U29006 (N_29006,N_28468,N_28831);
xnor U29007 (N_29007,N_28690,N_28217);
xor U29008 (N_29008,N_28765,N_28242);
nor U29009 (N_29009,N_28413,N_28119);
nor U29010 (N_29010,N_28757,N_28820);
nand U29011 (N_29011,N_28044,N_28279);
and U29012 (N_29012,N_28483,N_28889);
nand U29013 (N_29013,N_28449,N_28902);
nor U29014 (N_29014,N_28750,N_28373);
nor U29015 (N_29015,N_28879,N_28367);
nand U29016 (N_29016,N_28937,N_28725);
nor U29017 (N_29017,N_28997,N_28743);
nand U29018 (N_29018,N_28385,N_28768);
nand U29019 (N_29019,N_28507,N_28543);
nand U29020 (N_29020,N_28633,N_28846);
nor U29021 (N_29021,N_28362,N_28695);
xnor U29022 (N_29022,N_28460,N_28288);
xnor U29023 (N_29023,N_28450,N_28090);
nor U29024 (N_29024,N_28262,N_28297);
or U29025 (N_29025,N_28307,N_28710);
nand U29026 (N_29026,N_28587,N_28230);
nor U29027 (N_29027,N_28303,N_28542);
or U29028 (N_29028,N_28920,N_28799);
nor U29029 (N_29029,N_28766,N_28216);
xor U29030 (N_29030,N_28443,N_28667);
and U29031 (N_29031,N_28065,N_28479);
and U29032 (N_29032,N_28179,N_28722);
nand U29033 (N_29033,N_28513,N_28595);
nand U29034 (N_29034,N_28323,N_28210);
or U29035 (N_29035,N_28068,N_28211);
xnor U29036 (N_29036,N_28576,N_28173);
nand U29037 (N_29037,N_28239,N_28036);
or U29038 (N_29038,N_28448,N_28337);
nor U29039 (N_29039,N_28097,N_28165);
nor U29040 (N_29040,N_28635,N_28559);
nand U29041 (N_29041,N_28991,N_28704);
and U29042 (N_29042,N_28347,N_28356);
and U29043 (N_29043,N_28907,N_28045);
or U29044 (N_29044,N_28678,N_28838);
xnor U29045 (N_29045,N_28687,N_28209);
or U29046 (N_29046,N_28748,N_28284);
or U29047 (N_29047,N_28258,N_28266);
and U29048 (N_29048,N_28594,N_28478);
and U29049 (N_29049,N_28446,N_28011);
xnor U29050 (N_29050,N_28095,N_28291);
xnor U29051 (N_29051,N_28277,N_28379);
nand U29052 (N_29052,N_28228,N_28653);
and U29053 (N_29053,N_28380,N_28520);
or U29054 (N_29054,N_28548,N_28160);
nor U29055 (N_29055,N_28490,N_28968);
nor U29056 (N_29056,N_28663,N_28855);
xnor U29057 (N_29057,N_28213,N_28295);
nand U29058 (N_29058,N_28453,N_28661);
and U29059 (N_29059,N_28959,N_28572);
and U29060 (N_29060,N_28568,N_28925);
nor U29061 (N_29061,N_28703,N_28618);
or U29062 (N_29062,N_28116,N_28694);
xor U29063 (N_29063,N_28523,N_28797);
or U29064 (N_29064,N_28192,N_28943);
nor U29065 (N_29065,N_28714,N_28254);
nor U29066 (N_29066,N_28016,N_28923);
nand U29067 (N_29067,N_28330,N_28252);
or U29068 (N_29068,N_28940,N_28175);
nor U29069 (N_29069,N_28405,N_28030);
xor U29070 (N_29070,N_28600,N_28958);
or U29071 (N_29071,N_28432,N_28435);
and U29072 (N_29072,N_28391,N_28382);
or U29073 (N_29073,N_28359,N_28221);
nand U29074 (N_29074,N_28904,N_28790);
xor U29075 (N_29075,N_28880,N_28628);
nor U29076 (N_29076,N_28128,N_28070);
or U29077 (N_29077,N_28234,N_28939);
nor U29078 (N_29078,N_28951,N_28801);
and U29079 (N_29079,N_28871,N_28434);
and U29080 (N_29080,N_28538,N_28433);
nor U29081 (N_29081,N_28321,N_28220);
and U29082 (N_29082,N_28477,N_28194);
nor U29083 (N_29083,N_28643,N_28806);
xnor U29084 (N_29084,N_28821,N_28418);
and U29085 (N_29085,N_28229,N_28668);
or U29086 (N_29086,N_28199,N_28584);
or U29087 (N_29087,N_28028,N_28426);
or U29088 (N_29088,N_28047,N_28143);
xor U29089 (N_29089,N_28488,N_28440);
nor U29090 (N_29090,N_28980,N_28280);
or U29091 (N_29091,N_28203,N_28816);
xnor U29092 (N_29092,N_28464,N_28058);
and U29093 (N_29093,N_28341,N_28121);
xor U29094 (N_29094,N_28749,N_28112);
or U29095 (N_29095,N_28412,N_28442);
nand U29096 (N_29096,N_28161,N_28073);
nand U29097 (N_29097,N_28961,N_28499);
xnor U29098 (N_29098,N_28334,N_28540);
and U29099 (N_29099,N_28053,N_28616);
xnor U29100 (N_29100,N_28527,N_28098);
and U29101 (N_29101,N_28076,N_28004);
nor U29102 (N_29102,N_28086,N_28832);
nand U29103 (N_29103,N_28979,N_28569);
and U29104 (N_29104,N_28934,N_28567);
xor U29105 (N_29105,N_28914,N_28580);
and U29106 (N_29106,N_28311,N_28401);
nand U29107 (N_29107,N_28952,N_28894);
xor U29108 (N_29108,N_28500,N_28287);
and U29109 (N_29109,N_28172,N_28219);
xor U29110 (N_29110,N_28973,N_28746);
nand U29111 (N_29111,N_28593,N_28544);
and U29112 (N_29112,N_28985,N_28241);
nor U29113 (N_29113,N_28787,N_28555);
xnor U29114 (N_29114,N_28530,N_28429);
nor U29115 (N_29115,N_28808,N_28636);
nand U29116 (N_29116,N_28942,N_28897);
nand U29117 (N_29117,N_28759,N_28273);
nand U29118 (N_29118,N_28899,N_28737);
xnor U29119 (N_29119,N_28551,N_28982);
and U29120 (N_29120,N_28471,N_28320);
nor U29121 (N_29121,N_28463,N_28487);
and U29122 (N_29122,N_28532,N_28726);
nor U29123 (N_29123,N_28993,N_28769);
or U29124 (N_29124,N_28105,N_28908);
and U29125 (N_29125,N_28676,N_28627);
xor U29126 (N_29126,N_28840,N_28340);
nand U29127 (N_29127,N_28778,N_28553);
and U29128 (N_29128,N_28510,N_28657);
xor U29129 (N_29129,N_28240,N_28718);
and U29130 (N_29130,N_28854,N_28949);
nor U29131 (N_29131,N_28163,N_28850);
or U29132 (N_29132,N_28461,N_28884);
nand U29133 (N_29133,N_28779,N_28550);
nor U29134 (N_29134,N_28866,N_28802);
or U29135 (N_29135,N_28462,N_28063);
nor U29136 (N_29136,N_28706,N_28204);
nor U29137 (N_29137,N_28995,N_28604);
nor U29138 (N_29138,N_28729,N_28422);
nor U29139 (N_29139,N_28767,N_28954);
and U29140 (N_29140,N_28862,N_28794);
nor U29141 (N_29141,N_28132,N_28868);
xnor U29142 (N_29142,N_28282,N_28411);
nor U29143 (N_29143,N_28989,N_28827);
xor U29144 (N_29144,N_28648,N_28717);
and U29145 (N_29145,N_28976,N_28579);
nor U29146 (N_29146,N_28005,N_28339);
or U29147 (N_29147,N_28508,N_28384);
xnor U29148 (N_29148,N_28275,N_28823);
nor U29149 (N_29149,N_28589,N_28296);
xnor U29150 (N_29150,N_28346,N_28699);
nand U29151 (N_29151,N_28171,N_28541);
nor U29152 (N_29152,N_28197,N_28521);
xnor U29153 (N_29153,N_28360,N_28861);
nand U29154 (N_29154,N_28629,N_28145);
nor U29155 (N_29155,N_28534,N_28670);
xnor U29156 (N_29156,N_28564,N_28484);
or U29157 (N_29157,N_28813,N_28333);
nand U29158 (N_29158,N_28134,N_28114);
or U29159 (N_29159,N_28304,N_28911);
or U29160 (N_29160,N_28673,N_28793);
or U29161 (N_29161,N_28263,N_28822);
nor U29162 (N_29162,N_28100,N_28099);
and U29163 (N_29163,N_28582,N_28101);
and U29164 (N_29164,N_28238,N_28646);
nor U29165 (N_29165,N_28233,N_28399);
nor U29166 (N_29166,N_28392,N_28415);
nand U29167 (N_29167,N_28136,N_28118);
xnor U29168 (N_29168,N_28972,N_28046);
xnor U29169 (N_29169,N_28547,N_28519);
and U29170 (N_29170,N_28772,N_28738);
nor U29171 (N_29171,N_28721,N_28560);
xnor U29172 (N_29172,N_28141,N_28588);
xor U29173 (N_29173,N_28844,N_28692);
and U29174 (N_29174,N_28231,N_28083);
nor U29175 (N_29175,N_28208,N_28366);
nand U29176 (N_29176,N_28060,N_28039);
or U29177 (N_29177,N_28990,N_28810);
xor U29178 (N_29178,N_28404,N_28506);
xor U29179 (N_29179,N_28421,N_28509);
or U29180 (N_29180,N_28955,N_28744);
or U29181 (N_29181,N_28267,N_28901);
nand U29182 (N_29182,N_28124,N_28454);
nand U29183 (N_29183,N_28496,N_28470);
or U29184 (N_29184,N_28182,N_28913);
or U29185 (N_29185,N_28087,N_28697);
nand U29186 (N_29186,N_28394,N_28009);
xor U29187 (N_29187,N_28864,N_28410);
or U29188 (N_29188,N_28089,N_28873);
or U29189 (N_29189,N_28396,N_28938);
nand U29190 (N_29190,N_28518,N_28155);
nor U29191 (N_29191,N_28860,N_28876);
nand U29192 (N_29192,N_28785,N_28041);
xor U29193 (N_29193,N_28457,N_28368);
or U29194 (N_29194,N_28056,N_28125);
xnor U29195 (N_29195,N_28256,N_28023);
and U29196 (N_29196,N_28994,N_28592);
nor U29197 (N_29197,N_28851,N_28102);
nand U29198 (N_29198,N_28571,N_28049);
or U29199 (N_29199,N_28257,N_28666);
or U29200 (N_29200,N_28222,N_28857);
nand U29201 (N_29201,N_28875,N_28445);
nor U29202 (N_29202,N_28186,N_28818);
and U29203 (N_29203,N_28245,N_28887);
or U29204 (N_29204,N_28299,N_28107);
or U29205 (N_29205,N_28716,N_28158);
nor U29206 (N_29206,N_28650,N_28162);
nand U29207 (N_29207,N_28611,N_28919);
nor U29208 (N_29208,N_28789,N_28269);
or U29209 (N_29209,N_28498,N_28363);
nor U29210 (N_29210,N_28127,N_28189);
xor U29211 (N_29211,N_28685,N_28218);
xnor U29212 (N_29212,N_28067,N_28671);
nand U29213 (N_29213,N_28586,N_28027);
or U29214 (N_29214,N_28042,N_28085);
nand U29215 (N_29215,N_28615,N_28933);
xnor U29216 (N_29216,N_28927,N_28515);
nand U29217 (N_29217,N_28549,N_28565);
and U29218 (N_29218,N_28617,N_28686);
nor U29219 (N_29219,N_28645,N_28578);
or U29220 (N_29220,N_28620,N_28688);
nand U29221 (N_29221,N_28906,N_28308);
or U29222 (N_29222,N_28946,N_28679);
nand U29223 (N_29223,N_28557,N_28265);
nand U29224 (N_29224,N_28014,N_28184);
nor U29225 (N_29225,N_28585,N_28909);
nand U29226 (N_29226,N_28178,N_28803);
nand U29227 (N_29227,N_28596,N_28764);
and U29228 (N_29228,N_28828,N_28079);
or U29229 (N_29229,N_28581,N_28003);
nand U29230 (N_29230,N_28815,N_28669);
and U29231 (N_29231,N_28377,N_28935);
xor U29232 (N_29232,N_28892,N_28886);
and U29233 (N_29233,N_28293,N_28093);
nor U29234 (N_29234,N_28357,N_28225);
and U29235 (N_29235,N_28351,N_28358);
or U29236 (N_29236,N_28109,N_28224);
and U29237 (N_29237,N_28074,N_28482);
or U29238 (N_29238,N_28640,N_28409);
nand U29239 (N_29239,N_28408,N_28271);
nand U29240 (N_29240,N_28371,N_28177);
and U29241 (N_29241,N_28169,N_28264);
xor U29242 (N_29242,N_28066,N_28807);
nor U29243 (N_29243,N_28999,N_28031);
nand U29244 (N_29244,N_28314,N_28190);
and U29245 (N_29245,N_28051,N_28981);
and U29246 (N_29246,N_28932,N_28013);
nor U29247 (N_29247,N_28259,N_28372);
xor U29248 (N_29248,N_28774,N_28804);
or U29249 (N_29249,N_28122,N_28497);
xnor U29250 (N_29250,N_28270,N_28104);
xor U29251 (N_29251,N_28856,N_28071);
nor U29252 (N_29252,N_28841,N_28459);
and U29253 (N_29253,N_28261,N_28709);
nor U29254 (N_29254,N_28511,N_28950);
or U29255 (N_29255,N_28719,N_28969);
xor U29256 (N_29256,N_28055,N_28237);
xnor U29257 (N_29257,N_28425,N_28888);
nand U29258 (N_29258,N_28151,N_28423);
or U29259 (N_29259,N_28285,N_28419);
and U29260 (N_29260,N_28536,N_28452);
nand U29261 (N_29261,N_28370,N_28281);
or U29262 (N_29262,N_28361,N_28365);
nor U29263 (N_29263,N_28733,N_28406);
nand U29264 (N_29264,N_28400,N_28763);
nor U29265 (N_29265,N_28930,N_28654);
and U29266 (N_29266,N_28614,N_28021);
nor U29267 (N_29267,N_28395,N_28910);
xor U29268 (N_29268,N_28978,N_28852);
or U29269 (N_29269,N_28660,N_28010);
xor U29270 (N_29270,N_28130,N_28438);
nor U29271 (N_29271,N_28561,N_28953);
and U29272 (N_29272,N_28754,N_28847);
or U29273 (N_29273,N_28147,N_28247);
nor U29274 (N_29274,N_28554,N_28369);
nor U29275 (N_29275,N_28342,N_28701);
or U29276 (N_29276,N_28019,N_28251);
xor U29277 (N_29277,N_28845,N_28784);
and U29278 (N_29278,N_28632,N_28563);
nor U29279 (N_29279,N_28712,N_28798);
xor U29280 (N_29280,N_28226,N_28492);
nor U29281 (N_29281,N_28002,N_28665);
nand U29282 (N_29282,N_28108,N_28032);
xor U29283 (N_29283,N_28174,N_28428);
or U29284 (N_29284,N_28150,N_28469);
or U29285 (N_29285,N_28393,N_28863);
xnor U29286 (N_29286,N_28417,N_28691);
and U29287 (N_29287,N_28825,N_28276);
nor U29288 (N_29288,N_28133,N_28613);
xor U29289 (N_29289,N_28651,N_28877);
and U29290 (N_29290,N_28327,N_28191);
or U29291 (N_29291,N_28786,N_28062);
or U29292 (N_29292,N_28975,N_28292);
nor U29293 (N_29293,N_28967,N_28606);
xnor U29294 (N_29294,N_28715,N_28962);
and U29295 (N_29295,N_28146,N_28290);
and U29296 (N_29296,N_28659,N_28000);
or U29297 (N_29297,N_28987,N_28501);
nand U29298 (N_29298,N_28905,N_28782);
nor U29299 (N_29299,N_28072,N_28159);
nor U29300 (N_29300,N_28612,N_28300);
nand U29301 (N_29301,N_28773,N_28514);
and U29302 (N_29302,N_28388,N_28672);
and U29303 (N_29303,N_28964,N_28619);
or U29304 (N_29304,N_28517,N_28020);
xnor U29305 (N_29305,N_28064,N_28753);
nor U29306 (N_29306,N_28941,N_28148);
xnor U29307 (N_29307,N_28268,N_28957);
and U29308 (N_29308,N_28120,N_28664);
and U29309 (N_29309,N_28248,N_28796);
and U29310 (N_29310,N_28447,N_28526);
and U29311 (N_29311,N_28332,N_28837);
nand U29312 (N_29312,N_28545,N_28867);
xor U29313 (N_29313,N_28111,N_28986);
xnor U29314 (N_29314,N_28310,N_28139);
and U29315 (N_29315,N_28075,N_28882);
nand U29316 (N_29316,N_28631,N_28577);
nand U29317 (N_29317,N_28170,N_28931);
and U29318 (N_29318,N_28775,N_28006);
nor U29319 (N_29319,N_28081,N_28723);
or U29320 (N_29320,N_28922,N_28702);
and U29321 (N_29321,N_28728,N_28947);
nor U29322 (N_29322,N_28998,N_28811);
nor U29323 (N_29323,N_28326,N_28494);
nand U29324 (N_29324,N_28033,N_28878);
xor U29325 (N_29325,N_28791,N_28834);
nand U29326 (N_29326,N_28819,N_28476);
or U29327 (N_29327,N_28720,N_28260);
or U29328 (N_29328,N_28336,N_28558);
nor U29329 (N_29329,N_28278,N_28157);
nor U29330 (N_29330,N_28928,N_28912);
or U29331 (N_29331,N_28770,N_28921);
xor U29332 (N_29332,N_28414,N_28539);
and U29333 (N_29333,N_28355,N_28865);
nand U29334 (N_29334,N_28250,N_28842);
or U29335 (N_29335,N_28895,N_28641);
nand U29336 (N_29336,N_28971,N_28570);
and U29337 (N_29337,N_28349,N_28486);
nand U29338 (N_29338,N_28504,N_28137);
nor U29339 (N_29339,N_28397,N_28007);
nor U29340 (N_29340,N_28298,N_28736);
nand U29341 (N_29341,N_28809,N_28180);
xor U29342 (N_29342,N_28590,N_28652);
nor U29343 (N_29343,N_28383,N_28647);
nor U29344 (N_29344,N_28724,N_28129);
nand U29345 (N_29345,N_28624,N_28839);
and U29346 (N_29346,N_28605,N_28974);
nand U29347 (N_29347,N_28286,N_28187);
nor U29348 (N_29348,N_28598,N_28531);
and U29349 (N_29349,N_28849,N_28528);
xnor U29350 (N_29350,N_28830,N_28444);
nor U29351 (N_29351,N_28313,N_28138);
nor U29352 (N_29352,N_28591,N_28700);
and U29353 (N_29353,N_28693,N_28420);
nand U29354 (N_29354,N_28350,N_28924);
xnor U29355 (N_29355,N_28574,N_28963);
nand U29356 (N_29356,N_28929,N_28630);
and U29357 (N_29357,N_28376,N_28752);
or U29358 (N_29358,N_28140,N_28325);
xor U29359 (N_29359,N_28088,N_28727);
or U29360 (N_29360,N_28215,N_28289);
xor U29361 (N_29361,N_28198,N_28185);
nor U29362 (N_29362,N_28788,N_28708);
xor U29363 (N_29363,N_28301,N_28078);
xor U29364 (N_29364,N_28742,N_28966);
or U29365 (N_29365,N_28236,N_28338);
xor U29366 (N_29366,N_28826,N_28205);
nor U29367 (N_29367,N_28253,N_28546);
xor U29368 (N_29368,N_28917,N_28029);
and U29369 (N_29369,N_28481,N_28069);
xnor U29370 (N_29370,N_28437,N_28018);
xor U29371 (N_29371,N_28623,N_28183);
nor U29372 (N_29372,N_28034,N_28348);
or U29373 (N_29373,N_28493,N_28048);
and U29374 (N_29374,N_28610,N_28883);
and U29375 (N_29375,N_28603,N_28677);
nand U29376 (N_29376,N_28622,N_28680);
nor U29377 (N_29377,N_28681,N_28683);
or U29378 (N_29378,N_28761,N_28731);
or U29379 (N_29379,N_28689,N_28364);
or U29380 (N_29380,N_28575,N_28829);
and U29381 (N_29381,N_28573,N_28200);
and U29382 (N_29382,N_28080,N_28243);
nor U29383 (N_29383,N_28008,N_28201);
nand U29384 (N_29384,N_28552,N_28037);
xnor U29385 (N_29385,N_28485,N_28747);
nor U29386 (N_29386,N_28235,N_28638);
or U29387 (N_29387,N_28084,N_28126);
nor U29388 (N_29388,N_28472,N_28345);
or U29389 (N_29389,N_28096,N_28335);
nor U29390 (N_29390,N_28777,N_28996);
nor U29391 (N_29391,N_28024,N_28698);
xnor U29392 (N_29392,N_28232,N_28696);
nand U29393 (N_29393,N_28607,N_28781);
nand U29394 (N_29394,N_28077,N_28082);
nand U29395 (N_29395,N_28430,N_28792);
nor U29396 (N_29396,N_28043,N_28142);
nand U29397 (N_29397,N_28025,N_28012);
nor U29398 (N_29398,N_28168,N_28050);
nor U29399 (N_29399,N_28115,N_28322);
or U29400 (N_29400,N_28312,N_28926);
nor U29401 (N_29401,N_28092,N_28983);
nor U29402 (N_29402,N_28918,N_28059);
or U29403 (N_29403,N_28283,N_28783);
or U29404 (N_29404,N_28776,N_28890);
xor U29405 (N_29405,N_28202,N_28853);
nor U29406 (N_29406,N_28835,N_28212);
nor U29407 (N_29407,N_28473,N_28316);
or U29408 (N_29408,N_28272,N_28398);
or U29409 (N_29409,N_28317,N_28467);
and U29410 (N_29410,N_28711,N_28386);
xnor U29411 (N_29411,N_28732,N_28318);
nand U29412 (N_29412,N_28780,N_28156);
nor U29413 (N_29413,N_28328,N_28948);
nand U29414 (N_29414,N_28294,N_28502);
or U29415 (N_29415,N_28431,N_28489);
nor U29416 (N_29416,N_28378,N_28735);
and U29417 (N_29417,N_28945,N_28249);
nand U29418 (N_29418,N_28512,N_28858);
xor U29419 (N_29419,N_28131,N_28817);
xnor U29420 (N_29420,N_28869,N_28756);
nor U29421 (N_29421,N_28319,N_28387);
or U29422 (N_29422,N_28814,N_28166);
or U29423 (N_29423,N_28505,N_28599);
nand U29424 (N_29424,N_28956,N_28758);
nand U29425 (N_29425,N_28374,N_28244);
and U29426 (N_29426,N_28893,N_28524);
xnor U29427 (N_29427,N_28903,N_28495);
nand U29428 (N_29428,N_28977,N_28441);
and U29429 (N_29429,N_28306,N_28188);
nand U29430 (N_29430,N_28566,N_28329);
nand U29431 (N_29431,N_28965,N_28988);
or U29432 (N_29432,N_28436,N_28656);
xnor U29433 (N_29433,N_28302,N_28621);
or U29434 (N_29434,N_28439,N_28730);
nor U29435 (N_29435,N_28533,N_28117);
nand U29436 (N_29436,N_28848,N_28103);
nand U29437 (N_29437,N_28639,N_28760);
nor U29438 (N_29438,N_28874,N_28535);
xnor U29439 (N_29439,N_28196,N_28529);
xnor U29440 (N_29440,N_28152,N_28193);
nand U29441 (N_29441,N_28824,N_28537);
or U29442 (N_29442,N_28491,N_28164);
nand U29443 (N_29443,N_28608,N_28455);
and U29444 (N_29444,N_28655,N_28682);
nand U29445 (N_29445,N_28896,N_28352);
nand U29446 (N_29446,N_28135,N_28181);
xor U29447 (N_29447,N_28480,N_28707);
xor U29448 (N_29448,N_28206,N_28644);
or U29449 (N_29449,N_28734,N_28389);
xor U29450 (N_29450,N_28424,N_28403);
nand U29451 (N_29451,N_28390,N_28755);
and U29452 (N_29452,N_28381,N_28601);
nand U29453 (N_29453,N_28214,N_28451);
xor U29454 (N_29454,N_28771,N_28891);
and U29455 (N_29455,N_28057,N_28110);
nand U29456 (N_29456,N_28154,N_28805);
or U29457 (N_29457,N_28833,N_28207);
nand U29458 (N_29458,N_28713,N_28223);
xor U29459 (N_29459,N_28970,N_28870);
nand U29460 (N_29460,N_28992,N_28407);
or U29461 (N_29461,N_28458,N_28475);
nor U29462 (N_29462,N_28344,N_28739);
xor U29463 (N_29463,N_28343,N_28227);
nor U29464 (N_29464,N_28900,N_28026);
nand U29465 (N_29465,N_28674,N_28556);
or U29466 (N_29466,N_28751,N_28740);
nand U29467 (N_29467,N_28602,N_28741);
xor U29468 (N_29468,N_28255,N_28015);
xnor U29469 (N_29469,N_28195,N_28123);
and U29470 (N_29470,N_28054,N_28503);
nor U29471 (N_29471,N_28675,N_28658);
and U29472 (N_29472,N_28583,N_28525);
xnor U29473 (N_29473,N_28522,N_28516);
nor U29474 (N_29474,N_28562,N_28898);
or U29475 (N_29475,N_28859,N_28038);
or U29476 (N_29476,N_28944,N_28812);
and U29477 (N_29477,N_28416,N_28022);
nand U29478 (N_29478,N_28106,N_28331);
nor U29479 (N_29479,N_28167,N_28466);
or U29480 (N_29480,N_28153,N_28843);
and U29481 (N_29481,N_28375,N_28705);
or U29482 (N_29482,N_28246,N_28885);
and U29483 (N_29483,N_28915,N_28634);
nand U29484 (N_29484,N_28094,N_28984);
nor U29485 (N_29485,N_28061,N_28427);
nand U29486 (N_29486,N_28465,N_28626);
or U29487 (N_29487,N_28176,N_28474);
or U29488 (N_29488,N_28353,N_28625);
xnor U29489 (N_29489,N_28597,N_28113);
and U29490 (N_29490,N_28324,N_28872);
nand U29491 (N_29491,N_28035,N_28936);
xor U29492 (N_29492,N_28745,N_28309);
and U29493 (N_29493,N_28684,N_28800);
xnor U29494 (N_29494,N_28274,N_28315);
and U29495 (N_29495,N_28960,N_28402);
xor U29496 (N_29496,N_28762,N_28916);
xor U29497 (N_29497,N_28609,N_28354);
and U29498 (N_29498,N_28836,N_28052);
and U29499 (N_29499,N_28881,N_28637);
xnor U29500 (N_29500,N_28965,N_28426);
or U29501 (N_29501,N_28382,N_28014);
nor U29502 (N_29502,N_28364,N_28206);
xnor U29503 (N_29503,N_28253,N_28093);
and U29504 (N_29504,N_28721,N_28780);
and U29505 (N_29505,N_28824,N_28685);
nor U29506 (N_29506,N_28322,N_28688);
nand U29507 (N_29507,N_28426,N_28279);
nor U29508 (N_29508,N_28111,N_28843);
and U29509 (N_29509,N_28495,N_28444);
or U29510 (N_29510,N_28075,N_28704);
nor U29511 (N_29511,N_28963,N_28840);
nand U29512 (N_29512,N_28650,N_28681);
or U29513 (N_29513,N_28413,N_28856);
or U29514 (N_29514,N_28974,N_28187);
and U29515 (N_29515,N_28707,N_28440);
xor U29516 (N_29516,N_28034,N_28459);
or U29517 (N_29517,N_28551,N_28366);
and U29518 (N_29518,N_28376,N_28620);
and U29519 (N_29519,N_28929,N_28483);
and U29520 (N_29520,N_28205,N_28495);
xor U29521 (N_29521,N_28467,N_28940);
xnor U29522 (N_29522,N_28734,N_28934);
or U29523 (N_29523,N_28900,N_28472);
or U29524 (N_29524,N_28371,N_28879);
xnor U29525 (N_29525,N_28381,N_28939);
or U29526 (N_29526,N_28771,N_28012);
nor U29527 (N_29527,N_28319,N_28238);
or U29528 (N_29528,N_28850,N_28885);
or U29529 (N_29529,N_28261,N_28363);
nand U29530 (N_29530,N_28251,N_28581);
xnor U29531 (N_29531,N_28177,N_28325);
nand U29532 (N_29532,N_28309,N_28918);
nand U29533 (N_29533,N_28438,N_28887);
nor U29534 (N_29534,N_28915,N_28198);
xor U29535 (N_29535,N_28468,N_28697);
and U29536 (N_29536,N_28776,N_28999);
and U29537 (N_29537,N_28257,N_28774);
or U29538 (N_29538,N_28036,N_28469);
or U29539 (N_29539,N_28005,N_28208);
nand U29540 (N_29540,N_28367,N_28275);
nor U29541 (N_29541,N_28986,N_28521);
xnor U29542 (N_29542,N_28600,N_28755);
nand U29543 (N_29543,N_28851,N_28059);
and U29544 (N_29544,N_28527,N_28993);
nor U29545 (N_29545,N_28579,N_28272);
xnor U29546 (N_29546,N_28073,N_28136);
or U29547 (N_29547,N_28784,N_28021);
xnor U29548 (N_29548,N_28895,N_28640);
nor U29549 (N_29549,N_28660,N_28277);
or U29550 (N_29550,N_28787,N_28853);
xor U29551 (N_29551,N_28040,N_28117);
or U29552 (N_29552,N_28524,N_28746);
and U29553 (N_29553,N_28387,N_28474);
nor U29554 (N_29554,N_28313,N_28110);
and U29555 (N_29555,N_28841,N_28129);
nor U29556 (N_29556,N_28550,N_28725);
and U29557 (N_29557,N_28965,N_28728);
and U29558 (N_29558,N_28281,N_28477);
xnor U29559 (N_29559,N_28123,N_28016);
nand U29560 (N_29560,N_28605,N_28896);
nand U29561 (N_29561,N_28363,N_28942);
nor U29562 (N_29562,N_28589,N_28625);
and U29563 (N_29563,N_28812,N_28405);
nor U29564 (N_29564,N_28346,N_28805);
or U29565 (N_29565,N_28797,N_28702);
or U29566 (N_29566,N_28050,N_28251);
nand U29567 (N_29567,N_28240,N_28321);
nand U29568 (N_29568,N_28359,N_28706);
nor U29569 (N_29569,N_28561,N_28571);
or U29570 (N_29570,N_28201,N_28732);
or U29571 (N_29571,N_28228,N_28728);
nand U29572 (N_29572,N_28784,N_28426);
and U29573 (N_29573,N_28483,N_28747);
nand U29574 (N_29574,N_28370,N_28557);
xor U29575 (N_29575,N_28665,N_28314);
nor U29576 (N_29576,N_28467,N_28933);
nand U29577 (N_29577,N_28625,N_28795);
or U29578 (N_29578,N_28207,N_28345);
xor U29579 (N_29579,N_28945,N_28911);
and U29580 (N_29580,N_28111,N_28580);
and U29581 (N_29581,N_28162,N_28139);
nor U29582 (N_29582,N_28821,N_28828);
or U29583 (N_29583,N_28303,N_28894);
nor U29584 (N_29584,N_28895,N_28792);
xnor U29585 (N_29585,N_28550,N_28074);
and U29586 (N_29586,N_28181,N_28616);
xnor U29587 (N_29587,N_28920,N_28044);
xor U29588 (N_29588,N_28975,N_28339);
nand U29589 (N_29589,N_28291,N_28656);
nand U29590 (N_29590,N_28247,N_28443);
nand U29591 (N_29591,N_28868,N_28469);
nand U29592 (N_29592,N_28467,N_28339);
nand U29593 (N_29593,N_28582,N_28506);
xor U29594 (N_29594,N_28389,N_28857);
nor U29595 (N_29595,N_28221,N_28663);
nor U29596 (N_29596,N_28801,N_28784);
nor U29597 (N_29597,N_28486,N_28635);
nor U29598 (N_29598,N_28753,N_28178);
xnor U29599 (N_29599,N_28721,N_28750);
or U29600 (N_29600,N_28526,N_28323);
nand U29601 (N_29601,N_28726,N_28448);
xor U29602 (N_29602,N_28508,N_28227);
or U29603 (N_29603,N_28720,N_28904);
nor U29604 (N_29604,N_28410,N_28109);
xnor U29605 (N_29605,N_28830,N_28763);
and U29606 (N_29606,N_28025,N_28399);
nand U29607 (N_29607,N_28739,N_28969);
or U29608 (N_29608,N_28571,N_28267);
nand U29609 (N_29609,N_28464,N_28809);
nor U29610 (N_29610,N_28280,N_28541);
nand U29611 (N_29611,N_28211,N_28358);
nor U29612 (N_29612,N_28900,N_28425);
nor U29613 (N_29613,N_28142,N_28913);
nand U29614 (N_29614,N_28063,N_28732);
nor U29615 (N_29615,N_28711,N_28906);
xnor U29616 (N_29616,N_28621,N_28628);
xor U29617 (N_29617,N_28757,N_28855);
nand U29618 (N_29618,N_28485,N_28268);
and U29619 (N_29619,N_28145,N_28742);
xor U29620 (N_29620,N_28048,N_28152);
or U29621 (N_29621,N_28696,N_28870);
or U29622 (N_29622,N_28099,N_28793);
and U29623 (N_29623,N_28924,N_28020);
nor U29624 (N_29624,N_28136,N_28054);
or U29625 (N_29625,N_28693,N_28433);
nand U29626 (N_29626,N_28648,N_28234);
xnor U29627 (N_29627,N_28723,N_28276);
nand U29628 (N_29628,N_28907,N_28151);
nor U29629 (N_29629,N_28631,N_28578);
and U29630 (N_29630,N_28929,N_28957);
xor U29631 (N_29631,N_28010,N_28986);
or U29632 (N_29632,N_28697,N_28195);
nand U29633 (N_29633,N_28321,N_28143);
and U29634 (N_29634,N_28713,N_28281);
or U29635 (N_29635,N_28360,N_28768);
and U29636 (N_29636,N_28014,N_28195);
nand U29637 (N_29637,N_28354,N_28103);
xnor U29638 (N_29638,N_28166,N_28840);
and U29639 (N_29639,N_28795,N_28738);
xnor U29640 (N_29640,N_28415,N_28397);
nor U29641 (N_29641,N_28703,N_28655);
nor U29642 (N_29642,N_28689,N_28116);
xor U29643 (N_29643,N_28911,N_28784);
nand U29644 (N_29644,N_28825,N_28077);
xnor U29645 (N_29645,N_28517,N_28378);
and U29646 (N_29646,N_28827,N_28902);
nand U29647 (N_29647,N_28644,N_28325);
and U29648 (N_29648,N_28796,N_28156);
nand U29649 (N_29649,N_28081,N_28856);
xor U29650 (N_29650,N_28505,N_28598);
nor U29651 (N_29651,N_28777,N_28757);
or U29652 (N_29652,N_28517,N_28550);
nand U29653 (N_29653,N_28552,N_28712);
nand U29654 (N_29654,N_28932,N_28050);
xnor U29655 (N_29655,N_28715,N_28418);
nand U29656 (N_29656,N_28230,N_28803);
xnor U29657 (N_29657,N_28213,N_28259);
or U29658 (N_29658,N_28406,N_28616);
and U29659 (N_29659,N_28425,N_28286);
nand U29660 (N_29660,N_28404,N_28819);
nand U29661 (N_29661,N_28875,N_28954);
xor U29662 (N_29662,N_28671,N_28179);
nand U29663 (N_29663,N_28958,N_28699);
or U29664 (N_29664,N_28423,N_28097);
or U29665 (N_29665,N_28395,N_28136);
xnor U29666 (N_29666,N_28166,N_28546);
or U29667 (N_29667,N_28763,N_28245);
or U29668 (N_29668,N_28485,N_28588);
or U29669 (N_29669,N_28305,N_28826);
nand U29670 (N_29670,N_28148,N_28292);
nand U29671 (N_29671,N_28650,N_28827);
and U29672 (N_29672,N_28508,N_28371);
nor U29673 (N_29673,N_28826,N_28771);
or U29674 (N_29674,N_28567,N_28507);
or U29675 (N_29675,N_28253,N_28594);
nor U29676 (N_29676,N_28927,N_28923);
nor U29677 (N_29677,N_28407,N_28156);
and U29678 (N_29678,N_28652,N_28833);
nor U29679 (N_29679,N_28829,N_28202);
or U29680 (N_29680,N_28064,N_28775);
and U29681 (N_29681,N_28975,N_28867);
nor U29682 (N_29682,N_28122,N_28976);
xor U29683 (N_29683,N_28282,N_28563);
nand U29684 (N_29684,N_28434,N_28358);
or U29685 (N_29685,N_28552,N_28035);
nor U29686 (N_29686,N_28251,N_28213);
or U29687 (N_29687,N_28681,N_28132);
or U29688 (N_29688,N_28832,N_28291);
or U29689 (N_29689,N_28856,N_28340);
or U29690 (N_29690,N_28473,N_28299);
and U29691 (N_29691,N_28520,N_28723);
xnor U29692 (N_29692,N_28842,N_28653);
and U29693 (N_29693,N_28610,N_28511);
and U29694 (N_29694,N_28366,N_28141);
or U29695 (N_29695,N_28788,N_28564);
and U29696 (N_29696,N_28603,N_28479);
and U29697 (N_29697,N_28064,N_28417);
nor U29698 (N_29698,N_28083,N_28054);
or U29699 (N_29699,N_28285,N_28516);
nand U29700 (N_29700,N_28785,N_28636);
nor U29701 (N_29701,N_28329,N_28843);
nand U29702 (N_29702,N_28237,N_28771);
or U29703 (N_29703,N_28207,N_28904);
xnor U29704 (N_29704,N_28481,N_28984);
and U29705 (N_29705,N_28098,N_28854);
nor U29706 (N_29706,N_28177,N_28091);
xnor U29707 (N_29707,N_28605,N_28410);
and U29708 (N_29708,N_28989,N_28325);
nor U29709 (N_29709,N_28729,N_28736);
and U29710 (N_29710,N_28174,N_28909);
and U29711 (N_29711,N_28558,N_28535);
or U29712 (N_29712,N_28381,N_28848);
nor U29713 (N_29713,N_28975,N_28393);
and U29714 (N_29714,N_28462,N_28951);
nand U29715 (N_29715,N_28803,N_28214);
nand U29716 (N_29716,N_28056,N_28018);
or U29717 (N_29717,N_28425,N_28402);
xor U29718 (N_29718,N_28445,N_28968);
or U29719 (N_29719,N_28473,N_28031);
or U29720 (N_29720,N_28387,N_28156);
nor U29721 (N_29721,N_28486,N_28603);
xnor U29722 (N_29722,N_28453,N_28759);
or U29723 (N_29723,N_28755,N_28665);
nand U29724 (N_29724,N_28862,N_28550);
or U29725 (N_29725,N_28968,N_28066);
or U29726 (N_29726,N_28947,N_28471);
xnor U29727 (N_29727,N_28684,N_28504);
nand U29728 (N_29728,N_28355,N_28007);
nor U29729 (N_29729,N_28483,N_28859);
nor U29730 (N_29730,N_28295,N_28328);
nor U29731 (N_29731,N_28020,N_28577);
and U29732 (N_29732,N_28514,N_28499);
nor U29733 (N_29733,N_28814,N_28664);
xnor U29734 (N_29734,N_28191,N_28257);
and U29735 (N_29735,N_28540,N_28582);
or U29736 (N_29736,N_28618,N_28141);
nand U29737 (N_29737,N_28970,N_28930);
and U29738 (N_29738,N_28508,N_28615);
nor U29739 (N_29739,N_28067,N_28294);
or U29740 (N_29740,N_28534,N_28716);
nor U29741 (N_29741,N_28225,N_28766);
xor U29742 (N_29742,N_28304,N_28401);
nor U29743 (N_29743,N_28998,N_28828);
nor U29744 (N_29744,N_28633,N_28794);
nor U29745 (N_29745,N_28262,N_28771);
nand U29746 (N_29746,N_28414,N_28329);
xor U29747 (N_29747,N_28613,N_28586);
nand U29748 (N_29748,N_28246,N_28006);
xnor U29749 (N_29749,N_28061,N_28539);
or U29750 (N_29750,N_28055,N_28897);
nor U29751 (N_29751,N_28545,N_28052);
nand U29752 (N_29752,N_28493,N_28893);
and U29753 (N_29753,N_28485,N_28897);
xnor U29754 (N_29754,N_28994,N_28618);
nor U29755 (N_29755,N_28246,N_28891);
and U29756 (N_29756,N_28760,N_28958);
xnor U29757 (N_29757,N_28920,N_28977);
or U29758 (N_29758,N_28480,N_28699);
xnor U29759 (N_29759,N_28014,N_28035);
and U29760 (N_29760,N_28335,N_28958);
and U29761 (N_29761,N_28696,N_28183);
nand U29762 (N_29762,N_28929,N_28490);
nand U29763 (N_29763,N_28304,N_28543);
nand U29764 (N_29764,N_28397,N_28882);
or U29765 (N_29765,N_28940,N_28956);
nor U29766 (N_29766,N_28025,N_28895);
xor U29767 (N_29767,N_28100,N_28130);
nand U29768 (N_29768,N_28498,N_28847);
xor U29769 (N_29769,N_28250,N_28792);
and U29770 (N_29770,N_28967,N_28138);
or U29771 (N_29771,N_28710,N_28709);
xnor U29772 (N_29772,N_28631,N_28135);
or U29773 (N_29773,N_28236,N_28911);
nand U29774 (N_29774,N_28734,N_28629);
or U29775 (N_29775,N_28173,N_28706);
or U29776 (N_29776,N_28405,N_28488);
nor U29777 (N_29777,N_28394,N_28007);
xor U29778 (N_29778,N_28153,N_28862);
nand U29779 (N_29779,N_28607,N_28390);
nand U29780 (N_29780,N_28492,N_28776);
xor U29781 (N_29781,N_28127,N_28622);
nor U29782 (N_29782,N_28107,N_28276);
and U29783 (N_29783,N_28679,N_28661);
nand U29784 (N_29784,N_28246,N_28795);
and U29785 (N_29785,N_28854,N_28662);
or U29786 (N_29786,N_28386,N_28190);
nand U29787 (N_29787,N_28345,N_28595);
and U29788 (N_29788,N_28232,N_28638);
nand U29789 (N_29789,N_28380,N_28546);
and U29790 (N_29790,N_28973,N_28082);
or U29791 (N_29791,N_28305,N_28792);
or U29792 (N_29792,N_28816,N_28402);
xor U29793 (N_29793,N_28054,N_28398);
nand U29794 (N_29794,N_28852,N_28669);
nor U29795 (N_29795,N_28955,N_28337);
xor U29796 (N_29796,N_28733,N_28718);
or U29797 (N_29797,N_28388,N_28569);
nand U29798 (N_29798,N_28448,N_28552);
or U29799 (N_29799,N_28417,N_28776);
nand U29800 (N_29800,N_28270,N_28730);
nor U29801 (N_29801,N_28431,N_28217);
nor U29802 (N_29802,N_28673,N_28761);
nor U29803 (N_29803,N_28779,N_28724);
and U29804 (N_29804,N_28648,N_28528);
and U29805 (N_29805,N_28695,N_28361);
nor U29806 (N_29806,N_28961,N_28928);
or U29807 (N_29807,N_28622,N_28299);
nor U29808 (N_29808,N_28018,N_28540);
or U29809 (N_29809,N_28061,N_28675);
xor U29810 (N_29810,N_28827,N_28429);
nand U29811 (N_29811,N_28389,N_28228);
or U29812 (N_29812,N_28852,N_28796);
or U29813 (N_29813,N_28794,N_28319);
nor U29814 (N_29814,N_28871,N_28197);
xnor U29815 (N_29815,N_28370,N_28454);
xnor U29816 (N_29816,N_28874,N_28246);
nor U29817 (N_29817,N_28051,N_28289);
xor U29818 (N_29818,N_28456,N_28000);
and U29819 (N_29819,N_28238,N_28372);
and U29820 (N_29820,N_28732,N_28648);
nor U29821 (N_29821,N_28590,N_28654);
nor U29822 (N_29822,N_28426,N_28718);
and U29823 (N_29823,N_28922,N_28877);
nand U29824 (N_29824,N_28317,N_28529);
nor U29825 (N_29825,N_28862,N_28728);
or U29826 (N_29826,N_28958,N_28315);
xnor U29827 (N_29827,N_28030,N_28886);
nor U29828 (N_29828,N_28512,N_28156);
xor U29829 (N_29829,N_28968,N_28294);
nand U29830 (N_29830,N_28195,N_28269);
and U29831 (N_29831,N_28203,N_28675);
xnor U29832 (N_29832,N_28490,N_28212);
and U29833 (N_29833,N_28244,N_28071);
xnor U29834 (N_29834,N_28765,N_28412);
xor U29835 (N_29835,N_28238,N_28800);
xor U29836 (N_29836,N_28431,N_28854);
or U29837 (N_29837,N_28008,N_28182);
xor U29838 (N_29838,N_28342,N_28722);
and U29839 (N_29839,N_28715,N_28402);
or U29840 (N_29840,N_28960,N_28720);
xor U29841 (N_29841,N_28815,N_28780);
or U29842 (N_29842,N_28274,N_28752);
and U29843 (N_29843,N_28717,N_28595);
xnor U29844 (N_29844,N_28040,N_28336);
or U29845 (N_29845,N_28643,N_28087);
and U29846 (N_29846,N_28547,N_28598);
nor U29847 (N_29847,N_28379,N_28705);
nand U29848 (N_29848,N_28800,N_28886);
xnor U29849 (N_29849,N_28516,N_28512);
nor U29850 (N_29850,N_28940,N_28840);
nand U29851 (N_29851,N_28016,N_28534);
xor U29852 (N_29852,N_28975,N_28690);
nand U29853 (N_29853,N_28826,N_28679);
and U29854 (N_29854,N_28786,N_28194);
and U29855 (N_29855,N_28104,N_28230);
or U29856 (N_29856,N_28500,N_28036);
nand U29857 (N_29857,N_28439,N_28661);
xnor U29858 (N_29858,N_28739,N_28643);
nand U29859 (N_29859,N_28271,N_28249);
nand U29860 (N_29860,N_28305,N_28626);
or U29861 (N_29861,N_28238,N_28579);
or U29862 (N_29862,N_28718,N_28627);
or U29863 (N_29863,N_28977,N_28226);
nor U29864 (N_29864,N_28581,N_28809);
and U29865 (N_29865,N_28157,N_28603);
and U29866 (N_29866,N_28502,N_28393);
nor U29867 (N_29867,N_28787,N_28322);
nand U29868 (N_29868,N_28448,N_28089);
nand U29869 (N_29869,N_28805,N_28468);
or U29870 (N_29870,N_28052,N_28811);
or U29871 (N_29871,N_28460,N_28382);
or U29872 (N_29872,N_28970,N_28830);
and U29873 (N_29873,N_28651,N_28737);
or U29874 (N_29874,N_28313,N_28795);
or U29875 (N_29875,N_28947,N_28382);
and U29876 (N_29876,N_28142,N_28219);
and U29877 (N_29877,N_28421,N_28781);
xnor U29878 (N_29878,N_28976,N_28341);
and U29879 (N_29879,N_28649,N_28575);
nor U29880 (N_29880,N_28968,N_28299);
nor U29881 (N_29881,N_28347,N_28156);
and U29882 (N_29882,N_28313,N_28783);
xnor U29883 (N_29883,N_28295,N_28983);
or U29884 (N_29884,N_28261,N_28008);
nor U29885 (N_29885,N_28223,N_28818);
nor U29886 (N_29886,N_28915,N_28695);
and U29887 (N_29887,N_28302,N_28427);
nand U29888 (N_29888,N_28842,N_28536);
nor U29889 (N_29889,N_28964,N_28641);
nor U29890 (N_29890,N_28758,N_28876);
xnor U29891 (N_29891,N_28391,N_28519);
and U29892 (N_29892,N_28799,N_28578);
nand U29893 (N_29893,N_28502,N_28975);
xor U29894 (N_29894,N_28290,N_28324);
xor U29895 (N_29895,N_28323,N_28998);
nor U29896 (N_29896,N_28305,N_28170);
nor U29897 (N_29897,N_28113,N_28236);
xor U29898 (N_29898,N_28833,N_28005);
nor U29899 (N_29899,N_28039,N_28212);
xor U29900 (N_29900,N_28029,N_28712);
and U29901 (N_29901,N_28678,N_28416);
and U29902 (N_29902,N_28276,N_28722);
nor U29903 (N_29903,N_28055,N_28743);
xnor U29904 (N_29904,N_28633,N_28735);
nand U29905 (N_29905,N_28641,N_28341);
or U29906 (N_29906,N_28082,N_28920);
nor U29907 (N_29907,N_28782,N_28804);
nor U29908 (N_29908,N_28287,N_28729);
and U29909 (N_29909,N_28708,N_28111);
and U29910 (N_29910,N_28956,N_28182);
nor U29911 (N_29911,N_28815,N_28750);
xor U29912 (N_29912,N_28428,N_28763);
nand U29913 (N_29913,N_28465,N_28691);
and U29914 (N_29914,N_28628,N_28565);
or U29915 (N_29915,N_28841,N_28204);
or U29916 (N_29916,N_28182,N_28691);
nand U29917 (N_29917,N_28810,N_28076);
nor U29918 (N_29918,N_28137,N_28718);
or U29919 (N_29919,N_28378,N_28334);
and U29920 (N_29920,N_28210,N_28242);
nor U29921 (N_29921,N_28637,N_28331);
nand U29922 (N_29922,N_28274,N_28746);
nor U29923 (N_29923,N_28044,N_28034);
nor U29924 (N_29924,N_28407,N_28744);
xnor U29925 (N_29925,N_28328,N_28393);
and U29926 (N_29926,N_28986,N_28476);
xnor U29927 (N_29927,N_28900,N_28786);
xor U29928 (N_29928,N_28569,N_28381);
nor U29929 (N_29929,N_28227,N_28982);
xnor U29930 (N_29930,N_28563,N_28885);
nand U29931 (N_29931,N_28740,N_28530);
nor U29932 (N_29932,N_28664,N_28091);
nand U29933 (N_29933,N_28954,N_28961);
nor U29934 (N_29934,N_28807,N_28761);
and U29935 (N_29935,N_28819,N_28240);
xor U29936 (N_29936,N_28314,N_28680);
and U29937 (N_29937,N_28105,N_28270);
nor U29938 (N_29938,N_28650,N_28904);
or U29939 (N_29939,N_28671,N_28580);
or U29940 (N_29940,N_28660,N_28849);
xnor U29941 (N_29941,N_28352,N_28053);
nand U29942 (N_29942,N_28124,N_28849);
xor U29943 (N_29943,N_28084,N_28927);
nor U29944 (N_29944,N_28594,N_28125);
nor U29945 (N_29945,N_28323,N_28097);
xor U29946 (N_29946,N_28269,N_28714);
and U29947 (N_29947,N_28549,N_28632);
or U29948 (N_29948,N_28304,N_28034);
and U29949 (N_29949,N_28167,N_28135);
nor U29950 (N_29950,N_28000,N_28979);
xor U29951 (N_29951,N_28619,N_28614);
or U29952 (N_29952,N_28531,N_28408);
or U29953 (N_29953,N_28637,N_28308);
nor U29954 (N_29954,N_28683,N_28062);
and U29955 (N_29955,N_28404,N_28244);
nor U29956 (N_29956,N_28719,N_28460);
nor U29957 (N_29957,N_28708,N_28676);
nand U29958 (N_29958,N_28791,N_28992);
xor U29959 (N_29959,N_28147,N_28176);
or U29960 (N_29960,N_28851,N_28489);
and U29961 (N_29961,N_28562,N_28058);
nor U29962 (N_29962,N_28979,N_28663);
xor U29963 (N_29963,N_28202,N_28779);
nand U29964 (N_29964,N_28948,N_28157);
nand U29965 (N_29965,N_28500,N_28955);
xnor U29966 (N_29966,N_28363,N_28989);
xnor U29967 (N_29967,N_28486,N_28453);
or U29968 (N_29968,N_28459,N_28003);
nand U29969 (N_29969,N_28829,N_28644);
xor U29970 (N_29970,N_28171,N_28087);
nand U29971 (N_29971,N_28553,N_28525);
nor U29972 (N_29972,N_28563,N_28387);
nor U29973 (N_29973,N_28105,N_28233);
xnor U29974 (N_29974,N_28363,N_28655);
or U29975 (N_29975,N_28151,N_28618);
or U29976 (N_29976,N_28727,N_28604);
or U29977 (N_29977,N_28024,N_28945);
nand U29978 (N_29978,N_28490,N_28576);
nand U29979 (N_29979,N_28227,N_28746);
nor U29980 (N_29980,N_28524,N_28634);
and U29981 (N_29981,N_28569,N_28591);
nor U29982 (N_29982,N_28976,N_28532);
xnor U29983 (N_29983,N_28961,N_28316);
nor U29984 (N_29984,N_28483,N_28955);
nor U29985 (N_29985,N_28662,N_28557);
and U29986 (N_29986,N_28010,N_28785);
nand U29987 (N_29987,N_28549,N_28103);
nor U29988 (N_29988,N_28094,N_28859);
nand U29989 (N_29989,N_28561,N_28890);
xnor U29990 (N_29990,N_28913,N_28934);
or U29991 (N_29991,N_28198,N_28786);
and U29992 (N_29992,N_28454,N_28365);
xnor U29993 (N_29993,N_28819,N_28499);
nand U29994 (N_29994,N_28603,N_28537);
and U29995 (N_29995,N_28847,N_28681);
xor U29996 (N_29996,N_28741,N_28556);
and U29997 (N_29997,N_28935,N_28769);
xnor U29998 (N_29998,N_28571,N_28569);
or U29999 (N_29999,N_28344,N_28427);
xor UO_0 (O_0,N_29514,N_29087);
nand UO_1 (O_1,N_29509,N_29807);
nor UO_2 (O_2,N_29838,N_29898);
nor UO_3 (O_3,N_29887,N_29129);
nand UO_4 (O_4,N_29960,N_29348);
or UO_5 (O_5,N_29506,N_29248);
nand UO_6 (O_6,N_29830,N_29632);
nor UO_7 (O_7,N_29667,N_29569);
nor UO_8 (O_8,N_29567,N_29237);
nand UO_9 (O_9,N_29730,N_29521);
or UO_10 (O_10,N_29800,N_29902);
nand UO_11 (O_11,N_29221,N_29616);
nand UO_12 (O_12,N_29552,N_29818);
nand UO_13 (O_13,N_29401,N_29640);
nand UO_14 (O_14,N_29613,N_29454);
and UO_15 (O_15,N_29903,N_29549);
or UO_16 (O_16,N_29125,N_29490);
nor UO_17 (O_17,N_29264,N_29469);
and UO_18 (O_18,N_29048,N_29097);
or UO_19 (O_19,N_29849,N_29657);
xnor UO_20 (O_20,N_29741,N_29932);
and UO_21 (O_21,N_29132,N_29115);
or UO_22 (O_22,N_29277,N_29750);
or UO_23 (O_23,N_29540,N_29359);
nor UO_24 (O_24,N_29376,N_29899);
and UO_25 (O_25,N_29319,N_29833);
xor UO_26 (O_26,N_29166,N_29980);
nor UO_27 (O_27,N_29752,N_29385);
or UO_28 (O_28,N_29735,N_29679);
and UO_29 (O_29,N_29421,N_29607);
xor UO_30 (O_30,N_29384,N_29590);
or UO_31 (O_31,N_29988,N_29497);
and UO_32 (O_32,N_29227,N_29229);
and UO_33 (O_33,N_29949,N_29621);
or UO_34 (O_34,N_29892,N_29714);
and UO_35 (O_35,N_29769,N_29772);
xor UO_36 (O_36,N_29163,N_29969);
nand UO_37 (O_37,N_29910,N_29940);
or UO_38 (O_38,N_29602,N_29516);
or UO_39 (O_39,N_29245,N_29456);
and UO_40 (O_40,N_29099,N_29395);
xor UO_41 (O_41,N_29620,N_29782);
xnor UO_42 (O_42,N_29909,N_29143);
xnor UO_43 (O_43,N_29146,N_29022);
or UO_44 (O_44,N_29071,N_29976);
nor UO_45 (O_45,N_29078,N_29826);
xnor UO_46 (O_46,N_29234,N_29530);
and UO_47 (O_47,N_29130,N_29236);
nand UO_48 (O_48,N_29536,N_29811);
nand UO_49 (O_49,N_29825,N_29339);
nor UO_50 (O_50,N_29795,N_29770);
xor UO_51 (O_51,N_29928,N_29799);
xor UO_52 (O_52,N_29453,N_29803);
nor UO_53 (O_53,N_29559,N_29832);
or UO_54 (O_54,N_29983,N_29990);
nand UO_55 (O_55,N_29513,N_29879);
nor UO_56 (O_56,N_29089,N_29161);
or UO_57 (O_57,N_29318,N_29011);
nand UO_58 (O_58,N_29193,N_29827);
and UO_59 (O_59,N_29324,N_29634);
or UO_60 (O_60,N_29953,N_29205);
xnor UO_61 (O_61,N_29499,N_29906);
and UO_62 (O_62,N_29583,N_29578);
nor UO_63 (O_63,N_29045,N_29950);
xnor UO_64 (O_64,N_29758,N_29177);
xor UO_65 (O_65,N_29995,N_29265);
or UO_66 (O_66,N_29195,N_29939);
xnor UO_67 (O_67,N_29186,N_29968);
nor UO_68 (O_68,N_29785,N_29472);
or UO_69 (O_69,N_29531,N_29542);
nand UO_70 (O_70,N_29481,N_29656);
and UO_71 (O_71,N_29780,N_29343);
nor UO_72 (O_72,N_29076,N_29913);
and UO_73 (O_73,N_29996,N_29432);
and UO_74 (O_74,N_29669,N_29708);
or UO_75 (O_75,N_29707,N_29209);
nor UO_76 (O_76,N_29912,N_29415);
nand UO_77 (O_77,N_29659,N_29035);
and UO_78 (O_78,N_29031,N_29337);
xor UO_79 (O_79,N_29926,N_29523);
or UO_80 (O_80,N_29214,N_29680);
and UO_81 (O_81,N_29283,N_29999);
nand UO_82 (O_82,N_29139,N_29352);
xor UO_83 (O_83,N_29170,N_29500);
xnor UO_84 (O_84,N_29331,N_29231);
nor UO_85 (O_85,N_29055,N_29353);
or UO_86 (O_86,N_29340,N_29576);
xor UO_87 (O_87,N_29965,N_29548);
or UO_88 (O_88,N_29649,N_29654);
or UO_89 (O_89,N_29298,N_29972);
or UO_90 (O_90,N_29003,N_29515);
nor UO_91 (O_91,N_29777,N_29639);
xnor UO_92 (O_92,N_29183,N_29273);
nor UO_93 (O_93,N_29922,N_29042);
and UO_94 (O_94,N_29646,N_29451);
xnor UO_95 (O_95,N_29225,N_29062);
nor UO_96 (O_96,N_29437,N_29554);
nor UO_97 (O_97,N_29598,N_29282);
and UO_98 (O_98,N_29582,N_29916);
xnor UO_99 (O_99,N_29556,N_29094);
or UO_100 (O_100,N_29762,N_29550);
xnor UO_101 (O_101,N_29893,N_29368);
or UO_102 (O_102,N_29495,N_29105);
xor UO_103 (O_103,N_29661,N_29109);
nor UO_104 (O_104,N_29015,N_29030);
nor UO_105 (O_105,N_29502,N_29178);
xor UO_106 (O_106,N_29993,N_29631);
nor UO_107 (O_107,N_29058,N_29781);
nor UO_108 (O_108,N_29285,N_29301);
or UO_109 (O_109,N_29111,N_29459);
or UO_110 (O_110,N_29036,N_29216);
or UO_111 (O_111,N_29617,N_29788);
nand UO_112 (O_112,N_29180,N_29921);
or UO_113 (O_113,N_29256,N_29544);
nand UO_114 (O_114,N_29737,N_29215);
xor UO_115 (O_115,N_29624,N_29837);
nor UO_116 (O_116,N_29822,N_29228);
nor UO_117 (O_117,N_29140,N_29270);
or UO_118 (O_118,N_29528,N_29239);
nand UO_119 (O_119,N_29619,N_29450);
or UO_120 (O_120,N_29158,N_29241);
and UO_121 (O_121,N_29464,N_29846);
or UO_122 (O_122,N_29424,N_29056);
nand UO_123 (O_123,N_29573,N_29683);
and UO_124 (O_124,N_29745,N_29038);
xnor UO_125 (O_125,N_29079,N_29476);
or UO_126 (O_126,N_29757,N_29753);
xnor UO_127 (O_127,N_29244,N_29606);
and UO_128 (O_128,N_29179,N_29853);
nor UO_129 (O_129,N_29806,N_29703);
nand UO_130 (O_130,N_29915,N_29650);
nor UO_131 (O_131,N_29726,N_29756);
xor UO_132 (O_132,N_29603,N_29059);
or UO_133 (O_133,N_29314,N_29964);
and UO_134 (O_134,N_29175,N_29819);
and UO_135 (O_135,N_29197,N_29802);
nand UO_136 (O_136,N_29086,N_29439);
nand UO_137 (O_137,N_29941,N_29392);
xor UO_138 (O_138,N_29814,N_29411);
xor UO_139 (O_139,N_29103,N_29057);
nor UO_140 (O_140,N_29355,N_29841);
nand UO_141 (O_141,N_29615,N_29463);
and UO_142 (O_142,N_29890,N_29959);
nor UO_143 (O_143,N_29191,N_29749);
or UO_144 (O_144,N_29519,N_29108);
and UO_145 (O_145,N_29370,N_29151);
xor UO_146 (O_146,N_29759,N_29026);
xor UO_147 (O_147,N_29341,N_29627);
xnor UO_148 (O_148,N_29865,N_29309);
xor UO_149 (O_149,N_29718,N_29091);
xor UO_150 (O_150,N_29958,N_29378);
and UO_151 (O_151,N_29250,N_29660);
nand UO_152 (O_152,N_29075,N_29564);
or UO_153 (O_153,N_29110,N_29520);
xnor UO_154 (O_154,N_29375,N_29966);
and UO_155 (O_155,N_29860,N_29948);
nand UO_156 (O_156,N_29678,N_29013);
nor UO_157 (O_157,N_29389,N_29755);
nor UO_158 (O_158,N_29297,N_29347);
or UO_159 (O_159,N_29713,N_29494);
and UO_160 (O_160,N_29073,N_29754);
or UO_161 (O_161,N_29246,N_29586);
xnor UO_162 (O_162,N_29824,N_29532);
nor UO_163 (O_163,N_29066,N_29695);
and UO_164 (O_164,N_29417,N_29278);
xor UO_165 (O_165,N_29374,N_29033);
or UO_166 (O_166,N_29380,N_29767);
nor UO_167 (O_167,N_29206,N_29700);
xnor UO_168 (O_168,N_29449,N_29570);
and UO_169 (O_169,N_29200,N_29484);
and UO_170 (O_170,N_29687,N_29396);
and UO_171 (O_171,N_29652,N_29252);
or UO_172 (O_172,N_29302,N_29159);
nor UO_173 (O_173,N_29386,N_29409);
nand UO_174 (O_174,N_29367,N_29369);
nand UO_175 (O_175,N_29203,N_29346);
nand UO_176 (O_176,N_29560,N_29051);
nand UO_177 (O_177,N_29247,N_29333);
nand UO_178 (O_178,N_29118,N_29230);
and UO_179 (O_179,N_29381,N_29072);
nand UO_180 (O_180,N_29723,N_29611);
nor UO_181 (O_181,N_29082,N_29039);
nand UO_182 (O_182,N_29303,N_29740);
xnor UO_183 (O_183,N_29967,N_29731);
and UO_184 (O_184,N_29190,N_29300);
nand UO_185 (O_185,N_29345,N_29223);
nand UO_186 (O_186,N_29208,N_29350);
or UO_187 (O_187,N_29947,N_29291);
nor UO_188 (O_188,N_29771,N_29383);
nor UO_189 (O_189,N_29642,N_29336);
and UO_190 (O_190,N_29496,N_29946);
xor UO_191 (O_191,N_29222,N_29101);
xnor UO_192 (O_192,N_29522,N_29594);
nand UO_193 (O_193,N_29169,N_29761);
or UO_194 (O_194,N_29982,N_29287);
nor UO_195 (O_195,N_29410,N_29002);
nand UO_196 (O_196,N_29435,N_29334);
and UO_197 (O_197,N_29828,N_29263);
nor UO_198 (O_198,N_29775,N_29877);
or UO_199 (O_199,N_29136,N_29307);
and UO_200 (O_200,N_29942,N_29486);
xor UO_201 (O_201,N_29455,N_29153);
and UO_202 (O_202,N_29474,N_29004);
xor UO_203 (O_203,N_29801,N_29870);
nand UO_204 (O_204,N_29604,N_29275);
xor UO_205 (O_205,N_29137,N_29407);
and UO_206 (O_206,N_29693,N_29400);
and UO_207 (O_207,N_29212,N_29167);
nand UO_208 (O_208,N_29905,N_29581);
nand UO_209 (O_209,N_29289,N_29473);
nor UO_210 (O_210,N_29671,N_29371);
nand UO_211 (O_211,N_29356,N_29290);
and UO_212 (O_212,N_29238,N_29043);
and UO_213 (O_213,N_29557,N_29629);
or UO_214 (O_214,N_29046,N_29120);
xor UO_215 (O_215,N_29638,N_29738);
xor UO_216 (O_216,N_29975,N_29468);
xor UO_217 (O_217,N_29416,N_29147);
and UO_218 (O_218,N_29269,N_29413);
xnor UO_219 (O_219,N_29460,N_29436);
nand UO_220 (O_220,N_29483,N_29839);
xor UO_221 (O_221,N_29872,N_29406);
xnor UO_222 (O_222,N_29106,N_29719);
and UO_223 (O_223,N_29251,N_29171);
xnor UO_224 (O_224,N_29390,N_29475);
xnor UO_225 (O_225,N_29000,N_29527);
and UO_226 (O_226,N_29834,N_29794);
nor UO_227 (O_227,N_29694,N_29024);
nor UO_228 (O_228,N_29956,N_29253);
nor UO_229 (O_229,N_29541,N_29973);
nor UO_230 (O_230,N_29875,N_29373);
and UO_231 (O_231,N_29842,N_29596);
nor UO_232 (O_232,N_29701,N_29864);
and UO_233 (O_233,N_29697,N_29847);
and UO_234 (O_234,N_29600,N_29776);
nand UO_235 (O_235,N_29280,N_29243);
xnor UO_236 (O_236,N_29081,N_29744);
nand UO_237 (O_237,N_29260,N_29836);
nor UO_238 (O_238,N_29722,N_29595);
nor UO_239 (O_239,N_29618,N_29927);
nor UO_240 (O_240,N_29562,N_29812);
xnor UO_241 (O_241,N_29665,N_29907);
nor UO_242 (O_242,N_29991,N_29187);
or UO_243 (O_243,N_29485,N_29420);
nor UO_244 (O_244,N_29461,N_29001);
xor UO_245 (O_245,N_29335,N_29168);
nand UO_246 (O_246,N_29891,N_29878);
nand UO_247 (O_247,N_29090,N_29625);
and UO_248 (O_248,N_29537,N_29050);
or UO_249 (O_249,N_29184,N_29571);
nor UO_250 (O_250,N_29820,N_29119);
nor UO_251 (O_251,N_29141,N_29746);
nor UO_252 (O_252,N_29085,N_29018);
and UO_253 (O_253,N_29696,N_29635);
nor UO_254 (O_254,N_29428,N_29725);
nand UO_255 (O_255,N_29561,N_29778);
xnor UO_256 (O_256,N_29023,N_29342);
or UO_257 (O_257,N_29447,N_29831);
or UO_258 (O_258,N_29816,N_29008);
nand UO_259 (O_259,N_29391,N_29142);
and UO_260 (O_260,N_29525,N_29242);
xnor UO_261 (O_261,N_29405,N_29255);
nand UO_262 (O_262,N_29543,N_29354);
and UO_263 (O_263,N_29492,N_29313);
xnor UO_264 (O_264,N_29727,N_29845);
nor UO_265 (O_265,N_29507,N_29937);
or UO_266 (O_266,N_29226,N_29176);
xnor UO_267 (O_267,N_29053,N_29107);
xnor UO_268 (O_268,N_29419,N_29123);
nand UO_269 (O_269,N_29423,N_29064);
xnor UO_270 (O_270,N_29539,N_29458);
nor UO_271 (O_271,N_29095,N_29029);
or UO_272 (O_272,N_29593,N_29686);
or UO_273 (O_273,N_29098,N_29565);
and UO_274 (O_274,N_29936,N_29148);
nand UO_275 (O_275,N_29360,N_29729);
or UO_276 (O_276,N_29466,N_29007);
nor UO_277 (O_277,N_29052,N_29633);
or UO_278 (O_278,N_29597,N_29970);
xor UO_279 (O_279,N_29526,N_29124);
and UO_280 (O_280,N_29572,N_29470);
nor UO_281 (O_281,N_29145,N_29551);
nand UO_282 (O_282,N_29293,N_29317);
and UO_283 (O_283,N_29808,N_29897);
and UO_284 (O_284,N_29748,N_29358);
or UO_285 (O_285,N_29404,N_29612);
and UO_286 (O_286,N_29135,N_29773);
nor UO_287 (O_287,N_29249,N_29900);
nor UO_288 (O_288,N_29357,N_29880);
and UO_289 (O_289,N_29784,N_29764);
and UO_290 (O_290,N_29403,N_29152);
xnor UO_291 (O_291,N_29288,N_29935);
nor UO_292 (O_292,N_29173,N_29259);
or UO_293 (O_293,N_29911,N_29217);
nor UO_294 (O_294,N_29019,N_29889);
nand UO_295 (O_295,N_29194,N_29568);
or UO_296 (O_296,N_29821,N_29804);
xor UO_297 (O_297,N_29920,N_29306);
and UO_298 (O_298,N_29235,N_29041);
nor UO_299 (O_299,N_29080,N_29524);
or UO_300 (O_300,N_29162,N_29813);
and UO_301 (O_301,N_29016,N_29295);
or UO_302 (O_302,N_29862,N_29742);
nand UO_303 (O_303,N_29734,N_29711);
and UO_304 (O_304,N_29704,N_29427);
and UO_305 (O_305,N_29326,N_29365);
nor UO_306 (O_306,N_29866,N_29692);
or UO_307 (O_307,N_29533,N_29330);
and UO_308 (O_308,N_29589,N_29442);
nand UO_309 (O_309,N_29279,N_29088);
nand UO_310 (O_310,N_29211,N_29857);
xnor UO_311 (O_311,N_29257,N_29321);
or UO_312 (O_312,N_29299,N_29553);
or UO_313 (O_313,N_29637,N_29272);
and UO_314 (O_314,N_29308,N_29848);
and UO_315 (O_315,N_29823,N_29732);
and UO_316 (O_316,N_29883,N_29805);
nor UO_317 (O_317,N_29724,N_29363);
nand UO_318 (O_318,N_29651,N_29418);
nor UO_319 (O_319,N_29009,N_29760);
nor UO_320 (O_320,N_29574,N_29869);
nand UO_321 (O_321,N_29325,N_29316);
xor UO_322 (O_322,N_29233,N_29037);
xor UO_323 (O_323,N_29083,N_29093);
xnor UO_324 (O_324,N_29944,N_29546);
and UO_325 (O_325,N_29266,N_29643);
or UO_326 (O_326,N_29471,N_29793);
or UO_327 (O_327,N_29685,N_29599);
and UO_328 (O_328,N_29786,N_29955);
xor UO_329 (O_329,N_29957,N_29438);
nor UO_330 (O_330,N_29116,N_29709);
or UO_331 (O_331,N_29763,N_29684);
nand UO_332 (O_332,N_29622,N_29224);
and UO_333 (O_333,N_29917,N_29240);
xnor UO_334 (O_334,N_29010,N_29479);
xnor UO_335 (O_335,N_29677,N_29859);
and UO_336 (O_336,N_29382,N_29322);
and UO_337 (O_337,N_29498,N_29305);
or UO_338 (O_338,N_29992,N_29923);
nor UO_339 (O_339,N_29127,N_29338);
xnor UO_340 (O_340,N_29219,N_29663);
xor UO_341 (O_341,N_29610,N_29207);
and UO_342 (O_342,N_29017,N_29518);
xnor UO_343 (O_343,N_29943,N_29394);
or UO_344 (O_344,N_29901,N_29854);
and UO_345 (O_345,N_29133,N_29810);
xor UO_346 (O_346,N_29580,N_29096);
nor UO_347 (O_347,N_29431,N_29443);
and UO_348 (O_348,N_29362,N_29210);
xnor UO_349 (O_349,N_29710,N_29626);
nor UO_350 (O_350,N_29452,N_29480);
and UO_351 (O_351,N_29579,N_29886);
nor UO_352 (O_352,N_29274,N_29204);
nor UO_353 (O_353,N_29032,N_29112);
nor UO_354 (O_354,N_29715,N_29962);
and UO_355 (O_355,N_29605,N_29320);
nor UO_356 (O_356,N_29681,N_29070);
or UO_357 (O_357,N_29065,N_29790);
and UO_358 (O_358,N_29164,N_29863);
or UO_359 (O_359,N_29402,N_29998);
and UO_360 (O_360,N_29733,N_29014);
or UO_361 (O_361,N_29121,N_29284);
nand UO_362 (O_362,N_29930,N_29844);
and UO_363 (O_363,N_29858,N_29344);
and UO_364 (O_364,N_29867,N_29489);
and UO_365 (O_365,N_29575,N_29766);
and UO_366 (O_366,N_29961,N_29262);
xor UO_367 (O_367,N_29792,N_29304);
xor UO_368 (O_368,N_29994,N_29444);
nor UO_369 (O_369,N_29670,N_29645);
xnor UO_370 (O_370,N_29768,N_29851);
and UO_371 (O_371,N_29312,N_29448);
and UO_372 (O_372,N_29717,N_29914);
or UO_373 (O_373,N_29020,N_29063);
xnor UO_374 (O_374,N_29393,N_29218);
nand UO_375 (O_375,N_29918,N_29829);
and UO_376 (O_376,N_29465,N_29084);
nor UO_377 (O_377,N_29798,N_29868);
nand UO_378 (O_378,N_29276,N_29895);
or UO_379 (O_379,N_29372,N_29566);
nor UO_380 (O_380,N_29462,N_29888);
xnor UO_381 (O_381,N_29232,N_29478);
nor UO_382 (O_382,N_29351,N_29328);
nand UO_383 (O_383,N_29641,N_29074);
nor UO_384 (O_384,N_29584,N_29315);
xnor UO_385 (O_385,N_29706,N_29765);
nor UO_386 (O_386,N_29835,N_29267);
nand UO_387 (O_387,N_29477,N_29924);
and UO_388 (O_388,N_29510,N_29102);
or UO_389 (O_389,N_29198,N_29987);
nand UO_390 (O_390,N_29412,N_29558);
or UO_391 (O_391,N_29155,N_29672);
or UO_392 (O_392,N_29188,N_29311);
xnor UO_393 (O_393,N_29213,N_29664);
nor UO_394 (O_394,N_29329,N_29908);
nor UO_395 (O_395,N_29588,N_29931);
nand UO_396 (O_396,N_29743,N_29220);
xor UO_397 (O_397,N_29429,N_29666);
nor UO_398 (O_398,N_29154,N_29690);
nand UO_399 (O_399,N_29736,N_29774);
and UO_400 (O_400,N_29281,N_29012);
and UO_401 (O_401,N_29387,N_29934);
nor UO_402 (O_402,N_29545,N_29332);
or UO_403 (O_403,N_29815,N_29861);
and UO_404 (O_404,N_29491,N_29655);
and UO_405 (O_405,N_29535,N_29529);
xor UO_406 (O_406,N_29150,N_29658);
or UO_407 (O_407,N_29682,N_29985);
nor UO_408 (O_408,N_29201,N_29113);
nor UO_409 (O_409,N_29508,N_29587);
nor UO_410 (O_410,N_29720,N_29636);
nor UO_411 (O_411,N_29712,N_29292);
and UO_412 (O_412,N_29034,N_29430);
and UO_413 (O_413,N_29268,N_29377);
and UO_414 (O_414,N_29702,N_29182);
nor UO_415 (O_415,N_29885,N_29441);
nand UO_416 (O_416,N_29981,N_29873);
nor UO_417 (O_417,N_29027,N_29676);
nor UO_418 (O_418,N_29871,N_29675);
nand UO_419 (O_419,N_29894,N_29047);
nor UO_420 (O_420,N_29467,N_29555);
nand UO_421 (O_421,N_29172,N_29060);
and UO_422 (O_422,N_29399,N_29104);
xnor UO_423 (O_423,N_29006,N_29261);
or UO_424 (O_424,N_29196,N_29185);
xor UO_425 (O_425,N_29986,N_29054);
or UO_426 (O_426,N_29971,N_29876);
nand UO_427 (O_427,N_29850,N_29379);
nand UO_428 (O_428,N_29563,N_29644);
or UO_429 (O_429,N_29787,N_29904);
and UO_430 (O_430,N_29126,N_29747);
or UO_431 (O_431,N_29323,N_29271);
and UO_432 (O_432,N_29978,N_29601);
nor UO_433 (O_433,N_29577,N_29585);
nand UO_434 (O_434,N_29843,N_29397);
and UO_435 (O_435,N_29174,N_29364);
xor UO_436 (O_436,N_29791,N_29673);
nand UO_437 (O_437,N_29092,N_29789);
nand UO_438 (O_438,N_29534,N_29979);
nor UO_439 (O_439,N_29408,N_29614);
nand UO_440 (O_440,N_29751,N_29881);
and UO_441 (O_441,N_29933,N_29705);
xor UO_442 (O_442,N_29067,N_29286);
and UO_443 (O_443,N_29202,N_29128);
xor UO_444 (O_444,N_29440,N_29797);
or UO_445 (O_445,N_29425,N_29852);
and UO_446 (O_446,N_29882,N_29945);
or UO_447 (O_447,N_29258,N_29134);
nand UO_448 (O_448,N_29457,N_29192);
nor UO_449 (O_449,N_29061,N_29504);
nor UO_450 (O_450,N_29840,N_29668);
xnor UO_451 (O_451,N_29779,N_29426);
nand UO_452 (O_452,N_29925,N_29517);
or UO_453 (O_453,N_29310,N_29254);
nand UO_454 (O_454,N_29938,N_29157);
nand UO_455 (O_455,N_29954,N_29422);
and UO_456 (O_456,N_29783,N_29688);
or UO_457 (O_457,N_29855,N_29691);
and UO_458 (O_458,N_29398,N_29538);
nand UO_459 (O_459,N_29974,N_29591);
nand UO_460 (O_460,N_29896,N_29199);
and UO_461 (O_461,N_29989,N_29156);
or UO_462 (O_462,N_29349,N_29653);
and UO_463 (O_463,N_29487,N_29952);
or UO_464 (O_464,N_29433,N_29963);
and UO_465 (O_465,N_29608,N_29716);
nor UO_466 (O_466,N_29294,N_29984);
nand UO_467 (O_467,N_29131,N_29388);
or UO_468 (O_468,N_29144,N_29628);
and UO_469 (O_469,N_29796,N_29434);
or UO_470 (O_470,N_29077,N_29728);
nor UO_471 (O_471,N_29511,N_29856);
xnor UO_472 (O_472,N_29181,N_29025);
nand UO_473 (O_473,N_29446,N_29630);
or UO_474 (O_474,N_29414,N_29997);
and UO_475 (O_475,N_29296,N_29100);
and UO_476 (O_476,N_29040,N_29919);
nor UO_477 (O_477,N_29044,N_29874);
nor UO_478 (O_478,N_29361,N_29817);
or UO_479 (O_479,N_29609,N_29138);
nand UO_480 (O_480,N_29809,N_29699);
nor UO_481 (O_481,N_29068,N_29488);
and UO_482 (O_482,N_29648,N_29122);
xor UO_483 (O_483,N_29623,N_29028);
or UO_484 (O_484,N_29114,N_29592);
and UO_485 (O_485,N_29977,N_29049);
xnor UO_486 (O_486,N_29884,N_29503);
or UO_487 (O_487,N_29165,N_29189);
xor UO_488 (O_488,N_29721,N_29501);
nand UO_489 (O_489,N_29951,N_29069);
or UO_490 (O_490,N_29493,N_29505);
and UO_491 (O_491,N_29149,N_29482);
xor UO_492 (O_492,N_29327,N_29698);
or UO_493 (O_493,N_29647,N_29547);
xor UO_494 (O_494,N_29445,N_29512);
nor UO_495 (O_495,N_29021,N_29366);
or UO_496 (O_496,N_29929,N_29005);
nand UO_497 (O_497,N_29662,N_29674);
nand UO_498 (O_498,N_29739,N_29160);
nand UO_499 (O_499,N_29117,N_29689);
or UO_500 (O_500,N_29336,N_29295);
xnor UO_501 (O_501,N_29367,N_29964);
or UO_502 (O_502,N_29809,N_29343);
or UO_503 (O_503,N_29710,N_29729);
or UO_504 (O_504,N_29194,N_29487);
xor UO_505 (O_505,N_29730,N_29913);
or UO_506 (O_506,N_29279,N_29832);
xor UO_507 (O_507,N_29270,N_29956);
or UO_508 (O_508,N_29931,N_29030);
xnor UO_509 (O_509,N_29555,N_29299);
and UO_510 (O_510,N_29071,N_29241);
and UO_511 (O_511,N_29602,N_29418);
nand UO_512 (O_512,N_29812,N_29727);
xnor UO_513 (O_513,N_29901,N_29531);
xor UO_514 (O_514,N_29184,N_29361);
and UO_515 (O_515,N_29799,N_29054);
or UO_516 (O_516,N_29446,N_29869);
xnor UO_517 (O_517,N_29488,N_29134);
nand UO_518 (O_518,N_29058,N_29878);
and UO_519 (O_519,N_29715,N_29196);
nor UO_520 (O_520,N_29650,N_29553);
xnor UO_521 (O_521,N_29000,N_29991);
nor UO_522 (O_522,N_29443,N_29029);
and UO_523 (O_523,N_29522,N_29912);
or UO_524 (O_524,N_29425,N_29108);
nor UO_525 (O_525,N_29635,N_29970);
nor UO_526 (O_526,N_29024,N_29311);
and UO_527 (O_527,N_29764,N_29054);
nor UO_528 (O_528,N_29546,N_29122);
nor UO_529 (O_529,N_29182,N_29039);
xor UO_530 (O_530,N_29461,N_29861);
and UO_531 (O_531,N_29721,N_29162);
nor UO_532 (O_532,N_29837,N_29946);
or UO_533 (O_533,N_29400,N_29383);
and UO_534 (O_534,N_29180,N_29951);
nand UO_535 (O_535,N_29338,N_29349);
and UO_536 (O_536,N_29911,N_29814);
xnor UO_537 (O_537,N_29530,N_29150);
xor UO_538 (O_538,N_29771,N_29420);
or UO_539 (O_539,N_29154,N_29472);
or UO_540 (O_540,N_29700,N_29994);
nor UO_541 (O_541,N_29452,N_29526);
xnor UO_542 (O_542,N_29393,N_29126);
or UO_543 (O_543,N_29429,N_29811);
nand UO_544 (O_544,N_29412,N_29624);
nor UO_545 (O_545,N_29750,N_29770);
nor UO_546 (O_546,N_29385,N_29042);
and UO_547 (O_547,N_29459,N_29864);
and UO_548 (O_548,N_29383,N_29131);
nor UO_549 (O_549,N_29316,N_29356);
or UO_550 (O_550,N_29550,N_29196);
and UO_551 (O_551,N_29874,N_29025);
or UO_552 (O_552,N_29432,N_29082);
and UO_553 (O_553,N_29290,N_29730);
nand UO_554 (O_554,N_29587,N_29355);
xor UO_555 (O_555,N_29853,N_29537);
nand UO_556 (O_556,N_29239,N_29009);
xor UO_557 (O_557,N_29405,N_29951);
nor UO_558 (O_558,N_29828,N_29095);
nand UO_559 (O_559,N_29052,N_29568);
and UO_560 (O_560,N_29116,N_29096);
nor UO_561 (O_561,N_29050,N_29502);
xor UO_562 (O_562,N_29782,N_29223);
nor UO_563 (O_563,N_29856,N_29356);
or UO_564 (O_564,N_29689,N_29681);
and UO_565 (O_565,N_29336,N_29516);
nand UO_566 (O_566,N_29675,N_29754);
nor UO_567 (O_567,N_29470,N_29248);
nand UO_568 (O_568,N_29969,N_29129);
and UO_569 (O_569,N_29124,N_29083);
and UO_570 (O_570,N_29580,N_29544);
or UO_571 (O_571,N_29604,N_29914);
or UO_572 (O_572,N_29819,N_29843);
or UO_573 (O_573,N_29340,N_29448);
nor UO_574 (O_574,N_29993,N_29514);
and UO_575 (O_575,N_29066,N_29158);
xor UO_576 (O_576,N_29177,N_29292);
nand UO_577 (O_577,N_29977,N_29655);
nand UO_578 (O_578,N_29048,N_29870);
and UO_579 (O_579,N_29720,N_29826);
nor UO_580 (O_580,N_29277,N_29627);
nor UO_581 (O_581,N_29461,N_29634);
nor UO_582 (O_582,N_29527,N_29213);
and UO_583 (O_583,N_29195,N_29644);
or UO_584 (O_584,N_29577,N_29579);
and UO_585 (O_585,N_29119,N_29675);
and UO_586 (O_586,N_29019,N_29795);
nor UO_587 (O_587,N_29318,N_29639);
nor UO_588 (O_588,N_29251,N_29719);
nor UO_589 (O_589,N_29932,N_29435);
xor UO_590 (O_590,N_29913,N_29784);
or UO_591 (O_591,N_29811,N_29583);
nor UO_592 (O_592,N_29054,N_29740);
or UO_593 (O_593,N_29097,N_29792);
xnor UO_594 (O_594,N_29340,N_29769);
nand UO_595 (O_595,N_29513,N_29226);
nor UO_596 (O_596,N_29160,N_29581);
or UO_597 (O_597,N_29053,N_29196);
xnor UO_598 (O_598,N_29188,N_29083);
nor UO_599 (O_599,N_29747,N_29911);
or UO_600 (O_600,N_29295,N_29424);
xnor UO_601 (O_601,N_29905,N_29706);
xor UO_602 (O_602,N_29910,N_29594);
and UO_603 (O_603,N_29323,N_29740);
nand UO_604 (O_604,N_29587,N_29238);
or UO_605 (O_605,N_29816,N_29298);
nand UO_606 (O_606,N_29788,N_29943);
xnor UO_607 (O_607,N_29658,N_29135);
and UO_608 (O_608,N_29717,N_29175);
and UO_609 (O_609,N_29640,N_29853);
or UO_610 (O_610,N_29352,N_29848);
nor UO_611 (O_611,N_29200,N_29015);
nand UO_612 (O_612,N_29427,N_29774);
and UO_613 (O_613,N_29299,N_29414);
xor UO_614 (O_614,N_29341,N_29867);
nor UO_615 (O_615,N_29037,N_29049);
and UO_616 (O_616,N_29606,N_29628);
or UO_617 (O_617,N_29341,N_29691);
and UO_618 (O_618,N_29317,N_29796);
nand UO_619 (O_619,N_29381,N_29882);
nand UO_620 (O_620,N_29327,N_29913);
and UO_621 (O_621,N_29316,N_29990);
nand UO_622 (O_622,N_29979,N_29831);
or UO_623 (O_623,N_29757,N_29384);
nor UO_624 (O_624,N_29523,N_29685);
and UO_625 (O_625,N_29960,N_29192);
nor UO_626 (O_626,N_29632,N_29233);
and UO_627 (O_627,N_29766,N_29242);
xor UO_628 (O_628,N_29045,N_29235);
nand UO_629 (O_629,N_29400,N_29235);
or UO_630 (O_630,N_29342,N_29948);
nor UO_631 (O_631,N_29374,N_29590);
and UO_632 (O_632,N_29666,N_29156);
xnor UO_633 (O_633,N_29795,N_29306);
nor UO_634 (O_634,N_29942,N_29983);
xnor UO_635 (O_635,N_29416,N_29334);
xor UO_636 (O_636,N_29526,N_29037);
nor UO_637 (O_637,N_29624,N_29221);
xnor UO_638 (O_638,N_29477,N_29424);
or UO_639 (O_639,N_29267,N_29984);
nor UO_640 (O_640,N_29465,N_29202);
and UO_641 (O_641,N_29598,N_29447);
or UO_642 (O_642,N_29024,N_29071);
nand UO_643 (O_643,N_29864,N_29786);
nand UO_644 (O_644,N_29561,N_29670);
nor UO_645 (O_645,N_29634,N_29664);
nand UO_646 (O_646,N_29242,N_29992);
and UO_647 (O_647,N_29858,N_29127);
nand UO_648 (O_648,N_29376,N_29127);
nor UO_649 (O_649,N_29809,N_29791);
or UO_650 (O_650,N_29228,N_29740);
nor UO_651 (O_651,N_29735,N_29586);
or UO_652 (O_652,N_29664,N_29216);
nor UO_653 (O_653,N_29150,N_29419);
nand UO_654 (O_654,N_29783,N_29533);
nor UO_655 (O_655,N_29896,N_29785);
nand UO_656 (O_656,N_29887,N_29764);
or UO_657 (O_657,N_29459,N_29646);
or UO_658 (O_658,N_29582,N_29815);
or UO_659 (O_659,N_29700,N_29650);
and UO_660 (O_660,N_29811,N_29205);
nand UO_661 (O_661,N_29658,N_29846);
nor UO_662 (O_662,N_29312,N_29849);
nor UO_663 (O_663,N_29040,N_29021);
and UO_664 (O_664,N_29497,N_29640);
nand UO_665 (O_665,N_29547,N_29257);
nand UO_666 (O_666,N_29467,N_29739);
nor UO_667 (O_667,N_29821,N_29227);
xnor UO_668 (O_668,N_29598,N_29805);
and UO_669 (O_669,N_29313,N_29619);
xor UO_670 (O_670,N_29272,N_29325);
or UO_671 (O_671,N_29613,N_29682);
and UO_672 (O_672,N_29871,N_29551);
nand UO_673 (O_673,N_29295,N_29970);
xnor UO_674 (O_674,N_29838,N_29310);
or UO_675 (O_675,N_29177,N_29920);
nand UO_676 (O_676,N_29851,N_29518);
nor UO_677 (O_677,N_29238,N_29108);
nand UO_678 (O_678,N_29975,N_29920);
or UO_679 (O_679,N_29324,N_29266);
nand UO_680 (O_680,N_29891,N_29605);
nand UO_681 (O_681,N_29005,N_29824);
or UO_682 (O_682,N_29670,N_29834);
nor UO_683 (O_683,N_29404,N_29905);
xor UO_684 (O_684,N_29412,N_29442);
xor UO_685 (O_685,N_29261,N_29170);
nor UO_686 (O_686,N_29586,N_29388);
nand UO_687 (O_687,N_29192,N_29498);
nand UO_688 (O_688,N_29455,N_29334);
or UO_689 (O_689,N_29048,N_29703);
xor UO_690 (O_690,N_29158,N_29596);
nand UO_691 (O_691,N_29202,N_29759);
xnor UO_692 (O_692,N_29659,N_29855);
nand UO_693 (O_693,N_29843,N_29446);
or UO_694 (O_694,N_29821,N_29124);
nor UO_695 (O_695,N_29909,N_29837);
nand UO_696 (O_696,N_29345,N_29960);
nor UO_697 (O_697,N_29737,N_29046);
and UO_698 (O_698,N_29675,N_29407);
nand UO_699 (O_699,N_29057,N_29348);
nor UO_700 (O_700,N_29266,N_29223);
or UO_701 (O_701,N_29459,N_29850);
and UO_702 (O_702,N_29744,N_29217);
or UO_703 (O_703,N_29070,N_29307);
and UO_704 (O_704,N_29694,N_29804);
or UO_705 (O_705,N_29060,N_29814);
or UO_706 (O_706,N_29471,N_29814);
and UO_707 (O_707,N_29616,N_29587);
xor UO_708 (O_708,N_29350,N_29256);
nor UO_709 (O_709,N_29438,N_29209);
nand UO_710 (O_710,N_29226,N_29321);
nor UO_711 (O_711,N_29839,N_29381);
xnor UO_712 (O_712,N_29467,N_29057);
xor UO_713 (O_713,N_29857,N_29292);
xnor UO_714 (O_714,N_29226,N_29533);
or UO_715 (O_715,N_29572,N_29010);
xnor UO_716 (O_716,N_29046,N_29862);
xor UO_717 (O_717,N_29037,N_29787);
xor UO_718 (O_718,N_29761,N_29139);
nand UO_719 (O_719,N_29514,N_29872);
and UO_720 (O_720,N_29688,N_29105);
or UO_721 (O_721,N_29134,N_29113);
nor UO_722 (O_722,N_29916,N_29592);
xor UO_723 (O_723,N_29494,N_29560);
or UO_724 (O_724,N_29060,N_29776);
nor UO_725 (O_725,N_29952,N_29188);
or UO_726 (O_726,N_29167,N_29882);
nor UO_727 (O_727,N_29621,N_29950);
xor UO_728 (O_728,N_29509,N_29716);
or UO_729 (O_729,N_29554,N_29288);
xnor UO_730 (O_730,N_29898,N_29916);
nor UO_731 (O_731,N_29692,N_29792);
nor UO_732 (O_732,N_29621,N_29233);
nand UO_733 (O_733,N_29327,N_29895);
and UO_734 (O_734,N_29908,N_29805);
and UO_735 (O_735,N_29837,N_29072);
nor UO_736 (O_736,N_29234,N_29283);
or UO_737 (O_737,N_29599,N_29025);
and UO_738 (O_738,N_29790,N_29580);
or UO_739 (O_739,N_29484,N_29509);
xor UO_740 (O_740,N_29950,N_29138);
xor UO_741 (O_741,N_29212,N_29169);
xnor UO_742 (O_742,N_29697,N_29487);
xor UO_743 (O_743,N_29133,N_29707);
and UO_744 (O_744,N_29731,N_29203);
or UO_745 (O_745,N_29913,N_29191);
or UO_746 (O_746,N_29072,N_29005);
xor UO_747 (O_747,N_29334,N_29818);
xor UO_748 (O_748,N_29347,N_29036);
or UO_749 (O_749,N_29639,N_29471);
xnor UO_750 (O_750,N_29810,N_29568);
nand UO_751 (O_751,N_29732,N_29155);
and UO_752 (O_752,N_29938,N_29495);
or UO_753 (O_753,N_29690,N_29997);
nand UO_754 (O_754,N_29468,N_29912);
nand UO_755 (O_755,N_29620,N_29051);
xnor UO_756 (O_756,N_29351,N_29305);
and UO_757 (O_757,N_29232,N_29335);
and UO_758 (O_758,N_29316,N_29826);
nor UO_759 (O_759,N_29334,N_29370);
or UO_760 (O_760,N_29928,N_29179);
nand UO_761 (O_761,N_29840,N_29065);
nand UO_762 (O_762,N_29808,N_29717);
and UO_763 (O_763,N_29744,N_29251);
or UO_764 (O_764,N_29558,N_29092);
nand UO_765 (O_765,N_29773,N_29248);
and UO_766 (O_766,N_29243,N_29639);
nor UO_767 (O_767,N_29522,N_29911);
nand UO_768 (O_768,N_29483,N_29068);
and UO_769 (O_769,N_29148,N_29736);
xor UO_770 (O_770,N_29442,N_29468);
nand UO_771 (O_771,N_29490,N_29113);
xor UO_772 (O_772,N_29777,N_29183);
nand UO_773 (O_773,N_29805,N_29458);
and UO_774 (O_774,N_29465,N_29825);
nor UO_775 (O_775,N_29750,N_29034);
nand UO_776 (O_776,N_29237,N_29719);
nand UO_777 (O_777,N_29887,N_29593);
or UO_778 (O_778,N_29159,N_29982);
nor UO_779 (O_779,N_29199,N_29211);
or UO_780 (O_780,N_29400,N_29012);
or UO_781 (O_781,N_29024,N_29668);
and UO_782 (O_782,N_29724,N_29675);
or UO_783 (O_783,N_29003,N_29509);
nor UO_784 (O_784,N_29032,N_29503);
or UO_785 (O_785,N_29478,N_29192);
xor UO_786 (O_786,N_29608,N_29404);
nand UO_787 (O_787,N_29917,N_29050);
and UO_788 (O_788,N_29169,N_29435);
nand UO_789 (O_789,N_29356,N_29888);
or UO_790 (O_790,N_29493,N_29387);
and UO_791 (O_791,N_29582,N_29184);
or UO_792 (O_792,N_29221,N_29897);
nor UO_793 (O_793,N_29308,N_29207);
or UO_794 (O_794,N_29562,N_29542);
nor UO_795 (O_795,N_29446,N_29633);
or UO_796 (O_796,N_29814,N_29330);
and UO_797 (O_797,N_29992,N_29989);
or UO_798 (O_798,N_29557,N_29006);
nand UO_799 (O_799,N_29516,N_29036);
and UO_800 (O_800,N_29663,N_29246);
or UO_801 (O_801,N_29847,N_29130);
nand UO_802 (O_802,N_29027,N_29465);
xor UO_803 (O_803,N_29272,N_29322);
nand UO_804 (O_804,N_29501,N_29479);
xor UO_805 (O_805,N_29082,N_29071);
and UO_806 (O_806,N_29641,N_29696);
nand UO_807 (O_807,N_29945,N_29156);
nand UO_808 (O_808,N_29801,N_29499);
or UO_809 (O_809,N_29541,N_29605);
nor UO_810 (O_810,N_29013,N_29109);
and UO_811 (O_811,N_29323,N_29554);
and UO_812 (O_812,N_29948,N_29598);
xor UO_813 (O_813,N_29553,N_29841);
or UO_814 (O_814,N_29851,N_29852);
nand UO_815 (O_815,N_29436,N_29634);
and UO_816 (O_816,N_29041,N_29684);
nor UO_817 (O_817,N_29414,N_29740);
nand UO_818 (O_818,N_29564,N_29898);
nand UO_819 (O_819,N_29105,N_29036);
and UO_820 (O_820,N_29266,N_29697);
nand UO_821 (O_821,N_29705,N_29520);
and UO_822 (O_822,N_29470,N_29839);
xnor UO_823 (O_823,N_29842,N_29346);
or UO_824 (O_824,N_29171,N_29701);
and UO_825 (O_825,N_29466,N_29088);
nand UO_826 (O_826,N_29762,N_29508);
and UO_827 (O_827,N_29242,N_29372);
nand UO_828 (O_828,N_29887,N_29197);
and UO_829 (O_829,N_29801,N_29718);
xnor UO_830 (O_830,N_29347,N_29249);
nor UO_831 (O_831,N_29002,N_29944);
or UO_832 (O_832,N_29001,N_29717);
or UO_833 (O_833,N_29230,N_29405);
nor UO_834 (O_834,N_29636,N_29694);
nand UO_835 (O_835,N_29504,N_29508);
xnor UO_836 (O_836,N_29012,N_29543);
nand UO_837 (O_837,N_29961,N_29228);
nand UO_838 (O_838,N_29432,N_29628);
and UO_839 (O_839,N_29367,N_29984);
or UO_840 (O_840,N_29380,N_29294);
xor UO_841 (O_841,N_29118,N_29635);
or UO_842 (O_842,N_29279,N_29313);
xnor UO_843 (O_843,N_29992,N_29442);
nor UO_844 (O_844,N_29308,N_29021);
nor UO_845 (O_845,N_29554,N_29892);
and UO_846 (O_846,N_29250,N_29765);
nand UO_847 (O_847,N_29269,N_29802);
xnor UO_848 (O_848,N_29368,N_29776);
nor UO_849 (O_849,N_29271,N_29109);
nor UO_850 (O_850,N_29669,N_29233);
and UO_851 (O_851,N_29864,N_29540);
or UO_852 (O_852,N_29444,N_29751);
xnor UO_853 (O_853,N_29964,N_29592);
nor UO_854 (O_854,N_29448,N_29251);
nor UO_855 (O_855,N_29110,N_29443);
nor UO_856 (O_856,N_29086,N_29884);
or UO_857 (O_857,N_29684,N_29811);
or UO_858 (O_858,N_29373,N_29485);
xnor UO_859 (O_859,N_29882,N_29848);
nor UO_860 (O_860,N_29462,N_29673);
or UO_861 (O_861,N_29994,N_29377);
or UO_862 (O_862,N_29481,N_29285);
xnor UO_863 (O_863,N_29227,N_29881);
and UO_864 (O_864,N_29949,N_29238);
nand UO_865 (O_865,N_29913,N_29088);
or UO_866 (O_866,N_29227,N_29296);
and UO_867 (O_867,N_29379,N_29692);
xnor UO_868 (O_868,N_29647,N_29843);
nand UO_869 (O_869,N_29352,N_29532);
or UO_870 (O_870,N_29552,N_29029);
or UO_871 (O_871,N_29128,N_29923);
nor UO_872 (O_872,N_29785,N_29875);
nand UO_873 (O_873,N_29020,N_29961);
nor UO_874 (O_874,N_29897,N_29567);
nor UO_875 (O_875,N_29285,N_29323);
nor UO_876 (O_876,N_29141,N_29098);
and UO_877 (O_877,N_29251,N_29055);
nand UO_878 (O_878,N_29228,N_29889);
nand UO_879 (O_879,N_29150,N_29868);
nor UO_880 (O_880,N_29465,N_29372);
or UO_881 (O_881,N_29024,N_29657);
or UO_882 (O_882,N_29868,N_29486);
nand UO_883 (O_883,N_29860,N_29713);
nor UO_884 (O_884,N_29964,N_29623);
nor UO_885 (O_885,N_29579,N_29468);
or UO_886 (O_886,N_29889,N_29764);
nor UO_887 (O_887,N_29148,N_29513);
xor UO_888 (O_888,N_29879,N_29128);
and UO_889 (O_889,N_29920,N_29007);
xnor UO_890 (O_890,N_29124,N_29345);
nor UO_891 (O_891,N_29073,N_29283);
and UO_892 (O_892,N_29861,N_29190);
nand UO_893 (O_893,N_29881,N_29006);
or UO_894 (O_894,N_29628,N_29892);
nor UO_895 (O_895,N_29150,N_29278);
and UO_896 (O_896,N_29777,N_29848);
or UO_897 (O_897,N_29663,N_29216);
nand UO_898 (O_898,N_29077,N_29469);
xnor UO_899 (O_899,N_29180,N_29422);
nor UO_900 (O_900,N_29052,N_29946);
xor UO_901 (O_901,N_29421,N_29457);
nor UO_902 (O_902,N_29096,N_29353);
nand UO_903 (O_903,N_29141,N_29704);
nand UO_904 (O_904,N_29920,N_29240);
nand UO_905 (O_905,N_29908,N_29158);
or UO_906 (O_906,N_29785,N_29947);
nand UO_907 (O_907,N_29050,N_29306);
nand UO_908 (O_908,N_29471,N_29257);
nand UO_909 (O_909,N_29038,N_29620);
nand UO_910 (O_910,N_29428,N_29523);
xnor UO_911 (O_911,N_29811,N_29659);
nand UO_912 (O_912,N_29488,N_29383);
xor UO_913 (O_913,N_29888,N_29632);
xor UO_914 (O_914,N_29763,N_29873);
or UO_915 (O_915,N_29022,N_29448);
and UO_916 (O_916,N_29599,N_29639);
nand UO_917 (O_917,N_29656,N_29708);
or UO_918 (O_918,N_29066,N_29748);
xor UO_919 (O_919,N_29755,N_29341);
nand UO_920 (O_920,N_29196,N_29541);
nand UO_921 (O_921,N_29189,N_29041);
nand UO_922 (O_922,N_29460,N_29262);
xor UO_923 (O_923,N_29534,N_29010);
nor UO_924 (O_924,N_29873,N_29193);
and UO_925 (O_925,N_29684,N_29898);
nor UO_926 (O_926,N_29480,N_29614);
nand UO_927 (O_927,N_29994,N_29465);
xnor UO_928 (O_928,N_29921,N_29545);
or UO_929 (O_929,N_29335,N_29773);
and UO_930 (O_930,N_29801,N_29906);
or UO_931 (O_931,N_29629,N_29021);
nor UO_932 (O_932,N_29636,N_29265);
nand UO_933 (O_933,N_29078,N_29679);
nand UO_934 (O_934,N_29734,N_29233);
nor UO_935 (O_935,N_29645,N_29193);
nor UO_936 (O_936,N_29328,N_29043);
xnor UO_937 (O_937,N_29014,N_29133);
nor UO_938 (O_938,N_29009,N_29240);
nand UO_939 (O_939,N_29389,N_29140);
nand UO_940 (O_940,N_29277,N_29084);
xor UO_941 (O_941,N_29271,N_29669);
and UO_942 (O_942,N_29060,N_29445);
or UO_943 (O_943,N_29548,N_29338);
and UO_944 (O_944,N_29434,N_29595);
or UO_945 (O_945,N_29921,N_29102);
or UO_946 (O_946,N_29818,N_29715);
xnor UO_947 (O_947,N_29210,N_29452);
and UO_948 (O_948,N_29356,N_29762);
or UO_949 (O_949,N_29049,N_29166);
xor UO_950 (O_950,N_29328,N_29876);
or UO_951 (O_951,N_29639,N_29230);
nor UO_952 (O_952,N_29433,N_29127);
nand UO_953 (O_953,N_29133,N_29706);
xor UO_954 (O_954,N_29740,N_29297);
nor UO_955 (O_955,N_29133,N_29795);
and UO_956 (O_956,N_29719,N_29888);
or UO_957 (O_957,N_29161,N_29158);
nand UO_958 (O_958,N_29329,N_29328);
nand UO_959 (O_959,N_29326,N_29246);
or UO_960 (O_960,N_29445,N_29067);
nor UO_961 (O_961,N_29631,N_29227);
or UO_962 (O_962,N_29298,N_29800);
xnor UO_963 (O_963,N_29119,N_29888);
nand UO_964 (O_964,N_29703,N_29040);
nand UO_965 (O_965,N_29050,N_29296);
or UO_966 (O_966,N_29400,N_29366);
xnor UO_967 (O_967,N_29078,N_29943);
nor UO_968 (O_968,N_29279,N_29883);
xnor UO_969 (O_969,N_29960,N_29702);
nand UO_970 (O_970,N_29847,N_29472);
xnor UO_971 (O_971,N_29057,N_29822);
nand UO_972 (O_972,N_29021,N_29818);
xnor UO_973 (O_973,N_29854,N_29006);
or UO_974 (O_974,N_29658,N_29255);
xnor UO_975 (O_975,N_29487,N_29466);
xor UO_976 (O_976,N_29684,N_29900);
nor UO_977 (O_977,N_29938,N_29788);
xor UO_978 (O_978,N_29307,N_29297);
nor UO_979 (O_979,N_29436,N_29086);
nor UO_980 (O_980,N_29588,N_29587);
nand UO_981 (O_981,N_29076,N_29747);
nand UO_982 (O_982,N_29834,N_29153);
nor UO_983 (O_983,N_29807,N_29207);
xnor UO_984 (O_984,N_29998,N_29612);
nor UO_985 (O_985,N_29751,N_29118);
and UO_986 (O_986,N_29320,N_29245);
or UO_987 (O_987,N_29910,N_29603);
nand UO_988 (O_988,N_29493,N_29096);
or UO_989 (O_989,N_29881,N_29430);
xor UO_990 (O_990,N_29418,N_29756);
or UO_991 (O_991,N_29265,N_29690);
or UO_992 (O_992,N_29917,N_29441);
and UO_993 (O_993,N_29400,N_29164);
or UO_994 (O_994,N_29302,N_29902);
nor UO_995 (O_995,N_29374,N_29155);
and UO_996 (O_996,N_29895,N_29717);
nand UO_997 (O_997,N_29213,N_29733);
and UO_998 (O_998,N_29657,N_29787);
nand UO_999 (O_999,N_29313,N_29762);
nand UO_1000 (O_1000,N_29014,N_29485);
nand UO_1001 (O_1001,N_29035,N_29615);
nor UO_1002 (O_1002,N_29067,N_29590);
or UO_1003 (O_1003,N_29271,N_29244);
and UO_1004 (O_1004,N_29601,N_29772);
xnor UO_1005 (O_1005,N_29303,N_29019);
nor UO_1006 (O_1006,N_29652,N_29683);
xnor UO_1007 (O_1007,N_29433,N_29739);
nand UO_1008 (O_1008,N_29446,N_29609);
and UO_1009 (O_1009,N_29824,N_29319);
nor UO_1010 (O_1010,N_29592,N_29673);
nand UO_1011 (O_1011,N_29690,N_29776);
or UO_1012 (O_1012,N_29961,N_29548);
or UO_1013 (O_1013,N_29343,N_29549);
or UO_1014 (O_1014,N_29810,N_29910);
or UO_1015 (O_1015,N_29941,N_29837);
and UO_1016 (O_1016,N_29404,N_29998);
and UO_1017 (O_1017,N_29916,N_29293);
or UO_1018 (O_1018,N_29072,N_29532);
and UO_1019 (O_1019,N_29841,N_29593);
nor UO_1020 (O_1020,N_29393,N_29435);
or UO_1021 (O_1021,N_29534,N_29950);
nor UO_1022 (O_1022,N_29544,N_29546);
nand UO_1023 (O_1023,N_29108,N_29510);
or UO_1024 (O_1024,N_29230,N_29119);
and UO_1025 (O_1025,N_29271,N_29982);
nand UO_1026 (O_1026,N_29179,N_29270);
or UO_1027 (O_1027,N_29463,N_29793);
nor UO_1028 (O_1028,N_29805,N_29310);
and UO_1029 (O_1029,N_29214,N_29480);
nand UO_1030 (O_1030,N_29746,N_29300);
or UO_1031 (O_1031,N_29806,N_29493);
and UO_1032 (O_1032,N_29793,N_29092);
and UO_1033 (O_1033,N_29724,N_29313);
xor UO_1034 (O_1034,N_29078,N_29496);
nor UO_1035 (O_1035,N_29853,N_29726);
or UO_1036 (O_1036,N_29283,N_29727);
nor UO_1037 (O_1037,N_29001,N_29964);
nor UO_1038 (O_1038,N_29581,N_29681);
xnor UO_1039 (O_1039,N_29041,N_29839);
xnor UO_1040 (O_1040,N_29389,N_29853);
and UO_1041 (O_1041,N_29026,N_29326);
and UO_1042 (O_1042,N_29507,N_29067);
and UO_1043 (O_1043,N_29059,N_29319);
xnor UO_1044 (O_1044,N_29411,N_29440);
xnor UO_1045 (O_1045,N_29920,N_29602);
or UO_1046 (O_1046,N_29645,N_29119);
xnor UO_1047 (O_1047,N_29757,N_29659);
xnor UO_1048 (O_1048,N_29961,N_29079);
or UO_1049 (O_1049,N_29137,N_29405);
nand UO_1050 (O_1050,N_29006,N_29179);
and UO_1051 (O_1051,N_29591,N_29408);
nor UO_1052 (O_1052,N_29566,N_29602);
or UO_1053 (O_1053,N_29716,N_29653);
xor UO_1054 (O_1054,N_29091,N_29762);
and UO_1055 (O_1055,N_29301,N_29407);
nand UO_1056 (O_1056,N_29415,N_29337);
nand UO_1057 (O_1057,N_29592,N_29719);
or UO_1058 (O_1058,N_29245,N_29388);
xor UO_1059 (O_1059,N_29761,N_29124);
nor UO_1060 (O_1060,N_29356,N_29345);
nor UO_1061 (O_1061,N_29556,N_29992);
or UO_1062 (O_1062,N_29210,N_29721);
xnor UO_1063 (O_1063,N_29266,N_29587);
and UO_1064 (O_1064,N_29063,N_29524);
nand UO_1065 (O_1065,N_29808,N_29430);
xnor UO_1066 (O_1066,N_29490,N_29936);
nand UO_1067 (O_1067,N_29463,N_29586);
xnor UO_1068 (O_1068,N_29853,N_29010);
or UO_1069 (O_1069,N_29698,N_29217);
or UO_1070 (O_1070,N_29200,N_29758);
nor UO_1071 (O_1071,N_29411,N_29102);
xnor UO_1072 (O_1072,N_29694,N_29900);
and UO_1073 (O_1073,N_29166,N_29116);
xor UO_1074 (O_1074,N_29600,N_29959);
or UO_1075 (O_1075,N_29714,N_29704);
and UO_1076 (O_1076,N_29474,N_29376);
nand UO_1077 (O_1077,N_29984,N_29559);
nor UO_1078 (O_1078,N_29038,N_29815);
nor UO_1079 (O_1079,N_29047,N_29893);
nor UO_1080 (O_1080,N_29226,N_29352);
or UO_1081 (O_1081,N_29730,N_29899);
nand UO_1082 (O_1082,N_29571,N_29052);
or UO_1083 (O_1083,N_29276,N_29861);
and UO_1084 (O_1084,N_29690,N_29388);
nand UO_1085 (O_1085,N_29650,N_29669);
nor UO_1086 (O_1086,N_29724,N_29571);
and UO_1087 (O_1087,N_29339,N_29453);
and UO_1088 (O_1088,N_29890,N_29271);
nand UO_1089 (O_1089,N_29442,N_29010);
and UO_1090 (O_1090,N_29380,N_29996);
nor UO_1091 (O_1091,N_29415,N_29763);
xor UO_1092 (O_1092,N_29531,N_29771);
or UO_1093 (O_1093,N_29659,N_29276);
nand UO_1094 (O_1094,N_29830,N_29196);
or UO_1095 (O_1095,N_29373,N_29814);
nor UO_1096 (O_1096,N_29961,N_29582);
xnor UO_1097 (O_1097,N_29719,N_29214);
nor UO_1098 (O_1098,N_29439,N_29759);
nor UO_1099 (O_1099,N_29730,N_29701);
and UO_1100 (O_1100,N_29436,N_29691);
nand UO_1101 (O_1101,N_29021,N_29971);
xnor UO_1102 (O_1102,N_29109,N_29869);
and UO_1103 (O_1103,N_29289,N_29270);
xnor UO_1104 (O_1104,N_29361,N_29876);
nand UO_1105 (O_1105,N_29287,N_29022);
nand UO_1106 (O_1106,N_29376,N_29249);
nor UO_1107 (O_1107,N_29764,N_29870);
or UO_1108 (O_1108,N_29269,N_29195);
xnor UO_1109 (O_1109,N_29338,N_29593);
xor UO_1110 (O_1110,N_29011,N_29221);
or UO_1111 (O_1111,N_29705,N_29413);
or UO_1112 (O_1112,N_29384,N_29369);
and UO_1113 (O_1113,N_29982,N_29110);
nand UO_1114 (O_1114,N_29896,N_29904);
nand UO_1115 (O_1115,N_29275,N_29273);
nor UO_1116 (O_1116,N_29899,N_29054);
or UO_1117 (O_1117,N_29032,N_29327);
or UO_1118 (O_1118,N_29777,N_29361);
nand UO_1119 (O_1119,N_29963,N_29450);
xnor UO_1120 (O_1120,N_29679,N_29052);
nor UO_1121 (O_1121,N_29495,N_29926);
nand UO_1122 (O_1122,N_29187,N_29107);
xor UO_1123 (O_1123,N_29089,N_29162);
xor UO_1124 (O_1124,N_29384,N_29889);
or UO_1125 (O_1125,N_29529,N_29846);
nand UO_1126 (O_1126,N_29016,N_29628);
xnor UO_1127 (O_1127,N_29529,N_29361);
nand UO_1128 (O_1128,N_29376,N_29042);
xnor UO_1129 (O_1129,N_29095,N_29067);
and UO_1130 (O_1130,N_29075,N_29166);
or UO_1131 (O_1131,N_29266,N_29721);
nor UO_1132 (O_1132,N_29236,N_29520);
xor UO_1133 (O_1133,N_29707,N_29258);
nand UO_1134 (O_1134,N_29173,N_29233);
or UO_1135 (O_1135,N_29112,N_29467);
or UO_1136 (O_1136,N_29710,N_29360);
nor UO_1137 (O_1137,N_29720,N_29135);
xor UO_1138 (O_1138,N_29206,N_29403);
or UO_1139 (O_1139,N_29472,N_29509);
nor UO_1140 (O_1140,N_29396,N_29026);
nand UO_1141 (O_1141,N_29121,N_29869);
xnor UO_1142 (O_1142,N_29563,N_29800);
xor UO_1143 (O_1143,N_29886,N_29247);
and UO_1144 (O_1144,N_29932,N_29513);
nor UO_1145 (O_1145,N_29619,N_29252);
xnor UO_1146 (O_1146,N_29526,N_29861);
nor UO_1147 (O_1147,N_29384,N_29276);
xnor UO_1148 (O_1148,N_29610,N_29582);
nand UO_1149 (O_1149,N_29982,N_29305);
nand UO_1150 (O_1150,N_29499,N_29342);
nand UO_1151 (O_1151,N_29311,N_29869);
nand UO_1152 (O_1152,N_29449,N_29005);
nand UO_1153 (O_1153,N_29309,N_29207);
nor UO_1154 (O_1154,N_29730,N_29088);
and UO_1155 (O_1155,N_29318,N_29314);
xor UO_1156 (O_1156,N_29958,N_29006);
xor UO_1157 (O_1157,N_29474,N_29496);
or UO_1158 (O_1158,N_29464,N_29899);
nor UO_1159 (O_1159,N_29474,N_29323);
xor UO_1160 (O_1160,N_29293,N_29539);
xor UO_1161 (O_1161,N_29781,N_29235);
or UO_1162 (O_1162,N_29746,N_29308);
or UO_1163 (O_1163,N_29492,N_29462);
nor UO_1164 (O_1164,N_29864,N_29161);
and UO_1165 (O_1165,N_29259,N_29171);
xnor UO_1166 (O_1166,N_29401,N_29188);
nor UO_1167 (O_1167,N_29612,N_29928);
or UO_1168 (O_1168,N_29997,N_29831);
and UO_1169 (O_1169,N_29834,N_29068);
nand UO_1170 (O_1170,N_29222,N_29167);
nor UO_1171 (O_1171,N_29759,N_29780);
and UO_1172 (O_1172,N_29252,N_29787);
nor UO_1173 (O_1173,N_29398,N_29587);
xor UO_1174 (O_1174,N_29847,N_29715);
nand UO_1175 (O_1175,N_29008,N_29715);
or UO_1176 (O_1176,N_29763,N_29166);
nand UO_1177 (O_1177,N_29640,N_29826);
nor UO_1178 (O_1178,N_29269,N_29872);
nand UO_1179 (O_1179,N_29324,N_29999);
nor UO_1180 (O_1180,N_29223,N_29841);
nor UO_1181 (O_1181,N_29858,N_29385);
nand UO_1182 (O_1182,N_29729,N_29438);
or UO_1183 (O_1183,N_29440,N_29218);
xor UO_1184 (O_1184,N_29708,N_29502);
nor UO_1185 (O_1185,N_29643,N_29840);
xor UO_1186 (O_1186,N_29232,N_29309);
nor UO_1187 (O_1187,N_29408,N_29321);
or UO_1188 (O_1188,N_29460,N_29495);
or UO_1189 (O_1189,N_29475,N_29396);
nand UO_1190 (O_1190,N_29454,N_29871);
xnor UO_1191 (O_1191,N_29057,N_29410);
xnor UO_1192 (O_1192,N_29116,N_29792);
nand UO_1193 (O_1193,N_29580,N_29878);
xor UO_1194 (O_1194,N_29459,N_29744);
or UO_1195 (O_1195,N_29371,N_29960);
xnor UO_1196 (O_1196,N_29515,N_29244);
nand UO_1197 (O_1197,N_29062,N_29121);
nor UO_1198 (O_1198,N_29847,N_29150);
nand UO_1199 (O_1199,N_29968,N_29649);
xor UO_1200 (O_1200,N_29923,N_29959);
nand UO_1201 (O_1201,N_29708,N_29260);
and UO_1202 (O_1202,N_29878,N_29328);
and UO_1203 (O_1203,N_29937,N_29901);
xor UO_1204 (O_1204,N_29686,N_29896);
and UO_1205 (O_1205,N_29605,N_29380);
nor UO_1206 (O_1206,N_29884,N_29232);
or UO_1207 (O_1207,N_29735,N_29802);
nand UO_1208 (O_1208,N_29942,N_29957);
xnor UO_1209 (O_1209,N_29495,N_29813);
nand UO_1210 (O_1210,N_29666,N_29750);
or UO_1211 (O_1211,N_29170,N_29212);
or UO_1212 (O_1212,N_29179,N_29789);
and UO_1213 (O_1213,N_29062,N_29025);
and UO_1214 (O_1214,N_29373,N_29502);
or UO_1215 (O_1215,N_29285,N_29447);
xnor UO_1216 (O_1216,N_29226,N_29552);
xor UO_1217 (O_1217,N_29375,N_29618);
xnor UO_1218 (O_1218,N_29048,N_29568);
nand UO_1219 (O_1219,N_29885,N_29331);
and UO_1220 (O_1220,N_29836,N_29726);
or UO_1221 (O_1221,N_29003,N_29566);
xor UO_1222 (O_1222,N_29162,N_29387);
xor UO_1223 (O_1223,N_29811,N_29731);
or UO_1224 (O_1224,N_29515,N_29366);
nand UO_1225 (O_1225,N_29906,N_29018);
xor UO_1226 (O_1226,N_29489,N_29908);
nand UO_1227 (O_1227,N_29294,N_29435);
xnor UO_1228 (O_1228,N_29691,N_29502);
or UO_1229 (O_1229,N_29356,N_29618);
xor UO_1230 (O_1230,N_29343,N_29240);
xnor UO_1231 (O_1231,N_29311,N_29152);
nand UO_1232 (O_1232,N_29836,N_29123);
and UO_1233 (O_1233,N_29256,N_29197);
and UO_1234 (O_1234,N_29998,N_29735);
or UO_1235 (O_1235,N_29075,N_29958);
or UO_1236 (O_1236,N_29546,N_29288);
xnor UO_1237 (O_1237,N_29603,N_29463);
nand UO_1238 (O_1238,N_29390,N_29456);
or UO_1239 (O_1239,N_29211,N_29055);
nor UO_1240 (O_1240,N_29933,N_29542);
and UO_1241 (O_1241,N_29033,N_29662);
nand UO_1242 (O_1242,N_29537,N_29192);
or UO_1243 (O_1243,N_29244,N_29424);
xnor UO_1244 (O_1244,N_29341,N_29024);
nand UO_1245 (O_1245,N_29472,N_29475);
nor UO_1246 (O_1246,N_29555,N_29739);
or UO_1247 (O_1247,N_29521,N_29581);
xnor UO_1248 (O_1248,N_29908,N_29889);
and UO_1249 (O_1249,N_29061,N_29798);
and UO_1250 (O_1250,N_29343,N_29516);
xor UO_1251 (O_1251,N_29405,N_29082);
xor UO_1252 (O_1252,N_29983,N_29070);
and UO_1253 (O_1253,N_29726,N_29768);
nand UO_1254 (O_1254,N_29219,N_29008);
nand UO_1255 (O_1255,N_29425,N_29146);
xnor UO_1256 (O_1256,N_29560,N_29752);
xor UO_1257 (O_1257,N_29256,N_29385);
xnor UO_1258 (O_1258,N_29058,N_29106);
nor UO_1259 (O_1259,N_29536,N_29474);
nor UO_1260 (O_1260,N_29032,N_29437);
or UO_1261 (O_1261,N_29952,N_29147);
and UO_1262 (O_1262,N_29256,N_29406);
nor UO_1263 (O_1263,N_29907,N_29524);
and UO_1264 (O_1264,N_29972,N_29760);
or UO_1265 (O_1265,N_29569,N_29450);
nor UO_1266 (O_1266,N_29544,N_29533);
nand UO_1267 (O_1267,N_29521,N_29537);
xnor UO_1268 (O_1268,N_29715,N_29283);
nor UO_1269 (O_1269,N_29900,N_29443);
nor UO_1270 (O_1270,N_29818,N_29066);
xor UO_1271 (O_1271,N_29756,N_29573);
xor UO_1272 (O_1272,N_29788,N_29733);
nand UO_1273 (O_1273,N_29352,N_29900);
xor UO_1274 (O_1274,N_29912,N_29710);
nand UO_1275 (O_1275,N_29955,N_29051);
nor UO_1276 (O_1276,N_29810,N_29215);
nand UO_1277 (O_1277,N_29711,N_29637);
nand UO_1278 (O_1278,N_29834,N_29712);
and UO_1279 (O_1279,N_29445,N_29760);
or UO_1280 (O_1280,N_29865,N_29266);
nand UO_1281 (O_1281,N_29858,N_29254);
xor UO_1282 (O_1282,N_29149,N_29170);
xnor UO_1283 (O_1283,N_29342,N_29755);
or UO_1284 (O_1284,N_29228,N_29727);
and UO_1285 (O_1285,N_29683,N_29449);
xor UO_1286 (O_1286,N_29898,N_29160);
nand UO_1287 (O_1287,N_29946,N_29443);
nor UO_1288 (O_1288,N_29333,N_29160);
nor UO_1289 (O_1289,N_29680,N_29038);
nor UO_1290 (O_1290,N_29027,N_29162);
nor UO_1291 (O_1291,N_29436,N_29717);
or UO_1292 (O_1292,N_29254,N_29896);
and UO_1293 (O_1293,N_29739,N_29518);
or UO_1294 (O_1294,N_29099,N_29287);
or UO_1295 (O_1295,N_29148,N_29106);
nand UO_1296 (O_1296,N_29478,N_29221);
xor UO_1297 (O_1297,N_29829,N_29687);
or UO_1298 (O_1298,N_29782,N_29152);
xnor UO_1299 (O_1299,N_29161,N_29771);
xnor UO_1300 (O_1300,N_29987,N_29385);
or UO_1301 (O_1301,N_29809,N_29646);
and UO_1302 (O_1302,N_29874,N_29601);
xor UO_1303 (O_1303,N_29190,N_29535);
and UO_1304 (O_1304,N_29819,N_29289);
nor UO_1305 (O_1305,N_29490,N_29252);
nand UO_1306 (O_1306,N_29970,N_29354);
xnor UO_1307 (O_1307,N_29730,N_29079);
or UO_1308 (O_1308,N_29914,N_29248);
nand UO_1309 (O_1309,N_29908,N_29905);
or UO_1310 (O_1310,N_29204,N_29649);
xnor UO_1311 (O_1311,N_29511,N_29268);
nand UO_1312 (O_1312,N_29519,N_29861);
and UO_1313 (O_1313,N_29781,N_29722);
nor UO_1314 (O_1314,N_29071,N_29587);
or UO_1315 (O_1315,N_29590,N_29379);
or UO_1316 (O_1316,N_29833,N_29187);
and UO_1317 (O_1317,N_29885,N_29187);
and UO_1318 (O_1318,N_29488,N_29197);
nand UO_1319 (O_1319,N_29623,N_29704);
xnor UO_1320 (O_1320,N_29995,N_29690);
or UO_1321 (O_1321,N_29853,N_29470);
or UO_1322 (O_1322,N_29379,N_29520);
and UO_1323 (O_1323,N_29864,N_29062);
xnor UO_1324 (O_1324,N_29488,N_29090);
nor UO_1325 (O_1325,N_29072,N_29997);
or UO_1326 (O_1326,N_29807,N_29562);
xor UO_1327 (O_1327,N_29725,N_29071);
or UO_1328 (O_1328,N_29390,N_29599);
xor UO_1329 (O_1329,N_29604,N_29816);
nor UO_1330 (O_1330,N_29801,N_29230);
xor UO_1331 (O_1331,N_29657,N_29793);
and UO_1332 (O_1332,N_29863,N_29015);
or UO_1333 (O_1333,N_29219,N_29511);
nand UO_1334 (O_1334,N_29408,N_29740);
and UO_1335 (O_1335,N_29043,N_29679);
nand UO_1336 (O_1336,N_29635,N_29233);
xnor UO_1337 (O_1337,N_29656,N_29289);
nor UO_1338 (O_1338,N_29163,N_29557);
or UO_1339 (O_1339,N_29623,N_29141);
nor UO_1340 (O_1340,N_29490,N_29084);
or UO_1341 (O_1341,N_29140,N_29098);
xor UO_1342 (O_1342,N_29620,N_29362);
and UO_1343 (O_1343,N_29613,N_29572);
or UO_1344 (O_1344,N_29562,N_29398);
or UO_1345 (O_1345,N_29968,N_29722);
or UO_1346 (O_1346,N_29021,N_29936);
nor UO_1347 (O_1347,N_29315,N_29526);
nand UO_1348 (O_1348,N_29048,N_29044);
xnor UO_1349 (O_1349,N_29539,N_29227);
or UO_1350 (O_1350,N_29499,N_29704);
xnor UO_1351 (O_1351,N_29327,N_29798);
or UO_1352 (O_1352,N_29439,N_29939);
or UO_1353 (O_1353,N_29543,N_29449);
nor UO_1354 (O_1354,N_29280,N_29214);
nor UO_1355 (O_1355,N_29875,N_29938);
nand UO_1356 (O_1356,N_29895,N_29306);
nor UO_1357 (O_1357,N_29197,N_29352);
and UO_1358 (O_1358,N_29336,N_29963);
or UO_1359 (O_1359,N_29483,N_29415);
or UO_1360 (O_1360,N_29459,N_29705);
or UO_1361 (O_1361,N_29596,N_29632);
nor UO_1362 (O_1362,N_29198,N_29401);
and UO_1363 (O_1363,N_29488,N_29712);
nor UO_1364 (O_1364,N_29145,N_29708);
nand UO_1365 (O_1365,N_29095,N_29513);
xnor UO_1366 (O_1366,N_29511,N_29030);
and UO_1367 (O_1367,N_29313,N_29275);
or UO_1368 (O_1368,N_29085,N_29686);
or UO_1369 (O_1369,N_29738,N_29774);
and UO_1370 (O_1370,N_29151,N_29791);
nor UO_1371 (O_1371,N_29796,N_29478);
or UO_1372 (O_1372,N_29167,N_29454);
or UO_1373 (O_1373,N_29210,N_29832);
and UO_1374 (O_1374,N_29382,N_29080);
or UO_1375 (O_1375,N_29496,N_29376);
nor UO_1376 (O_1376,N_29069,N_29455);
and UO_1377 (O_1377,N_29572,N_29153);
nand UO_1378 (O_1378,N_29091,N_29617);
and UO_1379 (O_1379,N_29911,N_29673);
or UO_1380 (O_1380,N_29072,N_29043);
or UO_1381 (O_1381,N_29279,N_29860);
xor UO_1382 (O_1382,N_29066,N_29328);
nor UO_1383 (O_1383,N_29273,N_29585);
nor UO_1384 (O_1384,N_29026,N_29852);
nor UO_1385 (O_1385,N_29802,N_29838);
xor UO_1386 (O_1386,N_29053,N_29533);
nor UO_1387 (O_1387,N_29830,N_29839);
nor UO_1388 (O_1388,N_29189,N_29650);
or UO_1389 (O_1389,N_29737,N_29256);
nor UO_1390 (O_1390,N_29145,N_29602);
or UO_1391 (O_1391,N_29115,N_29849);
nand UO_1392 (O_1392,N_29510,N_29348);
and UO_1393 (O_1393,N_29190,N_29357);
xor UO_1394 (O_1394,N_29298,N_29260);
nor UO_1395 (O_1395,N_29533,N_29837);
nor UO_1396 (O_1396,N_29123,N_29327);
or UO_1397 (O_1397,N_29559,N_29340);
or UO_1398 (O_1398,N_29768,N_29467);
and UO_1399 (O_1399,N_29838,N_29323);
nor UO_1400 (O_1400,N_29969,N_29280);
nand UO_1401 (O_1401,N_29213,N_29095);
or UO_1402 (O_1402,N_29412,N_29417);
xnor UO_1403 (O_1403,N_29147,N_29733);
xnor UO_1404 (O_1404,N_29455,N_29749);
or UO_1405 (O_1405,N_29509,N_29566);
and UO_1406 (O_1406,N_29143,N_29939);
and UO_1407 (O_1407,N_29328,N_29833);
xnor UO_1408 (O_1408,N_29875,N_29119);
and UO_1409 (O_1409,N_29724,N_29239);
or UO_1410 (O_1410,N_29056,N_29527);
nand UO_1411 (O_1411,N_29473,N_29876);
and UO_1412 (O_1412,N_29675,N_29191);
nand UO_1413 (O_1413,N_29057,N_29645);
nand UO_1414 (O_1414,N_29731,N_29010);
and UO_1415 (O_1415,N_29753,N_29175);
xor UO_1416 (O_1416,N_29978,N_29135);
and UO_1417 (O_1417,N_29370,N_29612);
or UO_1418 (O_1418,N_29361,N_29580);
nor UO_1419 (O_1419,N_29269,N_29510);
nand UO_1420 (O_1420,N_29026,N_29483);
nor UO_1421 (O_1421,N_29177,N_29996);
nand UO_1422 (O_1422,N_29189,N_29620);
or UO_1423 (O_1423,N_29428,N_29297);
xnor UO_1424 (O_1424,N_29303,N_29789);
nor UO_1425 (O_1425,N_29365,N_29756);
and UO_1426 (O_1426,N_29341,N_29975);
xor UO_1427 (O_1427,N_29888,N_29333);
and UO_1428 (O_1428,N_29074,N_29198);
nor UO_1429 (O_1429,N_29285,N_29952);
xnor UO_1430 (O_1430,N_29627,N_29133);
or UO_1431 (O_1431,N_29498,N_29625);
or UO_1432 (O_1432,N_29751,N_29397);
and UO_1433 (O_1433,N_29132,N_29149);
or UO_1434 (O_1434,N_29957,N_29968);
nor UO_1435 (O_1435,N_29885,N_29927);
or UO_1436 (O_1436,N_29891,N_29515);
nand UO_1437 (O_1437,N_29727,N_29761);
xnor UO_1438 (O_1438,N_29927,N_29249);
and UO_1439 (O_1439,N_29725,N_29373);
nand UO_1440 (O_1440,N_29867,N_29063);
nor UO_1441 (O_1441,N_29120,N_29304);
nand UO_1442 (O_1442,N_29406,N_29900);
or UO_1443 (O_1443,N_29137,N_29037);
xor UO_1444 (O_1444,N_29701,N_29789);
and UO_1445 (O_1445,N_29904,N_29546);
nor UO_1446 (O_1446,N_29927,N_29908);
nor UO_1447 (O_1447,N_29030,N_29775);
or UO_1448 (O_1448,N_29118,N_29763);
nand UO_1449 (O_1449,N_29186,N_29472);
nor UO_1450 (O_1450,N_29749,N_29953);
xnor UO_1451 (O_1451,N_29986,N_29306);
nand UO_1452 (O_1452,N_29857,N_29054);
or UO_1453 (O_1453,N_29088,N_29026);
and UO_1454 (O_1454,N_29109,N_29495);
nor UO_1455 (O_1455,N_29126,N_29057);
and UO_1456 (O_1456,N_29307,N_29156);
and UO_1457 (O_1457,N_29924,N_29255);
nand UO_1458 (O_1458,N_29837,N_29374);
xnor UO_1459 (O_1459,N_29233,N_29476);
nand UO_1460 (O_1460,N_29510,N_29540);
nand UO_1461 (O_1461,N_29352,N_29239);
xnor UO_1462 (O_1462,N_29704,N_29874);
and UO_1463 (O_1463,N_29709,N_29982);
and UO_1464 (O_1464,N_29854,N_29975);
or UO_1465 (O_1465,N_29352,N_29150);
nor UO_1466 (O_1466,N_29061,N_29123);
nand UO_1467 (O_1467,N_29589,N_29370);
nor UO_1468 (O_1468,N_29633,N_29409);
nor UO_1469 (O_1469,N_29066,N_29776);
or UO_1470 (O_1470,N_29248,N_29204);
nor UO_1471 (O_1471,N_29679,N_29177);
or UO_1472 (O_1472,N_29501,N_29032);
xnor UO_1473 (O_1473,N_29233,N_29300);
nand UO_1474 (O_1474,N_29519,N_29696);
or UO_1475 (O_1475,N_29177,N_29571);
nand UO_1476 (O_1476,N_29831,N_29002);
or UO_1477 (O_1477,N_29431,N_29184);
xnor UO_1478 (O_1478,N_29620,N_29658);
or UO_1479 (O_1479,N_29489,N_29146);
nor UO_1480 (O_1480,N_29542,N_29301);
nor UO_1481 (O_1481,N_29022,N_29178);
nor UO_1482 (O_1482,N_29420,N_29956);
xor UO_1483 (O_1483,N_29191,N_29438);
or UO_1484 (O_1484,N_29681,N_29163);
or UO_1485 (O_1485,N_29838,N_29544);
nand UO_1486 (O_1486,N_29428,N_29643);
nand UO_1487 (O_1487,N_29468,N_29015);
xnor UO_1488 (O_1488,N_29022,N_29183);
nand UO_1489 (O_1489,N_29392,N_29563);
nand UO_1490 (O_1490,N_29402,N_29254);
nor UO_1491 (O_1491,N_29439,N_29440);
nor UO_1492 (O_1492,N_29159,N_29701);
nor UO_1493 (O_1493,N_29648,N_29538);
nand UO_1494 (O_1494,N_29883,N_29066);
xnor UO_1495 (O_1495,N_29344,N_29070);
xnor UO_1496 (O_1496,N_29571,N_29466);
and UO_1497 (O_1497,N_29456,N_29654);
and UO_1498 (O_1498,N_29779,N_29325);
or UO_1499 (O_1499,N_29730,N_29338);
nor UO_1500 (O_1500,N_29129,N_29949);
nand UO_1501 (O_1501,N_29510,N_29935);
xor UO_1502 (O_1502,N_29277,N_29653);
xor UO_1503 (O_1503,N_29847,N_29450);
and UO_1504 (O_1504,N_29199,N_29434);
or UO_1505 (O_1505,N_29288,N_29361);
nand UO_1506 (O_1506,N_29857,N_29239);
or UO_1507 (O_1507,N_29598,N_29672);
and UO_1508 (O_1508,N_29273,N_29022);
nor UO_1509 (O_1509,N_29883,N_29635);
nand UO_1510 (O_1510,N_29223,N_29757);
xnor UO_1511 (O_1511,N_29602,N_29620);
or UO_1512 (O_1512,N_29276,N_29613);
and UO_1513 (O_1513,N_29345,N_29888);
nor UO_1514 (O_1514,N_29213,N_29826);
and UO_1515 (O_1515,N_29299,N_29489);
nor UO_1516 (O_1516,N_29301,N_29127);
and UO_1517 (O_1517,N_29049,N_29479);
xor UO_1518 (O_1518,N_29623,N_29953);
nor UO_1519 (O_1519,N_29712,N_29221);
or UO_1520 (O_1520,N_29792,N_29812);
nor UO_1521 (O_1521,N_29967,N_29175);
xnor UO_1522 (O_1522,N_29624,N_29388);
and UO_1523 (O_1523,N_29817,N_29568);
or UO_1524 (O_1524,N_29164,N_29647);
nand UO_1525 (O_1525,N_29550,N_29597);
xnor UO_1526 (O_1526,N_29643,N_29834);
xnor UO_1527 (O_1527,N_29541,N_29553);
xor UO_1528 (O_1528,N_29311,N_29782);
or UO_1529 (O_1529,N_29799,N_29051);
nand UO_1530 (O_1530,N_29762,N_29185);
and UO_1531 (O_1531,N_29643,N_29425);
xor UO_1532 (O_1532,N_29729,N_29127);
nand UO_1533 (O_1533,N_29524,N_29270);
and UO_1534 (O_1534,N_29478,N_29448);
and UO_1535 (O_1535,N_29669,N_29761);
xor UO_1536 (O_1536,N_29687,N_29177);
nor UO_1537 (O_1537,N_29231,N_29990);
nand UO_1538 (O_1538,N_29159,N_29222);
nand UO_1539 (O_1539,N_29069,N_29195);
and UO_1540 (O_1540,N_29447,N_29854);
or UO_1541 (O_1541,N_29551,N_29193);
nand UO_1542 (O_1542,N_29280,N_29853);
nand UO_1543 (O_1543,N_29898,N_29410);
and UO_1544 (O_1544,N_29071,N_29075);
and UO_1545 (O_1545,N_29313,N_29769);
nand UO_1546 (O_1546,N_29168,N_29708);
nor UO_1547 (O_1547,N_29685,N_29386);
nor UO_1548 (O_1548,N_29740,N_29384);
nor UO_1549 (O_1549,N_29392,N_29815);
nor UO_1550 (O_1550,N_29402,N_29932);
and UO_1551 (O_1551,N_29282,N_29047);
nor UO_1552 (O_1552,N_29428,N_29302);
xnor UO_1553 (O_1553,N_29150,N_29262);
or UO_1554 (O_1554,N_29564,N_29010);
or UO_1555 (O_1555,N_29019,N_29971);
nand UO_1556 (O_1556,N_29241,N_29616);
or UO_1557 (O_1557,N_29060,N_29447);
nand UO_1558 (O_1558,N_29559,N_29741);
xnor UO_1559 (O_1559,N_29544,N_29569);
nor UO_1560 (O_1560,N_29554,N_29728);
and UO_1561 (O_1561,N_29977,N_29133);
and UO_1562 (O_1562,N_29707,N_29245);
nand UO_1563 (O_1563,N_29076,N_29341);
or UO_1564 (O_1564,N_29554,N_29739);
and UO_1565 (O_1565,N_29493,N_29376);
nand UO_1566 (O_1566,N_29509,N_29799);
and UO_1567 (O_1567,N_29488,N_29096);
and UO_1568 (O_1568,N_29671,N_29192);
nor UO_1569 (O_1569,N_29856,N_29044);
nand UO_1570 (O_1570,N_29491,N_29321);
nand UO_1571 (O_1571,N_29936,N_29733);
xor UO_1572 (O_1572,N_29844,N_29052);
or UO_1573 (O_1573,N_29954,N_29046);
nor UO_1574 (O_1574,N_29661,N_29395);
nand UO_1575 (O_1575,N_29484,N_29899);
nand UO_1576 (O_1576,N_29151,N_29958);
and UO_1577 (O_1577,N_29400,N_29415);
xor UO_1578 (O_1578,N_29237,N_29102);
nor UO_1579 (O_1579,N_29005,N_29491);
nor UO_1580 (O_1580,N_29766,N_29808);
xnor UO_1581 (O_1581,N_29428,N_29309);
nor UO_1582 (O_1582,N_29179,N_29876);
nand UO_1583 (O_1583,N_29002,N_29629);
or UO_1584 (O_1584,N_29565,N_29320);
nor UO_1585 (O_1585,N_29417,N_29549);
nand UO_1586 (O_1586,N_29463,N_29439);
nand UO_1587 (O_1587,N_29781,N_29811);
and UO_1588 (O_1588,N_29054,N_29605);
nand UO_1589 (O_1589,N_29963,N_29849);
xnor UO_1590 (O_1590,N_29993,N_29194);
xor UO_1591 (O_1591,N_29643,N_29525);
nand UO_1592 (O_1592,N_29807,N_29115);
or UO_1593 (O_1593,N_29301,N_29147);
and UO_1594 (O_1594,N_29064,N_29833);
nand UO_1595 (O_1595,N_29810,N_29110);
nand UO_1596 (O_1596,N_29019,N_29597);
nand UO_1597 (O_1597,N_29515,N_29638);
nor UO_1598 (O_1598,N_29797,N_29519);
xnor UO_1599 (O_1599,N_29776,N_29194);
nor UO_1600 (O_1600,N_29598,N_29433);
or UO_1601 (O_1601,N_29355,N_29876);
or UO_1602 (O_1602,N_29732,N_29929);
nand UO_1603 (O_1603,N_29069,N_29221);
nor UO_1604 (O_1604,N_29185,N_29506);
or UO_1605 (O_1605,N_29304,N_29638);
nor UO_1606 (O_1606,N_29119,N_29732);
and UO_1607 (O_1607,N_29562,N_29134);
nor UO_1608 (O_1608,N_29649,N_29443);
nor UO_1609 (O_1609,N_29267,N_29000);
and UO_1610 (O_1610,N_29630,N_29723);
nor UO_1611 (O_1611,N_29254,N_29252);
nand UO_1612 (O_1612,N_29633,N_29999);
or UO_1613 (O_1613,N_29567,N_29924);
or UO_1614 (O_1614,N_29771,N_29986);
and UO_1615 (O_1615,N_29125,N_29005);
and UO_1616 (O_1616,N_29747,N_29449);
nor UO_1617 (O_1617,N_29762,N_29942);
nand UO_1618 (O_1618,N_29947,N_29046);
nor UO_1619 (O_1619,N_29238,N_29291);
nand UO_1620 (O_1620,N_29076,N_29860);
xor UO_1621 (O_1621,N_29335,N_29766);
or UO_1622 (O_1622,N_29021,N_29436);
xnor UO_1623 (O_1623,N_29009,N_29785);
nor UO_1624 (O_1624,N_29904,N_29994);
or UO_1625 (O_1625,N_29640,N_29603);
xnor UO_1626 (O_1626,N_29173,N_29186);
or UO_1627 (O_1627,N_29426,N_29270);
nand UO_1628 (O_1628,N_29426,N_29224);
xor UO_1629 (O_1629,N_29232,N_29297);
and UO_1630 (O_1630,N_29365,N_29227);
or UO_1631 (O_1631,N_29578,N_29483);
xor UO_1632 (O_1632,N_29093,N_29863);
nor UO_1633 (O_1633,N_29504,N_29474);
and UO_1634 (O_1634,N_29671,N_29279);
xor UO_1635 (O_1635,N_29944,N_29749);
nand UO_1636 (O_1636,N_29013,N_29133);
xor UO_1637 (O_1637,N_29328,N_29860);
xor UO_1638 (O_1638,N_29881,N_29190);
or UO_1639 (O_1639,N_29463,N_29139);
nor UO_1640 (O_1640,N_29670,N_29792);
or UO_1641 (O_1641,N_29234,N_29827);
and UO_1642 (O_1642,N_29949,N_29044);
and UO_1643 (O_1643,N_29884,N_29139);
or UO_1644 (O_1644,N_29284,N_29108);
xor UO_1645 (O_1645,N_29811,N_29628);
or UO_1646 (O_1646,N_29905,N_29259);
xnor UO_1647 (O_1647,N_29807,N_29182);
nor UO_1648 (O_1648,N_29247,N_29846);
nor UO_1649 (O_1649,N_29789,N_29428);
nand UO_1650 (O_1650,N_29680,N_29313);
nand UO_1651 (O_1651,N_29788,N_29497);
nor UO_1652 (O_1652,N_29450,N_29809);
or UO_1653 (O_1653,N_29486,N_29507);
and UO_1654 (O_1654,N_29788,N_29456);
xor UO_1655 (O_1655,N_29546,N_29881);
xnor UO_1656 (O_1656,N_29551,N_29206);
xor UO_1657 (O_1657,N_29282,N_29781);
nor UO_1658 (O_1658,N_29289,N_29640);
nor UO_1659 (O_1659,N_29148,N_29015);
and UO_1660 (O_1660,N_29863,N_29741);
and UO_1661 (O_1661,N_29984,N_29504);
xnor UO_1662 (O_1662,N_29390,N_29083);
or UO_1663 (O_1663,N_29667,N_29341);
nor UO_1664 (O_1664,N_29719,N_29137);
nand UO_1665 (O_1665,N_29978,N_29015);
xor UO_1666 (O_1666,N_29550,N_29818);
or UO_1667 (O_1667,N_29592,N_29716);
xnor UO_1668 (O_1668,N_29674,N_29808);
nand UO_1669 (O_1669,N_29045,N_29677);
xnor UO_1670 (O_1670,N_29034,N_29166);
nor UO_1671 (O_1671,N_29087,N_29757);
nor UO_1672 (O_1672,N_29267,N_29444);
nand UO_1673 (O_1673,N_29937,N_29585);
and UO_1674 (O_1674,N_29902,N_29841);
nand UO_1675 (O_1675,N_29335,N_29634);
and UO_1676 (O_1676,N_29366,N_29206);
xnor UO_1677 (O_1677,N_29150,N_29577);
and UO_1678 (O_1678,N_29440,N_29226);
nand UO_1679 (O_1679,N_29120,N_29394);
nand UO_1680 (O_1680,N_29393,N_29283);
and UO_1681 (O_1681,N_29892,N_29090);
nand UO_1682 (O_1682,N_29525,N_29041);
or UO_1683 (O_1683,N_29800,N_29092);
xnor UO_1684 (O_1684,N_29223,N_29080);
and UO_1685 (O_1685,N_29523,N_29881);
nand UO_1686 (O_1686,N_29883,N_29161);
nor UO_1687 (O_1687,N_29396,N_29918);
or UO_1688 (O_1688,N_29087,N_29920);
nor UO_1689 (O_1689,N_29980,N_29175);
and UO_1690 (O_1690,N_29336,N_29532);
and UO_1691 (O_1691,N_29839,N_29348);
nand UO_1692 (O_1692,N_29843,N_29005);
nand UO_1693 (O_1693,N_29929,N_29838);
xor UO_1694 (O_1694,N_29198,N_29961);
xnor UO_1695 (O_1695,N_29342,N_29270);
xnor UO_1696 (O_1696,N_29127,N_29206);
xor UO_1697 (O_1697,N_29920,N_29346);
xnor UO_1698 (O_1698,N_29485,N_29182);
nor UO_1699 (O_1699,N_29360,N_29815);
or UO_1700 (O_1700,N_29307,N_29914);
nand UO_1701 (O_1701,N_29316,N_29326);
nand UO_1702 (O_1702,N_29449,N_29839);
or UO_1703 (O_1703,N_29322,N_29723);
nand UO_1704 (O_1704,N_29701,N_29907);
nand UO_1705 (O_1705,N_29436,N_29761);
nand UO_1706 (O_1706,N_29111,N_29896);
nand UO_1707 (O_1707,N_29192,N_29690);
and UO_1708 (O_1708,N_29436,N_29030);
xnor UO_1709 (O_1709,N_29482,N_29471);
or UO_1710 (O_1710,N_29031,N_29144);
nand UO_1711 (O_1711,N_29377,N_29975);
nor UO_1712 (O_1712,N_29132,N_29640);
and UO_1713 (O_1713,N_29167,N_29606);
or UO_1714 (O_1714,N_29664,N_29925);
xor UO_1715 (O_1715,N_29489,N_29062);
and UO_1716 (O_1716,N_29033,N_29942);
or UO_1717 (O_1717,N_29057,N_29585);
and UO_1718 (O_1718,N_29176,N_29529);
nor UO_1719 (O_1719,N_29170,N_29214);
or UO_1720 (O_1720,N_29920,N_29856);
or UO_1721 (O_1721,N_29162,N_29902);
and UO_1722 (O_1722,N_29474,N_29822);
or UO_1723 (O_1723,N_29925,N_29154);
xor UO_1724 (O_1724,N_29663,N_29863);
or UO_1725 (O_1725,N_29282,N_29248);
nand UO_1726 (O_1726,N_29533,N_29326);
xor UO_1727 (O_1727,N_29412,N_29983);
and UO_1728 (O_1728,N_29134,N_29417);
or UO_1729 (O_1729,N_29267,N_29737);
or UO_1730 (O_1730,N_29269,N_29061);
nor UO_1731 (O_1731,N_29554,N_29049);
and UO_1732 (O_1732,N_29693,N_29822);
or UO_1733 (O_1733,N_29832,N_29923);
or UO_1734 (O_1734,N_29402,N_29698);
and UO_1735 (O_1735,N_29408,N_29085);
and UO_1736 (O_1736,N_29708,N_29849);
or UO_1737 (O_1737,N_29325,N_29334);
and UO_1738 (O_1738,N_29250,N_29551);
and UO_1739 (O_1739,N_29818,N_29034);
and UO_1740 (O_1740,N_29467,N_29115);
nor UO_1741 (O_1741,N_29692,N_29564);
xor UO_1742 (O_1742,N_29707,N_29290);
xor UO_1743 (O_1743,N_29412,N_29804);
nor UO_1744 (O_1744,N_29608,N_29193);
nand UO_1745 (O_1745,N_29600,N_29837);
xor UO_1746 (O_1746,N_29347,N_29770);
and UO_1747 (O_1747,N_29229,N_29522);
or UO_1748 (O_1748,N_29328,N_29929);
nor UO_1749 (O_1749,N_29518,N_29848);
nand UO_1750 (O_1750,N_29563,N_29106);
nand UO_1751 (O_1751,N_29254,N_29323);
nand UO_1752 (O_1752,N_29075,N_29167);
xnor UO_1753 (O_1753,N_29954,N_29828);
nor UO_1754 (O_1754,N_29269,N_29232);
xor UO_1755 (O_1755,N_29955,N_29589);
nand UO_1756 (O_1756,N_29074,N_29927);
and UO_1757 (O_1757,N_29826,N_29828);
nand UO_1758 (O_1758,N_29484,N_29978);
nand UO_1759 (O_1759,N_29028,N_29380);
or UO_1760 (O_1760,N_29164,N_29652);
nand UO_1761 (O_1761,N_29057,N_29123);
or UO_1762 (O_1762,N_29599,N_29466);
xor UO_1763 (O_1763,N_29577,N_29792);
nor UO_1764 (O_1764,N_29906,N_29703);
xnor UO_1765 (O_1765,N_29492,N_29780);
nor UO_1766 (O_1766,N_29389,N_29526);
or UO_1767 (O_1767,N_29420,N_29017);
nand UO_1768 (O_1768,N_29659,N_29502);
xnor UO_1769 (O_1769,N_29038,N_29084);
nand UO_1770 (O_1770,N_29283,N_29976);
or UO_1771 (O_1771,N_29375,N_29334);
xnor UO_1772 (O_1772,N_29181,N_29579);
xnor UO_1773 (O_1773,N_29690,N_29858);
xor UO_1774 (O_1774,N_29461,N_29293);
or UO_1775 (O_1775,N_29605,N_29706);
nand UO_1776 (O_1776,N_29533,N_29921);
and UO_1777 (O_1777,N_29240,N_29175);
or UO_1778 (O_1778,N_29036,N_29802);
or UO_1779 (O_1779,N_29016,N_29987);
xnor UO_1780 (O_1780,N_29961,N_29338);
or UO_1781 (O_1781,N_29483,N_29423);
nor UO_1782 (O_1782,N_29364,N_29328);
nand UO_1783 (O_1783,N_29968,N_29859);
xnor UO_1784 (O_1784,N_29366,N_29450);
nor UO_1785 (O_1785,N_29315,N_29766);
xnor UO_1786 (O_1786,N_29350,N_29922);
or UO_1787 (O_1787,N_29508,N_29899);
xnor UO_1788 (O_1788,N_29496,N_29080);
nand UO_1789 (O_1789,N_29527,N_29935);
or UO_1790 (O_1790,N_29387,N_29441);
or UO_1791 (O_1791,N_29472,N_29607);
nand UO_1792 (O_1792,N_29852,N_29378);
or UO_1793 (O_1793,N_29576,N_29433);
and UO_1794 (O_1794,N_29248,N_29681);
nor UO_1795 (O_1795,N_29873,N_29992);
or UO_1796 (O_1796,N_29175,N_29321);
or UO_1797 (O_1797,N_29049,N_29385);
and UO_1798 (O_1798,N_29341,N_29333);
and UO_1799 (O_1799,N_29352,N_29966);
nand UO_1800 (O_1800,N_29071,N_29731);
nor UO_1801 (O_1801,N_29030,N_29800);
nand UO_1802 (O_1802,N_29816,N_29410);
nor UO_1803 (O_1803,N_29401,N_29949);
and UO_1804 (O_1804,N_29416,N_29449);
nor UO_1805 (O_1805,N_29343,N_29785);
and UO_1806 (O_1806,N_29659,N_29637);
and UO_1807 (O_1807,N_29671,N_29472);
nand UO_1808 (O_1808,N_29155,N_29619);
and UO_1809 (O_1809,N_29318,N_29479);
or UO_1810 (O_1810,N_29473,N_29379);
xnor UO_1811 (O_1811,N_29663,N_29432);
xnor UO_1812 (O_1812,N_29105,N_29569);
nand UO_1813 (O_1813,N_29476,N_29193);
nand UO_1814 (O_1814,N_29651,N_29678);
and UO_1815 (O_1815,N_29275,N_29207);
or UO_1816 (O_1816,N_29888,N_29548);
nand UO_1817 (O_1817,N_29367,N_29595);
nand UO_1818 (O_1818,N_29139,N_29882);
xnor UO_1819 (O_1819,N_29189,N_29156);
and UO_1820 (O_1820,N_29792,N_29290);
nand UO_1821 (O_1821,N_29644,N_29421);
or UO_1822 (O_1822,N_29014,N_29557);
nand UO_1823 (O_1823,N_29722,N_29811);
nor UO_1824 (O_1824,N_29115,N_29707);
or UO_1825 (O_1825,N_29595,N_29146);
and UO_1826 (O_1826,N_29984,N_29809);
nor UO_1827 (O_1827,N_29025,N_29020);
and UO_1828 (O_1828,N_29910,N_29397);
nand UO_1829 (O_1829,N_29913,N_29002);
nand UO_1830 (O_1830,N_29851,N_29887);
nor UO_1831 (O_1831,N_29768,N_29186);
nor UO_1832 (O_1832,N_29956,N_29280);
nor UO_1833 (O_1833,N_29248,N_29070);
nor UO_1834 (O_1834,N_29419,N_29644);
and UO_1835 (O_1835,N_29127,N_29937);
or UO_1836 (O_1836,N_29350,N_29666);
and UO_1837 (O_1837,N_29747,N_29514);
nand UO_1838 (O_1838,N_29562,N_29685);
nor UO_1839 (O_1839,N_29353,N_29599);
nand UO_1840 (O_1840,N_29348,N_29120);
or UO_1841 (O_1841,N_29956,N_29881);
or UO_1842 (O_1842,N_29794,N_29713);
xor UO_1843 (O_1843,N_29500,N_29906);
nor UO_1844 (O_1844,N_29406,N_29040);
or UO_1845 (O_1845,N_29936,N_29791);
xnor UO_1846 (O_1846,N_29146,N_29005);
xnor UO_1847 (O_1847,N_29736,N_29317);
nor UO_1848 (O_1848,N_29035,N_29222);
or UO_1849 (O_1849,N_29290,N_29961);
xnor UO_1850 (O_1850,N_29318,N_29954);
and UO_1851 (O_1851,N_29239,N_29381);
nand UO_1852 (O_1852,N_29039,N_29216);
nand UO_1853 (O_1853,N_29631,N_29987);
and UO_1854 (O_1854,N_29048,N_29391);
xnor UO_1855 (O_1855,N_29013,N_29896);
nor UO_1856 (O_1856,N_29649,N_29961);
or UO_1857 (O_1857,N_29994,N_29353);
xor UO_1858 (O_1858,N_29459,N_29462);
or UO_1859 (O_1859,N_29906,N_29796);
or UO_1860 (O_1860,N_29740,N_29715);
or UO_1861 (O_1861,N_29866,N_29874);
xnor UO_1862 (O_1862,N_29405,N_29143);
or UO_1863 (O_1863,N_29638,N_29882);
and UO_1864 (O_1864,N_29109,N_29350);
and UO_1865 (O_1865,N_29428,N_29165);
and UO_1866 (O_1866,N_29076,N_29122);
nand UO_1867 (O_1867,N_29686,N_29525);
xor UO_1868 (O_1868,N_29958,N_29129);
or UO_1869 (O_1869,N_29832,N_29545);
nor UO_1870 (O_1870,N_29288,N_29121);
and UO_1871 (O_1871,N_29319,N_29180);
and UO_1872 (O_1872,N_29296,N_29279);
or UO_1873 (O_1873,N_29107,N_29748);
or UO_1874 (O_1874,N_29691,N_29126);
or UO_1875 (O_1875,N_29315,N_29399);
or UO_1876 (O_1876,N_29635,N_29586);
nor UO_1877 (O_1877,N_29613,N_29130);
and UO_1878 (O_1878,N_29768,N_29528);
and UO_1879 (O_1879,N_29421,N_29749);
nand UO_1880 (O_1880,N_29229,N_29772);
and UO_1881 (O_1881,N_29162,N_29796);
nand UO_1882 (O_1882,N_29679,N_29636);
or UO_1883 (O_1883,N_29021,N_29860);
or UO_1884 (O_1884,N_29564,N_29910);
and UO_1885 (O_1885,N_29746,N_29064);
nand UO_1886 (O_1886,N_29008,N_29529);
or UO_1887 (O_1887,N_29736,N_29809);
nor UO_1888 (O_1888,N_29863,N_29980);
xnor UO_1889 (O_1889,N_29514,N_29512);
nor UO_1890 (O_1890,N_29265,N_29662);
and UO_1891 (O_1891,N_29046,N_29237);
or UO_1892 (O_1892,N_29133,N_29848);
and UO_1893 (O_1893,N_29214,N_29523);
nand UO_1894 (O_1894,N_29764,N_29836);
nand UO_1895 (O_1895,N_29362,N_29933);
or UO_1896 (O_1896,N_29024,N_29155);
xnor UO_1897 (O_1897,N_29736,N_29409);
nand UO_1898 (O_1898,N_29944,N_29266);
nand UO_1899 (O_1899,N_29576,N_29742);
and UO_1900 (O_1900,N_29615,N_29590);
and UO_1901 (O_1901,N_29628,N_29502);
or UO_1902 (O_1902,N_29428,N_29847);
or UO_1903 (O_1903,N_29136,N_29141);
nand UO_1904 (O_1904,N_29539,N_29456);
or UO_1905 (O_1905,N_29242,N_29834);
nand UO_1906 (O_1906,N_29928,N_29503);
and UO_1907 (O_1907,N_29237,N_29147);
and UO_1908 (O_1908,N_29786,N_29439);
nand UO_1909 (O_1909,N_29286,N_29296);
nand UO_1910 (O_1910,N_29180,N_29131);
and UO_1911 (O_1911,N_29825,N_29377);
or UO_1912 (O_1912,N_29135,N_29701);
and UO_1913 (O_1913,N_29365,N_29471);
and UO_1914 (O_1914,N_29123,N_29618);
nand UO_1915 (O_1915,N_29504,N_29751);
or UO_1916 (O_1916,N_29467,N_29812);
or UO_1917 (O_1917,N_29391,N_29318);
and UO_1918 (O_1918,N_29088,N_29491);
xnor UO_1919 (O_1919,N_29057,N_29754);
nor UO_1920 (O_1920,N_29241,N_29040);
nand UO_1921 (O_1921,N_29545,N_29040);
nand UO_1922 (O_1922,N_29428,N_29877);
nand UO_1923 (O_1923,N_29614,N_29088);
nand UO_1924 (O_1924,N_29754,N_29263);
xnor UO_1925 (O_1925,N_29145,N_29968);
nand UO_1926 (O_1926,N_29030,N_29588);
nor UO_1927 (O_1927,N_29908,N_29246);
or UO_1928 (O_1928,N_29787,N_29997);
nand UO_1929 (O_1929,N_29499,N_29360);
xor UO_1930 (O_1930,N_29302,N_29069);
nor UO_1931 (O_1931,N_29525,N_29088);
or UO_1932 (O_1932,N_29069,N_29444);
xnor UO_1933 (O_1933,N_29068,N_29248);
nand UO_1934 (O_1934,N_29278,N_29023);
or UO_1935 (O_1935,N_29808,N_29673);
xor UO_1936 (O_1936,N_29661,N_29728);
xor UO_1937 (O_1937,N_29574,N_29679);
nor UO_1938 (O_1938,N_29018,N_29186);
nand UO_1939 (O_1939,N_29296,N_29104);
nor UO_1940 (O_1940,N_29986,N_29467);
and UO_1941 (O_1941,N_29228,N_29402);
or UO_1942 (O_1942,N_29037,N_29215);
or UO_1943 (O_1943,N_29999,N_29486);
and UO_1944 (O_1944,N_29641,N_29666);
nor UO_1945 (O_1945,N_29334,N_29852);
nand UO_1946 (O_1946,N_29489,N_29398);
or UO_1947 (O_1947,N_29039,N_29702);
nor UO_1948 (O_1948,N_29228,N_29975);
and UO_1949 (O_1949,N_29581,N_29083);
and UO_1950 (O_1950,N_29527,N_29312);
xnor UO_1951 (O_1951,N_29315,N_29555);
xnor UO_1952 (O_1952,N_29188,N_29501);
nor UO_1953 (O_1953,N_29380,N_29124);
or UO_1954 (O_1954,N_29898,N_29252);
nor UO_1955 (O_1955,N_29188,N_29712);
and UO_1956 (O_1956,N_29327,N_29144);
xor UO_1957 (O_1957,N_29335,N_29405);
and UO_1958 (O_1958,N_29970,N_29186);
and UO_1959 (O_1959,N_29204,N_29796);
or UO_1960 (O_1960,N_29877,N_29592);
or UO_1961 (O_1961,N_29904,N_29955);
nand UO_1962 (O_1962,N_29588,N_29384);
nor UO_1963 (O_1963,N_29944,N_29020);
and UO_1964 (O_1964,N_29697,N_29880);
nand UO_1965 (O_1965,N_29848,N_29878);
and UO_1966 (O_1966,N_29833,N_29572);
and UO_1967 (O_1967,N_29211,N_29390);
and UO_1968 (O_1968,N_29625,N_29411);
nand UO_1969 (O_1969,N_29637,N_29269);
or UO_1970 (O_1970,N_29701,N_29283);
nor UO_1971 (O_1971,N_29966,N_29041);
or UO_1972 (O_1972,N_29226,N_29662);
nand UO_1973 (O_1973,N_29037,N_29163);
and UO_1974 (O_1974,N_29231,N_29994);
and UO_1975 (O_1975,N_29553,N_29631);
and UO_1976 (O_1976,N_29816,N_29725);
xnor UO_1977 (O_1977,N_29089,N_29613);
or UO_1978 (O_1978,N_29556,N_29221);
nor UO_1979 (O_1979,N_29295,N_29299);
xnor UO_1980 (O_1980,N_29994,N_29396);
xor UO_1981 (O_1981,N_29669,N_29405);
or UO_1982 (O_1982,N_29505,N_29079);
or UO_1983 (O_1983,N_29473,N_29573);
nor UO_1984 (O_1984,N_29259,N_29564);
or UO_1985 (O_1985,N_29681,N_29803);
and UO_1986 (O_1986,N_29856,N_29820);
and UO_1987 (O_1987,N_29766,N_29090);
nand UO_1988 (O_1988,N_29907,N_29294);
or UO_1989 (O_1989,N_29907,N_29358);
and UO_1990 (O_1990,N_29715,N_29751);
nand UO_1991 (O_1991,N_29591,N_29685);
or UO_1992 (O_1992,N_29595,N_29389);
nor UO_1993 (O_1993,N_29821,N_29852);
nor UO_1994 (O_1994,N_29059,N_29308);
and UO_1995 (O_1995,N_29407,N_29431);
or UO_1996 (O_1996,N_29064,N_29405);
nand UO_1997 (O_1997,N_29610,N_29341);
nor UO_1998 (O_1998,N_29936,N_29802);
or UO_1999 (O_1999,N_29027,N_29970);
nor UO_2000 (O_2000,N_29419,N_29960);
or UO_2001 (O_2001,N_29609,N_29181);
nor UO_2002 (O_2002,N_29985,N_29657);
or UO_2003 (O_2003,N_29033,N_29258);
nand UO_2004 (O_2004,N_29843,N_29349);
or UO_2005 (O_2005,N_29766,N_29193);
nand UO_2006 (O_2006,N_29299,N_29564);
xor UO_2007 (O_2007,N_29068,N_29756);
xor UO_2008 (O_2008,N_29154,N_29716);
or UO_2009 (O_2009,N_29005,N_29251);
nand UO_2010 (O_2010,N_29234,N_29395);
nand UO_2011 (O_2011,N_29265,N_29613);
and UO_2012 (O_2012,N_29239,N_29137);
xnor UO_2013 (O_2013,N_29804,N_29646);
and UO_2014 (O_2014,N_29693,N_29826);
and UO_2015 (O_2015,N_29526,N_29906);
and UO_2016 (O_2016,N_29464,N_29712);
and UO_2017 (O_2017,N_29257,N_29481);
xor UO_2018 (O_2018,N_29271,N_29950);
nor UO_2019 (O_2019,N_29430,N_29514);
and UO_2020 (O_2020,N_29441,N_29218);
xnor UO_2021 (O_2021,N_29300,N_29430);
nand UO_2022 (O_2022,N_29789,N_29692);
or UO_2023 (O_2023,N_29501,N_29583);
nor UO_2024 (O_2024,N_29973,N_29117);
or UO_2025 (O_2025,N_29105,N_29091);
or UO_2026 (O_2026,N_29858,N_29329);
nor UO_2027 (O_2027,N_29593,N_29410);
or UO_2028 (O_2028,N_29530,N_29669);
nand UO_2029 (O_2029,N_29475,N_29255);
or UO_2030 (O_2030,N_29219,N_29853);
or UO_2031 (O_2031,N_29851,N_29072);
or UO_2032 (O_2032,N_29100,N_29429);
xnor UO_2033 (O_2033,N_29106,N_29364);
or UO_2034 (O_2034,N_29591,N_29607);
and UO_2035 (O_2035,N_29009,N_29142);
and UO_2036 (O_2036,N_29658,N_29661);
nor UO_2037 (O_2037,N_29720,N_29742);
and UO_2038 (O_2038,N_29554,N_29640);
nor UO_2039 (O_2039,N_29050,N_29461);
xor UO_2040 (O_2040,N_29165,N_29069);
nand UO_2041 (O_2041,N_29544,N_29043);
or UO_2042 (O_2042,N_29199,N_29035);
or UO_2043 (O_2043,N_29869,N_29646);
nor UO_2044 (O_2044,N_29896,N_29172);
or UO_2045 (O_2045,N_29063,N_29538);
nand UO_2046 (O_2046,N_29215,N_29820);
and UO_2047 (O_2047,N_29258,N_29318);
and UO_2048 (O_2048,N_29115,N_29555);
xor UO_2049 (O_2049,N_29034,N_29009);
nand UO_2050 (O_2050,N_29271,N_29989);
nor UO_2051 (O_2051,N_29249,N_29348);
nor UO_2052 (O_2052,N_29186,N_29500);
or UO_2053 (O_2053,N_29953,N_29896);
nand UO_2054 (O_2054,N_29477,N_29794);
and UO_2055 (O_2055,N_29690,N_29306);
or UO_2056 (O_2056,N_29520,N_29799);
or UO_2057 (O_2057,N_29177,N_29542);
nand UO_2058 (O_2058,N_29493,N_29837);
nand UO_2059 (O_2059,N_29475,N_29760);
xnor UO_2060 (O_2060,N_29080,N_29454);
nand UO_2061 (O_2061,N_29563,N_29716);
nand UO_2062 (O_2062,N_29095,N_29456);
and UO_2063 (O_2063,N_29121,N_29736);
or UO_2064 (O_2064,N_29488,N_29764);
xnor UO_2065 (O_2065,N_29530,N_29455);
or UO_2066 (O_2066,N_29191,N_29993);
nor UO_2067 (O_2067,N_29472,N_29508);
nand UO_2068 (O_2068,N_29390,N_29622);
nand UO_2069 (O_2069,N_29655,N_29596);
xnor UO_2070 (O_2070,N_29010,N_29801);
and UO_2071 (O_2071,N_29586,N_29017);
or UO_2072 (O_2072,N_29392,N_29932);
and UO_2073 (O_2073,N_29619,N_29894);
and UO_2074 (O_2074,N_29552,N_29966);
and UO_2075 (O_2075,N_29536,N_29579);
xnor UO_2076 (O_2076,N_29481,N_29767);
and UO_2077 (O_2077,N_29636,N_29321);
xor UO_2078 (O_2078,N_29573,N_29768);
or UO_2079 (O_2079,N_29363,N_29535);
nand UO_2080 (O_2080,N_29088,N_29494);
and UO_2081 (O_2081,N_29424,N_29604);
xnor UO_2082 (O_2082,N_29909,N_29902);
xor UO_2083 (O_2083,N_29690,N_29509);
or UO_2084 (O_2084,N_29344,N_29509);
xnor UO_2085 (O_2085,N_29587,N_29186);
nor UO_2086 (O_2086,N_29118,N_29043);
or UO_2087 (O_2087,N_29353,N_29920);
and UO_2088 (O_2088,N_29192,N_29673);
or UO_2089 (O_2089,N_29704,N_29219);
nand UO_2090 (O_2090,N_29779,N_29387);
or UO_2091 (O_2091,N_29007,N_29843);
and UO_2092 (O_2092,N_29885,N_29797);
or UO_2093 (O_2093,N_29339,N_29626);
and UO_2094 (O_2094,N_29141,N_29411);
or UO_2095 (O_2095,N_29315,N_29681);
or UO_2096 (O_2096,N_29888,N_29793);
xnor UO_2097 (O_2097,N_29447,N_29026);
or UO_2098 (O_2098,N_29758,N_29696);
or UO_2099 (O_2099,N_29535,N_29882);
and UO_2100 (O_2100,N_29008,N_29804);
nor UO_2101 (O_2101,N_29131,N_29483);
nor UO_2102 (O_2102,N_29500,N_29580);
xnor UO_2103 (O_2103,N_29943,N_29346);
or UO_2104 (O_2104,N_29341,N_29283);
nand UO_2105 (O_2105,N_29689,N_29377);
or UO_2106 (O_2106,N_29566,N_29502);
xnor UO_2107 (O_2107,N_29803,N_29986);
nand UO_2108 (O_2108,N_29059,N_29852);
xor UO_2109 (O_2109,N_29940,N_29618);
xnor UO_2110 (O_2110,N_29160,N_29548);
or UO_2111 (O_2111,N_29848,N_29235);
xor UO_2112 (O_2112,N_29849,N_29907);
nor UO_2113 (O_2113,N_29134,N_29047);
and UO_2114 (O_2114,N_29021,N_29192);
and UO_2115 (O_2115,N_29644,N_29385);
nor UO_2116 (O_2116,N_29360,N_29672);
xnor UO_2117 (O_2117,N_29832,N_29607);
and UO_2118 (O_2118,N_29806,N_29521);
xor UO_2119 (O_2119,N_29840,N_29303);
nor UO_2120 (O_2120,N_29283,N_29313);
xor UO_2121 (O_2121,N_29464,N_29765);
nor UO_2122 (O_2122,N_29645,N_29579);
and UO_2123 (O_2123,N_29884,N_29922);
and UO_2124 (O_2124,N_29260,N_29892);
and UO_2125 (O_2125,N_29556,N_29516);
or UO_2126 (O_2126,N_29419,N_29035);
xnor UO_2127 (O_2127,N_29269,N_29857);
nor UO_2128 (O_2128,N_29885,N_29692);
nor UO_2129 (O_2129,N_29915,N_29985);
and UO_2130 (O_2130,N_29593,N_29261);
nor UO_2131 (O_2131,N_29632,N_29044);
and UO_2132 (O_2132,N_29607,N_29413);
and UO_2133 (O_2133,N_29362,N_29999);
nand UO_2134 (O_2134,N_29468,N_29514);
nand UO_2135 (O_2135,N_29006,N_29029);
nand UO_2136 (O_2136,N_29070,N_29608);
or UO_2137 (O_2137,N_29055,N_29455);
and UO_2138 (O_2138,N_29415,N_29784);
and UO_2139 (O_2139,N_29034,N_29437);
xor UO_2140 (O_2140,N_29953,N_29929);
xor UO_2141 (O_2141,N_29538,N_29956);
nor UO_2142 (O_2142,N_29708,N_29142);
nor UO_2143 (O_2143,N_29972,N_29527);
xor UO_2144 (O_2144,N_29844,N_29675);
or UO_2145 (O_2145,N_29911,N_29021);
nand UO_2146 (O_2146,N_29668,N_29876);
and UO_2147 (O_2147,N_29358,N_29506);
and UO_2148 (O_2148,N_29703,N_29792);
nor UO_2149 (O_2149,N_29551,N_29813);
and UO_2150 (O_2150,N_29776,N_29522);
and UO_2151 (O_2151,N_29682,N_29033);
nor UO_2152 (O_2152,N_29515,N_29542);
nor UO_2153 (O_2153,N_29862,N_29795);
nand UO_2154 (O_2154,N_29835,N_29532);
xor UO_2155 (O_2155,N_29313,N_29237);
and UO_2156 (O_2156,N_29186,N_29607);
or UO_2157 (O_2157,N_29012,N_29366);
and UO_2158 (O_2158,N_29688,N_29073);
xnor UO_2159 (O_2159,N_29640,N_29727);
or UO_2160 (O_2160,N_29495,N_29099);
or UO_2161 (O_2161,N_29252,N_29899);
nand UO_2162 (O_2162,N_29429,N_29749);
or UO_2163 (O_2163,N_29495,N_29089);
or UO_2164 (O_2164,N_29486,N_29044);
or UO_2165 (O_2165,N_29899,N_29834);
and UO_2166 (O_2166,N_29213,N_29054);
nor UO_2167 (O_2167,N_29884,N_29131);
nor UO_2168 (O_2168,N_29355,N_29200);
and UO_2169 (O_2169,N_29070,N_29157);
and UO_2170 (O_2170,N_29269,N_29634);
or UO_2171 (O_2171,N_29699,N_29942);
xor UO_2172 (O_2172,N_29836,N_29178);
nor UO_2173 (O_2173,N_29158,N_29523);
nand UO_2174 (O_2174,N_29794,N_29439);
nand UO_2175 (O_2175,N_29183,N_29601);
and UO_2176 (O_2176,N_29568,N_29144);
and UO_2177 (O_2177,N_29946,N_29351);
and UO_2178 (O_2178,N_29912,N_29320);
nor UO_2179 (O_2179,N_29525,N_29355);
xnor UO_2180 (O_2180,N_29847,N_29383);
or UO_2181 (O_2181,N_29104,N_29866);
nand UO_2182 (O_2182,N_29933,N_29026);
and UO_2183 (O_2183,N_29087,N_29567);
nand UO_2184 (O_2184,N_29786,N_29580);
nor UO_2185 (O_2185,N_29170,N_29645);
nand UO_2186 (O_2186,N_29410,N_29821);
and UO_2187 (O_2187,N_29811,N_29181);
xor UO_2188 (O_2188,N_29836,N_29342);
nand UO_2189 (O_2189,N_29308,N_29775);
xor UO_2190 (O_2190,N_29512,N_29487);
or UO_2191 (O_2191,N_29322,N_29504);
and UO_2192 (O_2192,N_29912,N_29631);
or UO_2193 (O_2193,N_29312,N_29073);
and UO_2194 (O_2194,N_29846,N_29950);
xor UO_2195 (O_2195,N_29815,N_29850);
or UO_2196 (O_2196,N_29466,N_29048);
xnor UO_2197 (O_2197,N_29501,N_29643);
nand UO_2198 (O_2198,N_29881,N_29852);
or UO_2199 (O_2199,N_29797,N_29510);
nor UO_2200 (O_2200,N_29431,N_29131);
and UO_2201 (O_2201,N_29492,N_29717);
and UO_2202 (O_2202,N_29445,N_29758);
or UO_2203 (O_2203,N_29509,N_29694);
nor UO_2204 (O_2204,N_29287,N_29944);
xor UO_2205 (O_2205,N_29278,N_29745);
xnor UO_2206 (O_2206,N_29456,N_29171);
nor UO_2207 (O_2207,N_29617,N_29361);
and UO_2208 (O_2208,N_29240,N_29869);
and UO_2209 (O_2209,N_29402,N_29648);
xnor UO_2210 (O_2210,N_29362,N_29220);
and UO_2211 (O_2211,N_29177,N_29100);
nor UO_2212 (O_2212,N_29895,N_29447);
and UO_2213 (O_2213,N_29247,N_29964);
or UO_2214 (O_2214,N_29298,N_29012);
nand UO_2215 (O_2215,N_29887,N_29106);
nand UO_2216 (O_2216,N_29834,N_29516);
xor UO_2217 (O_2217,N_29999,N_29917);
and UO_2218 (O_2218,N_29331,N_29344);
and UO_2219 (O_2219,N_29294,N_29548);
nand UO_2220 (O_2220,N_29317,N_29034);
and UO_2221 (O_2221,N_29516,N_29306);
or UO_2222 (O_2222,N_29042,N_29568);
or UO_2223 (O_2223,N_29530,N_29686);
nand UO_2224 (O_2224,N_29871,N_29199);
or UO_2225 (O_2225,N_29943,N_29707);
nor UO_2226 (O_2226,N_29626,N_29795);
and UO_2227 (O_2227,N_29633,N_29954);
nor UO_2228 (O_2228,N_29753,N_29713);
and UO_2229 (O_2229,N_29844,N_29603);
nor UO_2230 (O_2230,N_29117,N_29241);
or UO_2231 (O_2231,N_29374,N_29461);
xor UO_2232 (O_2232,N_29568,N_29947);
and UO_2233 (O_2233,N_29532,N_29817);
nand UO_2234 (O_2234,N_29630,N_29337);
and UO_2235 (O_2235,N_29118,N_29930);
or UO_2236 (O_2236,N_29890,N_29665);
or UO_2237 (O_2237,N_29521,N_29681);
or UO_2238 (O_2238,N_29312,N_29177);
nand UO_2239 (O_2239,N_29657,N_29733);
nor UO_2240 (O_2240,N_29847,N_29077);
xor UO_2241 (O_2241,N_29163,N_29331);
or UO_2242 (O_2242,N_29796,N_29113);
nand UO_2243 (O_2243,N_29325,N_29143);
nand UO_2244 (O_2244,N_29967,N_29954);
nor UO_2245 (O_2245,N_29775,N_29496);
nand UO_2246 (O_2246,N_29285,N_29127);
or UO_2247 (O_2247,N_29395,N_29801);
nand UO_2248 (O_2248,N_29906,N_29326);
and UO_2249 (O_2249,N_29651,N_29861);
nand UO_2250 (O_2250,N_29031,N_29165);
nor UO_2251 (O_2251,N_29825,N_29159);
and UO_2252 (O_2252,N_29608,N_29524);
xor UO_2253 (O_2253,N_29535,N_29424);
nand UO_2254 (O_2254,N_29517,N_29174);
nand UO_2255 (O_2255,N_29653,N_29433);
or UO_2256 (O_2256,N_29084,N_29402);
and UO_2257 (O_2257,N_29231,N_29139);
and UO_2258 (O_2258,N_29228,N_29967);
nand UO_2259 (O_2259,N_29555,N_29950);
nor UO_2260 (O_2260,N_29563,N_29522);
nand UO_2261 (O_2261,N_29783,N_29624);
or UO_2262 (O_2262,N_29242,N_29444);
nor UO_2263 (O_2263,N_29270,N_29492);
nor UO_2264 (O_2264,N_29801,N_29116);
xor UO_2265 (O_2265,N_29181,N_29428);
nand UO_2266 (O_2266,N_29572,N_29829);
or UO_2267 (O_2267,N_29942,N_29005);
nand UO_2268 (O_2268,N_29344,N_29527);
or UO_2269 (O_2269,N_29238,N_29520);
and UO_2270 (O_2270,N_29553,N_29989);
and UO_2271 (O_2271,N_29985,N_29300);
or UO_2272 (O_2272,N_29115,N_29402);
nor UO_2273 (O_2273,N_29564,N_29505);
nand UO_2274 (O_2274,N_29055,N_29375);
and UO_2275 (O_2275,N_29020,N_29607);
nand UO_2276 (O_2276,N_29296,N_29336);
and UO_2277 (O_2277,N_29828,N_29027);
and UO_2278 (O_2278,N_29586,N_29865);
and UO_2279 (O_2279,N_29061,N_29258);
nor UO_2280 (O_2280,N_29324,N_29997);
and UO_2281 (O_2281,N_29663,N_29043);
or UO_2282 (O_2282,N_29511,N_29540);
nand UO_2283 (O_2283,N_29555,N_29830);
nor UO_2284 (O_2284,N_29100,N_29342);
and UO_2285 (O_2285,N_29116,N_29939);
or UO_2286 (O_2286,N_29788,N_29804);
and UO_2287 (O_2287,N_29428,N_29815);
nand UO_2288 (O_2288,N_29020,N_29952);
nand UO_2289 (O_2289,N_29903,N_29870);
and UO_2290 (O_2290,N_29540,N_29207);
or UO_2291 (O_2291,N_29243,N_29424);
or UO_2292 (O_2292,N_29218,N_29955);
nand UO_2293 (O_2293,N_29787,N_29434);
nand UO_2294 (O_2294,N_29650,N_29935);
and UO_2295 (O_2295,N_29996,N_29456);
or UO_2296 (O_2296,N_29705,N_29773);
xnor UO_2297 (O_2297,N_29441,N_29026);
and UO_2298 (O_2298,N_29939,N_29084);
or UO_2299 (O_2299,N_29980,N_29758);
xnor UO_2300 (O_2300,N_29924,N_29503);
and UO_2301 (O_2301,N_29645,N_29127);
xnor UO_2302 (O_2302,N_29331,N_29266);
nand UO_2303 (O_2303,N_29863,N_29500);
xor UO_2304 (O_2304,N_29994,N_29209);
nand UO_2305 (O_2305,N_29913,N_29993);
nor UO_2306 (O_2306,N_29860,N_29127);
nor UO_2307 (O_2307,N_29157,N_29912);
and UO_2308 (O_2308,N_29807,N_29701);
nand UO_2309 (O_2309,N_29325,N_29434);
nor UO_2310 (O_2310,N_29314,N_29056);
and UO_2311 (O_2311,N_29712,N_29635);
and UO_2312 (O_2312,N_29730,N_29415);
or UO_2313 (O_2313,N_29852,N_29320);
xnor UO_2314 (O_2314,N_29464,N_29345);
nand UO_2315 (O_2315,N_29412,N_29286);
or UO_2316 (O_2316,N_29286,N_29661);
and UO_2317 (O_2317,N_29274,N_29934);
nor UO_2318 (O_2318,N_29152,N_29146);
or UO_2319 (O_2319,N_29578,N_29360);
nand UO_2320 (O_2320,N_29700,N_29400);
and UO_2321 (O_2321,N_29674,N_29190);
nand UO_2322 (O_2322,N_29502,N_29203);
nor UO_2323 (O_2323,N_29881,N_29589);
or UO_2324 (O_2324,N_29115,N_29749);
xnor UO_2325 (O_2325,N_29118,N_29677);
and UO_2326 (O_2326,N_29172,N_29049);
xnor UO_2327 (O_2327,N_29523,N_29067);
and UO_2328 (O_2328,N_29672,N_29532);
nor UO_2329 (O_2329,N_29669,N_29333);
nand UO_2330 (O_2330,N_29536,N_29277);
xor UO_2331 (O_2331,N_29885,N_29402);
xor UO_2332 (O_2332,N_29522,N_29554);
and UO_2333 (O_2333,N_29060,N_29781);
nor UO_2334 (O_2334,N_29997,N_29886);
nand UO_2335 (O_2335,N_29634,N_29102);
nor UO_2336 (O_2336,N_29211,N_29906);
xnor UO_2337 (O_2337,N_29493,N_29911);
nor UO_2338 (O_2338,N_29929,N_29137);
nor UO_2339 (O_2339,N_29285,N_29876);
or UO_2340 (O_2340,N_29725,N_29117);
or UO_2341 (O_2341,N_29014,N_29366);
nor UO_2342 (O_2342,N_29109,N_29775);
nor UO_2343 (O_2343,N_29475,N_29077);
nor UO_2344 (O_2344,N_29603,N_29159);
nand UO_2345 (O_2345,N_29912,N_29557);
nand UO_2346 (O_2346,N_29708,N_29128);
nand UO_2347 (O_2347,N_29623,N_29016);
or UO_2348 (O_2348,N_29249,N_29018);
or UO_2349 (O_2349,N_29992,N_29809);
nand UO_2350 (O_2350,N_29168,N_29283);
nand UO_2351 (O_2351,N_29793,N_29599);
and UO_2352 (O_2352,N_29191,N_29294);
and UO_2353 (O_2353,N_29574,N_29450);
and UO_2354 (O_2354,N_29136,N_29185);
xor UO_2355 (O_2355,N_29338,N_29486);
xnor UO_2356 (O_2356,N_29354,N_29640);
nand UO_2357 (O_2357,N_29954,N_29111);
nor UO_2358 (O_2358,N_29470,N_29005);
nand UO_2359 (O_2359,N_29618,N_29718);
and UO_2360 (O_2360,N_29177,N_29440);
xnor UO_2361 (O_2361,N_29700,N_29862);
xnor UO_2362 (O_2362,N_29224,N_29692);
and UO_2363 (O_2363,N_29647,N_29773);
or UO_2364 (O_2364,N_29677,N_29928);
xnor UO_2365 (O_2365,N_29305,N_29558);
or UO_2366 (O_2366,N_29412,N_29568);
or UO_2367 (O_2367,N_29151,N_29650);
or UO_2368 (O_2368,N_29660,N_29083);
or UO_2369 (O_2369,N_29865,N_29513);
or UO_2370 (O_2370,N_29542,N_29257);
nor UO_2371 (O_2371,N_29423,N_29173);
and UO_2372 (O_2372,N_29358,N_29837);
xor UO_2373 (O_2373,N_29480,N_29735);
and UO_2374 (O_2374,N_29020,N_29526);
nor UO_2375 (O_2375,N_29802,N_29016);
nor UO_2376 (O_2376,N_29862,N_29683);
xor UO_2377 (O_2377,N_29952,N_29905);
or UO_2378 (O_2378,N_29174,N_29981);
nor UO_2379 (O_2379,N_29181,N_29848);
xnor UO_2380 (O_2380,N_29111,N_29223);
nor UO_2381 (O_2381,N_29116,N_29149);
or UO_2382 (O_2382,N_29370,N_29698);
or UO_2383 (O_2383,N_29444,N_29112);
and UO_2384 (O_2384,N_29595,N_29003);
and UO_2385 (O_2385,N_29598,N_29793);
nand UO_2386 (O_2386,N_29080,N_29278);
nor UO_2387 (O_2387,N_29651,N_29119);
nor UO_2388 (O_2388,N_29703,N_29898);
and UO_2389 (O_2389,N_29477,N_29419);
or UO_2390 (O_2390,N_29885,N_29621);
xnor UO_2391 (O_2391,N_29031,N_29396);
xnor UO_2392 (O_2392,N_29925,N_29974);
xnor UO_2393 (O_2393,N_29423,N_29410);
nand UO_2394 (O_2394,N_29588,N_29341);
xnor UO_2395 (O_2395,N_29779,N_29454);
nand UO_2396 (O_2396,N_29156,N_29045);
or UO_2397 (O_2397,N_29474,N_29408);
nor UO_2398 (O_2398,N_29210,N_29936);
xnor UO_2399 (O_2399,N_29155,N_29068);
nand UO_2400 (O_2400,N_29382,N_29616);
or UO_2401 (O_2401,N_29972,N_29163);
nand UO_2402 (O_2402,N_29255,N_29854);
and UO_2403 (O_2403,N_29183,N_29841);
or UO_2404 (O_2404,N_29248,N_29348);
or UO_2405 (O_2405,N_29341,N_29976);
nor UO_2406 (O_2406,N_29110,N_29637);
or UO_2407 (O_2407,N_29352,N_29288);
and UO_2408 (O_2408,N_29015,N_29571);
and UO_2409 (O_2409,N_29749,N_29008);
or UO_2410 (O_2410,N_29613,N_29758);
and UO_2411 (O_2411,N_29888,N_29107);
or UO_2412 (O_2412,N_29895,N_29786);
and UO_2413 (O_2413,N_29062,N_29484);
or UO_2414 (O_2414,N_29247,N_29182);
and UO_2415 (O_2415,N_29288,N_29604);
nor UO_2416 (O_2416,N_29609,N_29739);
nand UO_2417 (O_2417,N_29812,N_29124);
xor UO_2418 (O_2418,N_29670,N_29572);
xnor UO_2419 (O_2419,N_29808,N_29828);
nand UO_2420 (O_2420,N_29692,N_29328);
nand UO_2421 (O_2421,N_29390,N_29757);
and UO_2422 (O_2422,N_29141,N_29977);
and UO_2423 (O_2423,N_29237,N_29701);
and UO_2424 (O_2424,N_29693,N_29040);
xnor UO_2425 (O_2425,N_29679,N_29061);
xor UO_2426 (O_2426,N_29223,N_29267);
or UO_2427 (O_2427,N_29757,N_29063);
xor UO_2428 (O_2428,N_29509,N_29183);
nand UO_2429 (O_2429,N_29296,N_29273);
nor UO_2430 (O_2430,N_29741,N_29506);
xnor UO_2431 (O_2431,N_29337,N_29684);
nor UO_2432 (O_2432,N_29945,N_29672);
xor UO_2433 (O_2433,N_29028,N_29876);
nor UO_2434 (O_2434,N_29310,N_29239);
nand UO_2435 (O_2435,N_29934,N_29241);
xor UO_2436 (O_2436,N_29468,N_29793);
and UO_2437 (O_2437,N_29094,N_29259);
and UO_2438 (O_2438,N_29076,N_29485);
nor UO_2439 (O_2439,N_29575,N_29019);
and UO_2440 (O_2440,N_29385,N_29012);
or UO_2441 (O_2441,N_29618,N_29939);
or UO_2442 (O_2442,N_29290,N_29592);
xnor UO_2443 (O_2443,N_29793,N_29730);
xor UO_2444 (O_2444,N_29553,N_29350);
nor UO_2445 (O_2445,N_29745,N_29819);
nor UO_2446 (O_2446,N_29555,N_29624);
or UO_2447 (O_2447,N_29178,N_29089);
nor UO_2448 (O_2448,N_29606,N_29502);
nand UO_2449 (O_2449,N_29795,N_29838);
or UO_2450 (O_2450,N_29571,N_29734);
nand UO_2451 (O_2451,N_29893,N_29351);
or UO_2452 (O_2452,N_29414,N_29521);
and UO_2453 (O_2453,N_29615,N_29844);
nor UO_2454 (O_2454,N_29692,N_29394);
and UO_2455 (O_2455,N_29902,N_29321);
and UO_2456 (O_2456,N_29235,N_29769);
nor UO_2457 (O_2457,N_29140,N_29513);
nor UO_2458 (O_2458,N_29576,N_29519);
or UO_2459 (O_2459,N_29079,N_29178);
nand UO_2460 (O_2460,N_29596,N_29162);
xnor UO_2461 (O_2461,N_29309,N_29095);
xnor UO_2462 (O_2462,N_29415,N_29631);
nand UO_2463 (O_2463,N_29591,N_29633);
nand UO_2464 (O_2464,N_29237,N_29532);
nand UO_2465 (O_2465,N_29988,N_29014);
and UO_2466 (O_2466,N_29778,N_29732);
xor UO_2467 (O_2467,N_29644,N_29648);
xnor UO_2468 (O_2468,N_29107,N_29227);
nand UO_2469 (O_2469,N_29453,N_29914);
and UO_2470 (O_2470,N_29438,N_29004);
xnor UO_2471 (O_2471,N_29347,N_29436);
and UO_2472 (O_2472,N_29263,N_29578);
nand UO_2473 (O_2473,N_29902,N_29362);
nor UO_2474 (O_2474,N_29525,N_29223);
or UO_2475 (O_2475,N_29345,N_29882);
nand UO_2476 (O_2476,N_29168,N_29490);
xnor UO_2477 (O_2477,N_29506,N_29684);
xnor UO_2478 (O_2478,N_29419,N_29165);
xor UO_2479 (O_2479,N_29374,N_29035);
nor UO_2480 (O_2480,N_29001,N_29918);
nor UO_2481 (O_2481,N_29286,N_29459);
nor UO_2482 (O_2482,N_29238,N_29292);
xor UO_2483 (O_2483,N_29374,N_29101);
nor UO_2484 (O_2484,N_29201,N_29143);
or UO_2485 (O_2485,N_29176,N_29631);
xnor UO_2486 (O_2486,N_29150,N_29397);
nor UO_2487 (O_2487,N_29374,N_29721);
nand UO_2488 (O_2488,N_29365,N_29969);
and UO_2489 (O_2489,N_29121,N_29021);
or UO_2490 (O_2490,N_29243,N_29315);
and UO_2491 (O_2491,N_29509,N_29322);
and UO_2492 (O_2492,N_29768,N_29384);
xnor UO_2493 (O_2493,N_29535,N_29840);
xor UO_2494 (O_2494,N_29917,N_29515);
and UO_2495 (O_2495,N_29302,N_29765);
nor UO_2496 (O_2496,N_29671,N_29378);
and UO_2497 (O_2497,N_29100,N_29889);
and UO_2498 (O_2498,N_29114,N_29879);
nand UO_2499 (O_2499,N_29143,N_29127);
nor UO_2500 (O_2500,N_29292,N_29075);
or UO_2501 (O_2501,N_29060,N_29596);
or UO_2502 (O_2502,N_29195,N_29518);
nor UO_2503 (O_2503,N_29338,N_29168);
nand UO_2504 (O_2504,N_29797,N_29623);
nor UO_2505 (O_2505,N_29320,N_29378);
xnor UO_2506 (O_2506,N_29716,N_29316);
nor UO_2507 (O_2507,N_29209,N_29731);
xnor UO_2508 (O_2508,N_29192,N_29670);
nand UO_2509 (O_2509,N_29262,N_29495);
or UO_2510 (O_2510,N_29662,N_29912);
and UO_2511 (O_2511,N_29007,N_29163);
xnor UO_2512 (O_2512,N_29503,N_29495);
nor UO_2513 (O_2513,N_29724,N_29112);
nand UO_2514 (O_2514,N_29172,N_29620);
and UO_2515 (O_2515,N_29594,N_29394);
and UO_2516 (O_2516,N_29195,N_29704);
nor UO_2517 (O_2517,N_29874,N_29319);
xnor UO_2518 (O_2518,N_29239,N_29254);
or UO_2519 (O_2519,N_29543,N_29229);
and UO_2520 (O_2520,N_29110,N_29043);
and UO_2521 (O_2521,N_29186,N_29712);
and UO_2522 (O_2522,N_29033,N_29879);
xnor UO_2523 (O_2523,N_29525,N_29543);
nand UO_2524 (O_2524,N_29224,N_29241);
and UO_2525 (O_2525,N_29536,N_29405);
nand UO_2526 (O_2526,N_29561,N_29173);
nor UO_2527 (O_2527,N_29466,N_29431);
nor UO_2528 (O_2528,N_29768,N_29915);
or UO_2529 (O_2529,N_29699,N_29944);
xor UO_2530 (O_2530,N_29040,N_29867);
nor UO_2531 (O_2531,N_29513,N_29986);
and UO_2532 (O_2532,N_29857,N_29682);
and UO_2533 (O_2533,N_29009,N_29321);
xor UO_2534 (O_2534,N_29395,N_29341);
and UO_2535 (O_2535,N_29122,N_29295);
nand UO_2536 (O_2536,N_29898,N_29422);
and UO_2537 (O_2537,N_29649,N_29430);
xor UO_2538 (O_2538,N_29019,N_29760);
or UO_2539 (O_2539,N_29510,N_29058);
nor UO_2540 (O_2540,N_29981,N_29485);
nand UO_2541 (O_2541,N_29560,N_29421);
xor UO_2542 (O_2542,N_29309,N_29586);
nand UO_2543 (O_2543,N_29704,N_29238);
or UO_2544 (O_2544,N_29996,N_29114);
nor UO_2545 (O_2545,N_29915,N_29127);
or UO_2546 (O_2546,N_29281,N_29823);
nand UO_2547 (O_2547,N_29406,N_29414);
or UO_2548 (O_2548,N_29379,N_29132);
nor UO_2549 (O_2549,N_29058,N_29084);
or UO_2550 (O_2550,N_29864,N_29150);
or UO_2551 (O_2551,N_29640,N_29305);
xnor UO_2552 (O_2552,N_29877,N_29861);
nand UO_2553 (O_2553,N_29119,N_29433);
or UO_2554 (O_2554,N_29029,N_29724);
xnor UO_2555 (O_2555,N_29119,N_29989);
and UO_2556 (O_2556,N_29419,N_29761);
and UO_2557 (O_2557,N_29865,N_29006);
nor UO_2558 (O_2558,N_29512,N_29693);
xor UO_2559 (O_2559,N_29370,N_29753);
nor UO_2560 (O_2560,N_29191,N_29679);
or UO_2561 (O_2561,N_29228,N_29878);
xor UO_2562 (O_2562,N_29603,N_29939);
nor UO_2563 (O_2563,N_29315,N_29840);
xor UO_2564 (O_2564,N_29287,N_29851);
and UO_2565 (O_2565,N_29026,N_29898);
nor UO_2566 (O_2566,N_29632,N_29540);
nor UO_2567 (O_2567,N_29204,N_29680);
or UO_2568 (O_2568,N_29021,N_29614);
or UO_2569 (O_2569,N_29007,N_29918);
nor UO_2570 (O_2570,N_29433,N_29898);
xor UO_2571 (O_2571,N_29454,N_29267);
nand UO_2572 (O_2572,N_29571,N_29660);
nand UO_2573 (O_2573,N_29450,N_29149);
or UO_2574 (O_2574,N_29917,N_29535);
xnor UO_2575 (O_2575,N_29242,N_29348);
or UO_2576 (O_2576,N_29471,N_29679);
and UO_2577 (O_2577,N_29270,N_29726);
or UO_2578 (O_2578,N_29872,N_29781);
xnor UO_2579 (O_2579,N_29765,N_29330);
and UO_2580 (O_2580,N_29341,N_29802);
xnor UO_2581 (O_2581,N_29815,N_29511);
and UO_2582 (O_2582,N_29375,N_29189);
or UO_2583 (O_2583,N_29070,N_29483);
and UO_2584 (O_2584,N_29254,N_29515);
nor UO_2585 (O_2585,N_29591,N_29446);
nor UO_2586 (O_2586,N_29332,N_29791);
nand UO_2587 (O_2587,N_29850,N_29993);
nor UO_2588 (O_2588,N_29273,N_29708);
xor UO_2589 (O_2589,N_29758,N_29165);
nand UO_2590 (O_2590,N_29144,N_29601);
or UO_2591 (O_2591,N_29083,N_29962);
or UO_2592 (O_2592,N_29008,N_29866);
and UO_2593 (O_2593,N_29289,N_29942);
or UO_2594 (O_2594,N_29310,N_29577);
nand UO_2595 (O_2595,N_29292,N_29031);
or UO_2596 (O_2596,N_29420,N_29669);
and UO_2597 (O_2597,N_29595,N_29861);
nand UO_2598 (O_2598,N_29277,N_29220);
nand UO_2599 (O_2599,N_29324,N_29814);
and UO_2600 (O_2600,N_29601,N_29865);
nand UO_2601 (O_2601,N_29414,N_29480);
nor UO_2602 (O_2602,N_29759,N_29336);
xor UO_2603 (O_2603,N_29067,N_29272);
nor UO_2604 (O_2604,N_29087,N_29446);
xnor UO_2605 (O_2605,N_29038,N_29788);
nor UO_2606 (O_2606,N_29393,N_29273);
and UO_2607 (O_2607,N_29488,N_29066);
nand UO_2608 (O_2608,N_29277,N_29911);
xnor UO_2609 (O_2609,N_29525,N_29137);
nor UO_2610 (O_2610,N_29223,N_29343);
and UO_2611 (O_2611,N_29970,N_29439);
or UO_2612 (O_2612,N_29647,N_29182);
and UO_2613 (O_2613,N_29439,N_29959);
or UO_2614 (O_2614,N_29756,N_29604);
xor UO_2615 (O_2615,N_29343,N_29882);
nand UO_2616 (O_2616,N_29849,N_29080);
or UO_2617 (O_2617,N_29156,N_29845);
nor UO_2618 (O_2618,N_29948,N_29729);
nor UO_2619 (O_2619,N_29603,N_29385);
xor UO_2620 (O_2620,N_29668,N_29234);
nand UO_2621 (O_2621,N_29834,N_29547);
nand UO_2622 (O_2622,N_29698,N_29971);
or UO_2623 (O_2623,N_29829,N_29461);
or UO_2624 (O_2624,N_29700,N_29961);
nor UO_2625 (O_2625,N_29607,N_29353);
nor UO_2626 (O_2626,N_29814,N_29028);
xor UO_2627 (O_2627,N_29859,N_29744);
xor UO_2628 (O_2628,N_29697,N_29647);
nand UO_2629 (O_2629,N_29571,N_29168);
xor UO_2630 (O_2630,N_29685,N_29784);
xnor UO_2631 (O_2631,N_29729,N_29015);
nand UO_2632 (O_2632,N_29658,N_29398);
nand UO_2633 (O_2633,N_29033,N_29527);
xor UO_2634 (O_2634,N_29501,N_29124);
and UO_2635 (O_2635,N_29975,N_29692);
or UO_2636 (O_2636,N_29621,N_29995);
nand UO_2637 (O_2637,N_29052,N_29044);
xor UO_2638 (O_2638,N_29480,N_29052);
and UO_2639 (O_2639,N_29282,N_29076);
nor UO_2640 (O_2640,N_29564,N_29855);
xnor UO_2641 (O_2641,N_29902,N_29190);
nand UO_2642 (O_2642,N_29959,N_29363);
xnor UO_2643 (O_2643,N_29065,N_29651);
xor UO_2644 (O_2644,N_29594,N_29328);
or UO_2645 (O_2645,N_29104,N_29345);
xor UO_2646 (O_2646,N_29870,N_29755);
and UO_2647 (O_2647,N_29955,N_29264);
or UO_2648 (O_2648,N_29418,N_29970);
nor UO_2649 (O_2649,N_29108,N_29102);
nor UO_2650 (O_2650,N_29316,N_29644);
nor UO_2651 (O_2651,N_29109,N_29165);
nand UO_2652 (O_2652,N_29504,N_29715);
nor UO_2653 (O_2653,N_29294,N_29329);
nand UO_2654 (O_2654,N_29478,N_29334);
or UO_2655 (O_2655,N_29045,N_29137);
or UO_2656 (O_2656,N_29374,N_29431);
xor UO_2657 (O_2657,N_29806,N_29421);
xor UO_2658 (O_2658,N_29465,N_29211);
and UO_2659 (O_2659,N_29082,N_29239);
nor UO_2660 (O_2660,N_29993,N_29964);
or UO_2661 (O_2661,N_29188,N_29029);
and UO_2662 (O_2662,N_29768,N_29637);
or UO_2663 (O_2663,N_29699,N_29486);
xor UO_2664 (O_2664,N_29716,N_29547);
or UO_2665 (O_2665,N_29703,N_29321);
xor UO_2666 (O_2666,N_29285,N_29690);
nand UO_2667 (O_2667,N_29394,N_29836);
or UO_2668 (O_2668,N_29398,N_29617);
nand UO_2669 (O_2669,N_29839,N_29246);
xnor UO_2670 (O_2670,N_29361,N_29749);
and UO_2671 (O_2671,N_29203,N_29234);
and UO_2672 (O_2672,N_29952,N_29220);
nand UO_2673 (O_2673,N_29430,N_29541);
nor UO_2674 (O_2674,N_29834,N_29860);
nand UO_2675 (O_2675,N_29268,N_29900);
and UO_2676 (O_2676,N_29912,N_29053);
nand UO_2677 (O_2677,N_29472,N_29811);
xnor UO_2678 (O_2678,N_29366,N_29410);
xor UO_2679 (O_2679,N_29749,N_29626);
nor UO_2680 (O_2680,N_29624,N_29901);
xnor UO_2681 (O_2681,N_29601,N_29155);
nand UO_2682 (O_2682,N_29371,N_29306);
nand UO_2683 (O_2683,N_29070,N_29480);
or UO_2684 (O_2684,N_29151,N_29491);
xor UO_2685 (O_2685,N_29317,N_29558);
nor UO_2686 (O_2686,N_29128,N_29528);
and UO_2687 (O_2687,N_29305,N_29470);
and UO_2688 (O_2688,N_29897,N_29241);
nor UO_2689 (O_2689,N_29770,N_29243);
nor UO_2690 (O_2690,N_29858,N_29148);
or UO_2691 (O_2691,N_29369,N_29648);
nand UO_2692 (O_2692,N_29081,N_29350);
or UO_2693 (O_2693,N_29314,N_29803);
nand UO_2694 (O_2694,N_29592,N_29053);
and UO_2695 (O_2695,N_29724,N_29424);
xnor UO_2696 (O_2696,N_29588,N_29396);
nor UO_2697 (O_2697,N_29478,N_29689);
or UO_2698 (O_2698,N_29386,N_29067);
nand UO_2699 (O_2699,N_29158,N_29354);
or UO_2700 (O_2700,N_29144,N_29779);
or UO_2701 (O_2701,N_29184,N_29421);
nor UO_2702 (O_2702,N_29127,N_29191);
nand UO_2703 (O_2703,N_29760,N_29423);
and UO_2704 (O_2704,N_29120,N_29132);
nor UO_2705 (O_2705,N_29686,N_29972);
or UO_2706 (O_2706,N_29132,N_29704);
nor UO_2707 (O_2707,N_29898,N_29964);
xnor UO_2708 (O_2708,N_29273,N_29604);
xnor UO_2709 (O_2709,N_29011,N_29801);
and UO_2710 (O_2710,N_29645,N_29435);
and UO_2711 (O_2711,N_29007,N_29326);
nand UO_2712 (O_2712,N_29815,N_29502);
or UO_2713 (O_2713,N_29206,N_29764);
xor UO_2714 (O_2714,N_29916,N_29547);
nor UO_2715 (O_2715,N_29840,N_29943);
xor UO_2716 (O_2716,N_29814,N_29013);
and UO_2717 (O_2717,N_29773,N_29756);
nand UO_2718 (O_2718,N_29462,N_29345);
nand UO_2719 (O_2719,N_29570,N_29486);
xnor UO_2720 (O_2720,N_29242,N_29133);
and UO_2721 (O_2721,N_29655,N_29549);
nor UO_2722 (O_2722,N_29560,N_29750);
or UO_2723 (O_2723,N_29506,N_29920);
xnor UO_2724 (O_2724,N_29276,N_29633);
and UO_2725 (O_2725,N_29451,N_29181);
and UO_2726 (O_2726,N_29653,N_29225);
and UO_2727 (O_2727,N_29893,N_29397);
or UO_2728 (O_2728,N_29642,N_29167);
nand UO_2729 (O_2729,N_29761,N_29995);
or UO_2730 (O_2730,N_29891,N_29948);
xor UO_2731 (O_2731,N_29722,N_29020);
and UO_2732 (O_2732,N_29029,N_29419);
nor UO_2733 (O_2733,N_29305,N_29814);
nand UO_2734 (O_2734,N_29354,N_29914);
or UO_2735 (O_2735,N_29764,N_29256);
xor UO_2736 (O_2736,N_29967,N_29521);
or UO_2737 (O_2737,N_29554,N_29472);
or UO_2738 (O_2738,N_29704,N_29642);
nand UO_2739 (O_2739,N_29307,N_29808);
xor UO_2740 (O_2740,N_29605,N_29757);
nand UO_2741 (O_2741,N_29243,N_29951);
or UO_2742 (O_2742,N_29512,N_29283);
nor UO_2743 (O_2743,N_29438,N_29914);
xnor UO_2744 (O_2744,N_29790,N_29538);
nor UO_2745 (O_2745,N_29293,N_29099);
nand UO_2746 (O_2746,N_29876,N_29617);
and UO_2747 (O_2747,N_29406,N_29101);
nor UO_2748 (O_2748,N_29424,N_29460);
xnor UO_2749 (O_2749,N_29065,N_29172);
nand UO_2750 (O_2750,N_29175,N_29090);
and UO_2751 (O_2751,N_29300,N_29781);
xor UO_2752 (O_2752,N_29231,N_29400);
xor UO_2753 (O_2753,N_29442,N_29928);
or UO_2754 (O_2754,N_29838,N_29450);
or UO_2755 (O_2755,N_29866,N_29318);
nand UO_2756 (O_2756,N_29295,N_29836);
or UO_2757 (O_2757,N_29163,N_29403);
or UO_2758 (O_2758,N_29281,N_29249);
and UO_2759 (O_2759,N_29663,N_29038);
and UO_2760 (O_2760,N_29266,N_29085);
or UO_2761 (O_2761,N_29244,N_29511);
nor UO_2762 (O_2762,N_29094,N_29857);
nand UO_2763 (O_2763,N_29256,N_29363);
xor UO_2764 (O_2764,N_29590,N_29129);
and UO_2765 (O_2765,N_29806,N_29694);
nand UO_2766 (O_2766,N_29770,N_29936);
nor UO_2767 (O_2767,N_29943,N_29576);
nand UO_2768 (O_2768,N_29234,N_29393);
nor UO_2769 (O_2769,N_29768,N_29112);
or UO_2770 (O_2770,N_29980,N_29248);
xor UO_2771 (O_2771,N_29616,N_29990);
xor UO_2772 (O_2772,N_29685,N_29296);
xnor UO_2773 (O_2773,N_29360,N_29230);
xor UO_2774 (O_2774,N_29235,N_29518);
nor UO_2775 (O_2775,N_29492,N_29728);
or UO_2776 (O_2776,N_29730,N_29371);
nand UO_2777 (O_2777,N_29934,N_29685);
or UO_2778 (O_2778,N_29371,N_29427);
xor UO_2779 (O_2779,N_29591,N_29650);
nor UO_2780 (O_2780,N_29859,N_29985);
nor UO_2781 (O_2781,N_29613,N_29596);
nand UO_2782 (O_2782,N_29717,N_29823);
nor UO_2783 (O_2783,N_29676,N_29658);
and UO_2784 (O_2784,N_29080,N_29755);
or UO_2785 (O_2785,N_29687,N_29458);
nand UO_2786 (O_2786,N_29418,N_29103);
or UO_2787 (O_2787,N_29600,N_29429);
or UO_2788 (O_2788,N_29759,N_29172);
nor UO_2789 (O_2789,N_29288,N_29125);
nor UO_2790 (O_2790,N_29101,N_29126);
or UO_2791 (O_2791,N_29877,N_29482);
and UO_2792 (O_2792,N_29410,N_29456);
and UO_2793 (O_2793,N_29743,N_29777);
or UO_2794 (O_2794,N_29000,N_29969);
xor UO_2795 (O_2795,N_29290,N_29263);
nand UO_2796 (O_2796,N_29708,N_29282);
or UO_2797 (O_2797,N_29513,N_29218);
or UO_2798 (O_2798,N_29313,N_29732);
nor UO_2799 (O_2799,N_29203,N_29522);
nand UO_2800 (O_2800,N_29525,N_29279);
nor UO_2801 (O_2801,N_29098,N_29627);
or UO_2802 (O_2802,N_29217,N_29238);
nand UO_2803 (O_2803,N_29736,N_29160);
nand UO_2804 (O_2804,N_29405,N_29189);
nand UO_2805 (O_2805,N_29366,N_29586);
nor UO_2806 (O_2806,N_29828,N_29483);
or UO_2807 (O_2807,N_29600,N_29692);
nand UO_2808 (O_2808,N_29436,N_29015);
xor UO_2809 (O_2809,N_29518,N_29938);
or UO_2810 (O_2810,N_29900,N_29279);
nor UO_2811 (O_2811,N_29045,N_29532);
xnor UO_2812 (O_2812,N_29310,N_29569);
nand UO_2813 (O_2813,N_29045,N_29640);
xor UO_2814 (O_2814,N_29656,N_29949);
nor UO_2815 (O_2815,N_29924,N_29823);
xnor UO_2816 (O_2816,N_29753,N_29318);
xor UO_2817 (O_2817,N_29384,N_29929);
xnor UO_2818 (O_2818,N_29415,N_29956);
nor UO_2819 (O_2819,N_29396,N_29038);
nor UO_2820 (O_2820,N_29626,N_29011);
nor UO_2821 (O_2821,N_29787,N_29864);
xnor UO_2822 (O_2822,N_29108,N_29207);
or UO_2823 (O_2823,N_29668,N_29060);
and UO_2824 (O_2824,N_29039,N_29289);
and UO_2825 (O_2825,N_29810,N_29380);
nand UO_2826 (O_2826,N_29391,N_29115);
nor UO_2827 (O_2827,N_29348,N_29548);
or UO_2828 (O_2828,N_29518,N_29005);
xnor UO_2829 (O_2829,N_29497,N_29690);
nor UO_2830 (O_2830,N_29207,N_29647);
nand UO_2831 (O_2831,N_29945,N_29281);
xor UO_2832 (O_2832,N_29455,N_29991);
and UO_2833 (O_2833,N_29470,N_29833);
or UO_2834 (O_2834,N_29161,N_29657);
nor UO_2835 (O_2835,N_29467,N_29760);
or UO_2836 (O_2836,N_29044,N_29184);
or UO_2837 (O_2837,N_29189,N_29968);
xor UO_2838 (O_2838,N_29523,N_29180);
and UO_2839 (O_2839,N_29459,N_29040);
nand UO_2840 (O_2840,N_29027,N_29380);
or UO_2841 (O_2841,N_29256,N_29009);
xor UO_2842 (O_2842,N_29021,N_29501);
nand UO_2843 (O_2843,N_29019,N_29617);
xor UO_2844 (O_2844,N_29026,N_29328);
nor UO_2845 (O_2845,N_29177,N_29602);
xor UO_2846 (O_2846,N_29098,N_29175);
and UO_2847 (O_2847,N_29815,N_29578);
xor UO_2848 (O_2848,N_29066,N_29472);
xor UO_2849 (O_2849,N_29225,N_29456);
and UO_2850 (O_2850,N_29048,N_29948);
xnor UO_2851 (O_2851,N_29452,N_29219);
or UO_2852 (O_2852,N_29955,N_29927);
and UO_2853 (O_2853,N_29521,N_29575);
nand UO_2854 (O_2854,N_29798,N_29143);
nor UO_2855 (O_2855,N_29554,N_29456);
xnor UO_2856 (O_2856,N_29127,N_29356);
nor UO_2857 (O_2857,N_29812,N_29709);
or UO_2858 (O_2858,N_29917,N_29208);
or UO_2859 (O_2859,N_29712,N_29288);
or UO_2860 (O_2860,N_29326,N_29591);
or UO_2861 (O_2861,N_29959,N_29294);
nor UO_2862 (O_2862,N_29629,N_29359);
or UO_2863 (O_2863,N_29697,N_29203);
or UO_2864 (O_2864,N_29509,N_29641);
nand UO_2865 (O_2865,N_29626,N_29404);
nand UO_2866 (O_2866,N_29618,N_29575);
and UO_2867 (O_2867,N_29513,N_29216);
and UO_2868 (O_2868,N_29761,N_29433);
nand UO_2869 (O_2869,N_29679,N_29133);
nand UO_2870 (O_2870,N_29142,N_29566);
xnor UO_2871 (O_2871,N_29765,N_29017);
xor UO_2872 (O_2872,N_29316,N_29581);
nand UO_2873 (O_2873,N_29317,N_29549);
nor UO_2874 (O_2874,N_29807,N_29972);
or UO_2875 (O_2875,N_29115,N_29632);
and UO_2876 (O_2876,N_29221,N_29723);
xnor UO_2877 (O_2877,N_29363,N_29762);
and UO_2878 (O_2878,N_29032,N_29061);
or UO_2879 (O_2879,N_29614,N_29947);
nor UO_2880 (O_2880,N_29635,N_29805);
nand UO_2881 (O_2881,N_29261,N_29734);
nor UO_2882 (O_2882,N_29825,N_29794);
nor UO_2883 (O_2883,N_29878,N_29139);
or UO_2884 (O_2884,N_29901,N_29320);
nand UO_2885 (O_2885,N_29688,N_29269);
xnor UO_2886 (O_2886,N_29361,N_29029);
xor UO_2887 (O_2887,N_29810,N_29641);
xor UO_2888 (O_2888,N_29183,N_29553);
or UO_2889 (O_2889,N_29382,N_29476);
xor UO_2890 (O_2890,N_29263,N_29171);
or UO_2891 (O_2891,N_29615,N_29504);
and UO_2892 (O_2892,N_29483,N_29054);
and UO_2893 (O_2893,N_29392,N_29992);
or UO_2894 (O_2894,N_29207,N_29918);
and UO_2895 (O_2895,N_29774,N_29362);
or UO_2896 (O_2896,N_29428,N_29751);
and UO_2897 (O_2897,N_29398,N_29115);
nor UO_2898 (O_2898,N_29489,N_29343);
or UO_2899 (O_2899,N_29092,N_29062);
or UO_2900 (O_2900,N_29970,N_29236);
or UO_2901 (O_2901,N_29653,N_29798);
or UO_2902 (O_2902,N_29202,N_29496);
xor UO_2903 (O_2903,N_29093,N_29749);
nor UO_2904 (O_2904,N_29163,N_29648);
and UO_2905 (O_2905,N_29989,N_29842);
nor UO_2906 (O_2906,N_29263,N_29259);
nor UO_2907 (O_2907,N_29877,N_29448);
and UO_2908 (O_2908,N_29070,N_29164);
and UO_2909 (O_2909,N_29119,N_29053);
and UO_2910 (O_2910,N_29324,N_29182);
or UO_2911 (O_2911,N_29688,N_29896);
or UO_2912 (O_2912,N_29606,N_29270);
nand UO_2913 (O_2913,N_29064,N_29114);
or UO_2914 (O_2914,N_29008,N_29086);
nor UO_2915 (O_2915,N_29605,N_29459);
and UO_2916 (O_2916,N_29039,N_29044);
and UO_2917 (O_2917,N_29327,N_29566);
nand UO_2918 (O_2918,N_29836,N_29505);
nand UO_2919 (O_2919,N_29560,N_29057);
nand UO_2920 (O_2920,N_29325,N_29067);
and UO_2921 (O_2921,N_29985,N_29118);
xnor UO_2922 (O_2922,N_29578,N_29364);
and UO_2923 (O_2923,N_29706,N_29716);
and UO_2924 (O_2924,N_29859,N_29764);
nor UO_2925 (O_2925,N_29670,N_29793);
xnor UO_2926 (O_2926,N_29560,N_29229);
and UO_2927 (O_2927,N_29273,N_29217);
xnor UO_2928 (O_2928,N_29795,N_29376);
nor UO_2929 (O_2929,N_29990,N_29424);
nand UO_2930 (O_2930,N_29987,N_29384);
or UO_2931 (O_2931,N_29202,N_29966);
nor UO_2932 (O_2932,N_29486,N_29376);
xnor UO_2933 (O_2933,N_29636,N_29287);
nand UO_2934 (O_2934,N_29829,N_29265);
and UO_2935 (O_2935,N_29847,N_29361);
and UO_2936 (O_2936,N_29869,N_29862);
xor UO_2937 (O_2937,N_29635,N_29420);
xor UO_2938 (O_2938,N_29296,N_29408);
xor UO_2939 (O_2939,N_29622,N_29579);
and UO_2940 (O_2940,N_29234,N_29402);
nor UO_2941 (O_2941,N_29201,N_29280);
or UO_2942 (O_2942,N_29709,N_29181);
and UO_2943 (O_2943,N_29978,N_29996);
or UO_2944 (O_2944,N_29571,N_29561);
nand UO_2945 (O_2945,N_29843,N_29885);
and UO_2946 (O_2946,N_29495,N_29135);
xnor UO_2947 (O_2947,N_29919,N_29785);
or UO_2948 (O_2948,N_29927,N_29075);
xnor UO_2949 (O_2949,N_29181,N_29289);
nor UO_2950 (O_2950,N_29625,N_29510);
nor UO_2951 (O_2951,N_29223,N_29445);
nand UO_2952 (O_2952,N_29179,N_29070);
xor UO_2953 (O_2953,N_29202,N_29533);
xnor UO_2954 (O_2954,N_29775,N_29209);
or UO_2955 (O_2955,N_29431,N_29990);
and UO_2956 (O_2956,N_29804,N_29736);
nand UO_2957 (O_2957,N_29978,N_29523);
nor UO_2958 (O_2958,N_29223,N_29246);
or UO_2959 (O_2959,N_29137,N_29827);
nor UO_2960 (O_2960,N_29141,N_29819);
and UO_2961 (O_2961,N_29110,N_29169);
nand UO_2962 (O_2962,N_29150,N_29110);
or UO_2963 (O_2963,N_29230,N_29214);
nand UO_2964 (O_2964,N_29369,N_29246);
and UO_2965 (O_2965,N_29240,N_29303);
nor UO_2966 (O_2966,N_29482,N_29848);
xor UO_2967 (O_2967,N_29791,N_29202);
nor UO_2968 (O_2968,N_29968,N_29481);
xnor UO_2969 (O_2969,N_29492,N_29151);
nand UO_2970 (O_2970,N_29904,N_29805);
xor UO_2971 (O_2971,N_29748,N_29502);
xor UO_2972 (O_2972,N_29002,N_29401);
or UO_2973 (O_2973,N_29698,N_29994);
xor UO_2974 (O_2974,N_29712,N_29630);
or UO_2975 (O_2975,N_29784,N_29515);
nand UO_2976 (O_2976,N_29418,N_29302);
xor UO_2977 (O_2977,N_29256,N_29691);
nor UO_2978 (O_2978,N_29907,N_29109);
or UO_2979 (O_2979,N_29406,N_29113);
nor UO_2980 (O_2980,N_29105,N_29934);
nor UO_2981 (O_2981,N_29582,N_29564);
and UO_2982 (O_2982,N_29265,N_29708);
xnor UO_2983 (O_2983,N_29723,N_29712);
and UO_2984 (O_2984,N_29195,N_29163);
and UO_2985 (O_2985,N_29616,N_29595);
nand UO_2986 (O_2986,N_29927,N_29155);
and UO_2987 (O_2987,N_29777,N_29303);
nand UO_2988 (O_2988,N_29803,N_29217);
and UO_2989 (O_2989,N_29515,N_29439);
xor UO_2990 (O_2990,N_29201,N_29395);
nand UO_2991 (O_2991,N_29172,N_29130);
nor UO_2992 (O_2992,N_29175,N_29925);
xor UO_2993 (O_2993,N_29898,N_29503);
nand UO_2994 (O_2994,N_29323,N_29938);
or UO_2995 (O_2995,N_29311,N_29760);
and UO_2996 (O_2996,N_29990,N_29055);
xnor UO_2997 (O_2997,N_29683,N_29941);
or UO_2998 (O_2998,N_29080,N_29668);
and UO_2999 (O_2999,N_29982,N_29799);
nand UO_3000 (O_3000,N_29579,N_29626);
xnor UO_3001 (O_3001,N_29198,N_29981);
xnor UO_3002 (O_3002,N_29812,N_29601);
and UO_3003 (O_3003,N_29399,N_29245);
and UO_3004 (O_3004,N_29687,N_29276);
or UO_3005 (O_3005,N_29816,N_29724);
nor UO_3006 (O_3006,N_29533,N_29190);
and UO_3007 (O_3007,N_29436,N_29256);
nor UO_3008 (O_3008,N_29501,N_29112);
and UO_3009 (O_3009,N_29347,N_29520);
nor UO_3010 (O_3010,N_29533,N_29659);
nor UO_3011 (O_3011,N_29196,N_29314);
nor UO_3012 (O_3012,N_29430,N_29708);
nand UO_3013 (O_3013,N_29861,N_29832);
xor UO_3014 (O_3014,N_29305,N_29288);
and UO_3015 (O_3015,N_29931,N_29160);
and UO_3016 (O_3016,N_29346,N_29149);
and UO_3017 (O_3017,N_29158,N_29979);
or UO_3018 (O_3018,N_29527,N_29387);
nand UO_3019 (O_3019,N_29439,N_29841);
nor UO_3020 (O_3020,N_29369,N_29211);
or UO_3021 (O_3021,N_29120,N_29465);
xor UO_3022 (O_3022,N_29097,N_29471);
nand UO_3023 (O_3023,N_29601,N_29090);
nand UO_3024 (O_3024,N_29792,N_29718);
and UO_3025 (O_3025,N_29571,N_29127);
and UO_3026 (O_3026,N_29391,N_29137);
nand UO_3027 (O_3027,N_29659,N_29681);
nand UO_3028 (O_3028,N_29682,N_29054);
or UO_3029 (O_3029,N_29822,N_29293);
nor UO_3030 (O_3030,N_29951,N_29177);
and UO_3031 (O_3031,N_29571,N_29174);
and UO_3032 (O_3032,N_29744,N_29866);
or UO_3033 (O_3033,N_29756,N_29907);
nand UO_3034 (O_3034,N_29251,N_29274);
nor UO_3035 (O_3035,N_29967,N_29870);
and UO_3036 (O_3036,N_29392,N_29455);
nand UO_3037 (O_3037,N_29791,N_29874);
and UO_3038 (O_3038,N_29238,N_29634);
nand UO_3039 (O_3039,N_29131,N_29588);
or UO_3040 (O_3040,N_29490,N_29796);
nand UO_3041 (O_3041,N_29265,N_29465);
or UO_3042 (O_3042,N_29455,N_29107);
nor UO_3043 (O_3043,N_29335,N_29985);
xnor UO_3044 (O_3044,N_29822,N_29991);
nor UO_3045 (O_3045,N_29600,N_29135);
nor UO_3046 (O_3046,N_29393,N_29431);
or UO_3047 (O_3047,N_29688,N_29568);
nand UO_3048 (O_3048,N_29557,N_29627);
xnor UO_3049 (O_3049,N_29724,N_29019);
or UO_3050 (O_3050,N_29070,N_29573);
and UO_3051 (O_3051,N_29735,N_29904);
or UO_3052 (O_3052,N_29997,N_29700);
and UO_3053 (O_3053,N_29619,N_29427);
xor UO_3054 (O_3054,N_29945,N_29242);
or UO_3055 (O_3055,N_29588,N_29392);
nor UO_3056 (O_3056,N_29549,N_29535);
xnor UO_3057 (O_3057,N_29203,N_29517);
or UO_3058 (O_3058,N_29418,N_29893);
xor UO_3059 (O_3059,N_29423,N_29204);
nor UO_3060 (O_3060,N_29834,N_29878);
nand UO_3061 (O_3061,N_29282,N_29624);
and UO_3062 (O_3062,N_29476,N_29667);
nand UO_3063 (O_3063,N_29164,N_29877);
xnor UO_3064 (O_3064,N_29243,N_29793);
or UO_3065 (O_3065,N_29796,N_29623);
xor UO_3066 (O_3066,N_29840,N_29230);
and UO_3067 (O_3067,N_29659,N_29229);
xnor UO_3068 (O_3068,N_29657,N_29283);
or UO_3069 (O_3069,N_29565,N_29422);
nand UO_3070 (O_3070,N_29810,N_29774);
nand UO_3071 (O_3071,N_29230,N_29674);
nand UO_3072 (O_3072,N_29166,N_29885);
and UO_3073 (O_3073,N_29964,N_29498);
xnor UO_3074 (O_3074,N_29362,N_29982);
and UO_3075 (O_3075,N_29091,N_29587);
xor UO_3076 (O_3076,N_29640,N_29397);
and UO_3077 (O_3077,N_29473,N_29591);
nor UO_3078 (O_3078,N_29926,N_29696);
nor UO_3079 (O_3079,N_29928,N_29234);
xnor UO_3080 (O_3080,N_29819,N_29770);
nand UO_3081 (O_3081,N_29785,N_29348);
and UO_3082 (O_3082,N_29263,N_29571);
nand UO_3083 (O_3083,N_29219,N_29924);
nor UO_3084 (O_3084,N_29866,N_29439);
nand UO_3085 (O_3085,N_29800,N_29094);
and UO_3086 (O_3086,N_29373,N_29235);
or UO_3087 (O_3087,N_29150,N_29858);
xnor UO_3088 (O_3088,N_29482,N_29007);
nand UO_3089 (O_3089,N_29112,N_29407);
nand UO_3090 (O_3090,N_29949,N_29012);
and UO_3091 (O_3091,N_29885,N_29565);
and UO_3092 (O_3092,N_29669,N_29107);
xnor UO_3093 (O_3093,N_29192,N_29272);
and UO_3094 (O_3094,N_29752,N_29310);
or UO_3095 (O_3095,N_29446,N_29723);
nand UO_3096 (O_3096,N_29029,N_29487);
nor UO_3097 (O_3097,N_29059,N_29398);
and UO_3098 (O_3098,N_29677,N_29151);
and UO_3099 (O_3099,N_29775,N_29637);
or UO_3100 (O_3100,N_29947,N_29814);
and UO_3101 (O_3101,N_29976,N_29413);
xor UO_3102 (O_3102,N_29538,N_29732);
xor UO_3103 (O_3103,N_29029,N_29200);
or UO_3104 (O_3104,N_29128,N_29335);
xnor UO_3105 (O_3105,N_29073,N_29217);
nor UO_3106 (O_3106,N_29438,N_29394);
nor UO_3107 (O_3107,N_29035,N_29558);
or UO_3108 (O_3108,N_29113,N_29111);
and UO_3109 (O_3109,N_29805,N_29397);
or UO_3110 (O_3110,N_29516,N_29731);
xnor UO_3111 (O_3111,N_29447,N_29190);
xnor UO_3112 (O_3112,N_29535,N_29942);
and UO_3113 (O_3113,N_29321,N_29164);
nand UO_3114 (O_3114,N_29364,N_29511);
xor UO_3115 (O_3115,N_29437,N_29122);
xor UO_3116 (O_3116,N_29010,N_29874);
or UO_3117 (O_3117,N_29906,N_29320);
and UO_3118 (O_3118,N_29052,N_29091);
and UO_3119 (O_3119,N_29268,N_29949);
xor UO_3120 (O_3120,N_29165,N_29744);
and UO_3121 (O_3121,N_29276,N_29130);
and UO_3122 (O_3122,N_29644,N_29322);
nor UO_3123 (O_3123,N_29175,N_29662);
nor UO_3124 (O_3124,N_29070,N_29469);
or UO_3125 (O_3125,N_29778,N_29482);
xor UO_3126 (O_3126,N_29744,N_29485);
and UO_3127 (O_3127,N_29800,N_29592);
or UO_3128 (O_3128,N_29950,N_29348);
nand UO_3129 (O_3129,N_29300,N_29519);
and UO_3130 (O_3130,N_29577,N_29642);
xor UO_3131 (O_3131,N_29781,N_29519);
or UO_3132 (O_3132,N_29271,N_29113);
nor UO_3133 (O_3133,N_29708,N_29657);
xnor UO_3134 (O_3134,N_29009,N_29417);
xnor UO_3135 (O_3135,N_29796,N_29922);
xor UO_3136 (O_3136,N_29060,N_29928);
or UO_3137 (O_3137,N_29309,N_29767);
xor UO_3138 (O_3138,N_29979,N_29242);
nor UO_3139 (O_3139,N_29684,N_29609);
xor UO_3140 (O_3140,N_29407,N_29539);
nor UO_3141 (O_3141,N_29608,N_29232);
nor UO_3142 (O_3142,N_29540,N_29482);
nor UO_3143 (O_3143,N_29908,N_29307);
and UO_3144 (O_3144,N_29626,N_29532);
nor UO_3145 (O_3145,N_29834,N_29840);
and UO_3146 (O_3146,N_29871,N_29630);
and UO_3147 (O_3147,N_29478,N_29953);
nor UO_3148 (O_3148,N_29807,N_29527);
xor UO_3149 (O_3149,N_29295,N_29643);
nor UO_3150 (O_3150,N_29077,N_29215);
or UO_3151 (O_3151,N_29873,N_29867);
and UO_3152 (O_3152,N_29299,N_29712);
or UO_3153 (O_3153,N_29125,N_29062);
and UO_3154 (O_3154,N_29818,N_29420);
or UO_3155 (O_3155,N_29672,N_29955);
xnor UO_3156 (O_3156,N_29041,N_29644);
xnor UO_3157 (O_3157,N_29112,N_29520);
or UO_3158 (O_3158,N_29000,N_29135);
nand UO_3159 (O_3159,N_29541,N_29336);
nand UO_3160 (O_3160,N_29989,N_29390);
or UO_3161 (O_3161,N_29839,N_29889);
or UO_3162 (O_3162,N_29751,N_29369);
nor UO_3163 (O_3163,N_29007,N_29615);
nand UO_3164 (O_3164,N_29969,N_29035);
nor UO_3165 (O_3165,N_29736,N_29139);
or UO_3166 (O_3166,N_29794,N_29045);
nor UO_3167 (O_3167,N_29821,N_29088);
xor UO_3168 (O_3168,N_29115,N_29564);
nor UO_3169 (O_3169,N_29230,N_29385);
nand UO_3170 (O_3170,N_29175,N_29083);
nor UO_3171 (O_3171,N_29156,N_29004);
and UO_3172 (O_3172,N_29375,N_29058);
xnor UO_3173 (O_3173,N_29596,N_29195);
or UO_3174 (O_3174,N_29164,N_29404);
xnor UO_3175 (O_3175,N_29443,N_29292);
nand UO_3176 (O_3176,N_29898,N_29841);
nand UO_3177 (O_3177,N_29833,N_29793);
and UO_3178 (O_3178,N_29579,N_29589);
or UO_3179 (O_3179,N_29643,N_29599);
nand UO_3180 (O_3180,N_29895,N_29703);
nand UO_3181 (O_3181,N_29114,N_29211);
xor UO_3182 (O_3182,N_29744,N_29488);
xor UO_3183 (O_3183,N_29807,N_29452);
nand UO_3184 (O_3184,N_29329,N_29706);
nor UO_3185 (O_3185,N_29400,N_29332);
nor UO_3186 (O_3186,N_29090,N_29121);
or UO_3187 (O_3187,N_29571,N_29104);
xnor UO_3188 (O_3188,N_29119,N_29715);
nand UO_3189 (O_3189,N_29121,N_29888);
xnor UO_3190 (O_3190,N_29019,N_29343);
xor UO_3191 (O_3191,N_29100,N_29211);
xor UO_3192 (O_3192,N_29657,N_29951);
or UO_3193 (O_3193,N_29837,N_29121);
xnor UO_3194 (O_3194,N_29929,N_29883);
and UO_3195 (O_3195,N_29008,N_29109);
nor UO_3196 (O_3196,N_29401,N_29596);
and UO_3197 (O_3197,N_29709,N_29483);
and UO_3198 (O_3198,N_29115,N_29941);
and UO_3199 (O_3199,N_29846,N_29015);
xor UO_3200 (O_3200,N_29637,N_29293);
or UO_3201 (O_3201,N_29108,N_29359);
and UO_3202 (O_3202,N_29611,N_29498);
nor UO_3203 (O_3203,N_29782,N_29944);
nor UO_3204 (O_3204,N_29630,N_29150);
or UO_3205 (O_3205,N_29429,N_29731);
nand UO_3206 (O_3206,N_29194,N_29443);
nand UO_3207 (O_3207,N_29500,N_29334);
or UO_3208 (O_3208,N_29051,N_29475);
and UO_3209 (O_3209,N_29817,N_29259);
and UO_3210 (O_3210,N_29177,N_29126);
and UO_3211 (O_3211,N_29205,N_29165);
and UO_3212 (O_3212,N_29943,N_29785);
and UO_3213 (O_3213,N_29371,N_29818);
xnor UO_3214 (O_3214,N_29841,N_29776);
xnor UO_3215 (O_3215,N_29736,N_29869);
nor UO_3216 (O_3216,N_29028,N_29182);
nand UO_3217 (O_3217,N_29031,N_29515);
xor UO_3218 (O_3218,N_29373,N_29919);
xnor UO_3219 (O_3219,N_29329,N_29178);
nor UO_3220 (O_3220,N_29256,N_29578);
nand UO_3221 (O_3221,N_29424,N_29190);
nand UO_3222 (O_3222,N_29365,N_29051);
nand UO_3223 (O_3223,N_29936,N_29322);
xor UO_3224 (O_3224,N_29746,N_29437);
and UO_3225 (O_3225,N_29093,N_29560);
or UO_3226 (O_3226,N_29278,N_29073);
nand UO_3227 (O_3227,N_29619,N_29807);
nor UO_3228 (O_3228,N_29293,N_29619);
and UO_3229 (O_3229,N_29279,N_29897);
xor UO_3230 (O_3230,N_29439,N_29811);
or UO_3231 (O_3231,N_29326,N_29399);
or UO_3232 (O_3232,N_29823,N_29290);
nand UO_3233 (O_3233,N_29750,N_29996);
nand UO_3234 (O_3234,N_29390,N_29089);
nor UO_3235 (O_3235,N_29866,N_29366);
nand UO_3236 (O_3236,N_29062,N_29311);
and UO_3237 (O_3237,N_29998,N_29015);
nand UO_3238 (O_3238,N_29276,N_29568);
xnor UO_3239 (O_3239,N_29350,N_29152);
xor UO_3240 (O_3240,N_29949,N_29620);
nor UO_3241 (O_3241,N_29275,N_29110);
or UO_3242 (O_3242,N_29387,N_29777);
or UO_3243 (O_3243,N_29850,N_29598);
xor UO_3244 (O_3244,N_29837,N_29635);
xor UO_3245 (O_3245,N_29253,N_29550);
and UO_3246 (O_3246,N_29149,N_29430);
or UO_3247 (O_3247,N_29252,N_29869);
nor UO_3248 (O_3248,N_29675,N_29704);
and UO_3249 (O_3249,N_29353,N_29170);
nand UO_3250 (O_3250,N_29872,N_29786);
and UO_3251 (O_3251,N_29639,N_29548);
or UO_3252 (O_3252,N_29439,N_29932);
xnor UO_3253 (O_3253,N_29744,N_29951);
nor UO_3254 (O_3254,N_29024,N_29116);
nor UO_3255 (O_3255,N_29457,N_29258);
or UO_3256 (O_3256,N_29604,N_29316);
nand UO_3257 (O_3257,N_29320,N_29798);
nand UO_3258 (O_3258,N_29502,N_29788);
or UO_3259 (O_3259,N_29164,N_29844);
and UO_3260 (O_3260,N_29647,N_29993);
nand UO_3261 (O_3261,N_29045,N_29733);
xnor UO_3262 (O_3262,N_29602,N_29099);
or UO_3263 (O_3263,N_29506,N_29575);
xor UO_3264 (O_3264,N_29464,N_29248);
xnor UO_3265 (O_3265,N_29603,N_29879);
and UO_3266 (O_3266,N_29786,N_29644);
nand UO_3267 (O_3267,N_29018,N_29844);
or UO_3268 (O_3268,N_29948,N_29541);
nand UO_3269 (O_3269,N_29224,N_29397);
nand UO_3270 (O_3270,N_29362,N_29727);
or UO_3271 (O_3271,N_29859,N_29203);
xnor UO_3272 (O_3272,N_29210,N_29571);
and UO_3273 (O_3273,N_29965,N_29833);
or UO_3274 (O_3274,N_29030,N_29314);
or UO_3275 (O_3275,N_29081,N_29461);
nor UO_3276 (O_3276,N_29790,N_29959);
and UO_3277 (O_3277,N_29181,N_29310);
xor UO_3278 (O_3278,N_29103,N_29889);
or UO_3279 (O_3279,N_29252,N_29256);
nand UO_3280 (O_3280,N_29200,N_29096);
and UO_3281 (O_3281,N_29075,N_29514);
and UO_3282 (O_3282,N_29400,N_29356);
xor UO_3283 (O_3283,N_29776,N_29955);
xor UO_3284 (O_3284,N_29137,N_29084);
xnor UO_3285 (O_3285,N_29610,N_29968);
nor UO_3286 (O_3286,N_29786,N_29024);
nor UO_3287 (O_3287,N_29269,N_29496);
and UO_3288 (O_3288,N_29088,N_29084);
and UO_3289 (O_3289,N_29183,N_29674);
or UO_3290 (O_3290,N_29050,N_29133);
nand UO_3291 (O_3291,N_29709,N_29599);
or UO_3292 (O_3292,N_29069,N_29230);
or UO_3293 (O_3293,N_29535,N_29711);
and UO_3294 (O_3294,N_29347,N_29839);
or UO_3295 (O_3295,N_29494,N_29391);
xnor UO_3296 (O_3296,N_29849,N_29231);
nor UO_3297 (O_3297,N_29748,N_29103);
and UO_3298 (O_3298,N_29988,N_29073);
nor UO_3299 (O_3299,N_29359,N_29104);
and UO_3300 (O_3300,N_29951,N_29895);
xnor UO_3301 (O_3301,N_29968,N_29707);
and UO_3302 (O_3302,N_29102,N_29359);
nand UO_3303 (O_3303,N_29169,N_29393);
nor UO_3304 (O_3304,N_29831,N_29242);
xor UO_3305 (O_3305,N_29217,N_29424);
xor UO_3306 (O_3306,N_29343,N_29946);
or UO_3307 (O_3307,N_29851,N_29234);
nor UO_3308 (O_3308,N_29561,N_29514);
or UO_3309 (O_3309,N_29157,N_29155);
nor UO_3310 (O_3310,N_29938,N_29133);
xnor UO_3311 (O_3311,N_29270,N_29552);
nand UO_3312 (O_3312,N_29300,N_29416);
and UO_3313 (O_3313,N_29521,N_29988);
xor UO_3314 (O_3314,N_29019,N_29064);
nand UO_3315 (O_3315,N_29389,N_29331);
and UO_3316 (O_3316,N_29168,N_29562);
and UO_3317 (O_3317,N_29915,N_29335);
nor UO_3318 (O_3318,N_29830,N_29315);
xor UO_3319 (O_3319,N_29828,N_29821);
nand UO_3320 (O_3320,N_29670,N_29603);
xor UO_3321 (O_3321,N_29320,N_29416);
or UO_3322 (O_3322,N_29481,N_29586);
nor UO_3323 (O_3323,N_29508,N_29369);
xor UO_3324 (O_3324,N_29224,N_29447);
or UO_3325 (O_3325,N_29568,N_29469);
xor UO_3326 (O_3326,N_29365,N_29609);
or UO_3327 (O_3327,N_29511,N_29427);
and UO_3328 (O_3328,N_29112,N_29600);
and UO_3329 (O_3329,N_29074,N_29439);
nor UO_3330 (O_3330,N_29826,N_29905);
xor UO_3331 (O_3331,N_29668,N_29549);
xnor UO_3332 (O_3332,N_29277,N_29528);
xnor UO_3333 (O_3333,N_29916,N_29534);
nand UO_3334 (O_3334,N_29560,N_29646);
and UO_3335 (O_3335,N_29365,N_29251);
xor UO_3336 (O_3336,N_29885,N_29384);
and UO_3337 (O_3337,N_29604,N_29809);
xnor UO_3338 (O_3338,N_29388,N_29505);
nor UO_3339 (O_3339,N_29123,N_29178);
or UO_3340 (O_3340,N_29247,N_29138);
and UO_3341 (O_3341,N_29921,N_29657);
xnor UO_3342 (O_3342,N_29976,N_29701);
nand UO_3343 (O_3343,N_29097,N_29287);
or UO_3344 (O_3344,N_29581,N_29289);
nor UO_3345 (O_3345,N_29316,N_29020);
or UO_3346 (O_3346,N_29341,N_29351);
and UO_3347 (O_3347,N_29082,N_29021);
nand UO_3348 (O_3348,N_29431,N_29705);
and UO_3349 (O_3349,N_29134,N_29833);
nor UO_3350 (O_3350,N_29669,N_29909);
nand UO_3351 (O_3351,N_29387,N_29292);
nor UO_3352 (O_3352,N_29251,N_29326);
nor UO_3353 (O_3353,N_29046,N_29219);
or UO_3354 (O_3354,N_29691,N_29190);
nand UO_3355 (O_3355,N_29065,N_29188);
nand UO_3356 (O_3356,N_29391,N_29540);
or UO_3357 (O_3357,N_29523,N_29682);
or UO_3358 (O_3358,N_29819,N_29164);
or UO_3359 (O_3359,N_29069,N_29963);
or UO_3360 (O_3360,N_29004,N_29109);
or UO_3361 (O_3361,N_29569,N_29285);
nand UO_3362 (O_3362,N_29574,N_29116);
xnor UO_3363 (O_3363,N_29328,N_29323);
nand UO_3364 (O_3364,N_29740,N_29879);
nor UO_3365 (O_3365,N_29209,N_29119);
nand UO_3366 (O_3366,N_29260,N_29051);
nor UO_3367 (O_3367,N_29509,N_29816);
xor UO_3368 (O_3368,N_29059,N_29984);
or UO_3369 (O_3369,N_29047,N_29870);
nor UO_3370 (O_3370,N_29603,N_29226);
xor UO_3371 (O_3371,N_29191,N_29319);
nand UO_3372 (O_3372,N_29668,N_29003);
nand UO_3373 (O_3373,N_29168,N_29469);
nand UO_3374 (O_3374,N_29161,N_29943);
nand UO_3375 (O_3375,N_29454,N_29662);
or UO_3376 (O_3376,N_29726,N_29035);
and UO_3377 (O_3377,N_29907,N_29729);
xor UO_3378 (O_3378,N_29422,N_29128);
and UO_3379 (O_3379,N_29518,N_29473);
and UO_3380 (O_3380,N_29649,N_29858);
nand UO_3381 (O_3381,N_29806,N_29222);
xor UO_3382 (O_3382,N_29066,N_29290);
nor UO_3383 (O_3383,N_29014,N_29087);
nor UO_3384 (O_3384,N_29056,N_29652);
nand UO_3385 (O_3385,N_29780,N_29964);
or UO_3386 (O_3386,N_29889,N_29714);
nand UO_3387 (O_3387,N_29876,N_29307);
or UO_3388 (O_3388,N_29033,N_29225);
nand UO_3389 (O_3389,N_29951,N_29486);
nor UO_3390 (O_3390,N_29058,N_29811);
or UO_3391 (O_3391,N_29603,N_29354);
and UO_3392 (O_3392,N_29168,N_29762);
or UO_3393 (O_3393,N_29299,N_29665);
nor UO_3394 (O_3394,N_29083,N_29185);
and UO_3395 (O_3395,N_29763,N_29406);
xor UO_3396 (O_3396,N_29088,N_29102);
or UO_3397 (O_3397,N_29561,N_29138);
xnor UO_3398 (O_3398,N_29674,N_29628);
or UO_3399 (O_3399,N_29846,N_29467);
and UO_3400 (O_3400,N_29854,N_29568);
or UO_3401 (O_3401,N_29565,N_29012);
nor UO_3402 (O_3402,N_29049,N_29193);
and UO_3403 (O_3403,N_29524,N_29305);
xor UO_3404 (O_3404,N_29153,N_29977);
and UO_3405 (O_3405,N_29362,N_29465);
nor UO_3406 (O_3406,N_29397,N_29448);
nor UO_3407 (O_3407,N_29345,N_29040);
xor UO_3408 (O_3408,N_29612,N_29933);
xor UO_3409 (O_3409,N_29859,N_29990);
nor UO_3410 (O_3410,N_29663,N_29668);
nor UO_3411 (O_3411,N_29586,N_29615);
nand UO_3412 (O_3412,N_29701,N_29002);
or UO_3413 (O_3413,N_29651,N_29960);
nand UO_3414 (O_3414,N_29495,N_29600);
xor UO_3415 (O_3415,N_29775,N_29726);
and UO_3416 (O_3416,N_29256,N_29774);
and UO_3417 (O_3417,N_29098,N_29734);
and UO_3418 (O_3418,N_29595,N_29830);
and UO_3419 (O_3419,N_29069,N_29511);
xnor UO_3420 (O_3420,N_29588,N_29032);
and UO_3421 (O_3421,N_29036,N_29524);
and UO_3422 (O_3422,N_29111,N_29671);
and UO_3423 (O_3423,N_29026,N_29056);
and UO_3424 (O_3424,N_29497,N_29556);
nand UO_3425 (O_3425,N_29868,N_29366);
nor UO_3426 (O_3426,N_29778,N_29627);
nand UO_3427 (O_3427,N_29499,N_29579);
or UO_3428 (O_3428,N_29876,N_29718);
xnor UO_3429 (O_3429,N_29028,N_29659);
and UO_3430 (O_3430,N_29314,N_29946);
nand UO_3431 (O_3431,N_29285,N_29893);
nor UO_3432 (O_3432,N_29735,N_29451);
nor UO_3433 (O_3433,N_29069,N_29507);
nor UO_3434 (O_3434,N_29458,N_29763);
and UO_3435 (O_3435,N_29729,N_29846);
xor UO_3436 (O_3436,N_29058,N_29246);
nand UO_3437 (O_3437,N_29424,N_29615);
and UO_3438 (O_3438,N_29422,N_29735);
and UO_3439 (O_3439,N_29089,N_29900);
nand UO_3440 (O_3440,N_29370,N_29275);
nor UO_3441 (O_3441,N_29941,N_29178);
or UO_3442 (O_3442,N_29719,N_29742);
and UO_3443 (O_3443,N_29640,N_29569);
nand UO_3444 (O_3444,N_29890,N_29732);
nand UO_3445 (O_3445,N_29663,N_29971);
xor UO_3446 (O_3446,N_29566,N_29633);
and UO_3447 (O_3447,N_29934,N_29769);
or UO_3448 (O_3448,N_29864,N_29333);
and UO_3449 (O_3449,N_29769,N_29644);
xnor UO_3450 (O_3450,N_29086,N_29134);
xor UO_3451 (O_3451,N_29153,N_29176);
nand UO_3452 (O_3452,N_29746,N_29394);
nor UO_3453 (O_3453,N_29652,N_29213);
and UO_3454 (O_3454,N_29221,N_29075);
nor UO_3455 (O_3455,N_29968,N_29918);
xnor UO_3456 (O_3456,N_29258,N_29170);
and UO_3457 (O_3457,N_29136,N_29895);
and UO_3458 (O_3458,N_29160,N_29391);
nor UO_3459 (O_3459,N_29418,N_29477);
xnor UO_3460 (O_3460,N_29857,N_29497);
and UO_3461 (O_3461,N_29965,N_29384);
nand UO_3462 (O_3462,N_29039,N_29944);
and UO_3463 (O_3463,N_29053,N_29991);
xnor UO_3464 (O_3464,N_29141,N_29331);
nand UO_3465 (O_3465,N_29800,N_29070);
nand UO_3466 (O_3466,N_29509,N_29659);
and UO_3467 (O_3467,N_29392,N_29841);
nand UO_3468 (O_3468,N_29034,N_29580);
and UO_3469 (O_3469,N_29286,N_29989);
nor UO_3470 (O_3470,N_29655,N_29756);
and UO_3471 (O_3471,N_29404,N_29354);
nand UO_3472 (O_3472,N_29629,N_29797);
or UO_3473 (O_3473,N_29401,N_29415);
and UO_3474 (O_3474,N_29187,N_29430);
or UO_3475 (O_3475,N_29988,N_29730);
nand UO_3476 (O_3476,N_29004,N_29911);
nor UO_3477 (O_3477,N_29148,N_29251);
nand UO_3478 (O_3478,N_29130,N_29617);
nand UO_3479 (O_3479,N_29430,N_29645);
nand UO_3480 (O_3480,N_29980,N_29163);
nor UO_3481 (O_3481,N_29918,N_29702);
and UO_3482 (O_3482,N_29993,N_29081);
xnor UO_3483 (O_3483,N_29294,N_29832);
nor UO_3484 (O_3484,N_29860,N_29692);
xor UO_3485 (O_3485,N_29674,N_29273);
nand UO_3486 (O_3486,N_29053,N_29581);
or UO_3487 (O_3487,N_29901,N_29415);
or UO_3488 (O_3488,N_29085,N_29095);
or UO_3489 (O_3489,N_29649,N_29524);
nand UO_3490 (O_3490,N_29876,N_29054);
xor UO_3491 (O_3491,N_29571,N_29826);
and UO_3492 (O_3492,N_29421,N_29183);
nand UO_3493 (O_3493,N_29155,N_29206);
nor UO_3494 (O_3494,N_29912,N_29041);
nand UO_3495 (O_3495,N_29681,N_29825);
xor UO_3496 (O_3496,N_29227,N_29602);
or UO_3497 (O_3497,N_29611,N_29969);
or UO_3498 (O_3498,N_29929,N_29402);
or UO_3499 (O_3499,N_29760,N_29139);
endmodule