module basic_500_3000_500_40_levels_5xor_9(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
and U0 (N_0,In_341,In_409);
or U1 (N_1,In_374,In_470);
nor U2 (N_2,In_455,In_175);
or U3 (N_3,In_130,In_284);
nor U4 (N_4,In_437,In_400);
or U5 (N_5,In_469,In_5);
and U6 (N_6,In_414,In_210);
and U7 (N_7,In_264,In_166);
or U8 (N_8,In_156,In_74);
xor U9 (N_9,In_191,In_221);
and U10 (N_10,In_267,In_295);
nor U11 (N_11,In_381,In_336);
or U12 (N_12,In_215,In_200);
and U13 (N_13,In_230,In_289);
and U14 (N_14,In_9,In_79);
nand U15 (N_15,In_199,In_116);
or U16 (N_16,In_61,In_26);
and U17 (N_17,In_340,In_386);
nor U18 (N_18,In_112,In_485);
and U19 (N_19,In_178,In_316);
nor U20 (N_20,In_350,In_356);
nor U21 (N_21,In_369,In_206);
nor U22 (N_22,In_355,In_47);
and U23 (N_23,In_128,In_225);
nand U24 (N_24,In_330,In_67);
or U25 (N_25,In_313,In_59);
nand U26 (N_26,In_32,In_242);
and U27 (N_27,In_357,In_496);
or U28 (N_28,In_413,In_382);
xnor U29 (N_29,In_124,In_245);
and U30 (N_30,In_379,In_105);
nand U31 (N_31,In_183,In_464);
nand U32 (N_32,In_387,In_41);
nand U33 (N_33,In_232,In_450);
nand U34 (N_34,In_270,In_127);
nand U35 (N_35,In_351,In_332);
or U36 (N_36,In_309,In_474);
and U37 (N_37,In_261,In_222);
nand U38 (N_38,In_160,In_172);
nor U39 (N_39,In_354,In_296);
nor U40 (N_40,In_233,In_337);
xor U41 (N_41,In_12,In_248);
nand U42 (N_42,In_93,In_275);
and U43 (N_43,In_151,In_83);
xnor U44 (N_44,In_104,In_147);
nor U45 (N_45,In_235,In_461);
or U46 (N_46,In_489,In_228);
or U47 (N_47,In_158,In_258);
nand U48 (N_48,In_34,In_82);
and U49 (N_49,In_111,In_177);
or U50 (N_50,In_198,In_283);
nand U51 (N_51,In_179,In_118);
nand U52 (N_52,In_494,In_481);
nand U53 (N_53,In_287,In_407);
nor U54 (N_54,In_133,In_6);
nor U55 (N_55,In_168,In_68);
or U56 (N_56,In_72,In_152);
and U57 (N_57,In_85,In_138);
nor U58 (N_58,In_285,In_323);
nor U59 (N_59,In_203,In_227);
nand U60 (N_60,In_273,In_57);
nor U61 (N_61,In_466,In_184);
and U62 (N_62,In_364,In_398);
or U63 (N_63,In_439,In_218);
or U64 (N_64,In_463,In_266);
or U65 (N_65,In_395,In_148);
nand U66 (N_66,In_63,In_446);
xnor U67 (N_67,In_176,In_243);
or U68 (N_68,In_171,In_484);
xnor U69 (N_69,In_102,In_333);
nor U70 (N_70,In_317,In_327);
nor U71 (N_71,In_58,In_107);
or U72 (N_72,In_87,In_373);
nor U73 (N_73,In_402,In_231);
nor U74 (N_74,In_119,In_475);
and U75 (N_75,In_279,In_54);
nor U76 (N_76,In_89,In_318);
or U77 (N_77,N_15,In_299);
nand U78 (N_78,In_346,In_165);
nor U79 (N_79,In_77,In_23);
or U80 (N_80,In_43,N_22);
nand U81 (N_81,In_201,In_181);
nor U82 (N_82,In_277,In_433);
nand U83 (N_83,N_8,In_10);
nand U84 (N_84,In_448,In_249);
and U85 (N_85,In_352,In_189);
or U86 (N_86,In_305,In_390);
nand U87 (N_87,In_281,In_126);
nor U88 (N_88,In_39,N_56);
and U89 (N_89,N_33,N_38);
and U90 (N_90,In_211,In_367);
or U91 (N_91,In_55,In_456);
or U92 (N_92,In_223,In_343);
nand U93 (N_93,In_239,In_458);
xnor U94 (N_94,In_292,N_2);
and U95 (N_95,In_38,In_302);
and U96 (N_96,In_457,In_92);
and U97 (N_97,In_88,In_94);
xnor U98 (N_98,N_25,In_120);
nor U99 (N_99,N_44,In_27);
and U100 (N_100,In_440,N_24);
nor U101 (N_101,N_20,In_271);
nor U102 (N_102,In_384,N_43);
nand U103 (N_103,In_197,In_146);
or U104 (N_104,In_453,In_306);
xor U105 (N_105,In_194,N_9);
and U106 (N_106,In_28,In_49);
nand U107 (N_107,In_0,In_399);
and U108 (N_108,In_434,In_263);
or U109 (N_109,N_31,N_55);
nor U110 (N_110,In_91,In_1);
xor U111 (N_111,In_52,In_62);
nand U112 (N_112,In_244,In_497);
nand U113 (N_113,In_108,In_449);
and U114 (N_114,N_69,In_408);
or U115 (N_115,In_412,In_321);
or U116 (N_116,In_425,In_269);
nor U117 (N_117,In_100,In_159);
or U118 (N_118,In_491,N_13);
xor U119 (N_119,In_220,In_44);
nand U120 (N_120,In_103,In_265);
and U121 (N_121,In_372,In_334);
nor U122 (N_122,N_1,In_46);
or U123 (N_123,In_472,In_136);
or U124 (N_124,In_335,In_297);
nor U125 (N_125,In_375,In_149);
xor U126 (N_126,In_213,In_143);
and U127 (N_127,N_52,In_417);
or U128 (N_128,N_4,In_262);
xnor U129 (N_129,In_288,In_25);
nand U130 (N_130,In_473,In_393);
nand U131 (N_131,In_14,N_42);
xor U132 (N_132,In_422,In_345);
or U133 (N_133,In_445,In_274);
xor U134 (N_134,N_35,In_421);
nor U135 (N_135,In_349,In_234);
or U136 (N_136,In_339,N_57);
or U137 (N_137,In_17,N_61);
nand U138 (N_138,In_430,N_12);
or U139 (N_139,In_250,In_362);
nand U140 (N_140,N_49,In_388);
nand U141 (N_141,In_499,In_174);
xnor U142 (N_142,In_256,N_47);
and U143 (N_143,In_212,In_33);
or U144 (N_144,In_122,N_40);
nor U145 (N_145,In_442,In_188);
nor U146 (N_146,In_224,In_76);
nand U147 (N_147,In_241,In_348);
or U148 (N_148,In_467,In_110);
and U149 (N_149,In_483,In_29);
nor U150 (N_150,In_65,In_361);
nand U151 (N_151,N_16,N_109);
or U152 (N_152,In_180,In_479);
xor U153 (N_153,In_278,In_240);
and U154 (N_154,In_419,In_8);
nand U155 (N_155,In_157,N_96);
or U156 (N_156,In_385,N_53);
nand U157 (N_157,In_161,N_28);
nor U158 (N_158,N_6,In_99);
and U159 (N_159,In_209,In_435);
and U160 (N_160,N_97,In_308);
and U161 (N_161,N_36,In_319);
or U162 (N_162,N_60,In_202);
nand U163 (N_163,N_115,In_314);
xor U164 (N_164,N_82,In_193);
nor U165 (N_165,In_251,In_182);
and U166 (N_166,In_404,N_21);
nand U167 (N_167,In_150,In_84);
xor U168 (N_168,In_252,In_31);
nor U169 (N_169,N_144,In_490);
or U170 (N_170,In_95,In_298);
nand U171 (N_171,In_492,N_107);
and U172 (N_172,In_392,In_286);
nor U173 (N_173,N_37,In_42);
nand U174 (N_174,In_56,N_72);
or U175 (N_175,N_100,N_75);
xnor U176 (N_176,In_410,In_66);
or U177 (N_177,N_67,In_344);
or U178 (N_178,In_301,In_80);
and U179 (N_179,N_79,In_71);
nand U180 (N_180,N_126,In_98);
or U181 (N_181,N_84,In_24);
or U182 (N_182,N_102,N_135);
nor U183 (N_183,N_128,In_64);
nand U184 (N_184,In_69,In_73);
nor U185 (N_185,N_32,In_13);
or U186 (N_186,In_377,In_101);
and U187 (N_187,N_106,In_363);
and U188 (N_188,N_85,In_78);
and U189 (N_189,In_238,In_324);
nor U190 (N_190,In_204,N_71);
nor U191 (N_191,In_476,In_145);
xnor U192 (N_192,In_229,In_257);
nor U193 (N_193,N_95,In_423);
xnor U194 (N_194,In_81,In_358);
and U195 (N_195,In_125,In_429);
and U196 (N_196,In_187,In_115);
or U197 (N_197,In_4,N_54);
nor U198 (N_198,N_46,In_15);
or U199 (N_199,In_163,In_405);
xnor U200 (N_200,N_124,In_438);
or U201 (N_201,In_451,In_291);
or U202 (N_202,In_22,In_452);
nand U203 (N_203,In_406,In_394);
and U204 (N_204,In_311,N_108);
or U205 (N_205,In_331,In_154);
and U206 (N_206,In_236,N_10);
or U207 (N_207,In_418,In_131);
xor U208 (N_208,N_103,N_139);
or U209 (N_209,In_460,N_39);
and U210 (N_210,In_282,N_125);
nor U211 (N_211,In_444,In_376);
nor U212 (N_212,N_149,In_214);
or U213 (N_213,In_35,In_416);
or U214 (N_214,N_81,In_135);
and U215 (N_215,N_63,In_370);
xnor U216 (N_216,N_17,In_359);
nor U217 (N_217,N_26,In_253);
nor U218 (N_218,In_487,N_59);
nand U219 (N_219,In_190,In_139);
and U220 (N_220,In_328,N_89);
or U221 (N_221,In_132,N_23);
and U222 (N_222,N_127,In_217);
and U223 (N_223,In_97,In_36);
and U224 (N_224,In_259,In_255);
and U225 (N_225,In_186,In_325);
nor U226 (N_226,N_99,N_150);
and U227 (N_227,N_122,In_424);
nor U228 (N_228,N_206,In_498);
nand U229 (N_229,In_30,N_216);
nand U230 (N_230,In_342,N_200);
nor U231 (N_231,N_188,In_162);
and U232 (N_232,In_48,In_276);
nor U233 (N_233,In_195,N_147);
and U234 (N_234,N_155,N_164);
or U235 (N_235,In_300,N_189);
nand U236 (N_236,In_427,In_478);
and U237 (N_237,N_11,N_65);
nand U238 (N_238,N_76,In_468);
nand U239 (N_239,In_268,In_431);
or U240 (N_240,N_90,N_166);
and U241 (N_241,In_420,N_172);
nor U242 (N_242,In_219,N_142);
or U243 (N_243,In_304,N_130);
and U244 (N_244,N_113,In_3);
nand U245 (N_245,In_389,N_119);
xor U246 (N_246,N_80,N_198);
and U247 (N_247,In_428,In_226);
and U248 (N_248,N_215,In_216);
nand U249 (N_249,N_160,N_211);
or U250 (N_250,In_353,In_482);
or U251 (N_251,N_116,N_214);
nand U252 (N_252,N_121,N_94);
or U253 (N_253,N_104,In_205);
and U254 (N_254,In_155,N_145);
or U255 (N_255,In_365,In_169);
nand U256 (N_256,In_51,In_477);
nand U257 (N_257,N_201,N_171);
or U258 (N_258,N_62,In_164);
nand U259 (N_259,In_96,N_123);
and U260 (N_260,In_170,In_109);
nor U261 (N_261,In_134,In_436);
nor U262 (N_262,In_123,In_45);
nand U263 (N_263,N_179,In_53);
nor U264 (N_264,In_303,N_202);
xor U265 (N_265,N_30,In_153);
xnor U266 (N_266,In_16,N_41);
xor U267 (N_267,In_167,In_454);
and U268 (N_268,N_77,N_87);
or U269 (N_269,N_70,In_480);
and U270 (N_270,N_209,N_18);
nand U271 (N_271,In_142,In_60);
nor U272 (N_272,N_111,In_307);
or U273 (N_273,N_140,N_138);
and U274 (N_274,N_173,N_205);
and U275 (N_275,N_213,N_45);
and U276 (N_276,N_180,N_165);
nor U277 (N_277,N_212,N_78);
nand U278 (N_278,In_397,N_158);
nand U279 (N_279,N_153,N_88);
xor U280 (N_280,N_137,In_21);
and U281 (N_281,In_315,In_310);
and U282 (N_282,In_20,N_3);
nor U283 (N_283,N_182,In_192);
nor U284 (N_284,N_162,N_91);
nand U285 (N_285,N_34,N_156);
nand U286 (N_286,In_141,In_50);
nand U287 (N_287,In_432,N_51);
nand U288 (N_288,In_459,N_148);
nor U289 (N_289,In_173,In_488);
and U290 (N_290,N_132,N_157);
nand U291 (N_291,N_220,N_83);
nand U292 (N_292,N_152,In_144);
or U293 (N_293,N_151,N_110);
and U294 (N_294,In_86,In_75);
nor U295 (N_295,N_185,N_203);
nor U296 (N_296,In_106,In_129);
or U297 (N_297,In_90,N_193);
and U298 (N_298,N_141,In_207);
and U299 (N_299,In_18,In_247);
xor U300 (N_300,N_258,N_181);
or U301 (N_301,In_293,N_222);
nor U302 (N_302,N_133,N_273);
or U303 (N_303,N_221,N_262);
nor U304 (N_304,N_272,N_264);
nor U305 (N_305,N_19,N_73);
nor U306 (N_306,In_465,N_256);
or U307 (N_307,In_383,In_447);
and U308 (N_308,N_282,N_295);
or U309 (N_309,N_208,N_283);
nand U310 (N_310,N_240,N_58);
nand U311 (N_311,In_280,N_86);
nand U312 (N_312,N_187,N_217);
nand U313 (N_313,In_411,In_326);
and U314 (N_314,N_199,N_292);
nor U315 (N_315,In_117,In_208);
nor U316 (N_316,N_218,N_279);
xnor U317 (N_317,N_249,N_259);
xnor U318 (N_318,N_252,N_197);
nor U319 (N_319,N_219,In_70);
nor U320 (N_320,N_177,N_114);
or U321 (N_321,In_19,In_371);
or U322 (N_322,In_401,N_183);
or U323 (N_323,N_266,N_268);
and U324 (N_324,In_7,N_0);
and U325 (N_325,N_296,In_396);
nor U326 (N_326,N_168,N_233);
nand U327 (N_327,N_261,N_143);
and U328 (N_328,In_380,N_297);
or U329 (N_329,In_246,N_207);
nand U330 (N_330,N_248,In_137);
xnor U331 (N_331,N_294,N_178);
nand U332 (N_332,N_284,N_254);
nand U333 (N_333,N_7,N_299);
and U334 (N_334,In_260,N_257);
or U335 (N_335,N_280,In_471);
nor U336 (N_336,N_134,N_191);
nand U337 (N_337,N_270,In_196);
and U338 (N_338,In_113,In_2);
nand U339 (N_339,In_378,N_289);
nand U340 (N_340,N_242,N_192);
or U341 (N_341,N_29,N_255);
nand U342 (N_342,N_290,N_64);
and U343 (N_343,N_234,In_360);
xor U344 (N_344,N_271,In_495);
or U345 (N_345,N_239,In_347);
nand U346 (N_346,N_170,N_174);
nor U347 (N_347,In_272,N_260);
or U348 (N_348,N_226,N_246);
or U349 (N_349,N_167,N_291);
xnor U350 (N_350,N_210,N_204);
nand U351 (N_351,N_175,N_278);
or U352 (N_352,N_276,N_154);
and U353 (N_353,N_269,N_245);
or U354 (N_354,N_232,N_223);
and U355 (N_355,N_68,N_93);
nand U356 (N_356,N_92,N_190);
and U357 (N_357,N_267,N_163);
or U358 (N_358,In_441,In_426);
nand U359 (N_359,In_237,In_329);
nor U360 (N_360,In_40,N_288);
xor U361 (N_361,N_237,In_254);
nand U362 (N_362,N_244,N_227);
nor U363 (N_363,In_140,N_236);
xnor U364 (N_364,N_275,N_27);
nor U365 (N_365,In_294,N_231);
and U366 (N_366,In_462,In_185);
xnor U367 (N_367,In_320,In_322);
nand U368 (N_368,N_228,In_486);
nor U369 (N_369,N_263,N_285);
xor U370 (N_370,N_136,N_14);
xnor U371 (N_371,In_415,N_229);
nand U372 (N_372,N_281,N_131);
and U373 (N_373,N_169,N_277);
nand U374 (N_374,N_265,In_338);
and U375 (N_375,N_235,N_331);
nor U376 (N_376,In_443,In_403);
or U377 (N_377,N_330,N_230);
xnor U378 (N_378,N_332,N_184);
nor U379 (N_379,In_368,N_105);
nand U380 (N_380,N_176,N_118);
and U381 (N_381,N_359,N_370);
and U382 (N_382,N_306,N_161);
and U383 (N_383,N_329,N_350);
or U384 (N_384,N_324,N_243);
or U385 (N_385,N_363,N_374);
xnor U386 (N_386,N_310,N_354);
or U387 (N_387,N_314,N_101);
nor U388 (N_388,N_336,N_318);
nand U389 (N_389,N_50,N_301);
or U390 (N_390,N_326,N_305);
nor U391 (N_391,N_333,N_186);
or U392 (N_392,N_319,N_274);
nor U393 (N_393,N_347,N_308);
or U394 (N_394,N_304,N_241);
nor U395 (N_395,N_341,N_335);
and U396 (N_396,In_11,N_364);
xnor U397 (N_397,In_114,N_5);
nor U398 (N_398,N_112,N_348);
nand U399 (N_399,N_195,N_365);
nor U400 (N_400,N_74,In_121);
or U401 (N_401,N_194,N_117);
nor U402 (N_402,N_303,N_307);
or U403 (N_403,N_321,In_391);
and U404 (N_404,N_372,N_361);
and U405 (N_405,N_146,N_251);
and U406 (N_406,N_327,N_367);
and U407 (N_407,N_343,N_371);
nand U408 (N_408,N_309,N_316);
nand U409 (N_409,N_224,N_120);
or U410 (N_410,N_373,N_346);
or U411 (N_411,N_313,N_302);
or U412 (N_412,N_66,N_300);
or U413 (N_413,N_98,In_37);
or U414 (N_414,N_357,N_356);
xnor U415 (N_415,N_325,N_48);
nor U416 (N_416,N_286,N_334);
nand U417 (N_417,N_337,N_159);
and U418 (N_418,N_312,N_358);
nand U419 (N_419,N_315,N_353);
or U420 (N_420,N_311,N_328);
nand U421 (N_421,In_493,N_293);
and U422 (N_422,N_345,N_238);
and U423 (N_423,N_355,N_225);
nor U424 (N_424,In_366,N_322);
xnor U425 (N_425,N_360,N_287);
or U426 (N_426,N_339,N_368);
nand U427 (N_427,N_196,N_253);
or U428 (N_428,N_351,N_250);
xnor U429 (N_429,N_344,N_342);
nor U430 (N_430,In_312,N_366);
nand U431 (N_431,N_129,In_290);
nor U432 (N_432,N_323,N_247);
nor U433 (N_433,N_349,N_338);
or U434 (N_434,N_317,N_340);
nor U435 (N_435,N_298,N_362);
and U436 (N_436,N_369,N_352);
and U437 (N_437,N_320,N_327);
or U438 (N_438,N_186,N_351);
and U439 (N_439,N_274,N_243);
nor U440 (N_440,N_238,N_348);
nor U441 (N_441,N_105,N_332);
xnor U442 (N_442,N_337,N_324);
nand U443 (N_443,N_320,N_120);
or U444 (N_444,N_251,N_48);
or U445 (N_445,N_319,N_331);
or U446 (N_446,N_340,N_186);
or U447 (N_447,N_66,N_50);
and U448 (N_448,N_48,N_194);
nand U449 (N_449,N_371,N_293);
nand U450 (N_450,N_389,N_404);
or U451 (N_451,N_427,N_418);
and U452 (N_452,N_432,N_433);
nor U453 (N_453,N_428,N_436);
and U454 (N_454,N_414,N_443);
or U455 (N_455,N_441,N_385);
nor U456 (N_456,N_383,N_382);
nand U457 (N_457,N_381,N_415);
nor U458 (N_458,N_417,N_391);
nand U459 (N_459,N_384,N_424);
nor U460 (N_460,N_406,N_430);
nor U461 (N_461,N_425,N_379);
nand U462 (N_462,N_402,N_449);
and U463 (N_463,N_405,N_407);
or U464 (N_464,N_378,N_412);
xor U465 (N_465,N_392,N_437);
xor U466 (N_466,N_400,N_442);
nor U467 (N_467,N_390,N_419);
and U468 (N_468,N_396,N_440);
or U469 (N_469,N_397,N_387);
or U470 (N_470,N_408,N_380);
and U471 (N_471,N_438,N_426);
or U472 (N_472,N_403,N_399);
nand U473 (N_473,N_416,N_446);
xnor U474 (N_474,N_444,N_411);
and U475 (N_475,N_422,N_435);
or U476 (N_476,N_377,N_409);
or U477 (N_477,N_413,N_393);
nand U478 (N_478,N_395,N_431);
or U479 (N_479,N_410,N_386);
nor U480 (N_480,N_394,N_447);
and U481 (N_481,N_388,N_423);
xnor U482 (N_482,N_434,N_439);
nor U483 (N_483,N_448,N_375);
and U484 (N_484,N_420,N_429);
xnor U485 (N_485,N_398,N_445);
nand U486 (N_486,N_376,N_421);
nand U487 (N_487,N_401,N_424);
or U488 (N_488,N_386,N_442);
or U489 (N_489,N_417,N_400);
nor U490 (N_490,N_447,N_423);
nor U491 (N_491,N_426,N_420);
nor U492 (N_492,N_391,N_411);
xnor U493 (N_493,N_441,N_429);
or U494 (N_494,N_429,N_394);
and U495 (N_495,N_409,N_392);
and U496 (N_496,N_382,N_421);
nor U497 (N_497,N_445,N_441);
nor U498 (N_498,N_424,N_382);
nand U499 (N_499,N_392,N_395);
or U500 (N_500,N_403,N_398);
xnor U501 (N_501,N_424,N_398);
nand U502 (N_502,N_447,N_444);
nor U503 (N_503,N_434,N_416);
and U504 (N_504,N_397,N_445);
nand U505 (N_505,N_400,N_443);
nand U506 (N_506,N_380,N_391);
nand U507 (N_507,N_383,N_381);
nor U508 (N_508,N_431,N_400);
nand U509 (N_509,N_431,N_399);
nor U510 (N_510,N_427,N_398);
nor U511 (N_511,N_416,N_414);
nor U512 (N_512,N_439,N_411);
nor U513 (N_513,N_387,N_449);
and U514 (N_514,N_426,N_398);
nor U515 (N_515,N_396,N_381);
and U516 (N_516,N_397,N_380);
nand U517 (N_517,N_425,N_404);
nor U518 (N_518,N_439,N_416);
and U519 (N_519,N_430,N_425);
or U520 (N_520,N_425,N_402);
and U521 (N_521,N_447,N_417);
and U522 (N_522,N_401,N_395);
and U523 (N_523,N_436,N_438);
or U524 (N_524,N_437,N_394);
nand U525 (N_525,N_502,N_488);
nand U526 (N_526,N_506,N_521);
nand U527 (N_527,N_523,N_504);
nor U528 (N_528,N_483,N_497);
and U529 (N_529,N_505,N_491);
xor U530 (N_530,N_492,N_509);
nor U531 (N_531,N_501,N_463);
nor U532 (N_532,N_519,N_462);
nor U533 (N_533,N_469,N_478);
nor U534 (N_534,N_461,N_477);
nor U535 (N_535,N_485,N_511);
and U536 (N_536,N_470,N_512);
nand U537 (N_537,N_494,N_472);
nand U538 (N_538,N_503,N_522);
xnor U539 (N_539,N_476,N_475);
and U540 (N_540,N_513,N_493);
nor U541 (N_541,N_452,N_474);
and U542 (N_542,N_458,N_450);
nand U543 (N_543,N_465,N_466);
nand U544 (N_544,N_482,N_464);
or U545 (N_545,N_473,N_467);
nor U546 (N_546,N_496,N_516);
nand U547 (N_547,N_514,N_520);
or U548 (N_548,N_518,N_487);
nor U549 (N_549,N_498,N_468);
and U550 (N_550,N_479,N_507);
or U551 (N_551,N_486,N_454);
and U552 (N_552,N_451,N_471);
or U553 (N_553,N_484,N_457);
nand U554 (N_554,N_453,N_524);
xnor U555 (N_555,N_490,N_489);
nor U556 (N_556,N_515,N_499);
or U557 (N_557,N_481,N_500);
nand U558 (N_558,N_460,N_510);
or U559 (N_559,N_495,N_508);
nand U560 (N_560,N_480,N_456);
or U561 (N_561,N_517,N_459);
and U562 (N_562,N_455,N_490);
and U563 (N_563,N_494,N_481);
or U564 (N_564,N_470,N_489);
xor U565 (N_565,N_509,N_499);
and U566 (N_566,N_468,N_479);
nand U567 (N_567,N_493,N_450);
nand U568 (N_568,N_487,N_519);
and U569 (N_569,N_523,N_516);
and U570 (N_570,N_484,N_473);
nand U571 (N_571,N_454,N_508);
nor U572 (N_572,N_472,N_490);
nor U573 (N_573,N_467,N_455);
nor U574 (N_574,N_452,N_473);
and U575 (N_575,N_494,N_524);
xnor U576 (N_576,N_459,N_516);
nand U577 (N_577,N_497,N_522);
and U578 (N_578,N_471,N_477);
nor U579 (N_579,N_472,N_457);
nor U580 (N_580,N_490,N_460);
nor U581 (N_581,N_463,N_508);
xor U582 (N_582,N_498,N_510);
or U583 (N_583,N_523,N_511);
or U584 (N_584,N_499,N_516);
nand U585 (N_585,N_453,N_470);
or U586 (N_586,N_455,N_520);
nor U587 (N_587,N_497,N_521);
nor U588 (N_588,N_494,N_492);
nor U589 (N_589,N_461,N_480);
nand U590 (N_590,N_486,N_459);
and U591 (N_591,N_522,N_451);
nand U592 (N_592,N_464,N_507);
or U593 (N_593,N_490,N_476);
nor U594 (N_594,N_464,N_478);
or U595 (N_595,N_488,N_521);
or U596 (N_596,N_480,N_451);
nand U597 (N_597,N_456,N_502);
and U598 (N_598,N_502,N_494);
nand U599 (N_599,N_479,N_452);
nor U600 (N_600,N_526,N_590);
nand U601 (N_601,N_581,N_551);
or U602 (N_602,N_592,N_571);
xnor U603 (N_603,N_548,N_595);
nand U604 (N_604,N_553,N_554);
nor U605 (N_605,N_579,N_536);
nand U606 (N_606,N_550,N_538);
and U607 (N_607,N_563,N_528);
nor U608 (N_608,N_573,N_566);
or U609 (N_609,N_546,N_570);
nand U610 (N_610,N_586,N_575);
and U611 (N_611,N_558,N_545);
or U612 (N_612,N_582,N_547);
xnor U613 (N_613,N_529,N_543);
nand U614 (N_614,N_576,N_557);
and U615 (N_615,N_585,N_569);
and U616 (N_616,N_532,N_584);
nor U617 (N_617,N_561,N_597);
nor U618 (N_618,N_580,N_591);
xnor U619 (N_619,N_589,N_527);
or U620 (N_620,N_572,N_531);
xor U621 (N_621,N_544,N_596);
xor U622 (N_622,N_530,N_555);
nor U623 (N_623,N_598,N_574);
or U624 (N_624,N_542,N_560);
or U625 (N_625,N_534,N_593);
xnor U626 (N_626,N_577,N_578);
nor U627 (N_627,N_533,N_583);
nand U628 (N_628,N_535,N_568);
nand U629 (N_629,N_537,N_540);
or U630 (N_630,N_565,N_559);
nand U631 (N_631,N_541,N_594);
and U632 (N_632,N_556,N_567);
xnor U633 (N_633,N_525,N_552);
or U634 (N_634,N_564,N_588);
and U635 (N_635,N_562,N_549);
nand U636 (N_636,N_539,N_599);
nor U637 (N_637,N_587,N_542);
nor U638 (N_638,N_589,N_583);
and U639 (N_639,N_582,N_571);
and U640 (N_640,N_560,N_590);
nor U641 (N_641,N_561,N_567);
and U642 (N_642,N_593,N_544);
nor U643 (N_643,N_569,N_534);
nand U644 (N_644,N_525,N_566);
nor U645 (N_645,N_586,N_561);
xnor U646 (N_646,N_537,N_571);
xnor U647 (N_647,N_527,N_578);
xor U648 (N_648,N_555,N_525);
xor U649 (N_649,N_564,N_526);
xor U650 (N_650,N_591,N_554);
nor U651 (N_651,N_539,N_593);
nand U652 (N_652,N_534,N_570);
or U653 (N_653,N_552,N_536);
or U654 (N_654,N_599,N_585);
xor U655 (N_655,N_560,N_579);
nor U656 (N_656,N_570,N_582);
and U657 (N_657,N_548,N_534);
or U658 (N_658,N_579,N_546);
xor U659 (N_659,N_536,N_566);
and U660 (N_660,N_566,N_547);
and U661 (N_661,N_538,N_590);
and U662 (N_662,N_597,N_557);
nor U663 (N_663,N_571,N_588);
and U664 (N_664,N_578,N_531);
nor U665 (N_665,N_542,N_548);
xor U666 (N_666,N_530,N_542);
and U667 (N_667,N_582,N_538);
xor U668 (N_668,N_567,N_537);
or U669 (N_669,N_594,N_570);
nand U670 (N_670,N_538,N_589);
nor U671 (N_671,N_546,N_589);
nor U672 (N_672,N_564,N_596);
or U673 (N_673,N_567,N_564);
and U674 (N_674,N_589,N_565);
or U675 (N_675,N_606,N_625);
nand U676 (N_676,N_670,N_639);
nand U677 (N_677,N_628,N_646);
or U678 (N_678,N_616,N_602);
or U679 (N_679,N_601,N_612);
nor U680 (N_680,N_656,N_643);
or U681 (N_681,N_659,N_604);
nand U682 (N_682,N_610,N_623);
nand U683 (N_683,N_600,N_609);
or U684 (N_684,N_627,N_634);
nor U685 (N_685,N_631,N_648);
and U686 (N_686,N_647,N_674);
nand U687 (N_687,N_671,N_669);
or U688 (N_688,N_649,N_663);
xor U689 (N_689,N_621,N_641);
nor U690 (N_690,N_603,N_629);
nor U691 (N_691,N_662,N_660);
nand U692 (N_692,N_622,N_624);
nand U693 (N_693,N_657,N_658);
or U694 (N_694,N_608,N_630);
nand U695 (N_695,N_650,N_617);
and U696 (N_696,N_655,N_651);
nand U697 (N_697,N_652,N_636);
and U698 (N_698,N_626,N_638);
nand U699 (N_699,N_614,N_618);
or U700 (N_700,N_633,N_611);
nand U701 (N_701,N_654,N_619);
or U702 (N_702,N_642,N_672);
or U703 (N_703,N_640,N_668);
nand U704 (N_704,N_653,N_667);
nand U705 (N_705,N_673,N_664);
xnor U706 (N_706,N_644,N_637);
nor U707 (N_707,N_666,N_632);
or U708 (N_708,N_620,N_615);
nor U709 (N_709,N_645,N_613);
nor U710 (N_710,N_665,N_635);
nand U711 (N_711,N_607,N_605);
and U712 (N_712,N_661,N_622);
nand U713 (N_713,N_666,N_640);
nor U714 (N_714,N_640,N_667);
or U715 (N_715,N_638,N_657);
and U716 (N_716,N_648,N_627);
nor U717 (N_717,N_621,N_606);
or U718 (N_718,N_613,N_669);
nand U719 (N_719,N_625,N_627);
nor U720 (N_720,N_612,N_658);
or U721 (N_721,N_620,N_647);
or U722 (N_722,N_611,N_613);
or U723 (N_723,N_641,N_662);
nor U724 (N_724,N_672,N_614);
and U725 (N_725,N_673,N_614);
or U726 (N_726,N_626,N_667);
nand U727 (N_727,N_626,N_610);
and U728 (N_728,N_637,N_617);
nand U729 (N_729,N_638,N_631);
nor U730 (N_730,N_604,N_616);
and U731 (N_731,N_638,N_623);
and U732 (N_732,N_671,N_674);
nand U733 (N_733,N_648,N_625);
and U734 (N_734,N_660,N_673);
and U735 (N_735,N_662,N_636);
and U736 (N_736,N_613,N_658);
xnor U737 (N_737,N_640,N_661);
nor U738 (N_738,N_640,N_673);
nor U739 (N_739,N_658,N_668);
or U740 (N_740,N_621,N_600);
and U741 (N_741,N_617,N_672);
and U742 (N_742,N_618,N_627);
nor U743 (N_743,N_627,N_602);
or U744 (N_744,N_656,N_650);
and U745 (N_745,N_655,N_661);
nor U746 (N_746,N_651,N_626);
nor U747 (N_747,N_654,N_648);
xnor U748 (N_748,N_614,N_626);
nor U749 (N_749,N_673,N_616);
nor U750 (N_750,N_679,N_710);
xnor U751 (N_751,N_720,N_740);
xnor U752 (N_752,N_692,N_735);
and U753 (N_753,N_737,N_678);
nor U754 (N_754,N_742,N_707);
or U755 (N_755,N_726,N_686);
or U756 (N_756,N_687,N_731);
nor U757 (N_757,N_748,N_722);
nand U758 (N_758,N_729,N_709);
nand U759 (N_759,N_714,N_683);
xnor U760 (N_760,N_702,N_705);
or U761 (N_761,N_747,N_684);
or U762 (N_762,N_718,N_682);
and U763 (N_763,N_703,N_715);
nand U764 (N_764,N_739,N_676);
and U765 (N_765,N_711,N_749);
nor U766 (N_766,N_681,N_738);
and U767 (N_767,N_698,N_733);
nor U768 (N_768,N_734,N_725);
and U769 (N_769,N_685,N_728);
nand U770 (N_770,N_694,N_732);
nand U771 (N_771,N_704,N_696);
nor U772 (N_772,N_744,N_713);
xor U773 (N_773,N_719,N_712);
nand U774 (N_774,N_697,N_700);
and U775 (N_775,N_717,N_736);
nor U776 (N_776,N_680,N_706);
nor U777 (N_777,N_699,N_741);
and U778 (N_778,N_691,N_727);
or U779 (N_779,N_701,N_693);
or U780 (N_780,N_689,N_675);
nor U781 (N_781,N_743,N_688);
or U782 (N_782,N_677,N_721);
and U783 (N_783,N_716,N_723);
nor U784 (N_784,N_730,N_724);
or U785 (N_785,N_746,N_708);
xor U786 (N_786,N_695,N_745);
or U787 (N_787,N_690,N_736);
nor U788 (N_788,N_675,N_687);
and U789 (N_789,N_738,N_675);
or U790 (N_790,N_734,N_733);
and U791 (N_791,N_688,N_722);
nand U792 (N_792,N_723,N_698);
or U793 (N_793,N_692,N_696);
nor U794 (N_794,N_701,N_713);
xor U795 (N_795,N_714,N_680);
or U796 (N_796,N_693,N_740);
xnor U797 (N_797,N_697,N_740);
nor U798 (N_798,N_749,N_705);
and U799 (N_799,N_678,N_677);
or U800 (N_800,N_735,N_738);
or U801 (N_801,N_724,N_734);
nor U802 (N_802,N_709,N_745);
nor U803 (N_803,N_708,N_723);
or U804 (N_804,N_705,N_745);
nand U805 (N_805,N_731,N_698);
or U806 (N_806,N_715,N_729);
or U807 (N_807,N_740,N_721);
nor U808 (N_808,N_731,N_702);
and U809 (N_809,N_707,N_740);
nor U810 (N_810,N_734,N_714);
nand U811 (N_811,N_676,N_685);
nand U812 (N_812,N_702,N_706);
or U813 (N_813,N_723,N_736);
nor U814 (N_814,N_700,N_739);
and U815 (N_815,N_687,N_706);
nand U816 (N_816,N_721,N_688);
nand U817 (N_817,N_695,N_709);
nor U818 (N_818,N_709,N_684);
nand U819 (N_819,N_707,N_702);
nor U820 (N_820,N_707,N_703);
or U821 (N_821,N_723,N_696);
nor U822 (N_822,N_709,N_691);
or U823 (N_823,N_737,N_699);
or U824 (N_824,N_715,N_679);
nor U825 (N_825,N_791,N_762);
nand U826 (N_826,N_781,N_810);
nand U827 (N_827,N_757,N_807);
and U828 (N_828,N_759,N_761);
and U829 (N_829,N_769,N_806);
nor U830 (N_830,N_782,N_798);
nand U831 (N_831,N_805,N_787);
and U832 (N_832,N_754,N_767);
xor U833 (N_833,N_758,N_776);
xnor U834 (N_834,N_760,N_779);
or U835 (N_835,N_768,N_770);
and U836 (N_836,N_772,N_788);
or U837 (N_837,N_751,N_793);
xor U838 (N_838,N_765,N_816);
nor U839 (N_839,N_773,N_764);
xnor U840 (N_840,N_778,N_797);
nand U841 (N_841,N_795,N_802);
or U842 (N_842,N_771,N_820);
and U843 (N_843,N_766,N_821);
and U844 (N_844,N_799,N_811);
nand U845 (N_845,N_750,N_824);
and U846 (N_846,N_775,N_804);
and U847 (N_847,N_783,N_809);
or U848 (N_848,N_808,N_815);
nand U849 (N_849,N_813,N_819);
nand U850 (N_850,N_814,N_817);
or U851 (N_851,N_763,N_818);
and U852 (N_852,N_755,N_756);
nand U853 (N_853,N_801,N_780);
and U854 (N_854,N_777,N_784);
nand U855 (N_855,N_785,N_800);
nand U856 (N_856,N_794,N_774);
and U857 (N_857,N_753,N_790);
nor U858 (N_858,N_823,N_822);
nand U859 (N_859,N_789,N_812);
or U860 (N_860,N_786,N_792);
nor U861 (N_861,N_752,N_796);
or U862 (N_862,N_803,N_794);
xnor U863 (N_863,N_817,N_753);
nand U864 (N_864,N_801,N_769);
nand U865 (N_865,N_764,N_822);
nor U866 (N_866,N_774,N_771);
xor U867 (N_867,N_793,N_816);
nor U868 (N_868,N_801,N_751);
or U869 (N_869,N_764,N_750);
or U870 (N_870,N_788,N_819);
nor U871 (N_871,N_767,N_816);
nand U872 (N_872,N_776,N_792);
and U873 (N_873,N_762,N_754);
and U874 (N_874,N_765,N_783);
or U875 (N_875,N_751,N_750);
xor U876 (N_876,N_777,N_795);
xnor U877 (N_877,N_764,N_760);
nand U878 (N_878,N_809,N_801);
and U879 (N_879,N_786,N_805);
nor U880 (N_880,N_782,N_807);
nand U881 (N_881,N_813,N_768);
nor U882 (N_882,N_799,N_768);
or U883 (N_883,N_772,N_777);
xor U884 (N_884,N_793,N_809);
and U885 (N_885,N_808,N_809);
or U886 (N_886,N_797,N_757);
nor U887 (N_887,N_815,N_786);
or U888 (N_888,N_796,N_820);
and U889 (N_889,N_795,N_775);
and U890 (N_890,N_816,N_809);
nor U891 (N_891,N_794,N_802);
and U892 (N_892,N_757,N_794);
nor U893 (N_893,N_812,N_783);
xnor U894 (N_894,N_755,N_798);
nor U895 (N_895,N_766,N_780);
or U896 (N_896,N_791,N_764);
nand U897 (N_897,N_786,N_794);
xor U898 (N_898,N_778,N_801);
or U899 (N_899,N_812,N_813);
nor U900 (N_900,N_884,N_899);
or U901 (N_901,N_896,N_844);
nor U902 (N_902,N_825,N_859);
or U903 (N_903,N_846,N_882);
and U904 (N_904,N_860,N_848);
xor U905 (N_905,N_864,N_829);
or U906 (N_906,N_894,N_838);
or U907 (N_907,N_836,N_843);
nor U908 (N_908,N_827,N_876);
nor U909 (N_909,N_847,N_873);
nand U910 (N_910,N_886,N_851);
nand U911 (N_911,N_875,N_853);
and U912 (N_912,N_845,N_891);
or U913 (N_913,N_870,N_826);
and U914 (N_914,N_897,N_858);
nor U915 (N_915,N_893,N_895);
or U916 (N_916,N_833,N_879);
and U917 (N_917,N_830,N_890);
nand U918 (N_918,N_863,N_831);
nor U919 (N_919,N_857,N_856);
and U920 (N_920,N_855,N_832);
or U921 (N_921,N_877,N_872);
or U922 (N_922,N_878,N_880);
and U923 (N_923,N_862,N_828);
or U924 (N_924,N_871,N_852);
and U925 (N_925,N_840,N_834);
nand U926 (N_926,N_869,N_892);
and U927 (N_927,N_889,N_854);
or U928 (N_928,N_883,N_867);
and U929 (N_929,N_865,N_868);
nor U930 (N_930,N_887,N_861);
xor U931 (N_931,N_837,N_874);
nand U932 (N_932,N_866,N_850);
and U933 (N_933,N_885,N_881);
or U934 (N_934,N_839,N_842);
nand U935 (N_935,N_841,N_898);
nand U936 (N_936,N_849,N_888);
nor U937 (N_937,N_835,N_862);
nor U938 (N_938,N_863,N_871);
nor U939 (N_939,N_831,N_865);
and U940 (N_940,N_851,N_892);
nand U941 (N_941,N_878,N_842);
nand U942 (N_942,N_890,N_884);
or U943 (N_943,N_849,N_883);
and U944 (N_944,N_853,N_898);
or U945 (N_945,N_830,N_841);
or U946 (N_946,N_847,N_877);
and U947 (N_947,N_858,N_852);
and U948 (N_948,N_832,N_863);
or U949 (N_949,N_874,N_862);
or U950 (N_950,N_846,N_849);
nand U951 (N_951,N_851,N_867);
nand U952 (N_952,N_882,N_877);
and U953 (N_953,N_853,N_865);
nand U954 (N_954,N_831,N_853);
nand U955 (N_955,N_889,N_893);
xnor U956 (N_956,N_876,N_832);
and U957 (N_957,N_899,N_896);
nand U958 (N_958,N_887,N_874);
nand U959 (N_959,N_829,N_860);
nand U960 (N_960,N_848,N_871);
nand U961 (N_961,N_838,N_874);
or U962 (N_962,N_825,N_830);
nand U963 (N_963,N_879,N_877);
or U964 (N_964,N_894,N_876);
nor U965 (N_965,N_892,N_850);
nand U966 (N_966,N_860,N_897);
nor U967 (N_967,N_877,N_851);
or U968 (N_968,N_847,N_856);
and U969 (N_969,N_879,N_857);
xor U970 (N_970,N_842,N_864);
nand U971 (N_971,N_883,N_829);
and U972 (N_972,N_837,N_853);
nand U973 (N_973,N_886,N_870);
nor U974 (N_974,N_897,N_879);
and U975 (N_975,N_970,N_974);
nand U976 (N_976,N_960,N_912);
nand U977 (N_977,N_930,N_958);
and U978 (N_978,N_917,N_959);
nor U979 (N_979,N_916,N_921);
or U980 (N_980,N_910,N_940);
nor U981 (N_981,N_943,N_911);
nand U982 (N_982,N_939,N_957);
or U983 (N_983,N_938,N_901);
nand U984 (N_984,N_918,N_903);
and U985 (N_985,N_936,N_961);
or U986 (N_986,N_949,N_919);
or U987 (N_987,N_955,N_956);
nand U988 (N_988,N_929,N_966);
or U989 (N_989,N_933,N_923);
or U990 (N_990,N_972,N_934);
nand U991 (N_991,N_927,N_915);
or U992 (N_992,N_945,N_900);
xnor U993 (N_993,N_904,N_969);
nor U994 (N_994,N_909,N_964);
nand U995 (N_995,N_944,N_967);
or U996 (N_996,N_935,N_920);
nor U997 (N_997,N_953,N_926);
and U998 (N_998,N_907,N_973);
and U999 (N_999,N_925,N_913);
nand U1000 (N_1000,N_937,N_946);
nor U1001 (N_1001,N_950,N_914);
or U1002 (N_1002,N_931,N_908);
nand U1003 (N_1003,N_905,N_928);
nand U1004 (N_1004,N_968,N_963);
or U1005 (N_1005,N_922,N_906);
nor U1006 (N_1006,N_971,N_954);
or U1007 (N_1007,N_952,N_965);
or U1008 (N_1008,N_924,N_951);
xor U1009 (N_1009,N_947,N_962);
and U1010 (N_1010,N_932,N_902);
nand U1011 (N_1011,N_948,N_941);
nor U1012 (N_1012,N_942,N_949);
nor U1013 (N_1013,N_951,N_945);
nand U1014 (N_1014,N_932,N_911);
nand U1015 (N_1015,N_942,N_945);
nor U1016 (N_1016,N_950,N_924);
or U1017 (N_1017,N_954,N_909);
or U1018 (N_1018,N_965,N_958);
xnor U1019 (N_1019,N_963,N_902);
xnor U1020 (N_1020,N_952,N_932);
nor U1021 (N_1021,N_901,N_904);
and U1022 (N_1022,N_959,N_908);
nor U1023 (N_1023,N_919,N_935);
or U1024 (N_1024,N_968,N_970);
nor U1025 (N_1025,N_929,N_911);
nor U1026 (N_1026,N_918,N_974);
nor U1027 (N_1027,N_930,N_963);
or U1028 (N_1028,N_952,N_918);
nor U1029 (N_1029,N_953,N_969);
and U1030 (N_1030,N_934,N_964);
or U1031 (N_1031,N_901,N_958);
xnor U1032 (N_1032,N_937,N_908);
and U1033 (N_1033,N_935,N_903);
and U1034 (N_1034,N_955,N_930);
nand U1035 (N_1035,N_906,N_945);
nand U1036 (N_1036,N_954,N_923);
nand U1037 (N_1037,N_965,N_917);
or U1038 (N_1038,N_902,N_952);
and U1039 (N_1039,N_973,N_928);
nor U1040 (N_1040,N_915,N_974);
xor U1041 (N_1041,N_916,N_959);
nor U1042 (N_1042,N_930,N_918);
or U1043 (N_1043,N_957,N_959);
and U1044 (N_1044,N_927,N_930);
nor U1045 (N_1045,N_907,N_931);
or U1046 (N_1046,N_950,N_965);
or U1047 (N_1047,N_951,N_910);
nand U1048 (N_1048,N_968,N_958);
xor U1049 (N_1049,N_901,N_937);
nor U1050 (N_1050,N_1007,N_1025);
and U1051 (N_1051,N_992,N_1018);
nand U1052 (N_1052,N_989,N_994);
and U1053 (N_1053,N_1006,N_1032);
nand U1054 (N_1054,N_1043,N_1003);
nand U1055 (N_1055,N_1005,N_997);
xor U1056 (N_1056,N_980,N_1029);
and U1057 (N_1057,N_998,N_982);
nand U1058 (N_1058,N_1000,N_1024);
nor U1059 (N_1059,N_976,N_1047);
or U1060 (N_1060,N_983,N_1049);
nand U1061 (N_1061,N_1014,N_1040);
nor U1062 (N_1062,N_1033,N_1027);
nand U1063 (N_1063,N_975,N_979);
or U1064 (N_1064,N_1001,N_1026);
nand U1065 (N_1065,N_1039,N_1048);
nand U1066 (N_1066,N_1010,N_1021);
or U1067 (N_1067,N_1016,N_1020);
and U1068 (N_1068,N_987,N_1045);
xnor U1069 (N_1069,N_1004,N_1002);
and U1070 (N_1070,N_1012,N_986);
nand U1071 (N_1071,N_1008,N_978);
and U1072 (N_1072,N_977,N_993);
nand U1073 (N_1073,N_1023,N_990);
and U1074 (N_1074,N_988,N_1028);
or U1075 (N_1075,N_1038,N_1044);
and U1076 (N_1076,N_995,N_981);
and U1077 (N_1077,N_996,N_1041);
nand U1078 (N_1078,N_1037,N_1031);
or U1079 (N_1079,N_1017,N_984);
and U1080 (N_1080,N_1046,N_999);
nor U1081 (N_1081,N_1009,N_1019);
and U1082 (N_1082,N_1035,N_1042);
and U1083 (N_1083,N_1030,N_1011);
nand U1084 (N_1084,N_1015,N_991);
nand U1085 (N_1085,N_1022,N_1013);
or U1086 (N_1086,N_985,N_1036);
nand U1087 (N_1087,N_1034,N_988);
nand U1088 (N_1088,N_996,N_981);
nor U1089 (N_1089,N_1004,N_989);
nor U1090 (N_1090,N_1041,N_1032);
or U1091 (N_1091,N_996,N_1035);
nand U1092 (N_1092,N_1006,N_991);
or U1093 (N_1093,N_1012,N_1001);
or U1094 (N_1094,N_1047,N_1033);
and U1095 (N_1095,N_1044,N_1036);
nand U1096 (N_1096,N_1008,N_985);
xnor U1097 (N_1097,N_1015,N_987);
nand U1098 (N_1098,N_977,N_998);
and U1099 (N_1099,N_1026,N_1008);
and U1100 (N_1100,N_1048,N_1032);
nand U1101 (N_1101,N_980,N_1045);
nand U1102 (N_1102,N_989,N_984);
xnor U1103 (N_1103,N_1043,N_1021);
xnor U1104 (N_1104,N_988,N_994);
nor U1105 (N_1105,N_1042,N_1033);
or U1106 (N_1106,N_980,N_1007);
and U1107 (N_1107,N_1029,N_989);
nand U1108 (N_1108,N_1046,N_1027);
nor U1109 (N_1109,N_1011,N_1029);
or U1110 (N_1110,N_982,N_1023);
or U1111 (N_1111,N_981,N_1026);
nor U1112 (N_1112,N_999,N_976);
nor U1113 (N_1113,N_1040,N_1007);
and U1114 (N_1114,N_1043,N_996);
or U1115 (N_1115,N_1011,N_1017);
xnor U1116 (N_1116,N_1044,N_1046);
nor U1117 (N_1117,N_1046,N_1015);
nand U1118 (N_1118,N_1033,N_1046);
or U1119 (N_1119,N_1008,N_1036);
xnor U1120 (N_1120,N_990,N_1037);
and U1121 (N_1121,N_1036,N_1002);
or U1122 (N_1122,N_1046,N_979);
xor U1123 (N_1123,N_1016,N_1005);
and U1124 (N_1124,N_1042,N_1045);
xnor U1125 (N_1125,N_1095,N_1096);
nor U1126 (N_1126,N_1058,N_1076);
and U1127 (N_1127,N_1078,N_1097);
nand U1128 (N_1128,N_1052,N_1118);
xnor U1129 (N_1129,N_1074,N_1050);
or U1130 (N_1130,N_1094,N_1064);
and U1131 (N_1131,N_1086,N_1116);
nand U1132 (N_1132,N_1087,N_1108);
nor U1133 (N_1133,N_1112,N_1106);
and U1134 (N_1134,N_1120,N_1062);
or U1135 (N_1135,N_1059,N_1091);
or U1136 (N_1136,N_1079,N_1082);
nand U1137 (N_1137,N_1115,N_1107);
and U1138 (N_1138,N_1098,N_1089);
xnor U1139 (N_1139,N_1071,N_1123);
or U1140 (N_1140,N_1105,N_1119);
nand U1141 (N_1141,N_1075,N_1068);
and U1142 (N_1142,N_1104,N_1066);
and U1143 (N_1143,N_1109,N_1088);
nand U1144 (N_1144,N_1061,N_1051);
and U1145 (N_1145,N_1073,N_1080);
nor U1146 (N_1146,N_1111,N_1067);
or U1147 (N_1147,N_1085,N_1100);
or U1148 (N_1148,N_1077,N_1072);
xnor U1149 (N_1149,N_1084,N_1124);
or U1150 (N_1150,N_1093,N_1110);
and U1151 (N_1151,N_1099,N_1102);
and U1152 (N_1152,N_1069,N_1057);
and U1153 (N_1153,N_1056,N_1092);
nor U1154 (N_1154,N_1101,N_1060);
or U1155 (N_1155,N_1063,N_1083);
nand U1156 (N_1156,N_1122,N_1070);
or U1157 (N_1157,N_1065,N_1081);
or U1158 (N_1158,N_1121,N_1054);
nand U1159 (N_1159,N_1113,N_1103);
nand U1160 (N_1160,N_1055,N_1090);
nand U1161 (N_1161,N_1117,N_1053);
and U1162 (N_1162,N_1114,N_1090);
nor U1163 (N_1163,N_1088,N_1069);
or U1164 (N_1164,N_1051,N_1120);
and U1165 (N_1165,N_1109,N_1054);
and U1166 (N_1166,N_1118,N_1092);
nor U1167 (N_1167,N_1053,N_1096);
xor U1168 (N_1168,N_1055,N_1109);
and U1169 (N_1169,N_1075,N_1113);
nor U1170 (N_1170,N_1111,N_1097);
or U1171 (N_1171,N_1069,N_1050);
nand U1172 (N_1172,N_1091,N_1056);
nor U1173 (N_1173,N_1072,N_1074);
and U1174 (N_1174,N_1097,N_1064);
nor U1175 (N_1175,N_1050,N_1079);
nand U1176 (N_1176,N_1102,N_1052);
and U1177 (N_1177,N_1091,N_1077);
or U1178 (N_1178,N_1084,N_1082);
nor U1179 (N_1179,N_1080,N_1076);
or U1180 (N_1180,N_1072,N_1084);
nor U1181 (N_1181,N_1106,N_1114);
nand U1182 (N_1182,N_1050,N_1117);
and U1183 (N_1183,N_1096,N_1112);
nand U1184 (N_1184,N_1121,N_1104);
nand U1185 (N_1185,N_1123,N_1056);
or U1186 (N_1186,N_1065,N_1067);
nor U1187 (N_1187,N_1050,N_1104);
nor U1188 (N_1188,N_1123,N_1124);
or U1189 (N_1189,N_1087,N_1124);
or U1190 (N_1190,N_1122,N_1072);
or U1191 (N_1191,N_1085,N_1072);
and U1192 (N_1192,N_1063,N_1090);
nand U1193 (N_1193,N_1093,N_1097);
xor U1194 (N_1194,N_1099,N_1079);
and U1195 (N_1195,N_1064,N_1091);
and U1196 (N_1196,N_1120,N_1096);
and U1197 (N_1197,N_1073,N_1051);
nor U1198 (N_1198,N_1104,N_1116);
xor U1199 (N_1199,N_1070,N_1077);
nand U1200 (N_1200,N_1146,N_1150);
nand U1201 (N_1201,N_1192,N_1135);
nor U1202 (N_1202,N_1125,N_1174);
or U1203 (N_1203,N_1189,N_1129);
nor U1204 (N_1204,N_1173,N_1130);
and U1205 (N_1205,N_1158,N_1191);
or U1206 (N_1206,N_1142,N_1127);
and U1207 (N_1207,N_1166,N_1139);
or U1208 (N_1208,N_1134,N_1196);
nor U1209 (N_1209,N_1137,N_1143);
and U1210 (N_1210,N_1177,N_1136);
nand U1211 (N_1211,N_1179,N_1147);
and U1212 (N_1212,N_1155,N_1167);
nor U1213 (N_1213,N_1128,N_1140);
and U1214 (N_1214,N_1156,N_1170);
or U1215 (N_1215,N_1153,N_1132);
nand U1216 (N_1216,N_1171,N_1190);
nand U1217 (N_1217,N_1160,N_1141);
and U1218 (N_1218,N_1178,N_1185);
xor U1219 (N_1219,N_1194,N_1154);
and U1220 (N_1220,N_1186,N_1161);
or U1221 (N_1221,N_1133,N_1188);
and U1222 (N_1222,N_1131,N_1164);
nor U1223 (N_1223,N_1168,N_1152);
nor U1224 (N_1224,N_1145,N_1165);
nor U1225 (N_1225,N_1199,N_1187);
or U1226 (N_1226,N_1126,N_1175);
nor U1227 (N_1227,N_1148,N_1151);
nor U1228 (N_1228,N_1198,N_1183);
or U1229 (N_1229,N_1172,N_1176);
nand U1230 (N_1230,N_1138,N_1184);
and U1231 (N_1231,N_1157,N_1159);
nand U1232 (N_1232,N_1195,N_1163);
or U1233 (N_1233,N_1181,N_1197);
and U1234 (N_1234,N_1180,N_1149);
nor U1235 (N_1235,N_1162,N_1144);
nand U1236 (N_1236,N_1182,N_1193);
nand U1237 (N_1237,N_1169,N_1166);
and U1238 (N_1238,N_1183,N_1138);
and U1239 (N_1239,N_1136,N_1134);
nor U1240 (N_1240,N_1180,N_1125);
or U1241 (N_1241,N_1195,N_1128);
nand U1242 (N_1242,N_1140,N_1150);
nand U1243 (N_1243,N_1198,N_1188);
nand U1244 (N_1244,N_1179,N_1195);
or U1245 (N_1245,N_1183,N_1156);
or U1246 (N_1246,N_1185,N_1183);
nand U1247 (N_1247,N_1194,N_1184);
or U1248 (N_1248,N_1193,N_1187);
nand U1249 (N_1249,N_1147,N_1185);
nor U1250 (N_1250,N_1192,N_1136);
nand U1251 (N_1251,N_1142,N_1172);
and U1252 (N_1252,N_1151,N_1181);
and U1253 (N_1253,N_1183,N_1187);
and U1254 (N_1254,N_1154,N_1187);
nand U1255 (N_1255,N_1153,N_1145);
xnor U1256 (N_1256,N_1132,N_1187);
nand U1257 (N_1257,N_1171,N_1154);
nand U1258 (N_1258,N_1138,N_1161);
xor U1259 (N_1259,N_1138,N_1186);
or U1260 (N_1260,N_1180,N_1179);
nor U1261 (N_1261,N_1181,N_1196);
or U1262 (N_1262,N_1131,N_1144);
and U1263 (N_1263,N_1138,N_1162);
nor U1264 (N_1264,N_1155,N_1143);
and U1265 (N_1265,N_1164,N_1184);
and U1266 (N_1266,N_1184,N_1157);
and U1267 (N_1267,N_1160,N_1163);
nand U1268 (N_1268,N_1189,N_1157);
nand U1269 (N_1269,N_1167,N_1196);
or U1270 (N_1270,N_1143,N_1125);
xnor U1271 (N_1271,N_1190,N_1168);
and U1272 (N_1272,N_1175,N_1125);
or U1273 (N_1273,N_1169,N_1134);
nor U1274 (N_1274,N_1148,N_1174);
xnor U1275 (N_1275,N_1212,N_1260);
nand U1276 (N_1276,N_1221,N_1270);
nor U1277 (N_1277,N_1257,N_1248);
nor U1278 (N_1278,N_1269,N_1255);
and U1279 (N_1279,N_1252,N_1208);
nand U1280 (N_1280,N_1215,N_1202);
or U1281 (N_1281,N_1216,N_1239);
nand U1282 (N_1282,N_1220,N_1271);
and U1283 (N_1283,N_1218,N_1235);
nand U1284 (N_1284,N_1272,N_1200);
xor U1285 (N_1285,N_1263,N_1224);
xor U1286 (N_1286,N_1228,N_1227);
and U1287 (N_1287,N_1249,N_1201);
nand U1288 (N_1288,N_1274,N_1259);
xor U1289 (N_1289,N_1223,N_1240);
nand U1290 (N_1290,N_1254,N_1217);
nor U1291 (N_1291,N_1251,N_1262);
nor U1292 (N_1292,N_1245,N_1226);
nor U1293 (N_1293,N_1231,N_1247);
nand U1294 (N_1294,N_1211,N_1265);
nor U1295 (N_1295,N_1213,N_1203);
nor U1296 (N_1296,N_1250,N_1266);
and U1297 (N_1297,N_1205,N_1233);
or U1298 (N_1298,N_1258,N_1206);
or U1299 (N_1299,N_1230,N_1256);
nor U1300 (N_1300,N_1219,N_1210);
and U1301 (N_1301,N_1268,N_1225);
and U1302 (N_1302,N_1234,N_1214);
or U1303 (N_1303,N_1207,N_1209);
and U1304 (N_1304,N_1204,N_1244);
and U1305 (N_1305,N_1236,N_1261);
nor U1306 (N_1306,N_1232,N_1273);
xor U1307 (N_1307,N_1264,N_1237);
xnor U1308 (N_1308,N_1246,N_1253);
xnor U1309 (N_1309,N_1241,N_1238);
or U1310 (N_1310,N_1267,N_1222);
nor U1311 (N_1311,N_1242,N_1243);
nor U1312 (N_1312,N_1229,N_1240);
xnor U1313 (N_1313,N_1247,N_1211);
or U1314 (N_1314,N_1220,N_1248);
nand U1315 (N_1315,N_1224,N_1249);
or U1316 (N_1316,N_1204,N_1211);
xnor U1317 (N_1317,N_1209,N_1228);
nor U1318 (N_1318,N_1226,N_1235);
and U1319 (N_1319,N_1227,N_1232);
nand U1320 (N_1320,N_1265,N_1256);
nand U1321 (N_1321,N_1237,N_1205);
or U1322 (N_1322,N_1245,N_1241);
or U1323 (N_1323,N_1201,N_1216);
and U1324 (N_1324,N_1247,N_1210);
nand U1325 (N_1325,N_1265,N_1220);
or U1326 (N_1326,N_1259,N_1266);
or U1327 (N_1327,N_1251,N_1256);
nor U1328 (N_1328,N_1226,N_1249);
or U1329 (N_1329,N_1273,N_1215);
nand U1330 (N_1330,N_1230,N_1249);
or U1331 (N_1331,N_1231,N_1236);
xnor U1332 (N_1332,N_1210,N_1270);
and U1333 (N_1333,N_1233,N_1273);
and U1334 (N_1334,N_1237,N_1274);
nor U1335 (N_1335,N_1246,N_1245);
nor U1336 (N_1336,N_1227,N_1207);
and U1337 (N_1337,N_1213,N_1227);
or U1338 (N_1338,N_1229,N_1256);
nand U1339 (N_1339,N_1265,N_1248);
nand U1340 (N_1340,N_1242,N_1211);
or U1341 (N_1341,N_1240,N_1274);
nor U1342 (N_1342,N_1235,N_1214);
or U1343 (N_1343,N_1202,N_1213);
or U1344 (N_1344,N_1203,N_1256);
xor U1345 (N_1345,N_1221,N_1225);
and U1346 (N_1346,N_1224,N_1223);
or U1347 (N_1347,N_1239,N_1202);
xor U1348 (N_1348,N_1224,N_1209);
xnor U1349 (N_1349,N_1240,N_1247);
nor U1350 (N_1350,N_1341,N_1289);
and U1351 (N_1351,N_1306,N_1279);
and U1352 (N_1352,N_1311,N_1290);
nand U1353 (N_1353,N_1280,N_1283);
and U1354 (N_1354,N_1313,N_1320);
nand U1355 (N_1355,N_1310,N_1319);
nor U1356 (N_1356,N_1284,N_1348);
xor U1357 (N_1357,N_1305,N_1322);
nor U1358 (N_1358,N_1349,N_1288);
nor U1359 (N_1359,N_1299,N_1278);
and U1360 (N_1360,N_1275,N_1314);
or U1361 (N_1361,N_1287,N_1316);
or U1362 (N_1362,N_1293,N_1345);
or U1363 (N_1363,N_1342,N_1282);
nand U1364 (N_1364,N_1315,N_1325);
and U1365 (N_1365,N_1309,N_1302);
nand U1366 (N_1366,N_1286,N_1336);
and U1367 (N_1367,N_1335,N_1327);
or U1368 (N_1368,N_1347,N_1332);
nand U1369 (N_1369,N_1329,N_1312);
xor U1370 (N_1370,N_1308,N_1296);
nand U1371 (N_1371,N_1331,N_1334);
or U1372 (N_1372,N_1291,N_1292);
or U1373 (N_1373,N_1276,N_1324);
or U1374 (N_1374,N_1298,N_1300);
nand U1375 (N_1375,N_1346,N_1343);
and U1376 (N_1376,N_1328,N_1307);
nand U1377 (N_1377,N_1330,N_1318);
nor U1378 (N_1378,N_1321,N_1301);
nor U1379 (N_1379,N_1326,N_1303);
and U1380 (N_1380,N_1285,N_1297);
xnor U1381 (N_1381,N_1281,N_1295);
xnor U1382 (N_1382,N_1338,N_1277);
or U1383 (N_1383,N_1317,N_1344);
or U1384 (N_1384,N_1294,N_1304);
or U1385 (N_1385,N_1337,N_1340);
nor U1386 (N_1386,N_1333,N_1323);
and U1387 (N_1387,N_1339,N_1327);
or U1388 (N_1388,N_1280,N_1340);
and U1389 (N_1389,N_1290,N_1286);
or U1390 (N_1390,N_1279,N_1335);
nand U1391 (N_1391,N_1346,N_1288);
or U1392 (N_1392,N_1343,N_1302);
or U1393 (N_1393,N_1303,N_1310);
and U1394 (N_1394,N_1304,N_1324);
and U1395 (N_1395,N_1316,N_1323);
xor U1396 (N_1396,N_1321,N_1317);
and U1397 (N_1397,N_1327,N_1346);
or U1398 (N_1398,N_1336,N_1292);
nand U1399 (N_1399,N_1291,N_1304);
nand U1400 (N_1400,N_1319,N_1302);
and U1401 (N_1401,N_1317,N_1338);
nor U1402 (N_1402,N_1329,N_1295);
and U1403 (N_1403,N_1276,N_1343);
xnor U1404 (N_1404,N_1280,N_1315);
nor U1405 (N_1405,N_1299,N_1337);
nor U1406 (N_1406,N_1331,N_1335);
nor U1407 (N_1407,N_1278,N_1320);
and U1408 (N_1408,N_1345,N_1288);
or U1409 (N_1409,N_1331,N_1288);
and U1410 (N_1410,N_1286,N_1289);
or U1411 (N_1411,N_1310,N_1343);
or U1412 (N_1412,N_1275,N_1294);
nand U1413 (N_1413,N_1292,N_1307);
or U1414 (N_1414,N_1312,N_1314);
and U1415 (N_1415,N_1328,N_1337);
xor U1416 (N_1416,N_1314,N_1349);
or U1417 (N_1417,N_1277,N_1298);
or U1418 (N_1418,N_1308,N_1288);
or U1419 (N_1419,N_1287,N_1293);
xor U1420 (N_1420,N_1288,N_1280);
nand U1421 (N_1421,N_1330,N_1296);
or U1422 (N_1422,N_1331,N_1345);
and U1423 (N_1423,N_1320,N_1279);
or U1424 (N_1424,N_1310,N_1295);
or U1425 (N_1425,N_1406,N_1404);
nand U1426 (N_1426,N_1358,N_1353);
xor U1427 (N_1427,N_1384,N_1395);
nand U1428 (N_1428,N_1391,N_1381);
xnor U1429 (N_1429,N_1397,N_1371);
or U1430 (N_1430,N_1403,N_1377);
xor U1431 (N_1431,N_1376,N_1411);
or U1432 (N_1432,N_1415,N_1412);
xor U1433 (N_1433,N_1399,N_1402);
nor U1434 (N_1434,N_1408,N_1378);
or U1435 (N_1435,N_1416,N_1385);
or U1436 (N_1436,N_1387,N_1356);
nor U1437 (N_1437,N_1405,N_1424);
nor U1438 (N_1438,N_1394,N_1365);
xor U1439 (N_1439,N_1392,N_1360);
nand U1440 (N_1440,N_1350,N_1374);
or U1441 (N_1441,N_1357,N_1369);
and U1442 (N_1442,N_1355,N_1409);
nand U1443 (N_1443,N_1361,N_1373);
or U1444 (N_1444,N_1421,N_1368);
nand U1445 (N_1445,N_1422,N_1401);
nor U1446 (N_1446,N_1364,N_1418);
nor U1447 (N_1447,N_1417,N_1380);
nand U1448 (N_1448,N_1352,N_1390);
nand U1449 (N_1449,N_1423,N_1379);
and U1450 (N_1450,N_1388,N_1372);
or U1451 (N_1451,N_1389,N_1398);
and U1452 (N_1452,N_1351,N_1413);
or U1453 (N_1453,N_1359,N_1383);
xor U1454 (N_1454,N_1363,N_1354);
nand U1455 (N_1455,N_1396,N_1420);
and U1456 (N_1456,N_1410,N_1367);
nor U1457 (N_1457,N_1419,N_1386);
xnor U1458 (N_1458,N_1375,N_1414);
nand U1459 (N_1459,N_1400,N_1366);
nor U1460 (N_1460,N_1407,N_1362);
nor U1461 (N_1461,N_1370,N_1393);
nor U1462 (N_1462,N_1382,N_1389);
or U1463 (N_1463,N_1422,N_1370);
nor U1464 (N_1464,N_1415,N_1353);
and U1465 (N_1465,N_1423,N_1400);
nand U1466 (N_1466,N_1413,N_1368);
nand U1467 (N_1467,N_1387,N_1409);
and U1468 (N_1468,N_1389,N_1387);
and U1469 (N_1469,N_1358,N_1393);
nor U1470 (N_1470,N_1417,N_1419);
nand U1471 (N_1471,N_1391,N_1379);
or U1472 (N_1472,N_1401,N_1417);
xor U1473 (N_1473,N_1357,N_1402);
and U1474 (N_1474,N_1356,N_1354);
or U1475 (N_1475,N_1362,N_1357);
and U1476 (N_1476,N_1393,N_1373);
nand U1477 (N_1477,N_1413,N_1385);
or U1478 (N_1478,N_1387,N_1398);
nor U1479 (N_1479,N_1402,N_1373);
or U1480 (N_1480,N_1412,N_1354);
nor U1481 (N_1481,N_1396,N_1406);
xnor U1482 (N_1482,N_1420,N_1358);
and U1483 (N_1483,N_1374,N_1411);
nor U1484 (N_1484,N_1357,N_1419);
nor U1485 (N_1485,N_1387,N_1370);
or U1486 (N_1486,N_1367,N_1370);
and U1487 (N_1487,N_1419,N_1406);
nand U1488 (N_1488,N_1398,N_1355);
or U1489 (N_1489,N_1422,N_1352);
or U1490 (N_1490,N_1392,N_1380);
or U1491 (N_1491,N_1400,N_1367);
or U1492 (N_1492,N_1356,N_1371);
nor U1493 (N_1493,N_1413,N_1367);
nor U1494 (N_1494,N_1393,N_1364);
nand U1495 (N_1495,N_1373,N_1372);
nand U1496 (N_1496,N_1388,N_1400);
xnor U1497 (N_1497,N_1374,N_1418);
or U1498 (N_1498,N_1410,N_1372);
and U1499 (N_1499,N_1363,N_1352);
and U1500 (N_1500,N_1446,N_1479);
xnor U1501 (N_1501,N_1470,N_1482);
nor U1502 (N_1502,N_1476,N_1471);
and U1503 (N_1503,N_1468,N_1495);
and U1504 (N_1504,N_1463,N_1447);
nor U1505 (N_1505,N_1459,N_1445);
xnor U1506 (N_1506,N_1449,N_1480);
or U1507 (N_1507,N_1430,N_1475);
and U1508 (N_1508,N_1456,N_1436);
xor U1509 (N_1509,N_1438,N_1461);
nor U1510 (N_1510,N_1481,N_1457);
or U1511 (N_1511,N_1465,N_1490);
nor U1512 (N_1512,N_1444,N_1473);
and U1513 (N_1513,N_1434,N_1498);
xnor U1514 (N_1514,N_1452,N_1492);
and U1515 (N_1515,N_1497,N_1441);
nand U1516 (N_1516,N_1450,N_1455);
nand U1517 (N_1517,N_1426,N_1433);
nor U1518 (N_1518,N_1477,N_1484);
nand U1519 (N_1519,N_1486,N_1453);
nand U1520 (N_1520,N_1462,N_1483);
nand U1521 (N_1521,N_1467,N_1496);
xnor U1522 (N_1522,N_1466,N_1442);
nor U1523 (N_1523,N_1439,N_1448);
xor U1524 (N_1524,N_1489,N_1440);
or U1525 (N_1525,N_1472,N_1431);
nor U1526 (N_1526,N_1494,N_1451);
nor U1527 (N_1527,N_1429,N_1485);
and U1528 (N_1528,N_1427,N_1488);
and U1529 (N_1529,N_1464,N_1432);
nor U1530 (N_1530,N_1474,N_1437);
or U1531 (N_1531,N_1487,N_1499);
nor U1532 (N_1532,N_1458,N_1478);
xor U1533 (N_1533,N_1493,N_1443);
nor U1534 (N_1534,N_1428,N_1435);
or U1535 (N_1535,N_1425,N_1491);
nand U1536 (N_1536,N_1469,N_1460);
nand U1537 (N_1537,N_1454,N_1432);
and U1538 (N_1538,N_1426,N_1453);
xor U1539 (N_1539,N_1427,N_1440);
nand U1540 (N_1540,N_1476,N_1426);
xnor U1541 (N_1541,N_1463,N_1462);
nor U1542 (N_1542,N_1427,N_1454);
and U1543 (N_1543,N_1482,N_1457);
or U1544 (N_1544,N_1439,N_1484);
xor U1545 (N_1545,N_1456,N_1484);
nand U1546 (N_1546,N_1480,N_1491);
xnor U1547 (N_1547,N_1439,N_1460);
or U1548 (N_1548,N_1458,N_1459);
or U1549 (N_1549,N_1426,N_1434);
or U1550 (N_1550,N_1466,N_1495);
nor U1551 (N_1551,N_1455,N_1499);
and U1552 (N_1552,N_1437,N_1489);
and U1553 (N_1553,N_1471,N_1499);
and U1554 (N_1554,N_1441,N_1462);
or U1555 (N_1555,N_1470,N_1437);
nand U1556 (N_1556,N_1428,N_1492);
nor U1557 (N_1557,N_1471,N_1438);
nand U1558 (N_1558,N_1480,N_1442);
xnor U1559 (N_1559,N_1469,N_1451);
nor U1560 (N_1560,N_1493,N_1483);
or U1561 (N_1561,N_1458,N_1471);
xnor U1562 (N_1562,N_1450,N_1438);
nand U1563 (N_1563,N_1433,N_1438);
nand U1564 (N_1564,N_1487,N_1432);
nand U1565 (N_1565,N_1477,N_1499);
and U1566 (N_1566,N_1450,N_1474);
and U1567 (N_1567,N_1485,N_1434);
and U1568 (N_1568,N_1449,N_1456);
and U1569 (N_1569,N_1463,N_1457);
nand U1570 (N_1570,N_1429,N_1491);
nor U1571 (N_1571,N_1468,N_1473);
nor U1572 (N_1572,N_1495,N_1442);
xor U1573 (N_1573,N_1461,N_1427);
and U1574 (N_1574,N_1456,N_1442);
and U1575 (N_1575,N_1528,N_1547);
nor U1576 (N_1576,N_1540,N_1574);
nand U1577 (N_1577,N_1541,N_1510);
nand U1578 (N_1578,N_1504,N_1572);
nand U1579 (N_1579,N_1567,N_1535);
and U1580 (N_1580,N_1551,N_1502);
xor U1581 (N_1581,N_1503,N_1518);
nor U1582 (N_1582,N_1519,N_1532);
or U1583 (N_1583,N_1554,N_1530);
nand U1584 (N_1584,N_1573,N_1569);
and U1585 (N_1585,N_1500,N_1566);
nor U1586 (N_1586,N_1539,N_1542);
nor U1587 (N_1587,N_1556,N_1522);
nand U1588 (N_1588,N_1537,N_1524);
and U1589 (N_1589,N_1513,N_1545);
nand U1590 (N_1590,N_1546,N_1516);
and U1591 (N_1591,N_1562,N_1552);
and U1592 (N_1592,N_1550,N_1520);
nor U1593 (N_1593,N_1544,N_1525);
nor U1594 (N_1594,N_1501,N_1559);
and U1595 (N_1595,N_1505,N_1507);
nor U1596 (N_1596,N_1536,N_1509);
and U1597 (N_1597,N_1548,N_1538);
nor U1598 (N_1598,N_1564,N_1571);
nor U1599 (N_1599,N_1531,N_1534);
and U1600 (N_1600,N_1527,N_1561);
and U1601 (N_1601,N_1529,N_1506);
nor U1602 (N_1602,N_1515,N_1526);
xor U1603 (N_1603,N_1560,N_1517);
or U1604 (N_1604,N_1511,N_1512);
or U1605 (N_1605,N_1543,N_1514);
or U1606 (N_1606,N_1508,N_1555);
or U1607 (N_1607,N_1521,N_1568);
and U1608 (N_1608,N_1565,N_1563);
or U1609 (N_1609,N_1570,N_1558);
xor U1610 (N_1610,N_1533,N_1557);
nand U1611 (N_1611,N_1553,N_1549);
xnor U1612 (N_1612,N_1523,N_1551);
nor U1613 (N_1613,N_1528,N_1556);
nor U1614 (N_1614,N_1564,N_1500);
and U1615 (N_1615,N_1525,N_1563);
nor U1616 (N_1616,N_1539,N_1517);
and U1617 (N_1617,N_1530,N_1533);
xnor U1618 (N_1618,N_1569,N_1524);
nor U1619 (N_1619,N_1501,N_1535);
nand U1620 (N_1620,N_1564,N_1517);
or U1621 (N_1621,N_1569,N_1559);
or U1622 (N_1622,N_1526,N_1542);
nand U1623 (N_1623,N_1547,N_1553);
or U1624 (N_1624,N_1551,N_1528);
or U1625 (N_1625,N_1540,N_1547);
xnor U1626 (N_1626,N_1538,N_1511);
nand U1627 (N_1627,N_1561,N_1504);
nand U1628 (N_1628,N_1519,N_1551);
and U1629 (N_1629,N_1569,N_1547);
and U1630 (N_1630,N_1539,N_1515);
and U1631 (N_1631,N_1541,N_1529);
nand U1632 (N_1632,N_1560,N_1547);
nand U1633 (N_1633,N_1529,N_1551);
nand U1634 (N_1634,N_1535,N_1528);
nand U1635 (N_1635,N_1501,N_1539);
nor U1636 (N_1636,N_1528,N_1557);
nor U1637 (N_1637,N_1505,N_1510);
and U1638 (N_1638,N_1524,N_1530);
nand U1639 (N_1639,N_1508,N_1547);
or U1640 (N_1640,N_1549,N_1545);
xnor U1641 (N_1641,N_1513,N_1556);
and U1642 (N_1642,N_1554,N_1522);
xor U1643 (N_1643,N_1552,N_1527);
nand U1644 (N_1644,N_1530,N_1546);
or U1645 (N_1645,N_1523,N_1501);
and U1646 (N_1646,N_1529,N_1549);
or U1647 (N_1647,N_1503,N_1513);
and U1648 (N_1648,N_1568,N_1500);
nand U1649 (N_1649,N_1572,N_1518);
xor U1650 (N_1650,N_1606,N_1585);
nand U1651 (N_1651,N_1611,N_1634);
and U1652 (N_1652,N_1642,N_1618);
or U1653 (N_1653,N_1591,N_1590);
and U1654 (N_1654,N_1605,N_1632);
and U1655 (N_1655,N_1646,N_1616);
or U1656 (N_1656,N_1622,N_1588);
nand U1657 (N_1657,N_1625,N_1578);
and U1658 (N_1658,N_1579,N_1582);
nor U1659 (N_1659,N_1589,N_1630);
nand U1660 (N_1660,N_1640,N_1636);
nor U1661 (N_1661,N_1626,N_1584);
and U1662 (N_1662,N_1592,N_1601);
or U1663 (N_1663,N_1598,N_1649);
and U1664 (N_1664,N_1599,N_1628);
nand U1665 (N_1665,N_1608,N_1575);
and U1666 (N_1666,N_1587,N_1638);
and U1667 (N_1667,N_1619,N_1648);
and U1668 (N_1668,N_1594,N_1593);
xor U1669 (N_1669,N_1580,N_1610);
nor U1670 (N_1670,N_1629,N_1577);
nand U1671 (N_1671,N_1612,N_1607);
nor U1672 (N_1672,N_1623,N_1639);
or U1673 (N_1673,N_1620,N_1604);
nor U1674 (N_1674,N_1633,N_1576);
and U1675 (N_1675,N_1627,N_1615);
nand U1676 (N_1676,N_1609,N_1613);
nand U1677 (N_1677,N_1643,N_1595);
or U1678 (N_1678,N_1600,N_1644);
nand U1679 (N_1679,N_1637,N_1602);
and U1680 (N_1680,N_1614,N_1635);
nor U1681 (N_1681,N_1581,N_1597);
xnor U1682 (N_1682,N_1583,N_1621);
or U1683 (N_1683,N_1586,N_1641);
nand U1684 (N_1684,N_1617,N_1603);
or U1685 (N_1685,N_1631,N_1647);
xor U1686 (N_1686,N_1624,N_1645);
or U1687 (N_1687,N_1596,N_1646);
nand U1688 (N_1688,N_1644,N_1592);
nor U1689 (N_1689,N_1615,N_1622);
and U1690 (N_1690,N_1617,N_1627);
nor U1691 (N_1691,N_1648,N_1585);
or U1692 (N_1692,N_1616,N_1648);
nand U1693 (N_1693,N_1648,N_1586);
nand U1694 (N_1694,N_1609,N_1633);
or U1695 (N_1695,N_1607,N_1604);
xor U1696 (N_1696,N_1628,N_1638);
nor U1697 (N_1697,N_1622,N_1616);
xor U1698 (N_1698,N_1614,N_1596);
and U1699 (N_1699,N_1643,N_1627);
and U1700 (N_1700,N_1589,N_1600);
nand U1701 (N_1701,N_1611,N_1609);
xor U1702 (N_1702,N_1612,N_1622);
nand U1703 (N_1703,N_1599,N_1646);
and U1704 (N_1704,N_1575,N_1597);
nand U1705 (N_1705,N_1576,N_1612);
or U1706 (N_1706,N_1601,N_1610);
and U1707 (N_1707,N_1625,N_1605);
nand U1708 (N_1708,N_1639,N_1593);
and U1709 (N_1709,N_1598,N_1618);
or U1710 (N_1710,N_1614,N_1581);
and U1711 (N_1711,N_1583,N_1602);
nand U1712 (N_1712,N_1610,N_1619);
and U1713 (N_1713,N_1634,N_1582);
and U1714 (N_1714,N_1637,N_1607);
and U1715 (N_1715,N_1588,N_1589);
xor U1716 (N_1716,N_1638,N_1609);
or U1717 (N_1717,N_1628,N_1575);
nand U1718 (N_1718,N_1627,N_1609);
nand U1719 (N_1719,N_1618,N_1600);
nand U1720 (N_1720,N_1599,N_1644);
nand U1721 (N_1721,N_1597,N_1617);
nand U1722 (N_1722,N_1590,N_1579);
nand U1723 (N_1723,N_1591,N_1621);
nand U1724 (N_1724,N_1596,N_1631);
or U1725 (N_1725,N_1675,N_1659);
or U1726 (N_1726,N_1712,N_1670);
nor U1727 (N_1727,N_1651,N_1702);
or U1728 (N_1728,N_1706,N_1703);
or U1729 (N_1729,N_1690,N_1698);
nor U1730 (N_1730,N_1653,N_1660);
nor U1731 (N_1731,N_1694,N_1701);
nand U1732 (N_1732,N_1685,N_1707);
nand U1733 (N_1733,N_1674,N_1665);
or U1734 (N_1734,N_1663,N_1713);
and U1735 (N_1735,N_1655,N_1709);
xnor U1736 (N_1736,N_1723,N_1719);
nand U1737 (N_1737,N_1688,N_1672);
nor U1738 (N_1738,N_1699,N_1724);
and U1739 (N_1739,N_1692,N_1661);
nand U1740 (N_1740,N_1697,N_1679);
nor U1741 (N_1741,N_1710,N_1652);
and U1742 (N_1742,N_1664,N_1716);
nand U1743 (N_1743,N_1704,N_1714);
or U1744 (N_1744,N_1693,N_1718);
nand U1745 (N_1745,N_1715,N_1691);
and U1746 (N_1746,N_1717,N_1700);
and U1747 (N_1747,N_1667,N_1683);
nor U1748 (N_1748,N_1671,N_1680);
nor U1749 (N_1749,N_1654,N_1705);
nor U1750 (N_1750,N_1708,N_1696);
xnor U1751 (N_1751,N_1695,N_1662);
and U1752 (N_1752,N_1682,N_1686);
and U1753 (N_1753,N_1678,N_1650);
nor U1754 (N_1754,N_1720,N_1687);
and U1755 (N_1755,N_1677,N_1722);
xnor U1756 (N_1756,N_1721,N_1657);
xnor U1757 (N_1757,N_1676,N_1669);
or U1758 (N_1758,N_1711,N_1656);
and U1759 (N_1759,N_1658,N_1668);
nor U1760 (N_1760,N_1681,N_1666);
or U1761 (N_1761,N_1684,N_1673);
or U1762 (N_1762,N_1689,N_1688);
or U1763 (N_1763,N_1722,N_1718);
nand U1764 (N_1764,N_1671,N_1653);
or U1765 (N_1765,N_1656,N_1651);
nor U1766 (N_1766,N_1715,N_1684);
or U1767 (N_1767,N_1675,N_1672);
nand U1768 (N_1768,N_1670,N_1681);
or U1769 (N_1769,N_1710,N_1694);
nand U1770 (N_1770,N_1676,N_1662);
nand U1771 (N_1771,N_1700,N_1716);
nor U1772 (N_1772,N_1703,N_1689);
or U1773 (N_1773,N_1653,N_1698);
nand U1774 (N_1774,N_1698,N_1651);
and U1775 (N_1775,N_1723,N_1671);
xor U1776 (N_1776,N_1714,N_1692);
or U1777 (N_1777,N_1672,N_1679);
nor U1778 (N_1778,N_1718,N_1720);
and U1779 (N_1779,N_1655,N_1712);
nor U1780 (N_1780,N_1659,N_1707);
nand U1781 (N_1781,N_1713,N_1697);
nand U1782 (N_1782,N_1690,N_1724);
xor U1783 (N_1783,N_1675,N_1701);
nor U1784 (N_1784,N_1713,N_1710);
or U1785 (N_1785,N_1672,N_1669);
and U1786 (N_1786,N_1665,N_1693);
or U1787 (N_1787,N_1715,N_1670);
and U1788 (N_1788,N_1650,N_1669);
or U1789 (N_1789,N_1720,N_1675);
nor U1790 (N_1790,N_1684,N_1696);
and U1791 (N_1791,N_1700,N_1708);
nand U1792 (N_1792,N_1658,N_1650);
and U1793 (N_1793,N_1707,N_1658);
nand U1794 (N_1794,N_1674,N_1720);
xnor U1795 (N_1795,N_1710,N_1708);
nand U1796 (N_1796,N_1697,N_1696);
and U1797 (N_1797,N_1708,N_1718);
or U1798 (N_1798,N_1674,N_1706);
nand U1799 (N_1799,N_1664,N_1668);
nand U1800 (N_1800,N_1777,N_1758);
nand U1801 (N_1801,N_1752,N_1734);
nand U1802 (N_1802,N_1779,N_1765);
or U1803 (N_1803,N_1728,N_1725);
nand U1804 (N_1804,N_1749,N_1726);
nor U1805 (N_1805,N_1743,N_1769);
and U1806 (N_1806,N_1763,N_1787);
and U1807 (N_1807,N_1762,N_1798);
and U1808 (N_1808,N_1748,N_1740);
nor U1809 (N_1809,N_1793,N_1754);
nor U1810 (N_1810,N_1785,N_1775);
or U1811 (N_1811,N_1786,N_1771);
xor U1812 (N_1812,N_1736,N_1790);
xnor U1813 (N_1813,N_1729,N_1750);
nor U1814 (N_1814,N_1746,N_1733);
nand U1815 (N_1815,N_1772,N_1796);
or U1816 (N_1816,N_1760,N_1739);
xor U1817 (N_1817,N_1757,N_1783);
nand U1818 (N_1818,N_1791,N_1747);
nor U1819 (N_1819,N_1745,N_1731);
or U1820 (N_1820,N_1797,N_1784);
nor U1821 (N_1821,N_1756,N_1737);
or U1822 (N_1822,N_1761,N_1778);
or U1823 (N_1823,N_1792,N_1744);
xor U1824 (N_1824,N_1753,N_1730);
nor U1825 (N_1825,N_1773,N_1782);
nand U1826 (N_1826,N_1751,N_1741);
xor U1827 (N_1827,N_1768,N_1767);
and U1828 (N_1828,N_1742,N_1794);
and U1829 (N_1829,N_1781,N_1735);
nor U1830 (N_1830,N_1764,N_1770);
and U1831 (N_1831,N_1774,N_1795);
and U1832 (N_1832,N_1766,N_1780);
or U1833 (N_1833,N_1738,N_1755);
and U1834 (N_1834,N_1788,N_1799);
nor U1835 (N_1835,N_1759,N_1732);
nor U1836 (N_1836,N_1727,N_1776);
or U1837 (N_1837,N_1789,N_1785);
xnor U1838 (N_1838,N_1729,N_1748);
xnor U1839 (N_1839,N_1757,N_1779);
nand U1840 (N_1840,N_1797,N_1775);
and U1841 (N_1841,N_1751,N_1748);
nor U1842 (N_1842,N_1729,N_1790);
and U1843 (N_1843,N_1734,N_1740);
nor U1844 (N_1844,N_1754,N_1762);
and U1845 (N_1845,N_1755,N_1782);
and U1846 (N_1846,N_1730,N_1785);
or U1847 (N_1847,N_1736,N_1787);
or U1848 (N_1848,N_1752,N_1759);
nor U1849 (N_1849,N_1798,N_1791);
or U1850 (N_1850,N_1751,N_1774);
nor U1851 (N_1851,N_1768,N_1796);
or U1852 (N_1852,N_1745,N_1767);
or U1853 (N_1853,N_1754,N_1778);
xnor U1854 (N_1854,N_1785,N_1780);
or U1855 (N_1855,N_1799,N_1766);
or U1856 (N_1856,N_1757,N_1789);
nor U1857 (N_1857,N_1743,N_1732);
nor U1858 (N_1858,N_1755,N_1727);
nor U1859 (N_1859,N_1786,N_1769);
or U1860 (N_1860,N_1746,N_1760);
nor U1861 (N_1861,N_1792,N_1777);
nor U1862 (N_1862,N_1742,N_1738);
nand U1863 (N_1863,N_1766,N_1753);
or U1864 (N_1864,N_1778,N_1799);
or U1865 (N_1865,N_1772,N_1764);
nand U1866 (N_1866,N_1727,N_1758);
or U1867 (N_1867,N_1798,N_1734);
nand U1868 (N_1868,N_1767,N_1738);
nand U1869 (N_1869,N_1751,N_1731);
nor U1870 (N_1870,N_1788,N_1790);
and U1871 (N_1871,N_1738,N_1750);
and U1872 (N_1872,N_1795,N_1748);
nand U1873 (N_1873,N_1729,N_1738);
and U1874 (N_1874,N_1726,N_1753);
and U1875 (N_1875,N_1802,N_1841);
xor U1876 (N_1876,N_1839,N_1803);
nand U1877 (N_1877,N_1834,N_1816);
nor U1878 (N_1878,N_1810,N_1874);
xnor U1879 (N_1879,N_1871,N_1823);
nor U1880 (N_1880,N_1865,N_1856);
nand U1881 (N_1881,N_1842,N_1827);
nor U1882 (N_1882,N_1858,N_1862);
or U1883 (N_1883,N_1811,N_1854);
nor U1884 (N_1884,N_1807,N_1815);
nor U1885 (N_1885,N_1873,N_1805);
or U1886 (N_1886,N_1831,N_1824);
or U1887 (N_1887,N_1808,N_1869);
and U1888 (N_1888,N_1825,N_1828);
nand U1889 (N_1889,N_1818,N_1846);
nor U1890 (N_1890,N_1837,N_1863);
and U1891 (N_1891,N_1832,N_1840);
nor U1892 (N_1892,N_1817,N_1872);
nand U1893 (N_1893,N_1830,N_1809);
nor U1894 (N_1894,N_1848,N_1868);
or U1895 (N_1895,N_1835,N_1833);
and U1896 (N_1896,N_1867,N_1801);
and U1897 (N_1897,N_1826,N_1870);
or U1898 (N_1898,N_1853,N_1861);
xnor U1899 (N_1899,N_1800,N_1857);
xnor U1900 (N_1900,N_1851,N_1819);
or U1901 (N_1901,N_1822,N_1820);
or U1902 (N_1902,N_1855,N_1821);
and U1903 (N_1903,N_1814,N_1813);
or U1904 (N_1904,N_1866,N_1843);
and U1905 (N_1905,N_1852,N_1812);
nor U1906 (N_1906,N_1804,N_1838);
or U1907 (N_1907,N_1829,N_1806);
or U1908 (N_1908,N_1844,N_1845);
nor U1909 (N_1909,N_1859,N_1860);
or U1910 (N_1910,N_1849,N_1836);
or U1911 (N_1911,N_1850,N_1864);
or U1912 (N_1912,N_1847,N_1834);
or U1913 (N_1913,N_1802,N_1824);
nor U1914 (N_1914,N_1821,N_1870);
nor U1915 (N_1915,N_1874,N_1803);
xnor U1916 (N_1916,N_1819,N_1852);
and U1917 (N_1917,N_1819,N_1800);
xnor U1918 (N_1918,N_1832,N_1804);
nand U1919 (N_1919,N_1827,N_1833);
nor U1920 (N_1920,N_1822,N_1867);
or U1921 (N_1921,N_1826,N_1864);
and U1922 (N_1922,N_1808,N_1849);
nor U1923 (N_1923,N_1826,N_1845);
and U1924 (N_1924,N_1832,N_1803);
nand U1925 (N_1925,N_1823,N_1825);
xor U1926 (N_1926,N_1814,N_1834);
and U1927 (N_1927,N_1857,N_1865);
nand U1928 (N_1928,N_1857,N_1841);
nor U1929 (N_1929,N_1845,N_1814);
or U1930 (N_1930,N_1839,N_1873);
nor U1931 (N_1931,N_1838,N_1818);
and U1932 (N_1932,N_1800,N_1804);
and U1933 (N_1933,N_1867,N_1830);
nor U1934 (N_1934,N_1808,N_1852);
and U1935 (N_1935,N_1856,N_1866);
xor U1936 (N_1936,N_1831,N_1803);
nand U1937 (N_1937,N_1829,N_1854);
and U1938 (N_1938,N_1858,N_1806);
nand U1939 (N_1939,N_1873,N_1820);
or U1940 (N_1940,N_1808,N_1827);
nor U1941 (N_1941,N_1814,N_1833);
and U1942 (N_1942,N_1848,N_1874);
and U1943 (N_1943,N_1818,N_1854);
and U1944 (N_1944,N_1807,N_1803);
and U1945 (N_1945,N_1870,N_1865);
xor U1946 (N_1946,N_1835,N_1842);
nor U1947 (N_1947,N_1856,N_1821);
and U1948 (N_1948,N_1843,N_1801);
and U1949 (N_1949,N_1814,N_1863);
nor U1950 (N_1950,N_1890,N_1889);
nand U1951 (N_1951,N_1882,N_1895);
xor U1952 (N_1952,N_1934,N_1898);
nand U1953 (N_1953,N_1940,N_1932);
or U1954 (N_1954,N_1906,N_1933);
nor U1955 (N_1955,N_1885,N_1880);
nor U1956 (N_1956,N_1894,N_1921);
or U1957 (N_1957,N_1916,N_1937);
or U1958 (N_1958,N_1920,N_1897);
xnor U1959 (N_1959,N_1919,N_1884);
nor U1960 (N_1960,N_1877,N_1939);
nor U1961 (N_1961,N_1887,N_1902);
nor U1962 (N_1962,N_1903,N_1904);
or U1963 (N_1963,N_1891,N_1943);
xnor U1964 (N_1964,N_1930,N_1929);
or U1965 (N_1965,N_1905,N_1881);
and U1966 (N_1966,N_1923,N_1896);
xor U1967 (N_1967,N_1888,N_1901);
and U1968 (N_1968,N_1922,N_1918);
xor U1969 (N_1969,N_1892,N_1878);
nand U1970 (N_1970,N_1917,N_1912);
or U1971 (N_1971,N_1926,N_1936);
nor U1972 (N_1972,N_1927,N_1908);
and U1973 (N_1973,N_1946,N_1900);
nor U1974 (N_1974,N_1893,N_1935);
nand U1975 (N_1975,N_1876,N_1907);
nor U1976 (N_1976,N_1938,N_1945);
xor U1977 (N_1977,N_1925,N_1913);
nand U1978 (N_1978,N_1942,N_1948);
and U1979 (N_1979,N_1924,N_1911);
or U1980 (N_1980,N_1914,N_1947);
nor U1981 (N_1981,N_1899,N_1941);
or U1982 (N_1982,N_1875,N_1915);
and U1983 (N_1983,N_1928,N_1879);
and U1984 (N_1984,N_1910,N_1949);
and U1985 (N_1985,N_1944,N_1883);
nand U1986 (N_1986,N_1909,N_1886);
or U1987 (N_1987,N_1931,N_1907);
and U1988 (N_1988,N_1918,N_1910);
nor U1989 (N_1989,N_1938,N_1921);
nor U1990 (N_1990,N_1923,N_1884);
nand U1991 (N_1991,N_1947,N_1944);
and U1992 (N_1992,N_1911,N_1887);
and U1993 (N_1993,N_1884,N_1945);
nand U1994 (N_1994,N_1924,N_1899);
nor U1995 (N_1995,N_1933,N_1905);
nor U1996 (N_1996,N_1897,N_1922);
nor U1997 (N_1997,N_1945,N_1914);
and U1998 (N_1998,N_1925,N_1899);
nand U1999 (N_1999,N_1900,N_1905);
and U2000 (N_2000,N_1917,N_1892);
or U2001 (N_2001,N_1894,N_1901);
nor U2002 (N_2002,N_1906,N_1913);
or U2003 (N_2003,N_1949,N_1878);
nor U2004 (N_2004,N_1880,N_1941);
and U2005 (N_2005,N_1890,N_1932);
or U2006 (N_2006,N_1923,N_1930);
nor U2007 (N_2007,N_1902,N_1913);
nand U2008 (N_2008,N_1920,N_1939);
and U2009 (N_2009,N_1890,N_1882);
or U2010 (N_2010,N_1920,N_1878);
and U2011 (N_2011,N_1948,N_1913);
nand U2012 (N_2012,N_1881,N_1889);
nor U2013 (N_2013,N_1932,N_1928);
nand U2014 (N_2014,N_1918,N_1912);
nor U2015 (N_2015,N_1913,N_1927);
nand U2016 (N_2016,N_1885,N_1949);
nor U2017 (N_2017,N_1897,N_1917);
nor U2018 (N_2018,N_1945,N_1893);
and U2019 (N_2019,N_1906,N_1922);
xor U2020 (N_2020,N_1924,N_1878);
or U2021 (N_2021,N_1948,N_1884);
and U2022 (N_2022,N_1899,N_1882);
nand U2023 (N_2023,N_1935,N_1932);
nand U2024 (N_2024,N_1936,N_1877);
nor U2025 (N_2025,N_2001,N_1954);
xnor U2026 (N_2026,N_1966,N_1962);
nand U2027 (N_2027,N_1959,N_1953);
nand U2028 (N_2028,N_2006,N_2024);
or U2029 (N_2029,N_1950,N_2007);
nor U2030 (N_2030,N_1971,N_1984);
nand U2031 (N_2031,N_1977,N_1968);
or U2032 (N_2032,N_1972,N_2009);
or U2033 (N_2033,N_2018,N_1952);
nand U2034 (N_2034,N_2023,N_1988);
nand U2035 (N_2035,N_1976,N_2011);
nand U2036 (N_2036,N_2022,N_1964);
and U2037 (N_2037,N_1981,N_2003);
or U2038 (N_2038,N_1985,N_2021);
nor U2039 (N_2039,N_2005,N_1979);
or U2040 (N_2040,N_1999,N_1991);
or U2041 (N_2041,N_2010,N_1989);
xnor U2042 (N_2042,N_1997,N_1996);
and U2043 (N_2043,N_1951,N_1974);
xor U2044 (N_2044,N_2004,N_1980);
xnor U2045 (N_2045,N_2015,N_1973);
xnor U2046 (N_2046,N_1978,N_2013);
or U2047 (N_2047,N_1998,N_1987);
nor U2048 (N_2048,N_1992,N_2002);
and U2049 (N_2049,N_2019,N_1958);
and U2050 (N_2050,N_1960,N_1982);
or U2051 (N_2051,N_2017,N_2000);
and U2052 (N_2052,N_1994,N_1967);
or U2053 (N_2053,N_2020,N_1995);
xor U2054 (N_2054,N_2008,N_1965);
and U2055 (N_2055,N_1963,N_2016);
nand U2056 (N_2056,N_1970,N_1956);
nor U2057 (N_2057,N_1957,N_1969);
nand U2058 (N_2058,N_1986,N_1990);
and U2059 (N_2059,N_1961,N_1993);
or U2060 (N_2060,N_1975,N_2012);
nand U2061 (N_2061,N_1955,N_1983);
and U2062 (N_2062,N_2014,N_2005);
nand U2063 (N_2063,N_1951,N_2003);
and U2064 (N_2064,N_1971,N_1957);
or U2065 (N_2065,N_1995,N_1993);
nand U2066 (N_2066,N_1953,N_1965);
and U2067 (N_2067,N_2009,N_1957);
nand U2068 (N_2068,N_1952,N_1994);
nand U2069 (N_2069,N_1984,N_1991);
or U2070 (N_2070,N_1993,N_2009);
nor U2071 (N_2071,N_1977,N_2018);
nor U2072 (N_2072,N_1968,N_2019);
nand U2073 (N_2073,N_1954,N_1950);
and U2074 (N_2074,N_2023,N_2003);
nand U2075 (N_2075,N_1974,N_2010);
nor U2076 (N_2076,N_2021,N_1955);
nor U2077 (N_2077,N_1985,N_1957);
or U2078 (N_2078,N_1984,N_1987);
or U2079 (N_2079,N_1962,N_1953);
nand U2080 (N_2080,N_2003,N_1974);
and U2081 (N_2081,N_1978,N_2017);
xor U2082 (N_2082,N_2003,N_1992);
or U2083 (N_2083,N_2008,N_1977);
or U2084 (N_2084,N_1981,N_1987);
nor U2085 (N_2085,N_1955,N_1968);
and U2086 (N_2086,N_2010,N_1966);
nor U2087 (N_2087,N_2014,N_2001);
nor U2088 (N_2088,N_2024,N_1998);
xor U2089 (N_2089,N_1950,N_1982);
nor U2090 (N_2090,N_1989,N_1956);
and U2091 (N_2091,N_1997,N_1953);
xnor U2092 (N_2092,N_1976,N_2012);
nor U2093 (N_2093,N_1988,N_1950);
nor U2094 (N_2094,N_1987,N_2020);
and U2095 (N_2095,N_1963,N_2023);
nor U2096 (N_2096,N_1987,N_1989);
nor U2097 (N_2097,N_1989,N_1988);
nand U2098 (N_2098,N_1968,N_1976);
and U2099 (N_2099,N_1998,N_1953);
or U2100 (N_2100,N_2035,N_2057);
nor U2101 (N_2101,N_2070,N_2086);
and U2102 (N_2102,N_2050,N_2067);
or U2103 (N_2103,N_2091,N_2084);
nor U2104 (N_2104,N_2099,N_2048);
or U2105 (N_2105,N_2038,N_2097);
or U2106 (N_2106,N_2092,N_2074);
nor U2107 (N_2107,N_2037,N_2029);
and U2108 (N_2108,N_2080,N_2025);
nor U2109 (N_2109,N_2085,N_2041);
nor U2110 (N_2110,N_2078,N_2071);
and U2111 (N_2111,N_2077,N_2090);
xnor U2112 (N_2112,N_2056,N_2026);
xor U2113 (N_2113,N_2094,N_2075);
nor U2114 (N_2114,N_2036,N_2051);
nand U2115 (N_2115,N_2032,N_2095);
nor U2116 (N_2116,N_2082,N_2081);
nor U2117 (N_2117,N_2028,N_2064);
nor U2118 (N_2118,N_2043,N_2049);
or U2119 (N_2119,N_2098,N_2093);
or U2120 (N_2120,N_2047,N_2044);
or U2121 (N_2121,N_2046,N_2060);
or U2122 (N_2122,N_2072,N_2083);
nor U2123 (N_2123,N_2052,N_2058);
and U2124 (N_2124,N_2045,N_2054);
nor U2125 (N_2125,N_2027,N_2059);
nor U2126 (N_2126,N_2055,N_2087);
or U2127 (N_2127,N_2079,N_2088);
or U2128 (N_2128,N_2063,N_2034);
and U2129 (N_2129,N_2066,N_2096);
xnor U2130 (N_2130,N_2073,N_2053);
nor U2131 (N_2131,N_2068,N_2076);
xnor U2132 (N_2132,N_2062,N_2061);
or U2133 (N_2133,N_2089,N_2069);
xor U2134 (N_2134,N_2065,N_2042);
nand U2135 (N_2135,N_2040,N_2031);
or U2136 (N_2136,N_2033,N_2039);
and U2137 (N_2137,N_2030,N_2058);
or U2138 (N_2138,N_2063,N_2095);
nor U2139 (N_2139,N_2056,N_2090);
nand U2140 (N_2140,N_2047,N_2093);
nor U2141 (N_2141,N_2062,N_2066);
nor U2142 (N_2142,N_2035,N_2044);
and U2143 (N_2143,N_2060,N_2035);
nand U2144 (N_2144,N_2078,N_2065);
or U2145 (N_2145,N_2038,N_2056);
and U2146 (N_2146,N_2084,N_2037);
or U2147 (N_2147,N_2096,N_2075);
nand U2148 (N_2148,N_2037,N_2073);
and U2149 (N_2149,N_2034,N_2090);
nor U2150 (N_2150,N_2076,N_2083);
nand U2151 (N_2151,N_2038,N_2034);
nand U2152 (N_2152,N_2083,N_2051);
xor U2153 (N_2153,N_2091,N_2067);
nand U2154 (N_2154,N_2089,N_2039);
or U2155 (N_2155,N_2094,N_2049);
or U2156 (N_2156,N_2072,N_2064);
nor U2157 (N_2157,N_2064,N_2057);
nand U2158 (N_2158,N_2061,N_2066);
nor U2159 (N_2159,N_2059,N_2045);
nand U2160 (N_2160,N_2033,N_2026);
nand U2161 (N_2161,N_2065,N_2050);
nand U2162 (N_2162,N_2071,N_2047);
nand U2163 (N_2163,N_2046,N_2048);
and U2164 (N_2164,N_2060,N_2039);
and U2165 (N_2165,N_2047,N_2096);
and U2166 (N_2166,N_2057,N_2099);
xnor U2167 (N_2167,N_2070,N_2089);
or U2168 (N_2168,N_2071,N_2050);
or U2169 (N_2169,N_2046,N_2036);
or U2170 (N_2170,N_2079,N_2025);
nand U2171 (N_2171,N_2086,N_2038);
nor U2172 (N_2172,N_2077,N_2092);
or U2173 (N_2173,N_2043,N_2084);
or U2174 (N_2174,N_2066,N_2048);
nand U2175 (N_2175,N_2170,N_2119);
or U2176 (N_2176,N_2161,N_2173);
nor U2177 (N_2177,N_2100,N_2121);
or U2178 (N_2178,N_2169,N_2112);
or U2179 (N_2179,N_2101,N_2129);
and U2180 (N_2180,N_2125,N_2124);
nor U2181 (N_2181,N_2118,N_2149);
xor U2182 (N_2182,N_2123,N_2160);
and U2183 (N_2183,N_2134,N_2145);
or U2184 (N_2184,N_2142,N_2106);
or U2185 (N_2185,N_2168,N_2164);
or U2186 (N_2186,N_2148,N_2154);
nor U2187 (N_2187,N_2163,N_2136);
and U2188 (N_2188,N_2171,N_2109);
nand U2189 (N_2189,N_2151,N_2130);
or U2190 (N_2190,N_2147,N_2152);
nor U2191 (N_2191,N_2165,N_2113);
nand U2192 (N_2192,N_2103,N_2155);
nor U2193 (N_2193,N_2153,N_2140);
nor U2194 (N_2194,N_2157,N_2115);
nor U2195 (N_2195,N_2127,N_2138);
and U2196 (N_2196,N_2126,N_2117);
and U2197 (N_2197,N_2102,N_2146);
xor U2198 (N_2198,N_2131,N_2156);
nand U2199 (N_2199,N_2122,N_2159);
and U2200 (N_2200,N_2128,N_2111);
nor U2201 (N_2201,N_2114,N_2137);
nor U2202 (N_2202,N_2166,N_2135);
or U2203 (N_2203,N_2107,N_2150);
nor U2204 (N_2204,N_2174,N_2105);
and U2205 (N_2205,N_2141,N_2104);
nand U2206 (N_2206,N_2120,N_2110);
or U2207 (N_2207,N_2162,N_2133);
nor U2208 (N_2208,N_2116,N_2143);
or U2209 (N_2209,N_2132,N_2172);
xor U2210 (N_2210,N_2158,N_2144);
nor U2211 (N_2211,N_2139,N_2167);
or U2212 (N_2212,N_2108,N_2172);
nand U2213 (N_2213,N_2108,N_2141);
nor U2214 (N_2214,N_2129,N_2167);
nor U2215 (N_2215,N_2160,N_2102);
nor U2216 (N_2216,N_2135,N_2112);
nand U2217 (N_2217,N_2164,N_2149);
and U2218 (N_2218,N_2165,N_2117);
nand U2219 (N_2219,N_2113,N_2123);
nor U2220 (N_2220,N_2115,N_2139);
and U2221 (N_2221,N_2162,N_2127);
or U2222 (N_2222,N_2101,N_2167);
and U2223 (N_2223,N_2148,N_2115);
nor U2224 (N_2224,N_2171,N_2122);
nand U2225 (N_2225,N_2143,N_2124);
and U2226 (N_2226,N_2127,N_2135);
nand U2227 (N_2227,N_2119,N_2101);
nand U2228 (N_2228,N_2162,N_2116);
or U2229 (N_2229,N_2109,N_2110);
xor U2230 (N_2230,N_2117,N_2166);
or U2231 (N_2231,N_2129,N_2124);
nand U2232 (N_2232,N_2128,N_2120);
and U2233 (N_2233,N_2121,N_2170);
or U2234 (N_2234,N_2142,N_2135);
or U2235 (N_2235,N_2137,N_2163);
or U2236 (N_2236,N_2147,N_2122);
and U2237 (N_2237,N_2119,N_2169);
or U2238 (N_2238,N_2103,N_2134);
nor U2239 (N_2239,N_2103,N_2120);
and U2240 (N_2240,N_2114,N_2171);
nand U2241 (N_2241,N_2158,N_2171);
or U2242 (N_2242,N_2105,N_2126);
nor U2243 (N_2243,N_2156,N_2158);
and U2244 (N_2244,N_2144,N_2169);
and U2245 (N_2245,N_2142,N_2111);
nor U2246 (N_2246,N_2142,N_2121);
nand U2247 (N_2247,N_2104,N_2166);
or U2248 (N_2248,N_2123,N_2144);
and U2249 (N_2249,N_2129,N_2159);
nand U2250 (N_2250,N_2175,N_2230);
nand U2251 (N_2251,N_2218,N_2202);
nor U2252 (N_2252,N_2190,N_2180);
and U2253 (N_2253,N_2212,N_2208);
nor U2254 (N_2254,N_2236,N_2201);
nor U2255 (N_2255,N_2211,N_2191);
nand U2256 (N_2256,N_2183,N_2195);
or U2257 (N_2257,N_2225,N_2199);
and U2258 (N_2258,N_2185,N_2224);
or U2259 (N_2259,N_2232,N_2245);
xnor U2260 (N_2260,N_2227,N_2178);
nor U2261 (N_2261,N_2177,N_2186);
xnor U2262 (N_2262,N_2246,N_2182);
or U2263 (N_2263,N_2192,N_2234);
and U2264 (N_2264,N_2228,N_2219);
and U2265 (N_2265,N_2214,N_2203);
or U2266 (N_2266,N_2210,N_2181);
nand U2267 (N_2267,N_2221,N_2204);
nand U2268 (N_2268,N_2220,N_2248);
or U2269 (N_2269,N_2249,N_2216);
or U2270 (N_2270,N_2179,N_2238);
xnor U2271 (N_2271,N_2194,N_2205);
xor U2272 (N_2272,N_2197,N_2187);
or U2273 (N_2273,N_2231,N_2243);
and U2274 (N_2274,N_2217,N_2247);
or U2275 (N_2275,N_2241,N_2196);
nand U2276 (N_2276,N_2198,N_2242);
nor U2277 (N_2277,N_2237,N_2222);
nand U2278 (N_2278,N_2240,N_2235);
and U2279 (N_2279,N_2206,N_2226);
nand U2280 (N_2280,N_2223,N_2213);
nor U2281 (N_2281,N_2239,N_2215);
and U2282 (N_2282,N_2244,N_2209);
or U2283 (N_2283,N_2233,N_2193);
xnor U2284 (N_2284,N_2176,N_2229);
nor U2285 (N_2285,N_2184,N_2200);
or U2286 (N_2286,N_2188,N_2207);
or U2287 (N_2287,N_2189,N_2241);
or U2288 (N_2288,N_2247,N_2228);
nand U2289 (N_2289,N_2238,N_2222);
nor U2290 (N_2290,N_2195,N_2186);
nor U2291 (N_2291,N_2218,N_2239);
xor U2292 (N_2292,N_2233,N_2201);
and U2293 (N_2293,N_2248,N_2193);
nand U2294 (N_2294,N_2180,N_2235);
or U2295 (N_2295,N_2241,N_2199);
or U2296 (N_2296,N_2188,N_2210);
and U2297 (N_2297,N_2179,N_2239);
nand U2298 (N_2298,N_2219,N_2246);
or U2299 (N_2299,N_2226,N_2229);
nor U2300 (N_2300,N_2212,N_2193);
and U2301 (N_2301,N_2239,N_2240);
nand U2302 (N_2302,N_2198,N_2245);
or U2303 (N_2303,N_2218,N_2211);
nor U2304 (N_2304,N_2207,N_2198);
or U2305 (N_2305,N_2235,N_2188);
nor U2306 (N_2306,N_2217,N_2230);
nand U2307 (N_2307,N_2191,N_2181);
and U2308 (N_2308,N_2219,N_2193);
nor U2309 (N_2309,N_2176,N_2195);
and U2310 (N_2310,N_2244,N_2215);
and U2311 (N_2311,N_2221,N_2228);
nand U2312 (N_2312,N_2203,N_2185);
or U2313 (N_2313,N_2194,N_2247);
and U2314 (N_2314,N_2192,N_2210);
xor U2315 (N_2315,N_2227,N_2230);
nor U2316 (N_2316,N_2211,N_2220);
nor U2317 (N_2317,N_2232,N_2178);
nor U2318 (N_2318,N_2217,N_2237);
nor U2319 (N_2319,N_2217,N_2181);
and U2320 (N_2320,N_2245,N_2179);
and U2321 (N_2321,N_2196,N_2219);
or U2322 (N_2322,N_2231,N_2219);
and U2323 (N_2323,N_2182,N_2202);
nand U2324 (N_2324,N_2213,N_2217);
or U2325 (N_2325,N_2250,N_2269);
nor U2326 (N_2326,N_2298,N_2296);
nor U2327 (N_2327,N_2251,N_2317);
nand U2328 (N_2328,N_2301,N_2321);
xor U2329 (N_2329,N_2306,N_2259);
nand U2330 (N_2330,N_2285,N_2308);
nor U2331 (N_2331,N_2300,N_2262);
or U2332 (N_2332,N_2261,N_2311);
or U2333 (N_2333,N_2256,N_2299);
nand U2334 (N_2334,N_2295,N_2279);
nor U2335 (N_2335,N_2322,N_2314);
or U2336 (N_2336,N_2255,N_2268);
nand U2337 (N_2337,N_2276,N_2278);
and U2338 (N_2338,N_2260,N_2304);
nand U2339 (N_2339,N_2252,N_2313);
xnor U2340 (N_2340,N_2270,N_2274);
nand U2341 (N_2341,N_2309,N_2312);
and U2342 (N_2342,N_2264,N_2310);
nor U2343 (N_2343,N_2282,N_2290);
nor U2344 (N_2344,N_2275,N_2266);
nor U2345 (N_2345,N_2253,N_2316);
nand U2346 (N_2346,N_2323,N_2280);
and U2347 (N_2347,N_2263,N_2283);
and U2348 (N_2348,N_2293,N_2288);
nor U2349 (N_2349,N_2273,N_2315);
nand U2350 (N_2350,N_2271,N_2320);
nor U2351 (N_2351,N_2257,N_2318);
nand U2352 (N_2352,N_2324,N_2254);
nand U2353 (N_2353,N_2292,N_2305);
nor U2354 (N_2354,N_2319,N_2284);
nor U2355 (N_2355,N_2291,N_2265);
nor U2356 (N_2356,N_2307,N_2272);
nand U2357 (N_2357,N_2297,N_2294);
nand U2358 (N_2358,N_2289,N_2267);
nor U2359 (N_2359,N_2287,N_2258);
and U2360 (N_2360,N_2281,N_2277);
nor U2361 (N_2361,N_2286,N_2302);
or U2362 (N_2362,N_2303,N_2292);
nor U2363 (N_2363,N_2298,N_2276);
or U2364 (N_2364,N_2270,N_2255);
nand U2365 (N_2365,N_2265,N_2281);
and U2366 (N_2366,N_2281,N_2250);
and U2367 (N_2367,N_2276,N_2280);
or U2368 (N_2368,N_2251,N_2290);
or U2369 (N_2369,N_2320,N_2251);
nor U2370 (N_2370,N_2316,N_2252);
and U2371 (N_2371,N_2260,N_2319);
and U2372 (N_2372,N_2313,N_2269);
nand U2373 (N_2373,N_2295,N_2321);
xor U2374 (N_2374,N_2272,N_2254);
or U2375 (N_2375,N_2319,N_2254);
nor U2376 (N_2376,N_2304,N_2280);
or U2377 (N_2377,N_2301,N_2294);
and U2378 (N_2378,N_2314,N_2271);
nor U2379 (N_2379,N_2272,N_2258);
and U2380 (N_2380,N_2314,N_2281);
or U2381 (N_2381,N_2323,N_2268);
or U2382 (N_2382,N_2255,N_2311);
or U2383 (N_2383,N_2315,N_2257);
nor U2384 (N_2384,N_2269,N_2262);
or U2385 (N_2385,N_2267,N_2287);
nand U2386 (N_2386,N_2253,N_2309);
or U2387 (N_2387,N_2285,N_2280);
xor U2388 (N_2388,N_2287,N_2285);
nor U2389 (N_2389,N_2321,N_2276);
and U2390 (N_2390,N_2296,N_2314);
and U2391 (N_2391,N_2258,N_2308);
xnor U2392 (N_2392,N_2272,N_2273);
nand U2393 (N_2393,N_2292,N_2257);
or U2394 (N_2394,N_2267,N_2301);
or U2395 (N_2395,N_2252,N_2309);
nor U2396 (N_2396,N_2251,N_2265);
nor U2397 (N_2397,N_2290,N_2257);
and U2398 (N_2398,N_2252,N_2288);
xor U2399 (N_2399,N_2324,N_2280);
or U2400 (N_2400,N_2372,N_2339);
and U2401 (N_2401,N_2392,N_2390);
or U2402 (N_2402,N_2333,N_2352);
nand U2403 (N_2403,N_2366,N_2389);
and U2404 (N_2404,N_2341,N_2325);
nand U2405 (N_2405,N_2386,N_2399);
nand U2406 (N_2406,N_2393,N_2355);
and U2407 (N_2407,N_2346,N_2363);
xor U2408 (N_2408,N_2376,N_2326);
nand U2409 (N_2409,N_2358,N_2336);
and U2410 (N_2410,N_2344,N_2388);
xor U2411 (N_2411,N_2396,N_2338);
nand U2412 (N_2412,N_2334,N_2345);
xnor U2413 (N_2413,N_2394,N_2375);
or U2414 (N_2414,N_2356,N_2382);
nor U2415 (N_2415,N_2350,N_2370);
and U2416 (N_2416,N_2385,N_2348);
nor U2417 (N_2417,N_2343,N_2395);
xnor U2418 (N_2418,N_2342,N_2383);
xnor U2419 (N_2419,N_2367,N_2328);
nor U2420 (N_2420,N_2360,N_2353);
nand U2421 (N_2421,N_2369,N_2384);
and U2422 (N_2422,N_2354,N_2398);
or U2423 (N_2423,N_2364,N_2357);
xor U2424 (N_2424,N_2381,N_2359);
nor U2425 (N_2425,N_2327,N_2374);
nor U2426 (N_2426,N_2332,N_2380);
nand U2427 (N_2427,N_2379,N_2373);
xnor U2428 (N_2428,N_2371,N_2347);
nor U2429 (N_2429,N_2330,N_2351);
or U2430 (N_2430,N_2387,N_2362);
and U2431 (N_2431,N_2365,N_2391);
nor U2432 (N_2432,N_2361,N_2349);
or U2433 (N_2433,N_2337,N_2331);
and U2434 (N_2434,N_2329,N_2335);
nand U2435 (N_2435,N_2397,N_2377);
nor U2436 (N_2436,N_2368,N_2378);
and U2437 (N_2437,N_2340,N_2355);
nand U2438 (N_2438,N_2325,N_2339);
nand U2439 (N_2439,N_2361,N_2358);
nor U2440 (N_2440,N_2342,N_2340);
nor U2441 (N_2441,N_2372,N_2369);
nor U2442 (N_2442,N_2334,N_2391);
and U2443 (N_2443,N_2361,N_2338);
and U2444 (N_2444,N_2362,N_2379);
and U2445 (N_2445,N_2368,N_2370);
xor U2446 (N_2446,N_2375,N_2371);
nor U2447 (N_2447,N_2327,N_2331);
or U2448 (N_2448,N_2363,N_2342);
xor U2449 (N_2449,N_2376,N_2328);
xnor U2450 (N_2450,N_2335,N_2362);
nand U2451 (N_2451,N_2342,N_2398);
nand U2452 (N_2452,N_2395,N_2396);
xor U2453 (N_2453,N_2389,N_2326);
xnor U2454 (N_2454,N_2375,N_2392);
nand U2455 (N_2455,N_2383,N_2370);
or U2456 (N_2456,N_2376,N_2358);
nand U2457 (N_2457,N_2394,N_2383);
nand U2458 (N_2458,N_2356,N_2387);
or U2459 (N_2459,N_2343,N_2367);
and U2460 (N_2460,N_2336,N_2394);
nand U2461 (N_2461,N_2370,N_2373);
nor U2462 (N_2462,N_2375,N_2328);
nor U2463 (N_2463,N_2358,N_2330);
nor U2464 (N_2464,N_2392,N_2341);
xnor U2465 (N_2465,N_2372,N_2366);
nor U2466 (N_2466,N_2384,N_2332);
or U2467 (N_2467,N_2359,N_2376);
and U2468 (N_2468,N_2383,N_2371);
xnor U2469 (N_2469,N_2384,N_2329);
or U2470 (N_2470,N_2350,N_2346);
nor U2471 (N_2471,N_2341,N_2342);
or U2472 (N_2472,N_2339,N_2348);
nor U2473 (N_2473,N_2394,N_2372);
nand U2474 (N_2474,N_2395,N_2367);
or U2475 (N_2475,N_2414,N_2429);
or U2476 (N_2476,N_2460,N_2463);
and U2477 (N_2477,N_2458,N_2472);
nand U2478 (N_2478,N_2455,N_2422);
nand U2479 (N_2479,N_2418,N_2438);
or U2480 (N_2480,N_2451,N_2426);
or U2481 (N_2481,N_2424,N_2403);
xor U2482 (N_2482,N_2419,N_2447);
xor U2483 (N_2483,N_2411,N_2412);
nand U2484 (N_2484,N_2456,N_2413);
xnor U2485 (N_2485,N_2410,N_2437);
or U2486 (N_2486,N_2465,N_2474);
and U2487 (N_2487,N_2462,N_2471);
xor U2488 (N_2488,N_2433,N_2452);
or U2489 (N_2489,N_2416,N_2407);
or U2490 (N_2490,N_2434,N_2466);
nand U2491 (N_2491,N_2409,N_2473);
nor U2492 (N_2492,N_2408,N_2468);
nor U2493 (N_2493,N_2402,N_2428);
nor U2494 (N_2494,N_2443,N_2430);
xnor U2495 (N_2495,N_2440,N_2401);
xnor U2496 (N_2496,N_2470,N_2454);
nand U2497 (N_2497,N_2449,N_2423);
or U2498 (N_2498,N_2425,N_2448);
or U2499 (N_2499,N_2446,N_2415);
and U2500 (N_2500,N_2405,N_2431);
or U2501 (N_2501,N_2406,N_2453);
or U2502 (N_2502,N_2461,N_2435);
nand U2503 (N_2503,N_2400,N_2444);
nand U2504 (N_2504,N_2420,N_2469);
and U2505 (N_2505,N_2459,N_2421);
nor U2506 (N_2506,N_2457,N_2464);
or U2507 (N_2507,N_2467,N_2432);
nand U2508 (N_2508,N_2404,N_2445);
nor U2509 (N_2509,N_2439,N_2441);
or U2510 (N_2510,N_2417,N_2436);
and U2511 (N_2511,N_2442,N_2450);
or U2512 (N_2512,N_2427,N_2410);
nand U2513 (N_2513,N_2437,N_2436);
nor U2514 (N_2514,N_2434,N_2436);
nand U2515 (N_2515,N_2447,N_2443);
or U2516 (N_2516,N_2449,N_2428);
nor U2517 (N_2517,N_2453,N_2410);
nor U2518 (N_2518,N_2402,N_2471);
or U2519 (N_2519,N_2472,N_2444);
xnor U2520 (N_2520,N_2432,N_2463);
nand U2521 (N_2521,N_2401,N_2472);
nor U2522 (N_2522,N_2474,N_2402);
and U2523 (N_2523,N_2418,N_2413);
xnor U2524 (N_2524,N_2451,N_2416);
nand U2525 (N_2525,N_2445,N_2453);
nand U2526 (N_2526,N_2459,N_2437);
nor U2527 (N_2527,N_2409,N_2470);
nor U2528 (N_2528,N_2464,N_2429);
nor U2529 (N_2529,N_2453,N_2449);
nor U2530 (N_2530,N_2443,N_2402);
or U2531 (N_2531,N_2433,N_2401);
nand U2532 (N_2532,N_2404,N_2451);
nand U2533 (N_2533,N_2408,N_2474);
nor U2534 (N_2534,N_2437,N_2412);
nand U2535 (N_2535,N_2454,N_2415);
nor U2536 (N_2536,N_2464,N_2419);
nand U2537 (N_2537,N_2474,N_2446);
and U2538 (N_2538,N_2447,N_2407);
nor U2539 (N_2539,N_2469,N_2431);
or U2540 (N_2540,N_2428,N_2418);
nor U2541 (N_2541,N_2463,N_2405);
nand U2542 (N_2542,N_2400,N_2448);
and U2543 (N_2543,N_2459,N_2436);
or U2544 (N_2544,N_2458,N_2421);
xnor U2545 (N_2545,N_2420,N_2441);
and U2546 (N_2546,N_2401,N_2471);
nor U2547 (N_2547,N_2422,N_2426);
nor U2548 (N_2548,N_2464,N_2469);
nand U2549 (N_2549,N_2411,N_2473);
nor U2550 (N_2550,N_2536,N_2544);
and U2551 (N_2551,N_2487,N_2497);
or U2552 (N_2552,N_2495,N_2532);
or U2553 (N_2553,N_2533,N_2488);
xnor U2554 (N_2554,N_2477,N_2547);
or U2555 (N_2555,N_2510,N_2520);
nand U2556 (N_2556,N_2475,N_2494);
nand U2557 (N_2557,N_2541,N_2522);
or U2558 (N_2558,N_2489,N_2492);
nor U2559 (N_2559,N_2525,N_2546);
nor U2560 (N_2560,N_2506,N_2485);
nor U2561 (N_2561,N_2545,N_2515);
xnor U2562 (N_2562,N_2540,N_2543);
nor U2563 (N_2563,N_2493,N_2476);
or U2564 (N_2564,N_2504,N_2512);
and U2565 (N_2565,N_2529,N_2549);
xor U2566 (N_2566,N_2513,N_2524);
nand U2567 (N_2567,N_2535,N_2480);
or U2568 (N_2568,N_2483,N_2537);
or U2569 (N_2569,N_2499,N_2490);
nor U2570 (N_2570,N_2517,N_2518);
nor U2571 (N_2571,N_2548,N_2496);
nand U2572 (N_2572,N_2530,N_2507);
or U2573 (N_2573,N_2508,N_2503);
or U2574 (N_2574,N_2500,N_2514);
nor U2575 (N_2575,N_2538,N_2526);
and U2576 (N_2576,N_2479,N_2505);
xnor U2577 (N_2577,N_2509,N_2531);
and U2578 (N_2578,N_2498,N_2542);
or U2579 (N_2579,N_2521,N_2511);
xor U2580 (N_2580,N_2527,N_2519);
and U2581 (N_2581,N_2539,N_2486);
or U2582 (N_2582,N_2491,N_2501);
nor U2583 (N_2583,N_2482,N_2502);
nand U2584 (N_2584,N_2523,N_2516);
nand U2585 (N_2585,N_2478,N_2481);
nand U2586 (N_2586,N_2484,N_2534);
and U2587 (N_2587,N_2528,N_2505);
nand U2588 (N_2588,N_2481,N_2514);
nand U2589 (N_2589,N_2539,N_2495);
xnor U2590 (N_2590,N_2540,N_2504);
xnor U2591 (N_2591,N_2518,N_2493);
nor U2592 (N_2592,N_2493,N_2494);
nor U2593 (N_2593,N_2548,N_2511);
and U2594 (N_2594,N_2482,N_2475);
and U2595 (N_2595,N_2514,N_2519);
and U2596 (N_2596,N_2522,N_2491);
or U2597 (N_2597,N_2477,N_2483);
and U2598 (N_2598,N_2548,N_2514);
or U2599 (N_2599,N_2487,N_2542);
and U2600 (N_2600,N_2515,N_2514);
nor U2601 (N_2601,N_2537,N_2542);
nand U2602 (N_2602,N_2534,N_2486);
or U2603 (N_2603,N_2515,N_2543);
or U2604 (N_2604,N_2495,N_2527);
nor U2605 (N_2605,N_2482,N_2481);
nand U2606 (N_2606,N_2505,N_2544);
or U2607 (N_2607,N_2540,N_2542);
nor U2608 (N_2608,N_2477,N_2518);
and U2609 (N_2609,N_2546,N_2533);
or U2610 (N_2610,N_2485,N_2507);
nand U2611 (N_2611,N_2545,N_2514);
xor U2612 (N_2612,N_2546,N_2536);
or U2613 (N_2613,N_2478,N_2526);
nor U2614 (N_2614,N_2508,N_2542);
xnor U2615 (N_2615,N_2501,N_2513);
or U2616 (N_2616,N_2536,N_2530);
nand U2617 (N_2617,N_2483,N_2480);
and U2618 (N_2618,N_2538,N_2494);
nor U2619 (N_2619,N_2479,N_2504);
xor U2620 (N_2620,N_2526,N_2534);
and U2621 (N_2621,N_2499,N_2538);
or U2622 (N_2622,N_2548,N_2502);
or U2623 (N_2623,N_2481,N_2487);
and U2624 (N_2624,N_2514,N_2498);
nand U2625 (N_2625,N_2557,N_2579);
nor U2626 (N_2626,N_2620,N_2589);
nor U2627 (N_2627,N_2610,N_2566);
nand U2628 (N_2628,N_2615,N_2619);
and U2629 (N_2629,N_2577,N_2587);
nand U2630 (N_2630,N_2569,N_2572);
and U2631 (N_2631,N_2601,N_2608);
nor U2632 (N_2632,N_2612,N_2554);
or U2633 (N_2633,N_2597,N_2624);
nor U2634 (N_2634,N_2564,N_2563);
nand U2635 (N_2635,N_2602,N_2586);
nand U2636 (N_2636,N_2604,N_2613);
nor U2637 (N_2637,N_2616,N_2559);
nor U2638 (N_2638,N_2603,N_2565);
nand U2639 (N_2639,N_2576,N_2575);
nor U2640 (N_2640,N_2598,N_2592);
and U2641 (N_2641,N_2617,N_2570);
nand U2642 (N_2642,N_2552,N_2584);
or U2643 (N_2643,N_2571,N_2574);
nor U2644 (N_2644,N_2556,N_2591);
nand U2645 (N_2645,N_2551,N_2558);
or U2646 (N_2646,N_2573,N_2555);
or U2647 (N_2647,N_2596,N_2560);
or U2648 (N_2648,N_2618,N_2578);
and U2649 (N_2649,N_2582,N_2567);
xnor U2650 (N_2650,N_2595,N_2568);
nand U2651 (N_2651,N_2580,N_2606);
or U2652 (N_2652,N_2623,N_2614);
nand U2653 (N_2653,N_2607,N_2593);
or U2654 (N_2654,N_2561,N_2588);
nand U2655 (N_2655,N_2605,N_2550);
nor U2656 (N_2656,N_2594,N_2553);
nand U2657 (N_2657,N_2609,N_2590);
and U2658 (N_2658,N_2611,N_2583);
or U2659 (N_2659,N_2622,N_2600);
and U2660 (N_2660,N_2581,N_2585);
nor U2661 (N_2661,N_2621,N_2562);
nor U2662 (N_2662,N_2599,N_2562);
nand U2663 (N_2663,N_2572,N_2592);
and U2664 (N_2664,N_2566,N_2571);
and U2665 (N_2665,N_2561,N_2557);
and U2666 (N_2666,N_2550,N_2568);
nor U2667 (N_2667,N_2563,N_2560);
nor U2668 (N_2668,N_2568,N_2587);
nand U2669 (N_2669,N_2587,N_2616);
or U2670 (N_2670,N_2562,N_2623);
xor U2671 (N_2671,N_2563,N_2575);
nor U2672 (N_2672,N_2559,N_2620);
xnor U2673 (N_2673,N_2584,N_2573);
nor U2674 (N_2674,N_2565,N_2601);
nor U2675 (N_2675,N_2591,N_2566);
nor U2676 (N_2676,N_2621,N_2587);
or U2677 (N_2677,N_2581,N_2616);
nand U2678 (N_2678,N_2609,N_2596);
nand U2679 (N_2679,N_2578,N_2567);
and U2680 (N_2680,N_2599,N_2575);
xor U2681 (N_2681,N_2577,N_2574);
and U2682 (N_2682,N_2557,N_2576);
nand U2683 (N_2683,N_2561,N_2605);
xor U2684 (N_2684,N_2618,N_2574);
nand U2685 (N_2685,N_2556,N_2573);
nor U2686 (N_2686,N_2620,N_2554);
and U2687 (N_2687,N_2623,N_2582);
nand U2688 (N_2688,N_2572,N_2607);
nand U2689 (N_2689,N_2560,N_2556);
nor U2690 (N_2690,N_2582,N_2581);
xnor U2691 (N_2691,N_2567,N_2594);
or U2692 (N_2692,N_2551,N_2592);
and U2693 (N_2693,N_2608,N_2596);
nor U2694 (N_2694,N_2607,N_2554);
and U2695 (N_2695,N_2609,N_2624);
or U2696 (N_2696,N_2578,N_2594);
and U2697 (N_2697,N_2608,N_2583);
nand U2698 (N_2698,N_2559,N_2553);
and U2699 (N_2699,N_2602,N_2618);
nor U2700 (N_2700,N_2662,N_2631);
nand U2701 (N_2701,N_2681,N_2650);
nand U2702 (N_2702,N_2644,N_2687);
nand U2703 (N_2703,N_2649,N_2684);
nand U2704 (N_2704,N_2635,N_2647);
nand U2705 (N_2705,N_2657,N_2690);
nand U2706 (N_2706,N_2651,N_2656);
or U2707 (N_2707,N_2627,N_2699);
or U2708 (N_2708,N_2645,N_2676);
or U2709 (N_2709,N_2679,N_2672);
or U2710 (N_2710,N_2685,N_2675);
and U2711 (N_2711,N_2669,N_2655);
nand U2712 (N_2712,N_2630,N_2643);
and U2713 (N_2713,N_2668,N_2692);
nor U2714 (N_2714,N_2674,N_2639);
or U2715 (N_2715,N_2683,N_2665);
and U2716 (N_2716,N_2660,N_2628);
nand U2717 (N_2717,N_2678,N_2663);
nor U2718 (N_2718,N_2637,N_2694);
or U2719 (N_2719,N_2688,N_2634);
nor U2720 (N_2720,N_2640,N_2696);
and U2721 (N_2721,N_2682,N_2695);
nor U2722 (N_2722,N_2680,N_2638);
nand U2723 (N_2723,N_2677,N_2654);
or U2724 (N_2724,N_2666,N_2664);
and U2725 (N_2725,N_2686,N_2641);
and U2726 (N_2726,N_2632,N_2673);
or U2727 (N_2727,N_2671,N_2653);
and U2728 (N_2728,N_2689,N_2625);
nor U2729 (N_2729,N_2698,N_2697);
nand U2730 (N_2730,N_2633,N_2646);
and U2731 (N_2731,N_2648,N_2659);
nor U2732 (N_2732,N_2626,N_2642);
nand U2733 (N_2733,N_2667,N_2691);
xnor U2734 (N_2734,N_2661,N_2658);
nor U2735 (N_2735,N_2629,N_2652);
and U2736 (N_2736,N_2693,N_2636);
and U2737 (N_2737,N_2670,N_2691);
and U2738 (N_2738,N_2626,N_2672);
and U2739 (N_2739,N_2647,N_2662);
and U2740 (N_2740,N_2644,N_2628);
or U2741 (N_2741,N_2644,N_2661);
or U2742 (N_2742,N_2694,N_2672);
or U2743 (N_2743,N_2636,N_2645);
or U2744 (N_2744,N_2640,N_2659);
nor U2745 (N_2745,N_2653,N_2638);
and U2746 (N_2746,N_2656,N_2676);
and U2747 (N_2747,N_2657,N_2672);
nor U2748 (N_2748,N_2634,N_2697);
nand U2749 (N_2749,N_2678,N_2653);
or U2750 (N_2750,N_2636,N_2692);
xor U2751 (N_2751,N_2648,N_2686);
nand U2752 (N_2752,N_2691,N_2656);
nand U2753 (N_2753,N_2689,N_2663);
nand U2754 (N_2754,N_2632,N_2655);
nand U2755 (N_2755,N_2698,N_2659);
nand U2756 (N_2756,N_2650,N_2699);
and U2757 (N_2757,N_2687,N_2628);
nand U2758 (N_2758,N_2659,N_2688);
nor U2759 (N_2759,N_2688,N_2671);
nand U2760 (N_2760,N_2669,N_2665);
nor U2761 (N_2761,N_2657,N_2637);
or U2762 (N_2762,N_2677,N_2665);
and U2763 (N_2763,N_2666,N_2629);
xnor U2764 (N_2764,N_2682,N_2672);
or U2765 (N_2765,N_2685,N_2630);
and U2766 (N_2766,N_2628,N_2626);
nand U2767 (N_2767,N_2635,N_2638);
or U2768 (N_2768,N_2638,N_2650);
nand U2769 (N_2769,N_2626,N_2676);
nand U2770 (N_2770,N_2678,N_2625);
or U2771 (N_2771,N_2697,N_2693);
xor U2772 (N_2772,N_2657,N_2640);
nand U2773 (N_2773,N_2698,N_2638);
nor U2774 (N_2774,N_2639,N_2689);
or U2775 (N_2775,N_2731,N_2755);
and U2776 (N_2776,N_2756,N_2763);
nand U2777 (N_2777,N_2760,N_2717);
nand U2778 (N_2778,N_2769,N_2773);
nor U2779 (N_2779,N_2710,N_2730);
and U2780 (N_2780,N_2707,N_2754);
and U2781 (N_2781,N_2718,N_2700);
and U2782 (N_2782,N_2747,N_2706);
or U2783 (N_2783,N_2757,N_2729);
nand U2784 (N_2784,N_2758,N_2750);
or U2785 (N_2785,N_2765,N_2744);
nand U2786 (N_2786,N_2702,N_2746);
xnor U2787 (N_2787,N_2745,N_2738);
and U2788 (N_2788,N_2711,N_2737);
and U2789 (N_2789,N_2725,N_2774);
nand U2790 (N_2790,N_2727,N_2719);
nand U2791 (N_2791,N_2726,N_2742);
nand U2792 (N_2792,N_2733,N_2766);
xor U2793 (N_2793,N_2741,N_2771);
or U2794 (N_2794,N_2770,N_2739);
nor U2795 (N_2795,N_2764,N_2736);
or U2796 (N_2796,N_2715,N_2703);
and U2797 (N_2797,N_2752,N_2748);
nor U2798 (N_2798,N_2743,N_2735);
nor U2799 (N_2799,N_2704,N_2712);
nor U2800 (N_2800,N_2716,N_2722);
and U2801 (N_2801,N_2772,N_2759);
nand U2802 (N_2802,N_2728,N_2768);
or U2803 (N_2803,N_2749,N_2708);
or U2804 (N_2804,N_2701,N_2762);
nor U2805 (N_2805,N_2721,N_2740);
or U2806 (N_2806,N_2767,N_2732);
or U2807 (N_2807,N_2724,N_2761);
and U2808 (N_2808,N_2734,N_2753);
or U2809 (N_2809,N_2751,N_2720);
nor U2810 (N_2810,N_2714,N_2705);
nor U2811 (N_2811,N_2713,N_2723);
or U2812 (N_2812,N_2709,N_2723);
and U2813 (N_2813,N_2724,N_2747);
nand U2814 (N_2814,N_2721,N_2758);
nor U2815 (N_2815,N_2765,N_2764);
nand U2816 (N_2816,N_2720,N_2723);
or U2817 (N_2817,N_2760,N_2754);
nand U2818 (N_2818,N_2715,N_2709);
nor U2819 (N_2819,N_2715,N_2757);
nand U2820 (N_2820,N_2741,N_2766);
or U2821 (N_2821,N_2740,N_2726);
or U2822 (N_2822,N_2725,N_2728);
or U2823 (N_2823,N_2729,N_2763);
or U2824 (N_2824,N_2728,N_2764);
and U2825 (N_2825,N_2751,N_2762);
nand U2826 (N_2826,N_2766,N_2705);
nor U2827 (N_2827,N_2754,N_2743);
nand U2828 (N_2828,N_2746,N_2755);
nand U2829 (N_2829,N_2767,N_2703);
xnor U2830 (N_2830,N_2726,N_2730);
nand U2831 (N_2831,N_2768,N_2702);
and U2832 (N_2832,N_2737,N_2758);
nand U2833 (N_2833,N_2720,N_2708);
and U2834 (N_2834,N_2707,N_2747);
or U2835 (N_2835,N_2739,N_2703);
nor U2836 (N_2836,N_2731,N_2757);
nand U2837 (N_2837,N_2770,N_2731);
or U2838 (N_2838,N_2700,N_2773);
nor U2839 (N_2839,N_2752,N_2730);
nor U2840 (N_2840,N_2723,N_2705);
nand U2841 (N_2841,N_2738,N_2720);
or U2842 (N_2842,N_2738,N_2713);
nor U2843 (N_2843,N_2754,N_2750);
nor U2844 (N_2844,N_2708,N_2724);
and U2845 (N_2845,N_2715,N_2716);
nand U2846 (N_2846,N_2751,N_2736);
or U2847 (N_2847,N_2741,N_2772);
nor U2848 (N_2848,N_2702,N_2750);
nor U2849 (N_2849,N_2711,N_2765);
and U2850 (N_2850,N_2826,N_2820);
and U2851 (N_2851,N_2818,N_2783);
nand U2852 (N_2852,N_2788,N_2787);
nand U2853 (N_2853,N_2800,N_2823);
nor U2854 (N_2854,N_2844,N_2815);
or U2855 (N_2855,N_2845,N_2849);
or U2856 (N_2856,N_2782,N_2778);
nor U2857 (N_2857,N_2840,N_2785);
or U2858 (N_2858,N_2821,N_2791);
or U2859 (N_2859,N_2808,N_2848);
and U2860 (N_2860,N_2781,N_2802);
and U2861 (N_2861,N_2841,N_2795);
or U2862 (N_2862,N_2811,N_2838);
nor U2863 (N_2863,N_2777,N_2837);
or U2864 (N_2864,N_2799,N_2789);
nor U2865 (N_2865,N_2779,N_2817);
and U2866 (N_2866,N_2797,N_2831);
nor U2867 (N_2867,N_2825,N_2806);
nor U2868 (N_2868,N_2835,N_2809);
nand U2869 (N_2869,N_2843,N_2847);
nand U2870 (N_2870,N_2776,N_2798);
xnor U2871 (N_2871,N_2805,N_2793);
or U2872 (N_2872,N_2828,N_2836);
nand U2873 (N_2873,N_2842,N_2813);
nor U2874 (N_2874,N_2814,N_2790);
nor U2875 (N_2875,N_2792,N_2829);
or U2876 (N_2876,N_2796,N_2812);
nor U2877 (N_2877,N_2822,N_2801);
nand U2878 (N_2878,N_2830,N_2827);
nor U2879 (N_2879,N_2816,N_2846);
nand U2880 (N_2880,N_2832,N_2784);
nor U2881 (N_2881,N_2834,N_2794);
nand U2882 (N_2882,N_2819,N_2804);
nor U2883 (N_2883,N_2807,N_2833);
or U2884 (N_2884,N_2780,N_2786);
nand U2885 (N_2885,N_2775,N_2824);
nor U2886 (N_2886,N_2803,N_2810);
nor U2887 (N_2887,N_2839,N_2831);
nand U2888 (N_2888,N_2803,N_2819);
or U2889 (N_2889,N_2824,N_2845);
or U2890 (N_2890,N_2821,N_2779);
nand U2891 (N_2891,N_2792,N_2791);
nand U2892 (N_2892,N_2788,N_2781);
and U2893 (N_2893,N_2805,N_2818);
nor U2894 (N_2894,N_2809,N_2839);
and U2895 (N_2895,N_2783,N_2787);
and U2896 (N_2896,N_2782,N_2786);
nand U2897 (N_2897,N_2794,N_2802);
or U2898 (N_2898,N_2797,N_2818);
nand U2899 (N_2899,N_2824,N_2807);
nor U2900 (N_2900,N_2810,N_2826);
xor U2901 (N_2901,N_2835,N_2830);
and U2902 (N_2902,N_2801,N_2788);
and U2903 (N_2903,N_2835,N_2814);
xnor U2904 (N_2904,N_2839,N_2775);
nand U2905 (N_2905,N_2828,N_2786);
and U2906 (N_2906,N_2782,N_2827);
nand U2907 (N_2907,N_2835,N_2798);
or U2908 (N_2908,N_2824,N_2826);
nand U2909 (N_2909,N_2812,N_2776);
nor U2910 (N_2910,N_2848,N_2810);
or U2911 (N_2911,N_2849,N_2803);
nor U2912 (N_2912,N_2801,N_2786);
nand U2913 (N_2913,N_2800,N_2776);
nor U2914 (N_2914,N_2849,N_2790);
nand U2915 (N_2915,N_2829,N_2777);
or U2916 (N_2916,N_2796,N_2825);
xor U2917 (N_2917,N_2822,N_2834);
and U2918 (N_2918,N_2787,N_2836);
nand U2919 (N_2919,N_2849,N_2805);
and U2920 (N_2920,N_2783,N_2842);
nand U2921 (N_2921,N_2840,N_2802);
or U2922 (N_2922,N_2830,N_2836);
nor U2923 (N_2923,N_2816,N_2841);
nand U2924 (N_2924,N_2788,N_2826);
and U2925 (N_2925,N_2857,N_2894);
or U2926 (N_2926,N_2911,N_2872);
or U2927 (N_2927,N_2861,N_2908);
xor U2928 (N_2928,N_2879,N_2866);
nor U2929 (N_2929,N_2891,N_2902);
xnor U2930 (N_2930,N_2889,N_2876);
nand U2931 (N_2931,N_2881,N_2853);
nor U2932 (N_2932,N_2920,N_2863);
and U2933 (N_2933,N_2873,N_2882);
and U2934 (N_2934,N_2918,N_2860);
and U2935 (N_2935,N_2895,N_2859);
or U2936 (N_2936,N_2878,N_2884);
or U2937 (N_2937,N_2923,N_2915);
or U2938 (N_2938,N_2914,N_2885);
or U2939 (N_2939,N_2850,N_2887);
nand U2940 (N_2940,N_2922,N_2909);
nor U2941 (N_2941,N_2869,N_2892);
or U2942 (N_2942,N_2874,N_2867);
nand U2943 (N_2943,N_2900,N_2907);
nand U2944 (N_2944,N_2910,N_2855);
nand U2945 (N_2945,N_2888,N_2890);
nor U2946 (N_2946,N_2899,N_2865);
or U2947 (N_2947,N_2877,N_2921);
nor U2948 (N_2948,N_2871,N_2893);
xnor U2949 (N_2949,N_2919,N_2854);
nand U2950 (N_2950,N_2917,N_2913);
xnor U2951 (N_2951,N_2880,N_2852);
or U2952 (N_2952,N_2896,N_2856);
and U2953 (N_2953,N_2886,N_2875);
or U2954 (N_2954,N_2906,N_2851);
nand U2955 (N_2955,N_2901,N_2870);
nor U2956 (N_2956,N_2897,N_2924);
and U2957 (N_2957,N_2858,N_2916);
nor U2958 (N_2958,N_2864,N_2903);
or U2959 (N_2959,N_2905,N_2912);
or U2960 (N_2960,N_2862,N_2904);
nand U2961 (N_2961,N_2883,N_2898);
and U2962 (N_2962,N_2868,N_2876);
nand U2963 (N_2963,N_2918,N_2851);
or U2964 (N_2964,N_2921,N_2918);
nor U2965 (N_2965,N_2920,N_2887);
and U2966 (N_2966,N_2911,N_2870);
or U2967 (N_2967,N_2869,N_2886);
or U2968 (N_2968,N_2893,N_2882);
nor U2969 (N_2969,N_2889,N_2897);
or U2970 (N_2970,N_2897,N_2894);
xnor U2971 (N_2971,N_2859,N_2873);
xnor U2972 (N_2972,N_2852,N_2865);
or U2973 (N_2973,N_2867,N_2871);
nor U2974 (N_2974,N_2879,N_2877);
or U2975 (N_2975,N_2868,N_2883);
or U2976 (N_2976,N_2887,N_2924);
nor U2977 (N_2977,N_2878,N_2858);
or U2978 (N_2978,N_2872,N_2921);
and U2979 (N_2979,N_2864,N_2908);
or U2980 (N_2980,N_2917,N_2865);
nand U2981 (N_2981,N_2920,N_2877);
and U2982 (N_2982,N_2924,N_2857);
and U2983 (N_2983,N_2852,N_2888);
and U2984 (N_2984,N_2867,N_2855);
and U2985 (N_2985,N_2870,N_2866);
xnor U2986 (N_2986,N_2866,N_2894);
nand U2987 (N_2987,N_2869,N_2885);
nand U2988 (N_2988,N_2855,N_2895);
and U2989 (N_2989,N_2852,N_2872);
or U2990 (N_2990,N_2893,N_2908);
nand U2991 (N_2991,N_2907,N_2861);
nor U2992 (N_2992,N_2913,N_2922);
and U2993 (N_2993,N_2912,N_2898);
or U2994 (N_2994,N_2904,N_2922);
nand U2995 (N_2995,N_2869,N_2859);
nor U2996 (N_2996,N_2917,N_2856);
and U2997 (N_2997,N_2870,N_2898);
nand U2998 (N_2998,N_2896,N_2871);
and U2999 (N_2999,N_2919,N_2866);
nand UO_0 (O_0,N_2951,N_2946);
or UO_1 (O_1,N_2995,N_2947);
nand UO_2 (O_2,N_2935,N_2934);
xnor UO_3 (O_3,N_2962,N_2939);
and UO_4 (O_4,N_2986,N_2966);
and UO_5 (O_5,N_2964,N_2987);
xor UO_6 (O_6,N_2925,N_2977);
xor UO_7 (O_7,N_2990,N_2950);
nand UO_8 (O_8,N_2994,N_2974);
nor UO_9 (O_9,N_2968,N_2989);
nor UO_10 (O_10,N_2953,N_2996);
nor UO_11 (O_11,N_2971,N_2973);
nand UO_12 (O_12,N_2937,N_2969);
nand UO_13 (O_13,N_2948,N_2941);
xnor UO_14 (O_14,N_2967,N_2954);
xnor UO_15 (O_15,N_2938,N_2979);
nand UO_16 (O_16,N_2943,N_2997);
nor UO_17 (O_17,N_2963,N_2982);
nor UO_18 (O_18,N_2958,N_2988);
nor UO_19 (O_19,N_2981,N_2932);
and UO_20 (O_20,N_2940,N_2959);
nor UO_21 (O_21,N_2972,N_2985);
and UO_22 (O_22,N_2945,N_2984);
nand UO_23 (O_23,N_2949,N_2992);
and UO_24 (O_24,N_2926,N_2999);
nor UO_25 (O_25,N_2961,N_2993);
and UO_26 (O_26,N_2975,N_2976);
xnor UO_27 (O_27,N_2991,N_2956);
nand UO_28 (O_28,N_2930,N_2952);
nor UO_29 (O_29,N_2998,N_2978);
nand UO_30 (O_30,N_2928,N_2927);
nand UO_31 (O_31,N_2957,N_2960);
and UO_32 (O_32,N_2980,N_2970);
and UO_33 (O_33,N_2965,N_2933);
or UO_34 (O_34,N_2931,N_2983);
nor UO_35 (O_35,N_2942,N_2929);
nor UO_36 (O_36,N_2936,N_2955);
or UO_37 (O_37,N_2944,N_2948);
nand UO_38 (O_38,N_2978,N_2946);
and UO_39 (O_39,N_2966,N_2934);
nand UO_40 (O_40,N_2928,N_2944);
nor UO_41 (O_41,N_2930,N_2994);
nand UO_42 (O_42,N_2986,N_2976);
nor UO_43 (O_43,N_2995,N_2992);
xnor UO_44 (O_44,N_2990,N_2997);
nand UO_45 (O_45,N_2993,N_2962);
and UO_46 (O_46,N_2968,N_2960);
xor UO_47 (O_47,N_2953,N_2968);
xor UO_48 (O_48,N_2973,N_2934);
nor UO_49 (O_49,N_2962,N_2956);
nand UO_50 (O_50,N_2966,N_2980);
and UO_51 (O_51,N_2935,N_2940);
nand UO_52 (O_52,N_2996,N_2990);
nor UO_53 (O_53,N_2988,N_2998);
nor UO_54 (O_54,N_2936,N_2961);
nand UO_55 (O_55,N_2993,N_2983);
or UO_56 (O_56,N_2933,N_2946);
or UO_57 (O_57,N_2990,N_2946);
or UO_58 (O_58,N_2954,N_2972);
nand UO_59 (O_59,N_2958,N_2959);
and UO_60 (O_60,N_2990,N_2999);
nand UO_61 (O_61,N_2995,N_2984);
or UO_62 (O_62,N_2951,N_2967);
and UO_63 (O_63,N_2941,N_2931);
and UO_64 (O_64,N_2984,N_2994);
or UO_65 (O_65,N_2967,N_2955);
nor UO_66 (O_66,N_2941,N_2946);
nand UO_67 (O_67,N_2997,N_2927);
or UO_68 (O_68,N_2957,N_2983);
and UO_69 (O_69,N_2927,N_2931);
nor UO_70 (O_70,N_2929,N_2975);
and UO_71 (O_71,N_2996,N_2992);
or UO_72 (O_72,N_2998,N_2932);
and UO_73 (O_73,N_2943,N_2947);
nor UO_74 (O_74,N_2986,N_2925);
nor UO_75 (O_75,N_2952,N_2986);
nor UO_76 (O_76,N_2966,N_2990);
nand UO_77 (O_77,N_2986,N_2997);
or UO_78 (O_78,N_2995,N_2965);
or UO_79 (O_79,N_2971,N_2952);
or UO_80 (O_80,N_2966,N_2970);
or UO_81 (O_81,N_2990,N_2930);
nand UO_82 (O_82,N_2948,N_2979);
or UO_83 (O_83,N_2946,N_2959);
and UO_84 (O_84,N_2990,N_2949);
nor UO_85 (O_85,N_2927,N_2952);
nand UO_86 (O_86,N_2934,N_2970);
nand UO_87 (O_87,N_2957,N_2958);
nand UO_88 (O_88,N_2936,N_2967);
nand UO_89 (O_89,N_2993,N_2939);
nor UO_90 (O_90,N_2962,N_2938);
or UO_91 (O_91,N_2928,N_2949);
or UO_92 (O_92,N_2956,N_2975);
nor UO_93 (O_93,N_2966,N_2964);
nor UO_94 (O_94,N_2937,N_2950);
nand UO_95 (O_95,N_2945,N_2951);
and UO_96 (O_96,N_2936,N_2988);
nor UO_97 (O_97,N_2974,N_2925);
xor UO_98 (O_98,N_2945,N_2998);
or UO_99 (O_99,N_2936,N_2933);
or UO_100 (O_100,N_2972,N_2970);
or UO_101 (O_101,N_2959,N_2994);
nor UO_102 (O_102,N_2958,N_2947);
and UO_103 (O_103,N_2981,N_2985);
nor UO_104 (O_104,N_2990,N_2978);
and UO_105 (O_105,N_2987,N_2975);
or UO_106 (O_106,N_2952,N_2977);
nand UO_107 (O_107,N_2952,N_2979);
nor UO_108 (O_108,N_2959,N_2939);
nor UO_109 (O_109,N_2961,N_2991);
or UO_110 (O_110,N_2994,N_2989);
or UO_111 (O_111,N_2981,N_2970);
and UO_112 (O_112,N_2988,N_2944);
nand UO_113 (O_113,N_2996,N_2975);
nor UO_114 (O_114,N_2971,N_2926);
nand UO_115 (O_115,N_2998,N_2985);
or UO_116 (O_116,N_2975,N_2952);
nand UO_117 (O_117,N_2944,N_2950);
nand UO_118 (O_118,N_2945,N_2993);
or UO_119 (O_119,N_2933,N_2925);
or UO_120 (O_120,N_2989,N_2946);
nor UO_121 (O_121,N_2926,N_2965);
and UO_122 (O_122,N_2933,N_2954);
and UO_123 (O_123,N_2959,N_2966);
and UO_124 (O_124,N_2986,N_2955);
or UO_125 (O_125,N_2931,N_2981);
and UO_126 (O_126,N_2977,N_2939);
nand UO_127 (O_127,N_2950,N_2966);
and UO_128 (O_128,N_2941,N_2952);
nand UO_129 (O_129,N_2974,N_2931);
nor UO_130 (O_130,N_2988,N_2932);
and UO_131 (O_131,N_2989,N_2987);
nor UO_132 (O_132,N_2968,N_2942);
and UO_133 (O_133,N_2960,N_2927);
nor UO_134 (O_134,N_2928,N_2968);
nand UO_135 (O_135,N_2966,N_2953);
and UO_136 (O_136,N_2955,N_2992);
nand UO_137 (O_137,N_2935,N_2968);
and UO_138 (O_138,N_2978,N_2930);
or UO_139 (O_139,N_2938,N_2927);
or UO_140 (O_140,N_2955,N_2960);
xnor UO_141 (O_141,N_2945,N_2937);
nor UO_142 (O_142,N_2981,N_2933);
or UO_143 (O_143,N_2985,N_2995);
nand UO_144 (O_144,N_2955,N_2987);
nand UO_145 (O_145,N_2989,N_2931);
or UO_146 (O_146,N_2999,N_2945);
or UO_147 (O_147,N_2992,N_2998);
nand UO_148 (O_148,N_2996,N_2969);
nor UO_149 (O_149,N_2982,N_2926);
nand UO_150 (O_150,N_2978,N_2970);
nor UO_151 (O_151,N_2998,N_2946);
or UO_152 (O_152,N_2953,N_2981);
or UO_153 (O_153,N_2973,N_2926);
and UO_154 (O_154,N_2980,N_2979);
and UO_155 (O_155,N_2991,N_2954);
or UO_156 (O_156,N_2940,N_2948);
xor UO_157 (O_157,N_2966,N_2928);
and UO_158 (O_158,N_2945,N_2932);
or UO_159 (O_159,N_2936,N_2969);
or UO_160 (O_160,N_2949,N_2935);
nand UO_161 (O_161,N_2986,N_2974);
nor UO_162 (O_162,N_2964,N_2995);
xor UO_163 (O_163,N_2968,N_2955);
nand UO_164 (O_164,N_2989,N_2947);
and UO_165 (O_165,N_2966,N_2973);
xor UO_166 (O_166,N_2960,N_2947);
nand UO_167 (O_167,N_2933,N_2971);
nand UO_168 (O_168,N_2968,N_2986);
or UO_169 (O_169,N_2995,N_2999);
nor UO_170 (O_170,N_2972,N_2986);
or UO_171 (O_171,N_2995,N_2974);
nand UO_172 (O_172,N_2952,N_2989);
or UO_173 (O_173,N_2949,N_2986);
and UO_174 (O_174,N_2962,N_2930);
xnor UO_175 (O_175,N_2930,N_2993);
and UO_176 (O_176,N_2935,N_2976);
or UO_177 (O_177,N_2968,N_2950);
nand UO_178 (O_178,N_2984,N_2971);
nand UO_179 (O_179,N_2966,N_2954);
or UO_180 (O_180,N_2937,N_2942);
and UO_181 (O_181,N_2967,N_2986);
nand UO_182 (O_182,N_2944,N_2939);
or UO_183 (O_183,N_2937,N_2925);
nor UO_184 (O_184,N_2992,N_2956);
or UO_185 (O_185,N_2956,N_2946);
xnor UO_186 (O_186,N_2968,N_2940);
nand UO_187 (O_187,N_2929,N_2932);
nor UO_188 (O_188,N_2943,N_2992);
and UO_189 (O_189,N_2996,N_2982);
nor UO_190 (O_190,N_2951,N_2925);
or UO_191 (O_191,N_2996,N_2943);
and UO_192 (O_192,N_2961,N_2962);
nand UO_193 (O_193,N_2986,N_2975);
or UO_194 (O_194,N_2958,N_2970);
nand UO_195 (O_195,N_2979,N_2967);
or UO_196 (O_196,N_2949,N_2987);
nor UO_197 (O_197,N_2942,N_2975);
nor UO_198 (O_198,N_2980,N_2964);
nor UO_199 (O_199,N_2927,N_2954);
nand UO_200 (O_200,N_2970,N_2960);
or UO_201 (O_201,N_2996,N_2965);
nor UO_202 (O_202,N_2992,N_2960);
nand UO_203 (O_203,N_2953,N_2988);
xor UO_204 (O_204,N_2946,N_2929);
nor UO_205 (O_205,N_2998,N_2973);
or UO_206 (O_206,N_2992,N_2988);
xor UO_207 (O_207,N_2937,N_2994);
xnor UO_208 (O_208,N_2983,N_2946);
nor UO_209 (O_209,N_2939,N_2957);
xnor UO_210 (O_210,N_2999,N_2981);
or UO_211 (O_211,N_2961,N_2971);
xnor UO_212 (O_212,N_2979,N_2996);
or UO_213 (O_213,N_2943,N_2950);
nand UO_214 (O_214,N_2989,N_2933);
nor UO_215 (O_215,N_2940,N_2969);
or UO_216 (O_216,N_2952,N_2994);
nand UO_217 (O_217,N_2967,N_2989);
or UO_218 (O_218,N_2978,N_2983);
xor UO_219 (O_219,N_2972,N_2958);
or UO_220 (O_220,N_2965,N_2964);
nand UO_221 (O_221,N_2953,N_2994);
and UO_222 (O_222,N_2976,N_2951);
nand UO_223 (O_223,N_2995,N_2940);
and UO_224 (O_224,N_2998,N_2970);
nor UO_225 (O_225,N_2960,N_2979);
nand UO_226 (O_226,N_2961,N_2941);
and UO_227 (O_227,N_2972,N_2993);
or UO_228 (O_228,N_2943,N_2931);
nor UO_229 (O_229,N_2989,N_2983);
or UO_230 (O_230,N_2937,N_2960);
and UO_231 (O_231,N_2958,N_2939);
nor UO_232 (O_232,N_2968,N_2996);
nor UO_233 (O_233,N_2961,N_2986);
nand UO_234 (O_234,N_2928,N_2960);
or UO_235 (O_235,N_2926,N_2953);
nand UO_236 (O_236,N_2977,N_2976);
and UO_237 (O_237,N_2956,N_2981);
xnor UO_238 (O_238,N_2971,N_2985);
and UO_239 (O_239,N_2990,N_2973);
nor UO_240 (O_240,N_2940,N_2954);
and UO_241 (O_241,N_2971,N_2969);
and UO_242 (O_242,N_2968,N_2983);
nand UO_243 (O_243,N_2995,N_2928);
and UO_244 (O_244,N_2925,N_2998);
xnor UO_245 (O_245,N_2951,N_2928);
or UO_246 (O_246,N_2978,N_2962);
nor UO_247 (O_247,N_2995,N_2962);
and UO_248 (O_248,N_2925,N_2989);
nor UO_249 (O_249,N_2961,N_2943);
xnor UO_250 (O_250,N_2925,N_2983);
or UO_251 (O_251,N_2937,N_2999);
nand UO_252 (O_252,N_2955,N_2971);
nor UO_253 (O_253,N_2956,N_2994);
and UO_254 (O_254,N_2953,N_2949);
and UO_255 (O_255,N_2977,N_2991);
or UO_256 (O_256,N_2987,N_2969);
nand UO_257 (O_257,N_2975,N_2989);
nor UO_258 (O_258,N_2992,N_2967);
nand UO_259 (O_259,N_2998,N_2999);
nand UO_260 (O_260,N_2932,N_2980);
or UO_261 (O_261,N_2956,N_2969);
nor UO_262 (O_262,N_2994,N_2927);
or UO_263 (O_263,N_2935,N_2984);
nor UO_264 (O_264,N_2984,N_2998);
nor UO_265 (O_265,N_2942,N_2939);
and UO_266 (O_266,N_2979,N_2951);
xor UO_267 (O_267,N_2938,N_2944);
nor UO_268 (O_268,N_2981,N_2963);
nor UO_269 (O_269,N_2926,N_2978);
nand UO_270 (O_270,N_2962,N_2946);
xor UO_271 (O_271,N_2928,N_2990);
and UO_272 (O_272,N_2970,N_2946);
and UO_273 (O_273,N_2982,N_2953);
or UO_274 (O_274,N_2995,N_2946);
and UO_275 (O_275,N_2996,N_2967);
xnor UO_276 (O_276,N_2941,N_2942);
nand UO_277 (O_277,N_2955,N_2930);
nand UO_278 (O_278,N_2938,N_2929);
nand UO_279 (O_279,N_2971,N_2945);
nor UO_280 (O_280,N_2986,N_2957);
nor UO_281 (O_281,N_2954,N_2988);
xnor UO_282 (O_282,N_2943,N_2971);
nor UO_283 (O_283,N_2950,N_2985);
nand UO_284 (O_284,N_2933,N_2977);
or UO_285 (O_285,N_2946,N_2955);
xor UO_286 (O_286,N_2954,N_2999);
and UO_287 (O_287,N_2952,N_2945);
nand UO_288 (O_288,N_2949,N_2929);
xor UO_289 (O_289,N_2974,N_2966);
and UO_290 (O_290,N_2947,N_2981);
xnor UO_291 (O_291,N_2939,N_2938);
nand UO_292 (O_292,N_2934,N_2942);
or UO_293 (O_293,N_2991,N_2925);
nor UO_294 (O_294,N_2930,N_2937);
nand UO_295 (O_295,N_2927,N_2962);
or UO_296 (O_296,N_2988,N_2960);
xnor UO_297 (O_297,N_2926,N_2962);
nor UO_298 (O_298,N_2952,N_2988);
nand UO_299 (O_299,N_2983,N_2949);
nor UO_300 (O_300,N_2953,N_2936);
and UO_301 (O_301,N_2953,N_2989);
xor UO_302 (O_302,N_2934,N_2957);
nor UO_303 (O_303,N_2928,N_2988);
nor UO_304 (O_304,N_2955,N_2998);
nor UO_305 (O_305,N_2947,N_2965);
or UO_306 (O_306,N_2976,N_2970);
nand UO_307 (O_307,N_2967,N_2956);
nor UO_308 (O_308,N_2929,N_2952);
and UO_309 (O_309,N_2928,N_2978);
nand UO_310 (O_310,N_2969,N_2976);
or UO_311 (O_311,N_2927,N_2991);
or UO_312 (O_312,N_2929,N_2925);
or UO_313 (O_313,N_2999,N_2982);
nor UO_314 (O_314,N_2963,N_2978);
and UO_315 (O_315,N_2999,N_2959);
nor UO_316 (O_316,N_2970,N_2956);
or UO_317 (O_317,N_2954,N_2971);
or UO_318 (O_318,N_2929,N_2955);
or UO_319 (O_319,N_2979,N_2972);
and UO_320 (O_320,N_2940,N_2965);
nor UO_321 (O_321,N_2974,N_2973);
and UO_322 (O_322,N_2976,N_2988);
or UO_323 (O_323,N_2995,N_2935);
or UO_324 (O_324,N_2995,N_2987);
or UO_325 (O_325,N_2978,N_2995);
xor UO_326 (O_326,N_2937,N_2989);
nor UO_327 (O_327,N_2932,N_2958);
nand UO_328 (O_328,N_2991,N_2990);
nand UO_329 (O_329,N_2973,N_2970);
or UO_330 (O_330,N_2960,N_2997);
nor UO_331 (O_331,N_2929,N_2976);
or UO_332 (O_332,N_2977,N_2926);
or UO_333 (O_333,N_2958,N_2951);
and UO_334 (O_334,N_2957,N_2925);
and UO_335 (O_335,N_2976,N_2983);
and UO_336 (O_336,N_2971,N_2950);
nand UO_337 (O_337,N_2954,N_2969);
or UO_338 (O_338,N_2955,N_2926);
nor UO_339 (O_339,N_2929,N_2956);
nor UO_340 (O_340,N_2983,N_2969);
nand UO_341 (O_341,N_2984,N_2951);
and UO_342 (O_342,N_2955,N_2959);
xor UO_343 (O_343,N_2974,N_2981);
or UO_344 (O_344,N_2934,N_2981);
or UO_345 (O_345,N_2982,N_2992);
xor UO_346 (O_346,N_2964,N_2981);
or UO_347 (O_347,N_2965,N_2968);
and UO_348 (O_348,N_2982,N_2941);
nand UO_349 (O_349,N_2947,N_2926);
and UO_350 (O_350,N_2951,N_2953);
nor UO_351 (O_351,N_2926,N_2937);
or UO_352 (O_352,N_2939,N_2946);
nor UO_353 (O_353,N_2952,N_2963);
nor UO_354 (O_354,N_2925,N_2987);
xnor UO_355 (O_355,N_2949,N_2952);
and UO_356 (O_356,N_2973,N_2987);
or UO_357 (O_357,N_2958,N_2953);
xnor UO_358 (O_358,N_2987,N_2929);
or UO_359 (O_359,N_2970,N_2937);
or UO_360 (O_360,N_2952,N_2951);
nor UO_361 (O_361,N_2933,N_2972);
and UO_362 (O_362,N_2960,N_2986);
nor UO_363 (O_363,N_2941,N_2945);
nand UO_364 (O_364,N_2984,N_2943);
and UO_365 (O_365,N_2933,N_2983);
or UO_366 (O_366,N_2992,N_2972);
and UO_367 (O_367,N_2947,N_2998);
nor UO_368 (O_368,N_2988,N_2957);
or UO_369 (O_369,N_2954,N_2981);
nor UO_370 (O_370,N_2992,N_2997);
and UO_371 (O_371,N_2977,N_2928);
nor UO_372 (O_372,N_2943,N_2989);
or UO_373 (O_373,N_2991,N_2940);
and UO_374 (O_374,N_2940,N_2950);
nand UO_375 (O_375,N_2953,N_2950);
or UO_376 (O_376,N_2996,N_2945);
or UO_377 (O_377,N_2962,N_2963);
nor UO_378 (O_378,N_2947,N_2985);
nor UO_379 (O_379,N_2939,N_2948);
and UO_380 (O_380,N_2993,N_2947);
and UO_381 (O_381,N_2997,N_2995);
nor UO_382 (O_382,N_2951,N_2988);
and UO_383 (O_383,N_2991,N_2970);
nand UO_384 (O_384,N_2944,N_2987);
and UO_385 (O_385,N_2997,N_2980);
nor UO_386 (O_386,N_2940,N_2996);
or UO_387 (O_387,N_2986,N_2931);
nor UO_388 (O_388,N_2940,N_2926);
nor UO_389 (O_389,N_2985,N_2927);
nor UO_390 (O_390,N_2939,N_2981);
nand UO_391 (O_391,N_2941,N_2986);
xor UO_392 (O_392,N_2973,N_2948);
and UO_393 (O_393,N_2926,N_2966);
nand UO_394 (O_394,N_2987,N_2963);
xnor UO_395 (O_395,N_2963,N_2941);
and UO_396 (O_396,N_2972,N_2982);
xnor UO_397 (O_397,N_2970,N_2929);
nand UO_398 (O_398,N_2995,N_2952);
nor UO_399 (O_399,N_2928,N_2963);
nand UO_400 (O_400,N_2983,N_2979);
nand UO_401 (O_401,N_2984,N_2973);
or UO_402 (O_402,N_2977,N_2988);
and UO_403 (O_403,N_2970,N_2935);
or UO_404 (O_404,N_2933,N_2999);
or UO_405 (O_405,N_2995,N_2958);
and UO_406 (O_406,N_2939,N_2954);
and UO_407 (O_407,N_2927,N_2945);
nor UO_408 (O_408,N_2982,N_2930);
nand UO_409 (O_409,N_2961,N_2949);
nand UO_410 (O_410,N_2969,N_2968);
and UO_411 (O_411,N_2938,N_2989);
and UO_412 (O_412,N_2989,N_2934);
and UO_413 (O_413,N_2997,N_2947);
nor UO_414 (O_414,N_2928,N_2931);
xnor UO_415 (O_415,N_2939,N_2991);
nor UO_416 (O_416,N_2971,N_2931);
and UO_417 (O_417,N_2941,N_2985);
nor UO_418 (O_418,N_2991,N_2950);
and UO_419 (O_419,N_2937,N_2946);
or UO_420 (O_420,N_2940,N_2979);
nor UO_421 (O_421,N_2926,N_2992);
and UO_422 (O_422,N_2927,N_2970);
nor UO_423 (O_423,N_2958,N_2992);
and UO_424 (O_424,N_2996,N_2927);
xor UO_425 (O_425,N_2964,N_2955);
nand UO_426 (O_426,N_2997,N_2931);
nand UO_427 (O_427,N_2979,N_2939);
or UO_428 (O_428,N_2973,N_2931);
nor UO_429 (O_429,N_2973,N_2983);
or UO_430 (O_430,N_2983,N_2997);
and UO_431 (O_431,N_2957,N_2932);
or UO_432 (O_432,N_2963,N_2953);
nor UO_433 (O_433,N_2928,N_2925);
nand UO_434 (O_434,N_2982,N_2959);
xnor UO_435 (O_435,N_2936,N_2945);
or UO_436 (O_436,N_2959,N_2972);
nor UO_437 (O_437,N_2981,N_2935);
and UO_438 (O_438,N_2959,N_2984);
or UO_439 (O_439,N_2980,N_2995);
xor UO_440 (O_440,N_2978,N_2945);
or UO_441 (O_441,N_2977,N_2955);
nand UO_442 (O_442,N_2954,N_2961);
nand UO_443 (O_443,N_2951,N_2998);
and UO_444 (O_444,N_2948,N_2970);
nand UO_445 (O_445,N_2948,N_2965);
nand UO_446 (O_446,N_2962,N_2999);
or UO_447 (O_447,N_2931,N_2956);
nand UO_448 (O_448,N_2984,N_2950);
or UO_449 (O_449,N_2990,N_2960);
or UO_450 (O_450,N_2927,N_2999);
xnor UO_451 (O_451,N_2936,N_2930);
or UO_452 (O_452,N_2944,N_2926);
or UO_453 (O_453,N_2987,N_2999);
nand UO_454 (O_454,N_2998,N_2954);
or UO_455 (O_455,N_2978,N_2947);
or UO_456 (O_456,N_2970,N_2957);
and UO_457 (O_457,N_2935,N_2989);
or UO_458 (O_458,N_2951,N_2974);
or UO_459 (O_459,N_2969,N_2995);
xnor UO_460 (O_460,N_2936,N_2942);
nand UO_461 (O_461,N_2970,N_2932);
nor UO_462 (O_462,N_2961,N_2999);
or UO_463 (O_463,N_2929,N_2995);
nor UO_464 (O_464,N_2987,N_2948);
nor UO_465 (O_465,N_2927,N_2977);
or UO_466 (O_466,N_2964,N_2984);
or UO_467 (O_467,N_2994,N_2958);
and UO_468 (O_468,N_2980,N_2936);
or UO_469 (O_469,N_2928,N_2936);
or UO_470 (O_470,N_2950,N_2963);
nand UO_471 (O_471,N_2942,N_2932);
and UO_472 (O_472,N_2998,N_2989);
xor UO_473 (O_473,N_2989,N_2976);
xnor UO_474 (O_474,N_2995,N_2933);
nor UO_475 (O_475,N_2936,N_2981);
nand UO_476 (O_476,N_2970,N_2952);
or UO_477 (O_477,N_2981,N_2973);
and UO_478 (O_478,N_2940,N_2974);
nor UO_479 (O_479,N_2981,N_2978);
or UO_480 (O_480,N_2972,N_2957);
nor UO_481 (O_481,N_2931,N_2952);
xor UO_482 (O_482,N_2947,N_2940);
or UO_483 (O_483,N_2941,N_2975);
nor UO_484 (O_484,N_2974,N_2976);
or UO_485 (O_485,N_2971,N_2946);
or UO_486 (O_486,N_2936,N_2974);
nor UO_487 (O_487,N_2991,N_2998);
and UO_488 (O_488,N_2977,N_2948);
or UO_489 (O_489,N_2975,N_2951);
xnor UO_490 (O_490,N_2986,N_2970);
and UO_491 (O_491,N_2965,N_2966);
nor UO_492 (O_492,N_2937,N_2940);
nor UO_493 (O_493,N_2989,N_2979);
nor UO_494 (O_494,N_2926,N_2979);
and UO_495 (O_495,N_2995,N_2942);
or UO_496 (O_496,N_2940,N_2932);
and UO_497 (O_497,N_2934,N_2962);
and UO_498 (O_498,N_2936,N_2947);
xor UO_499 (O_499,N_2946,N_2963);
endmodule