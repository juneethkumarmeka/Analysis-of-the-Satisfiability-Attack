module basic_500_3000_500_4_levels_5xor_1(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
nand U0 (N_0,In_83,In_384);
nor U1 (N_1,In_10,In_354);
nor U2 (N_2,In_357,In_163);
nand U3 (N_3,In_336,In_189);
nor U4 (N_4,In_402,In_362);
nor U5 (N_5,In_33,In_167);
and U6 (N_6,In_447,In_274);
and U7 (N_7,In_233,In_8);
or U8 (N_8,In_333,In_186);
or U9 (N_9,In_289,In_58);
xnor U10 (N_10,In_2,In_37);
and U11 (N_11,In_419,In_92);
or U12 (N_12,In_240,In_475);
and U13 (N_13,In_398,In_40);
and U14 (N_14,In_316,In_353);
nor U15 (N_15,In_0,In_349);
nor U16 (N_16,In_94,In_467);
or U17 (N_17,In_297,In_466);
xor U18 (N_18,In_25,In_389);
or U19 (N_19,In_247,In_110);
and U20 (N_20,In_174,In_457);
nand U21 (N_21,In_442,In_304);
xnor U22 (N_22,In_56,In_373);
nor U23 (N_23,In_77,In_291);
and U24 (N_24,In_99,In_427);
xor U25 (N_25,In_250,In_190);
or U26 (N_26,In_489,In_301);
xnor U27 (N_27,In_95,In_50);
nor U28 (N_28,In_148,In_135);
or U29 (N_29,In_175,In_363);
nor U30 (N_30,In_343,In_424);
or U31 (N_31,In_234,In_416);
or U32 (N_32,In_64,In_71);
xor U33 (N_33,In_111,In_317);
and U34 (N_34,In_196,In_144);
nor U35 (N_35,In_246,In_407);
nor U36 (N_36,In_391,In_472);
nor U37 (N_37,In_139,In_166);
nand U38 (N_38,In_367,In_102);
nand U39 (N_39,In_216,In_378);
nor U40 (N_40,In_370,In_218);
nor U41 (N_41,In_118,In_114);
or U42 (N_42,In_371,In_19);
and U43 (N_43,In_123,In_21);
or U44 (N_44,In_486,In_411);
nor U45 (N_45,In_68,In_23);
or U46 (N_46,In_75,In_482);
xor U47 (N_47,In_397,In_62);
and U48 (N_48,In_57,In_168);
xor U49 (N_49,In_206,In_326);
nand U50 (N_50,In_93,In_458);
or U51 (N_51,In_59,In_129);
and U52 (N_52,In_421,In_41);
and U53 (N_53,In_409,In_382);
and U54 (N_54,In_280,In_481);
and U55 (N_55,In_191,In_219);
or U56 (N_56,In_209,In_236);
or U57 (N_57,In_82,In_112);
and U58 (N_58,In_300,In_169);
nor U59 (N_59,In_42,In_423);
xor U60 (N_60,In_224,In_22);
nor U61 (N_61,In_446,In_51);
nor U62 (N_62,In_201,In_263);
or U63 (N_63,In_369,In_310);
and U64 (N_64,In_499,In_451);
nand U65 (N_65,In_393,In_117);
or U66 (N_66,In_115,In_335);
nand U67 (N_67,In_435,In_98);
nor U68 (N_68,In_249,In_330);
or U69 (N_69,In_165,In_376);
and U70 (N_70,In_264,In_328);
xnor U71 (N_71,In_130,In_368);
nand U72 (N_72,In_355,In_151);
nor U73 (N_73,In_388,In_154);
nand U74 (N_74,In_313,In_146);
xnor U75 (N_75,In_387,In_74);
nand U76 (N_76,In_90,In_431);
or U77 (N_77,In_137,In_78);
nand U78 (N_78,In_65,In_244);
and U79 (N_79,In_223,In_32);
nand U80 (N_80,In_484,In_488);
nand U81 (N_81,In_221,In_436);
and U82 (N_82,In_403,In_177);
nand U83 (N_83,In_76,In_284);
nand U84 (N_84,In_293,In_122);
nand U85 (N_85,In_243,In_286);
or U86 (N_86,In_379,In_360);
nand U87 (N_87,In_453,In_205);
and U88 (N_88,In_106,In_456);
or U89 (N_89,In_81,In_5);
nand U90 (N_90,In_296,In_452);
nand U91 (N_91,In_157,In_3);
xnor U92 (N_92,In_470,In_277);
xnor U93 (N_93,In_437,In_36);
or U94 (N_94,In_420,In_31);
nand U95 (N_95,In_12,In_422);
and U96 (N_96,In_17,In_131);
xnor U97 (N_97,In_63,In_107);
and U98 (N_98,In_152,In_198);
nand U99 (N_99,In_432,In_292);
nor U100 (N_100,In_268,In_39);
or U101 (N_101,In_390,In_288);
xnor U102 (N_102,In_322,In_430);
nor U103 (N_103,In_105,In_260);
or U104 (N_104,In_394,In_49);
nand U105 (N_105,In_460,In_171);
nor U106 (N_106,In_433,In_60);
nand U107 (N_107,In_235,In_66);
nand U108 (N_108,In_396,In_479);
or U109 (N_109,In_321,In_187);
nand U110 (N_110,In_279,In_256);
nor U111 (N_111,In_231,In_126);
nand U112 (N_112,In_241,In_327);
nor U113 (N_113,In_121,In_359);
and U114 (N_114,In_113,In_338);
nand U115 (N_115,In_104,In_444);
nand U116 (N_116,In_347,In_340);
and U117 (N_117,In_132,In_119);
nor U118 (N_118,In_438,In_401);
xnor U119 (N_119,In_140,In_381);
or U120 (N_120,In_232,In_54);
and U121 (N_121,In_298,In_459);
or U122 (N_122,In_332,In_414);
nor U123 (N_123,In_358,In_375);
nand U124 (N_124,In_141,In_125);
nor U125 (N_125,In_30,In_155);
or U126 (N_126,In_434,In_302);
nor U127 (N_127,In_15,In_120);
and U128 (N_128,In_348,In_9);
and U129 (N_129,In_342,In_67);
xnor U130 (N_130,In_366,In_440);
or U131 (N_131,In_226,In_73);
and U132 (N_132,In_473,In_46);
xor U133 (N_133,In_116,In_303);
and U134 (N_134,In_228,In_188);
nand U135 (N_135,In_283,In_266);
nor U136 (N_136,In_295,In_275);
or U137 (N_137,In_143,In_213);
nor U138 (N_138,In_305,In_461);
and U139 (N_139,In_487,In_24);
xor U140 (N_140,In_257,In_197);
xnor U141 (N_141,In_84,In_281);
nand U142 (N_142,In_43,In_173);
and U143 (N_143,In_346,In_153);
nor U144 (N_144,In_399,In_285);
and U145 (N_145,In_429,In_331);
xnor U146 (N_146,In_47,In_109);
nand U147 (N_147,In_306,In_267);
and U148 (N_148,In_127,In_372);
or U149 (N_149,In_194,In_253);
and U150 (N_150,In_408,In_45);
nor U151 (N_151,In_69,In_449);
nand U152 (N_152,In_465,In_149);
nor U153 (N_153,In_133,In_1);
nor U154 (N_154,In_242,In_160);
or U155 (N_155,In_377,In_150);
nor U156 (N_156,In_178,In_225);
and U157 (N_157,In_20,In_491);
nor U158 (N_158,In_195,In_28);
and U159 (N_159,In_34,In_276);
and U160 (N_160,In_245,In_392);
nor U161 (N_161,In_252,In_320);
and U162 (N_162,In_202,In_254);
nor U163 (N_163,In_258,In_294);
nand U164 (N_164,In_162,In_450);
nand U165 (N_165,In_383,In_352);
nand U166 (N_166,In_238,In_255);
nor U167 (N_167,In_183,In_380);
and U168 (N_168,In_159,In_485);
and U169 (N_169,In_334,In_490);
nor U170 (N_170,In_478,In_103);
nor U171 (N_171,In_192,In_350);
and U172 (N_172,In_441,In_464);
and U173 (N_173,In_483,In_147);
and U174 (N_174,In_18,In_287);
xor U175 (N_175,In_425,In_220);
nor U176 (N_176,In_469,In_138);
nand U177 (N_177,In_455,In_315);
or U178 (N_178,In_361,In_272);
xor U179 (N_179,In_214,In_428);
nor U180 (N_180,In_417,In_182);
or U181 (N_181,In_345,In_229);
nor U182 (N_182,In_323,In_299);
nand U183 (N_183,In_471,In_443);
and U184 (N_184,In_124,In_44);
nand U185 (N_185,In_200,In_204);
xor U186 (N_186,In_38,In_307);
nand U187 (N_187,In_96,In_410);
nor U188 (N_188,In_142,In_208);
nor U189 (N_189,In_364,In_100);
and U190 (N_190,In_259,In_27);
or U191 (N_191,In_445,In_314);
nand U192 (N_192,In_262,In_210);
or U193 (N_193,In_474,In_16);
nor U194 (N_194,In_351,In_70);
and U195 (N_195,In_207,In_468);
nand U196 (N_196,In_318,In_181);
nand U197 (N_197,In_136,In_215);
xnor U198 (N_198,In_230,In_497);
and U199 (N_199,In_311,In_309);
nand U200 (N_200,In_134,In_199);
and U201 (N_201,In_72,In_329);
and U202 (N_202,In_365,In_80);
xnor U203 (N_203,In_439,In_312);
and U204 (N_204,In_172,In_53);
nand U205 (N_205,In_222,In_237);
nand U206 (N_206,In_493,In_344);
xor U207 (N_207,In_217,In_324);
xor U208 (N_208,In_161,In_179);
nor U209 (N_209,In_319,In_88);
and U210 (N_210,In_477,In_185);
or U211 (N_211,In_463,In_341);
nor U212 (N_212,In_413,In_29);
nor U213 (N_213,In_415,In_239);
nand U214 (N_214,In_261,In_52);
and U215 (N_215,In_6,In_211);
and U216 (N_216,In_212,In_406);
or U217 (N_217,In_184,In_14);
and U218 (N_218,In_356,In_405);
xor U219 (N_219,In_35,In_386);
nor U220 (N_220,In_418,In_170);
nand U221 (N_221,In_7,In_180);
xnor U222 (N_222,In_87,In_97);
xnor U223 (N_223,In_11,In_404);
nor U224 (N_224,In_395,In_176);
nor U225 (N_225,In_290,In_108);
nand U226 (N_226,In_498,In_278);
and U227 (N_227,In_412,In_85);
xor U228 (N_228,In_156,In_325);
nor U229 (N_229,In_339,In_61);
xor U230 (N_230,In_480,In_269);
nor U231 (N_231,In_494,In_270);
nand U232 (N_232,In_128,In_55);
or U233 (N_233,In_79,In_251);
or U234 (N_234,In_271,In_203);
nor U235 (N_235,In_48,In_164);
and U236 (N_236,In_265,In_273);
and U237 (N_237,In_91,In_86);
nor U238 (N_238,In_492,In_462);
and U239 (N_239,In_248,In_13);
or U240 (N_240,In_89,In_101);
or U241 (N_241,In_476,In_496);
and U242 (N_242,In_193,In_454);
and U243 (N_243,In_385,In_26);
nor U244 (N_244,In_4,In_337);
and U245 (N_245,In_495,In_374);
and U246 (N_246,In_282,In_448);
nand U247 (N_247,In_145,In_158);
and U248 (N_248,In_308,In_426);
and U249 (N_249,In_400,In_227);
nand U250 (N_250,In_16,In_495);
and U251 (N_251,In_382,In_189);
and U252 (N_252,In_309,In_70);
nand U253 (N_253,In_218,In_333);
nand U254 (N_254,In_345,In_114);
nand U255 (N_255,In_383,In_488);
nor U256 (N_256,In_281,In_284);
and U257 (N_257,In_9,In_31);
nor U258 (N_258,In_432,In_37);
and U259 (N_259,In_116,In_132);
nor U260 (N_260,In_467,In_87);
or U261 (N_261,In_450,In_110);
xor U262 (N_262,In_87,In_151);
nand U263 (N_263,In_344,In_306);
nor U264 (N_264,In_50,In_44);
or U265 (N_265,In_296,In_116);
and U266 (N_266,In_315,In_260);
xnor U267 (N_267,In_271,In_89);
nand U268 (N_268,In_94,In_471);
nand U269 (N_269,In_143,In_434);
and U270 (N_270,In_50,In_86);
nor U271 (N_271,In_90,In_180);
xnor U272 (N_272,In_419,In_302);
nor U273 (N_273,In_380,In_293);
or U274 (N_274,In_188,In_53);
or U275 (N_275,In_337,In_118);
and U276 (N_276,In_4,In_351);
nand U277 (N_277,In_279,In_209);
or U278 (N_278,In_205,In_469);
nor U279 (N_279,In_123,In_332);
or U280 (N_280,In_268,In_184);
and U281 (N_281,In_255,In_347);
and U282 (N_282,In_401,In_404);
nand U283 (N_283,In_97,In_199);
or U284 (N_284,In_291,In_220);
and U285 (N_285,In_33,In_329);
or U286 (N_286,In_144,In_269);
and U287 (N_287,In_337,In_455);
and U288 (N_288,In_113,In_16);
or U289 (N_289,In_45,In_351);
or U290 (N_290,In_310,In_284);
nand U291 (N_291,In_496,In_4);
nand U292 (N_292,In_215,In_8);
and U293 (N_293,In_484,In_323);
xor U294 (N_294,In_68,In_235);
nand U295 (N_295,In_313,In_304);
nand U296 (N_296,In_303,In_175);
nand U297 (N_297,In_208,In_427);
nand U298 (N_298,In_22,In_390);
or U299 (N_299,In_445,In_330);
nor U300 (N_300,In_18,In_341);
or U301 (N_301,In_98,In_151);
nand U302 (N_302,In_18,In_31);
or U303 (N_303,In_131,In_457);
or U304 (N_304,In_361,In_289);
nand U305 (N_305,In_203,In_129);
nor U306 (N_306,In_362,In_50);
and U307 (N_307,In_102,In_44);
xnor U308 (N_308,In_361,In_358);
xnor U309 (N_309,In_164,In_165);
nand U310 (N_310,In_187,In_257);
and U311 (N_311,In_342,In_435);
xnor U312 (N_312,In_446,In_184);
xnor U313 (N_313,In_163,In_476);
and U314 (N_314,In_65,In_343);
or U315 (N_315,In_303,In_202);
nand U316 (N_316,In_488,In_234);
xnor U317 (N_317,In_117,In_372);
or U318 (N_318,In_277,In_471);
nor U319 (N_319,In_120,In_383);
xor U320 (N_320,In_242,In_36);
or U321 (N_321,In_115,In_407);
or U322 (N_322,In_306,In_104);
nand U323 (N_323,In_254,In_39);
nor U324 (N_324,In_410,In_47);
or U325 (N_325,In_242,In_395);
or U326 (N_326,In_411,In_3);
and U327 (N_327,In_49,In_466);
and U328 (N_328,In_256,In_231);
xor U329 (N_329,In_389,In_453);
nor U330 (N_330,In_49,In_358);
xor U331 (N_331,In_236,In_408);
or U332 (N_332,In_107,In_358);
nor U333 (N_333,In_322,In_406);
nor U334 (N_334,In_452,In_150);
or U335 (N_335,In_310,In_464);
xnor U336 (N_336,In_73,In_287);
xor U337 (N_337,In_398,In_322);
or U338 (N_338,In_361,In_321);
nand U339 (N_339,In_182,In_217);
and U340 (N_340,In_15,In_37);
or U341 (N_341,In_225,In_325);
and U342 (N_342,In_270,In_63);
nor U343 (N_343,In_160,In_277);
or U344 (N_344,In_181,In_58);
and U345 (N_345,In_65,In_212);
nor U346 (N_346,In_454,In_418);
or U347 (N_347,In_264,In_99);
xor U348 (N_348,In_72,In_12);
nor U349 (N_349,In_167,In_318);
nand U350 (N_350,In_366,In_145);
or U351 (N_351,In_285,In_393);
nor U352 (N_352,In_152,In_478);
nor U353 (N_353,In_208,In_122);
nor U354 (N_354,In_313,In_291);
and U355 (N_355,In_432,In_160);
nand U356 (N_356,In_378,In_472);
nor U357 (N_357,In_267,In_233);
nand U358 (N_358,In_204,In_418);
or U359 (N_359,In_456,In_132);
and U360 (N_360,In_51,In_409);
xnor U361 (N_361,In_307,In_309);
and U362 (N_362,In_430,In_286);
nand U363 (N_363,In_137,In_385);
nand U364 (N_364,In_453,In_81);
or U365 (N_365,In_83,In_490);
and U366 (N_366,In_342,In_279);
or U367 (N_367,In_493,In_51);
xnor U368 (N_368,In_407,In_390);
nand U369 (N_369,In_159,In_19);
or U370 (N_370,In_467,In_231);
and U371 (N_371,In_133,In_417);
nand U372 (N_372,In_173,In_293);
nor U373 (N_373,In_100,In_39);
nor U374 (N_374,In_306,In_3);
or U375 (N_375,In_165,In_37);
nand U376 (N_376,In_193,In_318);
and U377 (N_377,In_417,In_304);
xor U378 (N_378,In_17,In_279);
and U379 (N_379,In_254,In_81);
or U380 (N_380,In_164,In_394);
and U381 (N_381,In_113,In_292);
xnor U382 (N_382,In_273,In_43);
and U383 (N_383,In_383,In_162);
or U384 (N_384,In_231,In_454);
or U385 (N_385,In_332,In_262);
nor U386 (N_386,In_41,In_144);
xor U387 (N_387,In_351,In_345);
nor U388 (N_388,In_489,In_432);
nor U389 (N_389,In_357,In_270);
or U390 (N_390,In_172,In_68);
or U391 (N_391,In_494,In_160);
or U392 (N_392,In_394,In_124);
nand U393 (N_393,In_484,In_429);
nand U394 (N_394,In_326,In_78);
xnor U395 (N_395,In_365,In_190);
nor U396 (N_396,In_55,In_499);
xnor U397 (N_397,In_175,In_81);
or U398 (N_398,In_86,In_436);
and U399 (N_399,In_477,In_273);
and U400 (N_400,In_37,In_287);
nor U401 (N_401,In_112,In_200);
and U402 (N_402,In_235,In_483);
nor U403 (N_403,In_71,In_421);
xnor U404 (N_404,In_319,In_463);
nand U405 (N_405,In_491,In_297);
nand U406 (N_406,In_34,In_106);
nor U407 (N_407,In_238,In_417);
and U408 (N_408,In_202,In_105);
nand U409 (N_409,In_204,In_102);
nor U410 (N_410,In_140,In_311);
nor U411 (N_411,In_202,In_64);
and U412 (N_412,In_212,In_286);
or U413 (N_413,In_150,In_203);
nor U414 (N_414,In_477,In_365);
xnor U415 (N_415,In_470,In_419);
nand U416 (N_416,In_114,In_344);
or U417 (N_417,In_151,In_188);
and U418 (N_418,In_283,In_281);
xnor U419 (N_419,In_492,In_280);
nand U420 (N_420,In_201,In_141);
and U421 (N_421,In_323,In_425);
nor U422 (N_422,In_342,In_450);
xor U423 (N_423,In_335,In_113);
nor U424 (N_424,In_453,In_291);
nor U425 (N_425,In_318,In_498);
nand U426 (N_426,In_480,In_233);
or U427 (N_427,In_145,In_48);
or U428 (N_428,In_273,In_367);
and U429 (N_429,In_141,In_366);
nand U430 (N_430,In_120,In_214);
and U431 (N_431,In_208,In_340);
nand U432 (N_432,In_142,In_457);
or U433 (N_433,In_231,In_64);
and U434 (N_434,In_425,In_179);
nor U435 (N_435,In_294,In_21);
and U436 (N_436,In_469,In_324);
nor U437 (N_437,In_303,In_438);
and U438 (N_438,In_121,In_235);
nand U439 (N_439,In_421,In_468);
nand U440 (N_440,In_296,In_41);
and U441 (N_441,In_360,In_357);
nand U442 (N_442,In_118,In_236);
or U443 (N_443,In_114,In_133);
nand U444 (N_444,In_120,In_432);
or U445 (N_445,In_98,In_89);
nand U446 (N_446,In_268,In_294);
or U447 (N_447,In_138,In_227);
nand U448 (N_448,In_212,In_146);
nor U449 (N_449,In_0,In_126);
nor U450 (N_450,In_327,In_390);
and U451 (N_451,In_183,In_7);
nand U452 (N_452,In_163,In_171);
and U453 (N_453,In_108,In_314);
and U454 (N_454,In_78,In_100);
nor U455 (N_455,In_196,In_79);
nor U456 (N_456,In_118,In_181);
or U457 (N_457,In_310,In_271);
nand U458 (N_458,In_178,In_493);
and U459 (N_459,In_312,In_329);
nor U460 (N_460,In_283,In_38);
or U461 (N_461,In_331,In_378);
nor U462 (N_462,In_288,In_290);
or U463 (N_463,In_139,In_168);
nor U464 (N_464,In_301,In_0);
nand U465 (N_465,In_279,In_451);
nor U466 (N_466,In_225,In_414);
nand U467 (N_467,In_292,In_359);
nor U468 (N_468,In_70,In_416);
nor U469 (N_469,In_400,In_150);
and U470 (N_470,In_261,In_172);
and U471 (N_471,In_177,In_472);
nand U472 (N_472,In_37,In_304);
nand U473 (N_473,In_24,In_147);
nor U474 (N_474,In_286,In_491);
nand U475 (N_475,In_398,In_210);
and U476 (N_476,In_245,In_371);
nor U477 (N_477,In_478,In_295);
nand U478 (N_478,In_493,In_149);
nand U479 (N_479,In_57,In_260);
and U480 (N_480,In_334,In_386);
xnor U481 (N_481,In_163,In_147);
or U482 (N_482,In_189,In_240);
or U483 (N_483,In_52,In_36);
and U484 (N_484,In_78,In_204);
and U485 (N_485,In_385,In_419);
and U486 (N_486,In_94,In_114);
or U487 (N_487,In_182,In_224);
nand U488 (N_488,In_32,In_55);
or U489 (N_489,In_96,In_121);
nor U490 (N_490,In_492,In_68);
nor U491 (N_491,In_214,In_167);
nor U492 (N_492,In_68,In_470);
xor U493 (N_493,In_70,In_80);
or U494 (N_494,In_85,In_75);
nand U495 (N_495,In_11,In_227);
nand U496 (N_496,In_85,In_252);
and U497 (N_497,In_387,In_160);
or U498 (N_498,In_69,In_296);
nand U499 (N_499,In_256,In_470);
or U500 (N_500,In_334,In_210);
or U501 (N_501,In_44,In_478);
and U502 (N_502,In_105,In_219);
and U503 (N_503,In_483,In_439);
nor U504 (N_504,In_284,In_2);
nor U505 (N_505,In_400,In_14);
xnor U506 (N_506,In_297,In_145);
or U507 (N_507,In_431,In_492);
or U508 (N_508,In_377,In_452);
nor U509 (N_509,In_92,In_497);
or U510 (N_510,In_311,In_446);
nand U511 (N_511,In_405,In_480);
nor U512 (N_512,In_490,In_247);
or U513 (N_513,In_316,In_380);
nor U514 (N_514,In_30,In_45);
xor U515 (N_515,In_205,In_0);
nor U516 (N_516,In_300,In_94);
or U517 (N_517,In_371,In_490);
nor U518 (N_518,In_499,In_205);
and U519 (N_519,In_6,In_97);
and U520 (N_520,In_467,In_345);
nand U521 (N_521,In_168,In_233);
nor U522 (N_522,In_332,In_290);
and U523 (N_523,In_472,In_225);
or U524 (N_524,In_84,In_391);
and U525 (N_525,In_195,In_90);
nand U526 (N_526,In_175,In_179);
xor U527 (N_527,In_269,In_466);
nor U528 (N_528,In_398,In_2);
nor U529 (N_529,In_242,In_497);
xnor U530 (N_530,In_378,In_101);
or U531 (N_531,In_242,In_398);
and U532 (N_532,In_42,In_450);
or U533 (N_533,In_166,In_109);
nor U534 (N_534,In_178,In_372);
nor U535 (N_535,In_373,In_221);
nor U536 (N_536,In_276,In_231);
and U537 (N_537,In_421,In_442);
and U538 (N_538,In_165,In_317);
or U539 (N_539,In_333,In_381);
xnor U540 (N_540,In_27,In_289);
xor U541 (N_541,In_62,In_343);
nand U542 (N_542,In_323,In_344);
or U543 (N_543,In_254,In_79);
nor U544 (N_544,In_19,In_279);
and U545 (N_545,In_240,In_439);
nor U546 (N_546,In_110,In_104);
and U547 (N_547,In_441,In_94);
and U548 (N_548,In_108,In_367);
or U549 (N_549,In_119,In_219);
nand U550 (N_550,In_47,In_388);
and U551 (N_551,In_474,In_453);
xnor U552 (N_552,In_67,In_339);
and U553 (N_553,In_316,In_281);
and U554 (N_554,In_479,In_204);
nand U555 (N_555,In_40,In_370);
nand U556 (N_556,In_49,In_279);
and U557 (N_557,In_456,In_420);
nand U558 (N_558,In_399,In_316);
nor U559 (N_559,In_60,In_27);
nand U560 (N_560,In_165,In_324);
and U561 (N_561,In_410,In_465);
and U562 (N_562,In_283,In_204);
xnor U563 (N_563,In_313,In_351);
nor U564 (N_564,In_53,In_496);
and U565 (N_565,In_86,In_430);
xor U566 (N_566,In_243,In_104);
and U567 (N_567,In_384,In_269);
nand U568 (N_568,In_100,In_95);
nor U569 (N_569,In_158,In_37);
nor U570 (N_570,In_402,In_491);
nand U571 (N_571,In_267,In_445);
and U572 (N_572,In_394,In_184);
nor U573 (N_573,In_435,In_90);
or U574 (N_574,In_57,In_285);
and U575 (N_575,In_343,In_49);
and U576 (N_576,In_38,In_82);
nand U577 (N_577,In_282,In_237);
or U578 (N_578,In_383,In_272);
nand U579 (N_579,In_319,In_458);
xnor U580 (N_580,In_361,In_466);
xnor U581 (N_581,In_168,In_108);
or U582 (N_582,In_28,In_30);
nand U583 (N_583,In_243,In_444);
xnor U584 (N_584,In_470,In_393);
and U585 (N_585,In_377,In_308);
nand U586 (N_586,In_338,In_114);
nor U587 (N_587,In_261,In_107);
and U588 (N_588,In_332,In_35);
nand U589 (N_589,In_368,In_455);
and U590 (N_590,In_244,In_305);
or U591 (N_591,In_63,In_21);
nor U592 (N_592,In_141,In_185);
nand U593 (N_593,In_460,In_20);
nand U594 (N_594,In_360,In_372);
or U595 (N_595,In_301,In_377);
nand U596 (N_596,In_42,In_31);
nor U597 (N_597,In_377,In_120);
nor U598 (N_598,In_381,In_78);
xor U599 (N_599,In_453,In_375);
or U600 (N_600,In_447,In_44);
xor U601 (N_601,In_352,In_227);
or U602 (N_602,In_139,In_113);
nor U603 (N_603,In_461,In_418);
and U604 (N_604,In_68,In_337);
nor U605 (N_605,In_441,In_447);
or U606 (N_606,In_388,In_476);
nor U607 (N_607,In_323,In_469);
xnor U608 (N_608,In_488,In_204);
or U609 (N_609,In_10,In_482);
nor U610 (N_610,In_367,In_363);
nor U611 (N_611,In_102,In_256);
nor U612 (N_612,In_142,In_23);
and U613 (N_613,In_20,In_13);
nor U614 (N_614,In_460,In_405);
nor U615 (N_615,In_137,In_158);
xnor U616 (N_616,In_352,In_410);
or U617 (N_617,In_19,In_109);
nor U618 (N_618,In_133,In_262);
or U619 (N_619,In_397,In_24);
nand U620 (N_620,In_65,In_184);
nor U621 (N_621,In_447,In_238);
nor U622 (N_622,In_234,In_79);
nand U623 (N_623,In_173,In_140);
or U624 (N_624,In_283,In_80);
xor U625 (N_625,In_306,In_453);
xor U626 (N_626,In_55,In_87);
nand U627 (N_627,In_454,In_412);
and U628 (N_628,In_320,In_85);
nor U629 (N_629,In_5,In_313);
nand U630 (N_630,In_74,In_57);
xor U631 (N_631,In_11,In_419);
nor U632 (N_632,In_462,In_330);
or U633 (N_633,In_296,In_231);
nor U634 (N_634,In_29,In_282);
nor U635 (N_635,In_191,In_302);
nor U636 (N_636,In_372,In_138);
nand U637 (N_637,In_146,In_235);
xnor U638 (N_638,In_299,In_480);
and U639 (N_639,In_2,In_50);
nand U640 (N_640,In_242,In_177);
xor U641 (N_641,In_396,In_33);
xnor U642 (N_642,In_465,In_104);
nor U643 (N_643,In_190,In_449);
nand U644 (N_644,In_280,In_347);
nor U645 (N_645,In_482,In_305);
nor U646 (N_646,In_91,In_4);
and U647 (N_647,In_388,In_292);
and U648 (N_648,In_225,In_253);
nand U649 (N_649,In_363,In_78);
nand U650 (N_650,In_93,In_243);
and U651 (N_651,In_275,In_164);
or U652 (N_652,In_282,In_440);
nand U653 (N_653,In_133,In_190);
and U654 (N_654,In_149,In_187);
nand U655 (N_655,In_175,In_428);
and U656 (N_656,In_456,In_394);
nor U657 (N_657,In_385,In_470);
nor U658 (N_658,In_452,In_111);
and U659 (N_659,In_406,In_251);
nor U660 (N_660,In_184,In_88);
and U661 (N_661,In_357,In_207);
nor U662 (N_662,In_338,In_299);
xor U663 (N_663,In_363,In_324);
xnor U664 (N_664,In_312,In_158);
nor U665 (N_665,In_180,In_312);
nand U666 (N_666,In_301,In_68);
and U667 (N_667,In_322,In_243);
nand U668 (N_668,In_438,In_207);
or U669 (N_669,In_438,In_362);
nor U670 (N_670,In_260,In_322);
nand U671 (N_671,In_299,In_195);
or U672 (N_672,In_167,In_32);
xor U673 (N_673,In_491,In_248);
nand U674 (N_674,In_377,In_274);
and U675 (N_675,In_440,In_273);
or U676 (N_676,In_478,In_249);
nand U677 (N_677,In_134,In_224);
and U678 (N_678,In_450,In_418);
nand U679 (N_679,In_101,In_299);
nand U680 (N_680,In_283,In_222);
nand U681 (N_681,In_423,In_237);
and U682 (N_682,In_38,In_209);
or U683 (N_683,In_9,In_72);
and U684 (N_684,In_138,In_344);
or U685 (N_685,In_28,In_100);
nor U686 (N_686,In_234,In_30);
or U687 (N_687,In_12,In_131);
and U688 (N_688,In_114,In_355);
nor U689 (N_689,In_103,In_187);
and U690 (N_690,In_314,In_415);
or U691 (N_691,In_277,In_6);
and U692 (N_692,In_153,In_163);
and U693 (N_693,In_436,In_68);
and U694 (N_694,In_55,In_262);
nand U695 (N_695,In_177,In_406);
or U696 (N_696,In_405,In_424);
xor U697 (N_697,In_158,In_444);
and U698 (N_698,In_55,In_470);
or U699 (N_699,In_385,In_490);
xnor U700 (N_700,In_103,In_127);
and U701 (N_701,In_196,In_294);
and U702 (N_702,In_415,In_448);
nor U703 (N_703,In_489,In_423);
and U704 (N_704,In_37,In_212);
nor U705 (N_705,In_466,In_206);
xnor U706 (N_706,In_298,In_89);
or U707 (N_707,In_189,In_207);
nor U708 (N_708,In_263,In_45);
and U709 (N_709,In_127,In_146);
and U710 (N_710,In_401,In_83);
nand U711 (N_711,In_13,In_138);
and U712 (N_712,In_201,In_65);
nand U713 (N_713,In_15,In_320);
or U714 (N_714,In_490,In_176);
and U715 (N_715,In_215,In_372);
nand U716 (N_716,In_208,In_296);
and U717 (N_717,In_95,In_119);
nor U718 (N_718,In_412,In_376);
or U719 (N_719,In_388,In_194);
nand U720 (N_720,In_401,In_373);
and U721 (N_721,In_89,In_190);
and U722 (N_722,In_311,In_494);
nand U723 (N_723,In_221,In_200);
nand U724 (N_724,In_342,In_321);
nand U725 (N_725,In_288,In_446);
and U726 (N_726,In_490,In_126);
and U727 (N_727,In_257,In_125);
and U728 (N_728,In_327,In_267);
nor U729 (N_729,In_35,In_149);
and U730 (N_730,In_121,In_183);
and U731 (N_731,In_160,In_487);
nand U732 (N_732,In_31,In_347);
nand U733 (N_733,In_439,In_239);
or U734 (N_734,In_275,In_350);
nor U735 (N_735,In_247,In_77);
xnor U736 (N_736,In_465,In_274);
or U737 (N_737,In_434,In_185);
or U738 (N_738,In_29,In_27);
and U739 (N_739,In_190,In_81);
nand U740 (N_740,In_269,In_351);
nor U741 (N_741,In_379,In_47);
or U742 (N_742,In_178,In_385);
nor U743 (N_743,In_424,In_430);
xor U744 (N_744,In_134,In_298);
nand U745 (N_745,In_168,In_478);
nand U746 (N_746,In_82,In_311);
nand U747 (N_747,In_102,In_115);
xor U748 (N_748,In_50,In_358);
and U749 (N_749,In_361,In_417);
nand U750 (N_750,N_552,N_77);
nand U751 (N_751,N_386,N_633);
nor U752 (N_752,N_278,N_609);
or U753 (N_753,N_1,N_102);
xnor U754 (N_754,N_90,N_607);
nand U755 (N_755,N_747,N_524);
and U756 (N_756,N_119,N_113);
nor U757 (N_757,N_564,N_49);
and U758 (N_758,N_9,N_337);
nor U759 (N_759,N_247,N_594);
nand U760 (N_760,N_612,N_478);
or U761 (N_761,N_448,N_323);
and U762 (N_762,N_616,N_710);
or U763 (N_763,N_503,N_551);
nand U764 (N_764,N_212,N_365);
or U765 (N_765,N_249,N_675);
nand U766 (N_766,N_228,N_590);
or U767 (N_767,N_694,N_682);
nor U768 (N_768,N_719,N_38);
or U769 (N_769,N_68,N_192);
nand U770 (N_770,N_405,N_541);
xor U771 (N_771,N_341,N_651);
nor U772 (N_772,N_592,N_536);
nor U773 (N_773,N_573,N_387);
nor U774 (N_774,N_122,N_267);
or U775 (N_775,N_589,N_553);
nor U776 (N_776,N_545,N_596);
or U777 (N_777,N_304,N_356);
nand U778 (N_778,N_454,N_44);
nand U779 (N_779,N_438,N_168);
or U780 (N_780,N_29,N_588);
xor U781 (N_781,N_453,N_737);
and U782 (N_782,N_225,N_24);
nor U783 (N_783,N_209,N_123);
nand U784 (N_784,N_426,N_504);
or U785 (N_785,N_474,N_67);
or U786 (N_786,N_402,N_429);
xor U787 (N_787,N_557,N_692);
or U788 (N_788,N_208,N_650);
nand U789 (N_789,N_582,N_408);
nand U790 (N_790,N_574,N_189);
nor U791 (N_791,N_727,N_458);
nand U792 (N_792,N_668,N_734);
nor U793 (N_793,N_57,N_124);
and U794 (N_794,N_60,N_490);
and U795 (N_795,N_593,N_40);
nand U796 (N_796,N_657,N_342);
and U797 (N_797,N_731,N_262);
nor U798 (N_798,N_510,N_652);
nor U799 (N_799,N_647,N_41);
or U800 (N_800,N_374,N_463);
or U801 (N_801,N_540,N_667);
and U802 (N_802,N_255,N_94);
or U803 (N_803,N_706,N_39);
and U804 (N_804,N_360,N_210);
nand U805 (N_805,N_580,N_466);
and U806 (N_806,N_270,N_70);
nor U807 (N_807,N_696,N_404);
nand U808 (N_808,N_437,N_591);
xor U809 (N_809,N_598,N_717);
nand U810 (N_810,N_281,N_103);
and U811 (N_811,N_640,N_608);
nor U812 (N_812,N_492,N_266);
or U813 (N_813,N_641,N_296);
nand U814 (N_814,N_152,N_555);
nor U815 (N_815,N_235,N_544);
nor U816 (N_816,N_450,N_644);
nor U817 (N_817,N_321,N_72);
nor U818 (N_818,N_479,N_625);
nand U819 (N_819,N_193,N_283);
or U820 (N_820,N_234,N_314);
nand U821 (N_821,N_377,N_223);
and U822 (N_822,N_610,N_111);
or U823 (N_823,N_600,N_128);
nor U824 (N_824,N_711,N_568);
or U825 (N_825,N_280,N_579);
and U826 (N_826,N_654,N_338);
and U827 (N_827,N_166,N_664);
and U828 (N_828,N_489,N_459);
nand U829 (N_829,N_260,N_475);
nor U830 (N_830,N_271,N_491);
nand U831 (N_831,N_78,N_261);
nor U832 (N_832,N_132,N_96);
and U833 (N_833,N_53,N_221);
or U834 (N_834,N_398,N_37);
xor U835 (N_835,N_167,N_393);
or U836 (N_836,N_748,N_363);
nor U837 (N_837,N_332,N_316);
nor U838 (N_838,N_302,N_186);
nand U839 (N_839,N_101,N_483);
xnor U840 (N_840,N_54,N_645);
or U841 (N_841,N_198,N_13);
nand U842 (N_842,N_721,N_163);
nor U843 (N_843,N_643,N_361);
xor U844 (N_844,N_626,N_171);
nand U845 (N_845,N_403,N_36);
and U846 (N_846,N_354,N_521);
and U847 (N_847,N_415,N_118);
nor U848 (N_848,N_334,N_485);
and U849 (N_849,N_330,N_367);
nor U850 (N_850,N_732,N_71);
and U851 (N_851,N_100,N_563);
nor U852 (N_852,N_133,N_333);
nor U853 (N_853,N_22,N_435);
nand U854 (N_854,N_250,N_97);
nor U855 (N_855,N_130,N_134);
and U856 (N_856,N_389,N_507);
nand U857 (N_857,N_66,N_177);
xor U858 (N_858,N_81,N_172);
and U859 (N_859,N_31,N_497);
nand U860 (N_860,N_656,N_595);
nand U861 (N_861,N_233,N_547);
or U862 (N_862,N_526,N_529);
nor U863 (N_863,N_83,N_179);
nor U864 (N_864,N_371,N_197);
and U865 (N_865,N_251,N_274);
nand U866 (N_866,N_410,N_394);
or U867 (N_867,N_318,N_533);
xnor U868 (N_868,N_462,N_30);
or U869 (N_869,N_702,N_336);
nor U870 (N_870,N_701,N_421);
or U871 (N_871,N_704,N_350);
or U872 (N_872,N_95,N_542);
or U873 (N_873,N_181,N_185);
and U874 (N_874,N_213,N_423);
nand U875 (N_875,N_465,N_217);
and U876 (N_876,N_639,N_259);
nand U877 (N_877,N_246,N_433);
and U878 (N_878,N_382,N_617);
or U879 (N_879,N_455,N_680);
nand U880 (N_880,N_43,N_349);
xor U881 (N_881,N_401,N_476);
and U882 (N_882,N_722,N_297);
nor U883 (N_883,N_575,N_705);
or U884 (N_884,N_91,N_661);
nor U885 (N_885,N_419,N_290);
and U886 (N_886,N_88,N_12);
nor U887 (N_887,N_520,N_169);
or U888 (N_888,N_666,N_630);
nand U889 (N_889,N_581,N_413);
or U890 (N_890,N_121,N_556);
or U891 (N_891,N_58,N_190);
or U892 (N_892,N_665,N_681);
nand U893 (N_893,N_561,N_180);
nand U894 (N_894,N_275,N_187);
xor U895 (N_895,N_295,N_222);
nor U896 (N_896,N_471,N_372);
or U897 (N_897,N_139,N_370);
and U898 (N_898,N_601,N_576);
nor U899 (N_899,N_659,N_3);
nand U900 (N_900,N_170,N_147);
and U901 (N_901,N_265,N_5);
or U902 (N_902,N_514,N_369);
xor U903 (N_903,N_472,N_736);
xor U904 (N_904,N_344,N_375);
or U905 (N_905,N_570,N_106);
and U906 (N_906,N_324,N_182);
nor U907 (N_907,N_632,N_512);
nor U908 (N_908,N_707,N_390);
and U909 (N_909,N_137,N_519);
or U910 (N_910,N_715,N_740);
xnor U911 (N_911,N_117,N_535);
or U912 (N_912,N_373,N_328);
and U913 (N_913,N_467,N_456);
and U914 (N_914,N_460,N_143);
or U915 (N_915,N_619,N_352);
or U916 (N_916,N_257,N_464);
or U917 (N_917,N_534,N_219);
xor U918 (N_918,N_412,N_618);
or U919 (N_919,N_378,N_220);
xnor U920 (N_920,N_531,N_241);
or U921 (N_921,N_417,N_0);
xor U922 (N_922,N_599,N_291);
nand U923 (N_923,N_461,N_47);
and U924 (N_924,N_391,N_506);
xor U925 (N_925,N_688,N_516);
or U926 (N_926,N_145,N_549);
and U927 (N_927,N_495,N_194);
or U928 (N_928,N_428,N_331);
xor U929 (N_929,N_546,N_311);
nor U930 (N_930,N_470,N_380);
nor U931 (N_931,N_603,N_6);
nand U932 (N_932,N_305,N_624);
nand U933 (N_933,N_399,N_559);
nor U934 (N_934,N_62,N_200);
or U935 (N_935,N_204,N_345);
or U936 (N_936,N_439,N_244);
and U937 (N_937,N_277,N_87);
xnor U938 (N_938,N_42,N_744);
nand U939 (N_939,N_567,N_745);
nor U940 (N_940,N_499,N_55);
and U941 (N_941,N_469,N_376);
or U942 (N_942,N_714,N_724);
and U943 (N_943,N_184,N_712);
nor U944 (N_944,N_728,N_8);
nand U945 (N_945,N_154,N_725);
and U946 (N_946,N_35,N_310);
nand U947 (N_947,N_445,N_59);
and U948 (N_948,N_226,N_698);
and U949 (N_949,N_206,N_86);
nand U950 (N_950,N_205,N_15);
nor U951 (N_951,N_135,N_45);
and U952 (N_952,N_395,N_739);
xor U953 (N_953,N_585,N_730);
or U954 (N_954,N_115,N_73);
nor U955 (N_955,N_703,N_487);
nor U956 (N_956,N_396,N_420);
nor U957 (N_957,N_34,N_287);
and U958 (N_958,N_508,N_174);
nor U959 (N_959,N_319,N_343);
and U960 (N_960,N_597,N_92);
and U961 (N_961,N_443,N_315);
nand U962 (N_962,N_366,N_741);
or U963 (N_963,N_158,N_362);
nor U964 (N_964,N_566,N_713);
or U965 (N_965,N_648,N_543);
nand U966 (N_966,N_153,N_407);
or U967 (N_967,N_441,N_127);
or U968 (N_968,N_572,N_294);
or U969 (N_969,N_658,N_108);
and U970 (N_970,N_447,N_473);
or U971 (N_971,N_708,N_16);
and U972 (N_972,N_468,N_735);
or U973 (N_973,N_4,N_742);
nor U974 (N_974,N_2,N_511);
nor U975 (N_975,N_239,N_230);
and U976 (N_976,N_528,N_19);
or U977 (N_977,N_199,N_718);
nor U978 (N_978,N_571,N_638);
and U979 (N_979,N_669,N_379);
and U980 (N_980,N_339,N_700);
xnor U981 (N_981,N_52,N_74);
nor U982 (N_982,N_381,N_484);
and U983 (N_983,N_684,N_517);
and U984 (N_984,N_162,N_690);
and U985 (N_985,N_709,N_201);
xor U986 (N_986,N_203,N_82);
or U987 (N_987,N_355,N_409);
nor U988 (N_988,N_273,N_749);
or U989 (N_989,N_173,N_602);
nor U990 (N_990,N_240,N_28);
or U991 (N_991,N_149,N_326);
nor U992 (N_992,N_320,N_418);
nand U993 (N_993,N_146,N_129);
nor U994 (N_994,N_627,N_160);
nor U995 (N_995,N_288,N_27);
or U996 (N_996,N_631,N_32);
or U997 (N_997,N_486,N_422);
nor U998 (N_998,N_655,N_434);
nand U999 (N_999,N_364,N_79);
or U1000 (N_1000,N_673,N_232);
nand U1001 (N_1001,N_218,N_577);
nor U1002 (N_1002,N_432,N_646);
and U1003 (N_1003,N_23,N_628);
nor U1004 (N_1004,N_89,N_357);
or U1005 (N_1005,N_500,N_416);
and U1006 (N_1006,N_17,N_560);
or U1007 (N_1007,N_697,N_532);
or U1008 (N_1008,N_562,N_424);
nand U1009 (N_1009,N_522,N_629);
xor U1010 (N_1010,N_313,N_178);
nor U1011 (N_1011,N_527,N_346);
or U1012 (N_1012,N_126,N_442);
nand U1013 (N_1013,N_446,N_300);
or U1014 (N_1014,N_358,N_674);
nor U1015 (N_1015,N_317,N_347);
nor U1016 (N_1016,N_444,N_183);
xor U1017 (N_1017,N_502,N_105);
or U1018 (N_1018,N_440,N_340);
and U1019 (N_1019,N_537,N_642);
nor U1020 (N_1020,N_243,N_548);
and U1021 (N_1021,N_104,N_660);
nand U1022 (N_1022,N_269,N_530);
nor U1023 (N_1023,N_653,N_276);
nand U1024 (N_1024,N_348,N_85);
nand U1025 (N_1025,N_175,N_202);
or U1026 (N_1026,N_481,N_286);
or U1027 (N_1027,N_161,N_687);
nor U1028 (N_1028,N_256,N_33);
nand U1029 (N_1029,N_227,N_676);
xnor U1030 (N_1030,N_248,N_11);
xor U1031 (N_1031,N_729,N_65);
nor U1032 (N_1032,N_569,N_691);
nor U1033 (N_1033,N_292,N_615);
nand U1034 (N_1034,N_236,N_351);
nor U1035 (N_1035,N_207,N_148);
nor U1036 (N_1036,N_188,N_238);
nor U1037 (N_1037,N_623,N_98);
nor U1038 (N_1038,N_430,N_604);
or U1039 (N_1039,N_622,N_678);
nand U1040 (N_1040,N_621,N_141);
xnor U1041 (N_1041,N_289,N_488);
nor U1042 (N_1042,N_672,N_746);
and U1043 (N_1043,N_231,N_306);
or U1044 (N_1044,N_634,N_144);
or U1045 (N_1045,N_695,N_677);
nand U1046 (N_1046,N_663,N_620);
nand U1047 (N_1047,N_254,N_75);
or U1048 (N_1048,N_411,N_114);
or U1049 (N_1049,N_685,N_494);
nor U1050 (N_1050,N_264,N_699);
nand U1051 (N_1051,N_584,N_48);
nand U1052 (N_1052,N_263,N_406);
and U1053 (N_1053,N_109,N_303);
nand U1054 (N_1054,N_253,N_258);
or U1055 (N_1055,N_196,N_637);
nor U1056 (N_1056,N_307,N_157);
or U1057 (N_1057,N_578,N_299);
or U1058 (N_1058,N_480,N_51);
nor U1059 (N_1059,N_452,N_21);
or U1060 (N_1060,N_150,N_195);
or U1061 (N_1061,N_493,N_538);
or U1062 (N_1062,N_252,N_693);
nand U1063 (N_1063,N_689,N_312);
and U1064 (N_1064,N_550,N_301);
nand U1065 (N_1065,N_477,N_140);
or U1066 (N_1066,N_325,N_93);
xor U1067 (N_1067,N_322,N_383);
and U1068 (N_1068,N_309,N_397);
nor U1069 (N_1069,N_436,N_587);
nor U1070 (N_1070,N_99,N_61);
or U1071 (N_1071,N_686,N_558);
xor U1072 (N_1072,N_245,N_723);
xnor U1073 (N_1073,N_279,N_670);
and U1074 (N_1074,N_385,N_523);
and U1075 (N_1075,N_50,N_211);
xor U1076 (N_1076,N_414,N_46);
nor U1077 (N_1077,N_635,N_14);
xor U1078 (N_1078,N_214,N_125);
nand U1079 (N_1079,N_191,N_155);
nor U1080 (N_1080,N_63,N_498);
nor U1081 (N_1081,N_427,N_285);
nor U1082 (N_1082,N_720,N_679);
nand U1083 (N_1083,N_662,N_56);
xnor U1084 (N_1084,N_131,N_216);
or U1085 (N_1085,N_176,N_76);
nor U1086 (N_1086,N_7,N_112);
nor U1087 (N_1087,N_138,N_457);
nor U1088 (N_1088,N_451,N_505);
xor U1089 (N_1089,N_136,N_606);
nand U1090 (N_1090,N_242,N_359);
nor U1091 (N_1091,N_384,N_293);
or U1092 (N_1092,N_613,N_308);
xnor U1093 (N_1093,N_449,N_110);
nand U1094 (N_1094,N_26,N_284);
nand U1095 (N_1095,N_501,N_518);
or U1096 (N_1096,N_636,N_392);
nor U1097 (N_1097,N_215,N_400);
xnor U1098 (N_1098,N_10,N_18);
and U1099 (N_1099,N_116,N_649);
nand U1100 (N_1100,N_84,N_69);
nand U1101 (N_1101,N_431,N_329);
nor U1102 (N_1102,N_496,N_513);
or U1103 (N_1103,N_142,N_156);
nand U1104 (N_1104,N_509,N_743);
and U1105 (N_1105,N_482,N_237);
xor U1106 (N_1106,N_164,N_25);
nor U1107 (N_1107,N_107,N_353);
nand U1108 (N_1108,N_586,N_716);
xnor U1109 (N_1109,N_159,N_268);
nor U1110 (N_1110,N_20,N_229);
nand U1111 (N_1111,N_165,N_80);
nor U1112 (N_1112,N_525,N_335);
nand U1113 (N_1113,N_583,N_282);
and U1114 (N_1114,N_554,N_726);
nor U1115 (N_1115,N_539,N_64);
nand U1116 (N_1116,N_272,N_565);
nor U1117 (N_1117,N_120,N_738);
and U1118 (N_1118,N_151,N_611);
or U1119 (N_1119,N_671,N_515);
or U1120 (N_1120,N_733,N_605);
nor U1121 (N_1121,N_327,N_298);
and U1122 (N_1122,N_614,N_368);
xor U1123 (N_1123,N_388,N_224);
nand U1124 (N_1124,N_683,N_425);
nor U1125 (N_1125,N_628,N_468);
or U1126 (N_1126,N_582,N_12);
nand U1127 (N_1127,N_573,N_51);
and U1128 (N_1128,N_395,N_296);
or U1129 (N_1129,N_355,N_721);
nand U1130 (N_1130,N_53,N_14);
or U1131 (N_1131,N_94,N_378);
nor U1132 (N_1132,N_193,N_664);
and U1133 (N_1133,N_435,N_137);
or U1134 (N_1134,N_544,N_371);
nand U1135 (N_1135,N_417,N_369);
or U1136 (N_1136,N_99,N_103);
nor U1137 (N_1137,N_366,N_119);
or U1138 (N_1138,N_601,N_643);
nand U1139 (N_1139,N_287,N_578);
or U1140 (N_1140,N_686,N_80);
nand U1141 (N_1141,N_535,N_143);
nand U1142 (N_1142,N_716,N_481);
and U1143 (N_1143,N_471,N_192);
and U1144 (N_1144,N_658,N_310);
and U1145 (N_1145,N_729,N_612);
nor U1146 (N_1146,N_435,N_224);
xnor U1147 (N_1147,N_676,N_107);
xor U1148 (N_1148,N_479,N_185);
or U1149 (N_1149,N_547,N_165);
nand U1150 (N_1150,N_624,N_124);
nand U1151 (N_1151,N_302,N_719);
or U1152 (N_1152,N_738,N_200);
nor U1153 (N_1153,N_623,N_493);
nand U1154 (N_1154,N_574,N_428);
and U1155 (N_1155,N_457,N_643);
and U1156 (N_1156,N_116,N_722);
xor U1157 (N_1157,N_461,N_199);
or U1158 (N_1158,N_333,N_595);
and U1159 (N_1159,N_638,N_143);
and U1160 (N_1160,N_407,N_3);
nand U1161 (N_1161,N_689,N_269);
or U1162 (N_1162,N_354,N_690);
xor U1163 (N_1163,N_335,N_380);
and U1164 (N_1164,N_635,N_344);
and U1165 (N_1165,N_226,N_123);
xnor U1166 (N_1166,N_740,N_38);
xnor U1167 (N_1167,N_256,N_271);
nand U1168 (N_1168,N_649,N_317);
nand U1169 (N_1169,N_598,N_477);
nor U1170 (N_1170,N_365,N_516);
and U1171 (N_1171,N_296,N_672);
nor U1172 (N_1172,N_618,N_217);
or U1173 (N_1173,N_378,N_749);
nand U1174 (N_1174,N_151,N_138);
and U1175 (N_1175,N_73,N_631);
xor U1176 (N_1176,N_686,N_20);
xnor U1177 (N_1177,N_356,N_536);
xnor U1178 (N_1178,N_507,N_298);
nand U1179 (N_1179,N_382,N_502);
nand U1180 (N_1180,N_147,N_167);
nor U1181 (N_1181,N_287,N_569);
nor U1182 (N_1182,N_378,N_4);
xor U1183 (N_1183,N_420,N_205);
and U1184 (N_1184,N_605,N_250);
or U1185 (N_1185,N_209,N_155);
nand U1186 (N_1186,N_178,N_6);
nor U1187 (N_1187,N_468,N_119);
and U1188 (N_1188,N_321,N_366);
nor U1189 (N_1189,N_412,N_208);
nor U1190 (N_1190,N_37,N_672);
or U1191 (N_1191,N_82,N_414);
and U1192 (N_1192,N_414,N_502);
nand U1193 (N_1193,N_28,N_164);
and U1194 (N_1194,N_717,N_101);
nand U1195 (N_1195,N_655,N_67);
and U1196 (N_1196,N_206,N_194);
nor U1197 (N_1197,N_19,N_325);
and U1198 (N_1198,N_620,N_188);
nor U1199 (N_1199,N_113,N_288);
nand U1200 (N_1200,N_72,N_62);
nor U1201 (N_1201,N_257,N_101);
nand U1202 (N_1202,N_630,N_667);
and U1203 (N_1203,N_560,N_485);
nand U1204 (N_1204,N_660,N_311);
and U1205 (N_1205,N_128,N_599);
or U1206 (N_1206,N_427,N_548);
and U1207 (N_1207,N_556,N_198);
and U1208 (N_1208,N_460,N_78);
and U1209 (N_1209,N_245,N_286);
nand U1210 (N_1210,N_390,N_718);
and U1211 (N_1211,N_165,N_634);
xor U1212 (N_1212,N_227,N_125);
or U1213 (N_1213,N_296,N_398);
nand U1214 (N_1214,N_52,N_543);
or U1215 (N_1215,N_716,N_670);
or U1216 (N_1216,N_167,N_22);
nor U1217 (N_1217,N_662,N_493);
nor U1218 (N_1218,N_418,N_564);
nand U1219 (N_1219,N_543,N_595);
nor U1220 (N_1220,N_201,N_386);
nor U1221 (N_1221,N_319,N_210);
xnor U1222 (N_1222,N_184,N_129);
nand U1223 (N_1223,N_241,N_670);
nor U1224 (N_1224,N_369,N_505);
or U1225 (N_1225,N_620,N_512);
xor U1226 (N_1226,N_747,N_541);
nor U1227 (N_1227,N_465,N_632);
and U1228 (N_1228,N_393,N_375);
or U1229 (N_1229,N_282,N_272);
or U1230 (N_1230,N_735,N_296);
and U1231 (N_1231,N_434,N_508);
or U1232 (N_1232,N_107,N_102);
nand U1233 (N_1233,N_130,N_186);
nand U1234 (N_1234,N_165,N_11);
or U1235 (N_1235,N_512,N_672);
or U1236 (N_1236,N_693,N_450);
nor U1237 (N_1237,N_595,N_606);
nor U1238 (N_1238,N_268,N_622);
nand U1239 (N_1239,N_2,N_667);
nand U1240 (N_1240,N_108,N_89);
or U1241 (N_1241,N_692,N_192);
or U1242 (N_1242,N_118,N_425);
nor U1243 (N_1243,N_447,N_211);
nor U1244 (N_1244,N_595,N_226);
or U1245 (N_1245,N_219,N_135);
or U1246 (N_1246,N_705,N_441);
nand U1247 (N_1247,N_138,N_687);
nor U1248 (N_1248,N_659,N_89);
or U1249 (N_1249,N_169,N_652);
xor U1250 (N_1250,N_700,N_302);
or U1251 (N_1251,N_384,N_37);
and U1252 (N_1252,N_334,N_108);
nand U1253 (N_1253,N_370,N_539);
nand U1254 (N_1254,N_525,N_428);
nand U1255 (N_1255,N_114,N_550);
nor U1256 (N_1256,N_269,N_587);
xor U1257 (N_1257,N_294,N_436);
and U1258 (N_1258,N_6,N_220);
nor U1259 (N_1259,N_528,N_451);
nand U1260 (N_1260,N_415,N_337);
nor U1261 (N_1261,N_690,N_508);
or U1262 (N_1262,N_721,N_131);
nor U1263 (N_1263,N_287,N_418);
and U1264 (N_1264,N_574,N_656);
nand U1265 (N_1265,N_289,N_471);
or U1266 (N_1266,N_446,N_604);
and U1267 (N_1267,N_347,N_588);
and U1268 (N_1268,N_540,N_510);
and U1269 (N_1269,N_272,N_410);
nor U1270 (N_1270,N_620,N_553);
nor U1271 (N_1271,N_681,N_259);
nor U1272 (N_1272,N_56,N_98);
or U1273 (N_1273,N_259,N_343);
xor U1274 (N_1274,N_235,N_266);
nand U1275 (N_1275,N_558,N_109);
or U1276 (N_1276,N_20,N_65);
nand U1277 (N_1277,N_69,N_24);
nor U1278 (N_1278,N_674,N_347);
nand U1279 (N_1279,N_623,N_234);
and U1280 (N_1280,N_236,N_378);
or U1281 (N_1281,N_3,N_449);
nor U1282 (N_1282,N_630,N_383);
and U1283 (N_1283,N_113,N_610);
nor U1284 (N_1284,N_386,N_296);
nand U1285 (N_1285,N_470,N_309);
or U1286 (N_1286,N_181,N_740);
xor U1287 (N_1287,N_115,N_419);
nand U1288 (N_1288,N_642,N_293);
nor U1289 (N_1289,N_190,N_98);
and U1290 (N_1290,N_294,N_401);
and U1291 (N_1291,N_140,N_375);
nand U1292 (N_1292,N_204,N_117);
or U1293 (N_1293,N_365,N_641);
or U1294 (N_1294,N_507,N_212);
or U1295 (N_1295,N_58,N_667);
nor U1296 (N_1296,N_684,N_563);
or U1297 (N_1297,N_338,N_538);
nor U1298 (N_1298,N_473,N_418);
and U1299 (N_1299,N_196,N_80);
nand U1300 (N_1300,N_362,N_136);
and U1301 (N_1301,N_207,N_78);
nor U1302 (N_1302,N_705,N_392);
or U1303 (N_1303,N_195,N_634);
or U1304 (N_1304,N_699,N_497);
nand U1305 (N_1305,N_353,N_285);
and U1306 (N_1306,N_199,N_65);
and U1307 (N_1307,N_593,N_158);
nor U1308 (N_1308,N_212,N_570);
and U1309 (N_1309,N_582,N_462);
nand U1310 (N_1310,N_190,N_389);
nor U1311 (N_1311,N_513,N_266);
or U1312 (N_1312,N_162,N_197);
nand U1313 (N_1313,N_96,N_216);
or U1314 (N_1314,N_151,N_620);
or U1315 (N_1315,N_265,N_428);
nand U1316 (N_1316,N_559,N_195);
nor U1317 (N_1317,N_141,N_391);
nor U1318 (N_1318,N_641,N_285);
and U1319 (N_1319,N_379,N_537);
and U1320 (N_1320,N_334,N_211);
nand U1321 (N_1321,N_362,N_712);
nand U1322 (N_1322,N_23,N_355);
or U1323 (N_1323,N_466,N_510);
or U1324 (N_1324,N_393,N_564);
or U1325 (N_1325,N_411,N_622);
xnor U1326 (N_1326,N_538,N_647);
or U1327 (N_1327,N_251,N_476);
nand U1328 (N_1328,N_736,N_405);
and U1329 (N_1329,N_599,N_529);
nor U1330 (N_1330,N_312,N_731);
and U1331 (N_1331,N_440,N_481);
and U1332 (N_1332,N_52,N_236);
or U1333 (N_1333,N_650,N_635);
and U1334 (N_1334,N_327,N_150);
or U1335 (N_1335,N_357,N_163);
and U1336 (N_1336,N_143,N_200);
or U1337 (N_1337,N_55,N_361);
and U1338 (N_1338,N_666,N_512);
and U1339 (N_1339,N_619,N_379);
nor U1340 (N_1340,N_364,N_692);
xnor U1341 (N_1341,N_464,N_603);
and U1342 (N_1342,N_644,N_366);
nand U1343 (N_1343,N_193,N_520);
or U1344 (N_1344,N_525,N_396);
xnor U1345 (N_1345,N_285,N_462);
nor U1346 (N_1346,N_472,N_578);
or U1347 (N_1347,N_547,N_246);
xor U1348 (N_1348,N_747,N_201);
nand U1349 (N_1349,N_342,N_583);
nor U1350 (N_1350,N_381,N_64);
nand U1351 (N_1351,N_552,N_261);
nor U1352 (N_1352,N_101,N_411);
nor U1353 (N_1353,N_691,N_117);
xnor U1354 (N_1354,N_218,N_505);
or U1355 (N_1355,N_77,N_100);
and U1356 (N_1356,N_608,N_323);
or U1357 (N_1357,N_743,N_725);
nor U1358 (N_1358,N_314,N_217);
nor U1359 (N_1359,N_82,N_650);
nand U1360 (N_1360,N_676,N_261);
and U1361 (N_1361,N_595,N_472);
or U1362 (N_1362,N_17,N_197);
or U1363 (N_1363,N_135,N_341);
nor U1364 (N_1364,N_606,N_547);
or U1365 (N_1365,N_497,N_119);
nor U1366 (N_1366,N_202,N_59);
nand U1367 (N_1367,N_247,N_560);
and U1368 (N_1368,N_28,N_674);
nand U1369 (N_1369,N_606,N_498);
and U1370 (N_1370,N_28,N_647);
nand U1371 (N_1371,N_184,N_569);
and U1372 (N_1372,N_201,N_185);
nand U1373 (N_1373,N_612,N_375);
or U1374 (N_1374,N_613,N_86);
nand U1375 (N_1375,N_616,N_360);
nand U1376 (N_1376,N_333,N_467);
nand U1377 (N_1377,N_379,N_147);
nor U1378 (N_1378,N_115,N_661);
and U1379 (N_1379,N_273,N_7);
nor U1380 (N_1380,N_690,N_417);
nor U1381 (N_1381,N_630,N_61);
nand U1382 (N_1382,N_209,N_343);
or U1383 (N_1383,N_445,N_318);
nor U1384 (N_1384,N_33,N_12);
and U1385 (N_1385,N_67,N_467);
and U1386 (N_1386,N_670,N_171);
nor U1387 (N_1387,N_619,N_238);
and U1388 (N_1388,N_121,N_167);
nor U1389 (N_1389,N_246,N_421);
nand U1390 (N_1390,N_693,N_111);
nand U1391 (N_1391,N_119,N_594);
or U1392 (N_1392,N_401,N_443);
nor U1393 (N_1393,N_334,N_584);
nand U1394 (N_1394,N_192,N_631);
nor U1395 (N_1395,N_415,N_508);
and U1396 (N_1396,N_729,N_262);
nor U1397 (N_1397,N_733,N_263);
or U1398 (N_1398,N_51,N_741);
nor U1399 (N_1399,N_731,N_522);
and U1400 (N_1400,N_613,N_418);
nand U1401 (N_1401,N_392,N_32);
or U1402 (N_1402,N_16,N_302);
or U1403 (N_1403,N_381,N_243);
nand U1404 (N_1404,N_244,N_679);
xnor U1405 (N_1405,N_440,N_527);
or U1406 (N_1406,N_77,N_286);
xnor U1407 (N_1407,N_620,N_630);
or U1408 (N_1408,N_411,N_77);
nand U1409 (N_1409,N_73,N_556);
xor U1410 (N_1410,N_664,N_462);
and U1411 (N_1411,N_412,N_330);
xor U1412 (N_1412,N_188,N_114);
nand U1413 (N_1413,N_246,N_115);
nor U1414 (N_1414,N_253,N_495);
nand U1415 (N_1415,N_184,N_496);
and U1416 (N_1416,N_622,N_694);
nor U1417 (N_1417,N_540,N_433);
or U1418 (N_1418,N_364,N_721);
or U1419 (N_1419,N_650,N_236);
or U1420 (N_1420,N_224,N_449);
or U1421 (N_1421,N_216,N_184);
and U1422 (N_1422,N_141,N_622);
and U1423 (N_1423,N_38,N_652);
or U1424 (N_1424,N_470,N_393);
or U1425 (N_1425,N_738,N_383);
nand U1426 (N_1426,N_594,N_598);
nand U1427 (N_1427,N_134,N_579);
xnor U1428 (N_1428,N_417,N_19);
and U1429 (N_1429,N_219,N_648);
nand U1430 (N_1430,N_532,N_379);
nand U1431 (N_1431,N_721,N_68);
xnor U1432 (N_1432,N_635,N_181);
nand U1433 (N_1433,N_445,N_595);
nor U1434 (N_1434,N_479,N_76);
nor U1435 (N_1435,N_672,N_518);
xor U1436 (N_1436,N_312,N_49);
nor U1437 (N_1437,N_746,N_187);
nor U1438 (N_1438,N_680,N_431);
nand U1439 (N_1439,N_119,N_3);
and U1440 (N_1440,N_75,N_590);
nor U1441 (N_1441,N_296,N_635);
nand U1442 (N_1442,N_456,N_203);
and U1443 (N_1443,N_498,N_345);
nand U1444 (N_1444,N_402,N_366);
or U1445 (N_1445,N_22,N_563);
and U1446 (N_1446,N_456,N_130);
xor U1447 (N_1447,N_238,N_191);
nand U1448 (N_1448,N_612,N_366);
nand U1449 (N_1449,N_182,N_650);
or U1450 (N_1450,N_153,N_638);
or U1451 (N_1451,N_531,N_346);
or U1452 (N_1452,N_467,N_65);
nand U1453 (N_1453,N_749,N_462);
nor U1454 (N_1454,N_104,N_338);
xor U1455 (N_1455,N_375,N_383);
or U1456 (N_1456,N_477,N_633);
and U1457 (N_1457,N_14,N_52);
or U1458 (N_1458,N_466,N_58);
nand U1459 (N_1459,N_391,N_62);
and U1460 (N_1460,N_657,N_268);
or U1461 (N_1461,N_285,N_4);
nor U1462 (N_1462,N_501,N_118);
nor U1463 (N_1463,N_524,N_643);
or U1464 (N_1464,N_636,N_287);
or U1465 (N_1465,N_7,N_628);
nor U1466 (N_1466,N_419,N_657);
nor U1467 (N_1467,N_244,N_692);
or U1468 (N_1468,N_430,N_325);
nand U1469 (N_1469,N_511,N_326);
or U1470 (N_1470,N_697,N_647);
nor U1471 (N_1471,N_428,N_699);
xor U1472 (N_1472,N_362,N_655);
nand U1473 (N_1473,N_416,N_737);
nor U1474 (N_1474,N_702,N_303);
or U1475 (N_1475,N_705,N_116);
xnor U1476 (N_1476,N_296,N_713);
or U1477 (N_1477,N_234,N_338);
nand U1478 (N_1478,N_190,N_540);
or U1479 (N_1479,N_172,N_232);
or U1480 (N_1480,N_481,N_727);
nor U1481 (N_1481,N_304,N_646);
nor U1482 (N_1482,N_335,N_501);
nand U1483 (N_1483,N_451,N_222);
or U1484 (N_1484,N_502,N_328);
and U1485 (N_1485,N_340,N_506);
and U1486 (N_1486,N_320,N_326);
or U1487 (N_1487,N_152,N_241);
nor U1488 (N_1488,N_576,N_264);
xor U1489 (N_1489,N_140,N_245);
or U1490 (N_1490,N_683,N_202);
or U1491 (N_1491,N_647,N_195);
or U1492 (N_1492,N_516,N_54);
and U1493 (N_1493,N_326,N_665);
nor U1494 (N_1494,N_64,N_647);
nand U1495 (N_1495,N_77,N_559);
nor U1496 (N_1496,N_593,N_739);
and U1497 (N_1497,N_576,N_457);
and U1498 (N_1498,N_530,N_375);
and U1499 (N_1499,N_658,N_259);
nand U1500 (N_1500,N_1138,N_1434);
xnor U1501 (N_1501,N_1173,N_1134);
nor U1502 (N_1502,N_1277,N_1128);
nand U1503 (N_1503,N_1405,N_1337);
xnor U1504 (N_1504,N_1169,N_1211);
nand U1505 (N_1505,N_1376,N_1265);
nand U1506 (N_1506,N_961,N_786);
nor U1507 (N_1507,N_919,N_1175);
xor U1508 (N_1508,N_1327,N_962);
xnor U1509 (N_1509,N_1331,N_1329);
or U1510 (N_1510,N_772,N_1479);
and U1511 (N_1511,N_1308,N_1143);
nand U1512 (N_1512,N_1037,N_1170);
and U1513 (N_1513,N_1245,N_1416);
nand U1514 (N_1514,N_1412,N_1157);
nand U1515 (N_1515,N_1466,N_967);
nor U1516 (N_1516,N_872,N_1436);
nand U1517 (N_1517,N_1283,N_1088);
nor U1518 (N_1518,N_1156,N_1046);
or U1519 (N_1519,N_1125,N_1028);
xnor U1520 (N_1520,N_1368,N_1290);
or U1521 (N_1521,N_1340,N_1389);
or U1522 (N_1522,N_1034,N_1262);
nor U1523 (N_1523,N_1172,N_1094);
and U1524 (N_1524,N_750,N_911);
nor U1525 (N_1525,N_769,N_809);
nor U1526 (N_1526,N_802,N_1189);
xnor U1527 (N_1527,N_1190,N_878);
nand U1528 (N_1528,N_1375,N_1266);
or U1529 (N_1529,N_1067,N_1310);
and U1530 (N_1530,N_818,N_814);
and U1531 (N_1531,N_1196,N_1379);
and U1532 (N_1532,N_935,N_773);
nor U1533 (N_1533,N_965,N_850);
and U1534 (N_1534,N_885,N_980);
or U1535 (N_1535,N_867,N_1124);
or U1536 (N_1536,N_1394,N_1033);
nor U1537 (N_1537,N_797,N_1314);
nor U1538 (N_1538,N_763,N_1141);
nand U1539 (N_1539,N_1123,N_1309);
and U1540 (N_1540,N_842,N_1038);
and U1541 (N_1541,N_1035,N_1241);
nand U1542 (N_1542,N_1366,N_1261);
and U1543 (N_1543,N_1263,N_1027);
xnor U1544 (N_1544,N_1091,N_778);
nand U1545 (N_1545,N_1455,N_1364);
or U1546 (N_1546,N_840,N_959);
nor U1547 (N_1547,N_1470,N_790);
nand U1548 (N_1548,N_1185,N_1054);
or U1549 (N_1549,N_1361,N_906);
nand U1550 (N_1550,N_1279,N_1484);
nand U1551 (N_1551,N_875,N_1199);
or U1552 (N_1552,N_1163,N_1159);
nand U1553 (N_1553,N_1025,N_902);
nand U1554 (N_1554,N_1451,N_1116);
and U1555 (N_1555,N_1428,N_1312);
and U1556 (N_1556,N_836,N_1282);
or U1557 (N_1557,N_1139,N_1118);
nor U1558 (N_1558,N_1042,N_1306);
or U1559 (N_1559,N_981,N_1051);
nor U1560 (N_1560,N_1005,N_1435);
xnor U1561 (N_1561,N_1338,N_1256);
and U1562 (N_1562,N_1002,N_1334);
or U1563 (N_1563,N_1475,N_1017);
nand U1564 (N_1564,N_1465,N_1221);
and U1565 (N_1565,N_1131,N_1267);
nor U1566 (N_1566,N_939,N_1460);
nand U1567 (N_1567,N_1145,N_1235);
nor U1568 (N_1568,N_1212,N_1010);
xnor U1569 (N_1569,N_1358,N_1371);
xor U1570 (N_1570,N_1392,N_1083);
nand U1571 (N_1571,N_851,N_1127);
or U1572 (N_1572,N_1024,N_983);
nand U1573 (N_1573,N_1441,N_865);
nand U1574 (N_1574,N_1209,N_1430);
or U1575 (N_1575,N_1440,N_1233);
and U1576 (N_1576,N_1359,N_1050);
nor U1577 (N_1577,N_1158,N_990);
nand U1578 (N_1578,N_1437,N_770);
nor U1579 (N_1579,N_905,N_1087);
nor U1580 (N_1580,N_1365,N_776);
nor U1581 (N_1581,N_1213,N_1269);
xnor U1582 (N_1582,N_1275,N_1075);
nand U1583 (N_1583,N_751,N_1220);
or U1584 (N_1584,N_1286,N_1150);
nor U1585 (N_1585,N_1208,N_1008);
xor U1586 (N_1586,N_1488,N_1178);
nand U1587 (N_1587,N_799,N_767);
nand U1588 (N_1588,N_971,N_1302);
nand U1589 (N_1589,N_888,N_815);
nand U1590 (N_1590,N_958,N_1203);
nand U1591 (N_1591,N_995,N_1102);
or U1592 (N_1592,N_834,N_1106);
nor U1593 (N_1593,N_1298,N_1176);
or U1594 (N_1594,N_833,N_937);
nor U1595 (N_1595,N_1372,N_1278);
nand U1596 (N_1596,N_795,N_792);
and U1597 (N_1597,N_1003,N_1184);
or U1598 (N_1598,N_1179,N_774);
nand U1599 (N_1599,N_828,N_789);
nand U1600 (N_1600,N_942,N_869);
nor U1601 (N_1601,N_926,N_913);
or U1602 (N_1602,N_1093,N_1273);
nand U1603 (N_1603,N_994,N_1349);
nor U1604 (N_1604,N_1432,N_1036);
nor U1605 (N_1605,N_969,N_859);
or U1606 (N_1606,N_1154,N_783);
nand U1607 (N_1607,N_1360,N_963);
and U1608 (N_1608,N_825,N_811);
nor U1609 (N_1609,N_912,N_1070);
nand U1610 (N_1610,N_823,N_812);
nor U1611 (N_1611,N_1194,N_1201);
and U1612 (N_1612,N_1255,N_753);
nor U1613 (N_1613,N_1498,N_1121);
and U1614 (N_1614,N_1322,N_943);
or U1615 (N_1615,N_1226,N_766);
and U1616 (N_1616,N_1292,N_1272);
nand U1617 (N_1617,N_757,N_1369);
and U1618 (N_1618,N_1271,N_1490);
or U1619 (N_1619,N_793,N_866);
and U1620 (N_1620,N_982,N_1403);
nor U1621 (N_1621,N_1242,N_1231);
or U1622 (N_1622,N_1078,N_1107);
nand U1623 (N_1623,N_1096,N_1496);
and U1624 (N_1624,N_1210,N_1200);
nand U1625 (N_1625,N_827,N_987);
nand U1626 (N_1626,N_1223,N_803);
or U1627 (N_1627,N_1377,N_861);
nor U1628 (N_1628,N_1383,N_933);
and U1629 (N_1629,N_1120,N_1464);
or U1630 (N_1630,N_893,N_1069);
nor U1631 (N_1631,N_904,N_908);
and U1632 (N_1632,N_765,N_1165);
xor U1633 (N_1633,N_1487,N_1420);
xor U1634 (N_1634,N_1012,N_921);
and U1635 (N_1635,N_1296,N_1014);
and U1636 (N_1636,N_1022,N_974);
xnor U1637 (N_1637,N_1344,N_1135);
nand U1638 (N_1638,N_972,N_991);
or U1639 (N_1639,N_1300,N_891);
or U1640 (N_1640,N_1007,N_1459);
or U1641 (N_1641,N_1030,N_1342);
and U1642 (N_1642,N_1395,N_1324);
xor U1643 (N_1643,N_1063,N_1445);
or U1644 (N_1644,N_762,N_779);
nor U1645 (N_1645,N_955,N_1048);
nand U1646 (N_1646,N_1414,N_756);
xor U1647 (N_1647,N_1071,N_1187);
xnor U1648 (N_1648,N_1426,N_915);
nand U1649 (N_1649,N_1239,N_985);
xor U1650 (N_1650,N_929,N_1381);
or U1651 (N_1651,N_1077,N_761);
or U1652 (N_1652,N_832,N_1418);
xor U1653 (N_1653,N_830,N_1476);
or U1654 (N_1654,N_1080,N_852);
xnor U1655 (N_1655,N_1243,N_1444);
nor U1656 (N_1656,N_1152,N_816);
or U1657 (N_1657,N_973,N_979);
nand U1658 (N_1658,N_1164,N_1373);
nand U1659 (N_1659,N_1244,N_1061);
and U1660 (N_1660,N_1354,N_791);
or U1661 (N_1661,N_993,N_1076);
xor U1662 (N_1662,N_1313,N_794);
nand U1663 (N_1663,N_1317,N_1497);
or U1664 (N_1664,N_1227,N_1425);
or U1665 (N_1665,N_996,N_1055);
or U1666 (N_1666,N_934,N_1422);
nor U1667 (N_1667,N_847,N_1174);
nor U1668 (N_1668,N_1433,N_1264);
or U1669 (N_1669,N_1291,N_835);
nand U1670 (N_1670,N_1068,N_1204);
and U1671 (N_1671,N_810,N_1238);
or U1672 (N_1672,N_1029,N_1321);
and U1673 (N_1673,N_752,N_947);
nand U1674 (N_1674,N_1085,N_831);
nand U1675 (N_1675,N_760,N_1147);
nand U1676 (N_1676,N_1011,N_1251);
nor U1677 (N_1677,N_1463,N_821);
xor U1678 (N_1678,N_845,N_1431);
nand U1679 (N_1679,N_870,N_805);
nand U1680 (N_1680,N_1177,N_975);
or U1681 (N_1681,N_1452,N_1108);
nor U1682 (N_1682,N_1112,N_998);
or U1683 (N_1683,N_862,N_1016);
nor U1684 (N_1684,N_1316,N_1408);
nand U1685 (N_1685,N_978,N_820);
and U1686 (N_1686,N_1181,N_1253);
nor U1687 (N_1687,N_1350,N_1442);
or U1688 (N_1688,N_918,N_1393);
xor U1689 (N_1689,N_754,N_1319);
or U1690 (N_1690,N_1336,N_1396);
nand U1691 (N_1691,N_1443,N_1098);
nor U1692 (N_1692,N_1104,N_1215);
and U1693 (N_1693,N_1032,N_1473);
and U1694 (N_1694,N_819,N_1406);
nor U1695 (N_1695,N_1374,N_1402);
or U1696 (N_1696,N_1000,N_1191);
nor U1697 (N_1697,N_843,N_1391);
nor U1698 (N_1698,N_1398,N_1301);
nor U1699 (N_1699,N_922,N_1467);
xor U1700 (N_1700,N_1474,N_1031);
or U1701 (N_1701,N_1217,N_920);
nor U1702 (N_1702,N_804,N_1384);
and U1703 (N_1703,N_1260,N_1328);
or U1704 (N_1704,N_1456,N_1491);
nand U1705 (N_1705,N_829,N_780);
or U1706 (N_1706,N_1399,N_903);
nand U1707 (N_1707,N_964,N_781);
nor U1708 (N_1708,N_1045,N_1161);
or U1709 (N_1709,N_1224,N_857);
nor U1710 (N_1710,N_1285,N_1343);
and U1711 (N_1711,N_1400,N_916);
nand U1712 (N_1712,N_1348,N_1449);
nand U1713 (N_1713,N_1270,N_897);
or U1714 (N_1714,N_1424,N_1018);
or U1715 (N_1715,N_1132,N_989);
nand U1716 (N_1716,N_1198,N_1234);
or U1717 (N_1717,N_1380,N_1186);
or U1718 (N_1718,N_1295,N_940);
and U1719 (N_1719,N_1129,N_1142);
or U1720 (N_1720,N_1257,N_1289);
nand U1721 (N_1721,N_927,N_1228);
xor U1722 (N_1722,N_1304,N_945);
and U1723 (N_1723,N_1130,N_952);
nand U1724 (N_1724,N_1341,N_1356);
or U1725 (N_1725,N_1252,N_1081);
nor U1726 (N_1726,N_1240,N_1453);
nor U1727 (N_1727,N_1023,N_1280);
nor U1728 (N_1728,N_1494,N_907);
and U1729 (N_1729,N_1387,N_1458);
xnor U1730 (N_1730,N_1049,N_1472);
and U1731 (N_1731,N_1439,N_1237);
or U1732 (N_1732,N_1462,N_1345);
and U1733 (N_1733,N_1454,N_839);
nor U1734 (N_1734,N_1074,N_1183);
nand U1735 (N_1735,N_771,N_1318);
xor U1736 (N_1736,N_941,N_899);
nand U1737 (N_1737,N_1288,N_858);
and U1738 (N_1738,N_1407,N_1415);
or U1739 (N_1739,N_1307,N_1346);
nor U1740 (N_1740,N_1254,N_1044);
and U1741 (N_1741,N_854,N_1409);
nor U1742 (N_1742,N_1060,N_1249);
nor U1743 (N_1743,N_898,N_1362);
or U1744 (N_1744,N_1168,N_1079);
or U1745 (N_1745,N_889,N_853);
nand U1746 (N_1746,N_1137,N_1281);
xor U1747 (N_1747,N_1073,N_877);
and U1748 (N_1748,N_1485,N_1378);
or U1749 (N_1749,N_1248,N_838);
nand U1750 (N_1750,N_887,N_1493);
or U1751 (N_1751,N_1021,N_1353);
and U1752 (N_1752,N_1047,N_1097);
and U1753 (N_1753,N_879,N_1040);
nor U1754 (N_1754,N_844,N_1064);
xnor U1755 (N_1755,N_1390,N_1236);
or U1756 (N_1756,N_806,N_1122);
or U1757 (N_1757,N_928,N_1193);
nor U1758 (N_1758,N_1188,N_1020);
nand U1759 (N_1759,N_1155,N_1001);
nor U1760 (N_1760,N_1180,N_801);
xnor U1761 (N_1761,N_863,N_1438);
or U1762 (N_1762,N_1325,N_846);
nand U1763 (N_1763,N_1207,N_1065);
and U1764 (N_1764,N_1246,N_1268);
nor U1765 (N_1765,N_798,N_871);
nor U1766 (N_1766,N_1446,N_917);
or U1767 (N_1767,N_949,N_1043);
nand U1768 (N_1768,N_1410,N_759);
and U1769 (N_1769,N_1084,N_986);
nand U1770 (N_1770,N_1287,N_1388);
xor U1771 (N_1771,N_1166,N_1367);
xor U1772 (N_1772,N_785,N_824);
and U1773 (N_1773,N_1247,N_1101);
and U1774 (N_1774,N_923,N_1303);
or U1775 (N_1775,N_1009,N_1469);
nor U1776 (N_1776,N_884,N_1015);
and U1777 (N_1777,N_1053,N_953);
nand U1778 (N_1778,N_1481,N_807);
or U1779 (N_1779,N_1218,N_1330);
nand U1780 (N_1780,N_948,N_1423);
nor U1781 (N_1781,N_1052,N_1401);
or U1782 (N_1782,N_936,N_1447);
nand U1783 (N_1783,N_1105,N_873);
nand U1784 (N_1784,N_1417,N_1450);
or U1785 (N_1785,N_1089,N_868);
nand U1786 (N_1786,N_1351,N_970);
nor U1787 (N_1787,N_1113,N_1483);
xor U1788 (N_1788,N_1214,N_1144);
nor U1789 (N_1789,N_1250,N_896);
nand U1790 (N_1790,N_874,N_957);
and U1791 (N_1791,N_1146,N_1419);
xnor U1792 (N_1792,N_822,N_1352);
and U1793 (N_1793,N_1299,N_1404);
nand U1794 (N_1794,N_1110,N_784);
nand U1795 (N_1795,N_755,N_800);
or U1796 (N_1796,N_1117,N_900);
and U1797 (N_1797,N_880,N_1133);
and U1798 (N_1798,N_1480,N_1323);
or U1799 (N_1799,N_988,N_1222);
nand U1800 (N_1800,N_775,N_1149);
or U1801 (N_1801,N_938,N_1347);
nor U1802 (N_1802,N_1092,N_1284);
nor U1803 (N_1803,N_1039,N_1326);
and U1804 (N_1804,N_890,N_1216);
nor U1805 (N_1805,N_1370,N_1059);
nor U1806 (N_1806,N_1489,N_1206);
and U1807 (N_1807,N_1274,N_977);
and U1808 (N_1808,N_883,N_1448);
nand U1809 (N_1809,N_950,N_1151);
nor U1810 (N_1810,N_1363,N_1495);
and U1811 (N_1811,N_1100,N_910);
nand U1812 (N_1812,N_1357,N_1311);
and U1813 (N_1813,N_1386,N_1197);
or U1814 (N_1814,N_788,N_817);
nor U1815 (N_1815,N_1160,N_976);
nor U1816 (N_1816,N_1294,N_1355);
or U1817 (N_1817,N_1297,N_1192);
and U1818 (N_1818,N_1056,N_1095);
nor U1819 (N_1819,N_1167,N_1305);
xor U1820 (N_1820,N_1006,N_787);
nand U1821 (N_1821,N_1335,N_1195);
and U1822 (N_1822,N_1382,N_1041);
nand U1823 (N_1823,N_1109,N_960);
and U1824 (N_1824,N_1461,N_1468);
nor U1825 (N_1825,N_864,N_1471);
or U1826 (N_1826,N_848,N_1103);
xnor U1827 (N_1827,N_1119,N_1421);
xnor U1828 (N_1828,N_997,N_886);
or U1829 (N_1829,N_1111,N_881);
nor U1830 (N_1830,N_1411,N_1115);
or U1831 (N_1831,N_1230,N_909);
nor U1832 (N_1832,N_956,N_1004);
or U1833 (N_1833,N_1066,N_1232);
and U1834 (N_1834,N_951,N_930);
and U1835 (N_1835,N_1136,N_1153);
and U1836 (N_1836,N_777,N_892);
nor U1837 (N_1837,N_1072,N_1482);
or U1838 (N_1838,N_1333,N_895);
xor U1839 (N_1839,N_1478,N_1219);
and U1840 (N_1840,N_1429,N_1090);
nor U1841 (N_1841,N_1276,N_1332);
xor U1842 (N_1842,N_856,N_992);
or U1843 (N_1843,N_841,N_1019);
nand U1844 (N_1844,N_1140,N_1413);
xor U1845 (N_1845,N_882,N_837);
or U1846 (N_1846,N_966,N_1427);
or U1847 (N_1847,N_1320,N_999);
xor U1848 (N_1848,N_1499,N_1258);
xnor U1849 (N_1849,N_894,N_1385);
and U1850 (N_1850,N_1486,N_808);
nand U1851 (N_1851,N_1086,N_1099);
or U1852 (N_1852,N_925,N_901);
nor U1853 (N_1853,N_1058,N_876);
nand U1854 (N_1854,N_1492,N_1293);
or U1855 (N_1855,N_826,N_1477);
xnor U1856 (N_1856,N_1057,N_1339);
or U1857 (N_1857,N_796,N_1171);
nand U1858 (N_1858,N_782,N_1259);
nor U1859 (N_1859,N_1082,N_1148);
and U1860 (N_1860,N_932,N_855);
nand U1861 (N_1861,N_1114,N_968);
nand U1862 (N_1862,N_1225,N_914);
nand U1863 (N_1863,N_1013,N_1205);
and U1864 (N_1864,N_764,N_1457);
nor U1865 (N_1865,N_768,N_954);
or U1866 (N_1866,N_1026,N_1315);
nor U1867 (N_1867,N_1202,N_758);
and U1868 (N_1868,N_1182,N_946);
or U1869 (N_1869,N_1229,N_1397);
or U1870 (N_1870,N_813,N_1162);
nand U1871 (N_1871,N_924,N_931);
nor U1872 (N_1872,N_944,N_1126);
or U1873 (N_1873,N_860,N_1062);
xnor U1874 (N_1874,N_984,N_849);
nand U1875 (N_1875,N_1371,N_1385);
or U1876 (N_1876,N_843,N_816);
nor U1877 (N_1877,N_1200,N_1039);
and U1878 (N_1878,N_976,N_1130);
xnor U1879 (N_1879,N_1200,N_1010);
nor U1880 (N_1880,N_1219,N_844);
xnor U1881 (N_1881,N_803,N_1367);
or U1882 (N_1882,N_1331,N_1412);
xor U1883 (N_1883,N_1037,N_1151);
nand U1884 (N_1884,N_1474,N_871);
nor U1885 (N_1885,N_1086,N_1125);
nand U1886 (N_1886,N_1476,N_955);
nand U1887 (N_1887,N_1270,N_860);
nor U1888 (N_1888,N_851,N_1311);
or U1889 (N_1889,N_1091,N_1154);
and U1890 (N_1890,N_1126,N_1405);
xnor U1891 (N_1891,N_1172,N_924);
nor U1892 (N_1892,N_940,N_761);
or U1893 (N_1893,N_1259,N_1147);
xor U1894 (N_1894,N_1023,N_850);
nor U1895 (N_1895,N_1488,N_1041);
xor U1896 (N_1896,N_989,N_1384);
nand U1897 (N_1897,N_814,N_1104);
xor U1898 (N_1898,N_1421,N_822);
nor U1899 (N_1899,N_965,N_752);
or U1900 (N_1900,N_1408,N_1436);
nor U1901 (N_1901,N_957,N_792);
nand U1902 (N_1902,N_1212,N_1303);
or U1903 (N_1903,N_1087,N_973);
nand U1904 (N_1904,N_1411,N_996);
nand U1905 (N_1905,N_872,N_1204);
and U1906 (N_1906,N_1321,N_1108);
nor U1907 (N_1907,N_1285,N_1309);
xor U1908 (N_1908,N_1063,N_1242);
nor U1909 (N_1909,N_1076,N_1367);
and U1910 (N_1910,N_904,N_1041);
or U1911 (N_1911,N_984,N_1189);
nor U1912 (N_1912,N_854,N_930);
xnor U1913 (N_1913,N_1047,N_1022);
nand U1914 (N_1914,N_798,N_1332);
or U1915 (N_1915,N_1087,N_1483);
xor U1916 (N_1916,N_912,N_972);
nand U1917 (N_1917,N_969,N_785);
and U1918 (N_1918,N_953,N_976);
nor U1919 (N_1919,N_1468,N_877);
and U1920 (N_1920,N_968,N_863);
and U1921 (N_1921,N_1187,N_1116);
or U1922 (N_1922,N_1451,N_1266);
nor U1923 (N_1923,N_928,N_1208);
nand U1924 (N_1924,N_783,N_913);
nor U1925 (N_1925,N_1480,N_1314);
nor U1926 (N_1926,N_1457,N_935);
or U1927 (N_1927,N_1167,N_915);
and U1928 (N_1928,N_1485,N_838);
or U1929 (N_1929,N_883,N_798);
and U1930 (N_1930,N_1107,N_1124);
and U1931 (N_1931,N_1424,N_783);
nand U1932 (N_1932,N_1318,N_1354);
and U1933 (N_1933,N_874,N_1382);
nand U1934 (N_1934,N_935,N_1379);
xnor U1935 (N_1935,N_1337,N_893);
or U1936 (N_1936,N_1446,N_936);
nand U1937 (N_1937,N_938,N_830);
nor U1938 (N_1938,N_1372,N_1073);
nor U1939 (N_1939,N_996,N_1131);
nand U1940 (N_1940,N_1160,N_1239);
nand U1941 (N_1941,N_1058,N_1421);
and U1942 (N_1942,N_1153,N_859);
and U1943 (N_1943,N_1357,N_1367);
and U1944 (N_1944,N_1175,N_1077);
or U1945 (N_1945,N_986,N_982);
nand U1946 (N_1946,N_1011,N_1239);
nor U1947 (N_1947,N_756,N_1165);
nand U1948 (N_1948,N_1363,N_794);
and U1949 (N_1949,N_809,N_905);
nor U1950 (N_1950,N_935,N_1188);
nand U1951 (N_1951,N_1258,N_1068);
or U1952 (N_1952,N_1078,N_764);
or U1953 (N_1953,N_1121,N_960);
nand U1954 (N_1954,N_1006,N_803);
nand U1955 (N_1955,N_1199,N_983);
nand U1956 (N_1956,N_850,N_1288);
and U1957 (N_1957,N_1411,N_1386);
nand U1958 (N_1958,N_1442,N_1333);
or U1959 (N_1959,N_1397,N_1327);
xnor U1960 (N_1960,N_1194,N_1151);
nor U1961 (N_1961,N_1188,N_1414);
or U1962 (N_1962,N_875,N_1223);
nor U1963 (N_1963,N_1315,N_950);
nor U1964 (N_1964,N_1142,N_971);
nand U1965 (N_1965,N_1207,N_843);
and U1966 (N_1966,N_1101,N_880);
xnor U1967 (N_1967,N_763,N_1273);
nand U1968 (N_1968,N_835,N_1003);
or U1969 (N_1969,N_1495,N_893);
and U1970 (N_1970,N_1199,N_1388);
xor U1971 (N_1971,N_976,N_893);
nand U1972 (N_1972,N_1117,N_994);
xnor U1973 (N_1973,N_992,N_1260);
or U1974 (N_1974,N_1225,N_1170);
or U1975 (N_1975,N_1449,N_1311);
and U1976 (N_1976,N_1452,N_795);
and U1977 (N_1977,N_1333,N_990);
and U1978 (N_1978,N_1194,N_933);
or U1979 (N_1979,N_1102,N_1407);
nor U1980 (N_1980,N_1373,N_1400);
nand U1981 (N_1981,N_1419,N_937);
xor U1982 (N_1982,N_993,N_1305);
nor U1983 (N_1983,N_1393,N_1099);
or U1984 (N_1984,N_963,N_1221);
xor U1985 (N_1985,N_917,N_847);
or U1986 (N_1986,N_1047,N_995);
nor U1987 (N_1987,N_1396,N_1160);
nor U1988 (N_1988,N_1032,N_912);
or U1989 (N_1989,N_1372,N_796);
or U1990 (N_1990,N_1129,N_1170);
nor U1991 (N_1991,N_968,N_1296);
or U1992 (N_1992,N_931,N_964);
nor U1993 (N_1993,N_815,N_1366);
or U1994 (N_1994,N_1185,N_972);
nor U1995 (N_1995,N_1040,N_777);
xnor U1996 (N_1996,N_784,N_972);
nand U1997 (N_1997,N_1485,N_1227);
or U1998 (N_1998,N_1256,N_1193);
and U1999 (N_1999,N_1258,N_1292);
xor U2000 (N_2000,N_1188,N_1455);
and U2001 (N_2001,N_791,N_851);
nand U2002 (N_2002,N_1459,N_769);
nor U2003 (N_2003,N_933,N_789);
nand U2004 (N_2004,N_1206,N_873);
or U2005 (N_2005,N_847,N_891);
nor U2006 (N_2006,N_1046,N_1420);
nor U2007 (N_2007,N_1387,N_1016);
or U2008 (N_2008,N_1144,N_1053);
nor U2009 (N_2009,N_1351,N_1257);
nor U2010 (N_2010,N_1472,N_1312);
nand U2011 (N_2011,N_982,N_975);
nand U2012 (N_2012,N_1147,N_1198);
nand U2013 (N_2013,N_1341,N_885);
nand U2014 (N_2014,N_846,N_1196);
and U2015 (N_2015,N_1112,N_1332);
nand U2016 (N_2016,N_751,N_1485);
nor U2017 (N_2017,N_1219,N_1455);
and U2018 (N_2018,N_1436,N_1437);
nand U2019 (N_2019,N_1282,N_1173);
or U2020 (N_2020,N_1255,N_876);
or U2021 (N_2021,N_813,N_1265);
nor U2022 (N_2022,N_1005,N_838);
and U2023 (N_2023,N_1108,N_1264);
and U2024 (N_2024,N_1397,N_857);
and U2025 (N_2025,N_1053,N_1256);
or U2026 (N_2026,N_913,N_1052);
nor U2027 (N_2027,N_821,N_1445);
nand U2028 (N_2028,N_951,N_1428);
xnor U2029 (N_2029,N_1128,N_884);
xor U2030 (N_2030,N_962,N_937);
and U2031 (N_2031,N_1270,N_1209);
nor U2032 (N_2032,N_954,N_1288);
and U2033 (N_2033,N_1281,N_984);
or U2034 (N_2034,N_793,N_1021);
and U2035 (N_2035,N_1139,N_810);
xnor U2036 (N_2036,N_1186,N_1351);
xnor U2037 (N_2037,N_1084,N_966);
nor U2038 (N_2038,N_1425,N_874);
xnor U2039 (N_2039,N_907,N_1353);
and U2040 (N_2040,N_971,N_1232);
nand U2041 (N_2041,N_1097,N_1263);
nand U2042 (N_2042,N_1246,N_1214);
and U2043 (N_2043,N_1218,N_756);
and U2044 (N_2044,N_917,N_893);
nand U2045 (N_2045,N_979,N_782);
or U2046 (N_2046,N_1472,N_1341);
nand U2047 (N_2047,N_1093,N_1354);
nand U2048 (N_2048,N_1032,N_833);
nand U2049 (N_2049,N_1430,N_1054);
or U2050 (N_2050,N_873,N_1172);
and U2051 (N_2051,N_973,N_950);
nand U2052 (N_2052,N_1224,N_1154);
xor U2053 (N_2053,N_1468,N_826);
and U2054 (N_2054,N_801,N_1280);
nand U2055 (N_2055,N_1483,N_1075);
and U2056 (N_2056,N_1319,N_1133);
and U2057 (N_2057,N_1306,N_1071);
and U2058 (N_2058,N_1268,N_946);
or U2059 (N_2059,N_754,N_1074);
and U2060 (N_2060,N_1300,N_791);
nand U2061 (N_2061,N_1146,N_942);
nand U2062 (N_2062,N_825,N_881);
nand U2063 (N_2063,N_1466,N_825);
and U2064 (N_2064,N_766,N_762);
nand U2065 (N_2065,N_1366,N_965);
nand U2066 (N_2066,N_1463,N_1178);
or U2067 (N_2067,N_1376,N_1169);
nor U2068 (N_2068,N_810,N_1047);
or U2069 (N_2069,N_1236,N_1076);
or U2070 (N_2070,N_893,N_977);
and U2071 (N_2071,N_1071,N_1167);
nor U2072 (N_2072,N_1154,N_1068);
or U2073 (N_2073,N_968,N_940);
nor U2074 (N_2074,N_1029,N_784);
nor U2075 (N_2075,N_961,N_1209);
nand U2076 (N_2076,N_943,N_1253);
or U2077 (N_2077,N_1411,N_1458);
or U2078 (N_2078,N_1118,N_1091);
or U2079 (N_2079,N_1430,N_888);
nor U2080 (N_2080,N_1499,N_903);
and U2081 (N_2081,N_841,N_1048);
or U2082 (N_2082,N_1180,N_1304);
or U2083 (N_2083,N_986,N_909);
xor U2084 (N_2084,N_1488,N_1272);
xnor U2085 (N_2085,N_1124,N_1174);
xnor U2086 (N_2086,N_1228,N_1175);
and U2087 (N_2087,N_952,N_783);
nand U2088 (N_2088,N_1376,N_921);
nand U2089 (N_2089,N_1118,N_1425);
nor U2090 (N_2090,N_1196,N_1136);
nand U2091 (N_2091,N_1427,N_1221);
nand U2092 (N_2092,N_1452,N_1483);
and U2093 (N_2093,N_1041,N_941);
nor U2094 (N_2094,N_1172,N_945);
or U2095 (N_2095,N_1092,N_1303);
and U2096 (N_2096,N_863,N_1172);
and U2097 (N_2097,N_1332,N_1126);
and U2098 (N_2098,N_970,N_1474);
and U2099 (N_2099,N_1125,N_1115);
nand U2100 (N_2100,N_1406,N_940);
xnor U2101 (N_2101,N_1282,N_1360);
or U2102 (N_2102,N_863,N_800);
or U2103 (N_2103,N_1027,N_908);
nor U2104 (N_2104,N_946,N_918);
or U2105 (N_2105,N_1137,N_1041);
nand U2106 (N_2106,N_1086,N_815);
xnor U2107 (N_2107,N_974,N_1483);
and U2108 (N_2108,N_1247,N_1332);
nor U2109 (N_2109,N_1433,N_1321);
nor U2110 (N_2110,N_796,N_837);
or U2111 (N_2111,N_1194,N_1236);
nand U2112 (N_2112,N_1049,N_841);
xnor U2113 (N_2113,N_860,N_945);
nand U2114 (N_2114,N_1477,N_1356);
nor U2115 (N_2115,N_887,N_1301);
and U2116 (N_2116,N_1023,N_1078);
nor U2117 (N_2117,N_1455,N_1035);
and U2118 (N_2118,N_1025,N_1027);
and U2119 (N_2119,N_1161,N_1411);
nor U2120 (N_2120,N_1442,N_965);
nor U2121 (N_2121,N_1182,N_1261);
nor U2122 (N_2122,N_1120,N_930);
xor U2123 (N_2123,N_1060,N_1284);
nand U2124 (N_2124,N_1016,N_1258);
or U2125 (N_2125,N_1473,N_761);
and U2126 (N_2126,N_802,N_776);
and U2127 (N_2127,N_1488,N_1347);
xnor U2128 (N_2128,N_1050,N_863);
and U2129 (N_2129,N_784,N_1222);
nand U2130 (N_2130,N_1320,N_1184);
and U2131 (N_2131,N_913,N_902);
nand U2132 (N_2132,N_1208,N_1040);
nor U2133 (N_2133,N_859,N_1114);
or U2134 (N_2134,N_1121,N_1008);
and U2135 (N_2135,N_951,N_1080);
and U2136 (N_2136,N_759,N_1022);
nand U2137 (N_2137,N_1402,N_1425);
and U2138 (N_2138,N_1325,N_870);
nand U2139 (N_2139,N_782,N_960);
nand U2140 (N_2140,N_1297,N_1060);
or U2141 (N_2141,N_1132,N_1111);
nor U2142 (N_2142,N_1255,N_1439);
nand U2143 (N_2143,N_932,N_868);
xor U2144 (N_2144,N_1278,N_1382);
xnor U2145 (N_2145,N_1473,N_1279);
xnor U2146 (N_2146,N_788,N_1250);
nor U2147 (N_2147,N_856,N_961);
nor U2148 (N_2148,N_1035,N_1125);
and U2149 (N_2149,N_1466,N_1231);
nor U2150 (N_2150,N_839,N_1160);
nor U2151 (N_2151,N_1049,N_832);
nor U2152 (N_2152,N_1109,N_764);
and U2153 (N_2153,N_1132,N_1494);
or U2154 (N_2154,N_1260,N_1256);
and U2155 (N_2155,N_1179,N_1380);
and U2156 (N_2156,N_1041,N_1283);
nand U2157 (N_2157,N_1111,N_969);
and U2158 (N_2158,N_1235,N_1258);
nand U2159 (N_2159,N_781,N_889);
or U2160 (N_2160,N_1062,N_992);
xnor U2161 (N_2161,N_1409,N_1460);
nand U2162 (N_2162,N_1308,N_1093);
xor U2163 (N_2163,N_1498,N_828);
nor U2164 (N_2164,N_1474,N_1359);
xnor U2165 (N_2165,N_1158,N_1041);
nand U2166 (N_2166,N_1270,N_1228);
or U2167 (N_2167,N_1271,N_1371);
nor U2168 (N_2168,N_1185,N_1256);
or U2169 (N_2169,N_915,N_877);
nor U2170 (N_2170,N_1007,N_902);
nand U2171 (N_2171,N_1473,N_1253);
xor U2172 (N_2172,N_1341,N_773);
xnor U2173 (N_2173,N_1351,N_1317);
xnor U2174 (N_2174,N_1378,N_1119);
or U2175 (N_2175,N_1442,N_1363);
xnor U2176 (N_2176,N_863,N_1111);
nand U2177 (N_2177,N_1377,N_938);
and U2178 (N_2178,N_1157,N_1069);
nand U2179 (N_2179,N_1280,N_1275);
nand U2180 (N_2180,N_904,N_1397);
and U2181 (N_2181,N_1296,N_1035);
nand U2182 (N_2182,N_1410,N_1268);
and U2183 (N_2183,N_984,N_1106);
nor U2184 (N_2184,N_1233,N_815);
nor U2185 (N_2185,N_1115,N_1195);
and U2186 (N_2186,N_1046,N_1172);
and U2187 (N_2187,N_904,N_1283);
or U2188 (N_2188,N_1019,N_1412);
nand U2189 (N_2189,N_972,N_1437);
nor U2190 (N_2190,N_766,N_1022);
or U2191 (N_2191,N_1307,N_1051);
nand U2192 (N_2192,N_1223,N_1274);
or U2193 (N_2193,N_754,N_1073);
nor U2194 (N_2194,N_888,N_1481);
or U2195 (N_2195,N_813,N_1214);
nand U2196 (N_2196,N_1270,N_945);
and U2197 (N_2197,N_1407,N_1307);
xnor U2198 (N_2198,N_1309,N_1253);
nand U2199 (N_2199,N_1070,N_780);
nand U2200 (N_2200,N_1083,N_792);
and U2201 (N_2201,N_1078,N_1028);
nor U2202 (N_2202,N_1497,N_1098);
nand U2203 (N_2203,N_1418,N_1033);
or U2204 (N_2204,N_842,N_874);
nor U2205 (N_2205,N_1493,N_1216);
and U2206 (N_2206,N_952,N_1230);
nand U2207 (N_2207,N_1439,N_1250);
nand U2208 (N_2208,N_897,N_1067);
xor U2209 (N_2209,N_925,N_1132);
and U2210 (N_2210,N_1409,N_1339);
and U2211 (N_2211,N_1204,N_1233);
or U2212 (N_2212,N_1432,N_1425);
and U2213 (N_2213,N_1441,N_1044);
and U2214 (N_2214,N_1381,N_897);
and U2215 (N_2215,N_1462,N_1289);
or U2216 (N_2216,N_998,N_913);
nor U2217 (N_2217,N_1368,N_874);
or U2218 (N_2218,N_1067,N_1368);
or U2219 (N_2219,N_1397,N_1242);
nand U2220 (N_2220,N_1390,N_1275);
nand U2221 (N_2221,N_1342,N_1122);
nor U2222 (N_2222,N_1217,N_1194);
or U2223 (N_2223,N_1314,N_1202);
nand U2224 (N_2224,N_1019,N_1227);
nor U2225 (N_2225,N_1128,N_1241);
and U2226 (N_2226,N_1324,N_914);
and U2227 (N_2227,N_896,N_994);
or U2228 (N_2228,N_1156,N_1376);
nand U2229 (N_2229,N_1353,N_852);
nor U2230 (N_2230,N_1041,N_867);
or U2231 (N_2231,N_1297,N_810);
xnor U2232 (N_2232,N_754,N_1382);
and U2233 (N_2233,N_943,N_1300);
and U2234 (N_2234,N_829,N_1384);
xor U2235 (N_2235,N_1114,N_1188);
or U2236 (N_2236,N_1273,N_909);
nor U2237 (N_2237,N_1087,N_1239);
or U2238 (N_2238,N_1420,N_1159);
nand U2239 (N_2239,N_1181,N_976);
or U2240 (N_2240,N_1177,N_1377);
and U2241 (N_2241,N_1164,N_1030);
and U2242 (N_2242,N_774,N_759);
xor U2243 (N_2243,N_1131,N_968);
nand U2244 (N_2244,N_1238,N_1333);
nand U2245 (N_2245,N_1439,N_1343);
xnor U2246 (N_2246,N_1034,N_1036);
xnor U2247 (N_2247,N_1200,N_1155);
xnor U2248 (N_2248,N_1073,N_1418);
or U2249 (N_2249,N_1089,N_1368);
or U2250 (N_2250,N_1896,N_1878);
nand U2251 (N_2251,N_1611,N_2220);
nand U2252 (N_2252,N_1723,N_1979);
nand U2253 (N_2253,N_2120,N_1883);
or U2254 (N_2254,N_2238,N_2040);
nand U2255 (N_2255,N_2097,N_1625);
nand U2256 (N_2256,N_2160,N_1514);
or U2257 (N_2257,N_2043,N_1973);
nor U2258 (N_2258,N_2231,N_2065);
or U2259 (N_2259,N_1686,N_1811);
and U2260 (N_2260,N_1513,N_1732);
and U2261 (N_2261,N_1673,N_2016);
nor U2262 (N_2262,N_1537,N_2113);
or U2263 (N_2263,N_1738,N_1947);
nor U2264 (N_2264,N_1808,N_1755);
and U2265 (N_2265,N_2055,N_2123);
nor U2266 (N_2266,N_1785,N_1605);
and U2267 (N_2267,N_1781,N_1921);
nor U2268 (N_2268,N_1532,N_1610);
and U2269 (N_2269,N_2006,N_1580);
and U2270 (N_2270,N_1666,N_1671);
or U2271 (N_2271,N_1850,N_2083);
or U2272 (N_2272,N_1775,N_2102);
and U2273 (N_2273,N_2101,N_2186);
or U2274 (N_2274,N_2202,N_1680);
and U2275 (N_2275,N_2165,N_1710);
or U2276 (N_2276,N_1857,N_1578);
nand U2277 (N_2277,N_1750,N_1587);
nor U2278 (N_2278,N_2227,N_1980);
xnor U2279 (N_2279,N_2201,N_2214);
nor U2280 (N_2280,N_1915,N_1655);
and U2281 (N_2281,N_1676,N_1527);
nor U2282 (N_2282,N_2076,N_2094);
and U2283 (N_2283,N_2082,N_1562);
nand U2284 (N_2284,N_1839,N_2229);
and U2285 (N_2285,N_1830,N_1805);
nor U2286 (N_2286,N_1734,N_1862);
nand U2287 (N_2287,N_2012,N_1638);
nor U2288 (N_2288,N_2090,N_1739);
and U2289 (N_2289,N_1520,N_1909);
nand U2290 (N_2290,N_1692,N_1945);
nand U2291 (N_2291,N_1586,N_1913);
or U2292 (N_2292,N_1927,N_2169);
nor U2293 (N_2293,N_1563,N_1963);
xor U2294 (N_2294,N_2004,N_2206);
nor U2295 (N_2295,N_1847,N_2033);
and U2296 (N_2296,N_1794,N_1911);
and U2297 (N_2297,N_1737,N_2019);
xor U2298 (N_2298,N_1953,N_2026);
and U2299 (N_2299,N_2086,N_1841);
xnor U2300 (N_2300,N_2167,N_2177);
and U2301 (N_2301,N_2173,N_1869);
or U2302 (N_2302,N_1637,N_2152);
and U2303 (N_2303,N_1623,N_1541);
nand U2304 (N_2304,N_1659,N_2241);
nand U2305 (N_2305,N_1906,N_1925);
or U2306 (N_2306,N_1698,N_2091);
nor U2307 (N_2307,N_2014,N_1531);
nor U2308 (N_2308,N_2068,N_1974);
nand U2309 (N_2309,N_2158,N_1989);
and U2310 (N_2310,N_2081,N_2233);
and U2311 (N_2311,N_1622,N_1855);
or U2312 (N_2312,N_2045,N_1823);
or U2313 (N_2313,N_1860,N_2242);
nor U2314 (N_2314,N_2213,N_1813);
nor U2315 (N_2315,N_1842,N_2212);
and U2316 (N_2316,N_1929,N_1547);
nor U2317 (N_2317,N_1517,N_1505);
nand U2318 (N_2318,N_2017,N_2039);
nand U2319 (N_2319,N_1511,N_2168);
nand U2320 (N_2320,N_2072,N_1814);
or U2321 (N_2321,N_1589,N_1771);
nor U2322 (N_2322,N_1539,N_1669);
and U2323 (N_2323,N_1995,N_1590);
and U2324 (N_2324,N_1645,N_1624);
and U2325 (N_2325,N_2194,N_1566);
nand U2326 (N_2326,N_1954,N_2023);
nand U2327 (N_2327,N_1536,N_2042);
nor U2328 (N_2328,N_1978,N_2190);
nor U2329 (N_2329,N_1933,N_2125);
nand U2330 (N_2330,N_1772,N_1993);
and U2331 (N_2331,N_1728,N_1786);
nand U2332 (N_2332,N_1821,N_1962);
and U2333 (N_2333,N_1773,N_1957);
or U2334 (N_2334,N_1608,N_1903);
xnor U2335 (N_2335,N_2156,N_2003);
nor U2336 (N_2336,N_1678,N_1726);
xor U2337 (N_2337,N_1971,N_1573);
nor U2338 (N_2338,N_2029,N_1657);
and U2339 (N_2339,N_2216,N_1508);
nor U2340 (N_2340,N_2184,N_1658);
nand U2341 (N_2341,N_2185,N_1546);
or U2342 (N_2342,N_1932,N_1885);
nand U2343 (N_2343,N_2234,N_1717);
nor U2344 (N_2344,N_1549,N_2096);
or U2345 (N_2345,N_1618,N_1684);
nor U2346 (N_2346,N_1922,N_1572);
and U2347 (N_2347,N_1900,N_1583);
or U2348 (N_2348,N_1644,N_1631);
or U2349 (N_2349,N_2144,N_1790);
nor U2350 (N_2350,N_1606,N_2073);
and U2351 (N_2351,N_1747,N_1859);
or U2352 (N_2352,N_1822,N_1597);
or U2353 (N_2353,N_2232,N_2215);
and U2354 (N_2354,N_1665,N_1877);
xnor U2355 (N_2355,N_1695,N_2187);
xor U2356 (N_2356,N_2163,N_1970);
and U2357 (N_2357,N_1584,N_1554);
or U2358 (N_2358,N_1820,N_1891);
nor U2359 (N_2359,N_1735,N_1986);
and U2360 (N_2360,N_1565,N_2151);
or U2361 (N_2361,N_2209,N_1793);
nand U2362 (N_2362,N_1519,N_2041);
nand U2363 (N_2363,N_2075,N_1769);
and U2364 (N_2364,N_1512,N_1682);
xor U2365 (N_2365,N_1600,N_1670);
nor U2366 (N_2366,N_2219,N_1942);
nor U2367 (N_2367,N_1715,N_1708);
and U2368 (N_2368,N_2166,N_2188);
and U2369 (N_2369,N_1568,N_1705);
xor U2370 (N_2370,N_1592,N_1627);
or U2371 (N_2371,N_2221,N_1579);
nand U2372 (N_2372,N_1526,N_2106);
nand U2373 (N_2373,N_2007,N_1881);
nand U2374 (N_2374,N_2115,N_1588);
nor U2375 (N_2375,N_1540,N_1660);
and U2376 (N_2376,N_1843,N_1873);
nor U2377 (N_2377,N_1743,N_1742);
or U2378 (N_2378,N_2174,N_2074);
and U2379 (N_2379,N_1696,N_1902);
or U2380 (N_2380,N_1522,N_2189);
or U2381 (N_2381,N_2129,N_1654);
nor U2382 (N_2382,N_2009,N_1560);
nor U2383 (N_2383,N_2181,N_1690);
and U2384 (N_2384,N_1712,N_1809);
or U2385 (N_2385,N_2024,N_2226);
xor U2386 (N_2386,N_2248,N_2058);
nor U2387 (N_2387,N_2149,N_1762);
nor U2388 (N_2388,N_2103,N_1561);
xnor U2389 (N_2389,N_1817,N_2133);
xnor U2390 (N_2390,N_2031,N_2235);
nor U2391 (N_2391,N_1534,N_1949);
xor U2392 (N_2392,N_1761,N_2059);
nand U2393 (N_2393,N_2048,N_1567);
and U2394 (N_2394,N_1694,N_1509);
nand U2395 (N_2395,N_2228,N_2067);
nor U2396 (N_2396,N_2246,N_2161);
nor U2397 (N_2397,N_1754,N_2150);
nand U2398 (N_2398,N_2010,N_1888);
nand U2399 (N_2399,N_1577,N_2128);
and U2400 (N_2400,N_2092,N_2157);
and U2401 (N_2401,N_1550,N_1542);
nor U2402 (N_2402,N_1991,N_1864);
and U2403 (N_2403,N_1976,N_1685);
xor U2404 (N_2404,N_1713,N_1551);
and U2405 (N_2405,N_1535,N_1525);
and U2406 (N_2406,N_1866,N_1759);
nor U2407 (N_2407,N_1745,N_1730);
or U2408 (N_2408,N_2062,N_2028);
nor U2409 (N_2409,N_2047,N_2183);
nand U2410 (N_2410,N_2119,N_1961);
nand U2411 (N_2411,N_1760,N_1788);
or U2412 (N_2412,N_1722,N_2192);
nor U2413 (N_2413,N_1643,N_2105);
and U2414 (N_2414,N_1774,N_2225);
or U2415 (N_2415,N_1870,N_1581);
nor U2416 (N_2416,N_1634,N_1895);
and U2417 (N_2417,N_1603,N_2180);
nor U2418 (N_2418,N_1596,N_1765);
nand U2419 (N_2419,N_1854,N_2176);
or U2420 (N_2420,N_1867,N_1557);
or U2421 (N_2421,N_2222,N_1663);
or U2422 (N_2422,N_1683,N_1799);
xnor U2423 (N_2423,N_1832,N_2032);
and U2424 (N_2424,N_2104,N_1656);
xor U2425 (N_2425,N_1844,N_1751);
nor U2426 (N_2426,N_1829,N_1892);
xnor U2427 (N_2427,N_1714,N_2122);
nor U2428 (N_2428,N_1782,N_2138);
nand U2429 (N_2429,N_1770,N_1731);
and U2430 (N_2430,N_1604,N_1806);
xor U2431 (N_2431,N_1912,N_1894);
nor U2432 (N_2432,N_1803,N_1956);
and U2433 (N_2433,N_1601,N_2197);
and U2434 (N_2434,N_1516,N_1958);
or U2435 (N_2435,N_1836,N_1834);
or U2436 (N_2436,N_1874,N_2118);
or U2437 (N_2437,N_1530,N_2239);
and U2438 (N_2438,N_1727,N_2036);
nor U2439 (N_2439,N_1807,N_1648);
xnor U2440 (N_2440,N_2069,N_2063);
xnor U2441 (N_2441,N_1777,N_1640);
nand U2442 (N_2442,N_1649,N_1652);
and U2443 (N_2443,N_2098,N_1575);
nand U2444 (N_2444,N_1826,N_2143);
or U2445 (N_2445,N_1591,N_1865);
or U2446 (N_2446,N_1944,N_1545);
and U2447 (N_2447,N_1642,N_1987);
or U2448 (N_2448,N_2035,N_2095);
nand U2449 (N_2449,N_1948,N_1619);
xnor U2450 (N_2450,N_1917,N_1992);
nor U2451 (N_2451,N_1798,N_1897);
nor U2452 (N_2452,N_1964,N_1941);
nand U2453 (N_2453,N_1524,N_1982);
or U2454 (N_2454,N_1548,N_1898);
or U2455 (N_2455,N_1628,N_1981);
or U2456 (N_2456,N_1882,N_1975);
xor U2457 (N_2457,N_1521,N_1967);
nand U2458 (N_2458,N_1955,N_1620);
or U2459 (N_2459,N_2030,N_2005);
nor U2460 (N_2460,N_1688,N_1939);
or U2461 (N_2461,N_2205,N_1965);
nor U2462 (N_2462,N_1996,N_1776);
nand U2463 (N_2463,N_2175,N_1740);
and U2464 (N_2464,N_1585,N_2116);
or U2465 (N_2465,N_1647,N_1636);
and U2466 (N_2466,N_1543,N_2025);
and U2467 (N_2467,N_1752,N_2146);
and U2468 (N_2468,N_1852,N_2114);
or U2469 (N_2469,N_2085,N_1664);
and U2470 (N_2470,N_1691,N_2195);
or U2471 (N_2471,N_1693,N_2100);
xnor U2472 (N_2472,N_2211,N_1632);
nor U2473 (N_2473,N_2093,N_1923);
and U2474 (N_2474,N_1748,N_1880);
and U2475 (N_2475,N_1667,N_2162);
nand U2476 (N_2476,N_2132,N_1668);
or U2477 (N_2477,N_2008,N_2070);
and U2478 (N_2478,N_1582,N_1838);
nor U2479 (N_2479,N_2249,N_1950);
or U2480 (N_2480,N_2139,N_2134);
nand U2481 (N_2481,N_1598,N_1812);
nand U2482 (N_2482,N_1946,N_2053);
and U2483 (N_2483,N_1501,N_2049);
nor U2484 (N_2484,N_1746,N_1528);
and U2485 (N_2485,N_1884,N_1679);
and U2486 (N_2486,N_2204,N_1571);
and U2487 (N_2487,N_1818,N_1612);
or U2488 (N_2488,N_1661,N_2127);
nand U2489 (N_2489,N_1502,N_2099);
nand U2490 (N_2490,N_2145,N_1766);
nor U2491 (N_2491,N_1791,N_2038);
or U2492 (N_2492,N_1983,N_1633);
xor U2493 (N_2493,N_2223,N_1651);
nand U2494 (N_2494,N_1988,N_2247);
or U2495 (N_2495,N_2061,N_2018);
nand U2496 (N_2496,N_2137,N_2064);
nor U2497 (N_2497,N_1778,N_1675);
nand U2498 (N_2498,N_1700,N_1506);
or U2499 (N_2499,N_2140,N_2022);
and U2500 (N_2500,N_1699,N_1901);
nor U2501 (N_2501,N_1662,N_1890);
nor U2502 (N_2502,N_1827,N_1707);
or U2503 (N_2503,N_2046,N_1966);
and U2504 (N_2504,N_2027,N_1763);
and U2505 (N_2505,N_1926,N_2164);
xnor U2506 (N_2506,N_2142,N_1756);
nand U2507 (N_2507,N_1825,N_2111);
xnor U2508 (N_2508,N_1507,N_1599);
or U2509 (N_2509,N_1609,N_1614);
nand U2510 (N_2510,N_1630,N_1701);
or U2511 (N_2511,N_2131,N_1674);
xnor U2512 (N_2512,N_1984,N_1709);
or U2513 (N_2513,N_2178,N_1510);
nand U2514 (N_2514,N_1617,N_1783);
and U2515 (N_2515,N_1908,N_1621);
xor U2516 (N_2516,N_1990,N_2060);
or U2517 (N_2517,N_2191,N_2210);
or U2518 (N_2518,N_1943,N_2237);
nor U2519 (N_2519,N_1960,N_2208);
nor U2520 (N_2520,N_1515,N_1792);
xor U2521 (N_2521,N_1907,N_2148);
nor U2522 (N_2522,N_1780,N_2001);
xor U2523 (N_2523,N_2236,N_1858);
nor U2524 (N_2524,N_1576,N_1930);
nand U2525 (N_2525,N_1544,N_1729);
and U2526 (N_2526,N_1725,N_1997);
nand U2527 (N_2527,N_2089,N_1959);
and U2528 (N_2528,N_1845,N_2244);
nor U2529 (N_2529,N_2153,N_1999);
xor U2530 (N_2530,N_1886,N_1889);
and U2531 (N_2531,N_1559,N_2054);
nor U2532 (N_2532,N_1795,N_1744);
and U2533 (N_2533,N_2198,N_1937);
xor U2534 (N_2534,N_1828,N_1626);
nor U2535 (N_2535,N_2126,N_2057);
or U2536 (N_2536,N_1616,N_2112);
xnor U2537 (N_2537,N_2135,N_2088);
nor U2538 (N_2538,N_1564,N_2056);
or U2539 (N_2539,N_2034,N_1800);
or U2540 (N_2540,N_1768,N_2170);
nor U2541 (N_2541,N_1757,N_1851);
nor U2542 (N_2542,N_1736,N_2136);
nand U2543 (N_2543,N_2218,N_2182);
and U2544 (N_2544,N_2052,N_1741);
and U2545 (N_2545,N_1721,N_1969);
or U2546 (N_2546,N_2011,N_1569);
or U2547 (N_2547,N_1529,N_1810);
nand U2548 (N_2548,N_1556,N_1504);
nor U2549 (N_2549,N_1920,N_1934);
xor U2550 (N_2550,N_1687,N_1595);
or U2551 (N_2551,N_1871,N_1681);
nand U2552 (N_2552,N_1607,N_1500);
nor U2553 (N_2553,N_2147,N_1899);
or U2554 (N_2554,N_1831,N_1503);
and U2555 (N_2555,N_2021,N_2240);
nor U2556 (N_2556,N_2015,N_2203);
and U2557 (N_2557,N_1789,N_2155);
and U2558 (N_2558,N_1677,N_1875);
xnor U2559 (N_2559,N_1797,N_2108);
nor U2560 (N_2560,N_2217,N_1824);
xor U2561 (N_2561,N_2117,N_2080);
xnor U2562 (N_2562,N_1815,N_2020);
and U2563 (N_2563,N_1555,N_2050);
xnor U2564 (N_2564,N_1936,N_1533);
and U2565 (N_2565,N_2078,N_1977);
and U2566 (N_2566,N_1672,N_1706);
nor U2567 (N_2567,N_2079,N_1905);
nor U2568 (N_2568,N_2087,N_1863);
nand U2569 (N_2569,N_1764,N_2245);
or U2570 (N_2570,N_1704,N_1801);
nand U2571 (N_2571,N_1802,N_1719);
xor U2572 (N_2572,N_1553,N_1940);
nand U2573 (N_2573,N_2207,N_1846);
nand U2574 (N_2574,N_1904,N_2154);
and U2575 (N_2575,N_1951,N_1724);
or U2576 (N_2576,N_1985,N_2199);
nand U2577 (N_2577,N_1629,N_1876);
and U2578 (N_2578,N_1840,N_1749);
nor U2579 (N_2579,N_1994,N_1872);
nor U2580 (N_2580,N_2002,N_1835);
nor U2581 (N_2581,N_1833,N_2077);
and U2582 (N_2582,N_1849,N_1650);
and U2583 (N_2583,N_1919,N_1848);
or U2584 (N_2584,N_1868,N_1931);
nor U2585 (N_2585,N_2141,N_1753);
or U2586 (N_2586,N_2179,N_1938);
nor U2587 (N_2587,N_1703,N_1653);
nand U2588 (N_2588,N_1720,N_1879);
xnor U2589 (N_2589,N_1593,N_1523);
nor U2590 (N_2590,N_1613,N_1716);
or U2591 (N_2591,N_2196,N_1784);
and U2592 (N_2592,N_2109,N_1924);
nand U2593 (N_2593,N_1819,N_1787);
and U2594 (N_2594,N_2121,N_2000);
and U2595 (N_2595,N_2243,N_1914);
and U2596 (N_2596,N_1518,N_1910);
and U2597 (N_2597,N_1538,N_1968);
nor U2598 (N_2598,N_1935,N_2124);
and U2599 (N_2599,N_1861,N_1635);
nand U2600 (N_2600,N_2193,N_1918);
nand U2601 (N_2601,N_1758,N_1702);
nand U2602 (N_2602,N_1853,N_1856);
nand U2603 (N_2603,N_1689,N_2110);
or U2604 (N_2604,N_1641,N_2230);
nor U2605 (N_2605,N_1767,N_1552);
nand U2606 (N_2606,N_2066,N_1594);
nand U2607 (N_2607,N_2037,N_1796);
and U2608 (N_2608,N_1697,N_1804);
xor U2609 (N_2609,N_1570,N_1893);
or U2610 (N_2610,N_2051,N_1615);
nor U2611 (N_2611,N_2071,N_1558);
nor U2612 (N_2612,N_1916,N_2130);
nor U2613 (N_2613,N_2200,N_1837);
or U2614 (N_2614,N_1718,N_1639);
and U2615 (N_2615,N_1602,N_2224);
xor U2616 (N_2616,N_2044,N_2171);
or U2617 (N_2617,N_2084,N_1952);
xor U2618 (N_2618,N_2172,N_1779);
nor U2619 (N_2619,N_1711,N_1887);
or U2620 (N_2620,N_2159,N_1998);
or U2621 (N_2621,N_1816,N_2107);
nand U2622 (N_2622,N_2013,N_1574);
nand U2623 (N_2623,N_1928,N_1733);
nand U2624 (N_2624,N_1972,N_1646);
nand U2625 (N_2625,N_2221,N_1791);
and U2626 (N_2626,N_1602,N_1699);
xnor U2627 (N_2627,N_1914,N_1833);
nand U2628 (N_2628,N_1614,N_1914);
nor U2629 (N_2629,N_1667,N_2183);
or U2630 (N_2630,N_2224,N_1533);
or U2631 (N_2631,N_2030,N_2192);
or U2632 (N_2632,N_2177,N_2033);
nand U2633 (N_2633,N_1632,N_1660);
xnor U2634 (N_2634,N_1796,N_2109);
nor U2635 (N_2635,N_1583,N_1692);
or U2636 (N_2636,N_1770,N_1803);
or U2637 (N_2637,N_1789,N_2202);
xnor U2638 (N_2638,N_2108,N_1631);
or U2639 (N_2639,N_1796,N_1967);
or U2640 (N_2640,N_1902,N_2055);
nand U2641 (N_2641,N_1898,N_2023);
nand U2642 (N_2642,N_1556,N_1950);
and U2643 (N_2643,N_1748,N_2097);
nor U2644 (N_2644,N_1979,N_1798);
or U2645 (N_2645,N_1631,N_1752);
nand U2646 (N_2646,N_1630,N_1669);
and U2647 (N_2647,N_1725,N_1944);
nor U2648 (N_2648,N_1841,N_1780);
xnor U2649 (N_2649,N_1776,N_1555);
nor U2650 (N_2650,N_1974,N_1767);
xor U2651 (N_2651,N_2248,N_2051);
nand U2652 (N_2652,N_1957,N_2242);
nor U2653 (N_2653,N_1878,N_1737);
xor U2654 (N_2654,N_2061,N_1737);
nor U2655 (N_2655,N_1834,N_2110);
nand U2656 (N_2656,N_1615,N_1964);
nor U2657 (N_2657,N_1730,N_2145);
nand U2658 (N_2658,N_2015,N_1746);
nor U2659 (N_2659,N_2211,N_2125);
or U2660 (N_2660,N_1689,N_1849);
nand U2661 (N_2661,N_2046,N_1977);
or U2662 (N_2662,N_2239,N_2099);
or U2663 (N_2663,N_1856,N_1980);
and U2664 (N_2664,N_2021,N_1647);
and U2665 (N_2665,N_2006,N_2038);
or U2666 (N_2666,N_1918,N_1594);
xnor U2667 (N_2667,N_2082,N_1885);
nand U2668 (N_2668,N_1542,N_1757);
and U2669 (N_2669,N_1560,N_1830);
or U2670 (N_2670,N_1927,N_2157);
nand U2671 (N_2671,N_1678,N_1544);
and U2672 (N_2672,N_1789,N_1725);
xor U2673 (N_2673,N_1599,N_1674);
nand U2674 (N_2674,N_2138,N_2017);
xor U2675 (N_2675,N_2165,N_2042);
nand U2676 (N_2676,N_2069,N_1520);
and U2677 (N_2677,N_1852,N_1947);
and U2678 (N_2678,N_2008,N_1787);
nor U2679 (N_2679,N_2138,N_2082);
and U2680 (N_2680,N_2036,N_1574);
and U2681 (N_2681,N_1994,N_1738);
xor U2682 (N_2682,N_1771,N_2248);
and U2683 (N_2683,N_1855,N_1654);
nand U2684 (N_2684,N_1632,N_1905);
or U2685 (N_2685,N_2055,N_2084);
nand U2686 (N_2686,N_1659,N_2074);
nand U2687 (N_2687,N_1944,N_1937);
nand U2688 (N_2688,N_2033,N_1628);
nand U2689 (N_2689,N_2036,N_1518);
and U2690 (N_2690,N_2037,N_1909);
nor U2691 (N_2691,N_1660,N_1856);
and U2692 (N_2692,N_2079,N_1816);
nand U2693 (N_2693,N_1775,N_1538);
xor U2694 (N_2694,N_1769,N_2047);
and U2695 (N_2695,N_1647,N_1543);
or U2696 (N_2696,N_1853,N_2060);
nor U2697 (N_2697,N_2161,N_1977);
or U2698 (N_2698,N_1817,N_1772);
nor U2699 (N_2699,N_1542,N_1500);
or U2700 (N_2700,N_1944,N_1989);
and U2701 (N_2701,N_1587,N_1712);
and U2702 (N_2702,N_1654,N_2137);
or U2703 (N_2703,N_1658,N_1580);
nor U2704 (N_2704,N_2069,N_1996);
nand U2705 (N_2705,N_2211,N_2116);
nand U2706 (N_2706,N_2166,N_1797);
nor U2707 (N_2707,N_1742,N_2057);
nand U2708 (N_2708,N_1904,N_1553);
nor U2709 (N_2709,N_1831,N_1708);
nor U2710 (N_2710,N_2178,N_1655);
and U2711 (N_2711,N_2089,N_1998);
xor U2712 (N_2712,N_1567,N_1864);
or U2713 (N_2713,N_1991,N_1630);
and U2714 (N_2714,N_2110,N_1881);
nor U2715 (N_2715,N_1774,N_1739);
nor U2716 (N_2716,N_1992,N_2048);
nor U2717 (N_2717,N_1830,N_1715);
xnor U2718 (N_2718,N_1560,N_2214);
and U2719 (N_2719,N_1895,N_1547);
nor U2720 (N_2720,N_2236,N_1901);
nand U2721 (N_2721,N_1807,N_1915);
or U2722 (N_2722,N_2000,N_2249);
nand U2723 (N_2723,N_1719,N_2077);
nor U2724 (N_2724,N_2101,N_2194);
xnor U2725 (N_2725,N_2069,N_2154);
nand U2726 (N_2726,N_1947,N_2186);
or U2727 (N_2727,N_1742,N_2012);
or U2728 (N_2728,N_1717,N_2238);
nand U2729 (N_2729,N_2175,N_2150);
or U2730 (N_2730,N_1842,N_1892);
nor U2731 (N_2731,N_2179,N_2125);
and U2732 (N_2732,N_1509,N_1968);
nand U2733 (N_2733,N_1527,N_2171);
nor U2734 (N_2734,N_2161,N_1904);
and U2735 (N_2735,N_1843,N_2136);
nand U2736 (N_2736,N_1780,N_1935);
and U2737 (N_2737,N_1548,N_1779);
nand U2738 (N_2738,N_2131,N_1966);
or U2739 (N_2739,N_1560,N_2238);
nand U2740 (N_2740,N_1875,N_1870);
nand U2741 (N_2741,N_1722,N_1737);
and U2742 (N_2742,N_2154,N_2011);
nand U2743 (N_2743,N_1572,N_2143);
nand U2744 (N_2744,N_2008,N_1646);
nand U2745 (N_2745,N_1516,N_1555);
or U2746 (N_2746,N_1884,N_1810);
xor U2747 (N_2747,N_1842,N_1525);
or U2748 (N_2748,N_1530,N_1616);
nor U2749 (N_2749,N_2117,N_1627);
and U2750 (N_2750,N_1870,N_1522);
nand U2751 (N_2751,N_1934,N_1832);
or U2752 (N_2752,N_1601,N_1508);
and U2753 (N_2753,N_1548,N_1571);
or U2754 (N_2754,N_1544,N_1824);
or U2755 (N_2755,N_1923,N_1570);
or U2756 (N_2756,N_1960,N_1758);
and U2757 (N_2757,N_1782,N_1956);
and U2758 (N_2758,N_2090,N_1931);
nor U2759 (N_2759,N_1656,N_2050);
and U2760 (N_2760,N_1594,N_2111);
or U2761 (N_2761,N_1530,N_2015);
or U2762 (N_2762,N_1516,N_1655);
xor U2763 (N_2763,N_1847,N_1573);
and U2764 (N_2764,N_1554,N_1771);
or U2765 (N_2765,N_1968,N_1522);
nand U2766 (N_2766,N_2094,N_1716);
or U2767 (N_2767,N_1692,N_1590);
and U2768 (N_2768,N_2073,N_1913);
and U2769 (N_2769,N_1644,N_2217);
xor U2770 (N_2770,N_2182,N_2227);
and U2771 (N_2771,N_1667,N_1884);
nand U2772 (N_2772,N_1821,N_1581);
or U2773 (N_2773,N_1874,N_1615);
xnor U2774 (N_2774,N_2177,N_1771);
nand U2775 (N_2775,N_1583,N_2149);
nand U2776 (N_2776,N_1520,N_1783);
xnor U2777 (N_2777,N_2022,N_1768);
xnor U2778 (N_2778,N_1853,N_1923);
and U2779 (N_2779,N_1595,N_1903);
nand U2780 (N_2780,N_1658,N_1553);
nor U2781 (N_2781,N_1580,N_1572);
and U2782 (N_2782,N_1920,N_2150);
xnor U2783 (N_2783,N_1596,N_2014);
and U2784 (N_2784,N_2140,N_2069);
nand U2785 (N_2785,N_2084,N_2123);
nor U2786 (N_2786,N_1575,N_1557);
xnor U2787 (N_2787,N_1514,N_2065);
nand U2788 (N_2788,N_1579,N_2120);
nand U2789 (N_2789,N_1655,N_1665);
nor U2790 (N_2790,N_1855,N_1587);
and U2791 (N_2791,N_1973,N_2234);
or U2792 (N_2792,N_1953,N_1940);
nor U2793 (N_2793,N_1907,N_1837);
nor U2794 (N_2794,N_2077,N_1968);
nor U2795 (N_2795,N_1640,N_1879);
or U2796 (N_2796,N_1530,N_1698);
nor U2797 (N_2797,N_2129,N_1925);
or U2798 (N_2798,N_1532,N_2237);
nor U2799 (N_2799,N_1792,N_2123);
and U2800 (N_2800,N_1932,N_1950);
nor U2801 (N_2801,N_1985,N_2164);
nor U2802 (N_2802,N_1903,N_2051);
nor U2803 (N_2803,N_1618,N_1872);
nor U2804 (N_2804,N_1676,N_2122);
or U2805 (N_2805,N_1973,N_1689);
nor U2806 (N_2806,N_1851,N_2152);
or U2807 (N_2807,N_1838,N_1822);
or U2808 (N_2808,N_1598,N_1622);
nor U2809 (N_2809,N_1830,N_1653);
and U2810 (N_2810,N_2225,N_1731);
or U2811 (N_2811,N_2001,N_2152);
and U2812 (N_2812,N_1917,N_1528);
nor U2813 (N_2813,N_2015,N_1632);
or U2814 (N_2814,N_2010,N_2070);
xnor U2815 (N_2815,N_2046,N_2066);
xor U2816 (N_2816,N_1564,N_1781);
and U2817 (N_2817,N_2141,N_2149);
and U2818 (N_2818,N_2012,N_1610);
nor U2819 (N_2819,N_1780,N_2004);
nor U2820 (N_2820,N_2185,N_1956);
nor U2821 (N_2821,N_1685,N_1707);
or U2822 (N_2822,N_1817,N_2028);
and U2823 (N_2823,N_1733,N_1924);
and U2824 (N_2824,N_2150,N_1854);
xor U2825 (N_2825,N_2210,N_2182);
nand U2826 (N_2826,N_2039,N_1932);
nand U2827 (N_2827,N_1734,N_1929);
nand U2828 (N_2828,N_1736,N_2006);
or U2829 (N_2829,N_1578,N_2218);
or U2830 (N_2830,N_2112,N_1593);
and U2831 (N_2831,N_1945,N_1913);
nand U2832 (N_2832,N_2035,N_1883);
nand U2833 (N_2833,N_1867,N_2049);
and U2834 (N_2834,N_1535,N_1812);
nand U2835 (N_2835,N_1715,N_2043);
and U2836 (N_2836,N_1905,N_1527);
nor U2837 (N_2837,N_1578,N_1656);
or U2838 (N_2838,N_1762,N_1557);
and U2839 (N_2839,N_1794,N_1869);
or U2840 (N_2840,N_2022,N_1639);
and U2841 (N_2841,N_2210,N_1966);
xnor U2842 (N_2842,N_1916,N_1807);
nand U2843 (N_2843,N_1926,N_1927);
nor U2844 (N_2844,N_1978,N_1965);
nor U2845 (N_2845,N_1691,N_2148);
nor U2846 (N_2846,N_1534,N_1735);
nand U2847 (N_2847,N_1671,N_2223);
or U2848 (N_2848,N_2126,N_1608);
nand U2849 (N_2849,N_1983,N_2043);
and U2850 (N_2850,N_2146,N_2128);
nand U2851 (N_2851,N_2032,N_2217);
or U2852 (N_2852,N_1993,N_2045);
or U2853 (N_2853,N_1951,N_1543);
and U2854 (N_2854,N_1963,N_1987);
nor U2855 (N_2855,N_2227,N_1912);
nand U2856 (N_2856,N_1895,N_1726);
nand U2857 (N_2857,N_1970,N_1542);
nor U2858 (N_2858,N_1813,N_2072);
and U2859 (N_2859,N_1794,N_1716);
nor U2860 (N_2860,N_1727,N_1984);
or U2861 (N_2861,N_1736,N_1927);
xor U2862 (N_2862,N_2178,N_2018);
xnor U2863 (N_2863,N_2207,N_1659);
and U2864 (N_2864,N_2027,N_2223);
and U2865 (N_2865,N_1879,N_2107);
and U2866 (N_2866,N_2204,N_1930);
nor U2867 (N_2867,N_1537,N_2147);
nor U2868 (N_2868,N_1701,N_1864);
or U2869 (N_2869,N_1589,N_1522);
nor U2870 (N_2870,N_1794,N_1642);
and U2871 (N_2871,N_2002,N_1860);
and U2872 (N_2872,N_1952,N_1614);
nor U2873 (N_2873,N_2167,N_1621);
nand U2874 (N_2874,N_1834,N_1517);
or U2875 (N_2875,N_2037,N_1584);
and U2876 (N_2876,N_2146,N_1574);
nor U2877 (N_2877,N_1500,N_2032);
nand U2878 (N_2878,N_2245,N_1850);
nand U2879 (N_2879,N_2008,N_1556);
or U2880 (N_2880,N_1711,N_2017);
nor U2881 (N_2881,N_2061,N_1818);
nand U2882 (N_2882,N_2106,N_1993);
xnor U2883 (N_2883,N_2000,N_1908);
and U2884 (N_2884,N_1779,N_2023);
and U2885 (N_2885,N_1668,N_2021);
nand U2886 (N_2886,N_1619,N_1624);
or U2887 (N_2887,N_1905,N_1859);
or U2888 (N_2888,N_2081,N_1534);
nand U2889 (N_2889,N_1633,N_1748);
nor U2890 (N_2890,N_2093,N_2039);
or U2891 (N_2891,N_1630,N_1830);
or U2892 (N_2892,N_2161,N_1570);
and U2893 (N_2893,N_2238,N_1651);
nor U2894 (N_2894,N_1820,N_2180);
and U2895 (N_2895,N_2060,N_2006);
and U2896 (N_2896,N_2246,N_1943);
nand U2897 (N_2897,N_1806,N_1505);
nand U2898 (N_2898,N_1673,N_2013);
nand U2899 (N_2899,N_2032,N_1523);
and U2900 (N_2900,N_1949,N_1631);
nand U2901 (N_2901,N_1831,N_1561);
nor U2902 (N_2902,N_2016,N_2027);
nand U2903 (N_2903,N_1826,N_2086);
xor U2904 (N_2904,N_1793,N_1831);
or U2905 (N_2905,N_2101,N_2166);
nor U2906 (N_2906,N_1613,N_1532);
nand U2907 (N_2907,N_2036,N_1886);
and U2908 (N_2908,N_1944,N_2025);
and U2909 (N_2909,N_1714,N_1627);
nor U2910 (N_2910,N_1914,N_1519);
nor U2911 (N_2911,N_2067,N_1503);
xor U2912 (N_2912,N_2119,N_1981);
nor U2913 (N_2913,N_1597,N_1651);
nor U2914 (N_2914,N_2003,N_1794);
nand U2915 (N_2915,N_2085,N_2116);
nand U2916 (N_2916,N_1696,N_1612);
or U2917 (N_2917,N_1808,N_1767);
nand U2918 (N_2918,N_2180,N_1857);
and U2919 (N_2919,N_1963,N_2087);
or U2920 (N_2920,N_2072,N_2080);
nand U2921 (N_2921,N_1835,N_1570);
and U2922 (N_2922,N_1871,N_2027);
and U2923 (N_2923,N_1787,N_1788);
nor U2924 (N_2924,N_2097,N_1706);
nor U2925 (N_2925,N_2002,N_1992);
nor U2926 (N_2926,N_2170,N_2214);
or U2927 (N_2927,N_1604,N_2222);
nand U2928 (N_2928,N_2216,N_1827);
or U2929 (N_2929,N_1831,N_1917);
and U2930 (N_2930,N_1895,N_1676);
xor U2931 (N_2931,N_1761,N_1984);
xnor U2932 (N_2932,N_2041,N_1796);
nor U2933 (N_2933,N_2015,N_1806);
nand U2934 (N_2934,N_1814,N_2247);
nand U2935 (N_2935,N_1686,N_1561);
or U2936 (N_2936,N_2155,N_2135);
xor U2937 (N_2937,N_1901,N_1831);
nor U2938 (N_2938,N_1949,N_2232);
xor U2939 (N_2939,N_1900,N_1998);
nand U2940 (N_2940,N_2231,N_1637);
or U2941 (N_2941,N_1787,N_1693);
or U2942 (N_2942,N_1780,N_1983);
nor U2943 (N_2943,N_1895,N_2241);
or U2944 (N_2944,N_1566,N_2230);
or U2945 (N_2945,N_1981,N_1527);
nor U2946 (N_2946,N_1814,N_1776);
or U2947 (N_2947,N_2195,N_2245);
or U2948 (N_2948,N_1913,N_1766);
nand U2949 (N_2949,N_1761,N_2106);
nor U2950 (N_2950,N_2249,N_1530);
nand U2951 (N_2951,N_2009,N_1828);
nor U2952 (N_2952,N_1951,N_2073);
or U2953 (N_2953,N_2116,N_1910);
nor U2954 (N_2954,N_2161,N_1531);
nor U2955 (N_2955,N_1768,N_2087);
and U2956 (N_2956,N_1787,N_1998);
and U2957 (N_2957,N_1508,N_1877);
or U2958 (N_2958,N_2094,N_2001);
and U2959 (N_2959,N_2022,N_1556);
nand U2960 (N_2960,N_2179,N_1639);
or U2961 (N_2961,N_1750,N_1544);
nor U2962 (N_2962,N_2203,N_1950);
nor U2963 (N_2963,N_1646,N_1779);
nand U2964 (N_2964,N_1508,N_2232);
nor U2965 (N_2965,N_1947,N_2029);
nor U2966 (N_2966,N_2056,N_1577);
or U2967 (N_2967,N_1672,N_1659);
nor U2968 (N_2968,N_1977,N_2108);
and U2969 (N_2969,N_2158,N_2032);
or U2970 (N_2970,N_1678,N_2046);
and U2971 (N_2971,N_2234,N_2013);
nor U2972 (N_2972,N_1839,N_2017);
nor U2973 (N_2973,N_1543,N_1926);
nand U2974 (N_2974,N_1776,N_1530);
or U2975 (N_2975,N_2143,N_2185);
nor U2976 (N_2976,N_1782,N_2026);
and U2977 (N_2977,N_1813,N_1777);
nand U2978 (N_2978,N_1534,N_2011);
nor U2979 (N_2979,N_1690,N_1503);
or U2980 (N_2980,N_1887,N_2208);
nand U2981 (N_2981,N_2033,N_2105);
nor U2982 (N_2982,N_2089,N_1566);
or U2983 (N_2983,N_1968,N_1581);
or U2984 (N_2984,N_1595,N_1927);
and U2985 (N_2985,N_1666,N_2157);
and U2986 (N_2986,N_1613,N_1770);
or U2987 (N_2987,N_1910,N_1515);
nor U2988 (N_2988,N_2224,N_1613);
nand U2989 (N_2989,N_1554,N_1880);
nor U2990 (N_2990,N_2136,N_2041);
nor U2991 (N_2991,N_2105,N_2121);
nor U2992 (N_2992,N_1754,N_1921);
or U2993 (N_2993,N_2176,N_2094);
and U2994 (N_2994,N_1998,N_1692);
and U2995 (N_2995,N_1786,N_1593);
nor U2996 (N_2996,N_1700,N_2093);
xor U2997 (N_2997,N_2239,N_2104);
and U2998 (N_2998,N_2232,N_1908);
and U2999 (N_2999,N_1758,N_2182);
nand UO_0 (O_0,N_2770,N_2373);
or UO_1 (O_1,N_2355,N_2449);
and UO_2 (O_2,N_2756,N_2827);
nor UO_3 (O_3,N_2347,N_2587);
or UO_4 (O_4,N_2922,N_2268);
nand UO_5 (O_5,N_2512,N_2309);
nand UO_6 (O_6,N_2434,N_2916);
nand UO_7 (O_7,N_2340,N_2873);
nand UO_8 (O_8,N_2724,N_2799);
or UO_9 (O_9,N_2938,N_2531);
nand UO_10 (O_10,N_2689,N_2384);
xor UO_11 (O_11,N_2420,N_2297);
nand UO_12 (O_12,N_2358,N_2726);
or UO_13 (O_13,N_2598,N_2332);
or UO_14 (O_14,N_2655,N_2704);
and UO_15 (O_15,N_2363,N_2401);
and UO_16 (O_16,N_2290,N_2845);
and UO_17 (O_17,N_2254,N_2965);
nand UO_18 (O_18,N_2354,N_2285);
and UO_19 (O_19,N_2788,N_2472);
nor UO_20 (O_20,N_2262,N_2331);
nor UO_21 (O_21,N_2550,N_2630);
nand UO_22 (O_22,N_2283,N_2780);
or UO_23 (O_23,N_2641,N_2897);
nand UO_24 (O_24,N_2623,N_2576);
nand UO_25 (O_25,N_2733,N_2624);
nand UO_26 (O_26,N_2737,N_2446);
and UO_27 (O_27,N_2293,N_2350);
nor UO_28 (O_28,N_2761,N_2785);
nand UO_29 (O_29,N_2554,N_2977);
and UO_30 (O_30,N_2452,N_2742);
nand UO_31 (O_31,N_2383,N_2578);
and UO_32 (O_32,N_2498,N_2457);
nor UO_33 (O_33,N_2648,N_2351);
nand UO_34 (O_34,N_2691,N_2545);
xnor UO_35 (O_35,N_2859,N_2880);
xor UO_36 (O_36,N_2376,N_2805);
nand UO_37 (O_37,N_2701,N_2806);
and UO_38 (O_38,N_2687,N_2719);
nand UO_39 (O_39,N_2601,N_2964);
nand UO_40 (O_40,N_2517,N_2345);
nor UO_41 (O_41,N_2560,N_2636);
or UO_42 (O_42,N_2522,N_2365);
xnor UO_43 (O_43,N_2708,N_2782);
and UO_44 (O_44,N_2839,N_2769);
and UO_45 (O_45,N_2444,N_2926);
or UO_46 (O_46,N_2323,N_2903);
or UO_47 (O_47,N_2468,N_2454);
nand UO_48 (O_48,N_2798,N_2665);
and UO_49 (O_49,N_2296,N_2666);
nand UO_50 (O_50,N_2929,N_2651);
and UO_51 (O_51,N_2612,N_2842);
nand UO_52 (O_52,N_2727,N_2721);
nor UO_53 (O_53,N_2802,N_2277);
and UO_54 (O_54,N_2960,N_2824);
or UO_55 (O_55,N_2917,N_2319);
nor UO_56 (O_56,N_2690,N_2458);
nand UO_57 (O_57,N_2479,N_2962);
nor UO_58 (O_58,N_2432,N_2492);
and UO_59 (O_59,N_2489,N_2483);
nand UO_60 (O_60,N_2341,N_2318);
nand UO_61 (O_61,N_2966,N_2588);
nand UO_62 (O_62,N_2884,N_2694);
nor UO_63 (O_63,N_2301,N_2586);
and UO_64 (O_64,N_2344,N_2754);
nor UO_65 (O_65,N_2914,N_2900);
nand UO_66 (O_66,N_2652,N_2907);
and UO_67 (O_67,N_2543,N_2764);
nor UO_68 (O_68,N_2306,N_2534);
or UO_69 (O_69,N_2375,N_2382);
nor UO_70 (O_70,N_2553,N_2577);
nand UO_71 (O_71,N_2295,N_2933);
nor UO_72 (O_72,N_2431,N_2276);
or UO_73 (O_73,N_2503,N_2581);
nor UO_74 (O_74,N_2437,N_2524);
or UO_75 (O_75,N_2870,N_2759);
nand UO_76 (O_76,N_2608,N_2357);
nor UO_77 (O_77,N_2281,N_2564);
nand UO_78 (O_78,N_2846,N_2925);
or UO_79 (O_79,N_2312,N_2656);
or UO_80 (O_80,N_2414,N_2450);
nor UO_81 (O_81,N_2872,N_2519);
nand UO_82 (O_82,N_2279,N_2356);
or UO_83 (O_83,N_2867,N_2711);
nand UO_84 (O_84,N_2419,N_2749);
xor UO_85 (O_85,N_2703,N_2530);
nor UO_86 (O_86,N_2583,N_2407);
nand UO_87 (O_87,N_2958,N_2506);
nor UO_88 (O_88,N_2265,N_2795);
nand UO_89 (O_89,N_2705,N_2835);
or UO_90 (O_90,N_2546,N_2850);
nand UO_91 (O_91,N_2547,N_2322);
or UO_92 (O_92,N_2395,N_2275);
nor UO_93 (O_93,N_2307,N_2783);
nor UO_94 (O_94,N_2532,N_2616);
and UO_95 (O_95,N_2607,N_2669);
nand UO_96 (O_96,N_2954,N_2399);
nor UO_97 (O_97,N_2728,N_2902);
and UO_98 (O_98,N_2571,N_2700);
and UO_99 (O_99,N_2280,N_2858);
or UO_100 (O_100,N_2619,N_2699);
nor UO_101 (O_101,N_2948,N_2590);
or UO_102 (O_102,N_2896,N_2470);
xor UO_103 (O_103,N_2515,N_2342);
nand UO_104 (O_104,N_2818,N_2939);
and UO_105 (O_105,N_2533,N_2812);
nand UO_106 (O_106,N_2814,N_2360);
and UO_107 (O_107,N_2570,N_2716);
and UO_108 (O_108,N_2766,N_2843);
nand UO_109 (O_109,N_2398,N_2313);
nand UO_110 (O_110,N_2520,N_2288);
and UO_111 (O_111,N_2676,N_2603);
and UO_112 (O_112,N_2300,N_2287);
xor UO_113 (O_113,N_2421,N_2946);
nand UO_114 (O_114,N_2992,N_2540);
nand UO_115 (O_115,N_2516,N_2730);
or UO_116 (O_116,N_2881,N_2349);
nor UO_117 (O_117,N_2316,N_2695);
and UO_118 (O_118,N_2252,N_2626);
nand UO_119 (O_119,N_2679,N_2574);
or UO_120 (O_120,N_2717,N_2480);
nor UO_121 (O_121,N_2745,N_2777);
or UO_122 (O_122,N_2459,N_2836);
nor UO_123 (O_123,N_2575,N_2681);
nor UO_124 (O_124,N_2311,N_2928);
and UO_125 (O_125,N_2696,N_2819);
and UO_126 (O_126,N_2830,N_2505);
nor UO_127 (O_127,N_2847,N_2353);
and UO_128 (O_128,N_2582,N_2477);
and UO_129 (O_129,N_2453,N_2853);
nor UO_130 (O_130,N_2658,N_2561);
and UO_131 (O_131,N_2969,N_2289);
and UO_132 (O_132,N_2329,N_2986);
and UO_133 (O_133,N_2707,N_2611);
nand UO_134 (O_134,N_2396,N_2250);
xnor UO_135 (O_135,N_2370,N_2927);
and UO_136 (O_136,N_2408,N_2308);
and UO_137 (O_137,N_2486,N_2474);
nor UO_138 (O_138,N_2475,N_2998);
nor UO_139 (O_139,N_2768,N_2871);
or UO_140 (O_140,N_2748,N_2438);
and UO_141 (O_141,N_2990,N_2677);
or UO_142 (O_142,N_2565,N_2501);
or UO_143 (O_143,N_2469,N_2654);
nor UO_144 (O_144,N_2755,N_2481);
or UO_145 (O_145,N_2993,N_2807);
nand UO_146 (O_146,N_2367,N_2826);
or UO_147 (O_147,N_2649,N_2364);
or UO_148 (O_148,N_2580,N_2878);
nor UO_149 (O_149,N_2659,N_2298);
and UO_150 (O_150,N_2589,N_2465);
nor UO_151 (O_151,N_2251,N_2832);
nand UO_152 (O_152,N_2974,N_2326);
nor UO_153 (O_153,N_2821,N_2911);
or UO_154 (O_154,N_2678,N_2609);
nor UO_155 (O_155,N_2892,N_2646);
nand UO_156 (O_156,N_2815,N_2513);
and UO_157 (O_157,N_2291,N_2371);
xor UO_158 (O_158,N_2889,N_2810);
or UO_159 (O_159,N_2856,N_2792);
nor UO_160 (O_160,N_2418,N_2661);
nand UO_161 (O_161,N_2976,N_2941);
nor UO_162 (O_162,N_2668,N_2735);
or UO_163 (O_163,N_2910,N_2321);
nor UO_164 (O_164,N_2831,N_2467);
and UO_165 (O_165,N_2504,N_2294);
and UO_166 (O_166,N_2763,N_2264);
nor UO_167 (O_167,N_2725,N_2667);
and UO_168 (O_168,N_2614,N_2885);
and UO_169 (O_169,N_2428,N_2854);
and UO_170 (O_170,N_2338,N_2862);
and UO_171 (O_171,N_2409,N_2959);
or UO_172 (O_172,N_2278,N_2563);
or UO_173 (O_173,N_2698,N_2688);
nor UO_174 (O_174,N_2888,N_2915);
nand UO_175 (O_175,N_2899,N_2482);
nand UO_176 (O_176,N_2841,N_2267);
nand UO_177 (O_177,N_2377,N_2372);
nand UO_178 (O_178,N_2919,N_2299);
xnor UO_179 (O_179,N_2476,N_2790);
and UO_180 (O_180,N_2935,N_2573);
nor UO_181 (O_181,N_2877,N_2493);
nor UO_182 (O_182,N_2400,N_2988);
and UO_183 (O_183,N_2820,N_2529);
and UO_184 (O_184,N_2594,N_2855);
and UO_185 (O_185,N_2424,N_2789);
nor UO_186 (O_186,N_2392,N_2706);
and UO_187 (O_187,N_2741,N_2991);
nand UO_188 (O_188,N_2572,N_2876);
or UO_189 (O_189,N_2374,N_2593);
and UO_190 (O_190,N_2848,N_2809);
or UO_191 (O_191,N_2255,N_2585);
and UO_192 (O_192,N_2874,N_2447);
nand UO_193 (O_193,N_2464,N_2989);
xnor UO_194 (O_194,N_2963,N_2422);
or UO_195 (O_195,N_2496,N_2924);
nand UO_196 (O_196,N_2639,N_2260);
or UO_197 (O_197,N_2999,N_2787);
nand UO_198 (O_198,N_2542,N_2595);
nor UO_199 (O_199,N_2975,N_2932);
and UO_200 (O_200,N_2765,N_2747);
or UO_201 (O_201,N_2647,N_2822);
nand UO_202 (O_202,N_2793,N_2462);
and UO_203 (O_203,N_2697,N_2272);
or UO_204 (O_204,N_2936,N_2514);
nand UO_205 (O_205,N_2898,N_2718);
or UO_206 (O_206,N_2253,N_2642);
nand UO_207 (O_207,N_2567,N_2320);
and UO_208 (O_208,N_2863,N_2430);
xnor UO_209 (O_209,N_2304,N_2934);
nand UO_210 (O_210,N_2348,N_2388);
nor UO_211 (O_211,N_2713,N_2702);
or UO_212 (O_212,N_2602,N_2817);
nor UO_213 (O_213,N_2261,N_2852);
nor UO_214 (O_214,N_2971,N_2495);
and UO_215 (O_215,N_2500,N_2473);
and UO_216 (O_216,N_2983,N_2368);
and UO_217 (O_217,N_2961,N_2346);
nor UO_218 (O_218,N_2794,N_2995);
nor UO_219 (O_219,N_2629,N_2369);
nor UO_220 (O_220,N_2536,N_2606);
nor UO_221 (O_221,N_2439,N_2823);
or UO_222 (O_222,N_2552,N_2951);
nand UO_223 (O_223,N_2406,N_2451);
nor UO_224 (O_224,N_2786,N_2596);
xnor UO_225 (O_225,N_2597,N_2685);
or UO_226 (O_226,N_2394,N_2869);
and UO_227 (O_227,N_2569,N_2343);
nand UO_228 (O_228,N_2901,N_2861);
nand UO_229 (O_229,N_2610,N_2271);
and UO_230 (O_230,N_2851,N_2840);
xor UO_231 (O_231,N_2672,N_2633);
nor UO_232 (O_232,N_2539,N_2904);
xnor UO_233 (O_233,N_2987,N_2729);
and UO_234 (O_234,N_2441,N_2397);
or UO_235 (O_235,N_2838,N_2837);
nor UO_236 (O_236,N_2947,N_2890);
or UO_237 (O_237,N_2617,N_2772);
nand UO_238 (O_238,N_2541,N_2274);
or UO_239 (O_239,N_2709,N_2337);
nor UO_240 (O_240,N_2303,N_2968);
nand UO_241 (O_241,N_2499,N_2778);
nand UO_242 (O_242,N_2671,N_2762);
or UO_243 (O_243,N_2429,N_2945);
and UO_244 (O_244,N_2555,N_2548);
and UO_245 (O_245,N_2662,N_2411);
xor UO_246 (O_246,N_2967,N_2317);
and UO_247 (O_247,N_2996,N_2637);
and UO_248 (O_248,N_2605,N_2740);
nand UO_249 (O_249,N_2269,N_2791);
xnor UO_250 (O_250,N_2886,N_2361);
and UO_251 (O_251,N_2640,N_2891);
and UO_252 (O_252,N_2895,N_2875);
and UO_253 (O_253,N_2774,N_2883);
and UO_254 (O_254,N_2664,N_2921);
xor UO_255 (O_255,N_2402,N_2849);
and UO_256 (O_256,N_2628,N_2868);
nor UO_257 (O_257,N_2620,N_2525);
and UO_258 (O_258,N_2722,N_2282);
nor UO_259 (O_259,N_2270,N_2305);
nor UO_260 (O_260,N_2510,N_2913);
or UO_261 (O_261,N_2315,N_2436);
nor UO_262 (O_262,N_2714,N_2887);
nor UO_263 (O_263,N_2390,N_2710);
nand UO_264 (O_264,N_2621,N_2256);
and UO_265 (O_265,N_2334,N_2956);
or UO_266 (O_266,N_2751,N_2442);
nor UO_267 (O_267,N_2404,N_2273);
nand UO_268 (O_268,N_2405,N_2739);
or UO_269 (O_269,N_2937,N_2314);
nand UO_270 (O_270,N_2448,N_2757);
nand UO_271 (O_271,N_2663,N_2604);
or UO_272 (O_272,N_2744,N_2385);
or UO_273 (O_273,N_2923,N_2638);
nor UO_274 (O_274,N_2461,N_2487);
nor UO_275 (O_275,N_2389,N_2403);
and UO_276 (O_276,N_2352,N_2692);
nor UO_277 (O_277,N_2627,N_2644);
xor UO_278 (O_278,N_2440,N_2425);
or UO_279 (O_279,N_2734,N_2912);
nor UO_280 (O_280,N_2746,N_2776);
or UO_281 (O_281,N_2391,N_2781);
and UO_282 (O_282,N_2767,N_2328);
nor UO_283 (O_283,N_2981,N_2864);
nor UO_284 (O_284,N_2731,N_2518);
and UO_285 (O_285,N_2286,N_2797);
or UO_286 (O_286,N_2618,N_2335);
or UO_287 (O_287,N_2393,N_2615);
nor UO_288 (O_288,N_2538,N_2645);
or UO_289 (O_289,N_2359,N_2686);
or UO_290 (O_290,N_2433,N_2860);
nand UO_291 (O_291,N_2804,N_2456);
nand UO_292 (O_292,N_2634,N_2994);
xnor UO_293 (O_293,N_2879,N_2632);
and UO_294 (O_294,N_2327,N_2257);
or UO_295 (O_295,N_2978,N_2779);
or UO_296 (O_296,N_2362,N_2339);
or UO_297 (O_297,N_2775,N_2423);
nor UO_298 (O_298,N_2549,N_2882);
xor UO_299 (O_299,N_2680,N_2502);
or UO_300 (O_300,N_2412,N_2909);
and UO_301 (O_301,N_2684,N_2292);
or UO_302 (O_302,N_2950,N_2381);
nand UO_303 (O_303,N_2497,N_2738);
nor UO_304 (O_304,N_2490,N_2491);
and UO_305 (O_305,N_2478,N_2427);
nor UO_306 (O_306,N_2920,N_2803);
and UO_307 (O_307,N_2263,N_2972);
nand UO_308 (O_308,N_2484,N_2622);
nand UO_309 (O_309,N_2387,N_2918);
or UO_310 (O_310,N_2712,N_2258);
or UO_311 (O_311,N_2535,N_2984);
nand UO_312 (O_312,N_2386,N_2463);
nand UO_313 (O_313,N_2310,N_2715);
or UO_314 (O_314,N_2908,N_2723);
or UO_315 (O_315,N_2732,N_2566);
or UO_316 (O_316,N_2758,N_2736);
or UO_317 (O_317,N_2635,N_2526);
and UO_318 (O_318,N_2366,N_2544);
and UO_319 (O_319,N_2944,N_2556);
nor UO_320 (O_320,N_2557,N_2771);
and UO_321 (O_321,N_2930,N_2866);
nor UO_322 (O_322,N_2865,N_2488);
and UO_323 (O_323,N_2952,N_2940);
nor UO_324 (O_324,N_2833,N_2650);
nand UO_325 (O_325,N_2631,N_2284);
or UO_326 (O_326,N_2537,N_2825);
nand UO_327 (O_327,N_2509,N_2693);
nor UO_328 (O_328,N_2455,N_2333);
and UO_329 (O_329,N_2527,N_2813);
nand UO_330 (O_330,N_2266,N_2562);
and UO_331 (O_331,N_2753,N_2528);
or UO_332 (O_332,N_2325,N_2808);
nor UO_333 (O_333,N_2949,N_2931);
nor UO_334 (O_334,N_2955,N_2894);
nand UO_335 (O_335,N_2905,N_2568);
nor UO_336 (O_336,N_2796,N_2893);
and UO_337 (O_337,N_2600,N_2720);
nor UO_338 (O_338,N_2471,N_2643);
and UO_339 (O_339,N_2816,N_2957);
and UO_340 (O_340,N_2683,N_2625);
nor UO_341 (O_341,N_2445,N_2670);
xor UO_342 (O_342,N_2985,N_2380);
and UO_343 (O_343,N_2800,N_2980);
and UO_344 (O_344,N_2416,N_2844);
or UO_345 (O_345,N_2584,N_2752);
xor UO_346 (O_346,N_2521,N_2435);
nand UO_347 (O_347,N_2330,N_2551);
nor UO_348 (O_348,N_2970,N_2523);
or UO_349 (O_349,N_2953,N_2801);
or UO_350 (O_350,N_2507,N_2857);
nand UO_351 (O_351,N_2653,N_2415);
and UO_352 (O_352,N_2829,N_2811);
nor UO_353 (O_353,N_2613,N_2973);
or UO_354 (O_354,N_2784,N_2559);
xnor UO_355 (O_355,N_2675,N_2773);
and UO_356 (O_356,N_2302,N_2466);
and UO_357 (O_357,N_2592,N_2426);
and UO_358 (O_358,N_2336,N_2591);
and UO_359 (O_359,N_2379,N_2324);
nor UO_360 (O_360,N_2979,N_2760);
or UO_361 (O_361,N_2485,N_2942);
and UO_362 (O_362,N_2410,N_2943);
and UO_363 (O_363,N_2579,N_2511);
nand UO_364 (O_364,N_2259,N_2743);
or UO_365 (O_365,N_2828,N_2494);
and UO_366 (O_366,N_2508,N_2460);
or UO_367 (O_367,N_2997,N_2443);
nor UO_368 (O_368,N_2413,N_2657);
nor UO_369 (O_369,N_2674,N_2660);
nor UO_370 (O_370,N_2906,N_2417);
xnor UO_371 (O_371,N_2834,N_2982);
nor UO_372 (O_372,N_2599,N_2682);
and UO_373 (O_373,N_2750,N_2378);
nand UO_374 (O_374,N_2558,N_2673);
or UO_375 (O_375,N_2601,N_2698);
nor UO_376 (O_376,N_2628,N_2462);
and UO_377 (O_377,N_2725,N_2427);
and UO_378 (O_378,N_2809,N_2860);
nor UO_379 (O_379,N_2957,N_2974);
and UO_380 (O_380,N_2660,N_2256);
and UO_381 (O_381,N_2752,N_2516);
or UO_382 (O_382,N_2626,N_2704);
or UO_383 (O_383,N_2915,N_2733);
or UO_384 (O_384,N_2796,N_2355);
or UO_385 (O_385,N_2316,N_2303);
and UO_386 (O_386,N_2440,N_2280);
or UO_387 (O_387,N_2969,N_2367);
or UO_388 (O_388,N_2766,N_2810);
or UO_389 (O_389,N_2681,N_2958);
nor UO_390 (O_390,N_2678,N_2759);
and UO_391 (O_391,N_2470,N_2860);
or UO_392 (O_392,N_2695,N_2927);
or UO_393 (O_393,N_2877,N_2937);
nor UO_394 (O_394,N_2668,N_2304);
xor UO_395 (O_395,N_2719,N_2524);
and UO_396 (O_396,N_2597,N_2338);
nand UO_397 (O_397,N_2301,N_2523);
or UO_398 (O_398,N_2368,N_2875);
nor UO_399 (O_399,N_2355,N_2985);
xnor UO_400 (O_400,N_2314,N_2576);
and UO_401 (O_401,N_2356,N_2801);
nor UO_402 (O_402,N_2449,N_2740);
and UO_403 (O_403,N_2694,N_2475);
nand UO_404 (O_404,N_2680,N_2415);
nor UO_405 (O_405,N_2883,N_2791);
and UO_406 (O_406,N_2955,N_2370);
xnor UO_407 (O_407,N_2751,N_2913);
nand UO_408 (O_408,N_2652,N_2589);
nor UO_409 (O_409,N_2512,N_2648);
nand UO_410 (O_410,N_2589,N_2628);
nand UO_411 (O_411,N_2773,N_2613);
and UO_412 (O_412,N_2348,N_2964);
nor UO_413 (O_413,N_2373,N_2922);
nand UO_414 (O_414,N_2796,N_2551);
or UO_415 (O_415,N_2756,N_2269);
or UO_416 (O_416,N_2427,N_2967);
or UO_417 (O_417,N_2383,N_2488);
and UO_418 (O_418,N_2461,N_2628);
nand UO_419 (O_419,N_2803,N_2906);
or UO_420 (O_420,N_2930,N_2522);
or UO_421 (O_421,N_2767,N_2594);
nand UO_422 (O_422,N_2892,N_2457);
nand UO_423 (O_423,N_2374,N_2461);
nand UO_424 (O_424,N_2935,N_2355);
nor UO_425 (O_425,N_2763,N_2577);
or UO_426 (O_426,N_2723,N_2984);
xnor UO_427 (O_427,N_2777,N_2563);
nand UO_428 (O_428,N_2695,N_2596);
nand UO_429 (O_429,N_2839,N_2802);
or UO_430 (O_430,N_2713,N_2476);
and UO_431 (O_431,N_2391,N_2834);
nand UO_432 (O_432,N_2836,N_2806);
or UO_433 (O_433,N_2966,N_2937);
nand UO_434 (O_434,N_2368,N_2613);
or UO_435 (O_435,N_2866,N_2818);
or UO_436 (O_436,N_2327,N_2821);
nor UO_437 (O_437,N_2669,N_2451);
nand UO_438 (O_438,N_2365,N_2369);
xnor UO_439 (O_439,N_2250,N_2909);
xnor UO_440 (O_440,N_2276,N_2628);
or UO_441 (O_441,N_2742,N_2293);
nand UO_442 (O_442,N_2262,N_2487);
xnor UO_443 (O_443,N_2433,N_2970);
or UO_444 (O_444,N_2892,N_2342);
nand UO_445 (O_445,N_2327,N_2381);
or UO_446 (O_446,N_2383,N_2708);
nor UO_447 (O_447,N_2834,N_2557);
and UO_448 (O_448,N_2491,N_2737);
and UO_449 (O_449,N_2661,N_2751);
xnor UO_450 (O_450,N_2743,N_2392);
or UO_451 (O_451,N_2635,N_2805);
nand UO_452 (O_452,N_2495,N_2528);
xor UO_453 (O_453,N_2946,N_2554);
xor UO_454 (O_454,N_2375,N_2545);
nand UO_455 (O_455,N_2581,N_2609);
xor UO_456 (O_456,N_2380,N_2963);
and UO_457 (O_457,N_2904,N_2459);
nand UO_458 (O_458,N_2973,N_2444);
nor UO_459 (O_459,N_2989,N_2811);
and UO_460 (O_460,N_2716,N_2686);
and UO_461 (O_461,N_2348,N_2272);
nor UO_462 (O_462,N_2992,N_2373);
nor UO_463 (O_463,N_2583,N_2329);
or UO_464 (O_464,N_2761,N_2260);
or UO_465 (O_465,N_2969,N_2995);
nor UO_466 (O_466,N_2877,N_2337);
nand UO_467 (O_467,N_2421,N_2743);
and UO_468 (O_468,N_2382,N_2318);
nand UO_469 (O_469,N_2618,N_2877);
xnor UO_470 (O_470,N_2878,N_2391);
xnor UO_471 (O_471,N_2923,N_2765);
or UO_472 (O_472,N_2355,N_2949);
nand UO_473 (O_473,N_2561,N_2866);
and UO_474 (O_474,N_2607,N_2508);
xor UO_475 (O_475,N_2333,N_2693);
or UO_476 (O_476,N_2298,N_2971);
or UO_477 (O_477,N_2323,N_2913);
and UO_478 (O_478,N_2449,N_2531);
nand UO_479 (O_479,N_2925,N_2556);
or UO_480 (O_480,N_2277,N_2578);
nor UO_481 (O_481,N_2908,N_2934);
nand UO_482 (O_482,N_2445,N_2358);
nor UO_483 (O_483,N_2892,N_2374);
nand UO_484 (O_484,N_2317,N_2852);
nor UO_485 (O_485,N_2868,N_2979);
or UO_486 (O_486,N_2870,N_2317);
or UO_487 (O_487,N_2857,N_2985);
and UO_488 (O_488,N_2905,N_2488);
nor UO_489 (O_489,N_2783,N_2791);
and UO_490 (O_490,N_2984,N_2335);
xor UO_491 (O_491,N_2369,N_2637);
and UO_492 (O_492,N_2984,N_2352);
nand UO_493 (O_493,N_2419,N_2938);
or UO_494 (O_494,N_2762,N_2963);
and UO_495 (O_495,N_2601,N_2978);
nand UO_496 (O_496,N_2688,N_2739);
or UO_497 (O_497,N_2393,N_2419);
nor UO_498 (O_498,N_2711,N_2386);
nor UO_499 (O_499,N_2904,N_2607);
endmodule